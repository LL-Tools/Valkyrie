
module b17_C_2inp_gates_syn ( 
    P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
    DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
    DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
    DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
    DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
    DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
    P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
    P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
    P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
    P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
    P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
    P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
    P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
    P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
    P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
    P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
    P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
    P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
    P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
    P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
    P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
    P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
    P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
    P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN,
    P1_REIP_REG_6__SCAN_IN, P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
    P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN,
    P1_REIP_REG_0__SCAN_IN, P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
    P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN,
    P1_EBX_REG_26__SCAN_IN, P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
    P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN,
    P1_EBX_REG_20__SCAN_IN, P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
    P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN,
    P1_EBX_REG_14__SCAN_IN, P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
    P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
    P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
    P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
    P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
    P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN,
    P1_EAX_REG_28__SCAN_IN, P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
    P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN,
    P1_EAX_REG_22__SCAN_IN, P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
    P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN,
    P1_EAX_REG_16__SCAN_IN, P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
    P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN,
    P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN,
    P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN,
    P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN,
    P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN,
    P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
    P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
    P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
    P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
    P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
    P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
    P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
    P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
    P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
    P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
    P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
    P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
    P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
    P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
    P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
    P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN,
    P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN,
    P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN,
    P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN,
    P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN,
    P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN,
    P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN,
    P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN,
    P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN,
    P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN,
    P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN,
    P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN,
    P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN,
    P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN,
    P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN,
    P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN,
    P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN,
    P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN,
    P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN,
    P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN,
    P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN,
    P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN,
    P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN,
    P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN,
    P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN,
    P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN,
    P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN,
    P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN,
    P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN,
    P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN,
    P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN,
    P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN,
    P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN,
    P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN,
    P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN,
    P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN,
    P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN,
    P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN,
    P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN,
    P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN,
    P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN,
    P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN,
    P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN,
    P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN,
    P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN,
    P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN,
    P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN,
    P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN,
    P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
    P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
    P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
    P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
    P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
    P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN,
    P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN,
    P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN,
    P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN,
    P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN,
    P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN,
    P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN,
    P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN,
    P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN,
    P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN,
    P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN,
    P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN,
    P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN,
    P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN,
    P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN,
    P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN,
    P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN,
    BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN,
    BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN,
    BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN,
    BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN,
    BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN,
    BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN,
    BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN,
    BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN,
    BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN,
    BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN,
    BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN,
    BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN,
    BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN,
    BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN,
    BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN,
    BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN,
    BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN,
    BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN,
    BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN,
    BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN,
    BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN,
    READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN,
    READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN,
    P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN,
    P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN,
    P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN,
    P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN,
    P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN,
    P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN,
    P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN,
    P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN,
    P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN,
    P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN,
    P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN,
    P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN,
    P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN,
    P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN,
    P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN,
    P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN,
    P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN,
    P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN,
    P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN,
    P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN,
    P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN,
    P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN,
    P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN,
    P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN,
    P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN,
    P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN,
    P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN,
    P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN,
    P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN,
    P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN,
    P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN,
    P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN,
    P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN,
    P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN,
    P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN,
    P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN,
    P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN,
    P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN,
    P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN,
    P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN,
    P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN,
    P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN,
    P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN,
    P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN,
    P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN,
    P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN,
    P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN,
    P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN,
    P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN,
    P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN,
    P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN,
    P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN,
    P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN,
    P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN,
    P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN,
    P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN,
    P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN,
    P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN,
    P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN,
    P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN,
    P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN,
    P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN,
    P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN,
    P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN,
    P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN,
    P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN,
    P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN,
    P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN,
    P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN,
    P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN,
    P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN,
    P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN,
    P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN,
    P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN,
    P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN,
    P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN,
    P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN,
    P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN,
    P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN,
    P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN,
    P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN,
    P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN,
    P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN,
    P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN,
    P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN,
    P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN,
    P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN,
    P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN,
    P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN,
    P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN,
    P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN,
    P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN,
    P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN,
    P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN,
    P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN,
    P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN,
    P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN,
    P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN,
    P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN,
    P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
    P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
    P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
    P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
    P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
    P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
    P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
    P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
    P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
    P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
    P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
    P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN,
    P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN,
    P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN,
    P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN,
    P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN,
    P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN,
    P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN,
    P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN,
    P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN,
    P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN,
    P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
    P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
    P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
    P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
    P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
    P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
    P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
    P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
    P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
    P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
    P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
    P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
    P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
    P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
    P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
    P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
    P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
    P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
    P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
    P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
    P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
    P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
    P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
    P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
    P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
    P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
    P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
    P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
    P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
    P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
    P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
    P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
    P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
    P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
    P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
    P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
    P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
    P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
    P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
    P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
    P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
    P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
    P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
    P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
    P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
    P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
    P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
    P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
    P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
    P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
    P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
    P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
    P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN,
    P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
    P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN,
    P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
    P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN,
    P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
    P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
    P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
    P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
    P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
    P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN,
    P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
    P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN,
    P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
    P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN,
    P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
    P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN,
    P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
    P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN,
    P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
    P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
    P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
    P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
    P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
    P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
    P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
    P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
    P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
    P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
    P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
    P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
    P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
    P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
    P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
    P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
    P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
    P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
    P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
    P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
    P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN,
    P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN,
    P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN,
    P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN,
    P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN,
    P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN,
    P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN,
    P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN,
    P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN,
    P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN,
    P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN,
    P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN,
    P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN,
    P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN,
    P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN,
    P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN,
    P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN,
    P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN,
    P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN,
    P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN,
    P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN,
    P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN,
    P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN,
    P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN,
    P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN,
    P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN,
    P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN,
    P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN,
    P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN,
    P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN,
    P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN,
    P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN,
    P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN,
    P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN,
    P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN,
    P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN,
    P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN,
    P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN,
    P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN,
    P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN,
    P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN,
    P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN,
    P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN,
    P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN,
    P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN,
    P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN,
    P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN,
    P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN,
    P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN,
    P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN,
    P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN,
    P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN,
    P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN,
    P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN,
    P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN,
    P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN,
    P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN,
    P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN,
    P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN,
    P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN,
    P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN,
    P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN,
    P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN,
    P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN,
    P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN,
    P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN,
    P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN,
    P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN,
    P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN,
    P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN,
    P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN,
    P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN,
    P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN,
    P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN,
    P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN,
    P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN,
    P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN,
    P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN,
    P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN,
    P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN,
    P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN,
    P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN,
    P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN,
    P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN,
    P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN,
    P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN,
    P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN,
    P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN,
    P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN,
    P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN,
    P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN,
    P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN,
    P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN,
    P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN,
    P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN,
    P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN,
    P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN,
    P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN,
    P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN,
    P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
    P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
    P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
    P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
    P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
    P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
    P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
    P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
    P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
    P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
    P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
    P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN,
    P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN,
    P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN,
    P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN,
    P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN,
    P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN,
    P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN,
    P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN,
    P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN,
    P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN,
    P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
    P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
    P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
    P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
    P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
    P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
    P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
    P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
    P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
    P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
    P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
    P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
    P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
    P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
    P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
    P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
    P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
    P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
    P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
    P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
    P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
    P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
    P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
    P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
    P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
    P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
    P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
    P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
    P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
    P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
    P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
    P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
    P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
    P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
    P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
    P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
    P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
    P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
    P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
    P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
    P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
    P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
    P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
    P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
    P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
    P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
    P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
    P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
    P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
    P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
    P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
    P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
    P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN,
    P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
    P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN,
    P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
    P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN,
    P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
    P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
    P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
    P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
    P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
    P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN,
    P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
    P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN,
    P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
    P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN,
    P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
    P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN,
    P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
    P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN,
    P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
    P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
    P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
    P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
    P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
    P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
    P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
    P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
    P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
    P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
    P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
    P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
    P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
    P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
    P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
    P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
    P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
    P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
    P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
    P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
    P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN,
    P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN,
    P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN,
    P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN,
    P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN,
    P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN,
    P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN,
    P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN,
    P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN,
    P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN,
    P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN,
    P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN,
    P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN,
    P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN,
    P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN,
    P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN,
    P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN,
    P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN,
    P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN,
    P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN,
    P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN,
    P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN,
    P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN,
    P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN,
    P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN,
    P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN,
    P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN,
    P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN,
    P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN,
    P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN,
    P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN,
    P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN,
    P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN,
    P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN,
    P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN,
    P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN,
    P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN,
    P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN,
    P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN,
    P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN,
    P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN,
    P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN,
    P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN,
    P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN,
    P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN,
    P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN,
    P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN,
    P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN,
    P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN,
    P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN,
    P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN,
    P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN,
    P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN,
    P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN,
    P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN,
    P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN,
    P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN,
    P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN,
    P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN,
    P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN,
    P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN,
    P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN,
    P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN,
    P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN,
    P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN,
    P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN,
    P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN,
    P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN,
    P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN,
    P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN,
    P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN,
    P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN,
    P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN,
    P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN,
    P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN,
    P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN,
    P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN,
    P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN,
    P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN,
    P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN,
    P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN,
    P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN,
    P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN,
    U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366, U367,
    U368, U369, U370, U371, U372, U373, U374, U375, U347, U348, U349, U350,
    U351, U352, U353, U354, U365, U376, U247, U246, U245, U244, U243, U242,
    U241, U240, U239, U238, U237, U236, U235, U234, U233, U232, U231, U230,
    U229, U228, U227, U226, U225, U224, U223, U222, U221, U220, U219, U218,
    U217, U216, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260,
    U261, U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272,
    U273, U274, U275, U276, U277, U278, U279, U280, U281, U282, U212, U215,
    U213, U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060,
    P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053,
    P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046,
    P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039,
    P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032,
    P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027,
    P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020,
    P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013,
    P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006,
    P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999,
    P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993,
    P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986,
    P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979,
    P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972,
    P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965,
    P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958,
    P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951,
    P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944,
    P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937,
    P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930,
    P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923,
    P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916,
    P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909,
    P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902,
    P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895,
    P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888,
    P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881,
    P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874,
    P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284,
    P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865,
    P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858,
    P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851,
    P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844,
    P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837,
    P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830,
    P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823,
    P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816,
    P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809,
    P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802,
    P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795,
    P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788,
    P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781,
    P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774,
    P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767,
    P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760,
    P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753,
    P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746,
    P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739,
    P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732,
    P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725,
    P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718,
    P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711,
    P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704,
    P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697,
    P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690,
    P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683,
    P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676,
    P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669,
    P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662,
    P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655,
    P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648,
    P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641,
    P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637,
    P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633,
    P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241,
    P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
    P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
    P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
    P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213,
    P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208,
    P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201,
    P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194,
    P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187,
    P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180,
    P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174,
    P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167,
    P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160,
    P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153,
    P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146,
    P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139,
    P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132,
    P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125,
    P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118,
    P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111,
    P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104,
    P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097,
    P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090,
    P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083,
    P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076,
    P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069,
    P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062,
    P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055,
    P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048,
    P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602,
    P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043,
    P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036,
    P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029,
    P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022,
    P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015,
    P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008,
    P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001,
    P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994,
    P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987,
    P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980,
    P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973,
    P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966,
    P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959,
    P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952,
    P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945,
    P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938,
    P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931,
    P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924,
    P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917,
    P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910,
    P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903,
    P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896,
    P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889,
    P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882,
    P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875,
    P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868,
    P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861,
    P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854,
    P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847,
    P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840,
    P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833,
    P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826,
    P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608,
    P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816,
    P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461,
    P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220,
    P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213,
    P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206,
    P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199,
    P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465,
    P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187,
    P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180,
    P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173,
    P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166,
    P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160,
    P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153,
    P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146,
    P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139,
    P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132,
    P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125,
    P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118,
    P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111,
    P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104,
    P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097,
    P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090,
    P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083,
    P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076,
    P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069,
    P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062,
    P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055,
    P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048,
    P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041,
    P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034,
    P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032,
    P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029,
    P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022,
    P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015,
    P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008,
    P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001,
    P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994,
    P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987,
    P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980,
    P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973,
    P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966,
    P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959,
    P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952,
    P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945,
    P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938,
    P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931,
    P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924,
    P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917,
    P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910,
    P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903,
    P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896,
    P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889,
    P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882,
    P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875,
    P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868,
    P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861,
    P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854,
    P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847,
    P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840,
    P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833,
    P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826,
    P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819,
    P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812,
    P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482,
    P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486,
    P1_U2803, P1_U2802, P1_U3487, P1_U2801  );
  input  P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_,
    DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_,
    DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_,
    DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_,
    DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_,
    DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
    P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
    P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
    P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
    P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
    P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
    P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
    P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
    P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
    P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
    P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
    P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
    P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
    P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
    P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
    P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
    P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
    P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
    P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN,
    P1_REIP_REG_6__SCAN_IN, P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
    P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN,
    P1_REIP_REG_0__SCAN_IN, P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
    P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN,
    P1_EBX_REG_26__SCAN_IN, P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
    P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN,
    P1_EBX_REG_20__SCAN_IN, P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
    P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN,
    P1_EBX_REG_14__SCAN_IN, P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
    P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
    P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
    P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
    P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
    P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN,
    P1_EAX_REG_28__SCAN_IN, P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
    P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN,
    P1_EAX_REG_22__SCAN_IN, P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
    P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN,
    P1_EAX_REG_16__SCAN_IN, P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
    P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN,
    P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN,
    P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN,
    P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN,
    P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN,
    P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
    P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
    P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
    P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
    P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
    P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
    P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
    P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
    P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
    P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
    P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
    P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
    P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
    P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
    P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
    P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN,
    P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN,
    P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN,
    P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN,
    P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN,
    P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN,
    P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN,
    P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN,
    P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN,
    P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN,
    P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN,
    P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN,
    P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN,
    P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN,
    P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN,
    P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN,
    P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN,
    P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN,
    P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN,
    P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN,
    P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN,
    P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN,
    P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN,
    P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN,
    P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN,
    P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN,
    P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN,
    P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN,
    P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN,
    P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN,
    P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN,
    P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN,
    P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN,
    P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN,
    P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN,
    P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN,
    P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN,
    P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN,
    P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN,
    P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN,
    P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN,
    P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN,
    P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN,
    P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN,
    P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN,
    P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN,
    P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN,
    P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN,
    P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
    P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
    P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
    P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
    P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
    P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN,
    P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN,
    P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN,
    P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN,
    P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN,
    P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN,
    P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN,
    P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN,
    P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN,
    P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN,
    P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN,
    P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN,
    P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN,
    P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN,
    P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN,
    P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN,
    P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN,
    BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN,
    BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN,
    BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN,
    BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN,
    BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN,
    BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN,
    BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN,
    BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN,
    BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN,
    BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN,
    BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN,
    BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN,
    BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN,
    BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN,
    BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN,
    BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN,
    BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN,
    BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN,
    BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN,
    BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN,
    BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN,
    READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN,
    READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN,
    P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN,
    P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN,
    P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN,
    P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN,
    P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN,
    P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN,
    P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN,
    P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN,
    P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN,
    P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN,
    P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN,
    P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN,
    P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN,
    P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN,
    P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN,
    P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN,
    P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN,
    P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN,
    P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN,
    P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN,
    P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN,
    P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN,
    P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN,
    P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN,
    P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN,
    P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN,
    P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN,
    P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN,
    P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN,
    P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN,
    P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN,
    P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN,
    P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN,
    P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN,
    P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN,
    P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN,
    P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN,
    P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN,
    P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN,
    P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN,
    P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN,
    P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN,
    P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN,
    P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN,
    P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN,
    P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN,
    P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN,
    P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN,
    P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN,
    P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN,
    P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN,
    P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN,
    P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN,
    P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN,
    P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN,
    P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN,
    P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN,
    P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN,
    P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN,
    P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN,
    P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN,
    P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN,
    P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN,
    P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN,
    P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN,
    P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN,
    P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN,
    P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN,
    P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN,
    P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN,
    P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN,
    P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN,
    P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN,
    P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN,
    P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN,
    P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN,
    P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN,
    P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN,
    P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN,
    P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN,
    P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN,
    P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN,
    P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN,
    P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN,
    P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN,
    P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN,
    P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN,
    P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN,
    P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN,
    P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN,
    P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN,
    P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN,
    P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN,
    P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN,
    P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN,
    P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN,
    P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN,
    P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN,
    P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN,
    P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
    P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
    P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
    P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
    P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
    P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
    P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
    P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
    P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
    P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
    P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
    P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN,
    P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN,
    P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN,
    P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN,
    P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN,
    P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN,
    P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN,
    P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN,
    P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN,
    P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN,
    P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
    P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
    P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
    P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
    P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
    P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
    P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
    P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
    P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
    P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
    P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
    P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
    P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
    P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
    P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
    P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
    P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
    P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
    P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
    P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
    P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
    P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
    P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
    P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
    P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
    P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
    P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
    P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
    P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
    P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
    P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
    P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
    P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
    P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
    P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
    P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
    P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
    P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
    P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
    P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
    P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
    P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
    P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
    P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
    P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
    P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
    P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
    P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
    P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
    P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
    P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
    P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
    P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN,
    P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
    P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN,
    P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
    P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN,
    P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
    P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
    P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
    P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
    P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
    P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN,
    P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
    P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN,
    P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
    P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN,
    P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
    P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN,
    P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
    P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN,
    P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
    P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
    P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
    P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
    P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
    P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
    P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
    P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
    P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
    P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
    P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
    P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
    P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
    P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
    P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
    P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
    P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
    P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
    P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
    P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
    P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN,
    P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN,
    P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN,
    P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN,
    P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN,
    P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN,
    P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN,
    P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN,
    P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN,
    P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN,
    P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN,
    P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN,
    P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN,
    P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN,
    P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN,
    P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN,
    P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN,
    P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN,
    P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN,
    P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN,
    P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN,
    P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN,
    P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN,
    P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN,
    P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN,
    P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN,
    P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN,
    P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN,
    P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN,
    P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN,
    P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN,
    P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN,
    P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN,
    P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN,
    P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN,
    P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN,
    P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN,
    P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN,
    P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN,
    P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN,
    P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN,
    P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN,
    P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN,
    P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN,
    P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN,
    P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN,
    P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN,
    P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN,
    P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN,
    P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN,
    P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN,
    P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN,
    P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN,
    P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN,
    P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN,
    P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN,
    P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN,
    P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN,
    P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN,
    P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN,
    P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN,
    P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN,
    P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN,
    P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN,
    P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN,
    P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN,
    P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN,
    P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN,
    P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN,
    P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN,
    P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN,
    P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN,
    P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN,
    P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN,
    P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN,
    P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN,
    P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN,
    P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN,
    P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN,
    P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN,
    P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN,
    P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN,
    P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN,
    P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN,
    P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN,
    P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN,
    P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN,
    P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN,
    P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN,
    P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN,
    P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN,
    P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN,
    P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN,
    P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN,
    P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN,
    P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN,
    P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN,
    P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN,
    P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN,
    P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
    P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
    P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
    P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
    P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
    P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
    P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
    P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
    P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
    P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
    P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
    P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN,
    P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN,
    P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN,
    P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN,
    P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN,
    P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN,
    P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN,
    P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN,
    P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN,
    P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN,
    P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
    P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
    P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
    P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
    P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
    P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
    P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
    P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
    P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
    P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
    P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
    P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
    P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
    P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
    P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
    P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
    P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
    P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
    P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
    P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
    P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
    P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
    P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
    P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
    P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
    P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
    P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
    P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
    P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
    P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
    P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
    P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
    P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
    P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
    P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
    P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
    P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
    P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
    P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
    P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
    P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
    P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
    P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
    P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
    P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
    P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
    P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
    P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
    P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
    P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
    P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
    P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
    P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN,
    P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
    P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN,
    P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
    P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN,
    P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
    P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
    P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
    P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
    P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
    P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN,
    P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
    P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN,
    P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
    P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN,
    P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
    P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN,
    P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
    P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN,
    P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
    P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
    P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
    P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
    P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
    P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
    P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
    P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
    P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
    P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
    P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
    P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
    P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
    P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
    P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
    P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
    P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
    P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
    P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
    P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
    P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN,
    P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN,
    P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN,
    P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN,
    P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN,
    P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN,
    P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN,
    P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN,
    P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN,
    P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN,
    P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN,
    P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN,
    P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN,
    P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN,
    P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN,
    P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN,
    P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN,
    P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN,
    P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN,
    P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN,
    P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN,
    P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN,
    P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN,
    P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN,
    P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN,
    P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN,
    P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN,
    P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN,
    P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN,
    P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN,
    P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN,
    P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN,
    P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN,
    P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN,
    P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN,
    P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN,
    P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN,
    P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN,
    P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN,
    P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN,
    P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN,
    P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN,
    P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN,
    P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN,
    P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN,
    P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN,
    P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN,
    P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN,
    P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN,
    P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN,
    P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN,
    P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN,
    P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN,
    P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN,
    P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN,
    P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN,
    P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN,
    P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN,
    P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN,
    P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN,
    P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN,
    P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN,
    P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN,
    P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN,
    P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN,
    P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN,
    P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN,
    P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN,
    P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN,
    P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN,
    P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN,
    P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN,
    P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN,
    P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN,
    P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN,
    P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN,
    P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN,
    P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN,
    P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN,
    P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN,
    P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN,
    P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN,
    P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
    U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348, U349,
    U350, U351, U352, U353, U354, U365, U376, U247, U246, U245, U244, U243,
    U242, U241, U240, U239, U238, U237, U236, U235, U234, U233, U232, U231,
    U230, U229, U228, U227, U226, U225, U224, U223, U222, U221, U220, U219,
    U218, U217, U216, U251, U252, U253, U254, U255, U256, U257, U258, U259,
    U260, U261, U262, U263, U264, U265, U266, U267, U268, U269, U270, U271,
    U272, U273, U274, U275, U276, U277, U278, U279, U280, U281, U282, U212,
    U215, U213, U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061,
    P3_U3060, P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054,
    P3_U3053, P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047,
    P3_U3046, P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040,
    P3_U3039, P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033,
    P3_U3032, P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028,
    P3_U3027, P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021,
    P3_U3020, P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014,
    P3_U3013, P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007,
    P3_U3006, P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000,
    P3_U2999, P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994,
    P3_U2993, P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987,
    P3_U2986, P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980,
    P3_U2979, P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973,
    P3_U2972, P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966,
    P3_U2965, P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959,
    P3_U2958, P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952,
    P3_U2951, P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945,
    P3_U2944, P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938,
    P3_U2937, P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931,
    P3_U2930, P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924,
    P3_U2923, P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917,
    P3_U2916, P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910,
    P3_U2909, P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903,
    P3_U2902, P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896,
    P3_U2895, P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889,
    P3_U2888, P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882,
    P3_U2881, P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875,
    P3_U2874, P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868,
    P3_U3284, P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866,
    P3_U2865, P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859,
    P3_U2858, P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852,
    P3_U2851, P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845,
    P3_U2844, P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838,
    P3_U2837, P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831,
    P3_U2830, P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824,
    P3_U2823, P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817,
    P3_U2816, P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810,
    P3_U2809, P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803,
    P3_U2802, P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796,
    P3_U2795, P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789,
    P3_U2788, P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782,
    P3_U2781, P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775,
    P3_U2774, P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768,
    P3_U2767, P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761,
    P3_U2760, P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754,
    P3_U2753, P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747,
    P3_U2746, P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740,
    P3_U2739, P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733,
    P3_U2732, P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726,
    P3_U2725, P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719,
    P3_U2718, P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712,
    P3_U2711, P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705,
    P3_U2704, P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698,
    P3_U2697, P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691,
    P3_U2690, P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684,
    P3_U2683, P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677,
    P3_U2676, P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670,
    P3_U2669, P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663,
    P3_U2662, P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656,
    P3_U2655, P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649,
    P3_U2648, P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642,
    P3_U2641, P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294,
    P3_U2637, P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634,
    P3_U2633, P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588,
    P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
    P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
    P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
    P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214,
    P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592,
    P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202,
    P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195,
    P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188,
    P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181,
    P2_U3180, P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175,
    P2_U3174, P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168,
    P2_U3167, P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161,
    P2_U3160, P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154,
    P2_U3153, P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147,
    P2_U3146, P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140,
    P2_U3139, P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133,
    P2_U3132, P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126,
    P2_U3125, P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119,
    P2_U3118, P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112,
    P2_U3111, P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105,
    P2_U3104, P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098,
    P2_U3097, P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091,
    P2_U3090, P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084,
    P2_U3083, P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077,
    P2_U3076, P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070,
    P2_U3069, P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063,
    P2_U3062, P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056,
    P2_U3055, P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049,
    P2_U3048, P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047,
    P2_U3602, P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044,
    P2_U3043, P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037,
    P2_U3036, P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030,
    P2_U3029, P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023,
    P2_U3022, P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016,
    P2_U3015, P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009,
    P2_U3008, P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002,
    P2_U3001, P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995,
    P2_U2994, P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988,
    P2_U2987, P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981,
    P2_U2980, P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974,
    P2_U2973, P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967,
    P2_U2966, P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960,
    P2_U2959, P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953,
    P2_U2952, P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946,
    P2_U2945, P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939,
    P2_U2938, P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932,
    P2_U2931, P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925,
    P2_U2924, P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918,
    P2_U2917, P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911,
    P2_U2910, P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904,
    P2_U2903, P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897,
    P2_U2896, P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890,
    P2_U2889, P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883,
    P2_U2882, P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876,
    P2_U2875, P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869,
    P2_U2868, P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862,
    P2_U2861, P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855,
    P2_U2854, P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848,
    P2_U2847, P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841,
    P2_U2840, P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834,
    P2_U2833, P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827,
    P2_U2826, P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820,
    P2_U3608, P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611,
    P2_U2816, P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460,
    P1_U3461, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221,
    P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214,
    P1_U3213, P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207,
    P1_U3206, P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200,
    P1_U3199, P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464,
    P1_U3465, P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188,
    P1_U3187, P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181,
    P1_U3180, P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174,
    P1_U3173, P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167,
    P1_U3166, P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161,
    P1_U3160, P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154,
    P1_U3153, P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147,
    P1_U3146, P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140,
    P1_U3139, P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133,
    P1_U3132, P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126,
    P1_U3125, P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119,
    P1_U3118, P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112,
    P1_U3111, P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105,
    P1_U3104, P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098,
    P1_U3097, P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091,
    P1_U3090, P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084,
    P1_U3083, P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077,
    P1_U3076, P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070,
    P1_U3069, P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063,
    P1_U3062, P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056,
    P1_U3055, P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049,
    P1_U3048, P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042,
    P1_U3041, P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035,
    P1_U3034, P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474,
    P1_U3032, P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030,
    P1_U3029, P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023,
    P1_U3022, P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016,
    P1_U3015, P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009,
    P1_U3008, P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002,
    P1_U3001, P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995,
    P1_U2994, P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988,
    P1_U2987, P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981,
    P1_U2980, P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974,
    P1_U2973, P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967,
    P1_U2966, P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960,
    P1_U2959, P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953,
    P1_U2952, P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946,
    P1_U2945, P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939,
    P1_U2938, P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932,
    P1_U2931, P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925,
    P1_U2924, P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918,
    P1_U2917, P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911,
    P1_U2910, P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904,
    P1_U2903, P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897,
    P1_U2896, P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890,
    P1_U2889, P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883,
    P1_U2882, P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876,
    P1_U2875, P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869,
    P1_U2868, P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862,
    P1_U2861, P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855,
    P1_U2854, P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848,
    P1_U2847, P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841,
    P1_U2840, P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834,
    P1_U2833, P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827,
    P1_U2826, P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820,
    P1_U2819, P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813,
    P1_U2812, P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807,
    P1_U3482, P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804,
    P1_U3486, P1_U2803, P1_U2802, P1_U3487, P1_U2801;
  wire n43871, n36151, n41228, n41686, n43067, n43398, n40820, n41751,
    n25837, n23180, n32932, n38758, n41418, n23864, n29891, n24634, n37494,
    n37473, n37482, n28494, n27817, n42760, n26866, n29581, n22838, n35412,
    n28734, n29753, n43161, n39805, n24802, n26630, n24898, n24936, n24734,
    n29002, n40303, n22818, n22819, n22820, n22822, n22823, n22825, n28500,
    n25085, n38721, n26859, n27880, n28283, n23627, n27665, n24721, n24668,
    n24116, n24010, n28596, n28669, n28586, n24598, n38695, n24188, n38757,
    n30957, n28980, n39627, n41785, n24522, n22828, n35252, n42461, n44298,
    n31658, n23244, n23178, n23222, n40560, n27656, n34384, n34430, n24625,
    n22837, n40729, n41878, n34470, n34971, n36662, n37453, n39110, n43042,
    n39820, n42177, n32726, n34631, n22826, n22827, n26986, n23702, n27631,
    n30654, n30851, n26482, n28126, n27908, n30676, n22964, n31700, n23126,
    n27900, n31974, n23515, n27610, n37190, n27163, n27162, n42961, n23690,
    n25235, n22829, n28298, n24763, n24738, n28309, n22830, n36515, n25555,
    n34525, n22832, n22833, n26806, n36767, n34447, n33747, n37008, n22834,
    n38696, n27742, n23181, n23438, n23269, n32526, n23493, n23331, n43892,
    n22835, n30950, n25883, n23091, n27884, n27781, n42932, n25411, n25393,
    n28174, n27715, n25030, n29831, n37514, n25054, n23706, n25009, n24927,
    n22836, n40437, n22841, n24315, n27510, n29761, n24815, n25089, n27348,
    n29861, n23335, n23662, n32829, n23179, n23295, n32321, n23465, n32613,
    n32750, n23462, n32197, n23522, n32212, n32898, n32200, n30663, n32186,
    n32433, n29029, n30889, n23443, n30657, n23422, n31971, n23520, n30687,
    n26908, n23195, n38806, n30791, n30665, n23847, n23115, n29991, n44042,
    n43366, n32524, n32634, n23425, n23695, n41399, n23338, n29842, n38790,
    n23407, n28305, n23340, n23326, n41329, n28300, n28070, n31810, n36191,
    n23588, n22905, n35514, n30899, n29810, n42391, n27844, n42413, n41310,
    n41479, n42960, n42446, n25916, n23664, n42400, n30826, n43102, n43117,
    n23484, n30878, n43132, n33204, n27877, n26954, n26956, n43147, n29813,
    n30883, n42631, n41411, n41788, n42625, n30908, n41242, n23321, n36832,
    n41490, n42443, n23397, n23090, n27887, n29805, n39335, n42937, n40657,
    n32254, n27780, n39620, n42153, n40577, n27956, n27767, n31689, n42076,
    n23743, n29326, n23446, n39636, n23669, n31954, n25859, n44767, n25868,
    n22848, n31955, n23926, n28145, n27723, n23904, n28154, n39588, n24582,
    n23350, n27732, n23349, n23867, n34002, n34376, n26568, n23359, n38797,
    n27729, n26526, n23675, n27695, n27688, n29843, n25833, n23725, n25048,
    n23930, n23724, n27549, n24617, n23903, n23117, n34116, n28242, n23727,
    n23728, n36610, n27677, n39443, n25822, n25629, n25660, n23234, n28575,
    n28512, n27579, n22839, n25645, n25669, n25001, n28601, n24187, n26914,
    n25601, n31502, n25462, n25639, n23537, n33802, n25055, n25042, n43131,
    n28498, n24865, n28595, n25008, n35773, n25661, n43057, n25011, n39593,
    n42209, n43116, n43146, n28552, n43101, n35753, n25017, n25609, n40501,
    n33538, n27531, n24569, n24149, n40471, n40444, n24897, n22840, n27208,
    n24801, n24928, n23227, n27209, n24925, n24783, n24893, n24924, n24851,
    n29575, n29580, n33147, n41894, n27045, n22842, n24923, n24513, n24300,
    n24292, n27319, n24972, n24973, n24989, n25065, n25118, n27379, n27334,
    n42024, n41158, n27218, n27228, n36653, n29752, n44597, n44691, n22843,
    n23065, n24005, n24006, n22844, n24318, n44835, n23758, n31657, n38728,
    n23999, n25912, n25196, n31445, n31449, n24753, n31651, n25614, n42196,
    n38719, n42134, n34451, n38709, n34395, n24000, n22845, n22846, n33342,
    n22847, n27886, n23692, n41782, n27412, n30257, n22849, n23630, n27779,
    n24253, n23128, n23189, n29739, n23932, n36297, n26899, n23569, n31670,
    n31668, n31662, n27121, n27245, n27195, n27149, n27184, n27213, n27136,
    n22850, n23101, n22851, n22852, n22853, n22854, n22855, n23505, n29588,
    n27747, n31012, n39380, n22856, n22857, n22858, n42120, n23194, n22859,
    n23271, n23696, n24861, n31431, n22860, n39637, n23174, n32305, n22862,
    n27509, n30684, n31663, n43065, n23299, n23280, n43379, n22863, n22864,
    n33146, n31665, n31667, n31669, n31659, n31660, n31661, n23275, n25232,
    n25648, n25642, n25243, n23916, n23341, n23343, n29320, n23445, n28347,
    n23482, n23819, n23722, n23860, n28835, n23388, n29319, n23684, n23685,
    n23774, n23772, n23840, n23816, n31420, n43051, n23506, n23141, n25778,
    n43056, n32931, n28344, n23262, n23945, n23481, n23478, n23896, n23897,
    n34483, n34320, n36384, n23147, n25677, n25675, n29896, n23253, n23254,
    n31896, n32441, n32537, n23245, n23246, n29013, n23450, n25616, n23594,
    n24765, n23183, n23777, n23781, n23778, n23779, n23780, n25107, n24813,
    n24814, n23580, n25426, n25414, n23834, n23906, n23907, n23374, n23395,
    n28142, n23912, n23920, n23918, n27498, n29497, n23231, n23232, n38775,
    n23392, n23470, n23186, n25646, n25457, n23491, n25424, n23507, n25189,
    n25550, n24961, n24896, n25004, n23233, n23230, n28553, n23877, n23910,
    n23911, n23576, n28090, n23477, n23719, n23854, n23720, n23855, n23342,
    n32527, n28012, n28295, n27693, n27672, n23686, n27336, n27221, n34779,
    n24009, n38740, n23759, n24633, n31508, n25647, n25594, n25595, n25789,
    n23808, n23809, n25730, n42444, n25043, n23285, n26890, n23843, n23845,
    n23844, n23839, n23841, n23812, n29993, n23739, n23741, n30825, n23559,
    n23558, n23560, n23184, n23729, n30228, n23208, n23209, n30269, n25498,
    n31368, n23673, n23328, n23776, n25709, n43380, n23620, n43082, n25392,
    n44308, n31524, n23461, n23460, n28879, n23882, n23517, n23828, n23518,
    n23832, n23833, n29633, n23880, n23881, n32837, n33239, n23873, n23874,
    n27632, n23884, n29780, n31832, n23944, n23432, n23433, n23435, n23753,
    n23898, n29025, n23700, n23579, n39356, n23666, n32470, n28071, n31958,
    n42140, n27775, n40436, n23708, n27566, n33228, n27561, n27562, n23367,
    n24704, n23547, n33801, n23796, n23797, n24585, n23653, n23196, n33307,
    n33408, n23202, n38673, n24593, n24604, n31417, n23848, n30013, n30056,
    n23214, n23215, n23810, n30332, n31370, n23632, n23838, n23320, n42963,
    n27060, n31541, n43967, n44399, n44152, n43471, n43199, n44418, n31570,
    n31573, n23458, n23456, n39141, n33245, n29799, n31595, n23252, n32168,
    n28967, n32405, n23902, n32457, n23886, n23888, n23889, n23887, n23890,
    n23891, n32564, n23892, n23264, n23413, n23418, n23710, n40111, n39975,
    n23665, n23637, n23749, n23747, n23748, n32309, n29070, n32359, n23267,
    n23694, n40399, n27883, n41575, n40557, n41002, n41664, n33788, n24632,
    n35812, n33905, n34371, n23366, n24021, n35504, n33428, n23760, n23761,
    n33284, n23535, n37197, n39105, n38815, n43062, n23182, n23613, n23611,
    n23315, n31091, n23607, n23608, n39888, n31969, n40397, n23502, n23503,
    n40408, n39132, n35945, n35667, n35671, n23659, n23660, n23200, n23452,
    n25615, n23311, n27916, n23595, n27893, n23600, n27898, n27981, n27853,
    n26360, n26320, n24754, n25619, n24882, n29188, n29171, n27410, n27849,
    n27777, n27759, n29536, n23276, n27447, n24969, n26753, n23508, n23509,
    n23735, n25692, n23602, n24878, n23098, n29696, n29124, n23681, n29226,
    n29687, n29574, n29426, n23226, n27810, n23345, n23721, n23857, n23565,
    n23566, n23567, n23573, n23905, n23385, n23410, n23386, n23411, n23406,
    n28033, n23236, n23396, n23369, n29576, n29669, n27125, n27183, n27446,
    n27350, n27359, n24608, n23368, n34396, n25592, n25593, n24735, n24762,
    n26522, n25499, n23322, n25685, n23302, n23211, n23212, n25464, n23329,
    n23626, n25455, n25443, n25139, n23557, n31446, n25134, n43548, n29801,
    n23924, n23925, n23915, n28127, n28080, n28073, n28064, n28094, n23373,
    n29577, n27700, n23711, n29749, n29709, n23263, n23400, n29331, n29330,
    n29311, n28152, n28150, n23923, n28160, n23381, n23940, n23699, n23869,
    n23868, n32602, n27795, n23919, n23378, n27501, n28577, n23571, n23716,
    n23707, n23693, n23691, n27552, n23551, n23548, n23534, n23995, n35811,
    n38724, n23356, n23216, n23217, n26184, n23625, n23469, n23678, n25022,
    n23849, n30440, n26910, n26975, n26842, n26794, n26745, n26656, n26399,
    n26318, n26267, n23628, n26072, n26031, n25990, n23287, n23811, n30140,
    n23210, n30845, n23733, n23806, n23807, n25507, n30633, n25679, n23308,
    n23309, n31415, n23802, n23800, n42462, n42464, n25398, n23835, n25234,
    n43081, n44051, n25182, n44132, n44765, n44775, n31555, n23459, n42244,
    n28246, n29803, n23922, n23875, n23876, n23908, n23909, n39291, n28714,
    n28118, n23382, n23383, n31646, n23830, n23831, n28572, n39973, n31831,
    n31666, n31664, n23853, n23479, n23476, n29829, n32653, n23878, n23879,
    n31901, n29087, n23486, n32904, n23817, n23617, n32536, n23426, n32525,
    n23634, n23635, n23933, n29800, n33136, n28291, n28290, n23256, n29314,
    n33162, n23570, n33165, n27773, n41324, n41503, n27536, n41489, n27613,
    n24710, n33322, n38694, n38687, n36107, n36113, n36164, n36196, n36231,
    n23549, n23550, n36267, n23794, n36483, n37091, n36540, n36536, n36590,
    n36622, n36766, n24283, n36278, n36321, n23647, n23773, n37239, n36704,
    n37338, n30058, n25804, n23804, n27102, n30174, n26273, n23846, n42411,
    n30327, n26973, n23814, n42421, n43190, n26660, n26661, n42582, n30602,
    n42621, n42752, n42761, n30645, n30767, n30792, n30855, n30891, n30283,
    n30971, n30982, n31023, n42895, n23824, n23822, n42945, n23323, n30652,
    n42947, n23931, n23624, n30980, n30992, n31400, n23928, n42929, n44760,
    n31528, n44744, n43281, n43225, n43449, n43397, n44766, n43951, n44306,
    n44138, n44294, n44230, n44382, n44394, n44468, n44491, n44415, n44750,
    n44853, n44850, n33223, n23883, n31699, n31736, n31789, n31806, n31813,
    n31929, n23250, n29086, n23862, n23865, n39672, n32391, n23901, n39709,
    n32585, n23150, n39814, n27637, n33137, n23258, n23257, n23259, n31872,
    n23412, n32153, n23861, n32171, n31966, n23872, n39586, n39660, n40435,
    n32232, n23248, n23942, n23591, n40329, n40344, n23937, n23938, n32615,
    n23468, n32279, n23856, n32727, n23618, n23270, n23939, n32344, n32782,
    n31947, n32817, n23238, n23273, n32917, n28087, n33213, n40428, n40497,
    n40755, n40807, n40746, n40920, n41144, n42139, n41326, n41336, n41491,
    n29313, n41680, n41591, n41703, n41710, n41733, n40531, n41590, n41756,
    n41795, n40518, n33217, n42214, n42111, n27368, n42197, n38682, n33862,
    n23793, n23543, n23546, n23789, n23790, n33830, n23553, n34024, n34585,
    n35535, n23362, n37502, n35583, n35632, n35800, n36833, n36249, n36247,
    n36880, n36347, n36389, n36511, n36508, n37146, n37183, n37185, n36490,
    n23655, n23656, n35948, n36665, n36702, n36730, n23769, n33294, n33388,
    n33429, n23762, n23763, n23204, n23764, n23765, n37363, n38675, n38763,
    n38487, n39118, n44838, n23220, n23219, n42343, n42500, n23954, n42559,
    n42561, n30348, n30441, n26922, n42622, n42746, n30729, n23633, n30053,
    n30753, n23837, n42915, n43061, n31032, n23316, n23317, n23495, n23556,
    n31117, n23318, n31116, n23532, n30775, n43054, n44757, n43207, n43312,
    n43544, n43713, n43876, n44047, n44215, n44405, n44214, n44220, n44406,
    n44326, n44514, n23454, n40117, n31745, n23249, n32169, n39653, n32406,
    n32421, n32472, n32493, n32550, n42170, n39782, n32057, n31886, n39964,
    n39970, n40022, n40077, n40114, n40273, n32369, n23294, n23281, n29905,
    n23188, n23146, n32230, n32781, n23615, n32845, n23296, n32876, n32989,
    n33086, n42133, n40467, n40482, n40530, n40566, n40546, n40637, n40740,
    n40808, n40894, n41063, n41832, n41237, n41311, n41675, n41856, n41819,
    n41838, n41855, n41867, n41653, n41672, n41690, n41700, n41745, n41796,
    n41762, n41873, n41765, n41868, n42123, n33879, n33796, n35487, n35623,
    n35677, n23365, n24218, n24180, n35784, n27595, n24047, n35752, n36099,
    n35944, n33338, n37331, n36731, n36152, n37383, n37382, n39077, n39078,
    n33585, n23610, n23169, n32765, n23361, n33304, n23658, n23173, n22865,
    n22866, n22867, n32482, n34872, n23504, n22868, n29824, n27389, n22869,
    n43066, n27757, n23914, n24191, n24297, n22870, n22871, n22872, n22873,
    n27119, n22874, n31928, n22875, n30821, n23475, n22876, n22877, n22878,
    n22879, n22880, n22881, n22882, n22883, n22884, n22885, n28149, n22886,
    n22887, n22888, n22889, n22890, n22891, n22892, n22893, n22894, n22895,
    n22896, n22897, n40734, n34425, n22898, n34394, n23642, n22899, n27569,
    n22900, n22901, n22902, n22903, n22904, n25838, n43569, n28366, n25741,
    n26192, n22906, n40356, n23239, n34564, n30237, n28580, n30215, n22907,
    n22908, n22909, n22910, n22911, n22912, n22913, n22914, n22915, n22916,
    n22917, n22918, n22919, n22920, n22921, n27622, n22922, n22923, n22924,
    n22925, n22926, n22927, n22928, n22929, n22930, n22931, n22932, n22933,
    n22934, n22935, n22936, n22937, n22938, n29836, n23575, n30152, n22939,
    n30171, n27103, n22940, n29864, n22941, n22942, n28114, n22943, n28178,
    n22944, n28137, n22945, n22946, n22947, n22948, n22949, n22950, n22951,
    n30877, n22952, n22953, n30994, n22954, n22955, n22956, n31033, n22957,
    n22958, n22959, n22960, n22961, n22962, n22963, n28955, n22965, n22966,
    n22967, n22968, n32549, n22969, n22970, n22971, n22972, n22973, n22974,
    n22975, n22976, n22977, n22978, n23775, n23218, n25790, n23213, n22979,
    n22980, n23894, n22981, n27570, n22982, n27433, n36290, n22983, n22984,
    n22985, n22986, n22987, n22988, n22989, n22990, n23784, n22991, n22992,
    n22993, n22994, n22995, n22996, n34309, n22997, n22998, n22999, n23000,
    n23001, n23002, n23003, n23004, n23005, n23006, n23007, n23008, n23009,
    n23010, n30010, n23011, n23012, n23013, n23014, n23015, n23016, n28044,
    n23017, n23018, n23019, n27644, n23020, n23021, n23022, n23023, n23024,
    n23025, n23026, n23027, n28164, n23742, n23166, n29278, n29365, n29537,
    n29501, n23028, n29527, n23029, n28027, n35319, n42949, n23829, n28089,
    n30849, n29530, n23030, n36554, n26391, n23031, n40342, n32597, n23917,
    n23032, n23818, n23033, n23034, n32511, n23035, n23036, n23037, n23038,
    n23039, n23040, n23041, n23042, n23043, n23044, n23045, n23046, n23047,
    n23048, n32458, n23251, n25549, n44142, n23621, n23049, n40323, n40348,
    n23050, n23051, n23052, n30054, n23913, n23053, n23054, n23055, n25988,
    n23056, n23057, n23058, n23791, n31677, n23059, n23060, n23061, n23062,
    n23063, n23064, n35405, n34782, n35328, n34717, n23066, n23393, n23067,
    n33186, n23648, n23649, n23927, n23068, n23069, n37235, n23279, n29855,
    n23278, n23070, n23071, n23766, n23767, n23072, n23643, n33023, n23768,
    n23581, n29869, n33073, n23073, n44851, n23074, n29053, n23075, n23640,
    n23641, n23562, n23563, n23076, n23077, n23078, n31580, n32362, n23364,
    n32222, n23751, n23079, n23080, n23081, n32752, n23082, n33003, n28542,
    n27761, n36652, n23198, n24220, n24219, n23083, n42899, n29094, n23084,
    n23085, n28258, n23303, n30828, n44843, n25014, n23852, n23698, n23950,
    n23697, n27758, n23086, n23087, n27722, n27863, n27749, n36706, n36750,
    n23088, n23089, n39726, n23597, n23414, n23416, n27118, n23092, n36260,
    n24186, n26962, n42372, n42112, n23093, n25936, n30926, n30928, n23744,
    n23094, n23596, n23360, n32632, n23095, n41378, n23096, n23097, n23099,
    n23100, n27724, n23305, n38723, n30995, n23102, n23103, n29103, n27219,
    n24150, n23609, n23603, n31230, n23444, n42227, n31517, n23314, n24869,
    n24986, n43450, n23104, n23105, n23106, n28306, n30305, n28299, n23437,
    n23301, n41624, n23203, n27251, n27905, n27847, n27400, n27269, n26869,
    n23674, n24752, n39849, n34610, n30261, n23107, n27881, n36333, n39729,
    n23402, n23709, n30946, n28543, n42208, n23441, n23108, n23109, n27603,
    n23110, n23114, n23111, n23112, n44391, n44499, n36213, n36215, n34777,
    n24535, n23405, n27768, n23171, n23863, n23113, n27606, n31074, n43013,
    n43031, n23310, n25650, n23605, n25637, n31727, n31843, n32090, n27605,
    n31964, n23403, n27743, n23207, n23116, n23682, n23118, n23119, n23243,
    n23268, n31536, n23120, n23121, n39106, n23815, n23813, n31961, n23131,
    n27279, n27270, n23122, n23123, n27192, n23124, n23125, n23127, n23129,
    n23130, n23353, n23132, n23372, n23162, n23337, n27418, n27135, n27268,
    n27374, n27196, n27335, n27246, n27314, n27230, n27289, n27301, n27158,
    n23526, n23133, n28493, n27171, n27689, n23160, n23134, n24179, n23135,
    n23136, n23137, n27661, n29694, n25547, n27385, n28062, n23138, n23820,
    n27344, n23139, n23140, n23398, n42920, n23157, n23496, n27176, n23142,
    n27145, n23143, n27668, n25397, n27756, n27720, n23145, n27191, n23144,
    n27115, n23265, n27265, n27267, n23601, n23442, n27890, n27876, n23622,
    n32646, n28573, n23313, n25617, n31062, n25850, n23193, n23619, n23718,
    n28015, n32223, n27889, n24832, n23148, n23639, n23149, n27727, n28317,
    n32272, n27774, n32562, n23151, n27177, n23152, n27608, n27897, n23420,
    n27635, n23825, n23153, n27685, n27345, n23473, n23154, n23298, n23291,
    n23564, n23163, n23387, n23599, n23978, n23408, n28507, n27206, n23155,
    n28328, n23688, n27859, n23156, n27740, n23274, n27224, n23423, n23158,
    n23159, n32703, n32271, n42432, n23755, n23668, n23589, n23380, n23161,
    n28131, n32604, n28088, n23485, n28236, n27607, n23164, n27638, n23489,
    n23165, n23431, n23176, n31441, n23525, n28013, n23167, n27342, n23325,
    n31639, n31627, n31635, n31631, n39219, n23168, n29854, n23170, n32221,
    n28301, n23389, n23593, n23590, n23821, n23235, n23941, n23391, n32687,
    n23679, n23440, n23527, n24577, n23172, n24588, n28311, n23190, n23175,
    n28296, n23241, n23242, n23177, n32211, n32649, n32583, n32573, n30655,
    n23612, n23185, n23187, n28307, n23266, n32452, n32403, n23292, n29028,
    n32361, n23191, n23192, n27718, n27669, n23197, n23199, n24183, n33305,
    n33381, n23201, n36612, n23205, n23542, n36800, n33144, n23206, n39618,
    n39810, n23521, n30180, n29946, n31037, n23221, n28304, n32559, n30970,
    n23223, n23224, n23836, n23528, n23225, n27442, n23228, n23229, n27554,
    n27486, n27449, n23237, n28276, n29798, n23471, n23240, n32665, n39579,
    n39582, n31900, n23247, n31935, n27748, n29318, n33176, n23255, n27751,
    n29682, n23260, n23261, n31908, n27601, n28315, n23578, n30953, n23732,
    n30695, n23272, n23638, n27409, n23277, n27151, n27413, n39667, n27882,
    n32799, n27428, n23750, n32398, n25858, n23282, n23283, n23284, n30981,
    n23286, n23288, n23289, n23290, n27763, n27867, n23683, n23293, n32356,
    n32778, n32415, n23297, n32231, n43210, n23394, n32404, n32848, n25003,
    n25040, n25033, n25242, n25195, n23300, n25435, n23704, n31045, n23306,
    n23307, n23312, n23449, n31380, n23319, n25504, n30824, n23324, n23327,
    n23330, n28308, n23332, n23333, n23334, n32332, n29093, n29063, n29026,
    n23336, n23584, n32346, n23339, n32418, n23344, n23419, n23347, n28223,
    n23346, n31768, n28226, n23348, n28166, n23351, n23352, n23436, n23354,
    n23355, n35810, n38710, n23357, n23358, n35519, n35558, n35574, n23363,
    n24600, n24673, n38725, n27275, n23370, n23371, n32438, n23375, n27808,
    n23376, n23377, n23379, n23384, n23586, n32574, n23390, n43716, n39772,
    n39926, n27653, n23399, n23401, n31999, n31858, n23404, n32577, n32261,
    n32688, n29683, n32014, n23409, n23513, n23417, n23415, n32481, n23745,
    n23859, n23467, n32228, n32666, n23421, n32575, n32809, n32819, n28312,
    n23428, n23424, n23427, n23429, n23430, n32257, n23434, n23723, n23494,
    n23623, n30805, n23439, n27754, n27861, n27950, n40568, n31419, n25634,
    n23447, n23448, n25608, n23451, n23453, n44510, n23455, n23457, n44512,
    n44515, n23568, n23463, n23464, n29931, n23466, n26964, n25673, n26193,
    n40281, n23472, n23483, n27765, n27896, n40316, n23474, n23480, n32372,
    n23487, n23488, n23490, n23492, n30673, n23737, n25562, n23497, n23555,
    n31375, n23498, n23499, n23500, n28303, n28069, n23501, n25461, n23738,
    n23510, n23511, n23512, n23514, n23516, n23827, n23519, n31854, n23524,
    n23523, n29731, n27286, n27249, n27116, n27317, n27226, n27216, n27155,
    n23529, n23530, n25440, n25907, n23531, n36651, n23533, n36726, n24082,
    n23536, n24080, n36419, n36399, n23538, n24733, n23539, n23540, n23541,
    n24284, n23544, n23545, n36312, n23552, n33996, n23554, n25013, n23731,
    n23561, n27879, n27660, n29907, n23572, n28072, n23574, n29820, n29827,
    n23577, n29823, n32581, n23582, n23583, n32389, n23585, n23587, n28248,
    n23592, n28316, n33218, n23616, n32348, n27913, n23598, n24976, n31043,
    n23604, n23606, n23614, n23936, n43969, n26241, n25559, n25997, n25382,
    n31000, n23629, n42399, n23631, n30099, n30115, n30789, n28108, n29839,
    n23636, n36556, n23644, n23645, n23646, n36463, n24579, n37293, n23650,
    n23651, n23652, n23657, n23654, n24574, n23661, n29061, n32343, n23663,
    n23667, n23670, n23671, n23672, n31478, n30993, n23677, n23676, n25652,
    n31887, n23680, n29679, n31870, n23687, n27716, n23689, n27721, n28499,
    n33164, n23701, n23703, n25885, n39621, n23705, n27598, n27343, n23715,
    n23714, n23712, n27678, n23713, n23717, n25046, n25016, n25664, n23726,
    n30846, n23730, n23734, n24764, n24919, n23736, n25558, n23740, n25233,
    n25412, n23752, n23746, n32246, n32707, n36632, n23754, n24255, n36672,
    n23756, n24184, n23757, n33331, n23771, n33279, n23770, n36498, n23782,
    n23783, n31476, n25062, n23785, n23786, n33831, n23787, n23788, n23792,
    n36408, n23795, n31474, n24759, n23798, n23799, n23801, n31388, n23803,
    n23805, n30292, n29952, n25823, n29975, n29973, n32358, n32780, n31461,
    n42931, n25406, n31009, n23823, n31981, n23826, n31488, n44781, n25422,
    n31534, n25099, n31022, n31021, n30958, n23842, n30195, n29967, n29932,
    n29969, n23850, n23851, n27299, n23858, n32862, n32885, n33046, n23866,
    n28623, n23870, n23871, n32973, n32970, n31722, n31784, n23885, n23893,
    n23895, n29071, n23899, n23900, n27639, n27618, n28208, n28076, n27796,
    n31728, n29811, n23921, n28222, n28232, n31019, n23929, n30754, n25027,
    n25052, n23934, n40279, n23935, n27132, n27180, n27377, n27332, n23946,
    n23943, n25722, n31509, n42216, n33112, n30644, n30632, n26923, n25183,
    n27134, n27242, n41808, n27904, n27241, n24917, n24886, n24830, n24776,
    n23947, n26894, n23948, n23949, n23951, n42855, n23952, n23953, n23955,
    n23956, n23957, n23958, n23959, n23960, n38768, n23961, n33722, n23962,
    n23963, n40515, n23964, n42755, n23965, n23966, n23967, n28476, n23968,
    n24287, n23969, n23970, n39945, n31948, n25147, n23971, n23972, n23973,
    n23974, n23975, n23976, n39520, n40390, n32996, n33062, n23977, n24731,
    n26818, n23979, n27611, n25006, n27494, n26622, n24739, n26759, n25199,
    n24885, n27347, n24681, n25580, n26748, n25668, n24892, n27426, n27599,
    n27396, n25577, n25066, n25399, n25023, n29283, n28670, n29717, n27836,
    n29540, n28045, n27202, n27182, n25587, n25584, n25103, n25278, n27483,
    n29670, n29767, n29098, n29394, n27321, n28032, n27547, n34545, n42328,
    n24748, n44845, n26912, n31459, n25194, n43799, n27363, n28240, n29713,
    n29656, n28668, n31634, n28518, n33145, n27643, n26272, n25980, n26151,
    n25946, n26904, n26702, n25877, n26275, n25908, n25436, n25241, n43880,
    n31439, n33237, n28179, n31607, n29636, n32883, n33141, n29306, n38688,
    n36109, n24595, n24594, n36760, n37147, n25596, n25678, n26439, n26972,
    n26900, n25803, n31424, n30666, n30743, n30216, n30307, n25902, n25551,
    n25449, n31535, n43717, n44311, n44792, n43191, n27560, n31632, n29032,
    n31638, n31642, n39516, n28427, n31811, n32950, n29335, n33140, n32291,
    n32436, n41789, n41769, n40922, n40991, n41255, n27619, n40547, n24720,
    n36538, n33848, n38796, n27587, n38689, n36166, n36320, n36327, n34481,
    n38788, n37667, n26949, n42494, n30287, n42488, n30097, n42907, n43001,
    n44745, n43388, n43867, n31582, n44546, n39138, n33240, n32823, n31648,
    n39678, n39656, n39677, n31946, n39725, n39850, n32712, n32373, n33115,
    n33125, n42154, n40452, n40513, n40582, n40741, n40982, n40556, n41422,
    n41606, n41642, n41693, n41720, n41740, n42204, n41895, n38681, n38674,
    n34405, n34448, n34492, n35447, n35726, n36881, n36683, n36666, n36745,
    n38678, n37292, n24730, n38483, n39068, n39069, n37805, n37878, n38025,
    n38248, n38468, n38537, n38831, n33659, n44800, n26977, n42440, n42493,
    n31515, n42553, n30984, n42599, n43070, n42758, n42326, n42936, n43053,
    n43152, n43122, n43137, n43976, n43113, n44327, n44508, n44815, n39160,
    n29031, n39628, n39495, n32471, n39898, n40429, n40249, n40200, n29797,
    n40294, n40403, n27563, n39140, n40722, n40806, n40985, n41071, n41143,
    n41227, n41477, n41569, n41562, n41651, n41715, n41814, n41850, n41870,
    n39976, n39120, n36183, n34468, n34469, n34459, n35006, n35273, n35353,
    n35394, n35554, n35789, n37212, n35799, n35937, n36062, n35966, n36400,
    n37066, n36613, n36743, n37080, n37210, n37257, n37349, n38781, n38570,
    n37797, n37870, n37501, n37941, n38017, n38087, n38240, n38308, n38340,
    n38545, n38534, n38654, n38814, n38811, n39114, n38890, n38854, n33487,
    n33660, n42759, n42234, n42373, n42389, n42481, n42562, n42540, n42556,
    n30536, n42592, n42749, n42891, n43018, n44809, n44741, n43198, n43290,
    n43458, n43629, n43708, n43796, n43960, n44129, n44303, n44505, n42243,
    n42200, n42075, n39681, n39686, n39639, n39647, n39817, n39954, n40037,
    n42199, n40108, n40324, n40337, n41786, n40645, n40904, n40981, n41068,
    n41151, n41318, n41486, n41563, n41660, n42181, n41926, n42065, n38799,
    n34291, n34478, n34843, n35391, n35477, n35490, n35661, n35807, n35872,
    n35909, n36580, n36629, n36727, n37201, n37352, n38489, n38476, n37396,
    n39097, n39126, n33588, n44859, n43055, n44521, n39163, n39977, n40076,
    n33749, n35940, n38686, n43060, n23981, n24289, n23980, n23983, n24373,
    n23982, n23986, n23984, n23985, n23989, n23987, n23988, n23993, n34516,
    n23991, n34575, n23990, n23992, n23994, n24018, n23998, n23996, n34578,
    n23997, n24004, n24002, n34660, n24001, n24003, n24016, n24008, n24301,
    n24007, n24014, n34532, n24012, n24308, n24011, n24013, n24015, n24017,
    n36732, n24020, n24019, n24022, n24025, n24023, n24024, n24048, n24027,
    n24026, n24031, n24029, n24028, n24030, n24039, n24033, n24032, n24037,
    n24035, n24034, n24036, n24038, n24046, n24041, n24040, n24045, n24043,
    n24042, n24044, n36749, n35804, n24572, n24050, n24049, n24052, n24051,
    n24055, n24053, n24054, n24063, n24057, n24107, n35415, n24056, n24061,
    n24059, n24058, n24060, n24062, n24079, n24065, n24064, n24069, n24067,
    n24066, n24068, n24077, n24098, n35422, n24071, n24070, n24075, n24073,
    n24072, n24074, n24076, n24078, n24552, n24567, n24081, n36707, n24564,
    n24084, n24083, n24086, n24085, n24089, n24087, n24088, n24097, n24091,
    n24090, n24095, n24093, n24092, n24094, n24096, n24115, n24100, n24099,
    n24104, n24102, n24101, n24103, n24113, n24106, n24105, n24111, n24109,
    n24108, n24110, n24112, n24114, n35782, n24119, n24117, n24118, n36681,
    n24121, n24120, n24123, n24122, n24126, n24124, n24125, n24134, n24128,
    n24127, n24132, n24130, n24129, n24131, n24133, n24136, n24135, n24140,
    n24138, n24137, n24139, n24148, n24142, n35396, n24141, n24146, n24144,
    n24143, n24145, n24147, n24151, n36682, n24152, n24153, n24182, n24155,
    n24154, n24157, n24156, n24160, n24158, n24159, n24168, n24162, n24161,
    n24166, n24164, n24163, n24165, n24167, n24181, n24170, n24169, n24171,
    n24173, n24172, n24177, n24175, n24174, n24176, n24178, n35761, n24185,
    n24221, n24190, n24189, n24195, n24193, n24192, n24194, n24203, n24197,
    n24196, n24201, n24199, n24198, n24200, n24202, n24205, n24204, n24209,
    n24207, n24206, n24208, n24217, n24211, n24210, n24215, n24213, n24212,
    n24214, n24216, n24223, n24222, n24225, n24224, n24228, n24226, n24227,
    n24236, n24230, n24229, n24234, n24232, n24231, n24233, n24235, n24252,
    n24238, n24237, n24242, n24240, n24239, n24241, n24250, n24244, n24243,
    n24248, n24246, n24245, n24247, n24249, n24251, n24254, n24256, n24257,
    n37121, n37154, n37065, n24258, n36437, n24259, n24265, n36574, n36432,
    n24262, n24260, n24261, n24263, n24264, n24267, n24266, n24268, n24270,
    n24269, n24271, n24272, n24273, n36322, n24629, n36874, n24274, n24596,
    n36298, n24275, n24276, n36276, n24277, n24278, n24280, n24279, n24281,
    n36193, n24282, n36781, n24641, n36764, n24285, n36134, n33399, n33267,
    n33276, n33426, n24286, n33268, n24288, n33306, n24470, n24291, n24290,
    n24296, n24451, n24294, n24293, n24295, n24307, n24299, n24298, n24305,
    n24303, n24540, n24302, n24304, n24306, n24326, n24310, n24309, n24314,
    n24543, n24312, n24311, n24313, n24324, n24317, n24316, n24322, n24320,
    n24516, n24319, n24321, n24323, n24325, n24328, n24327, n24332, n24330,
    n24329, n24331, n24340, n24334, n24333, n24338, n24336, n24335, n24337,
    n24339, n24356, n24342, n24341, n24346, n24344, n24343, n24345, n24354,
    n24348, n24347, n24352, n24350, n24349, n24351, n24353, n24355, n24482,
    n24358, n24357, n24362, n24360, n24359, n24361, n24370, n24364, n24363,
    n24368, n24366, n24365, n24367, n24369, n24387, n24372, n24371, n24377,
    n24375, n24374, n24376, n24385, n24379, n24378, n24383, n24381, n24380,
    n24382, n24384, n24386, n24388, n24390, n34783, n24389, n24392, n24391,
    n24394, n34778, n24393, n24402, n24396, n24395, n24400, n24398, n24397,
    n24399, n24401, n24418, n24404, n24403, n24408, n24406, n24405, n24407,
    n24416, n24410, n24409, n24414, n24412, n24411, n24413, n24415, n24417,
    n24616, n24420, n24419, n24424, n24422, n24421, n24423, n24432, n24426,
    n24425, n24430, n24428, n24427, n24429, n24431, n24448, n24434, n24433,
    n24438, n24436, n24435, n24437, n24446, n24440, n24439, n24444, n24442,
    n24441, n24443, n24445, n24447, n24450, n24449, n24455, n24453, n24452,
    n24454, n24463, n24457, n24456, n24461, n24459, n24458, n24460, n24462,
    n24480, n24465, n24464, n24469, n24467, n24466, n24468, n24478, n24472,
    n24471, n24476, n24474, n24473, n24475, n24477, n24479, n24481, n24484,
    n24483, n24488, n24486, n24485, n24487, n24496, n24490, n24489, n24494,
    n24492, n24491, n24493, n24495, n24512, n24498, n24497, n24502, n24500,
    n24499, n24501, n24510, n24504, n24503, n24508, n24506, n24505, n24507,
    n24509, n24511, n24515, n24514, n24520, n24518, n24517, n24519, n24532,
    n24521, n24530, n24523, n24526, n24524, n24525, n24528, n24527, n24529,
    n24531, n24551, n24534, n24533, n24539, n24537, n24536, n24538, n24549,
    n24542, n24541, n24547, n24545, n24544, n24546, n24548, n24550, n33406,
    n24631, n24646, n36380, n36258, n33412, n37059, n37056, n35794, n24553,
    n24565, n24559, n24557, n24554, n24556, n24555, n24586, n24587, n24583,
    n24558, n24581, n36678, n24561, n24560, n24580, n36690, n24563, n24562,
    n24578, n36705, n24566, n24568, n24576, n36716, n24570, n24571, n24573,
    n36715, n24575, n36677, n24584, n24592, n24590, n36645, n24589, n36619,
    n24591, n36462, n36201, n24597, n37087, n37085, n24628, n37184, n33393,
    n24649, n24605, n24667, n24599, n24665, n38745, n24678, n33740, n24601,
    n24602, n24603, n35943, n24606, n27588, n24623, n24614, n38756, n24664,
    n24607, n24611, n24609, n24610, n24612, n24613, n24622, n24615, n24620,
    n27590, n24675, n24618, n24619, n24621, n38732, n24626, n24642, n24624,
    n27586, n24627, n38703, n27583, n36962, n37295, n37302, n37317, n37278,
    n37256, n37259, n37188, n37058, n24638, n37140, n37062, n36968, n36863,
    n36916, n36884, n33413, n36869, n36849, n36811, n24630, n33417, n33433,
    n24652, n33386, n39129, n24636, n24635, n38706, n27584, n38730, n36774,
    n37369, n24637, n37294, n37260, n37218, n37064, n36990, n37012, n24639,
    n36975, n36919, n36893, n36951, n36909, n24640, n36864, n36842, n36792,
    n24654, n33382, n38744, n38704, n38705, n24643, n24644, n37010, n36879,
    n36836, n36770, n24645, n24653, n33384, n33432, n24648, n33313, n36932,
    n37356, n24647, n33365, n24663, n24651, n24650, n24661, n24659, n24656,
    n24655, n33419, n24657, n24658, n33395, n33362, n24660, n24662, n24671,
    n24666, n24669, n24670, n24672, n24674, n24676, n24677, n38692, n24716,
    n24679, n24692, n24690, n24693, n37428, n24685, n24680, n24682, n24684,
    n24683, n24699, n24698, n24701, n24687, n24686, n24697, n24694, n24688,
    n24689, n24691, n24705, n24695, n24696, n24718, n24700, n24702, n24703,
    n33737, n24706, n39005, n39112, n24707, n33742, n24708, n24709, n24726,
    n24713, n24715, n24711, n38677, n24712, n24714, n24723, n24717, n24719,
    n24722, n24724, n24725, n24727, n24729, n24728, n39056, n38803, n38810,
    n24732, n33319, n25574, n24741, n24737, n24736, n24740, n24749, n24743,
    n24742, n24747, n26629, n24745, n24744, n24746, n24769, n24905, n24750,
    n24751, n24758, n25088, n24756, n24755, n24757, n24947, n24761, n24760,
    n24767, n24766, n24768, n24771, n24770, n24774, n24772, n24773, n24777,
    n24775, n24785, n24779, n24778, n24781, n24780, n24782, n24784, n24786,
    n24788, n24787, n24792, n24790, n24789, n24791, n24800, n24794, n24793,
    n24798, n24796, n24795, n24797, n24799, n24803, n24804, n25123, n24806,
    n24805, n24808, n24807, n24812, n26851, n24810, n24809, n24811, n24833,
    n25100, n24817, n24816, n24821, n24819, n24818, n24820, n24831, n24822,
    n24824, n24823, n24828, n24826, n24825, n24827, n24829, n24835, n24834,
    n24839, n24837, n24836, n24838, n24847, n24841, n24840, n24845, n24843,
    n24842, n24844, n24846, n24863, n24853, n24911, n24849, n24848, n24850,
    n24852, n24855, n24854, n24859, n24857, n24856, n24858, n24860, n24862,
    n25002, n24864, n24929, n24867, n24866, n24871, n24868, n24870, n24879,
    n24873, n24872, n24877, n24875, n24874, n24876, n24881, n24880, n24884,
    n24883, n24887, n24895, n24889, n24888, n24891, n24890, n24894, n24900,
    n24899, n24904, n24902, n24901, n24903, n24910, n24906, n24908, n24907,
    n24909, n24913, n24912, n24916, n24914, n24915, n24918, n24926, n24920,
    n24922, n24921, n24966, n24931, n24930, n24933, n25513, n24932, n24935,
    n24934, n24944, n24938, n24937, n24942, n24940, n24939, n24941, n24943,
    n24946, n24945, n24951, n24949, n24948, n24950, n24959, n24953, n24952,
    n24957, n24955, n24954, n24956, n24958, n24960, n24963, n24964, n25021,
    n24971, n24968, n24967, n24970, n24982, n24975, n24974, n24980, n24978,
    n24977, n24979, n24981, n24999, n24984, n24983, n24988, n24985, n24987,
    n24997, n24991, n24990, n24995, n24993, n24992, n24994, n24996, n24998,
    n25018, n25000, n25041, n25034, n25053, n25832, n25007, n25005, n25015,
    n25010, n25731, n25693, n25012, n31438, n25599, n25691, n31568, n25029,
    n25019, n25020, n25025, n25024, n25026, n25028, n30634, n25031, n25185,
    n25032, n25035, n25187, n25038, n25036, n25037, n25039, n25703, n42393,
    n44748, n25044, n25045, n25047, n25051, n25049, n25050, n25061, n25059,
    n25056, n25057, n31497, n25058, n25060, n25064, n25063, n25068, n25067,
    n25070, n26483, n25069, n25078, n25072, n26035, n25071, n25076, n25074,
    n26326, n25073, n25075, n25077, n25097, n25080, n25079, n25084, n25082,
    n31463, n25081, n25083, n25095, n25294, n25087, n25267, n25086, n25093,
    n25091, n26349, n25090, n25092, n25094, n25096, n25098, n25102, n25101,
    n25105, n25104, n26154, n25106, n25115, n25109, n25108, n25113, n25111,
    n25110, n25112, n25114, n25133, n25117, n25116, n25122, n25465, n25120,
    n25119, n25121, n25131, n25125, n25124, n25129, n25127, n25126, n25128,
    n25130, n25132, n25172, n25135, n25137, n25136, n25138, n25141, n25140,
    n25143, n25142, n25146, n25144, n25145, n25155, n25149, n25148, n25153,
    n25151, n25150, n25152, n25154, n25171, n25157, n25156, n25161, n25159,
    n25158, n25160, n25169, n25163, n25162, n25167, n25165, n25164, n25166,
    n25168, n25170, n25174, n25177, n25173, n25175, n25181, n25176, n25179,
    n25178, n25180, n25391, n25184, n25186, n25188, n25236, n25190, n25191,
    n25238, n25193, n25192, n25198, n26750, n26876, n25197, n25201, n25200,
    n25203, n26612, n25202, n25211, n25205, n25204, n25209, n25207, n25206,
    n25208, n25210, n25228, n25213, n25212, n25217, n25215, n25214, n25216,
    n25226, n25219, n25218, n25224, n25481, n25220, n25222, n25337, n25221,
    n25223, n25225, n25227, n25229, n25231, n25230, n44307, n43729, n43718,
    n25237, n44153, n25240, n25239, n25277, n25245, n25244, n25247, n25246,
    n25250, n25248, n25249, n25258, n25252, n25251, n25256, n25254, n25253,
    n25255, n25257, n25275, n25260, n25259, n25264, n25262, n26577, n25261,
    n25263, n25273, n25266, n25265, n25271, n25269, n25268, n25270, n25272,
    n25274, n25276, n25312, n25280, n25279, n25282, n25281, n25285, n25283,
    n25284, n25293, n25287, n25286, n25291, n25289, n25288, n25290, n25292,
    n25310, n26879, n25296, n25295, n25300, n25298, n25297, n25299, n25308,
    n25302, n25301, n25306, n25304, n25303, n25305, n25307, n25309, n25311,
    n25347, n25313, n25320, n25316, n25315, n25318, n25317, n25319, n25328,
    n25322, n25321, n25326, n25324, n25323, n25325, n25327, n25345, n25330,
    n26686, n25329, n25334, n25332, n25331, n25333, n25343, n25336, n25335,
    n25341, n25339, n25338, n25340, n25342, n25344, n25346, n25380, n25349,
    n25348, n25351, n25350, n25353, n26800, n25352, n25361, n25355, n25354,
    n25359, n26870, n25357, n25356, n25358, n25360, n25378, n25364, n25363,
    n25368, n25366, n26817, n25365, n25367, n25376, n25370, n26858, n25369,
    n25374, n25372, n25371, n25373, n25375, n25377, n25379, n25383, n25381,
    n25384, n25390, n25413, n25428, n25437, n25385, n25444, n25386, n25456,
    n25387, n25388, n25389, n25396, n25394, n25419, n25395, n42948, n25404,
    n25400, n25402, n25401, n25403, n25407, n25405, n25408, n25409, n31010,
    n25410, n25423, n25416, n25415, n25417, n25418, n25420, n25421, n25425,
    n25431, n25427, n25429, n25430, n25432, n25434, n25433, n25438, n25439,
    n25442, n25441, n25445, n25446, n25447, n25448, n25450, n25453, n25451,
    n25452, n25454, n25460, n25501, n25458, n25459, n30947, n25463, n25542,
    n25467, n25466, n25471, n26707, n25469, n25468, n25470, n25479, n25473,
    n25472, n25477, n25475, n25474, n25476, n25478, n25480, n25497, n25483,
    n25482, n25487, n25485, n25484, n25486, n25495, n25489, n25488, n25493,
    n26847, n25491, n25490, n25492, n25494, n25496, n25500, n25502, n30951,
    n25503, n30949, n25506, n31332, n25505, n25508, n25509, n25511, n26617,
    n25510, n25517, n25512, n25515, n25514, n25516, n25521, n26875, n25519,
    n25518, n25520, n25541, n25523, n25522, n25539, n25525, n25524, n25529,
    n25527, n25526, n25528, n25537, n25531, n25530, n25535, n25533, n25532,
    n25534, n25536, n25538, n25540, n25543, n30927, n25545, n31287, n25544,
    n30879, n31233, n25546, n30903, n31286, n30907, n31261, n25548, n31216,
    n25552, n30844, n30864, n31189, n30823, n30898, n25553, n25554, n30804,
    n31134, n25557, n25556, n25560, n31105, n30706, n31078, n31075, n30674,
    n25842, n25561, n31063, n30683, n31048, n25563, n31049, n31035, n25564,
    n25567, n25565, n25566, n25568, n25569, n25570, n44522, n44841, n25598,
    n25588, n25590, n25571, n25581, n25573, n25572, n25583, n25578, n25575,
    n25576, n25585, n25579, n25632, n25582, n25627, n25586, n25640, n25591,
    n25589, n25613, n31512, n26911, n25597, n25600, n25659, n25643, n25602,
    n25636, n25605, n25603, n25604, n25607, n25606, n25628, n25626, n25611,
    n25610, n25612, n25625, n25618, n25620, n25622, n25621, n25623, n25624,
    n25630, n25631, n25633, n25635, n25641, n25638, n25644, n25649, n25651,
    n26985, n25653, n25655, n25654, n25656, n25657, n25658, n25676, n31503,
    n25663, n25662, n25666, n25665, n25672, n25667, n25671, n25670, n25697,
    n25674, n31493, n31423, n25684, n25681, n25680, n31451, n31506, n25682,
    n25683, n25690, n25686, n25687, n25688, n25689, n25696, n44842, n25694,
    n25695, n25698, n25701, n25699, n25700, n31444, n25702, n25704, n25705,
    n25706, n27066, n25714, n25712, n27064, n31232, n25710, n31315, n44753,
    n42993, n42965, n42972, n31395, n31381, n31348, n31318, n31277, n31243,
    n31187, n31173, n25711, n31167, n27068, n27072, n27097, n25840, n25707,
    n43014, n25713, n25708, n43032, n31248, n42968, n31404, n31312, n31347,
    n31317, n31279, n27065, n31241, n31170, n27069, n27096, n25839, n25715,
    n43027, n25720, n25717, n31090, n25716, n31059, n25718, n25719, n25721,
    n25848, n25723, n25724, n25728, n25727, n25725, n25726, n42486, n25729,
    n42439, n42485, n25733, n25732, n25734, n42438, n25736, n25735, n25737,
    n42420, n42384, n25739, n25738, n25740, n42385, n25743, n25742, n25744,
    n31401, n25746, n25745, n25747, n25749, n25748, n25750, n31367, n25752,
    n25751, n25753, n31352, n25755, n25754, n25756, n31338, n25758, n25757,
    n25759, n30330, n25761, n25760, n25762, n30314, n25764, n25763, n25765,
    n30291, n25767, n25766, n25768, n30267, n25770, n25769, n25771, n30243,
    n25773, n25772, n25774, n30226, n25779, n25776, n25775, n25777, n30199,
    n30182, n25781, n25780, n25782, n30181, n25784, n25783, n25785, n30156,
    n25787, n25786, n25788, n30138, n25792, n25791, n25793, n27082, n25795,
    n25794, n25796, n27104, n25798, n25797, n25799, n30083, n25801, n25800,
    n25802, n30055, n25806, n25805, n25807, n30033, n25809, n25808, n25810,
    n30014, n25812, n25811, n25813, n29994, n25815, n25814, n25816, n29972,
    n25818, n25817, n25819, n29950, n25821, n25820, n29911, n29936, n29913,
    n25825, n25824, n29914, n25826, n25827, n25831, n25829, n25828, n25830,
    n42503, n25835, n25834, n25836, n25847, n43026, n31102, n25841, n31119,
    n31079, n31036, n31031, n25843, n25844, n25846, n30637, n25845, n25849,
    n25920, n25895, n25857, n25851, n25855, n25853, n42919, n25852, n25854,
    n25856, n25881, n25860, n25867, n25865, n25861, n25863, n25862, n25864,
    n25866, n42459, n44801, n25869, n25876, n25874, n25870, n25872, n25871,
    n25873, n25875, n42482, n25880, n25878, n25879, n42458, n25882, n25884,
    n43072, n25894, n25890, n25886, n25888, n25887, n25889, n25892, n25903,
    n42906, n25891, n25893, n42431, n25901, n25896, n25899, n25897, n25898,
    n25900, n25905, n42894, n25904, n25906, n25909, n25911, n25910, n25914,
    n25918, n42363, n25913, n25915, n25926, n25917, n25924, n25928, n25919,
    n42350, n25922, n25921, n25923, n25925, n30999, n25935, n25927, n25933,
    n25938, n25929, n42327, n25931, n25930, n25932, n25934, n25945, n25937,
    n25943, n25939, n42306, n25941, n25940, n25942, n25944, n25948, n25947,
    n25952, n25950, n25949, n25951, n25960, n25954, n25953, n25958, n25956,
    n25955, n25957, n25959, n25977, n25962, n25961, n25964, n26481, n25963,
    n25967, n25965, n25966, n25975, n25969, n25968, n25973, n25971, n25970,
    n25972, n25974, n25976, n25978, n25987, n25979, n25985, n25991, n25981,
    n42290, n25983, n25982, n25984, n25986, n30956, n25989, n25995, n25993,
    n30937, n25992, n25994, n25996, n30323, n25999, n25998, n26003, n26001,
    n26000, n26002, n26011, n26005, n26004, n26009, n26007, n26006, n26008,
    n26010, n26027, n26013, n26012, n26017, n26015, n26014, n26016, n26025,
    n26019, n26018, n26023, n26021, n26020, n26022, n26024, n26026, n26028,
    n26030, n26029, n26066, n30911, n26033, n42872, n26032, n26034, n26037,
    n26036, n26041, n26039, n26038, n26040, n26049, n26043, n26042, n26047,
    n26045, n26044, n26046, n26048, n26051, n26050, n26055, n26053, n26052,
    n26054, n26063, n26057, n26056, n26061, n26059, n26058, n26060, n26062,
    n26064, n26065, n30304, n30921, n26071, n26067, n26069, n26068, n26070,
    n30258, n26110, n26113, n30893, n26109, n26074, n26073, n26078, n26076,
    n26075, n26077, n26086, n26080, n26079, n26084, n26082, n26081, n26083,
    n26085, n26102, n26088, n26087, n26092, n26090, n26089, n26091, n26100,
    n26094, n26093, n26098, n26096, n26095, n26097, n26099, n26101, n26103,
    n26107, n42877, n26105, n26104, n26106, n26108, n26111, n26112, n30871,
    n26150, n26115, n26114, n26119, n26117, n26116, n26118, n26127, n26121,
    n26120, n26125, n26123, n26122, n26124, n26126, n26143, n26129, n26128,
    n26131, n26130, n26133, n26799, n26132, n26141, n26135, n26134, n26139,
    n26137, n26136, n26138, n26140, n26142, n26144, n26148, n42882, n26146,
    n26145, n26147, n26149, n30238, n26327, n26158, n26153, n26152, n26156,
    n26155, n26157, n26166, n26160, n26159, n26164, n26162, n26161, n26163,
    n26165, n26182, n26168, n26167, n26172, n26170, n26169, n26171, n26180,
    n26174, n26173, n26178, n26176, n26175, n26177, n26179, n26181, n26183,
    n26191, n30606, n26189, n26231, n26185, n30858, n26187, n26186, n26188,
    n26190, n26195, n26194, n26199, n26197, n26196, n26198, n26207, n26201,
    n26200, n26205, n26203, n26202, n26204, n26206, n26223, n26209, n26208,
    n26213, n26211, n26210, n26212, n26221, n26215, n26214, n26219, n26217,
    n26216, n26218, n26220, n26222, n26224, n26230, n26225, n26228, n26226,
    n26227, n26229, n26234, n26232, n30839, n26233, n30196, n26236, n26235,
    n26240, n26238, n26237, n26239, n26248, n26242, n26246, n26244, n26243,
    n26245, n26247, n26264, n26250, n26249, n26254, n26252, n26251, n26253,
    n26262, n26256, n26255, n26260, n26258, n26257, n26259, n26261, n26263,
    n26265, n26274, n26266, n26268, n30815, n26270, n26269, n26271, n30172,
    n30807, n26316, n26277, n26276, n26281, n26279, n26278, n26280, n26289,
    n26283, n26282, n26287, n26285, n26284, n26286, n26288, n26307, n26291,
    n26290, n26294, n26292, n26293, n26297, n26295, n26296, n26305, n26299,
    n26298, n26303, n26301, n26300, n26302, n26304, n26306, n26308, n26314,
    n26309, n26312, n26310, n26311, n26313, n26315, n30153, n26317, n30059,
    n26398, n26319, n26324, n26322, n26321, n26323, n26331, n26325, n26329,
    n26328, n26330, n26347, n26333, n26332, n26337, n26335, n26334, n26336,
    n26345, n26339, n26338, n26343, n26341, n26340, n26342, n26344, n26346,
    n26355, n26348, n26353, n26351, n26350, n26352, n26354, n26480, n26356,
    n26364, n26358, n26357, n26362, n26359, n26361, n26363, n26372, n26366,
    n26365, n26370, n26368, n26367, n26369, n26371, n26388, n26374, n26373,
    n26378, n26376, n26375, n26377, n26386, n26380, n26379, n26384, n26382,
    n26381, n26383, n26385, n26387, n26479, n26390, n26389, n26396, n26903,
    n26394, n26392, n26393, n26395, n26397, n30770, n26438, n26401, n26400,
    n26405, n26403, n26402, n26404, n26429, n26407, n26406, n26411, n26409,
    n26408, n26410, n26427, n26413, n26412, n26417, n26415, n26414, n26416,
    n26425, n26419, n26418, n26423, n26421, n26420, n26422, n26424, n26426,
    n26428, n26430, n26436, n26431, n26434, n26432, n26433, n26435, n26437,
    n30795, n26478, n26441, n26440, n26445, n26443, n26442, n26444, n26449,
    n26447, n26446, n26448, n26469, n26451, n26450, n26467, n26453, n26452,
    n26457, n26455, n26454, n26456, n26465, n26459, n26458, n26463, n26461,
    n26460, n26462, n26464, n26466, n26468, n26470, n26476, n26471, n26474,
    n26472, n26473, n26475, n26477, n30131, n26647, n26485, n26484, n26487,
    n26486, n26490, n26488, n26489, n26498, n26492, n26491, n26496, n26494,
    n26493, n26495, n26497, n26514, n26500, n26499, n26504, n26502, n26501,
    n26503, n26512, n26506, n26505, n26510, n26508, n26507, n26509, n26511,
    n26513, n26648, n26515, n26521, n26516, n26519, n26517, n26518, n26520,
    n26524, n30734, n26523, n30032, n26525, n26566, n30781, n26565, n26528,
    n26527, n26532, n26530, n26529, n26531, n26540, n26534, n26533, n26538,
    n26536, n26535, n26537, n26539, n26556, n26542, n26541, n26546, n26544,
    n26543, n26545, n26554, n26548, n26547, n26552, n26550, n26549, n26551,
    n26553, n26555, n26557, n26563, n26558, n26561, n26559, n26560, n26562,
    n26564, n30114, n26567, n26609, n30758, n26608, n26570, n26569, n26574,
    n26572, n26571, n26573, n26583, n26576, n26575, n26581, n26579, n26578,
    n26580, n26582, n26599, n26585, n26584, n26587, n26586, n26589, n26588,
    n26597, n26591, n26590, n26595, n26593, n26592, n26594, n26596, n26598,
    n26600, n26606, n26601, n26604, n26602, n26603, n26605, n26607, n30074,
    n26610, n26611, n26614, n26613, n26616, n26615, n26619, n26618, n26628,
    n26621, n26620, n26626, n26624, n26623, n26625, n26627, n26646, n26632,
    n26631, n26636, n26634, n26633, n26635, n26644, n26638, n26637, n26642,
    n26640, n26639, n26641, n26643, n26645, n26663, n26662, n26649, n26655,
    n26650, n26653, n26651, n26652, n26654, n26659, n26657, n30716, n26658,
    n30011, n26705, n26665, n26664, n26669, n26667, n26666, n26668, n26677,
    n26671, n26670, n26675, n26673, n26672, n26674, n26676, n26694, n26679,
    n26678, n26683, n26681, n26680, n26682, n26692, n26685, n26684, n26690,
    n26688, n26687, n26689, n26691, n26693, n26706, n26695, n26701, n26696,
    n26699, n26697, n26698, n26700, n26704, n30700, n26703, n29992, n26786,
    n26709, n26708, n26713, n26711, n26710, n26712, n26721, n26715, n26714,
    n26719, n26717, n26716, n26718, n26720, n26737, n26723, n26722, n26727,
    n26725, n26724, n26726, n26735, n26729, n26728, n26733, n26731, n26730,
    n26732, n26734, n26736, n26784, n26738, n26744, n26739, n26742, n26740,
    n26741, n26743, n26747, n30688, n26746, n29968, n26752, n26749, n26751,
    n26755, n26754, n26758, n26756, n26757, n26767, n26761, n26760, n26765,
    n26763, n26762, n26764, n26766, n26783, n26769, n26768, n26773, n26771,
    n26770, n26772, n26781, n26775, n26774, n26779, n26777, n26776, n26778,
    n26780, n26782, n26798, n26785, n26797, n26787, n26793, n26788, n26791,
    n26789, n26790, n26792, n26796, n30668, n26795, n29949, n26845, n26802,
    n26801, n26804, n26803, n26808, n26805, n26807, n26816, n26810, n26809,
    n26814, n26812, n26811, n26813, n26815, n26834, n26820, n26819, n26824,
    n26822, n26821, n26823, n26832, n26826, n26825, n26830, n26828, n26827,
    n26829, n26831, n26833, n26846, n26835, n26841, n26836, n26839, n26837,
    n26838, n26840, n26844, n30658, n26843, n29933, n26889, n26850, n26849,
    n26855, n26853, n26852, n26854, n26865, n26857, n26856, n26863, n26861,
    n26860, n26862, n26864, n26887, n26868, n26867, n26874, n26872, n26871,
    n26873, n26885, n26878, n26877, n26883, n26881, n26880, n26882, n26884,
    n26886, n26888, n26891, n26898, n26892, n26896, n26893, n26895, n26897,
    n26902, n30647, n26901, n29910, n26906, n26905, n26907, n26909, n26921,
    n26918, n26916, n26913, n26915, n30346, n26917, n26919, n26920, n26924,
    n26959, n26926, n26925, n26930, n26928, n26927, n26929, n26951, n26932,
    n26931, n26936, n26934, n26933, n26935, n26938, n26937, n26942, n26940,
    n26939, n26941, n26947, n26944, n26943, n26945, n26946, n26948, n26950,
    n26952, n26953, n26958, n26955, n26957, n26960, n26961, n26974, n27056,
    n26963, n26969, n26965, n26966, n26967, n26968, n26970, n26971, n42469,
    n26976, n30639, n31566, n26978, n26979, n26990, n44676, n44671, n26992,
    n26984, n30263, n44661, n30080, n30079, n44621, n44611, n44586, n44576,
    n44566, n26980, n42404, n42379, n42355, n42334, n42313, n42296, n30328,
    n30264, n30265, n26981, n30245, n30218, n30202, n30141, n26982, n30075,
    n26983, n30060, n30015, n30017, n26991, n29976, n26987, n26998, n26995,
    n29959, n44692, n44686, n26993, n26988, n29924, n26989, n27004, n44681,
    n30005, n29960, n29943, n26994, n27002, n26996, n26997, n27000, n42470,
    n26999, n27001, n27003, n27010, n27006, n27005, n27008, n27007, n27009,
    n27046, n27016, n27012, n27011, n27014, n27013, n27015, n27017, n27019,
    n27018, n27023, n27021, n27020, n27022, n27028, n27025, n27024, n27026,
    n27027, n27044, n27030, n27029, n27034, n27032, n27031, n27033, n27042,
    n27036, n27035, n27040, n27038, n27037, n27039, n27041, n27043, n33460,
    n42232, n27047, n44530, n27052, n41918, n27049, n27048, n27050, n27051,
    n27053, n27058, n27054, n27055, n27057, n27059, n30790, n27062, n31151,
    n27061, n27090, n27063, n30786, n27089, n31231, n31162, n31268, n31244,
    n27067, n31259, n27079, n27075, n31242, n27070, n31150, n27071, n27087,
    n27074, n42966, n27073, n27077, n27076, n27078, n31147, n27080, n27081,
    n27085, n30396, n27083, n30780, n27084, n27086, n27088, n27095, n27091,
    n27093, n27092, n27094, n27099, n27098, n27100, n31137, n27101, n27110,
    n27105, n30390, n27108, n30766, n31131, n27106, n27107, n27109, n29853,
    n27111, n33131, n27113, n41887, n27112, n27114, n33265, n42079, n27117,
    n27123, n27120, n27122, n27131, n29688, n27200, n27124, n27129, n27127,
    n27126, n27128, n27130, n27147, n27133, n27137, n27139, n27138, n27143,
    n27141, n27140, n27142, n27144, n27146, n27612, n27179, n27148, n27154,
    n27150, n27152, n27153, n27164, n27156, n27157, n27160, n27159, n27161,
    n27178, n27166, n27165, n27169, n27168, n27167, n27170, n27175, n27172,
    n27174, n27173, n27181, n27185, n27187, n27186, n27190, n27189, n27260,
    n27188, n27194, n27193, n27198, n27197, n27207, n27199, n27201, n27205,
    n27204, n27203, n40486, n27276, n27211, n27210, n27215, n27212, n27214,
    n27225, n28017, n27217, n27223, n27220, n27222, n28020, n27227, n27232,
    n27229, n27231, n27240, n27234, n27233, n27238, n40545, n27236, n27235,
    n27237, n27239, n27244, n27243, n27248, n27476, n29116, n27247, n27257,
    n29126, n27250, n27255, n27253, n27252, n27254, n27256, n27273, n27259,
    n27258, n27264, n27262, n27261, n27263, n27271, n27453, n27266, n29111,
    n27272, n27277, n27626, n27274, n40552, n27278, n40519, n27281, n27280,
    n27285, n27283, n27282, n27284, n27294, n29502, n27288, n27287, n27292,
    n27290, n29498, n27291, n27293, n27310, n27295, n27297, n27296, n27298,
    n27308, n27300, n27302, n27306, n27304, n27303, n27305, n27307, n27309,
    n27312, n27311, n27316, n27313, n27315, n27325, n27318, n27323, n27421,
    n27320, n27322, n27324, n27327, n27326, n27331, n27329, n27328, n27330,
    n27340, n27333, n27338, n27337, n27339, n27341, n27358, n27357, n27346,
    n27354, n27349, n27444, n27355, n27352, n27351, n27364, n27353, n27539,
    n27356, n27543, n27362, n27361, n27360, n27522, n27525, n27367, n27366,
    n27365, n27551, n27370, n39150, n27369, n27406, n27372, n27371, n27376,
    n27373, n27375, n27386, n27378, n27384, n27380, n27382, n27381, n27383,
    n27403, n27388, n27387, n27393, n27391, n27390, n27392, n27401, n27394,
    n27395, n27399, n27398, n27397, n27402, n27404, n27627, n27405, n27407,
    n42206, n27564, n27408, n27411, n27845, n27417, n29718, n29355, n27415,
    n29660, n27852, n27414, n27416, n27427, n27420, n27419, n27425, n29602,
    n27423, n29569, n28763, n27422, n27424, n27443, n29099, n27431, n27429,
    n29591, n27430, n27437, n27432, n29592, n27435, n27434, n27436, n27438,
    n29436, n27440, n27439, n27441, n31598, n27445, n27448, n27452, n27450,
    n27451, n27457, n29519, n27455, n27454, n27456, n27465, n27459, n27458,
    n27463, n27461, n29447, n27460, n27462, n27464, n27482, n27467, n27466,
    n27471, n27469, n27468, n27470, n27475, n27473, n29597, n27472, n27474,
    n27480, n27478, n27477, n27479, n27481, n27484, n27550, n27485, n28060,
    n28051, n28245, n27487, n27548, n27489, n27488, n27493, n27491, n27490,
    n27492, n27502, n27496, n27495, n27500, n29558, n27497, n27499, n27520,
    n27504, n27503, n27508, n27506, n27505, n27507, n27514, n27512, n27511,
    n27513, n27518, n27516, n28647, n27515, n27517, n27519, n28554, n28285,
    n27524, n27521, n27565, n27523, n28241, n27527, n27528, n27526, n27535,
    n27530, n27529, n27533, n27655, n27537, n27532, n27534, n27542, n40456,
    n27538, n27540, n28054, n27541, n27545, n27544, n27546, n27559, n27553,
    n27555, n27557, n27556, n27558, n27567, n27568, n27575, n27571, n27572,
    n27574, n27573, n42180, n27576, n27577, n42186, n27578, n27582, n27580,
    n27581, n27585, n27589, n35745, n27594, n27592, n27591, n27593, n27597,
    n27596, n27600, n27602, n27604, n27628, n28250, n27609, n28261, n27616,
    n27614, n27615, n27623, n27640, n27617, n27620, n27621, n27624, n28318,
    n27625, n27630, n27629, n27634, n27633, n27636, n27642, n27641, n27645,
    n27647, n27646, n27651, n27649, n27648, n27650, n27652, n27654, n27657,
    n27658, n27663, n27659, n27662, n27683, n27664, n27666, n27667, n40343,
    n27671, n27670, n27673, n27675, n27674, n27676, n33230, n27682, n28057,
    n27680, n27679, n27681, n27687, n27684, n27686, n27744, n27696, n27691,
    n27690, n27694, n27692, n27745, n27698, n27697, n27701, n27699, n27703,
    n27702, n27734, n27705, n27704, n27709, n27708, n27706, n27707, n27735,
    n27714, n27711, n27710, n27712, n28325, n27713, n27717, n27719, n28327,
    n27726, n27725, n27728, n28332, n27731, n27730, n28335, n27739, n27733,
    n27737, n27738, n27736, n27741, n27746, n27750, n28678, n27752, n29424,
    n27753, n27755, n27760, n27892, n28700, n28681, n27762, n27764, n29222,
    n41574, n28682, n27766, n27772, n27770, n27769, n27771, n27778, n27776,
    n27782, n27783, n29520, n27786, n27784, n27785, n27787, n27789, n27788,
    n27794, n27792, n27790, n27791, n27793, n27809, n27798, n27797, n27802,
    n27800, n27799, n27801, n27804, n27803, n27806, n27805, n27807, n33116,
    n27843, n27812, n27811, n27816, n27814, n27813, n27815, n27825, n29491,
    n27819, n27818, n27823, n27821, n27820, n27822, n27824, n27842, n27827,
    n27826, n27831, n27829, n27828, n27830, n27835, n27833, n27832, n27834,
    n27840, n27838, n27837, n27839, n27841, n28565, n28767, n27846, n27851,
    n27848, n27850, n27860, n40421, n27854, n27857, n27855, n27856, n27858,
    n27862, n27866, n27864, n27865, n27875, n27868, n28766, n27873, n27869,
    n27871, n27870, n27872, n27874, n27878, n27885, n27888, n27891, n29350,
    n27895, n29356, n27894, n28840, n27899, n28845, n27902, n28865, n27901,
    n27903, n29651, n27907, n27906, n27911, n41766, n27909, n27910, n27912,
    n27946, n27915, n27914, n27920, n27918, n27917, n27919, n27928, n27922,
    n27921, n27926, n27924, n27923, n27925, n27927, n27944, n27930, n27929,
    n27934, n27932, n27931, n27933, n27938, n27936, n27935, n27937, n27942,
    n27940, n27939, n27941, n27943, n28609, n27945, n27947, n27949, n28905,
    n27948, n27953, n27951, n27952, n27964, n27955, n27954, n27962, n27958,
    n27957, n27960, n27988, n27959, n27961, n27963, n27978, n27966, n27965,
    n27970, n27968, n27967, n27969, n27976, n29712, n27972, n27971, n27974,
    n28904, n27973, n27975, n27977, n27980, n27979, n27985, n27983, n27982,
    n27984, n27994, n27987, n27986, n27992, n27990, n27989, n27991, n27993,
    n28010, n27996, n27995, n28000, n27998, n27997, n27999, n28004, n28002,
    n28001, n28003, n28008, n28006, n28005, n28007, n28009, n28616, n28011,
    n28014, n28016, n28019, n29730, n28018, n28024, n28022, n28021, n28023,
    n28026, n28025, n28031, n28029, n28928, n28028, n28030, n28050, n28035,
    n28034, n28039, n28037, n28036, n28038, n28043, n28041, n28040, n28042,
    n28048, n28046, n28047, n28049, n28077, n28053, n28052, n28091, n28055,
    n28056, n28059, n28095, n28058, n28099, n28061, n28063, n39790, n28065,
    n28066, n28067, n28068, n39544, n28074, n39559, n28075, n28079, n28078,
    n28081, n28083, n28082, n28084, n39498, n28085, n32533, n32529, n32530,
    n28086, n28093, n28092, n39605, n39629, n40302, n28096, n39682, n33123,
    n28100, n28097, n28098, n28101, n40320, n42096, n28102, n33111, n39665,
    n40319, n40301, n28105, n28103, n28104, n40284, n39583, n40289, n28106,
    n28107, n28110, n40368, n28109, n28111, n28112, n32532, n39521, n28113,
    n32488, n28115, n28116, n39479, n28117, n32975, n32509, n28121, n28119,
    n39458, n28120, n32502, n32487, n28122, n28123, n32486, n28124, n32508,
    n28125, n28128, n39439, n28129, n32927, n32469, n28130, n32468, n28132,
    n28133, n28134, n39416, n28135, n32455, n28136, n32899, n32454, n28155,
    n28146, n28138, n28139, n28140, n28184, n28141, n32771, n32345, n28143,
    n39296, n28187, n32360, n28144, n29022, n28158, n28147, n39340, n28148,
    n32390, n28151, n39313, n28153, n32808, n32374, n28162, n28156, n28157,
    n28159, n32831, n32402, n28161, n39376, n28163, n32858, n32432, n28165,
    n28191, n28167, n32849, n32437, n28168, n28169, n28170, n28171, n28177,
    n28172, n28173, n28175, n39255, n29062, n28176, n28182, n28180, n28201,
    n28181, n29075, n29067, n28183, n29024, n28200, n39280, n28185, n28186,
    n28188, n29021, n28189, n32401, n28190, n32431, n39402, n28192, n28193,
    n28195, n28194, n29020, n28197, n28196, n28198, n28199, n28203, n39243,
    n28202, n29066, n28204, n28205, n39225, n28206, n32306, n28207, n32307,
    n28209, n28210, n28215, n28211, n28212, n31833, n28213, n28993, n32292,
    n28214, n28216, n28217, n31814, n28218, n28219, n28220, n32277, n28224,
    n28221, n29825, n32259, n28225, n31790, n28227, n29808, n28228, n32256,
    n28231, n28229, n28230, n28234, n28233, n31746, n32224, n28235, n28237,
    n28238, n28239, n28281, n28243, n28244, n28247, n33221, n28249, n28269,
    n28251, n28253, n28252, n28514, n28254, n28255, n28256, n28257, n28260,
    n28259, n28264, n28262, n28263, n28268, n41920, n39153, n28265, n41909,
    n31608, n33236, n28266, n28267, n28278, n28270, n28271, n28273, n28272,
    n28274, n28275, n28277, n28279, n28280, n28282, n28284, n29019, n28287,
    n28286, n28288, n40322, n28289, n28292, n40306, n40305, n40308, n28293,
    n28294, n28297, n28302, n28310, n32925, n32851, n32859, n32376, n28313,
    n32807, n29054, n28314, n33220, n29017, n28324, n28320, n28319, n28322,
    n42040, n28321, n28323, n28326, n28330, n28329, n28331, n28333, n28334,
    n28336, n28343, n28338, n28337, n28341, n28339, n28340, n28342, n39580,
    n28351, n28346, n28345, n28349, n32586, n28348, n28350, n28358, n28353,
    n28352, n28356, n28354, n28355, n28357, n32563, n28365, n28360, n28359,
    n28363, n28361, n28362, n28364, n28373, n28368, n28367, n28371, n28369,
    n28370, n28372, n28379, n28375, n28374, n28377, n32974, n28376, n28378,
    n32512, n28386, n28381, n28380, n28384, n28382, n28383, n28385, n32492,
    n28393, n28388, n28387, n28391, n28389, n28390, n28392, n28400, n28395,
    n28394, n28398, n28396, n28397, n28399, n28407, n28402, n28401, n28405,
    n28403, n28404, n28406, n32440, n28413, n28409, n28408, n28411, n32422,
    n28410, n28412, n32420, n28419, n28415, n28414, n28417, n41984, n28416,
    n28418, n28426, n28421, n28420, n28424, n28422, n28423, n28425, n28434,
    n28429, n28428, n28432, n28430, n28431, n28433, n28440, n28436, n28435,
    n28438, n41997, n28437, n28439, n31936, n28447, n28442, n28441, n28445,
    n28443, n28444, n28446, n28454, n28449, n28448, n28452, n28450, n28451,
    n28453, n28461, n28456, n28455, n28459, n28457, n28458, n28460, n29072,
    n28467, n28463, n28462, n28465, n32310, n28464, n28466, n28473, n28469,
    n28468, n28471, n42018, n28470, n28472, n28480, n28475, n28474, n28478,
    n42025, n28477, n28479, n31809, n31788, n28486, n28482, n28481, n28484,
    n42030, n28483, n28485, n28492, n28488, n28487, n28490, n42035, n28489,
    n28491, n31785, n33184, n28496, n28495, n28497, n28541, n28502, n28501,
    n28504, n28503, n28506, n28505, n28510, n31968, n28508, n28509, n28511,
    n28517, n28513, n28524, n28515, n28516, n33143, n32736, n28523, n29038,
    n29043, n28519, n29073, n33015, n28522, n33061, n40377, n33074, n33002,
    n28520, n32991, n32852, n29074, n32671, n28521, n28531, n28581, n33065,
    n32995, n29050, n29078, n29866, n32673, n28533, n28536, n33185, n28525,
    n28526, n33229, n28527, n28529, n28528, n40325, n33064, n28530, n29873,
    n32993, n28532, n32637, n29867, n28534, n28535, n28539, n32635, n28537,
    n32236, n28538, n28540, n29015, n28547, n28555, n29897, n28545, n29898,
    n28544, n28546, n29882, n28551, n28549, n40205, n28548, n28550, n28559,
    n28566, n42179, n28556, n28557, n28558, n28564, n28562, n28560, n28561,
    n28563, n33113, n28571, n28567, n28569, n28568, n28570, n39659, n28574,
    n28579, n28576, n28578, n28587, n28585, n28583, n40210, n28582, n28584,
    n39626, n28590, n28588, n28589, n33094, n28594, n33104, n28592, n28591,
    n28593, n28600, n28598, n40215, n28597, n28599, n33093, n28602, n28606,
    n28604, n40220, n28603, n28605, n28608, n28607, n39587, n28613, n28611,
    n40225, n28610, n28612, n28615, n28614, n33072, n28617, n28621, n28619,
    n40231, n28618, n28620, n33045, n28622, n33026, n28627, n28625, n40236,
    n28624, n28626, n33025, n33027, n28629, n28628, n28633, n29474, n28631,
    n28630, n28632, n28646, n28634, n28638, n28636, n28635, n28637, n28640,
    n29469, n28639, n28644, n29478, n28642, n29475, n28641, n28643, n28645,
    n28649, n28648, n28654, n28650, n28652, n28651, n28653, n28659, n28657,
    n28655, n28656, n28658, n28660, n29340, n28667, n28665, n28663, n28661,
    n28662, n28664, n28666, n33006, n28672, n28671, n28677, n28675, n28673,
    n28674, n28676, n28688, n28680, n29437, n28679, n28686, n28684, n28683,
    n28685, n28687, n28706, n28691, n28690, n28695, n28693, n28692, n28694,
    n28699, n28697, n28696, n28698, n28704, n28702, n28701, n28703, n28705,
    n39762, n28711, n28709, n28707, n28708, n28710, n28713, n28712, n32971,
    n28716, n28715, n28720, n28718, n28717, n28719, n28733, n28721, n28725,
    n28723, n28722, n28724, n28727, n28726, n28731, n29466, n28729, n29465,
    n28728, n28730, n28732, n28736, n28735, n28738, n28737, n28740, n28739,
    n28746, n28741, n28744, n28742, n28743, n28745, n28747, n39736, n28754,
    n28752, n28750, n28748, n28749, n28751, n28753, n32951, n28757, n28755,
    n28756, n28761, n28759, n28758, n28760, n28773, n28762, n28765, n28764,
    n28771, n28769, n28768, n28770, n28772, n28790, n28775, n28774, n28779,
    n28777, n28776, n28778, n28783, n28781, n28780, n28782, n28788, n28786,
    n28784, n28785, n28787, n28789, n39744, n28795, n28793, n28791, n28792,
    n28794, n28797, n28796, n32933, n28836, n28799, n28798, n28803, n28801,
    n28800, n28802, n28811, n28805, n28804, n28809, n28807, n28806, n28808,
    n28810, n28815, n28813, n28812, n28814, n28817, n28816, n28826, n29125,
    n28819, n28818, n28824, n29449, n28822, n28820, n28821, n28823, n28825,
    n28827, n39737, n28834, n28832, n28830, n28828, n28829, n28831, n28833,
    n32902, n28838, n28837, n28844, n28839, n28842, n28841, n28843, n28854,
    n28848, n28846, n28847, n28852, n28850, n28849, n28851, n28853, n28871,
    n28856, n28855, n28860, n28858, n28857, n28859, n28864, n28862, n28861,
    n28863, n28869, n28867, n28866, n28868, n28870, n29343, n28876, n28874,
    n28872, n28873, n28875, n28878, n28877, n28881, n28880, n28885, n28883,
    n28882, n28884, n28897, n29568, n28889, n28887, n28886, n28888, n28891,
    n28890, n28895, n28893, n28892, n28894, n28896, n28911, n28901, n28899,
    n28898, n28900, n28903, n28902, n28909, n28907, n28906, n28908, n28910,
    n39717, n28918, n28916, n28914, n28912, n28913, n28915, n28917, n32863,
    n28920, n28919, n28926, n28921, n28924, n28922, n28923, n28925, n28937,
    n28927, n28930, n28929, n28935, n28933, n28931, n28932, n28934, n28936,
    n28954, n28939, n28938, n28943, n28941, n28940, n28942, n28947, n28945,
    n28944, n28946, n28952, n28948, n28950, n28949, n28951, n28953, n29609,
    n28960, n28958, n28956, n28957, n28959, n28962, n28961, n32835, n28966,
    n32818, n28964, n40118, n28963, n28965, n28971, n28969, n40123, n28968,
    n28970, n28975, n28973, n40128, n28972, n28974, n32151, n28979, n28977,
    n40133, n28976, n28978, n32136, n29033, n28984, n28982, n40138, n28981,
    n28983, n28988, n28986, n40143, n28985, n28987, n28992, n28990, n40148,
    n28989, n28991, n32089, n28997, n28995, n40153, n28994, n28996, n31844,
    n29001, n28999, n40158, n28998, n29000, n31805, n29006, n29004, n40164,
    n29003, n29005, n31765, n29010, n32245, n29008, n40170, n29007, n29009,
    n31764, n31763, n32015, n29011, n29012, n29014, n29016, n29018, n29023,
    n29064, n29027, n29030, n32333, n29059, n39267, n31917, n29037, n29034,
    n39248, n29035, n32335, n29036, n29049, n29041, n32800, n29039, n29040,
    n29046, n29042, n32921, n29044, n29045, n32803, n32784, n29047, n32772,
    n29048, n29057, n29055, n29052, n29051, n32969, n32861, n32830, n32791,
    n32770, n29056, n29058, n29060, n29065, n29069, n29068, n29091, n39230,
    n29085, n32734, n29083, n29076, n29077, n29080, n29079, n32732, n29081,
    n32324, n29082, n29084, n29089, n32105, n29088, n29090, n29092, n29095,
    n29757, n29097, n29756, n29096, n29110, n29100, n29102, n29101, n29107,
    n29105, n29104, n29106, n29108, n29109, n29115, n29113, n29112, n29114,
    n29137, n29119, n29117, n29118, n29135, n29121, n29120, n29132, n29122,
    n29123, n29130, n29128, n29127, n29129, n29131, n29133, n29134, n29136,
    n29680, n29139, n29138, n29143, n29141, n29140, n29142, n29151, n29145,
    n29144, n29149, n29147, n29479, n29146, n29148, n29150, n29167, n29153,
    n29152, n29157, n29155, n29154, n29156, n29165, n29159, n29158, n29163,
    n29161, n29160, n29162, n29164, n29166, n29618, n29169, n29168, n29178,
    n29170, n29175, n29173, n29172, n29174, n29176, n29177, n29182, n29180,
    n29760, n29179, n29181, n29199, n29184, n29183, n29193, n29186, n29185,
    n29190, n29187, n29189, n29191, n29192, n29197, n29195, n29194, n29196,
    n29198, n29619, n29621, n29200, n29203, n29201, n29202, n29211, n29205,
    n29204, n29209, n29207, n29206, n29208, n29210, n29215, n29213, n29212,
    n29214, n29234, n29217, n29216, n29221, n29219, n29218, n29220, n29232,
    n29223, n29225, n29224, n29230, n29228, n29227, n29229, n29231, n29233,
    n29625, n29624, n29628, n29236, n29235, n29245, n29238, n29237, n29242,
    n29240, n29239, n29241, n29243, n29244, n29249, n29247, n29246, n29248,
    n29266, n29251, n29250, n29260, n29253, n29252, n29257, n29255, n29254,
    n29256, n29258, n29259, n29264, n29262, n29261, n29263, n29265, n29627,
    n29630, n29631, n29267, n29269, n29268, n29277, n29271, n29270, n29275,
    n29273, n29272, n29274, n29276, n29282, n29280, n29279, n29281, n29300,
    n29286, n29284, n29285, n29294, n29288, n29287, n29292, n29290, n29289,
    n29291, n29293, n29298, n29296, n29403, n29295, n29297, n29299, n29637,
    n29301, n29681, n29303, n29302, n29312, n29310, n41089, n29308, n40648,
    n40553, n41768, n29304, n29305, n41869, n40432, n29307, n41493, n29309,
    n29328, n29316, n40992, n29315, n29317, n29323, n29321, n40823, n29322,
    n29324, n29325, n29327, n29329, n29334, n29332, n29333, n29337, n29336,
    n29338, n29339, n39773, n29341, n29342, n29345, n29344, n29349, n29347,
    n29346, n29348, n29364, n29352, n29425, n29351, n29354, n29353, n29358,
    n29450, n29357, n29362, n29360, n29359, n29361, n29363, n29377, n29367,
    n29366, n29371, n29369, n29368, n29370, n29375, n29373, n29372, n29374,
    n29376, n31914, n29379, n29378, n29383, n29381, n29380, n29382, n29391,
    n29385, n29384, n29389, n29387, n29386, n29388, n29390, n29409, n29393,
    n29392, n29400, n29398, n29396, n29395, n29397, n29399, n29407, n29402,
    n29401, n29405, n29404, n29406, n29408, n31932, n29615, n29411, n29410,
    n29415, n29413, n29412, n29414, n29423, n29417, n29416, n29421, n29419,
    n29418, n29420, n29422, n29446, n29429, n29427, n29428, n29431, n29430,
    n29435, n29433, n29432, n29434, n29444, n29438, n29442, n29440, n29439,
    n29441, n29443, n29445, n31951, n29448, n29452, n29451, n29464, n29454,
    n29453, n29458, n29456, n29455, n29457, n29462, n29460, n29459, n29461,
    n29463, n29487, n29468, n29467, n29473, n29471, n29470, n29472, n29485,
    n29477, n29476, n29483, n29481, n29480, n29482, n29484, n29486, n31905,
    n29490, n29488, n29489, n29496, n29494, n29492, n29493, n29495, n29508,
    n29500, n29499, n29506, n29504, n29503, n29505, n29507, n29526, n29510,
    n29509, n29514, n29512, n29511, n29513, n29518, n29516, n29515, n29517,
    n29524, n29522, n29521, n29523, n29525, n31904, n29612, n29529, n29528,
    n29535, n29533, n29531, n29532, n29534, n29547, n29539, n29538, n29545,
    n29543, n29541, n29542, n29544, n29546, n29564, n29549, n29548, n29553,
    n29551, n29550, n29552, n29557, n29555, n29554, n29556, n29562, n29560,
    n29559, n29561, n29563, n39698, n29567, n29566, n29573, n29571, n29570,
    n29572, n29587, n29579, n29578, n29585, n29583, n29701, n29582, n29584,
    n29586, n29608, n29590, n29589, n29596, n29594, n29593, n29595, n29601,
    n29599, n29598, n29600, n29606, n29604, n29603, n29605, n29607, n31906,
    n29610, n39708, n29611, n29613, n29614, n29616, n29617, n29620, n31897,
    n29622, n29623, n31889, n31888, n29626, n29629, n31881, n29632, n29634,
    n29635, n29638, n31871, n29639, n29640, n29642, n29641, n29650, n29644,
    n29643, n29648, n29646, n29645, n29647, n29649, n29655, n29653, n29652,
    n29654, n29676, n29659, n29657, n29658, n29668, n29662, n29661, n29666,
    n29664, n29663, n29665, n29667, n29674, n29672, n29671, n29673, n29675,
    n29684, n29677, n31865, n29678, n31859, n29686, n31860, n29685, n29728,
    n29691, n29689, n29690, n29700, n29693, n29692, n29698, n29695, n29697,
    n29699, n29705, n29703, n29702, n29704, n29726, n29707, n29706, n29711,
    n29708, n29710, n29724, n29714, n29716, n29715, n29722, n29720, n29719,
    n29721, n29723, n29725, n29727, n29729, n29732, n29734, n29733, n29738,
    n29736, n29735, n29737, n29747, n29741, n29740, n29745, n29743, n29742,
    n29744, n29746, n29773, n29748, n29751, n29750, n29771, n29755, n29754,
    n29769, n29759, n29758, n29765, n29763, n29762, n29764, n29766, n29768,
    n29770, n29772, n29796, n29779, n29775, n29774, n29777, n42056, n29776,
    n29778, n29841, n29786, n29782, n29781, n29784, n42045, n29783, n29785,
    n31723, n29792, n29788, n29787, n29790, n42050, n29789, n29791, n31680,
    n29794, n31682, n29793, n29795, n32617, n29863, n29862, n29802, n29804,
    n32227, n29806, n29807, n29809, n29816, n29812, n29814, n29815, n29817,
    n29818, n29819, n29821, n31705, n32638, n32198, n29822, n31681, n32184,
    n29826, n31596, n29828, n29830, n32199, n29832, n29834, n29833, n29835,
    n29837, n29838, n29840, n29851, n29849, n29845, n29844, n29847, n42055,
    n29846, n29848, n29850, n42137, n42176, n29852, n29860, n31626, n31628,
    n31630, n31636, n31640, n31644, n31650, n31652, n31649, n31647, n31645,
    n31643, n31641, n31637, n31633, n31629, n31625, n31622, n31601, n40338,
    n40304, n40330, n29858, n29878, n29856, n29857, n29859, n29909, n29881,
    n29865, n29871, n29868, n32713, n32655, n32618, n29870, n29877, n33124,
    n29874, n29872, n32616, n29875, n29876, n29879, n29880, n31725, n29886,
    n29884, n40182, n29883, n29885, n31724, n31701, n29890, n29888, n29887,
    n29889, n31702, n29895, n29893, n40194, n29892, n29894, n31696, n29903,
    n29902, n29900, n29899, n29901, n29904, n29906, n29908, n29930, n29912,
    n29915, n29922, n30036, n30349, n29920, n29918, n29916, n29917, n29919,
    n29921, n29928, n29923, n29926, n29925, n29927, n29929, n29935, n29934,
    n29948, n29940, n29938, n29937, n29939, n29941, n29942, n29944, n29945,
    n29947, n29966, n29951, n31047, n29958, n29954, n29953, n29956, n29955,
    n29957, n29964, n29962, n29961, n29963, n29965, n29971, n29970, n29990,
    n29974, n31061, n29979, n29996, n29977, n29978, n29982, n29980, n29981,
    n29988, n29984, n29983, n29986, n29985, n29987, n29989, n30698, n30009,
    n31082, n30004, n29995, n30002, n30000, n29998, n29997, n29999, n30001,
    n30003, n30007, n30006, n30008, n30012, n30713, n30495, n30030, n31092,
    n30028, n30048, n44666, n30016, n30047, n30041, n30062, n30020, n30018,
    n30019, n30026, n30371, n30024, n30022, n30021, n30023, n30025, n30027,
    n30029, n30031, n30117, n30052, n30035, n30034, n31109, n30046, n30376,
    n30040, n30038, n30037, n30039, n30044, n30042, n30043, n30045, n30050,
    n30049, n30051, n30073, n30057, n31118, n30071, n30746, n30069, n30061,
    n30063, n30067, n30065, n30064, n30066, n30068, n30070, n30072, n30096,
    n44651, n30101, n30076, n30119, n44646, n30100, n30077, n30078, n30094,
    n30185, n30137, n30118, n30082, n30081, n30092, n30084, n31138, n30086,
    n30085, n30090, n30088, n30087, n30089, n30091, n30093, n30095, n30098,
    n30765, n30113, n30111, n30107, n30105, n30103, n30102, n30104, n30106,
    n30109, n30108, n30110, n30112, n30116, n30778, n30130, n44641, n30120,
    n30128, n30122, n30121, n30126, n30124, n30123, n30125, n30127, n30129,
    n30151, n30136, n30134, n42367, n30132, n30133, n30135, n30149, n44636,
    n30147, n30139, n31148, n30145, n30158, n30142, n30184, n30157, n30143,
    n30144, n30146, n30148, n30150, n30803, n30170, n30155, n30154, n30168,
    n31177, n30166, n30159, n30162, n30160, n30161, n30164, n30163, n30165,
    n30167, n30169, n30173, n30814, n30194, n30175, n30177, n30176, n30179,
    n30178, n30192, n30183, n31194, n30190, n30188, n30186, n30187, n30189,
    n30191, n30193, n30837, n30589, n30214, n30198, n30197, n30212, n31204,
    n30210, n44616, n30219, n30201, n30200, n30247, n30205, n30203, n30204,
    n30208, n30206, n30207, n30209, n30211, n30213, n30217, n30854, n30601,
    n30236, n30225, n30220, n30222, n30221, n30223, n30224, n30234, n30227,
    n31222, n30232, n30230, n30229, n30231, n30233, n30235, n30239, n30869,
    n30256, n30242, n30240, n30241, n30254, n31236, n30244, n30252, n30246,
    n30248, n30250, n30249, n30251, n30253, n30255, n30260, n30259, n30284,
    n30616, n30282, n30262, n30313, n30280, n30306, n30288, n30266, n30278,
    n30268, n31265, n30276, n30274, n30272, n30270, n30271, n30273, n30275,
    n30277, n30279, n30281, n30285, n30303, n30286, n44602, n30290, n30289,
    n30301, n31290, n30299, n30297, n30295, n30293, n30294, n30296, n30298,
    n30300, n30302, n30919, n30322, n30326, n44596, n30312, n30308, n30310,
    n30309, n30311, n30320, n30318, n31303, n30316, n30315, n30317, n30319,
    n30321, n30325, n30324, n42506, n30345, n44591, n30343, n30329, n30341,
    n30331, n42507, n30339, n30337, n30335, n30333, n30334, n30336, n30338,
    n30340, n30342, n30344, n30347, n30353, n30351, n30350, n30352, n30357,
    n30355, n30354, n30356, n30361, n30359, n30358, n30360, n30362, n30366,
    n30364, n30363, n30365, n30370, n30368, n30367, n30369, n30375, n30373,
    n30372, n30374, n30380, n30378, n30377, n30379, n30385, n30383, n30381,
    n30382, n30384, n30389, n30387, n30386, n30388, n30395, n30393, n30391,
    n30392, n30394, n30547, n30400, n30398, n30397, n30399, n30404, n30402,
    n30401, n30403, n30408, n30406, n30405, n30407, n30578, n30412, n30410,
    n30409, n30411, n30416, n30414, n30413, n30415, n30421, n30419, n30417,
    n30418, n30420, n30425, n30423, n30422, n30424, n30430, n30428, n30426,
    n30427, n30429, n30435, n30433, n30431, n30432, n30434, n30439, n30437,
    n30436, n30438, n30452, n30442, n30592, n30444, n30443, n42818, n30446,
    n30445, n30450, n30448, n30447, n30449, n30451, n30462, n30454, n30453,
    n30617, n30456, n30455, n30460, n30458, n30457, n30459, n30461, n30463,
    n30473, n30465, n30464, n30622, n30467, n30466, n30471, n30469, n30468,
    n30470, n30472, n30483, n30475, n30474, n42805, n30477, n30476, n30481,
    n30479, n30478, n30480, n30482, n30484, n30494, n30486, n30485, n42800,
    n30488, n30487, n30492, n30490, n30489, n30491, n30493, n30505, n30497,
    n30496, n42795, n30499, n30498, n30503, n30501, n30500, n30502, n30504,
    n30515, n30507, n30506, n42790, n30509, n30508, n30513, n30511, n30510,
    n30512, n30514, n30525, n30517, n30516, n42785, n30519, n30518, n30523,
    n30521, n30520, n30522, n30524, n30535, n30527, n30526, n42781, n30529,
    n30528, n30533, n30531, n30530, n30532, n30534, n30546, n30538, n30537,
    n42777, n30540, n30539, n30544, n30542, n30541, n30543, n30545, n30557,
    n30549, n30548, n42598, n30551, n30550, n30555, n30553, n30552, n30554,
    n30556, n30567, n30559, n30558, n42604, n30561, n30560, n30565, n30563,
    n30562, n30564, n30566, n30577, n30569, n30568, n42610, n30571, n30570,
    n30575, n30573, n30572, n30574, n30576, n30588, n30580, n30579, n42615,
    n30582, n30581, n30586, n30584, n30583, n30585, n30587, n30600, n30591,
    n30590, n42620, n30594, n30593, n30598, n30596, n30595, n30597, n30599,
    n30610, n30603, n30605, n30604, n42887, n30608, n30607, n30609, n30614,
    n30612, n30611, n30613, n30621, n42814, n30619, n30618, n30620, n30626,
    n42810, n30624, n30623, n30625, n30630, n30628, n30627, n30629, n44791,
    n30631, n30643, n44837, n30635, n30636, n30641, n31571, n30638, n42944,
    n30640, n30642, n30651, n31034, n30646, n30649, n30648, n30650, n30656,
    n30664, n30653, n30661, n31038, n30659, n30660, n30662, n30672, n31052,
    n30667, n30670, n30669, n30671, n30686, n30675, n30678, n30705, n30677,
    n30682, n30680, n30679, n30681, n31046, n30685, n30693, n30691, n31065,
    n30689, n30690, n30692, n30697, n30694, n31070, n30696, n30704, n31083,
    n30699, n30702, n30701, n30703, n30712, n30709, n30707, n30708, n30710,
    n31073, n30711, n30720, n31093, n30714, n30715, n30718, n30717, n30719,
    n30728, n30742, n30722, n30721, n30731, n30730, n30724, n30723, n30726,
    n30725, n31089, n30727, n30740, n31101, n30738, n31110, n30733, n30732,
    n30736, n30735, n30737, n30739, n30752, n30750, n31122, n30745, n30744,
    n30748, n30747, n30749, n30751, n30764, n31129, n30762, n31139, n30757,
    n30755, n30756, n30760, n30759, n30761, n30763, n30774, n30769, n30768,
    n30772, n30771, n30773, n30777, n30776, n30785, n30779, n30783, n30782,
    n30784, n30788, n30787, n30802, n31146, n30800, n31154, n30794, n30793,
    n30798, n30796, n30797, n30799, n30801, n30813, n31183, n30811, n31179,
    n30806, n30809, n30808, n30810, n30812, n30820, n30818, n31196, n30816,
    n30817, n30819, n30836, n30822, n30834, n30830, n30827, n30829, n30832,
    n30831, n30833, n31186, n30835, n30843, n31207, n30838, n30841, n30840,
    n30842, n30853, n30929, n30848, n30847, n30866, n30850, n31202, n30852,
    n30863, n31224, n30857, n30856, n30861, n30859, n30860, n30862, n30868,
    n30865, n31214, n30867, n30876, n31237, n30870, n30874, n30872, n30873,
    n30875, n30888, n30882, n30880, n30881, n30884, n30886, n30885, n31255,
    n30887, n30897, n30890, n31266, n30892, n30895, n30894, n30896, n30906,
    n30901, n30900, n30909, n30902, n30904, n31258, n30905, n30918, n30910,
    n31276, n30916, n30914, n31292, n30912, n30913, n30915, n30917, n30925,
    n31304, n30920, n30923, n30922, n30924, n30935, n30936, n30931, n30930,
    n30933, n30932, n31300, n30934, n31329, n30945, n30943, n30941, n31323,
    n30939, n30938, n30940, n30942, n30944, n30948, n30969, n30968, n30952,
    n30955, n30954, n31337, n30967, n30959, n42572, n30960, n30965, n30963,
    n31339, n30961, n30962, n30964, n30966, n31346, n30979, n42579, n30977,
    n30972, n30975, n31353, n30973, n30974, n30976, n30978, n30991, n30983,
    n30989, n30987, n31371, n30985, n30986, n30988, n30990, n30998, n30996,
    n30997, n31387, n31008, n31001, n42587, n31006, n31389, n31002, n31004,
    n31003, n31005, n31007, n42921, n31011, n31013, n42910, n31015, n31014,
    n31016, n42898, n31018, n31017, n31020, n31411, n31030, n42371, n31028,
    n31398, n31024, n31026, n31025, n31027, n31029, n31041, n31039, n31040,
    n31042, n31044, n31058, n31056, n31054, n31050, n31051, n31053, n31055,
    n31057, n31060, n31069, n31067, n31064, n31066, n31068, n31072, n31071,
    n31088, n31077, n31076, n31095, n31081, n31080, n31086, n31084, n31085,
    n31087, n31100, n31098, n31094, n31096, n31097, n31099, n31115, n31103,
    n31104, n31108, n31106, n31107, n31113, n31111, n31112, n31114, n31128,
    n31126, n31124, n31120, n31121, n31123, n31125, n31127, n31145, n31136,
    n31130, n31133, n31132, n31135, n31143, n31142, n31140, n31141, n31144,
    n31160, n31158, n31149, n31156, n31152, n31153, n31155, n31157, n31159,
    n42967, n31164, n31161, n31163, n31215, n31166, n31165, n31176, n31168,
    n31169, n31172, n31171, n31218, n31174, n31191, n31175, n31182, n31178,
    n31180, n31181, n31185, n31184, n31201, n31188, n31190, n31193, n31192,
    n31199, n31195, n31197, n31198, n31200, n31213, n31203, n31211, n31205,
    n31209, n31206, n31208, n31210, n31212, n31229, n31217, n31221, n31219,
    n31220, n31227, n31223, n31225, n31226, n31228, n31283, n31301, n31289,
    n31234, n31235, n31240, n31238, n31239, n31254, n31251, n31269, n31246,
    n31245, n31247, n31249, n31262, n31250, n31252, n31253, n31257, n31256,
    n31275, n31260, n31264, n31263, n31273, n31267, n31271, n31270, n31272,
    n31274, n31299, n31278, n31282, n31280, n31281, n31302, n31284, n31285,
    n31297, n31288, n31295, n31291, n31293, n31294, n31296, n31298, n31311,
    n31309, n31307, n31305, n31306, n31308, n31310, n31314, n31313, n31378,
    n31362, n31333, n31316, n31328, n31320, n31319, n31321, n31334, n31322,
    n31326, n31324, n31325, n31327, n31331, n31330, n31336, n31335, n31344,
    n31342, n42512, n31340, n31341, n31343, n31364, n31345, n31360, n31358,
    n31350, n31349, n31351, n31361, n31356, n42518, n31354, n31355, n31357,
    n31359, n31366, n31363, n31365, n31374, n31369, n42323, n31372, n31373,
    n31377, n31376, n31386, n31379, n31382, n31396, n31406, n31383, n31384,
    n31385, n31394, n31392, n42342, n31390, n31391, n31393, n31397, n31399,
    n31403, n42533, n31402, n31410, n31405, n31408, n31407, n31409, n31413,
    n31412, n31414, n31425, n31498, n31416, n31433, n31418, n31421, n31422,
    n31430, n31471, n31426, n31428, n31427, n31429, n31432, n42390, n31434,
    n31435, n31437, n31436, n31440, n31442, n31443, n31543, n31467, n31448,
    n31447, n31450, n31452, n31475, n31458, n31455, n31453, n31454, n31456,
    n31457, n31465, n31460, n31462, n44712, n31464, n31466, n44713, n31469,
    n31468, n31559, n31470, n31473, n31529, n31472, n31492, n31487, n44719,
    n31485, n31483, n31477, n31481, n31479, n44784, n31480, n31482, n31484,
    n44721, n31486, n31490, n31489, n31491, n43046, n31522, n31496, n42228,
    n31494, n31495, n42235, n31499, n31500, n42248, n31501, n31520, n31504,
    n31505, n31507, n31511, n31510, n31514, n31513, n31516, n44832, n31518,
    n31519, n31521, n31533, n31523, n31527, n31525, n31526, n31531, n31530,
    n43047, n31532, n31565, n31540, n31538, n44729, n31537, n31539, n44732,
    n31542, n31552, n31549, n31544, n31546, n31545, n44749, n31547, n31548,
    n31550, n31551, n31553, n31557, n31554, n31556, n31560, n31558, n31563,
    n31561, n31562, n31564, n31567, n31569, n31576, n31572, n31574, n31575,
    n31587, n44517, n31578, n31577, n31579, n31589, n31581, n31584, n31583,
    n31585, n44519, n31586, n31588, n31590, n31592, n31591, n43049, n31610,
    n31593, n31594, n31675, n31600, n31597, n31599, n39683, n31621, n31603,
    n31602, n41893, n31604, n31605, n33133, n31606, n31619, n31676, n31609,
    n31613, n31615, n31611, n31612, n31614, n31617, n31616, n31618, n31620,
    n31673, n31624, n31623, n42095, n32201, n32233, n32263, n32294, n39231,
    n39272, n39324, n39367, n39396, n39453, n39485, n39531, n39565, n39613,
    n31654, n31653, n39675, n31656, n31655, n39652, n39644, n39612, n39598,
    n40293, n39564, n39549, n39550, n39530, n39510, n39511, n39484, n39462,
    n39461, n39444, n39419, n39394, n39379, n39360, n39333, n39336, n39317,
    n39297, n39271, n39259, n39258, n39261, n39215, n39217, n31845, n31824,
    n32280, n31798, n31777, n32248, n31754, n32213, n31713, n32187, n31671,
    n31672, n31674, n31679, n33135, n31678, n31695, n31688, n31686, n31684,
    n31683, n31685, n31687, n31693, n42097, n31690, n31691, n31692, n31694,
    n31698, n32625, n31697, n32633, n31721, n31704, n31703, n31719, n31712,
    n31710, n31706, n31708, n31707, n31709, n31711, n31717, n31714, n31715,
    n31716, n31718, n31720, n32650, n31744, n31726, n32651, n31742, n31735,
    n31733, n31729, n31731, n31730, n31732, n31734, n31740, n31737, n31738,
    n31739, n31741, n31743, n31760, n31753, n31751, n31747, n31749, n31748,
    n31750, n31752, n31758, n31755, n31756, n31757, n31759, n31762, n31761,
    n31767, n31766, n32669, n32031, n31783, n31769, n31776, n31774, n31770,
    n31772, n31771, n31773, n31775, n31781, n31778, n31779, n31780, n31782,
    n31787, n32668, n31786, n32262, n32690, n31804, n31797, n31795, n31791,
    n31793, n31792, n31794, n31796, n31802, n31799, n31800, n31801, n31803,
    n31808, n32699, n31807, n32709, n31830, n31812, n32710, n31823, n31821,
    n31819, n31815, n31817, n31816, n31818, n31820, n31822, n31828, n31825,
    n31826, n31827, n31829, n32728, n31842, n31840, n31838, n31834, n31836,
    n31835, n31837, n31839, n31841, n31851, n32743, n31849, n31846, n31847,
    n31848, n31850, n31853, n31852, n31856, n31855, n31857, n32000, n31864,
    n31862, n31861, n31863, n31869, n31867, n31866, n31868, n31874, n31873,
    n32030, n31878, n31876, n31875, n31877, n31880, n31879, n31883, n31882,
    n31885, n31884, n31893, n31891, n31890, n32071, n31892, n31895, n31894,
    n31899, n32074, n31898, n39214, n31903, n31902, n31911, n39699, n39701,
    n31941, n31940, n31939, n31923, n31922, n31921, n31907, n31909, n32088,
    n31910, n31913, n31912, n31916, n32117, n31915, n31920, n31918, n31919,
    n31927, n31925, n31924, n32120, n31926, n39275, n31931, n31930, n31934,
    n32135, n31933, n39308, n31938, n31937, n31945, n31943, n31942, n32150,
    n31944, n39325, n31950, n31949, n31953, n32167, n31952, n31957, n31956,
    n31959, n31963, n31960, n31962, n31965, n31967, n33231, n31970, n31987,
    n31972, n31985, n39828, n31973, n31980, n39835, n31976, n31975, n40195,
    n31978, n31977, n31979, n31983, n39839, n31982, n31984, n31986, n31997,
    n31993, n31989, n31988, n40189, n31991, n31990, n31992, n31995, n31994,
    n31996, n31998, n32013, n32011, n32001, n32007, n32003, n32002, n40183,
    n32005, n32004, n32006, n32009, n32008, n32010, n32012, n32029, n32016,
    n32027, n32017, n32023, n32019, n32018, n40177, n32021, n32020, n32022,
    n32025, n32024, n32026, n32028, n32044, n32042, n32032, n32038, n32034,
    n32033, n40171, n32036, n32035, n32037, n32040, n32039, n32041, n32043,
    n32045, n32056, n32046, n32052, n32048, n32047, n40165, n32050, n32049,
    n32051, n32054, n32053, n32055, n32059, n32058, n32070, n32060, n32066,
    n32062, n32061, n40159, n32064, n32063, n32065, n32068, n32067, n32069,
    n32073, n32072, n32087, n32085, n32075, n32081, n32077, n32076, n40565,
    n32079, n32078, n32080, n32083, n32082, n32084, n32086, n32104, n32091,
    n39224, n32102, n32092, n32098, n32094, n32093, n40543, n32096, n32095,
    n32097, n32100, n32099, n32101, n32103, n39242, n32116, n32106, n32112,
    n32108, n32107, n40528, n32110, n32109, n32111, n32114, n32113, n32115,
    n32119, n32118, n32134, n32121, n32132, n32122, n32128, n32124, n32123,
    n40510, n32126, n32125, n32127, n32130, n32129, n32131, n32133, n32149,
    n39270, n32147, n32137, n32143, n32139, n32138, n40495, n32141, n32140,
    n32142, n32145, n32144, n32146, n32148, n32166, n32152, n39290, n32164,
    n32154, n32160, n32156, n32155, n40480, n32158, n32157, n32159, n32162,
    n32161, n32163, n32165, n32183, n39328, n32181, n32170, n32177, n32173,
    n32172, n40465, n32175, n32174, n32176, n32179, n32178, n32180, n32182,
    n32196, n32185, n32614, n32194, n32192, n32190, n32619, n32188, n32189,
    n32191, n32193, n32195, n32210, n32208, n32202, n32206, n32641, n32204,
    n32203, n32205, n32207, n32209, n32219, n32217, n32656, n32215, n32214,
    n32216, n32218, n32220, n32229, n32225, n32226, n32244, n32242, n32240,
    n32234, n32238, n32235, n32237, n32239, n32241, n32243, n32247, n32253,
    n32251, n32679, n32249, n32250, n32252, n32255, n32273, n32258, n32260,
    n32269, n32264, n32267, n32695, n32265, n32266, n32268, n32270, n32276,
    n32274, n32704, n32275, n32289, n32278, n32708, n32287, n32285, n32283,
    n32714, n32281, n32282, n32284, n32286, n32288, n32290, n32304, n32293,
    n32302, n32300, n32295, n32298, n32737, n32296, n32297, n32299, n32301,
    n32303, n32320, n32308, n32751, n32318, n32316, n32314, n32754, n32312,
    n32311, n32313, n32315, n32317, n32319, n32330, n32328, n32322, n32326,
    n32323, n32325, n32327, n32329, n32331, n32341, n32339, n32337, n32334,
    n32336, n32338, n32340, n32342, n32347, n32354, n32349, n32352, n32766,
    n32350, n32351, n32353, n32355, n32357, n32371, n32367, n32365, n32786,
    n32363, n32364, n32366, n32368, n32370, n32375, n32798, n32388, n32378,
    n32377, n32386, n32384, n32379, n32382, n32811, n32380, n32381, n32383,
    n32385, n32387, n32827, n32400, n39704, n32396, n32394, n32821, n32392,
    n32393, n32395, n32397, n32399, n32417, n39713, n32413, n32838, n32408,
    n32407, n32411, n32409, n32410, n32412, n32414, n32416, n32419, n32430,
    n39721, n32428, n32866, n32424, n32423, n32426, n32425, n32427, n32429,
    n32435, n32434, n32439, n32879, n32449, n39732, n32447, n32882, n32442,
    n32445, n32443, n32444, n32446, n32448, n32451, n32894, n32450, n32453,
    n32897, n32467, n32456, n32465, n39741, n32463, n32905, n32459, n32461,
    n32460, n32462, n32464, n32466, n32480, n39751, n32478, n32936, n32473,
    n32476, n32474, n32475, n32477, n32479, n32485, n32504, n32483, n32944,
    n32484, n32491, n32489, n32490, n32947, n32501, n39759, n32499, n32954,
    n32495, n32494, n32497, n32496, n32498, n32500, n32507, n32503, n32505,
    n32964, n32506, n32967, n32523, n32510, n32968, n32521, n39492, n32519,
    n32514, n32513, n32517, n32515, n32516, n32518, n32520, n32522, n32546,
    n32528, n32548, n32547, n32531, n32535, n32534, n32990, n32544, n39496,
    n32540, n33008, n32538, n32539, n32542, n32541, n32543, n32545, n33022,
    n32558, n39787, n32556, n33030, n32551, n32554, n32552, n32553, n32555,
    n32557, n32561, n33039, n32560, n33042, n32572, n39543, n39794, n32570,
    n33048, n32566, n32565, n32568, n32567, n32569, n32571, n32580, n32596,
    n32576, n32578, n33057, n32579, n32582, n32584, n33060, n32595, n39802,
    n32593, n33077, n32588, n32587, n32591, n32589, n32590, n32592, n32594,
    n32599, n33087, n32598, n32600, n33092, n32610, n32601, n32603, n40286,
    n40285, n33098, n32606, n33099, n32605, n32608, n32607, n32609, n32612,
    n32611, n32631, n32629, n32624, n32622, n32620, n32621, n32623, n32627,
    n32626, n32628, n32630, n32647, n32636, n32652, n32644, n32639, n32640,
    n32642, n32643, n32645, n32648, n32663, n32661, n32659, n32654, n32657,
    n32658, n32660, n32662, n32664, n32667, n32685, n32683, n32692, n32670,
    n32681, n32672, n32675, n32674, n32676, n32711, n32677, n32691, n32678,
    n32680, n32682, n32684, n32686, n32689, n32698, n32694, n32693, n32696,
    n32697, n32701, n32700, n32702, n32706, n32705, n32725, n32723, n32721,
    n32719, n32717, n32715, n32716, n32718, n32720, n32722, n32724, n32749,
    n32747, n32729, n32742, n32730, n32756, n32731, n32753, n32733, n32740,
    n32735, n32738, n32739, n32741, n32745, n32744, n32746, n32748, n32763,
    n32761, n32759, n32755, n32757, n32758, n32760, n32762, n32764, n32767,
    n32769, n32768, n32776, n32774, n32773, n32775, n32777, n32779, n32797,
    n32783, n32795, n32790, n32788, n32785, n32787, n32789, n32793, n32792,
    n32794, n32796, n32816, n32801, n32802, n32832, n40412, n32804, n32805,
    n32810, n32806, n32812, n32814, n32813, n32815, n32820, n32822, n32825,
    n39351, n32824, n32826, n32828, n32847, n32834, n32833, n32843, n32841,
    n32836, n39846, n32839, n32840, n32842, n32844, n32846, n32875, n32850,
    n32889, n32854, n32918, n32853, n32855, n32900, n32856, n32909, n32880,
    n32857, n32873, n32860, n32871, n32869, n32865, n32864, n39855, n32867,
    n32868, n32870, n32872, n32874, n32878, n32877, n32893, n32881, n32891,
    n32887, n32884, n39405, n32886, n32888, n32890, n32892, n32896, n32895,
    n32916, n32914, n32912, n32901, n32908, n32903, n39429, n32906, n32907,
    n32910, n32911, n32913, n32915, n32943, n32919, n32920, n32976, n32922,
    n32948, n32924, n32923, n32949, n32929, n32926, n32928, n32941, n32930,
    n32939, n32935, n32934, n39870, n32937, n32938, n32940, n32942, n32946,
    n32945, n32963, n32961, n32959, n32957, n32953, n32952, n39876, n32955,
    n32956, n32958, n32960, n32962, n32966, n32965, n32988, n32986, n32984,
    n32982, n32972, n39881, n32980, n32978, n32977, n32979, n32981, n32983,
    n32985, n32987, n33021, n33019, n32992, n32994, n32998, n32997, n33043,
    n32999, n33024, n40389, n33000, n33001, n33105, n33044, n33004, n33029,
    n33005, n33013, n33011, n33007, n39497, n33009, n33010, n33012, n33017,
    n33014, n33016, n33018, n33020, n33038, n33036, n33034, n33028, n39893,
    n33032, n33031, n33033, n33035, n33037, n33041, n33040, n33056, n33054,
    n33052, n33050, n39899, n33047, n33049, n33051, n33053, n33055, n33059,
    n33058, n33085, n33063, n40384, n33067, n40388, n40378, n33066, n33090,
    n33068, n40367, n33069, n40360, n33070, n33083, n33071, n33081, n39558,
    n33079, n33075, n33076, n33078, n33080, n33082, n33084, n33089, n33088,
    n33091, n33097, n33095, n42147, n33096, n33103, n33101, n33100, n33102,
    n33109, n33107, n33106, n33108, n33110, n40341, n33120, n33114, n39963,
    n33118, n40347, n33117, n33119, n33122, n33121, n33130, n33128, n33126,
    n40346, n33127, n33129, n41884, n33132, n33134, n33258, n33252, n33138,
    n33139, n33142, n33183, n33157, n33148, n33149, n33152, n33160, n33150,
    n33161, n33151, n33155, n33153, n33154, n33156, n42086, n33159, n33158,
    n33201, n33175, n33173, n33163, n33171, n33169, n33212, n33166, n33167,
    n33168, n33170, n33172, n42102, n33174, n33196, n33211, n33182, n33177,
    n33180, n33178, n33179, n33181, n42116, n33190, n33188, n33187, n33189,
    n42125, n33192, n33191, n33195, n33193, n33194, n33198, n33197, n33200,
    n33199, n33203, n33202, n33207, n33205, n33206, n33209, n33208, n33210,
    n33248, n33214, n33215, n33216, n42082, n33219, n33227, n33225, n33222,
    n33224, n33226, n33235, n33233, n33232, n33234, n42192, n33238, n33241,
    n39161, n33242, n33243, n33244, n33246, n33247, n33254, n33249, n33250,
    n33251, n41890, n33253, n33256, n33255, n33257, n33263, n33259, n33261,
    n41885, n33260, n33262, n33264, n33266, n33269, n33275, n39046, n33363,
    n33274, n33272, n33270, n33271, n33273, n33281, n33277, n33278, n33280,
    n33283, n33282, n38668, n33348, n36229, n34343, n36686, n33285, n36639,
    n33286, n36537, n33820, n33822, n33287, n36405, n33811, n36205, n33803,
    n33288, n36751, n33729, n39104, n33289, n36112, n33794, n33303, n33292,
    n37441, n39038, n33290, n37436, n38115, n34460, n36478, n36262, n33291,
    n36484, n33299, n33315, n33298, n33376, n33293, n33369, n33296, n36691,
    n33372, n33295, n33297, n33343, n33300, n33301, n33347, n36390, n33349,
    n33317, n33302, n33330, n33309, n33308, n33339, n33310, n33328, n33312,
    n33311, n36220, n36172, n36142, n33314, n33326, n33316, n33321, n33318,
    n33320, n33324, n33863, n33323, n33325, n33327, n33329, n33334, n33332,
    n33333, n33335, n33402, n33361, n33336, n33337, n33359, n33341, n33340,
    n33357, n33344, n33345, n33346, n33355, n33880, n33350, n33353, n33351,
    n33400, n33352, n33354, n33356, n33358, n33360, n33368, n37300, n33364,
    n33366, n33367, n33371, n33370, n33374, n33373, n33375, n33379, n33377,
    n33378, n33380, n33390, n36780, n33383, n33385, n33387, n33389, n33391,
    n33392, n33398, n33394, n33396, n33397, n33401, n37165, n33403, n36132,
    n33405, n33404, n36135, n33407, n33425, n33409, n33422, n33411, n33410,
    n36987, n33416, n33415, n33414, n36808, n33418, n33420, n33421, n33423,
    n33424, n33445, n33427, n33441, n33431, n33430, n33439, n36892, n33437,
    n33435, n33434, n33436, n33438, n33440, n33442, n33443, n33444, n33450,
    n33446, n33448, n33447, n36122, n33449, n33457, n33651, n33451, n33452,
    n33454, n33453, n33455, n33456, n33459, n33656, n33458, n33462, n33461,
    n33464, n40532, n33463, n33466, n33465, n33468, n40514, n33467, n33470,
    n33469, n33472, n40498, n33471, n33474, n33473, n33476, n40483, n33475,
    n33478, n33477, n33480, n40468, n33479, n33482, n33481, n33484, n40453,
    n33483, n33486, n33485, n33489, n40445, n33488, n33491, n33490, n33493,
    n33492, n33495, n33494, n33497, n33496, n33499, n33498, n33501, n33500,
    n33503, n33502, n33505, n33504, n33507, n33506, n33509, n33508, n33511,
    n33510, n33513, n33512, n33515, n33514, n33517, n33516, n33519, n33518,
    n33521, n33520, n33523, n33522, n40040, n33525, n33524, n33527, n33526,
    n40045, n33529, n33528, n33531, n33530, n40050, n33533, n33532, n33535,
    n33534, n40055, n33537, n33536, n33540, n33539, n40060, n33542, n33541,
    n33544, n33543, n40065, n33546, n33545, n33548, n33547, n40070, n33550,
    n33549, n33552, n33551, n40075, n33554, n33553, n33556, n33555, n33558,
    n33557, n33560, n33559, n33562, n33561, n33564, n33563, n33566, n33565,
    n33568, n33567, n33570, n33569, n33572, n33571, n33574, n33573, n33576,
    n33575, n33578, n33577, n33580, n33579, n33582, n33581, n33584, n33583,
    n33587, n33586, n33590, n33589, n33592, n33591, n33594, n33593, n33596,
    n33595, n33598, n33597, n33600, n33599, n33602, n33601, n33604, n33603,
    n33606, n33605, n33608, n33607, n33610, n33609, n33612, n33611, n33614,
    n33613, n33616, n33615, n33618, n33617, n33620, n33619, n33622, n33621,
    n33624, n33623, n33626, n33625, n33628, n33627, n33630, n33629, n33632,
    n33631, n33634, n33633, n33636, n33635, n33638, n33637, n33640, n33639,
    n33642, n33641, n33644, n33643, n33646, n33645, n33648, n33647, n33650,
    n33649, n33653, n33652, n33655, n33654, n33658, n33657, n33661, n33700,
    n33719, n33663, n33662, n33665, n33664, n33667, n33666, n33669, n33668,
    n33671, n33670, n33673, n33672, n33675, n33674, n33677, n33676, n33679,
    n33678, n33681, n33680, n33683, n33682, n33685, n33684, n33687, n33686,
    n33689, n33688, n33691, n33690, n33693, n33692, n33695, n33694, n33697,
    n33696, n33699, n33698, n33702, n33701, n33704, n33703, n33706, n33705,
    n33708, n33707, n33710, n33709, n33712, n33711, n33714, n33713, n33716,
    n33715, n33718, n33717, n33721, n33720, n33724, n33723, n33727, n38860,
    n33725, n33726, n39019, n33728, n39130, n33732, n33730, n33731, n33733,
    n33734, n33736, n33735, n33738, n39023, n33739, n38804, n33789, n33741,
    n33743, n33745, n33744, n33746, n38670, n39101, n33748, n33751, n33750,
    n33755, n33753, n33752, n33754, n33779, n33757, n33756, n33759, n33758,
    n33761, n33760, n33777, n33763, n33762, n33767, n33765, n33764, n33766,
    n33775, n33769, n33768, n33773, n33771, n33770, n33772, n33774, n33776,
    n33778, n39092, n33783, n39083, n39082, n33780, n33784, n33781, n33782,
    n33787, n39081, n33785, n33786, n39006, n33847, n34005, n38950, n38940,
    n38930, n38920, n38910, n38900, n38880, n39084, n33790, n34369, n34349,
    n34325, n34305, n34285, n34243, n34231, n34219, n34191, n34173, n34145,
    n34127, n34112, n34090, n34077, n34058, n34004, n33791, n33945, n33892,
    n33894, n33792, n33915, n33793, n33872, n33797, n33840, n33865, n33795,
    n38818, n38808, n33798, n33869, n33799, n33846, n33806, n33800, n36106,
    n33907, n36147, n36184, n33810, n36111, n33804, n33805, n36148, n33833,
    n33807, n33808, n36180, n33832, n36209, n33814, n36239, n33809, n36234,
    n36272, n33819, n36345, n36263, n33812, n33813, n36291, n36311, n33827,
    n36364, n33815, n33816, n36342, n33825, n33817, n33818, n36391, n36447,
    n36455, n33821, n34298, n36477, n34179, n36410, n36747, n34138, n34107,
    n36412, n33823, n33824, n36404, n34086, n34071, n36363, n34051, n33826,
    n34030, n33828, n33829, n33956, n33834, n33906, n33835, n34463, n34421,
    n33844, n33850, n33836, n34445, n33838, n33837, n33842, n33839, n33841,
    n33843, n33845, n33853, n34484, n34401, n34389, n34486, n34352, n34317,
    n34304, n34276, n34279, n34251, n34227, n34217, n34189, n34167, n34154,
    n35190, n34128, n35121, n34093, n34074, n34047, n34035, n34493, n34021,
    n34893, n33980, n33963, n34494, n33948, n33930, n34806, n33912, n33900,
    n33899, n33898, n33854, n33849, n33851, n33852, n34507, n33855, n33857,
    n33856, n33861, n33859, n33858, n33860, n33868, n33864, n33866, n33867,
    n33871, n33870, n33875, n33873, n33874, n33885, n33878, n33876, n33877,
    n33883, n33881, n33882, n33884, n33886, n33940, n33917, n33887, n33891,
    n33889, n33888, n33890, n33897, n33986, n33953, n33893, n33895, n33896,
    n33904, n33902, n33901, n33903, n33911, n33909, n33908, n33910, n34827,
    n33913, n33925, n33914, n33921, n33916, n33919, n33918, n33920, n33923,
    n33922, n33924, n33927, n33926, n33928, n33939, n33929, n33935, n33931,
    n33933, n33932, n33934, n33937, n33936, n33938, n33942, n33941, n33965,
    n33944, n33943, n33961, n33970, n33946, n33987, n33972, n33947, n38981,
    n33952, n34805, n33949, n33950, n33951, n33955, n33954, n33959, n33957,
    n33958, n33960, n33962, n33976, n33964, n33969, n33967, n33966, n33968,
    n33974, n33971, n33973, n33975, n33978, n33977, n33979, n33985, n34804,
    n33981, n33983, n33982, n33984, n33993, n33991, n33989, n33988, n33990,
    n33992, n33995, n33994, n33998, n33997, n34012, n34014, n33999, n34044,
    n38960, n34013, n34000, n34001, n38965, n34010, n34003, n34008, n34034,
    n34006, n34007, n34009, n34011, n34020, n34037, n34016, n34015, n34018,
    n34017, n34019, n34029, n34803, n34022, n34023, n34027, n34025, n34026,
    n34028, n34031, n34043, n34033, n34032, n34041, n34039, n34036, n34038,
    n34040, n34042, n34046, n34045, n34050, n34048, n34049, n34055, n34052,
    n34053, n34054, n34065, n34076, n34089, n34102, n34056, n34063, n34057,
    n34059, n34061, n34060, n34062, n34064, n34067, n34066, n34069, n34068,
    n34070, n34083, n34072, n34073, n34081, n34075, n34079, n34078, n34080,
    n34082, n35078, n34084, n34085, n34101, n34087, n34088, n34097, n34091,
    n34095, n34092, n34094, n34096, n34099, n34098, n34100, n34104, n34103,
    n34126, n34105, n34147, n34106, n34125, n34108, n34109, n34123, n34110,
    n34111, n34121, n34113, n34115, n34114, n34118, n34130, n34117, n34119,
    n34120, n34122, n34124, n34137, n34129, n34135, n34132, n34131, n34133,
    n34134, n34136, n34144, n34142, n36444, n34139, n34140, n34141, n34143,
    n34146, n38925, n34149, n34148, n34153, n34150, n34151, n34152, n34158,
    n34156, n34169, n34155, n34157, n34164, n36459, n34159, n34160, n34161,
    n34162, n34163, n38915, n34193, n34165, n34222, n34166, n34188, n34168,
    n34171, n34170, n34186, n34172, n34175, n34174, n34184, n34177, n34176,
    n34180, n34178, n36476, n34181, n34182, n34183, n34185, n34187, n34200,
    n34190, n34195, n34192, n34194, n34198, n34196, n34197, n34199, n34207,
    n34205, n36507, n34201, n34202, n34203, n34204, n34206, n34208, n34210,
    n34209, n34216, n34235, n34211, n36535, n34212, n34213, n34214, n34215,
    n34226, n35279, n34218, n34224, n34220, n34221, n34223, n34225, n34230,
    n34228, n34229, n34248, n34232, n34233, n34242, n36581, n34240, n34252,
    n34236, n34234, n36565, n34237, n34254, n34238, n34239, n34241, n34246,
    n38905, n34266, n34265, n34286, n34244, n34245, n34247, n35346, n34249,
    n34250, n34270, n34278, n34264, n36596, n34253, n34259, n34422, n34273,
    n34256, n34255, n34257, n34258, n34262, n34260, n34261, n34263, n34268,
    n34267, n34269, n34272, n34271, n36615, n34274, n34275, n34290, n34277,
    n34284, n34280, n34282, n34281, n34283, n34288, n34287, n34289, n34293,
    n34292, n35439, n34294, n34295, n34302, n34412, n34342, n34321, n34296,
    n34297, n36633, n34374, n34299, n34331, n34300, n34301, n34316, n34326,
    n34348, n34361, n34303, n34314, n34319, n34308, n34306, n34307, n34312,
    n34310, n34311, n34313, n34315, n34318, n34339, n34324, n36654, n36649,
    n34461, n34322, n34323, n34335, n34328, n34327, n34329, n34333, n34330,
    n34332, n34334, n34337, n34336, n34338, n34341, n34340, n36670, n34344,
    n34372, n34345, n34360, n35455, n34346, n34347, n34356, n34350, n34354,
    n34351, n34353, n34355, n34358, n34357, n34359, n34363, n34362, n35815,
    n39136, n37389, n34364, n34368, n34365, n34366, n34367, n34388, n38875,
    n34370, n34404, n34383, n36692, n34373, n34379, n34375, n34377, n34378,
    n34381, n34403, n34380, n34382, n34386, n34385, n34387, n34393, n34390,
    n34391, n34392, n36699, n34400, n38742, n38736, n39039, n34398, n34397,
    n34399, n34419, n34402, n34410, n38870, n34408, n34429, n34406, n34407,
    n34409, n34417, n36717, n34413, n34411, n36703, n34420, n34414, n34415,
    n34416, n34418, n34424, n36720, n34423, n34428, n34426, n34427, n34444,
    n38865, n34433, n34455, n34431, n34432, n34442, n34474, n39047, n34435,
    n34434, n34440, n34438, n34436, n34437, n34439, n34441, n34443, n34450,
    n35472, n34446, n35482, n34449, n34458, n34452, n39057, n34454, n34453,
    n34456, n34457, n34467, n34465, n34462, n34464, n34466, n34473, n34471,
    n34472, n34476, n34475, n34480, n39073, n34477, n34479, n34482, n35192,
    n35460, n34485, n35446, n34487, n35441, n34488, n35345, n35119, n35348,
    n34489, n35272, n35200, n34490, n35113, n35046, n35009, n34491, n34802,
    n34933, n34496, n34495, n34500, n34812, n34497, n34498, n34499, n34501,
    n34508, n34504, n34502, n34506, n34503, n34505, n34509, n34801, n34511,
    n34510, n34515, n34513, n34512, n34514, n34524, n34518, n34517, n34522,
    n34520, n34519, n34521, n34523, n34542, n34527, n34526, n34531, n34529,
    n34528, n34530, n34540, n34534, n34533, n34538, n34536, n34535, n34537,
    n34539, n34541, n34799, n34544, n34543, n34549, n34547, n34546, n34548,
    n34557, n34551, n34550, n34555, n34553, n34552, n34554, n34556, n34574,
    n34559, n34558, n34563, n34561, n34560, n34562, n34572, n34566, n34565,
    n34570, n34568, n34567, n34569, n34571, n34573, n34819, n34577, n34576,
    n34582, n34580, n34579, n34581, n34591, n34584, n34583, n34589, n34587,
    n35359, n34586, n34588, n34590, n34607, n34593, n34592, n34597, n34595,
    n34594, n34596, n34605, n34599, n34598, n34603, n34601, n34600, n34602,
    n34604, n34606, n34834, n34609, n34608, n34614, n34612, n34611, n34613,
    n34622, n34616, n34615, n34620, n35366, n34618, n34617, n34619, n34621,
    n34639, n34624, n34623, n34628, n34626, n34625, n34627, n34637, n34630,
    n34629, n34635, n34633, n34632, n34634, n34636, n34638, n34848, n34641,
    n34640, n34645, n34643, n34642, n34644, n34670, n34647, n34646, n34651,
    n34649, n34648, n34650, n34668, n34653, n34652, n34657, n34655, n34654,
    n34656, n34666, n34659, n34658, n34664, n34662, n34661, n34663, n34665,
    n34667, n34669, n34856, n34672, n34671, n34676, n34674, n34673, n34675,
    n34700, n34678, n34677, n34682, n34680, n34679, n34681, n34698, n34684,
    n34683, n34688, n34686, n34685, n34687, n34696, n34690, n34689, n34694,
    n34692, n34691, n34693, n34695, n34697, n34699, n34855, n34847, n34841,
    n34702, n34701, n34706, n34704, n34703, n34705, n34731, n34708, n34707,
    n34729, n34710, n34709, n34714, n34712, n34711, n34713, n34727, n34716,
    n34715, n34721, n34719, n34718, n34720, n34725, n34723, n34722, n34724,
    n34726, n34728, n34730, n34840, n34833, n34826, n34733, n34732, n34737,
    n34735, n34734, n34736, n34761, n34739, n34738, n34759, n34741, n34740,
    n34745, n34743, n34742, n34744, n34757, n34747, n34746, n34751, n34749,
    n34748, n34750, n34755, n34753, n34752, n34754, n34756, n34758, n34760,
    n34825, n34818, n34809, n34763, n34762, n34767, n34765, n34764, n34766,
    n34797, n34769, n34768, n34795, n34771, n34770, n34775, n34773, n34772,
    n34774, n34793, n34776, n34781, n34780, n34787, n37505, n34785, n34784,
    n34786, n34791, n34789, n34788, n34790, n34792, n34794, n34796, n34808,
    n34798, n35511, n34800, n34966, n34900, n34895, n34897, n34849, n34851,
    n34816, n34836, n34807, n34811, n35520, n34810, n34815, n34828, n35486,
    n35483, n34813, n34822, n34814, n34817, n34821, n35530, n34820, n34824,
    n34823, n35541, n34832, n34830, n34829, n34831, n35551, n34839, n34835,
    n34837, n34838, n35564, n34846, n34842, n34844, n34845, n35578, n34854,
    n34850, n34858, n34852, n34853, n35585, n34861, n34857, n34859, n34860,
    n34863, n34862, n34867, n34865, n34864, n34866, n34892, n34869, n34868,
    n34890, n34871, n34870, n34876, n34874, n34873, n34875, n34888, n34878,
    n34877, n34882, n34880, n34879, n34881, n34886, n34884, n34883, n34885,
    n34887, n34889, n34891, n35592, n34899, n34894, n34896, n34898, n34932,
    n34902, n34901, n34906, n34904, n34903, n34905, n34914, n34908, n34907,
    n34912, n34910, n34909, n34911, n34913, n34930, n34916, n34915, n34920,
    n34918, n34917, n34919, n34928, n34922, n34921, n34926, n34924, n34923,
    n34925, n34927, n34929, n35607, n34931, n34935, n34968, n34934, n34937,
    n34936, n34941, n34939, n34938, n34940, n34949, n34943, n34942, n34947,
    n34945, n34944, n34946, n34948, n34965, n34951, n34950, n34955, n34953,
    n34952, n34954, n34963, n34957, n34956, n34961, n34959, n34958, n34960,
    n34962, n34964, n35619, n34970, n34967, n34969, n34972, n35005, n34974,
    n34973, n34978, n34976, n34975, n34977, n34986, n34980, n34979, n34984,
    n34982, n34981, n34983, n34985, n35003, n34988, n34987, n34992, n34990,
    n34989, n34991, n35001, n34995, n34994, n34999, n34997, n34996, n34998,
    n35000, n35002, n35629, n35004, n35008, n35043, n35007, n35010, n35042,
    n35012, n35011, n35016, n35014, n35013, n35015, n35024, n35018, n35017,
    n35022, n35020, n35019, n35021, n35023, n35040, n35026, n35025, n35030,
    n35028, n35027, n35029, n35038, n35032, n35031, n35036, n35034, n35033,
    n35035, n35037, n35039, n35640, n35041, n35045, n35044, n35047, n35082,
    n35049, n35048, n35053, n35051, n35050, n35052, n35061, n35055, n35054,
    n35059, n35057, n35056, n35058, n35060, n35077, n35063, n35062, n35067,
    n35065, n35064, n35066, n35075, n35069, n35068, n35073, n35071, n35070,
    n35072, n35074, n35076, n35651, n35080, n35079, n35081, n35084, n35083,
    n35088, n35086, n35085, n35087, n35096, n35090, n35089, n35094, n35092,
    n35091, n35093, n35095, n35112, n35098, n35097, n35102, n35100, n35099,
    n35101, n35110, n35104, n35103, n35108, n35106, n35105, n35107, n35109,
    n35111, n35664, n35118, n35116, n35114, n35115, n35117, n35124, n35357,
    n35278, n35120, n35189, n35155, n35122, n35123, n35126, n35125, n35130,
    n35128, n35127, n35129, n35154, n35132, n35131, n35152, n35134, n35133,
    n35138, n35136, n35135, n35137, n35150, n35140, n35139, n35144, n35142,
    n35141, n35143, n35148, n35146, n35145, n35147, n35149, n35151, n35153,
    n35672, n35158, n35156, n35157, n35160, n35159, n35164, n35162, n35161,
    n35163, n35188, n35168, n35166, n35165, n35167, n35170, n35169, n35186,
    n35172, n35171, n35176, n35174, n35173, n35175, n35184, n35178, n35177,
    n35182, n35180, n35179, n35181, n35183, n35185, n35187, n35682, n35198,
    n35201, n35196, n35191, n35193, n35194, n35195, n35197, n35199, n35236,
    n35202, n35234, n35204, n35203, n35208, n35206, n35205, n35207, n35216,
    n35210, n35209, n35214, n35212, n35211, n35213, n35215, n35232, n35218,
    n35217, n35222, n35220, n35219, n35221, n35230, n35224, n35223, n35228,
    n35226, n35225, n35227, n35229, n35231, n35694, n35233, n35235, n35237,
    n35270, n35239, n35238, n35243, n35241, n35240, n35242, n35251, n35245,
    n35244, n35249, n35247, n35246, n35248, n35250, n35268, n35254, n35253,
    n35258, n35256, n35255, n35257, n35266, n35260, n35259, n35264, n35262,
    n35261, n35263, n35265, n35267, n35699, n35269, n35277, n35271, n35275,
    n35274, n35276, n35280, n35312, n35282, n35281, n35286, n35284, n35283,
    n35285, n35294, n35288, n35287, n35292, n35290, n35289, n35291, n35293,
    n35310, n35296, n35295, n35300, n35298, n35297, n35299, n35308, n35302,
    n35301, n35306, n35304, n35303, n35305, n35307, n35309, n35708, n35311,
    n35314, n35313, n35318, n35316, n35315, n35317, n35327, n35321, n35320,
    n35325, n35323, n35322, n35324, n35326, n35344, n35330, n35329, n35334,
    n35332, n35331, n35333, n35342, n35336, n35335, n35340, n35338, n35337,
    n35339, n35341, n35343, n35717, n35352, n35347, n35350, n35349, n35351,
    n35356, n35354, n35355, n35358, n35393, n35361, n35360, n35365, n35363,
    n35362, n35364, n35374, n35368, n35367, n35372, n35370, n35369, n35371,
    n35373, n35390, n35376, n35375, n35380, n35378, n35377, n35379, n35388,
    n35382, n35381, n35386, n35384, n35383, n35385, n35387, n35389, n35723,
    n35392, n35454, n35451, n35437, n35434, n35395, n35432, n35398, n35397,
    n35402, n35400, n35399, n35401, n35411, n35404, n35403, n35409, n35407,
    n35406, n35408, n35410, n35430, n35414, n35413, n35419, n35417, n35416,
    n35418, n35428, n35421, n35420, n35426, n35424, n35423, n35425, n35427,
    n35429, n35733, n35431, n35436, n35433, n35435, n35438, n35443, n35440,
    n35442, n35445, n35444, n35462, n35448, n35450, n35449, n35453, n35457,
    n35452, n35459, n35456, n35458, n35465, n35461, n35466, n35475, n35468,
    n35463, n35464, n35471, n35467, n35469, n35470, n35473, n35474, n35476,
    n35479, n35478, n35481, n37456, n35480, n35485, n35484, n35489, n37446,
    n35488, n35492, n35491, n36013, n36003, n35994, n36098, n35688, n35493,
    n35495, n35494, n35497, n35741, n35742, n35496, n35744, n35687, n35498,
    n35596, n35597, n35975, n35964, n35499, n35595, n35500, n35501, n35502,
    n35571, n35537, n35503, n35506, n40548, n35505, n35510, n36018, n35507,
    n35508, n35509, n35513, n35512, n35516, n35515, n35517, n35660, n35518,
    n35526, n35522, n35521, n35524, n35523, n35525, n35529, n35527, n35528,
    n35532, n35531, n35534, n35533, n35540, n35536, n35547, n35538, n35539,
    n35543, n35542, n35545, n35544, n35550, n35546, n35548, n35549, n35553,
    n35552, n35556, n35555, n35561, n35557, n35559, n35560, n35563, n35562,
    n35566, n35565, n35570, n35567, n35568, n35569, n35573, n35572, n35575,
    n35582, n35577, n35576, n35580, n35579, n35581, n35985, n35584, n35589,
    n35587, n35586, n35588, n35591, n35590, n35594, n35593, n35604, n35598,
    n35643, n35654, n35602, n35970, n35634, n35612, n35599, n35600, n35601,
    n35603, n35606, n35605, n35611, n35609, n35608, n35610, n35616, n35614,
    n35613, n35615, n35618, n35617, n35621, n35620, n35626, n35622, n35624,
    n35625, n35628, n35627, n35631, n35630, n35637, n35633, n35645, n35635,
    n35636, n35639, n35638, n35642, n35641, n35648, n35644, n35656, n35646,
    n35647, n35650, n35649, n35653, n35652, n35659, n35655, n35657, n35658,
    n35663, n35662, n35666, n35665, n35670, n35947, n35668, n35669, n35681,
    n35676, n35674, n35673, n35675, n35680, n35678, n35679, n36092, n35686,
    n35684, n35683, n35685, n35690, n36072, n35724, n35710, n35700, n35693,
    n35689, n36082, n35703, n36087, n35691, n35692, n35696, n35695, n35698,
    n35697, n35705, n35712, n35701, n35702, n35704, n35707, n35706, n35714,
    n36077, n35709, n35711, n35713, n35716, n35715, n35720, n35718, n35719,
    n35722, n35721, n35730, n35728, n36067, n35725, n35727, n35729, n35732,
    n35731, n35738, n35734, n35736, n35735, n35737, n35740, n35739, n35749,
    n36037, n35791, n35778, n35781, n35762, n35756, n36057, n35743, n35747,
    n35746, n35748, n35751, n35750, n35758, n36047, n35765, n36052, n35754,
    n35755, n35757, n35760, n35759, n35767, n35772, n35763, n35764, n35766,
    n35769, n35768, n36042, n35770, n35771, n35775, n35774, n35777, n35776,
    n35793, n35779, n35780, n35786, n35783, n35785, n35788, n35787, n36032,
    n35790, n35792, n35796, n35795, n35798, n35797, n35803, n36027, n35801,
    n35802, n35806, n35805, n35809, n35808, n35936, n35814, n35813, n35817,
    n35816, n35819, n35818, n35821, n35820, n35823, n35822, n35825, n35824,
    n35827, n35826, n35829, n35828, n35831, n35830, n35833, n35832, n35835,
    n35834, n35837, n35836, n35839, n35838, n35841, n35840, n35843, n35842,
    n35845, n35844, n35847, n35846, n35849, n35848, n35851, n35850, n35853,
    n35852, n35855, n35854, n35857, n35856, n35859, n35858, n35861, n35860,
    n35863, n35862, n35865, n35864, n35867, n35866, n35869, n35868, n35871,
    n35870, n35874, n35873, n35876, n35875, n35878, n35877, n35880, n35879,
    n35882, n35881, n35884, n35883, n35886, n35885, n35888, n35887, n35890,
    n35889, n35892, n35891, n35894, n35893, n35896, n35895, n35898, n35897,
    n35900, n35899, n35902, n35901, n35904, n35903, n35906, n35905, n35908,
    n35907, n35911, n35910, n35913, n35912, n35915, n35914, n35917, n35916,
    n35919, n35918, n35921, n35920, n35923, n35922, n35925, n35924, n35927,
    n35926, n35929, n35928, n35931, n35930, n35933, n35932, n35935, n35934,
    n35939, n35938, n35942, n35941, n35946, n36103, n35952, n36097, n35950,
    n35949, n36023, n35951, n35953, n36028, n35954, n35955, n35957, n35956,
    n35958, n36033, n35959, n35960, n35962, n35961, n35963, n36038, n35965,
    n35968, n35967, n35969, n36043, n35971, n35973, n35972, n35974, n36048,
    n35976, n35978, n35977, n35979, n36053, n35980, n35981, n35983, n35982,
    n35984, n36058, n35986, n35988, n35987, n35989, n36063, n35990, n35992,
    n35991, n35993, n36068, n35995, n35997, n35996, n35998, n36073, n35999,
    n36001, n36000, n36002, n36078, n36004, n36006, n36005, n36007, n36083,
    n36008, n36009, n36011, n36010, n36012, n36088, n36014, n36016, n36015,
    n36017, n36093, n36019, n36021, n36020, n36022, n36024, n36026, n36025,
    n36029, n36031, n36030, n36034, n36036, n36035, n36039, n36041, n36040,
    n36044, n36046, n36045, n36049, n36051, n36050, n36054, n36056, n36055,
    n36059, n36061, n36060, n36064, n36066, n36065, n36069, n36071, n36070,
    n36074, n36076, n36075, n36079, n36081, n36080, n36084, n36086, n36085,
    n36089, n36091, n36090, n36094, n36096, n36095, n36102, n36100, n36101,
    n36105, n36104, n36121, n36108, n36119, n36110, n36145, n36162, n36116,
    n37401, n38823, n36114, n36115, n36168, n36146, n36117, n36118, n36120,
    n36124, n36123, n36127, n36125, n36126, n36141, n36131, n36129, n36128,
    n36161, n36143, n36130, n36139, n36133, n36137, n36136, n36138, n36140,
    n36144, n36160, n36757, n36158, n36150, n36149, n36156, n36153, n36154,
    n36755, n36155, n36157, n36159, n36177, n36163, n36171, n36802, n36165,
    n36167, n36169, n36170, n36175, n36173, n36174, n36176, n36179, n36178,
    n36189, n36230, n36181, n36182, n36228, n36240, n36206, n36187, n36185,
    n36204, n36186, n36188, n36190, n36830, n36200, n36820, n36192, n36194,
    n36195, n36807, n36198, n36813, n36197, n36199, n36203, n36814, n36202,
    n36250, n36248, n36238, n36219, n36208, n36207, n36212, n36210, n36853,
    n36211, n36217, n36214, n36857, n36216, n36218, n36222, n36221, n36761,
    n36223, n36226, n36224, n36225, n36227, n36860, n36246, n38970, n36861,
    n36233, n36232, n36236, n36235, n36237, n36244, n36242, n36241, n36243,
    n36245, n36255, n36252, n36251, n36253, n36254, n37009, n36257, n36256,
    n36424, n36259, n36284, n36261, n36271, n36309, n36264, n36266, n36265,
    n36314, n36289, n36268, n36295, n36269, n36270, n36275, n36902, n36273,
    n36274, n36282, n36277, n36279, n36280, n36901, n36281, n36283, n36288,
    n36286, n36285, n36306, n36287, n36294, n36924, n36292, n36293, n36296,
    n36305, n36923, n36341, n36319, n36303, n36373, n36372, n36375, n36354,
    n36300, n36330, n36353, n36299, n36301, n36928, n36302, n36304, n36308,
    n36307, n36310, n36318, n36313, n36315, n36316, n36948, n36317, n36340,
    n36326, n36971, n36936, n36324, n36972, n36935, n36323, n36360, n36325,
    n36338, n36329, n36328, n36332, n36331, n36335, n36334, n36336, n36931,
    n36337, n36339, n36359, n36958, n36343, n36352, n36344, n36387, n36346,
    n36369, n36350, n36348, n36365, n36349, n36351, n36357, n36355, n36956,
    n36356, n36358, n36362, n36361, n36368, n36967, n36366, n36367, n36371,
    n36370, n36379, n36374, n36965, n36377, n36994, n36376, n36378, n36383,
    n36428, n36429, n36403, n36381, n36394, n36382, n37001, n36385, n36386,
    n36388, n36393, n36392, n36398, n36396, n37024, n37003, n36395, n36397,
    n36402, n37002, n36401, n36423, n36417, n36407, n36448, n36406, n36414,
    n36409, n36457, n36411, n36445, n36413, n36415, n37030, n36416, n36421,
    n36418, n37023, n36420, n36422, n36426, n36425, n37047, n36427, n37034,
    n36431, n36465, n37032, n36430, n36443, n36433, n36434, n36435, n36436,
    n36471, n36440, n36438, n36472, n36439, n36441, n37046, n36442, n36454,
    n36452, n36446, n37044, n36450, n36449, n36451, n36453, n36456, n36458,
    n36461, n36460, n36470, n37053, n36467, n36464, n37052, n36466, n36468,
    n37079, n36469, n36475, n36473, n37077, n36474, n36526, n37142, n37093,
    n36524, n36523, n36496, n36489, n36481, n36479, n36480, n36509, n36482,
    n37112, n36487, n36485, n36510, n36486, n36488, n36494, n37106, n36492,
    n36491, n36600, n36493, n36495, n36506, n36503, n36571, n36499, n36500,
    n36516, n37123, n36501, n36502, n36504, n37107, n36505, n36522, n36514,
    n37130, n36512, n36513, n36520, n36518, n36517, n37128, n36519, n36521,
    n36534, n36532, n36525, n36529, n36527, n36528, n36530, n36531, n36533,
    n36545, n37138, n36614, n36584, n36736, n36591, n36539, n36542, n36541,
    n36543, n36544, n36553, n36546, n36551, n36548, n36547, n36589, n36549,
    n36563, n36550, n36552, n36561, n36605, n36558, n36555, n36606, n36557,
    n36559, n37135, n36560, n37177, n36562, n37151, n36564, n36567, n36566,
    n36568, n36588, n36569, n36570, n36573, n37206, n36572, n36579, n37162,
    n36577, n36575, n36576, n36578, n37164, n36586, n36593, n36595, n36582,
    n36583, n36585, n36587, n36604, n36592, n36594, n36599, n37203, n36597,
    n36598, n36602, n36601, n36603, n36609, n36607, n37200, n36608, n36611,
    n37213, n36628, n36618, n37233, n36616, n36617, n36626, n37227, n36624,
    n36640, n36620, n36634, n36621, n36623, n36625, n36627, n36631, n36630,
    n37242, n36733, n36644, n36638, n37237, n36636, n36635, n36637, n36642,
    n36641, n36643, n36648, n36646, n37238, n36647, n37272, n36650, n36661,
    n37250, n36659, n36655, n36669, n36657, n36656, n36658, n36660, n36664,
    n37251, n36663, n36667, n36668, n36676, n36671, n37287, n36674, n37274,
    n36673, n36675, n36680, n37275, n36679, n37291, n37306, n36684, n36698,
    n36685, n36689, n36687, n36700, n36688, n36696, n36694, n36693, n36695,
    n36697, n36718, n36701, n36714, n37315, n36711, n37321, n36709, n37320,
    n36708, n36710, n36712, n36713, n37329, n36725, n36719, n36723, n36721,
    n37350, n36722, n36724, n36729, n36728, n36740, n37361, n36735, n37362,
    n36734, n36738, n36737, n36739, n36742, n37371, n36741, n36744, n36746,
    n36748, n37385, n36754, n37374, n36752, n36753, n36756, n36759, n36758,
    n36790, n36810, n36877, n36762, n36850, n36763, n36797, n36765, n36788,
    n36769, n36768, n36779, n36777, n36773, n36771, n36772, n36840, n36776,
    n36775, n36817, n36778, n36791, n36783, n36782, n36785, n36784, n36786,
    n36787, n36789, n36795, n36818, n36793, n36794, n36796, n36799, n36798,
    n36804, n36801, n36803, n36806, n36805, n36829, n36827, n36809, n36865,
    n36812, n36824, n36816, n36815, n36822, n36819, n36821, n36823, n36825,
    n36826, n36828, n36831, n36835, n36834, n36838, n36837, n36839, n36841,
    n36845, n36848, n36843, n36844, n36846, n36871, n36847, n36856, n36851,
    n36852, n36854, n36855, n36859, n36858, n36862, n36873, n36908, n36917,
    n36866, n36867, n36868, n36870, n36872, n36875, n36876, n36878, n36900,
    n36896, n36883, n36882, n36891, n36886, n36885, n36943, n36888, n36887,
    n36889, n36890, n36911, n36894, n36895, n36897, n36898, n36899, n36905,
    n36903, n36904, n36907, n36906, n36934, n36910, n36912, n36913, n36915,
    n36914, n36927, n37355, n36980, n37334, n36918, n36921, n36920, n36922,
    n36955, n36952, n36925, n36926, n36930, n36929, n36950, n37358, n36933,
    n36945, n36941, n36938, n36937, n36939, n36940, n36942, n36944, n36961,
    n36946, n36947, n36949, n36954, n36953, n36960, n36957, n36959, n36964,
    n36963, n36966, n36986, n37263, n37336, n36969, n36970, n36979, n36974,
    n36973, n36977, n36976, n36978, n36997, n36981, n36982, n36984, n36983,
    n36985, n36996, n36992, n36989, n36988, n37211, n37105, n37038, n36991,
    n36993, n37025, n36995, n36998, n36999, n37000, n37007, n37005, n37004,
    n37006, n37033, n37020, n37035, n37011, n37014, n37013, n37017, n37015,
    n37016, n37040, n37018, n37019, n37021, n37022, n37029, n37027, n37026,
    n37028, n37031, n37037, n37036, n37042, n37039, n37041, n37043, n37045,
    n37051, n37049, n37048, n37050, n37055, n37054, n37075, n37057, n37073,
    n37221, n37182, n37118, n37061, n37060, n37098, n37063, n37070, n37191,
    n37086, n37068, n37067, n37069, n37071, n37072, n37074, n37076, n37084,
    n37078, n37082, n37081, n37083, n37115, n37097, n37090, n37088, n37089,
    n37150, n37092, n37096, n37094, n37095, n37120, n37099, n37100, n37101,
    n37111, n37103, n37102, n37104, n37122, n37207, n37109, n37108, n37110,
    n37114, n37113, n37116, n37117, n37119, n37127, n37156, n37124, n37125,
    n37126, n37132, n37129, n37131, n37134, n37133, n37137, n37136, n37139,
    n37161, n37169, n37141, n37144, n37143, n37145, n37149, n37148, n37168,
    n37153, n37152, n37155, n37158, n37157, n37159, n37160, n37163, n37167,
    n37166, n37179, n37173, n37171, n37170, n37172, n37174, n37175, n37176,
    n37178, n37180, n37181, n37196, n37187, n37186, n37193, n37189, n37217,
    n37192, n37194, n37195, n37198, n37199, n37205, n37202, n37204, n37209,
    n37208, n37232, n37216, n37214, n37215, n37226, n37220, n37219, n37223,
    n37222, n37241, n37224, n37225, n37229, n37228, n37230, n37231, n37234,
    n37236, n37249, n37246, n37240, n37244, n37243, n37245, n37247, n37248,
    n37271, n37253, n37252, n37268, n37255, n37254, n37316, n37258, n37266,
    n37262, n37261, n37264, n37280, n37265, n37267, n37269, n37270, n37273,
    n37277, n37276, n37284, n37279, n37282, n37281, n37283, n37285, n37286,
    n37289, n37288, n37290, n37313, n37310, n37330, n37298, n37345, n37296,
    n37297, n37299, n37318, n37301, n37305, n37303, n37304, n37308, n37307,
    n37309, n37311, n37312, n37314, n37328, n37319, n37325, n37323, n37322,
    n37324, n37326, n37327, n37347, n37333, n37332, n37343, n37335, n37341,
    n37337, n37339, n37340, n37342, n37344, n37346, n37348, n37351, n37354,
    n37353, n37357, n37360, n37380, n37359, n37367, n37365, n37364, n37366,
    n37368, n37373, n37370, n37372, n37378, n37376, n37375, n37377, n37379,
    n37381, n37387, n37384, n37386, n37388, n39026, n39028, n37390, n38667,
    n37394, n37391, n37392, n37435, n37393, n37400, n37395, n38805, n37397,
    n37525, n37398, n37399, n37402, n37425, n37406, n38180, n37414, n37813,
    n37403, n37404, n37405, n37409, n37407, n37408, n37412, n37440, n37419,
    n37416, n37410, n38761, n37411, n37413, n37418, n37415, n37423, n37417,
    n37422, n37420, n37437, n37421, n37427, n37424, n37426, n37434, n38114,
    n37431, n37674, n37429, n38403, n38328, n37430, n37432, n37433, n39029,
    n38557, n38033, n37532, n37732, n37439, n38558, n38458, n37438, n37448,
    n38559, n38652, n38640, n37595, n38182, n38485, n37442, n37443, n37444,
    n37445, n37506, n37447, n37452, n38568, n38556, n37450, n38560, n37724,
    n37598, n37513, n37449, n37451, n38579, n37455, n38576, n37454, n37458,
    n37457, n37462, n38582, n37460, n38575, n37459, n37461, n38591, n37465,
    n38594, n37464, n37468, n37466, n37467, n37472, n38588, n37470, n38587,
    n37469, n37471, n38599, n37477, n38600, n37475, n38603, n37474, n37476,
    n37481, n37522, n37479, n38606, n37478, n37480, n38611, n37486, n38612,
    n37484, n38615, n37483, n37485, n37491, n37487, n37489, n38618, n37488,
    n37490, n38627, n37493, n37492, n37496, n37515, n38630, n37495, n37500,
    n38624, n37498, n38623, n37497, n37499, n38641, n37504, n38637, n37503,
    n37508, n37507, n37512, n38644, n37510, n38635, n37509, n37511, n38653,
    n37521, n38650, n37517, n38651, n37516, n37519, n38658, n37518, n37520,
    n37524, n37523, n37529, n38567, n37527, n37526, n37588, n37528, n37531,
    n37530, n37536, n37534, n37585, n37533, n37535, n37538, n37537, n37544,
    n37540, n37539, n37542, n37541, n37543, n37546, n37545, n37552, n37548,
    n37547, n37550, n37549, n37551, n37554, n37553, n37556, n37555, n37560,
    n37558, n37557, n37559, n37562, n37561, n37564, n37563, n37568, n37566,
    n37565, n37567, n37574, n37570, n37569, n37572, n37571, n37573, n37576,
    n37575, n37578, n37577, n37580, n37579, n37584, n37582, n37581, n37583,
    n37587, n37586, n37594, n37590, n37589, n37592, n37591, n37593, n37740,
    n37657, n37597, n37596, n37608, n37604, n37599, n37600, n37601, n37602,
    n37664, n37603, n37606, n37605, n37607, n37610, n37609, n37616, n37612,
    n37611, n37614, n37613, n37615, n37618, n37617, n37624, n37620, n37619,
    n37622, n37621, n37623, n37626, n37625, n37632, n37628, n37627, n37630,
    n37629, n37631, n37634, n37633, n37640, n37636, n37635, n37638, n37637,
    n37639, n37642, n37641, n37648, n37644, n37643, n37646, n37645, n37647,
    n37650, n37649, n37656, n37652, n37651, n37654, n37653, n37655, n37663,
    n37659, n37658, n37661, n37660, n37662, n37666, n37665, n37673, n37814,
    n37953, n37671, n37729, n37669, n37668, n37670, n37672, n37679, n37675,
    n37677, n37676, n37970, n37733, n37678, n37681, n37680, n37687, n37683,
    n37682, n37685, n37684, n37686, n37691, n37689, n37688, n37690, n37695,
    n37693, n37692, n37694, n37697, n37696, n37703, n37699, n37698, n37701,
    n37700, n37702, n37707, n37705, n37704, n37706, n37711, n37709, n37708,
    n37710, n37717, n37713, n37712, n37715, n37714, n37716, n37719, n37718,
    n37723, n37721, n37720, n37722, n37728, n37726, n37725, n37727, n37731,
    n37730, n37739, n37735, n37734, n37737, n37736, n37738, n38776, n37968,
    n37889, n37802, n37748, n37741, n37742, n37743, n37744, n37806, n37746,
    n37745, n37747, n37752, n37750, n37749, n37751, n37754, n37753, n37760,
    n37756, n37755, n37758, n37757, n37759, n37764, n37762, n37761, n37763,
    n37768, n37766, n37765, n37767, n37772, n37770, n37769, n37771, n37776,
    n37774, n37773, n37775, n37780, n37778, n37777, n37779, n37784, n37782,
    n37781, n37783, n37786, n37785, n37792, n37788, n37787, n37790, n37789,
    n37791, n37796, n37794, n37793, n37795, n37801, n37799, n37798, n37800,
    n37804, n37803, n37812, n37808, n37807, n37810, n37809, n37811, n38099,
    n37818, n37886, n37821, n37816, n37815, n37883, n37817, n37820, n37819,
    n37825, n37875, n37823, n37822, n37824, n37827, n37826, n37833, n37829,
    n37828, n37831, n37830, n37832, n37835, n37834, n37841, n37837, n37836,
    n37839, n37838, n37840, n37843, n37842, n37849, n37845, n37844, n37847,
    n37846, n37848, n37851, n37850, n37857, n37853, n37852, n37855, n37854,
    n37856, n37859, n37858, n37865, n37861, n37860, n37863, n37862, n37864,
    n37867, n37866, n37874, n37869, n37868, n37872, n37871, n37873, n37882,
    n37877, n37876, n37880, n37879, n37881, n37885, n37884, n37898, n37888,
    n37890, n38036, n37950, n37887, n37896, n37891, n37894, n38160, n38172,
    n37892, n37893, n37958, n37895, n37897, n37900, n37899, n37902, n37901,
    n37908, n37904, n37903, n37906, n37905, n37907, n37910, n37909, n37916,
    n37912, n37911, n37914, n37913, n37915, n37918, n37917, n37924, n37920,
    n37919, n37922, n37921, n37923, n37926, n37925, n37932, n37928, n37927,
    n37930, n37929, n37931, n37934, n37933, n37940, n37936, n37935, n37938,
    n37937, n37939, n37943, n37942, n37949, n37945, n37944, n37947, n37946,
    n37948, n37957, n37952, n37951, n37955, n37954, n37956, n37960, n37959,
    n37966, n37964, n38022, n37962, n37961, n37963, n37965, n37972, n37967,
    n37969, n38030, n37971, n37976, n37974, n37973, n37975, n37980, n37978,
    n37977, n37979, n37984, n37982, n37981, n37983, n37988, n37986, n37985,
    n37987, n37992, n37990, n37989, n37991, n37996, n37994, n37993, n37995,
    n37998, n37997, n38004, n38000, n37999, n38002, n38001, n38003, n38006,
    n38005, n38012, n38008, n38007, n38010, n38009, n38011, n38014, n38013,
    n38021, n38016, n38015, n38019, n38018, n38020, n38029, n38024, n38023,
    n38027, n38026, n38028, n38032, n38031, n38263, n38320, n38181, n38096,
    n38035, n38034, n38046, n38042, n38037, n38038, n38039, n38040, n38104,
    n38041, n38044, n38043, n38045, n38048, n38047, n38054, n38050, n38049,
    n38052, n38051, n38053, n38056, n38055, n38062, n38058, n38057, n38060,
    n38059, n38061, n38064, n38063, n38070, n38066, n38065, n38068, n38067,
    n38069, n38072, n38071, n38078, n38074, n38073, n38076, n38075, n38077,
    n38080, n38079, n38086, n38082, n38081, n38084, n38083, n38085, n38089,
    n38088, n38095, n38091, n38090, n38093, n38092, n38094, n38103, n38098,
    n38097, n38101, n38100, n38102, n38106, n38105, n38113, n38107, n38383,
    n38395, n38111, n38109, n38169, n38108, n38110, n38112, n38119, n38117,
    n38116, n38173, n38118, n38121, n38120, n38127, n38123, n38122, n38125,
    n38124, n38126, n38129, n38128, n38135, n38131, n38130, n38133, n38132,
    n38134, n38137, n38136, n38143, n38139, n38138, n38141, n38140, n38142,
    n38145, n38144, n38151, n38147, n38146, n38149, n38148, n38150, n38157,
    n38153, n38152, n38155, n38154, n38156, n38159, n38158, n38162, n38161,
    n38168, n38164, n38163, n38166, n38165, n38167, n38171, n38170, n38179,
    n38175, n38174, n38177, n38176, n38178, n38256, n38455, n38188, n38183,
    n38191, n38186, n38184, n38185, n38253, n38187, n38190, n38189, n38195,
    n38335, n38245, n38193, n38192, n38194, n38197, n38196, n38203, n38199,
    n38198, n38201, n38200, n38202, n38205, n38204, n38211, n38207, n38206,
    n38209, n38208, n38210, n38213, n38212, n38219, n38215, n38214, n38217,
    n38216, n38218, n38221, n38220, n38227, n38223, n38222, n38225, n38224,
    n38226, n38229, n38228, n38235, n38231, n38230, n38233, n38232, n38234,
    n38237, n38236, n38244, n38239, n38238, n38242, n38241, n38243, n38252,
    n38247, n38246, n38250, n38249, n38251, n38255, n38254, n38262, n38406,
    n38317, n38258, n38257, n38260, n38548, n38259, n38261, n38267, n38265,
    n38264, n38325, n38266, n38269, n38268, n38275, n38271, n38270, n38273,
    n38272, n38274, n38277, n38276, n38283, n38279, n38278, n38281, n38280,
    n38282, n38285, n38284, n38291, n38287, n38286, n38289, n38288, n38290,
    n38293, n38292, n38299, n38295, n38294, n38297, n38296, n38298, n38305,
    n38301, n38300, n38303, n38302, n38304, n38307, n38306, n38310, n38309,
    n38316, n38312, n38311, n38314, n38313, n38315, n38324, n38319, n38318,
    n38322, n38321, n38323, n38327, n38326, n38334, n38657, n38332, n38636,
    n38484, n38392, n38330, n38329, n38331, n38333, n38342, n38336, n38337,
    n38338, n38339, n38396, n38341, n38344, n38343, n38350, n38346, n38345,
    n38348, n38347, n38349, n38354, n38352, n38351, n38353, n38358, n38356,
    n38355, n38357, n38360, n38359, n38366, n38362, n38361, n38364, n38363,
    n38365, n38368, n38367, n38374, n38370, n38369, n38372, n38371, n38373,
    n38380, n38376, n38375, n38378, n38377, n38379, n38382, n38381, n38385,
    n38384, n38391, n38387, n38386, n38389, n38388, n38390, n38394, n38393,
    n38402, n38398, n38397, n38400, n38399, n38401, n38569, n38465, n38405,
    n38404, n38414, n38410, n38408, n38407, n38469, n38409, n38412, n38411,
    n38413, n38416, n38415, n38422, n38418, n38417, n38420, n38419, n38421,
    n38424, n38423, n38430, n38426, n38425, n38428, n38427, n38429, n38432,
    n38431, n38438, n38434, n38433, n38436, n38435, n38437, n38440, n38439,
    n38446, n38442, n38441, n38444, n38443, n38445, n38448, n38447, n38454,
    n38450, n38449, n38452, n38451, n38453, n38457, n38456, n38464, n38460,
    n38459, n38462, n38461, n38463, n38467, n38466, n38475, n38471, n38470,
    n38473, n38472, n38474, n38482, n38544, n38478, n38477, n38480, n38479,
    n38481, n38493, n38486, n38491, n38488, n38490, n38553, n38492, n38495,
    n38494, n38501, n38497, n38496, n38499, n38498, n38500, n38503, n38502,
    n38509, n38505, n38504, n38507, n38506, n38508, n38511, n38510, n38517,
    n38513, n38512, n38515, n38514, n38516, n38519, n38518, n38525, n38521,
    n38520, n38523, n38522, n38524, n38527, n38526, n38533, n38529, n38528,
    n38531, n38530, n38532, n38536, n38535, n38543, n38539, n38538, n38541,
    n38540, n38542, n38552, n38547, n38546, n38550, n38549, n38551, n38555,
    n38554, n38566, n38564, n38562, n38649, n38561, n38563, n38565, n38574,
    n38572, n38571, n38663, n38573, n38578, n38577, n38586, n38581, n38580,
    n38584, n38583, n38585, n38590, n38589, n38598, n38593, n38592, n38596,
    n38595, n38597, n38602, n38601, n38610, n38605, n38604, n38608, n38607,
    n38609, n38614, n38613, n38622, n38617, n38616, n38620, n38619, n38621,
    n38626, n38625, n38634, n38629, n38628, n38632, n38631, n38633, n38639,
    n38638, n38648, n38643, n38642, n38646, n38645, n38647, n38662, n38656,
    n38655, n38660, n38659, n38661, n38665, n38664, n38666, n39033, n38672,
    n38669, n38671, n38685, n38676, n38680, n38679, n38684, n38683, n39100,
    n38787, n38722, n38690, n38691, n38693, n38698, n38697, n38762, n38700,
    n38699, n38702, n38701, n38716, n38708, n38707, n38735, n38712, n38711,
    n38714, n38713, n38715, n38718, n38717, n39045, n38720, n38755, n38754,
    n38727, n38726, n38729, n38731, n38734, n38733, n38739, n38737, n38738,
    n38751, n38741, n38749, n38743, n38747, n38746, n38748, n38750, n39037,
    n39030, n38753, n38752, n38780, n38785, n38778, n38774, n38765, n38760,
    n38759, n39072, n38771, n38764, n38767, n38766, n39055, n38769, n38770,
    n38772, n38773, n38777, n38779, n38783, n38782, n38784, n38786, n38789,
    n38795, n38794, n38813, n38791, n38792, n38793, n38807, n38802, n38798,
    n38800, n38801, n39024, n38812, n38817, n38809, n38822, n38826, n38821,
    n38816, n38819, n38820, n38824, n38825, n38850, n38836, n38828, n38829,
    n38834, n44540, n38830, n38848, n38832, n38849, n38847, n38833, n38835,
    n38846, n38837, n38842, n38838, n38844, n38856, n38839, n38840, n38841,
    n38843, n38845, n38859, n38853, n38851, n38852, n38855, n38857, n38858,
    n38975, n38862, n38861, n38864, n38863, n38867, n38866, n38869, n39125,
    n38868, n38872, n38871, n38874, n38873, n38877, n38876, n38879, n38878,
    n38885, n38882, n38881, n38884, n38883, n38887, n38886, n38889, n38888,
    n38895, n38892, n38891, n38894, n38893, n38897, n38896, n38899, n38898,
    n38902, n38901, n38904, n38903, n38907, n38906, n38909, n38908, n38912,
    n38911, n38914, n38913, n38917, n38916, n38919, n38918, n38922, n38921,
    n38924, n38923, n38927, n38926, n38929, n38928, n38935, n38932, n38931,
    n38934, n38933, n38937, n38936, n38939, n38938, n38945, n38942, n38941,
    n38944, n38943, n38947, n38946, n38949, n38948, n38955, n38952, n38951,
    n38954, n38953, n38957, n38956, n38959, n38958, n38962, n38961, n38964,
    n38963, n38967, n38966, n38969, n38968, n38976, n38972, n38971, n38974,
    n38973, n38978, n38977, n38980, n38979, n38986, n38983, n38982, n38985,
    n38984, n38991, n38988, n38987, n38990, n38989, n38993, n38992, n38995,
    n38994, n38997, n38996, n38999, n38998, n39004, n39001, n39000, n39003,
    n39002, n39008, n39007, n39010, n39009, n39012, n39011, n39014, n39013,
    n39016, n39015, n39018, n39017, n39021, n39020, n39022, n39025, n39027,
    n39032, n39031, n39034, n39036, n39035, n39041, n39040, n39042, n39044,
    n39043, n39051, n39061, n39060, n39049, n39048, n39050, n39052, n39054,
    n39053, n39059, n39058, n39064, n39062, n39063, n39065, n39067, n39066,
    n39071, n39070, n39075, n39074, n39076, n39080, n39079, n39091, n39088,
    n39093, n39086, n39085, n39087, n39089, n39094, n39090, n39096, n39095,
    n39099, n39098, n39103, n39102, n39109, n39107, n39108, n39122, n39124,
    n39111, n39113, n39116, n39115, n39117, n39119, n39121, n39123, n39128,
    n39127, n39134, n39131, n39135, n39133, n39137, n39139, n39142, n39143,
    n39144, n39146, n39145, n39147, n39148, n41897, n42070, n39149, n39152,
    n39151, n42224, n42223, n39155, n41911, n39154, n39157, n39156, n42245,
    n39158, n42074, n39159, n42193, n42191, n39162, n39165, n39164, n39169,
    n39167, n39166, n39168, n39193, n39171, n39170, n39175, n39173, n39172,
    n39174, n39191, n39177, n39176, n39181, n39179, n39178, n39180, n39189,
    n39183, n39182, n39187, n39185, n39184, n39186, n39188, n39190, n39192,
    n39210, n39207, n39195, n39200, n39194, n39198, n39196, n39206, n39197,
    n39199, n39203, n39208, n39201, n39202, n39205, n39204, n39209, n39212,
    n39211, n39213, n39223, n39221, n39216, n39218, n39220, n39222, n39227,
    n39226, n39228, n39229, n39241, n39239, n39237, n39232, n39233, n39235,
    n39234, n39236, n39238, n39240, n39247, n39245, n39244, n39246, n39266,
    n39673, n39252, n39250, n39249, n39251, n39254, n39253, n39257, n39256,
    n39264, n39260, n39262, n39263, n39265, n39269, n39268, n39279, n39273,
    n39274, n39277, n39276, n39278, n39289, n39287, n39282, n39281, n39283,
    n39285, n39284, n39286, n39288, n39307, n39292, n39303, n39294, n39293,
    n39295, n39301, n39299, n39298, n39300, n39302, n39305, n39304, n39306,
    n39310, n39309, n39312, n39311, n39323, n39316, n39314, n39315, n39321,
    n39318, n39319, n39320, n39322, n39332, n39327, n39326, n39330, n39329,
    n39331, n39334, n39350, n39346, n39338, n39337, n39339, n39344, n39342,
    n39697, n39341, n39343, n39345, n39348, n39347, n39349, n39353, n39829,
    n39352, n39355, n39354, n39366, n39357, n39359, n39707, n39358, n39364,
    n39361, n39362, n39363, n39365, n39373, n39369, n39368, n39371, n39370,
    n39372, n39375, n39374, n39386, n39378, n39716, n39377, n39384, n39387,
    n39381, n39382, n39383, n39385, n39393, n39389, n39388, n39391, n39390,
    n39392, n39395, n39411, n39401, n39398, n39397, n39399, n39400, n39404,
    n39403, n39409, n39724, n39407, n39860, n39406, n39408, n39410, n39413,
    n39412, n39415, n39414, n39425, n39418, n39417, n39423, n39426, n39420,
    n39421, n39422, n39424, n39433, n39428, n39427, n39431, n39865, n39430,
    n39432, n39435, n39434, n39436, n39438, n39437, n39442, n39440, n39441,
    n39448, n39446, n39445, n39447, n39452, n39450, n39449, n39451, n39455,
    n39454, n39457, n39456, n39468, n39460, n39754, n39459, n39466, n39469,
    n39463, n39464, n39465, n39467, n39475, n39471, n39470, n39473, n39472,
    n39474, n39477, n39476, n39478, n39483, n39481, n39480, n39482, n39491,
    n39486, n39487, n39489, n39488, n39490, n39494, n39768, n39493, n39771,
    n39509, n39777, n39507, n39887, n39500, n39499, n39505, n39502, n39501,
    n39503, n39504, n39506, n39508, n39515, n39512, n39513, n39514, n39517,
    n39519, n39518, n39529, n39523, n39522, n39525, n39524, n39527, n39526,
    n39528, n39535, n39532, n39533, n39534, n39542, n39537, n39536, n39538,
    n39540, n39539, n39541, n39548, n39546, n39545, n39547, n39554, n39551,
    n39552, n39553, n39556, n39555, n39557, n39563, n39917, n39561, n39560,
    n39562, n39571, n39566, n39567, n39569, n39568, n39570, n39573, n39572,
    n39575, n39574, n39576, n39578, n39577, n39597, n39581, n40278, n39585,
    n39584, n39592, n39590, n39589, n40357, n39591, n39595, n39780, n39916,
    n39676, n39594, n39596, n39602, n39599, n39600, n39601, n39604, n39603,
    n39611, n39607, n39606, n39609, n39608, n39610, n39617, n39614, n39615,
    n39616, n39619, n39623, n42141, n39622, n39625, n39624, n39635, n39908,
    n42158, n39631, n39630, n39633, n39632, n39634, n39643, n42156, n39638,
    n39641, n39640, n39642, n39649, n39645, n39646, n39648, n39651, n39650,
    n39655, n42094, n39654, n39671, n39658, n39657, n39664, n39662, n39959,
    n39661, n39663, n39669, n39666, n39668, n39670, n39674, n39696, n42093,
    n39694, n39692, n39680, n39679, n39690, n39685, n39684, n39688, n39687,
    n39689, n39691, n39693, n39695, n39703, n39700, n39832, n39702, n39706,
    n39705, n39712, n39710, n39711, n39715, n39714, n39720, n39718, n39719,
    n39723, n39722, n39731, n39727, n39728, n39730, n39734, n39733, n39735,
    n39740, n39764, n39755, n39745, n39747, n39738, n39739, n39743, n39742,
    n39750, n39746, n39748, n39749, n39753, n39752, n39758, n39756, n39757,
    n39761, n39760, n39767, n39763, n39765, n39766, n39770, n39769, n39776,
    n39774, n39775, n39779, n39778, n39786, n39798, n39781, n39784, n39783,
    n39785, n39789, n39788, n39793, n39791, n39792, n39796, n39795, n39801,
    n39797, n39799, n39800, n39804, n39803, n39806, n39807, n39809, n39808,
    n39811, n39813, n39812, n39816, n39815, n39819, n39818, n39821, n39825,
    n39823, n39822, n39824, n39827, n39826, n39831, n39830, n39834, n39952,
    n39833, n39845, n39838, n39837, n39836, n39843, n39841, n39840, n39842,
    n39844, n39848, n39847, n39854, n39962, n39852, n39851, n40271, n39853,
    n39857, n39856, n39859, n39858, n39862, n39861, n39864, n39863, n39867,
    n39866, n39869, n39868, n39871, n39873, n39872, n39875, n39874, n39878,
    n39877, n39880, n39879, n39882, n39884, n39883, n39886, n39885, n39890,
    n39889, n39892, n39891, n39895, n40154, n39894, n39897, n39896, n39901,
    n40149, n39900, n39903, n39902, n39907, n39905, n39904, n39906, n39921,
    n39914, n39935, n39912, n39940, n42166, n39910, n39950, n39951, n39909,
    n39941, n39911, n39936, n39913, n39915, n39927, n39918, n39919, n39920,
    n39923, n39922, n39925, n39924, n39930, n39928, n39929, n39932, n39931,
    n39934, n39933, n39939, n39937, n39938, n39942, n39949, n39944, n39943,
    n39947, n39946, n39948, n39953, n39958, n39956, n39955, n39957, n39961,
    n39960, n39969, n39967, n39965, n39966, n39968, n39972, n39971, n39974,
    n42213, n39979, n39978, n39981, n39980, n39983, n39982, n39985, n39984,
    n39987, n39986, n39989, n39988, n39991, n39990, n39993, n39992, n39995,
    n39994, n39997, n39996, n39999, n39998, n40001, n40000, n40003, n40002,
    n40005, n40004, n40007, n40006, n40009, n40008, n40011, n40010, n40013,
    n40012, n40015, n40014, n40017, n40016, n40019, n40018, n40021, n40020,
    n40024, n40023, n40026, n40025, n40028, n40027, n40030, n40029, n40032,
    n40031, n40034, n40033, n40036, n40035, n40039, n40038, n40042, n40041,
    n40044, n40043, n40047, n40046, n40049, n40048, n40052, n40051, n40054,
    n40053, n40057, n40056, n40059, n40058, n40062, n40061, n40064, n40063,
    n40067, n40066, n40069, n40068, n40072, n40071, n40074, n40073, n40079,
    n40078, n40081, n40080, n40083, n40082, n40085, n40084, n40087, n40086,
    n40089, n40088, n40091, n40090, n40093, n40092, n40095, n40094, n40097,
    n40096, n40099, n40098, n40101, n40100, n40103, n40102, n40105, n40104,
    n40107, n40106, n40110, n40109, n40113, n40112, n40116, n40115, n40120,
    n40201, n40119, n40122, n40270, n40121, n40125, n40124, n40206, n40127,
    n40126, n40130, n40129, n40211, n40132, n40131, n40135, n40134, n40216,
    n40137, n40136, n40140, n40139, n40221, n40142, n40141, n40226, n40145,
    n40144, n40227, n40147, n40146, n40150, n40232, n40152, n40151, n40155,
    n40237, n40157, n40156, n40161, n40160, n40241, n40163, n40162, n40167,
    n40166, n40245, n40169, n40168, n40173, n40172, n40250, n40175, n40174,
    n40176, n40179, n40178, n40254, n40181, n40180, n40185, n40184, n40258,
    n40187, n40186, n40188, n40191, n40190, n40262, n40193, n40192, n40197,
    n40196, n40266, n40199, n40198, n40202, n40204, n40203, n40207, n40209,
    n40208, n40212, n40214, n40213, n40217, n40219, n40218, n40222, n40224,
    n40223, n40228, n40230, n40229, n40233, n40235, n40234, n40238, n40240,
    n40239, n40242, n40244, n40243, n40246, n40248, n40247, n40251, n40253,
    n40252, n40255, n40257, n40256, n40259, n40261, n40260, n40263, n40265,
    n40264, n40267, n40269, n40268, n40277, n40275, n40272, n40274, n40276,
    n40358, n40283, n40280, n40355, n40282, n40292, n40288, n40287, n40290,
    n40369, n40291, n40300, n40298, n40366, n40296, n40295, n40297, n40299,
    n40381, n40314, n40310, n40307, n40374, n40309, n40312, n40311, n40313,
    n40318, n40379, n40315, n40317, n40321, n40398, n40334, n40400, n40328,
    n40326, n40409, n40327, n40332, n40331, n40333, n40336, n40335, n40339,
    n40340, n40354, n40352, n40345, n40350, n40349, n40351, n40353, n40364,
    n40362, n40359, n40361, n40363, n40365, n40373, n40371, n40370, n40372,
    n40376, n40375, n40396, n40394, n40380, n40383, n40382, n40386, n40385,
    n40387, n40392, n40391, n40393, n40395, n40407, n40402, n40401, n40405,
    n40404, n40406, n40416, n40410, n40414, n40411, n40413, n40415, n40448,
    n41155, n40417, n40580, n40418, n40419, n40431, n40420, n40427, n40424,
    n40422, n40423, n40425, n40426, n40443, n41773, n40430, n40434, n40433,
    n40441, n40439, n40438, n40440, n40442, n41775, n40450, n40447, n40446,
    n41774, n40449, n40451, n40464, n40455, n40454, n41802, n40458, n41597,
    n40457, n40462, n40460, n40459, n40461, n40463, n41799, n40466, n40479,
    n40470, n40469, n41807, n40473, n40551, n40472, n40477, n40475, n40474,
    n40476, n40478, n41811, n40481, n40494, n40485, n40484, n41826, n40488,
    n41820, n40487, n40492, n40490, n40489, n40491, n40493, n41823, n40496,
    n40509, n40500, n40499, n41831, n40503, n40502, n40507, n40505, n40504,
    n40506, n40508, n40512, n41725, n41835, n40511, n40527, n40517, n40516,
    n41843, n40521, n41844, n40520, n40525, n40523, n40522, n40524, n40526,
    n41730, n41847, n40529, n40542, n40534, n40533, n41862, n40536, n40535,
    n40540, n40538, n40537, n40539, n40541, n41859, n40544, n40564, n40550,
    n40549, n41879, n40555, n40554, n40562, n40559, n40558, n40561, n40563,
    n41753, n41875, n40567, n40576, n40636, n40570, n40569, n40640, n40574,
    n40572, n40571, n40573, n40575, n40587, n40578, n40579, n40584, n40581,
    n40583, n40585, n40586, n40593, n40589, n40588, n40591, n40590, n40592,
    n40595, n40594, n40601, n40597, n40596, n40599, n40598, n40600, n40603,
    n40602, n40609, n40605, n40604, n40607, n40606, n40608, n40611, n40610,
    n40617, n40613, n40612, n40615, n40614, n40616, n40619, n40618, n40625,
    n40621, n40620, n40623, n40622, n40624, n40627, n40626, n40633, n40629,
    n40628, n40631, n40630, n40632, n40635, n40634, n40644, n40639, n40638,
    n40642, n40641, n40643, n40647, n40646, n40671, n40723, n40656, n40650,
    n40649, n40662, n40652, n40651, n40653, n40654, n40655, n40669, n40658,
    n40659, n40667, n40660, n40661, n40664, n40663, n40665, n40666, n40726,
    n40668, n40670, n40673, n40672, n40675, n40674, n40681, n40677, n40676,
    n40679, n40678, n40680, n40683, n40682, n40689, n40685, n40684, n40687,
    n40686, n40688, n40691, n40690, n40697, n40693, n40692, n40695, n40694,
    n40696, n40699, n40698, n40705, n40701, n40700, n40703, n40702, n40704,
    n40707, n40706, n40713, n40709, n40708, n40711, n40710, n40712, n40715,
    n40714, n40721, n40717, n40716, n40719, n40718, n40720, n40725, n40724,
    n40733, n40728, n40727, n40731, n40730, n40732, n40735, n40739, n40737,
    n40736, n40747, n40738, n40754, n40743, n40742, n40752, n40744, n40745,
    n40749, n40748, n40750, n40815, n40751, n40753, n40757, n40756, n40761,
    n40759, n40758, n40760, n40765, n40763, n40762, n40764, n40767, n40766,
    n40773, n40769, n40768, n40771, n40770, n40772, n40777, n40775, n40774,
    n40776, n40781, n40779, n40778, n40780, n40783, n40782, n40789, n40785,
    n40784, n40787, n40786, n40788, n40793, n40791, n40790, n40792, n40797,
    n40795, n40794, n40796, n40803, n40799, n40798, n40801, n40800, n40802,
    n40805, n40804, n40814, n40810, n40809, n40812, n40811, n40813, n40817,
    n40816, n40834, n40838, n40895, n40830, n40835, n40818, n40828, n40819,
    n40913, n40977, n40899, n40821, n40822, n40841, n40826, n40825, n40824,
    n41494, n40840, n40827, n40896, n40829, n40832, n40831, n40833, n40845,
    n40836, n40837, n40839, n40843, n40842, n40844, n40851, n40847, n40846,
    n40849, n40848, n40850, n40853, n40852, n40855, n40854, n40861, n40857,
    n40856, n40859, n40858, n40860, n40863, n40862, n40869, n40865, n40864,
    n40867, n40866, n40868, n40875, n40871, n40870, n40873, n40872, n40874,
    n40877, n40876, n40883, n40879, n40878, n40881, n40880, n40882, n40885,
    n40884, n40887, n40886, n40893, n40889, n40888, n40891, n40890, n40892,
    n40903, n40898, n40897, n40901, n40900, n40902, n40906, n40905, n40917,
    n40978, n40912, n40907, n40910, n40908, n40923, n40909, n40911, n40915,
    n40914, n40916, n40928, n40918, n40919, n40921, n40926, n40924, n40925,
    n40927, n40930, n40929, n40936, n40932, n40931, n40934, n40933, n40935,
    n40942, n40938, n40937, n40940, n40939, n40941, n40944, n40943, n40946,
    n40945, n40952, n40948, n40947, n40950, n40949, n40951, n40954, n40953,
    n40960, n40956, n40955, n40958, n40957, n40959, n40962, n40961, n40968,
    n40964, n40963, n40966, n40965, n40967, n40970, n40969, n40976, n40972,
    n40971, n40974, n40973, n40975, n40980, n40979, n40989, n40984, n40983,
    n40987, n40986, n40988, n41012, n41005, n41064, n40996, n41001, n40990,
    n40994, n40999, n40993, n40995, n41010, n40997, n40998, n41000, n41008,
    n41003, n41004, n41006, n41007, n41067, n41009, n41011, n41014, n41013,
    n41016, n41015, n41022, n41018, n41017, n41020, n41019, n41021, n41024,
    n41023, n41030, n41026, n41025, n41028, n41027, n41029, n41032, n41031,
    n41038, n41034, n41033, n41036, n41035, n41037, n41040, n41039, n41046,
    n41042, n41041, n41044, n41043, n41045, n41048, n41047, n41054, n41050,
    n41049, n41052, n41051, n41053, n41056, n41055, n41062, n41058, n41057,
    n41060, n41059, n41061, n41066, n41065, n41075, n41070, n41069, n41073,
    n41072, n41074, n41085, n41076, n41078, n41077, n41084, n41080, n41079,
    n41082, n41579, n41081, n41083, n41094, n41086, n41087, n41088, n41092,
    n41090, n41091, n41093, n41100, n41096, n41095, n41098, n41097, n41099,
    n41102, n41101, n41108, n41104, n41103, n41106, n41105, n41107, n41110,
    n41109, n41116, n41112, n41111, n41114, n41615, n41113, n41115, n41118,
    n41117, n41124, n41120, n41119, n41122, n41121, n41123, n41126, n41125,
    n41132, n41128, n41127, n41130, n41633, n41129, n41131, n41134, n41133,
    n41140, n41136, n41135, n41138, n41137, n41139, n41142, n41141, n41150,
    n41146, n41145, n41148, n41652, n41147, n41149, n41153, n41152, n41167,
    n41154, n41172, n41163, n41232, n41156, n41157, n41170, n41168, n41161,
    n41159, n41160, n41229, n41162, n41165, n41164, n41166, n41178, n41169,
    n41171, n41176, n41173, n41174, n41175, n41177, n41182, n41180, n41179,
    n41181, n41186, n41184, n41183, n41185, n41190, n41188, n41187, n41189,
    n41194, n41192, n41191, n41193, n41198, n41196, n41195, n41197, n41202,
    n41200, n41199, n41201, n41208, n41204, n41203, n41206, n41205, n41207,
    n41210, n41209, n41216, n41212, n41211, n41214, n41213, n41215, n41218,
    n41217, n41224, n41220, n41219, n41222, n41221, n41223, n41226, n41225,
    n41236, n41231, n41230, n41234, n41233, n41235, n41239, n41238, n41240,
    n41395, n41251, n41249, n41241, n41245, n41243, n41257, n41244, n41247,
    n41246, n41248, n41250, n41261, n41252, n41253, n41254, n41259, n41256,
    n41258, n41260, n41265, n41263, n41262, n41264, n41269, n41267, n41266,
    n41268, n41273, n41271, n41270, n41272, n41277, n41275, n41274, n41276,
    n41283, n41281, n41279, n41278, n41280, n41282, n41285, n41284, n41291,
    n41289, n41287, n41286, n41288, n41290, n41293, n41292, n41299, n41297,
    n41295, n41294, n41296, n41298, n41301, n41300, n41305, n41303, n41302,
    n41304, n41309, n41307, n41306, n41308, n41317, n41315, n41313, n41312,
    n41314, n41316, n41320, n41319, n41321, n41400, n41322, n41323, n41334,
    n41325, n41423, n41338, n41332, n41327, n41328, n41403, n41346, n41331,
    n41396, n41330, n41344, n41333, n41335, n41342, n41337, n41339, n41340,
    n41341, n41343, n41345, n41348, n41347, n41352, n41350, n41349, n41351,
    n41356, n41354, n41353, n41355, n41358, n41357, n41364, n41360, n41359,
    n41362, n41361, n41363, n41366, n41365, n41372, n41368, n41367, n41370,
    n41369, n41371, n41376, n41374, n41373, n41375, n41377, n41380, n41379,
    n41386, n41382, n41381, n41384, n41383, n41385, n41392, n41388, n41387,
    n41390, n41389, n41391, n41394, n41393, n41398, n41397, n41407, n41402,
    n41401, n41405, n41404, n41406, n41478, n41408, n41410, n41409, n41417,
    n41415, n41413, n41412, n41414, n41416, n41428, n41419, n41420, n41421,
    n41426, n41424, n41425, n41427, n41434, n41432, n41430, n41429, n41431,
    n41433, n41436, n41435, n41442, n41440, n41438, n41437, n41439, n41441,
    n41444, n41443, n41450, n41448, n41446, n41445, n41447, n41449, n41452,
    n41451, n41458, n41456, n41454, n41453, n41455, n41457, n41460, n41459,
    n41466, n41464, n41462, n41461, n41463, n41465, n41468, n41467, n41474,
    n41472, n41470, n41469, n41471, n41473, n41476, n41475, n41485, n41483,
    n41481, n41480, n41482, n41484, n41488, n41487, n41502, n41564, n41500,
    n41498, n41492, n41496, n41508, n41495, n41497, n41499, n41501, n41513,
    n41504, n41505, n41506, n41511, n41507, n41509, n41510, n41512, n41517,
    n41515, n41514, n41516, n41521, n41519, n41518, n41520, n41525, n41523,
    n41522, n41524, n41529, n41527, n41526, n41528, n41533, n41531, n41530,
    n41532, n41537, n41535, n41534, n41536, n41541, n41539, n41538, n41540,
    n41545, n41543, n41542, n41544, n41549, n41547, n41546, n41548, n41553,
    n41551, n41550, n41552, n41557, n41555, n41554, n41556, n41561, n41559,
    n41558, n41560, n41568, n41566, n41565, n41567, n41573, n41571, n41570,
    n41572, n41586, n41576, n41578, n41577, n41585, n41583, n41581, n41580,
    n41582, n41584, n41596, n41587, n41588, n41589, n41594, n41592, n41593,
    n41595, n41603, n41601, n41599, n41598, n41600, n41602, n41605, n41604,
    n41612, n41610, n41608, n41607, n41609, n41611, n41614, n41613, n41621,
    n41619, n41617, n41616, n41618, n41620, n41623, n41622, n41630, n41628,
    n41626, n41625, n41627, n41629, n41632, n41631, n41639, n41637, n41635,
    n41634, n41636, n41638, n41641, n41640, n41648, n41646, n41644, n41643,
    n41645, n41647, n41650, n41649, n41659, n41657, n41655, n41654, n41656,
    n41658, n41662, n41661, n41663, n41750, n41679, n41674, n41668, n41665,
    n41671, n41757, n41666, n41667, n41681, n41669, n41670, n41752, n41673,
    n41677, n41676, n41678, n41689, n41684, n41682, n41683, n41685, n41687,
    n41688, n41697, n41692, n41691, n41695, n41694, n41696, n41699, n41698,
    n41707, n41702, n41701, n41705, n41704, n41706, n41709, n41708, n41714,
    n41712, n41711, n41713, n41719, n41717, n41716, n41718, n41724, n41722,
    n41721, n41723, n41729, n41727, n41726, n41728, n41737, n41732, n41731,
    n41735, n41734, n41736, n41739, n41738, n41744, n41742, n41741, n41743,
    n41749, n41747, n41746, n41748, n41761, n41755, n41754, n41759, n41758,
    n41760, n41764, n41763, n41781, n41767, n41772, n41791, n41770, n41771,
    n41874, n41779, n41777, n41776, n41778, n41780, n41794, n41783, n41784,
    n41787, n41792, n41790, n41793, n41798, n41797, n41806, n41801, n41800,
    n41804, n41803, n41805, n41810, n41809, n41818, n41813, n41812, n41816,
    n41815, n41817, n41822, n41821, n41830, n41825, n41824, n41828, n41827,
    n41829, n41834, n41833, n41842, n41837, n41836, n41840, n41839, n41841,
    n41846, n41845, n41854, n41849, n41848, n41852, n41851, n41853, n41858,
    n41857, n41866, n41861, n41860, n41864, n41863, n41865, n41872, n41871,
    n41883, n41877, n41876, n41881, n41880, n41882, n41886, n41892, n41888,
    n41889, n41891, n41917, n41903, n41896, n41902, n41921, n41898, n41899,
    n41900, n41901, n41904, n41905, n41908, n41914, n41906, n41907, n41910,
    n41913, n41912, n41915, n41916, n41925, n41919, n41922, n41923, n41924,
    n41928, n42023, n41927, n41930, n41929, n41932, n41935, n41931, n41934,
    n41933, n41937, n41936, n41939, n41938, n41943, n41941, n41940, n41942,
    n41945, n41944, n41947, n41946, n41949, n41948, n41951, n41950, n41955,
    n41953, n41952, n41954, n41959, n41957, n41956, n41958, n41961, n41960,
    n41963, n41962, n41967, n41965, n41964, n41966, n41971, n41969, n41968,
    n41970, n41973, n41972, n41975, n41974, n41979, n41977, n41976, n41978,
    n41981, n41980, n41983, n41982, n41986, n41985, n41988, n41987, n41990,
    n41989, n41992, n41991, n41994, n41993, n41996, n41995, n41999, n41998,
    n42001, n42000, n42005, n42003, n42002, n42004, n42007, n42006, n42009,
    n42008, n42011, n42010, n42013, n42012, n42015, n42014, n42017, n42016,
    n42020, n42019, n42022, n42021, n42027, n42026, n42029, n42028, n42032,
    n42031, n42034, n42033, n42037, n42036, n42039, n42038, n42042, n42041,
    n42044, n42043, n42047, n42046, n42049, n42048, n42052, n42051, n42054,
    n42053, n42058, n42057, n42060, n42059, n42062, n42061, n42064, n42063,
    n42067, n42066, n42069, n42068, n42072, n42071, n42073, n42078, n42077,
    n42081, n42080, n42132, n42083, n42085, n42084, n42128, n42088, n42087,
    n42089, n42091, n42090, n42092, n42124, n42109, n42099, n42098, n42108,
    n42101, n42100, n42104, n42115, n42103, n42105, n42107, n42106, n42110,
    n42114, n42113, n42118, n42117, n42119, n42122, n42121, n42127, n42126,
    n42130, n42129, n42131, n42136, n42135, n42152, n42138, n42169, n42146,
    n42143, n42142, n42144, n42145, n42149, n42148, n42150, n42151, n42185,
    n42162, n42155, n42168, n42157, n42160, n42159, n42161, n42163, n42165,
    n42164, n42167, n42172, n42171, n42173, n42175, n42174, n42178, n42183,
    n42182, n42184, n42188, n42187, n42190, n42189, n42195, n42194, n42198,
    n42203, n42201, n42202, n42220, n42222, n42205, n42212, n42207, n42210,
    n42211, n42218, n42215, n42217, n42219, n42221, n42226, n42225, n42231,
    n42229, n42230, n42233, n42238, n42236, n42237, n42239, n42240, n42242,
    n44828, n42241, n44706, n44523, n42246, n44711, n44709, n42247, n44831,
    n42249, n42251, n42250, n42255, n42253, n42252, n42254, n42279, n42257,
    n42256, n42259, n42258, n42261, n42260, n42277, n42263, n42262, n42267,
    n42265, n42264, n42266, n42275, n42269, n42268, n42273, n42271, n42270,
    n42272, n42274, n42276, n42278, n44823, n42283, n44814, n44813, n42280,
    n42284, n42281, n42282, n42287, n44812, n42285, n42286, n42289, n42288,
    n42292, n42291, n42294, n42311, n42315, n42293, n42295, n42303, n42301,
    n42297, n42299, n42298, n42300, n42302, n42305, n42304, n42310, n42308,
    n42307, n42309, n42321, n42312, n42314, n42319, n42317, n42316, n42318,
    n42320, n42322, n42325, n42523, n42324, n42341, n42339, n42330, n42329,
    n42332, n42331, n42333, n42337, n42335, n42358, n42336, n42338, n42340,
    n42528, n42348, n42344, n42346, n42345, n42347, n42349, n42354, n42352,
    n42351, n42353, n42360, n44571, n42356, n42357, n42359, n42362, n42361,
    n42378, n42365, n42364, n42370, n42366, n42368, n42369, n42376, n42595,
    n42374, n42460, n42375, n42377, n42381, n42405, n42401, n42380, n42383,
    n42382, n42398, n42957, n42387, n42386, n42388, n42396, n42394, n42392,
    n42484, n42395, n42397, n42410, n42903, n42403, n42402, n42408, n42406,
    n42407, n42409, n44556, n42416, n42450, n42465, n42455, n42412, n42430,
    n42415, n42414, n42419, n44551, n42417, n42418, n42428, n42422, n42983,
    n42426, n42424, n42423, n42425, n42427, n42429, n42435, n42433, n42605,
    n42916, n42434, n42437, n42436, n42454, n43000, n42442, n42441, n42448,
    n42445, n42547, n42447, n42449, n42452, n42451, n42453, n42457, n42456,
    n42478, n42933, n42483, n42468, n42463, n43021, n42466, n42467, n42476,
    n42474, n42472, n42471, n42473, n42475, n42477, n42480, n42479, n42499,
    n42952, n42492, n42490, n42487, n43036, n42489, n42491, n42497, n42495,
    n42496, n42498, n42502, n42501, n42505, n42504, n42567, n42509, n42508,
    n42511, n42510, n42515, n42513, n42514, n42517, n42516, n42520, n42519,
    n42522, n42521, n42525, n42524, n42527, n42526, n42530, n42529, n42532,
    n42531, n42535, n42534, n42537, n42536, n42539, n42538, n42542, n42541,
    n42544, n42543, n42546, n42545, n42549, n42922, n42548, n42551, n42550,
    n42552, n42555, n42554, n42558, n42557, n42566, n42560, n42564, n42563,
    n42565, n42569, n42568, n42571, n42570, n42574, n42573, n42576, n42575,
    n42578, n42577, n42581, n42580, n42584, n42583, n42586, n42585, n42589,
    n42588, n42591, n42590, n42594, n42593, n42597, n42596, n42601, n42600,
    n42603, n42602, n42607, n42606, n42609, n42608, n42612, n42611, n42614,
    n42613, n42617, n42616, n42619, n42618, n42624, n42623, n42627, n42626,
    n42629, n42628, n42633, n42630, n42632, n42635, n42634, n42637, n42636,
    n42639, n42638, n42641, n42640, n42643, n42642, n42645, n42644, n42647,
    n42646, n42649, n42648, n42651, n42650, n42653, n42652, n42655, n42654,
    n42657, n42656, n42659, n42658, n42661, n42660, n42663, n42662, n42665,
    n42664, n42667, n42666, n42669, n42668, n42671, n42670, n42673, n42672,
    n42675, n42674, n42677, n42676, n42679, n42678, n42681, n42680, n42683,
    n42682, n42685, n42684, n42687, n42686, n42689, n42688, n42691, n42690,
    n42693, n42692, n42695, n42694, n42697, n42696, n42699, n42698, n42701,
    n42700, n42703, n42702, n42705, n42704, n42707, n42706, n42709, n42708,
    n42711, n42710, n42713, n42712, n42715, n42714, n42717, n42716, n42719,
    n42718, n42721, n42720, n42723, n42722, n42725, n42724, n42727, n42726,
    n42729, n42728, n42731, n42730, n42733, n42732, n42735, n42734, n42737,
    n42736, n42739, n42738, n42741, n42740, n42743, n42742, n42745, n42744,
    n42748, n42747, n42751, n42750, n42754, n42753, n42757, n42756, n42888,
    n42824, n42762, n42764, n42763, n42828, n42765, n42767, n42766, n42832,
    n42768, n42770, n42769, n42836, n42771, n42773, n42772, n42840, n42774,
    n42776, n42775, n43173, n42844, n42778, n42780, n42779, n43187, n42848,
    n42782, n42784, n42783, n43197, n42852, n42786, n42787, n42789, n42788,
    n42791, n42857, n42792, n42794, n42793, n42796, n42861, n42797, n42799,
    n42798, n42801, n42865, n42802, n42804, n42803, n42806, n42869, n42807,
    n42809, n42808, n42874, n42811, n42813, n42812, n42879, n42815, n42817,
    n42816, n42819, n42884, n42820, n42822, n42821, n42823, n42826, n42825,
    n42827, n42830, n42829, n42831, n42834, n42833, n42835, n42838, n42837,
    n42839, n42842, n42841, n42843, n42846, n42845, n42847, n42850, n42849,
    n42851, n42854, n42853, n42856, n42859, n42858, n42860, n42863, n42862,
    n42864, n42867, n42866, n42868, n42871, n42870, n42873, n42876, n42875,
    n42878, n42881, n42880, n42883, n42886, n42885, n42890, n42889, n42893,
    n42892, n42897, n42896, n42902, n42958, n42978, n42900, n42901, n42905,
    n42904, n42909, n42908, n42914, n42985, n42912, n42982, n42911, n42913,
    n42918, n42917, n42928, n43008, n42924, n42923, n42926, n42925, n42927,
    n42930, n43002, n43017, n42935, n42934, n42943, n42941, n43019, n42939,
    n42938, n42940, n42942, n42946, n42956, n43035, n42951, n43041, n42950,
    n42954, n42953, n42955, n42959, n42977, n42998, n42962, n42994, n42964,
    n43003, n42990, n42975, n42970, n42969, n42981, n42971, n42973, n42974,
    n42976, n42980, n42979, n42989, n42987, n42984, n42986, n42988, n42992,
    n42991, n42996, n42995, n42997, n43012, n42999, n43007, n43005, n43004,
    n43006, n43010, n43009, n43011, n43015, n43040, n43016, n43025, n43020,
    n43023, n43022, n43024, n43030, n43028, n43029, n43033, n43034, n43038,
    n43037, n43039, n43044, n43043, n43045, n43048, n44509, n43050, n43052,
    n44808, n43058, n43294, n43059, n43221, n43087, n43192, n43069, n43064,
    n43200, n43063, n44411, n44317, n43068, n43096, n44402, n43470, n43977,
    n43071, n43080, n43075, n43073, n43285, n43074, n43076, n43077, n43085,
    n43078, n43084, n43079, n43094, n43083, n43636, n43091, n44136, n43086,
    n43089, n43088, n43090, n43092, n43093, n43095, n43100, n43098, n43097,
    n43099, n43106, n43104, n43103, n44428, n43105, n43112, n43110, n43108,
    n43107, n44427, n43109, n43111, n43115, n44424, n43114, n43121, n43119,
    n43118, n44439, n43120, n43128, n44435, n43126, n43124, n43123, n44438,
    n43125, n43127, n43130, n43129, n43136, n43134, n43133, n44450, n43135,
    n43143, n44446, n43141, n43139, n43138, n44449, n43140, n43142, n43145,
    n43144, n43151, n43149, n43148, n44461, n43150, n43158, n44457, n43156,
    n43154, n43153, n44460, n43155, n43157, n43160, n43159, n43162, n43166,
    n43164, n43163, n44473, n43165, n43172, n43170, n43168, n43167, n44472,
    n43169, n43171, n43175, n44469, n43174, n43180, n43178, n43177, n44484,
    n43179, n43186, n43184, n43182, n43181, n44483, n43183, n43185, n43189,
    n44480, n43188, n44492, n43196, n43194, n43193, n44500, n43195, n43206,
    n44494, n43204, n43202, n43201, n44498, n43203, n43205, n43209, n43208,
    n43215, n43211, n43216, n43213, n43212, n43282, n43214, n43230, n43218,
    n43217, n43220, n43219, n43224, n43222, n43223, n43228, n43226, n43372,
    n43227, n43229, n43232, n43231, n43234, n43233, n43238, n43236, n43235,
    n43237, n43240, n43239, n43242, n43241, n43246, n43244, n43243, n43245,
    n43248, n43247, n43250, n43249, n43254, n43252, n43251, n43253, n43256,
    n43255, n43258, n43257, n43262, n43260, n43259, n43261, n43264, n43263,
    n43266, n43265, n43270, n43268, n43267, n43269, n43272, n43271, n43274,
    n43273, n43278, n43276, n43275, n43277, n43280, n43279, n43284, n43283,
    n43289, n43287, n43286, n43288, n43292, n43291, n43293, n43296, n43375,
    n43363, n43295, n43305, n43308, n43635, n43301, n43297, n43298, n43307,
    n43299, n43306, n43300, n43367, n43303, n43302, n43304, n43314, n43311,
    n43650, n43309, n43310, n43313, n43316, n43315, n43320, n43318, n43317,
    n43319, n43322, n43321, n43324, n43323, n43328, n43326, n43325, n43327,
    n43330, n43329, n43332, n43331, n43336, n43334, n43333, n43335, n43338,
    n43337, n43340, n43339, n43344, n43342, n43341, n43343, n43346, n43345,
    n43348, n43347, n43352, n43350, n43349, n43351, n43354, n43353, n43356,
    n43355, n43360, n43358, n43357, n43359, n43362, n43361, n43365, n43364,
    n43371, n43369, n43368, n43370, n43374, n43373, n43387, n43377, n43376,
    n43396, n43378, n43386, n43382, n43381, n43383, n43384, n43390, n43385,
    n43394, n43392, n43389, n43391, n43453, n43393, n43395, n43400, n43399,
    n43402, n43401, n43406, n43404, n43403, n43405, n43408, n43407, n43410,
    n43409, n43414, n43412, n43411, n43413, n43416, n43415, n43418, n43417,
    n43422, n43420, n43419, n43421, n43424, n43423, n43426, n43425, n43430,
    n43428, n43427, n43429, n43432, n43431, n43434, n43433, n43438, n43436,
    n43435, n43437, n43440, n43439, n43442, n43441, n43446, n43444, n43443,
    n43445, n43448, n43447, n43452, n43451, n43457, n43455, n43454, n43456,
    n43460, n43459, n43461, n43547, n43478, n43535, n43467, n44137, n43462,
    n43465, n43475, n43463, n43464, n43536, n43466, n43484, n43468, n43469,
    n44778, n43568, n43624, n43482, n43473, n43472, n43474, n43476, n43477,
    n43479, n43480, n43481, n43483, n43486, n43485, n43488, n43487, n43492,
    n43490, n43489, n43491, n43494, n43493, n43496, n43495, n43500, n43498,
    n43497, n43499, n43502, n43501, n43504, n43503, n43508, n43506, n43505,
    n43507, n43510, n43509, n43512, n43511, n43516, n43514, n43513, n43515,
    n43518, n43517, n43520, n43519, n43524, n43522, n43521, n43523, n43526,
    n43525, n43528, n43527, n43532, n43530, n43529, n43531, n43534, n43533,
    n43538, n43537, n43543, n43541, n43540, n43542, n43546, n43545, n43620,
    n43553, n43554, n43551, n43559, n43549, n43550, n43621, n43552, n43567,
    n43555, n43563, n43556, n43561, n43557, n43558, n43560, n43562, n43565,
    n43564, n43566, n43571, n43570, n43573, n43572, n43577, n43575, n43574,
    n43576, n43579, n43578, n43581, n43580, n43585, n43583, n43582, n43584,
    n43587, n43586, n43589, n43588, n43593, n43591, n43590, n43592, n43595,
    n43594, n43597, n43596, n43601, n43599, n43598, n43600, n43603, n43602,
    n43605, n43604, n43609, n43607, n43606, n43608, n43611, n43610, n43613,
    n43612, n43617, n43615, n43614, n43616, n43619, n43618, n43623, n43622,
    n43628, n43626, n43625, n43627, n43631, n43630, n43648, n43705, n43634,
    n43632, n43791, n43633, n43645, n43641, n43637, n43638, n43647, n43646,
    n43639, n43640, n43643, n43642, n43644, n43656, n43654, n43652, n43649,
    n43651, n43653, n43655, n43658, n43657, n43662, n43660, n43659, n43661,
    n43664, n43663, n43666, n43665, n43670, n43668, n43667, n43669, n43672,
    n43671, n43674, n43673, n43678, n43676, n43675, n43677, n43680, n43679,
    n43682, n43681, n43686, n43684, n43683, n43685, n43688, n43687, n43690,
    n43689, n43694, n43692, n43691, n43693, n43696, n43695, n43698, n43697,
    n43702, n43700, n43699, n43701, n43704, n43703, n43707, n43706, n43712,
    n43710, n43709, n43711, n43715, n43714, n43787, n43723, n44395, n43719,
    n43730, n43721, n43720, n43788, n43722, n43728, n43724, n43726, n43725,
    n43727, n43738, n43736, n43734, n43732, n43731, n43733, n43735, n43737,
    n43740, n43739, n43744, n43742, n43741, n43743, n43746, n43745, n43748,
    n43747, n43752, n43750, n43749, n43751, n43754, n43753, n43756, n43755,
    n43760, n43758, n43757, n43759, n43762, n43761, n43764, n43763, n43768,
    n43766, n43765, n43767, n43770, n43769, n43772, n43771, n43776, n43774,
    n43773, n43775, n43778, n43777, n43780, n43779, n43784, n43782, n43781,
    n43783, n43786, n43785, n43790, n43789, n43795, n43793, n43792, n43794,
    n43798, n43797, n44133, n43879, n43898, n43806, n43800, n43804, n43802,
    n43801, n43809, n43803, n43868, n43805, n43816, n44070, n43955, n43807,
    n43808, n43811, n43810, n43812, n43814, n43813, n43815, n43818, n43817,
    n43820, n43819, n43824, n43822, n43821, n43823, n43826, n43825, n43828,
    n43827, n43832, n43830, n43829, n43831, n43834, n43833, n43836, n43835,
    n43840, n43838, n43837, n43839, n43842, n43841, n43844, n43843, n43848,
    n43846, n43845, n43847, n43850, n43849, n43852, n43851, n43856, n43854,
    n43853, n43855, n43858, n43857, n43860, n43859, n43864, n43862, n43861,
    n43863, n43866, n43865, n43870, n43869, n43875, n43873, n43872, n43874,
    n43878, n43877, n43886, n43884, n44223, n43894, n43881, n43882, n43883,
    n43952, n43885, n43891, n43887, n44039, n43889, n43888, n43890, n43902,
    n43896, n43893, n43895, n43897, n43900, n43899, n43901, n43904, n43903,
    n43908, n43906, n43905, n43907, n43910, n43909, n43912, n43911, n43916,
    n43914, n43913, n43915, n43918, n43917, n43920, n43919, n43924, n43922,
    n43921, n43923, n43926, n43925, n43928, n43927, n43932, n43930, n43929,
    n43931, n43934, n43933, n43936, n43935, n43940, n43938, n43937, n43939,
    n43942, n43941, n43944, n43943, n43948, n43946, n43945, n43947, n43950,
    n43949, n43954, n43953, n43959, n43957, n43956, n43958, n43962, n43961,
    n43965, n43963, n44058, n43971, n44038, n43964, n43987, n43966, n43968,
    n43979, n43980, n43974, n43970, n44323, n43972, n43973, n43975, n43985,
    n43978, n44309, n43983, n43981, n43982, n43984, n43986, n43989, n43988,
    n43991, n43990, n43995, n43993, n43992, n43994, n43997, n43996, n43999,
    n43998, n44003, n44001, n44000, n44002, n44005, n44004, n44007, n44006,
    n44011, n44009, n44008, n44010, n44013, n44012, n44015, n44014, n44019,
    n44017, n44016, n44018, n44021, n44020, n44023, n44022, n44027, n44025,
    n44024, n44026, n44029, n44028, n44031, n44030, n44035, n44033, n44032,
    n44034, n44037, n44036, n44041, n44040, n44046, n44044, n44043, n44045,
    n44049, n44048, n44050, n44121, n44057, n44055, n44053, n44052, n44060,
    n44054, n44122, n44056, n44068, n44059, n44064, n44762, n44062, n44061,
    n44063, n44066, n44065, n44067, n44072, n44069, n44071, n44074, n44073,
    n44078, n44076, n44075, n44077, n44080, n44079, n44082, n44081, n44086,
    n44084, n44083, n44085, n44088, n44087, n44090, n44089, n44094, n44092,
    n44091, n44093, n44096, n44095, n44098, n44097, n44102, n44100, n44099,
    n44101, n44104, n44103, n44106, n44105, n44110, n44108, n44107, n44109,
    n44112, n44111, n44114, n44113, n44118, n44116, n44115, n44117, n44120,
    n44119, n44124, n44123, n44128, n44126, n44125, n44127, n44131, n44130,
    n44240, n44155, n44211, n44135, n44761, n44134, n44149, n44310, n44145,
    n44139, n44140, n44141, n44151, n44143, n44312, n44150, n44144, n44147,
    n44146, n44148, n44162, n44159, n44154, n44157, n44156, n44158, n44160,
    n44161, n44164, n44163, n44168, n44166, n44165, n44167, n44170, n44169,
    n44172, n44171, n44176, n44174, n44173, n44175, n44178, n44177, n44180,
    n44179, n44184, n44182, n44181, n44183, n44186, n44185, n44188, n44187,
    n44192, n44190, n44189, n44191, n44194, n44193, n44196, n44195, n44200,
    n44198, n44197, n44199, n44202, n44201, n44204, n44203, n44208, n44206,
    n44205, n44207, n44210, n44209, n44213, n44212, n44219, n44217, n44216,
    n44218, n44222, n44221, n44229, n44396, n44225, n44224, n44236, n44227,
    n44226, n44295, n44228, n44235, n44231, n44386, n44233, n44232, n44234,
    n44245, n44238, n44237, n44239, n44243, n44241, n44242, n44244, n44247,
    n44246, n44251, n44249, n44248, n44250, n44253, n44252, n44255, n44254,
    n44259, n44257, n44256, n44258, n44261, n44260, n44263, n44262, n44267,
    n44265, n44264, n44266, n44269, n44268, n44271, n44270, n44275, n44273,
    n44272, n44274, n44277, n44276, n44279, n44278, n44283, n44281, n44280,
    n44282, n44285, n44284, n44287, n44286, n44291, n44289, n44288, n44290,
    n44293, n44292, n44297, n44296, n44302, n44300, n44299, n44301, n44305,
    n44304, n44417, n44316, n44314, n44319, n44313, n44383, n44315, n44331,
    n44329, n44318, n44320, n44321, n44322, n44325, n44324, n44328, n44330,
    n44333, n44332, n44335, n44334, n44339, n44337, n44336, n44338, n44341,
    n44340, n44343, n44342, n44347, n44345, n44344, n44346, n44349, n44348,
    n44351, n44350, n44355, n44353, n44352, n44354, n44357, n44356, n44359,
    n44358, n44363, n44361, n44360, n44362, n44365, n44364, n44367, n44366,
    n44371, n44369, n44368, n44370, n44373, n44372, n44375, n44374, n44379,
    n44377, n44376, n44378, n44381, n44380, n44385, n44384, n44390, n44388,
    n44387, n44389, n44393, n44392, n44404, n44398, n44397, n44412, n44401,
    n44400, n44493, n44403, n44410, n44408, n44407, n44409, n44423, n44414,
    n44413, n44416, n44421, n44419, n44420, n44422, n44426, n44425, n44432,
    n44430, n44429, n44431, n44434, n44433, n44437, n44436, n44443, n44441,
    n44440, n44442, n44445, n44444, n44448, n44447, n44454, n44452, n44451,
    n44453, n44456, n44455, n44459, n44458, n44465, n44463, n44462, n44464,
    n44467, n44466, n44471, n44470, n44477, n44475, n44474, n44476, n44479,
    n44478, n44482, n44481, n44488, n44486, n44485, n44487, n44490, n44489,
    n44496, n44495, n44504, n44502, n44501, n44503, n44507, n44506, n44806,
    n44511, n44513, n44516, n44518, n44520, n44533, n44525, n44524, n44526,
    n44527, n44529, n44541, n44528, n44531, n44538, n44532, n44534, n44535,
    n44536, n44537, n44539, n44545, n44542, n44543, n44544, n44548, n44547,
    n44550, n44549, n44553, n44552, n44555, n44554, n44561, n44558, n44557,
    n44560, n44559, n44563, n44562, n44565, n44564, n44568, n44567, n44570,
    n44569, n44573, n44572, n44575, n44574, n44580, n44581, n44578, n44577,
    n44579, n44583, n44582, n44585, n44584, n44588, n44587, n44590, n44589,
    n44593, n44592, n44595, n44594, n44599, n44598, n44601, n44600, n44604,
    n44603, n44606, n44605, n44608, n44607, n44610, n44609, n44613, n44612,
    n44615, n44614, n44618, n44617, n44620, n44619, n44623, n44626, n44622,
    n44625, n44624, n44630, n44631, n44628, n44627, n44629, n44633, n44632,
    n44635, n44634, n44638, n44637, n44640, n44639, n44643, n44642, n44645,
    n44644, n44648, n44647, n44650, n44649, n44653, n44656, n44652, n44655,
    n44654, n44658, n44657, n44660, n44659, n44663, n44662, n44665, n44664,
    n44668, n44667, n44670, n44669, n44673, n44672, n44675, n44674, n44678,
    n44677, n44680, n44679, n44683, n44682, n44685, n44684, n44690, n44688,
    n44687, n44689, n44695, n44693, n44694, n44697, n44696, n44699, n44698,
    n44701, n44700, n44703, n44702, n44705, n44704, n44708, n44707, n44710,
    n44715, n44714, n44716, n44718, n44717, n44731, n44720, n44725, n44723,
    n44733, n44734, n44722, n44724, n44726, n44728, n44727, n44730, n44739,
    n44737, n44735, n44736, n44738, n44740, n44743, n44742, n44746, n44747,
    n44759, n44752, n44751, n44755, n44754, n44756, n44758, n44774, n44763,
    n44764, n44771, n44790, n44769, n44802, n44768, n44770, n44772, n44773,
    n44776, n44777, n44783, n44779, n44780, n44782, n44786, n44785, n44787,
    n44789, n44788, n44794, n44793, n44796, n44795, n44797, n44799, n44798,
    n44804, n44803, n44805, n44807, n44811, n44810, n44822, n44819, n44824,
    n44817, n44816, n44818, n44820, n44825, n44821, n44827, n44826, n44830,
    n44829, n44834, n44833, n44836, n44840, n44839, n44856, n44858, n44844,
    n44847, n44846, n44848, n44849, n44852, n44854, n44855, n44857, n44861,
    n44860, n34993, n36497, n23304, n37463, n30741, n44863, n44864, n44865,
    n30615;
  assign n43871 = n43724;
  assign n36151 = n24284 & P3_INSTADDRPOINTER_REG_27__SCAN_IN;
  assign n41228 = ~n42139 | ~n42177;
  assign n41686 = ~n41786;
  assign n43067 = ~n44317 & ~n44230;
  assign n43398 = ~n43397 & ~n44230;
  assign n40820 = n40755 & n42177;
  assign n41751 = ~n41590 | ~n42177;
  assign n25837 = ~n25677 | ~n44514;
  assign n23180 = ~n23407 | ~n28071;
  assign n32932 = n28669 & n23026;
  assign n38758 = ~n37190;
  assign n41418 = n27896;
  assign n23864 = n39660 | n39659;
  assign n29891 = n28555;
  assign n24634 = ~n37502;
  assign n37494 = ~n24625;
  assign n37473 = ~n24448 & ~n24447;
  assign n37482 = ~n24356 & ~n24355;
  assign n28494 = n27677 & n27622;
  assign n27817 = n29739 & n29098;
  assign n42760 = n25043;
  assign n26866 = ~n26035;
  assign n29581 = ~n23145 | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n22838 = ~n25652;
  assign n35412 = ~n24522;
  assign n28734 = ~n23277;
  assign n29753 = n27409;
  assign n43161 = n25004;
  assign n39805 = n27610;
  assign n24802 = ~n24785 & ~n24784;
  assign n26630 = ~n24815;
  assign n24898 = n24763 & n31461;
  assign n24936 = ~n31449 & ~n31474;
  assign n24734 = ~n31449;
  assign n29002 = ~n29086 & ~n23875;
  assign n40303 = ~P2_PHYADDRPOINTER_REG_2__SCAN_IN ^ P2_PHYADDRPOINTER_REG_1__SCAN_IN;
  assign n22818 = ~n41894;
  assign n22819 = ~n22818;
  assign n22820 = ~n22818;
  assign n22822 = ~n39019;
  assign n22823 = ~n39019;
  assign n22825 = ~n44863;
  assign n28500 = n39849 & n42208;
  assign n25085 = n24759 & n31461;
  assign n38721 = n38788 | n39045;
  assign n26859 = ~n25267;
  assign n27880 = n27879 & n23062;
  assign n28283 = ~n31598;
  assign n23627 = n23304 & n23446;
  assign n27665 = ~n28494 | ~P2_STATE2_REG_0__SCAN_IN;
  assign n24721 = ~n37494 | ~n24634;
  assign n24668 = ~n37473 & ~n34971;
  assign n24116 = ~n24564 ^ n35782;
  assign n24010 = ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n28596 = ~n40552 | ~n42196;
  assign n28669 = ~n33027;
  assign n28586 = ~n23864 | ~n28574;
  assign n24598 = n24665 | n24721;
  assign n38695 = ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN;
  assign n24188 = ~n24564 | ~n35782;
  assign n38757 = ~n38696;
  assign n30957 = ~n30970 | ~n25946;
  assign n28980 = n28580;
  assign n39627 = ~n28586 ^ n28587;
  assign n41785 = ~n41002;
  assign n24522 = ~n38740 | ~n38695;
  assign n22828 = n37190;
  assign n35252 = n24373;
  assign n42461 = ~n31415;
  assign n44298 = ~n44761 & ~n44801;
  assign n31658 = ~n31650 & ~n31649;
  assign n23244 = ~n27740 | ~n28331;
  assign n23178 = n23195 & n29053;
  assign n23222 = ~n23428 | ~n28303;
  assign n40560 = ~n40637;
  assign n27656 = n27607;
  assign n34384 = ~n34459;
  assign n34430 = ~n34405;
  assign n24625 = ~n24387 & ~n24386;
  assign n22837 = ~n23280;
  assign n40729 = n40580 | n41491;
  assign n41878 = ~n41757;
  assign n34470 = ~n34448;
  assign n34971 = ~n24480 & ~n24479;
  assign n36662 = n24583 ^ n24582;
  assign n37453 = ~n24512 & ~n24511;
  assign n39110 = ~n24551 & ~n24550;
  assign n43042 = ~n43018;
  assign n39820 = ~n29903 ^ n23960;
  assign n42177 = ~n41491;
  assign n32726 = ~n32290 & ~n22837;
  assign n34631 = ~n24292;
  assign n22826 = n24759 & n23602;
  assign n22827 = n27742 & n23206;
  assign n26986 = n24769 | n24768;
  assign n23702 = n23490 & n23703;
  assign n27631 = ~n27208 | ~n27209;
  assign n30654 = n23323 & n30664;
  assign n30851 = ~n30850 & ~n30864;
  assign n26482 = n24738 | n24754;
  assign n28126 = n28114 | n23907;
  assign n27908 = n23614 & n27757;
  assign n30676 = n23505 & n22910;
  assign n22964 = n23472 & n28305;
  assign n31700 = ~n31701 & ~n31702;
  assign n23126 = ~n23128 & ~n23127;
  assign n27900 = n27775 & n27774;
  assign n31974 = n28542;
  assign n23515 = ~n23511 | ~n23516;
  assign n27610 = ~n27613;
  assign n37190 = ~n33788 & ~n24627;
  assign n27163 = ~n27162 & ~n27161;
  assign n27162 = n23088 | n23089;
  assign n42961 = n43013 | n43031;
  assign n23690 = ~n28328 ^ n27735;
  assign n25235 = ~n23835 | ~n25188;
  assign n22829 = n24759 & n31461;
  assign n28298 = ~n23175 | ~n27880;
  assign n24763 = ~n24738;
  assign n24738 = ~n25183 | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN;
  assign n28309 = ~n23108 | ~n23472;
  assign n22830 = n35571;
  assign n36515 = n23774 & n23773;
  assign n25555 = ~n30825 & ~n25554;
  assign n34525 = ~n23643 | ~n23642;
  assign n22832 = n26806;
  assign n22833 = n26806;
  assign n26806 = ~n24734 | ~n24753;
  assign n36767 = ~n36201 & ~n36781;
  assign n34447 = ~P3_EBX_REG_0__SCAN_IN & ~P3_EBX_REG_1__SCAN_IN;
  assign n33747 = ~n24678 & ~n24603;
  assign n37008 = ~n36463 & ~n24628;
  assign n22834 = n38696;
  assign n38696 = ~n38732 & ~n24644;
  assign n27742 = ~n23978 | ~n27741;
  assign n23181 = ~n23266;
  assign n23438 = ~n32482;
  assign n23269 = ~n28302 | ~n28301;
  assign n32526 = ~n23389 | ~n22913;
  assign n23493 = n23331 & n30706;
  assign n23331 = ~n23622 | ~n23739;
  assign n43892 = n44070 | n43066;
  assign n22835 = ~n42413;
  assign n30950 = ~n23321 | ~n25502;
  assign n25883 = ~n23288 | ~n25920;
  assign n23091 = n27885 & n27884;
  assign n27884 = n27883 | n40513;
  assign n27781 = n27882 | n40452;
  assign n42932 = ~n31517 | ~n44514;
  assign n25411 = ~n23671 | ~n23669;
  assign n25393 = ~n23332 | ~n25175;
  assign n28174 = ~n28154 | ~n23576;
  assign n27715 = ~n27745 | ~n27744;
  assign n25030 = n25029 & n25028;
  assign n29831 = ~n28071;
  assign n37514 = ~n34971;
  assign n25054 = n25009;
  assign n23706 = ~n40471;
  assign n25009 = ~n24802 | ~n24801;
  assign n24927 = ~n24926 & ~n24925;
  assign n22836 = ~n27607;
  assign n40437 = ~P2_ADDRESS_REG_29__SCAN_IN | ~n27045;
  assign n22841 = n24898;
  assign n24315 = ~n34525;
  assign n27510 = n29761 & n29098;
  assign n29761 = ~n29731;
  assign n24815 = ~n31445 | ~n24764;
  assign n25089 = n23602 & n24764;
  assign n27348 = ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n29861 = n23463 & n22948;
  assign n23335 = ~n29069 ^ n29068;
  assign n23662 = ~n29027 ^ P2_INSTADDRPOINTER_REG_20__SCAN_IN;
  assign n32829 = ~n23462 ^ n23054;
  assign n23179 = n23188 & n32197;
  assign n23295 = ~n23522 | ~n23521;
  assign n32321 = ~n23270 | ~n29070;
  assign n23465 = n23636 & n22935;
  assign n32613 = ~n32197 ^ P2_INSTADDRPOINTER_REG_30__SCAN_IN;
  assign n32750 = n23503 & n23502;
  assign n23462 = ~n23946 | ~n32432;
  assign n32197 = ~n23181 | ~n23937;
  assign n23522 = n23524 & n23523;
  assign n32212 = ~n23181 | ~n23081;
  assign n32898 = ~n23273 ^ n32456;
  assign n32200 = ~n23481 | ~n23467;
  assign n30663 = ~n23323 | ~n30652;
  assign n32186 = n23852 & n32199;
  assign n32433 = n23663 & n23666;
  assign n29029 = ~n22873 | ~n22932;
  assign n30889 = ~n30261 | ~n30237;
  assign n23443 = n23269 & n22943;
  assign n30657 = ~n29935 & ~n29934;
  assign n23422 = n23178 & n23641;
  assign n31971 = ~n23520 ^ n23074;
  assign n23520 = ~n23519 | ~n23258;
  assign n30687 = ~n29971 & ~n29970;
  assign n26908 = n23847 & n23466;
  assign n23195 = ~n23617 | ~n23745;
  assign n38806 = P3_STATE2_REG_0__SCAN_IN & n23115;
  assign n30791 = n27060 & n27059;
  assign n30665 = ~n29967 ^ n29949;
  assign n23847 = ~n29991 & ~n23021;
  assign n23115 = n38805 | n38817;
  assign n29991 = ~n26661 | ~n26660;
  assign n44042 = ~n43983 | ~n43982;
  assign n43366 = ~n43976 | ~n43312;
  assign n32524 = ~n23425 | ~n23424;
  assign n32634 = ~n31703 | ~n31704;
  assign n23425 = n23427 & n23426;
  assign n23695 = n28016 & n28071;
  assign n41399 = ~n41342 | ~n41341;
  assign n23338 = n23339 & n23486;
  assign n29842 = ~n22869 & ~n31699;
  assign n38790 = ~n38787 & ~n38786;
  assign n23407 = ~n28300;
  assign n28305 = n28300;
  assign n23340 = n22870 & n23341;
  assign n23326 = n23327 & n23330;
  assign n41329 = n41323 & n23100;
  assign n28300 = ~n28298 ^ n28070;
  assign n28070 = ~n27946 | ~n27945;
  assign n31810 = ~n31832 & ~n31831;
  assign n36191 = n36215 & n23202;
  assign n23588 = n23589 & n23942;
  assign n22905 = ~n44070 & ~n43966;
  assign n35514 = ~n35537 & ~n36013;
  assign n30899 = ~n30926 | ~P1_INSTADDRPOINTER_REG_10__SCAN_IN;
  assign n29810 = n29809 & n32227;
  assign n42391 = n42469 & P1_STATE2_REG_2__SCAN_IN;
  assign n27844 = ~n23125 | ~n28575;
  assign n42413 = n42469 & n29916;
  assign n41310 = ~n41232;
  assign n41479 = ~n41400;
  assign n42960 = ~n42961;
  assign n42446 = ~n42444 | ~n42443;
  assign n25916 = n25384 & n23271;
  assign n23664 = n23379 & n23945;
  assign n42400 = n25907 & n25906;
  assign n30826 = n30844 | n30864;
  assign n43102 = ~n43191 & ~n43101;
  assign n43117 = ~n43191 & ~n43116;
  assign n23484 = n28228 & n32277;
  assign n30878 = n30903 & n30907;
  assign n43132 = ~n43191 & ~n43131;
  assign n33204 = n33200 | n33199;
  assign n27877 = n27859 & n27860;
  assign n26954 = ~n42625 & ~n26953;
  assign n26956 = ~n42625 & ~n26955;
  assign n43147 = ~n43191 & ~n43146;
  assign n29813 = n28231 & n28230;
  assign n30883 = n30953 | n31261;
  assign n42631 = ~n42630 & ~n43057;
  assign n41411 = n41321 | n41490;
  assign n41788 = n42140 | n41490;
  assign n42625 = ~n26922 | ~n44514;
  assign n30908 = n30953 | n31286;
  assign n41242 = n41490 | n41155;
  assign n23321 = n23470 | n23322;
  assign n36832 = ~n36881 & ~n24596;
  assign n41490 = n39621;
  assign n42443 = n42459 & n42458;
  assign n23397 = ~n23415 | ~n29335;
  assign n23090 = n27888 & n27887;
  assign n27887 = n40657 | n27916;
  assign n29805 = n31746 | n28071;
  assign n39335 = ~n39673;
  assign n42937 = n42932 & n30635;
  assign n40657 = n27886;
  assign n32254 = n31790 | n28071;
  assign n27780 = n27886 | n29426;
  assign n39620 = ~n29330 ^ n29328;
  assign n42153 = n42156 & n42170;
  assign n40577 = n23692 & n23693;
  assign n27956 = n27900;
  assign n27767 = n27904 | n29222;
  assign n31689 = ~n32201 & ~n31713;
  assign n42076 = ~n33142 & ~n33141;
  assign n23743 = ~n23136 | ~n23282;
  assign n29326 = ~n22883 | ~n23049;
  assign n23446 = ~n23510 | ~n23508;
  assign n39636 = n31958 & n29319;
  assign n23669 = ~n23670 | ~n22912;
  assign n31954 = n29314 & n29319;
  assign n25859 = n25182 & n25550;
  assign n44767 = ~n31431 ^ n23621;
  assign n25868 = ~n25393 ^ n25392;
  assign n22848 = ~n23206 & ~n22847;
  assign n31955 = n29318 & n29317;
  assign n23926 = n43210 & n44851;
  assign n28145 = n28154 & n28155;
  assign n27723 = ~n27718 | ~n27715;
  assign n23904 = n28114 | n23906;
  assign n28154 = ~n28166 & ~n28160;
  assign n39588 = n33094 | n33093;
  assign n24582 = ~n23172 | ~n24581;
  assign n23350 = ~n23349 & ~n23572;
  assign n27732 = n27735 | n27734;
  assign n23349 = n22865 | n28164;
  assign n23867 = ~n23869 & ~n23868;
  assign n34002 = ~P3_EBX_REG_21__SCAN_IN & ~n34021;
  assign n34376 = n34320;
  assign n26568 = ~n26399 & ~n30767;
  assign n23359 = ~n33747 | ~n24667;
  assign n38797 = ~n24604 | ~n24632;
  assign n27729 = ~n23243 | ~n23293;
  assign n26526 = ~n26439 & ~n30792;
  assign n23675 = n25833 & n23676;
  assign n27695 = ~n27694 & ~n27693;
  assign n27688 = n27687 & n27686;
  assign n29843 = ~n28318;
  assign n25833 = ~n23677 | ~n25678;
  assign n23725 = n25048 & n23728;
  assign n25048 = n22879 & n25007;
  assign n23930 = n25024 & n25026;
  assign n23724 = n23727 & n25693;
  assign n27549 = n27449 & n27448;
  assign n24617 = n24673 & n37463;
  assign n23903 = ~n27616 | ~n22956;
  assign n23117 = n23118 | P2_STATE2_REG_0__SCAN_IN;
  assign n34116 = ~P3_EBX_REG_15__SCAN_IN & ~n34128;
  assign n28242 = n23375 & n28054;
  assign n23727 = n31438 & n25691;
  assign n23728 = ~n25668 | ~n31568;
  assign n36610 = n33408 & n33284;
  assign n27677 = n27635 & n23137;
  assign n39443 = ~n39453 & ~n39444;
  assign n25822 = ~n27579;
  assign n25629 = ~n25645;
  assign n25660 = ~n25669 | ~n25023;
  assign n23234 = n23950 & n27445;
  assign n28575 = ~n27809 | ~n27808;
  assign n28512 = n28261 & n39805;
  assign n27579 = n25055;
  assign n22839 = ~n25041;
  assign n25645 = n25462 & n25243;
  assign n25669 = ~n25053;
  assign n25001 = ~n25000 & ~n25661;
  assign n28601 = n27482 & n27481;
  assign n24187 = n35773 | n35761;
  assign n26914 = ~n25014 | ~n25008;
  assign n25601 = n25609 & n42760;
  assign n31502 = n25004 & n25017;
  assign n25462 = ~n25134;
  assign n25639 = ~n25619 & ~n43146;
  assign n23537 = ~n24080 ^ P3_INSTADDRPOINTER_REG_2__SCAN_IN;
  assign n33802 = ~n36229 & ~n36231;
  assign n25055 = ~n25043 | ~n25054;
  assign n25042 = n25018;
  assign n43131 = n25008;
  assign n28498 = ~n23369 & ~n27614;
  assign n24865 = ~n26986 & ~n25054;
  assign n28595 = n27443 & n27442;
  assign n25008 = ~n25009;
  assign n35773 = n24150 & n24149;
  assign n25661 = ~n25014 | ~n25009;
  assign n43057 = ~n26986;
  assign n25011 = ~n25017 | ~n25609;
  assign n39593 = n27531;
  assign n42209 = ~n40444 | ~P2_STATE2_REG_0__SCAN_IN;
  assign n43116 = n25014;
  assign n43146 = n25017;
  assign n28552 = ~n40519;
  assign n43101 = ~n25043;
  assign n35753 = ~n22918 | ~n24218;
  assign n25017 = n24897 & n24896;
  assign n25609 = ~n24927 | ~n24928;
  assign n40501 = n27277;
  assign n33538 = ~U214;
  assign n27531 = ~n27536;
  assign n24569 = n24018 | n24017;
  assign n24149 = n24148 & n24147;
  assign n40471 = n27619;
  assign n40444 = n27536;
  assign n24897 = n24879 & n24878;
  assign n22840 = n27612;
  assign n27208 = ~n27207 | ~n27206;
  assign n24801 = n24800 & n24799;
  assign n24928 = n24910 & n23734;
  assign n23227 = n23229 & n23228;
  assign n27209 = ~n27192 | ~n27191;
  assign n24925 = ~n24924 | ~n24923;
  assign n24783 = n24779 & n24778;
  assign n24893 = n24889 & n24888;
  assign n24924 = n24920 & n24919;
  assign n24851 = n24849 & n24848;
  assign n29575 = ~n29660 | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n29580 = ~n29660 | ~n29098;
  assign n33147 = ~n23569 | ~n29098;
  assign n41894 = ~n42070;
  assign n27045 = n27044 | n27043;
  assign n22842 = ~n31463;
  assign n24923 = n24922 & n24921;
  assign n24513 = n34578;
  assign n24300 = n24006 & n24005;
  assign n24292 = n24006 & n24009;
  assign n27319 = n27317 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n24972 = n24936;
  assign n24973 = ~n24815;
  assign n24989 = ~n24905;
  assign n25065 = ~n24765 | ~n24763;
  assign n25118 = n24765 & n24764;
  assign n27379 = n27377 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n27334 = n27332 & n29098;
  assign n42024 = ~P2_STATE_REG_2__SCAN_IN | ~n42224;
  assign n41158 = ~n41089 & ~n41575;
  assign n27218 = n27216 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n27228 = n27226 & n29098;
  assign n36653 = ~n34343 & ~n36665;
  assign n29752 = ~n29718;
  assign n44597 = ~n44859 | ~n44546;
  assign n44691 = ~P1_STATE_REG_2__SCAN_IN | ~n44859;
  assign n22843 = ~n37197;
  assign n23065 = n24000 & n23758;
  assign n24005 = ~n38728;
  assign n24006 = ~n23999;
  assign n22844 = ~n24301;
  assign n24318 = n34451 & n23987;
  assign n44835 = ~n44508 & ~P1_STATE2_REG_0__SCAN_IN;
  assign n23758 = ~n23759 & ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN;
  assign n31657 = ~n31652 & ~n31651;
  assign n38728 = ~n34395 | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n23999 = ~n38709 | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN;
  assign n25912 = ~n25903 & ~n25902;
  assign n25196 = n24764 & n31461;
  assign n31445 = n23834 & P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n31449 = ~n25574 | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n24753 = n25614 & P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign n31651 = ~P2_PHYADDRPOINTER_REG_2__SCAN_IN | ~P2_PHYADDRPOINTER_REG_1__SCAN_IN;
  assign n25614 = ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN;
  assign n42196 = ~P2_STATE2_REG_3__SCAN_IN;
  assign n38719 = ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n42134 = P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN;
  assign n34451 = ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN & ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign n38709 = ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign n34395 = ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n24000 = ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN & ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n22845 = n23106;
  assign n22846 = ~n23407 | ~P2_INSTADDRPOINTER_REG_5__SCAN_IN;
  assign n33342 = ~n36107 & ~n36109;
  assign n22847 = ~n33176;
  assign n27886 = ~n23692 | ~n22848;
  assign n23692 = ~n23639;
  assign n41782 = n27908;
  assign n27412 = ~n27428 | ~n27348;
  assign n30257 = ~n23841 | ~n23840;
  assign n22849 = n23120 & n27947;
  assign n23630 = ~n23224 & ~n23631;
  assign n27779 = ~n23639 & ~n23206;
  assign n24253 = ~n24255 ^ n23754;
  assign n23128 = n27771 | n27782;
  assign n23189 = ~n23696;
  assign n29739 = ~n27418;
  assign n23932 = ~n28299 & ~n23933;
  assign n36297 = ~n36333 | ~n24273;
  assign n26899 = ~n26842 & ~n30666;
  assign n23569 = n22863;
  assign n31670 = ~n31625 & ~n31626;
  assign n31668 = ~n31630 & ~n31629;
  assign n31662 = ~n31642 & ~n31641;
  assign n27121 = n27412 | n29669;
  assign n27245 = n27412 | n29116;
  assign n27195 = n27412 | n40482;
  assign n27149 = n27412 | n29576;
  assign n27184 = n27412 | n29283;
  assign n27213 = n27412 | n29749;
  assign n27136 = n27412 | n40513;
  assign n22850 = ~n25382 | ~n25381;
  assign n23101 = ~n22850 | ~n22851;
  assign n22851 = n23103 & n23271;
  assign n22852 = n23671 & n23669;
  assign n22853 = ~n23835 | ~n25188;
  assign n22854 = n30695;
  assign n22855 = n23505;
  assign n23505 = ~n25559 | ~n23331;
  assign n29588 = n27119 & n27570;
  assign n27747 = n27744;
  assign n31012 = ~n25431 | ~n25430;
  assign n39380 = ~n39396 & ~n39394;
  assign n22856 = ~n42120;
  assign n22857 = ~n23276;
  assign n22858 = ~n22857;
  assign n42120 = P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign n23194 = n27743 & n22859;
  assign n22859 = n27742 & n40343;
  assign n23271 = ~n23445 | ~n23304;
  assign n23696 = ~n23501 | ~n28016;
  assign n24861 = ~n24853 & ~n24852;
  assign n31431 = ~n22853 | ~n25234;
  assign n22860 = ~n40552 | ~n42196;
  assign n39637 = ~n29326 ^ n29324;
  assign n23174 = ~n32562 | ~P2_INSTADDRPOINTER_REG_6__SCAN_IN;
  assign n32305 = ~n32482 & ~n23618;
  assign n22862 = ~n25065;
  assign n27509 = n29761 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n30684 = ~n30682 & ~n30681;
  assign n31663 = ~n31639 & ~n31640;
  assign n43065 = ~n23496 | ~n25424;
  assign n23299 = ~n25035 ^ n25187;
  assign n23280 = ~n23190 | ~n23422;
  assign n43379 = ~n23785 ^ n25139;
  assign n22863 = ~n33146;
  assign n22864 = ~n33146;
  assign n33146 = ~n27119 | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n31665 = ~n31635 & ~n31636;
  assign n31667 = ~n31631 & ~n31632;
  assign n31669 = ~n31627 & ~n31628;
  assign n31659 = ~n31648 & ~n31647;
  assign n31660 = ~n31646 & ~n31645;
  assign n31661 = ~n31644 & ~n31643;
  assign n23275 = n23638 & n23344;
  assign n25232 = n25231 & n25230;
  assign n25648 = n23606 & n23604;
  assign n25642 = ~P1_STATE2_REG_0__SCAN_IN & ~n31528;
  assign n25243 = ~n43146 | ~P1_STATE2_REG_0__SCAN_IN;
  assign n23916 = ~n28149 & ~n23917;
  assign n23341 = ~n23588 | ~n23343;
  assign n23343 = ~n23699;
  assign n29320 = ~n29331 | ~n42196;
  assign n23445 = n23446 & n23001;
  assign n28347 = n27647 & n27646;
  assign n23482 = ~n29810;
  assign n23819 = ~n23381;
  assign n23722 = n32292 & n32307;
  assign n23860 = n28183 & n32454;
  assign n28835 = ~n32902;
  assign n23388 = ~n23180 | ~n23430;
  assign n29319 = ~n23686 | ~n23684;
  assign n23684 = ~n22942 & ~n23685;
  assign n23685 = ~n27672;
  assign n23774 = ~n23203 | ~n23772;
  assign n23772 = n24256 & n22930;
  assign n23840 = n30323 & n23842;
  assign n23816 = n29972 | n29950;
  assign n31420 = ~n31508 & ~n27053;
  assign n43051 = ~n25650 | ~n25649;
  assign n23506 = n23331 & n22952;
  assign n23141 = n23185 & n23187;
  assign n25778 = ~n30199;
  assign n43056 = ~n43471;
  assign n32931 = ~n32932 | ~n32933;
  assign n28344 = ~n39580;
  assign n23262 = ~n23264 | ~n23263;
  assign n23945 = n32402 & n32432;
  assign n23481 = n23478 & n29817;
  assign n23478 = n23719 | n23482;
  assign n23896 = ~n31928 & ~n23019;
  assign n23897 = ~n29072;
  assign n34483 = ~n38689 & ~n27587;
  assign n34320 = P3_PHYADDRPOINTER_REG_31__SCAN_IN ^ n33288;
  assign n36384 = ~n36408 & ~n36405;
  assign n23147 = n43051;
  assign n25677 = ~n25676 | ~n25675;
  assign n25675 = n23310 & n31423;
  assign n29896 = ~n28580;
  assign n23253 = n23012 & n23254;
  assign n23254 = ~n32457;
  assign n31896 = n23517 | n23402;
  assign n32441 = ~n32458 & ~n32457;
  assign n32537 = ~n32564 | ~n23245;
  assign n23245 = ~n32549 & ~n23246;
  assign n23246 = ~n32563;
  assign n29013 = n28282 & n39160;
  assign n23450 = n23452 & n23451;
  assign n25616 = ~n25637 | ~n25613;
  assign n23594 = n41503 & P2_INSTQUEUE_REG_12__5__SCAN_IN;
  assign n24765 = ~n31449;
  assign n23183 = ~n25085 | ~P1_INSTQUEUE_REG_3__5__SCAN_IN;
  assign n23777 = ~n25232;
  assign n23781 = ~n25232 & ~n23782;
  assign n23778 = ~n22982 | ~n23779;
  assign n23779 = ~n25232 | ~n25229;
  assign n23780 = ~n23782 & ~n44851;
  assign n25107 = n25105 | n25104;
  assign n24813 = ~n24812 & ~n24811;
  assign n24814 = ~n23582 & ~n23580;
  assign n23580 = ~n24803 & ~n23581;
  assign n25426 = n25275 | n25274;
  assign n25414 = n25228 & n25227;
  assign n23834 = ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n23906 = n23907 | n28127;
  assign n23907 = n23040 | n28115;
  assign n23374 = ~n28242;
  assign n23395 = n27646 & P2_REIP_REG_2__SCAN_IN;
  assign n28142 = n28552 & P2_EBX_REG_18__SCAN_IN;
  assign n23912 = ~n23036;
  assign n23920 = ~n29753 | ~n23918;
  assign n23918 = n29098 & P2_INSTQUEUE_REG_6__2__SCAN_IN;
  assign n27498 = n29577 | n29558;
  assign n29497 = ~P2_INSTQUEUE_REG_8__2__SCAN_IN;
  assign n23231 = ~n31598 & ~n23232;
  assign n23232 = ~n27551;
  assign n38775 = ~n38774 & ~n38773;
  assign n23392 = ~n23494 & ~n30980;
  assign n23470 = ~n23271 | ~n25464;
  assign n23186 = ~n25506 | ~n25505;
  assign n25646 = n25648 | n25644;
  assign n25457 = ~n25499;
  assign n23491 = n23492 & n31010;
  assign n25424 = ~n23507 | ~n25278;
  assign n23507 = ~n44767 | ~n44851;
  assign n25189 = P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n25550 = n25243 | n25457;
  assign n24961 = ~n24944 & ~n24943;
  assign n24896 = ~n24895 & ~n24894;
  assign n25004 = ~n25609;
  assign n23233 = ~n23230 | ~n27550;
  assign n23230 = ~n27549;
  assign n28553 = ~n42208 | ~n42196;
  assign n23877 = ~n23878;
  assign n23910 = ~n23911 | ~n28172;
  assign n23911 = ~n28179;
  assign n23576 = n23004 & n28155;
  assign n28090 = ~n28094 | ~n28099;
  assign n23477 = ~n29817;
  assign n23719 = n23720 & n23854;
  assign n23854 = ~n23857 & ~n23855;
  assign n23720 = n22917 | n23721;
  assign n23855 = ~n32291;
  assign n23342 = ~n23588;
  assign n32527 = ~n28087 | ~n23387;
  assign n28012 = n27978 | n27977;
  assign n28295 = ~n28293 | ~P2_INSTADDRPOINTER_REG_3__SCAN_IN;
  assign n27693 = n27647 & n23396;
  assign n27672 = n27671 & n27670;
  assign n23686 = n40343 | n29855;
  assign n27336 = n27412 | n40428;
  assign n27221 = ~n27158 | ~P2_INSTQUEUE_REG_12__7__SCAN_IN;
  assign n34779 = ~n23065;
  assign n24009 = n38719 & P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n38740 = ~n34394 & ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n23759 = ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign n24633 = ~n24668 | ~n24617;
  assign n31508 = ~n43051;
  assign n25647 = ~n25595 & ~n25594;
  assign n25594 = ~n31528 & ~P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN;
  assign n25595 = ~n25593 & ~n25592;
  assign n25789 = ~n30138;
  assign n23808 = n23810 | n23809;
  assign n23809 = ~n30330;
  assign n25730 = n25728 | n42486;
  assign n42444 = ~n25883 ^ n25881;
  assign n25043 = n24999 | n24998;
  assign n23285 = n23628 & n23016;
  assign n26890 = n31459 & P1_STATE2_REG_0__SCAN_IN;
  assign n23843 = ~n23845 & ~n23844;
  assign n23845 = ~n23846;
  assign n23844 = ~n30172;
  assign n23839 = n23840 & n26112;
  assign n23841 = ~n30957;
  assign n23812 = ~n23816 & ~n23813;
  assign n29993 = n30013 & n30014;
  assign n23739 = n23741 & P1_INSTADDRPOINTER_REG_22__SCAN_IN;
  assign n23741 = n23931 | n23742;
  assign n30825 = ~n23558 | ~n23559;
  assign n23559 = ~n23561 & ~n23560;
  assign n23558 = n30898 & n30899;
  assign n23560 = ~n30908 | ~n23732;
  assign n23184 = ~n23731 & ~n23729;
  assign n23729 = ~n30883 | ~n23732;
  assign n30228 = n30292 | n23208;
  assign n23208 = n23210 | n23209;
  assign n23209 = ~n30226;
  assign n30269 = n30292 | n23211;
  assign n25498 = ~n23470;
  assign n31368 = ~n23802 & ~n23067;
  assign n23673 = ~n23702 | ~n23328;
  assign n23328 = n23329 & n23776;
  assign n23776 = ~n23528 | ~n22889;
  assign n25709 = ~n42393 & ~n23557;
  assign n43380 = ~n23620 | ~n31479;
  assign n23620 = ~n23619;
  assign n43082 = ~P1_STATE2_REG_2__SCAN_IN;
  assign n25392 = ~n25391;
  assign n44308 = ~P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n31524 = n23461 & n22995;
  assign n23461 = n31421 | n44850;
  assign n23460 = ~n31425 | ~n22969;
  assign n28879 = ~n32883;
  assign n23882 = ~n32951;
  assign n23517 = ~n23518 | ~n23828;
  assign n23828 = n23830 | n23829;
  assign n23518 = ~n23397 | ~n23014;
  assign n23832 = ~n39725 & ~n23833;
  assign n23833 = ~n39717;
  assign n29633 = ~n22922;
  assign n23880 = ~n23881 | ~n32089;
  assign n23881 = ~n29087;
  assign n32837 = ~n32862 | ~n32835;
  assign n33239 = n39140 & n39138;
  assign n23873 = ~n39587 & ~n23874;
  assign n23874 = ~n33072;
  assign n27632 = ~n27179 | ~n27607;
  assign n23884 = ~n31785 | ~n23885;
  assign n29780 = n28324 & n28323;
  assign n31832 = ~n23896 | ~n23247;
  assign n23944 = ~n32431;
  assign n23432 = n22917 & n23819;
  assign n23433 = n23434 & n23722;
  assign n23435 = ~n23860;
  assign n23753 = ~n22902 | ~P2_INSTADDRPOINTER_REG_23__SCAN_IN;
  assign n23898 = ~n23900 | ~n23899;
  assign n29025 = n39255 | n28071;
  assign n23700 = ~n29021;
  assign n23579 = ~n32832 & ~n23079;
  assign n39356 = n28158 & n28157;
  assign n23666 = n23667 & n32436;
  assign n32470 = ~n23162 | ~n28125;
  assign n28071 = ~n28077;
  assign n31958 = ~n31954 | ~n31955;
  assign n42140 = n42156 | n42112;
  assign n27775 = n23473 & n27752;
  assign n40436 = ~n42154 | ~n41686;
  assign n23708 = ~n23686 | ~n27672;
  assign n27566 = n27356 | n27543;
  assign n33228 = ~n27562 | ~n27561;
  assign n27561 = n27560 | n42209;
  assign n27562 = ~n27559 | ~n27558;
  assign n23367 = ~n37482 | ~n37502;
  assign n24704 = ~n24690 | ~n24689;
  assign n23547 = ~n23066 | ~n36180;
  assign n33801 = ~n33342 | ~P3_PHYADDRPOINTER_REG_1__SCAN_IN;
  assign n23796 = ~n36639 & ~n33287;
  assign n23797 = n33820 & P3_PHYADDRPOINTER_REG_7__SCAN_IN;
  assign n24585 = ~n23653 | ~n23652;
  assign n23653 = ~n23654 | ~P3_INSTADDRPOINTER_REG_7__SCAN_IN;
  assign n23196 = ~n24186 | ~n23534;
  assign n33307 = ~n33429 & ~n33399;
  assign n33408 = n24221 & n35753;
  assign n23202 = n36297 & n23766;
  assign n38673 = ~n38730;
  assign n24593 = ~n24482 & ~n24481;
  assign n24604 = ~n37494 & ~n24633;
  assign n31417 = ~n31512;
  assign n23848 = ~n29933;
  assign n30013 = ~n30058 & ~n30033;
  assign n30056 = n30182 | n23214;
  assign n23214 = ~n22981 | ~n23215;
  assign n23215 = ~n23216;
  assign n23810 = n31352 | n31338;
  assign n30332 = ~n31370 & ~n23808;
  assign n31370 = ~n31368 | ~n31367;
  assign n23632 = ~n30097;
  assign n23838 = ~n23836 | ~n25915;
  assign n23320 = ~n25839;
  assign n42963 = n25708 & n31248;
  assign n27060 = ~n30805 | ~n30804;
  assign n31541 = ~n31524;
  assign n43967 = n22905 | n44039;
  assign n44399 = ~P1_STATE2_REG_2__SCAN_IN & ~P1_STATE2_REG_3__SCAN_IN;
  assign n44152 = ~P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ^ P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n43471 = ~n43053 | ~n44851;
  assign n43199 = ~n43060 & ~n43061;
  assign n44418 = ~n44399;
  assign n31570 = n23147 & n22838;
  assign n31573 = ~n31580 | ~P1_STATE2_REG_2__SCAN_IN;
  assign n23458 = ~n23459 | ~P1_STATE2_REG_1__SCAN_IN;
  assign n23456 = n31565 & n22866;
  assign n39141 = n33240 & n39160;
  assign n33245 = ~n29800 & ~n29799;
  assign n29799 = ~n33217 & ~n33218;
  assign n31595 = ~n29864;
  assign n23252 = ~n31946;
  assign n32168 = n28971 & n28970;
  assign n28967 = ~n32823;
  assign n32405 = n28419 & n28418;
  assign n23902 = n32440 & n32420;
  assign n32457 = n28400 & n28399;
  assign n23886 = ~n32471;
  assign n23888 = ~n23889 & ~n23890;
  assign n23889 = ~n32492;
  assign n23887 = ~n32537;
  assign n23890 = ~n23891 | ~n32512;
  assign n23891 = ~n32536;
  assign n32564 = ~n23892 & ~n23895;
  assign n23892 = ~n23244 | ~n23893;
  assign n23264 = ~n23710 & ~n23829;
  assign n23413 = ~n23418 | ~n29335;
  assign n23418 = ~n39620;
  assign n23710 = ~n23830;
  assign n40111 = n39975 & n42213;
  assign n39975 = n39974 | n40200;
  assign n23665 = ~n32437;
  assign n23637 = n23853 & n23575;
  assign n23749 = ~n32712 & ~n23751;
  assign n23747 = ~n32712 & ~n23751;
  assign n23748 = ~n23280 | ~n23751;
  assign n32309 = n23859 & n28204;
  assign n29070 = ~n22932 | ~n22867;
  assign n32359 = ~n32346 | ~P2_INSTADDRPOINTER_REG_18__SCAN_IN;
  assign n23267 = ~n23222 | ~n33023;
  assign n23694 = n23269 & n28304;
  assign n40399 = ~n33115;
  assign n27883 = n27882;
  assign n41575 = ~P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n40557 = ~n40437 & ~n40436;
  assign n41002 = ~n41664 | ~n42196;
  assign n41664 = ~P2_STATE2_REG_2__SCAN_IN;
  assign n33788 = ~n38682;
  assign n24632 = ~n39110 & ~n35948;
  assign n35812 = ~n38681 | ~n39105;
  assign n33905 = ~n33906 & ~n33907;
  assign n34371 = ~n34478;
  assign n23366 = ~n35688;
  assign n24021 = n24315 & P3_INSTQUEUE_REG_15__0__SCAN_IN;
  assign n35504 = ~n23354 & ~n38799;
  assign n33428 = ~n36767 | ~n24646;
  assign n23760 = n23762 & n23761;
  assign n23761 = ~P3_INSTADDRPOINTER_REG_28__SCAN_IN;
  assign n33284 = n24252 | n24251;
  assign n23535 = ~n23536 | ~n24572;
  assign n37197 = n39056 | n38810;
  assign n39105 = ~n38799;
  assign n38815 = ~P3_STATE2_REG_1__SCAN_IN & ~n39118;
  assign n43062 = ~P1_ADDRESS_REG_29__SCAN_IN | ~n26952;
  assign n23182 = ~n23613 ^ P1_INSTADDRPOINTER_REG_30__SCAN_IN;
  assign n23613 = ~n30654 | ~n30653;
  assign n23611 = ~n23315 & ~n22915;
  assign n23315 = ~n31032;
  assign n31091 = ~n23607 & ~n31117;
  assign n23607 = n23608 | n25715;
  assign n23608 = n25714 | n22979;
  assign n39888 = n31969 & n39160;
  assign n31969 = ~n33140 | ~n31968;
  assign n40397 = ~n29013 | ~n28284;
  assign n23502 = ~n32305;
  assign n23503 = ~n29070 | ~n32752;
  assign n40408 = ~n33125;
  assign n39132 = ~n35945 | ~n33788;
  assign n35945 = ~n35812;
  assign n35667 = ~n36098 & ~n35677;
  assign n35671 = ~n37514 | ~n35504;
  assign n23659 = n33302 & n23660;
  assign n23660 = n33303 & n33376;
  assign n23200 = n33281 & n36629;
  assign n23452 = ~n25639 | ~n25613;
  assign n25615 = n25645 | n25618;
  assign n23311 = ~n25616;
  assign n27916 = ~P2_INSTQUEUE_REG_2__5__SCAN_IN;
  assign n23595 = ~n27903 | ~n27894;
  assign n27893 = n27892 | n28840;
  assign n23600 = n23601 & n27898;
  assign n27898 = n27897 | n28845;
  assign n27981 = ~P2_INSTQUEUE_REG_2__6__SCAN_IN;
  assign n27853 = n27886 | n27852;
  assign n26360 = n25065;
  assign n26320 = ~n26629;
  assign n24754 = ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n25619 = ~n26986 | ~P1_STATE2_REG_0__SCAN_IN;
  assign n24882 = ~P1_INSTQUEUE_REG_5__4__SCAN_IN;
  assign n29188 = ~n29756 | ~P2_INSTQUEUE_REG_3__0__SCAN_IN;
  assign n29171 = ~n29756 | ~P2_INSTQUEUE_REG_11__0__SCAN_IN;
  assign n27410 = n29577 | n27845;
  assign n27849 = n27905 | n29278;
  assign n27777 = n27776 & n40456;
  assign n27759 = n27892 | n28700;
  assign n29536 = ~P2_INSTQUEUE_REG_8__0__SCAN_IN;
  assign n23276 = n27569 & P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN;
  assign n27447 = n29306 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n24969 = ~P1_INSTQUEUE_REG_5__1__SCAN_IN;
  assign n26753 = n24972;
  assign n23508 = ~n22988 | ~n23509;
  assign n23509 = ~n25278;
  assign n23735 = ~n24906 | ~n23183;
  assign n25692 = ~n44842 | ~n23557;
  assign n23602 = ~n24754;
  assign n24878 = ~n24877 & ~n24876;
  assign n23098 = n23697 & n27624;
  assign n29696 = ~n29756 | ~P2_INSTQUEUE_REG_11__6__SCAN_IN;
  assign n29124 = n29753 & P2_INSTQUEUE_REG_9__4__SCAN_IN;
  assign n23681 = ~n31897;
  assign n29226 = ~P2_INSTQUEUE_REG_4__1__SCAN_IN;
  assign n29687 = ~P2_INSTQUEUE_REG_10__6__SCAN_IN;
  assign n29574 = ~P2_INSTQUEUE_REG_12__6__SCAN_IN;
  assign n29426 = ~P2_INSTQUEUE_REG_2__1__SCAN_IN;
  assign n23226 = ~n23227 | ~n27438;
  assign n27810 = ~P2_INSTQUEUE_REG_10__1__SCAN_IN;
  assign n23345 = ~n23565;
  assign n23721 = ~n23722;
  assign n23857 = ~n23043;
  assign n23565 = ~n23567 & ~n23566;
  assign n23566 = ~n32469;
  assign n23567 = ~n28122;
  assign n23573 = n22916 & n28081;
  assign n23905 = ~n23906;
  assign n23385 = ~n23386 | ~n23410;
  assign n23410 = ~n28086 | ~n23411;
  assign n23386 = ~n23180 | ~n22992;
  assign n23411 = ~n28075;
  assign n23406 = ~n29831 & ~n33073;
  assign n28033 = n28024 | n28023;
  assign n23236 = n28270 & n40456;
  assign n23396 = n27646 & P2_REIP_REG_1__SCAN_IN;
  assign n23369 = ~n27274 | ~n22836;
  assign n29576 = ~P2_INSTQUEUE_REG_8__6__SCAN_IN;
  assign n29669 = ~P2_INSTQUEUE_REG_8__5__SCAN_IN;
  assign n27125 = ~n27158 | ~P2_INSTQUEUE_REG_12__5__SCAN_IN;
  assign n27183 = ~n27158 | ~P2_INSTQUEUE_REG_12__3__SCAN_IN;
  assign n27446 = n27350 & n27349;
  assign n27350 = n27354 | n27347;
  assign n27359 = n41575 & n42134;
  assign n24608 = ~n24616 & ~n23368;
  assign n23368 = ~n23367;
  assign n34396 = ~n38695 | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n25592 = n25585 & n25584;
  assign n25593 = ~P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN & ~n43055;
  assign n24735 = ~P1_INSTQUEUE_REG_6__0__SCAN_IN;
  assign n24762 = ~n24758 & ~n24757;
  assign n26522 = ~n26568 | ~P1_PHYADDRPOINTER_REG_22__SCAN_IN;
  assign n25499 = n25133 | n25132;
  assign n23322 = ~n23971 | ~n25601;
  assign n25685 = n24833 | n24832;
  assign n23302 = n25503 & n25508;
  assign n23211 = ~n23212 | ~n23803;
  assign n23212 = ~n30291;
  assign n25464 = n25463 | n25542;
  assign n23329 = ~n25442 | ~n25441;
  assign n23626 = ~n22993;
  assign n25455 = n25378 | n25377;
  assign n25443 = n25345 | n25344;
  assign n25139 = ~n25061 | ~n25060;
  assign n23557 = n25011;
  assign n31446 = ~n31445;
  assign n25134 = ~n26986 & ~n44851;
  assign n43548 = n31479 | n23621;
  assign n29801 = ~n29803 & ~n29802;
  assign n23924 = ~n23925 | ~n28221;
  assign n23925 = ~n28216;
  assign n23915 = ~n28142;
  assign n28127 = n28552 & P2_EBX_REG_11__SCAN_IN;
  assign n28080 = ~n22865 & ~n23572;
  assign n28073 = n28064 & n28063;
  assign n28064 = n28609 | n28552;
  assign n28094 = ~n23373 | ~n28056;
  assign n23373 = ~n23374 | ~n29824;
  assign n29577 = ~n29753 | ~n29098;
  assign n27700 = n27647 & n23395;
  assign n23711 = n27606 & n27644;
  assign n29749 = ~P2_INSTQUEUE_REG_8__7__SCAN_IN;
  assign n29709 = ~n29756 | ~P2_INSTQUEUE_REG_3__6__SCAN_IN;
  assign n23263 = ~n29626;
  assign n23400 = ~n23517 | ~n23680;
  assign n29331 = n27656 | n42214;
  assign n29330 = ~n29312 | ~n29311;
  assign n29311 = n29310 & n29309;
  assign n28152 = ~n28145 | ~n23916;
  assign n28150 = ~n28145 | ~n28146;
  assign n23923 = n23924 | n23046;
  assign n28160 = n28552 & P2_EBX_REG_14__SCAN_IN;
  assign n23381 = ~n23380 | ~n23940;
  assign n23940 = ~n32455 & ~n23941;
  assign n23699 = n22985 & n28122;
  assign n23869 = ~n23873 & ~n23870;
  assign n23868 = ~n33045;
  assign n32602 = n28093 & n39605;
  assign n27795 = n27794 | n27793;
  assign n23919 = ~n27783 | ~n23920;
  assign n23378 = n27804 & n27803;
  assign n27501 = n27500 | n27499;
  assign n28577 = n39849 | n28555;
  assign n23571 = ~n23569;
  assign n23716 = n27601 & n39593;
  assign n23707 = ~n40519 | ~n23706;
  assign n23693 = n23206 & n27752;
  assign n23691 = ~n40343 & ~n27752;
  assign n27552 = n27364 | n27363;
  assign n23551 = ~n33811 & ~n23552;
  assign n23548 = ~n36347;
  assign n23534 = ~P3_INSTADDRPOINTER_REG_5__SCAN_IN;
  assign n23995 = ~n23986 & ~n23985;
  assign n35811 = ~n39112;
  assign n38724 = ~n24009;
  assign n23356 = ~n23358 & ~n23357;
  assign n23216 = ~n23217 | ~n30156;
  assign n23217 = ~n30181;
  assign n26184 = ~n26113 & ~n30891;
  assign n23625 = ~n23470 & ~n23469;
  assign n23469 = ~n23967;
  assign n23678 = ~n43057;
  assign n25022 = n24863 | n24862;
  assign n23849 = ~n29968 | ~n23850;
  assign n30440 = n25053;
  assign n26910 = n31459 & n25662;
  assign n26975 = n26899 & P1_PHYADDRPOINTER_REG_29__SCAN_IN;
  assign n26842 = ~n26794 | ~P1_PHYADDRPOINTER_REG_27__SCAN_IN;
  assign n26794 = n26745 & P1_PHYADDRPOINTER_REG_26__SCAN_IN;
  assign n26745 = P1_PHYADDRPOINTER_REG_25__SCAN_IN & n26702;
  assign n26656 = ~n26522 & ~n30743;
  assign n26399 = ~n26526 | ~P1_PHYADDRPOINTER_REG_20__SCAN_IN;
  assign n26318 = ~n26275 & ~n30174;
  assign n26267 = ~n26231 & ~n30855;
  assign n23628 = n23839 & n26151;
  assign n26072 = ~n26066 & ~n30307;
  assign n26031 = ~n25991 & ~n25990;
  assign n25990 = ~P1_PHYADDRPOINTER_REG_9__SCAN_IN;
  assign n23287 = n25412 & n25849;
  assign n23811 = ~n23813 & ~n29972;
  assign n30140 = ~n25790 | ~n25789;
  assign n23210 = n23211 | n30243;
  assign n30845 = ~n30878 | ~n25547;
  assign n23733 = n25551 & P1_INSTADDRPOINTER_REG_15__SCAN_IN;
  assign n23806 = ~n23808 & ~n23807;
  assign n23807 = ~n30314;
  assign n25507 = ~n23186;
  assign n30633 = n25679 & n25678;
  assign n25679 = ~n31503 & ~n23557;
  assign n23308 = ~n23309 & ~n22923;
  assign n23309 = ~n25649;
  assign n31415 = n25043 & n26986;
  assign n23802 = ~n23801 | ~n23800;
  assign n23800 = ~n42385 & ~n31401;
  assign n42462 = ~n25730 | ~n25729;
  assign n42464 = n42462 | n42461;
  assign n25398 = n25171 & n25170;
  assign n23835 = n23299 | n25062;
  assign n25234 = ~n25195 | ~n25194;
  assign n43081 = n25236 & n25191;
  assign n44051 = ~n43969;
  assign n25182 = ~n25393 | ~n25391;
  assign n44132 = ~P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign n44765 = ~P1_STATEBS16_REG_SCAN_IN;
  assign n44775 = n43066 & P1_STATEBS16_REG_SCAN_IN;
  assign n31555 = n31487 & n31486;
  assign n23459 = ~n31587;
  assign n42244 = ~P1_STATE_REG_1__SCAN_IN;
  assign n28246 = n23233 & n27551;
  assign n29803 = n28215 | n23922;
  assign n23922 = n23923 | n23045;
  assign n23875 = ~n23877 | ~n23876;
  assign n23876 = ~n31811;
  assign n23908 = ~n23910 & ~n23034;
  assign n23909 = ~n28174;
  assign n39291 = ~n39324 & ~n39317;
  assign n28714 = ~n32971;
  assign n28118 = ~n23383 | ~n23382;
  assign n23382 = ~n28115;
  assign n23383 = ~n28114;
  assign n31646 = ~P2_PHYADDRPOINTER_REG_9__SCAN_IN;
  assign n23830 = ~n29616 & ~n23831;
  assign n23831 = ~n23832;
  assign n28572 = n28551 & n28550;
  assign n39973 = n33136 | n39140;
  assign n31831 = n28473 & n28472;
  assign n31666 = ~n31634 & ~n31633;
  assign n31664 = ~n31638 & ~n31637;
  assign n23853 = ~n22939 & ~n23475;
  assign n23479 = ~n23474 | ~n23010;
  assign n23476 = ~n29810 & ~n23477;
  assign n29829 = n31705 | n28071;
  assign n32653 = ~P2_INSTADDRPOINTER_REG_28__SCAN_IN;
  assign n23878 = ~n23879 | ~n31844;
  assign n23879 = ~n23880;
  assign n31901 = n28467 & n28466;
  assign n29087 = n28988 & n28987;
  assign n23486 = n23487 & n32373;
  assign n32904 = ~n28836 | ~n28835;
  assign n23817 = ~n23381 | ~n32454;
  assign n23617 = ~n23267 | ~n32524;
  assign n32536 = n28373 & n28372;
  assign n23426 = n29831 | n23429;
  assign n32525 = ~n32573 | ~n28075;
  assign n23634 = ~n23635 & ~n22954;
  assign n23635 = ~n39605;
  assign n23933 = ~n28295;
  assign n29800 = ~n33221 & ~n28316;
  assign n33136 = ~n33228 | ~n40456;
  assign n28291 = n28288 & n23973;
  assign n28290 = ~n27843 | ~n28565;
  assign n23256 = ~n27746;
  assign n29314 = ~n23708 | ~n22942;
  assign n33162 = ~n23571 | ~n23570;
  assign n23570 = ~n33160;
  assign n33165 = ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign n27773 = n23194 & n23473;
  assign n41324 = ~P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign n41503 = n27761 & n23279;
  assign n27536 = n27341 & n27342;
  assign n41489 = n42156 | n42170;
  assign n27613 = ~n27241 | ~n27242;
  assign n24710 = ~n24720;
  assign n33322 = ~n33801 & ~n33348;
  assign n38694 = ~n23355 & ~n38688;
  assign n38687 = ~n35811 | ~n35810;
  assign n36107 = ~n36113 | ~P3_PHYADDRPOINTER_REG_27__SCAN_IN;
  assign n36113 = ~n36164 & ~n36166;
  assign n36164 = ~n33802 | ~n33803;
  assign n36196 = ~n36832 | ~P3_INSTADDRPOINTER_REG_24__SCAN_IN;
  assign n36231 = ~n23548 | ~n23549;
  assign n23549 = ~n22886 & ~n23550;
  assign n23550 = ~P3_PHYADDRPOINTER_REG_22__SCAN_IN;
  assign n36267 = ~n23548 | ~n23551;
  assign n23794 = n23797 & P3_PHYADDRPOINTER_REG_14__SCAN_IN;
  assign n36483 = ~P3_PHYADDRPOINTER_REG_13__SCAN_IN;
  assign n37091 = ~n24594 & ~n22899;
  assign n36540 = ~n23797 | ~n23795;
  assign n36536 = ~n36639 & ~n34309;
  assign n36590 = ~P3_PHYADDRPOINTER_REG_9__SCAN_IN;
  assign n36622 = ~P3_PHYADDRPOINTER_REG_8__SCAN_IN;
  assign n36766 = ~n36196 & ~n36781;
  assign n24283 = ~n36191 | ~n24641;
  assign n36278 = ~n36297 | ~n24274;
  assign n36321 = ~n36462 | ~n24595;
  assign n23647 = ~n22899 & ~n37066;
  assign n23773 = ~n23775 & ~n24258;
  assign n37239 = n36989 | n36988;
  assign n36704 = ~n24575 | ~n24576;
  assign n37338 = ~n38758 & ~n38757;
  assign n30058 = ~n25804 | ~n25803;
  assign n25804 = ~n30056;
  assign n23804 = ~n27082;
  assign n27102 = n25790 & n22888;
  assign n30174 = ~P1_PHYADDRPOINTER_REG_17__SCAN_IN;
  assign n26273 = n26272 & n26271;
  assign n23846 = ~n30196 & ~n30216;
  assign n42411 = ~n30327;
  assign n30327 = n26998 | n26995;
  assign n26973 = n26972 & n26971;
  assign n23814 = ~n23816 & ~n23815;
  assign n42421 = ~n42439 & ~n42438;
  assign n43190 = ~n31515;
  assign n26660 = ~n30011;
  assign n26661 = ~n30010;
  assign n42582 = ~n42326;
  assign n30602 = n30440 & n31515;
  assign n42621 = ~n42592;
  assign n42752 = ~n27058 | ~n27057;
  assign n42761 = ~n42891;
  assign n30645 = ~n29931 ^ n29910;
  assign n30767 = ~P1_PHYADDRPOINTER_REG_21__SCAN_IN;
  assign n30792 = ~P1_PHYADDRPOINTER_REG_19__SCAN_IN;
  assign n30855 = ~P1_PHYADDRPOINTER_REG_15__SCAN_IN;
  assign n30891 = ~P1_PHYADDRPOINTER_REG_13__SCAN_IN;
  assign n30283 = ~n23031 & ~n26034;
  assign n30971 = n25945 & n25944;
  assign n30982 = n25935 & n25934;
  assign n31023 = ~P1_PHYADDRPOINTER_REG_5__SCAN_IN;
  assign n42895 = n42907;
  assign n23824 = ~n25406 ^ n23822;
  assign n23822 = ~n25407;
  assign n42945 = ~n42937;
  assign n23323 = ~n23307 | ~n23742;
  assign n30652 = ~n30695 | ~n31049;
  assign n42947 = ~n42234 | ~n44851;
  assign n23931 = n30804 & n23957;
  assign n23624 = n23967 & n25601;
  assign n30980 = ~n25461 ^ P1_INSTADDRPOINTER_REG_7__SCAN_IN;
  assign n30992 = ~n23326 | ~n23673;
  assign n31400 = ~n23801 | ~n25741;
  assign n23928 = ~n23528 | ~n25446;
  assign n42929 = ~n42947;
  assign n44760 = n43632 | n44781;
  assign n31528 = ~P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN;
  assign n44744 = ~P1_STATE2_REG_1__SCAN_IN & ~P1_STATE2_REG_3__SCAN_IN;
  assign n43281 = n43221 & P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n43225 = n43072 | n43073;
  assign n43449 = P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & n43387;
  assign n43397 = n43072 | n43293;
  assign n44766 = ~P1_STATE2_REG_3__SCAN_IN;
  assign n43951 = n43879 & P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n44306 = ~P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN;
  assign n44138 = n44070 | n44069;
  assign n44294 = n44240 & P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n44230 = ~n44801;
  assign n44382 = n44417 & n44308;
  assign n44394 = n43058;
  assign n44468 = n43162;
  assign n44491 = n44417 & P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n44415 = n43471 | n43219;
  assign n44750 = ~n23147 | ~P1_STATE2_REG_3__SCAN_IN;
  assign n44853 = P1_STATE2_REG_2__SCAN_IN | P1_STATE2_REG_1__SCAN_IN;
  assign n44850 = ~n31582;
  assign n33223 = ~n33239;
  assign n23883 = ~n31723;
  assign n31699 = n29792 & n29791;
  assign n31736 = ~n32233 & ~n31754;
  assign n31789 = n28486 & n28485;
  assign n31806 = n29006 & n29005;
  assign n31813 = n31805;
  assign n31929 = n28447 & n28446;
  assign n23250 = n23253 & n23000;
  assign n29086 = n29033 | n29032;
  assign n23862 = ~n32168;
  assign n23865 = ~n32863;
  assign n39672 = ~n39677 & ~n42196;
  assign n32391 = n28426 & n28425;
  assign n23901 = ~n32405;
  assign n39709 = ~n23827 | ~n23832;
  assign n32585 = n28351 & n28350;
  assign n23150 = n27739 & n27732;
  assign n39814 = ~n39782;
  assign n27637 = n27665 & n27636;
  assign n33137 = ~n33228 & ~n33230;
  assign n23258 = ~n23257 & ~n29729;
  assign n23257 = ~n31859 & ~n23259;
  assign n23259 = ~n23035 | ~n23260;
  assign n31872 = ~n23515 ^ n23514;
  assign n23412 = ~n23058;
  assign n32153 = ~n32837 & ~n23861;
  assign n23861 = ~n22880 | ~n32151;
  assign n32171 = ~n39828;
  assign n31966 = n33229 | n33231;
  assign n23872 = ~n39588;
  assign n39586 = ~n39588 & ~n39587;
  assign n39660 = ~n28573 ^ n28572;
  assign n40435 = ~n40437;
  assign n32232 = ~n23248 ^ n29780;
  assign n23248 = ~n31788 & ~n23884;
  assign n23942 = n23943 & n32401;
  assign n23591 = ~n23372;
  assign n40329 = ~P2_PHYADDRPOINTER_REG_1__SCAN_IN;
  assign n40344 = n40337 | n29853;
  assign n23937 = ~n32653 & ~n23938;
  assign n23938 = ~P2_INSTADDRPOINTER_REG_27__SCAN_IN | ~P2_INSTADDRPOINTER_REG_29__SCAN_IN;
  assign n32615 = n29841 ^ n29842;
  assign n23468 = n23638 & n29810;
  assign n32279 = ~n23856 | ~n32291;
  assign n23856 = ~n23436 | ~n23433;
  assign n32727 = ~n23441 ^ n32293;
  assign n23618 = ~n23504 | ~n22902;
  assign n23270 = ~n29029 | ~n29075;
  assign n23939 = n29024 & n29023;
  assign n32344 = n39280 | n28185;
  assign n32782 = ~n32361 | ~n32362;
  assign n31947 = ~n23251 | ~n23253;
  assign n32817 = ~n23023 | ~n23578;
  assign n23238 = ~n40390 | ~n23239;
  assign n23273 = ~n28131 | ~n32468;
  assign n32917 = ~n32470 ^ n23047;
  assign n28087 = ~n28069 | ~n39544;
  assign n33213 = ~P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN;
  assign n40428 = ~P2_INSTQUEUE_REG_0__0__SCAN_IN;
  assign n40497 = ~P2_INSTQUEUE_REG_0__4__SCAN_IN;
  assign n40755 = n41490 & n42153;
  assign n40807 = ~n40740;
  assign n40746 = n40648 & P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN;
  assign n40920 = n40922 & P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n41144 = ~n41068;
  assign n42139 = n41490 & n40997;
  assign n41326 = n41255 & P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n41336 = n27773 & n33176;
  assign n41491 = ~n29313 | ~n27676;
  assign n29313 = ~n23708;
  assign n41680 = ~n41575 & ~n41591;
  assign n41591 = P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | n41768;
  assign n41703 = ~n40475 | ~n40474;
  assign n41710 = ~n40490 | ~n40489;
  assign n41733 = ~n40523 | ~n40522;
  assign n40531 = ~n40557;
  assign n41590 = ~n41490 & ~n41489;
  assign n41756 = ~n40559 | ~n40558;
  assign n41795 = ~n41693;
  assign n40518 = ~n41786 & ~n42196;
  assign n33217 = ~n27575 | ~n42180;
  assign n42214 = ~P2_STATE2_REG_0__SCAN_IN;
  assign n42111 = ~n33228 | ~P2_STATE2_REG_3__SCAN_IN;
  assign n27368 = n42123 & P2_STATE2_REG_0__SCAN_IN;
  assign n42197 = ~P2_STATE2_REG_0__SCAN_IN & ~P2_STATE2_REG_1__SCAN_IN;
  assign n38682 = ~n35810 & ~n27583;
  assign n33862 = n23792 & n23793;
  assign n23793 = ~n34376 & ~n23053;
  assign n23543 = n23545 | n34376;
  assign n23546 = ~n33956 & ~n23547;
  assign n23789 = ~n34376 & ~n23790;
  assign n23790 = n34376 & n23791;
  assign n33830 = n23554 & n23553;
  assign n23553 = ~n36272;
  assign n34024 = ~n33828 & ~n34376;
  assign n34585 = ~n24308;
  assign n35535 = n22830 & n23077;
  assign n23362 = ~n35994 & ~n23363;
  assign n37502 = ~n24418 & ~n24417;
  assign n35583 = ~n35596 & ~n35501;
  assign n35632 = ~n35597 & ~n35654;
  assign n35800 = ~n35745;
  assign n36833 = n36247 & n23768;
  assign n36249 = ~n36320 & ~n33412;
  assign n36247 = ~n36321 & ~n33412;
  assign n36880 = ~n36247;
  assign n36347 = ~n36384 | ~P3_PHYADDRPOINTER_REG_17__SCAN_IN;
  assign n36389 = ~n36666 & ~n33794;
  assign n36511 = ~P3_PHYADDRPOINTER_REG_12__SCAN_IN;
  assign n36508 = ~n36389;
  assign n37146 = ~n36554 | ~n23648;
  assign n37183 = ~n24594 & ~n37210;
  assign n37185 = ~n24592 | ~n24591;
  assign n36490 = n36727 & n37212;
  assign n23655 = n24584 & n23656;
  assign n23656 = ~n24587;
  assign n35948 = ~n37453;
  assign n36665 = ~n33285 | ~P3_PHYADDRPOINTER_REG_4__SCAN_IN;
  assign n36702 = ~n36730;
  assign n36730 = ~n36390 & ~n36389;
  assign n23769 = n23770 & n39046;
  assign n33294 = ~n33338 | ~P3_INSTADDRPOINTER_REG_30__SCAN_IN;
  assign n33388 = ~n24597 & ~n33393;
  assign n33429 = ~n36766 | ~n24646;
  assign n23762 = n24283 & n36764;
  assign n23763 = ~n23542 | ~n36497;
  assign n23204 = n36193 & n24282;
  assign n23764 = ~n23765 | ~n24278;
  assign n23765 = n24273 | n23767;
  assign n37363 = ~n38678;
  assign n38675 = ~n24720 | ~n24719;
  assign n38763 = ~n38745 | ~n38703;
  assign n38487 = ~P3_STATE2_REG_3__SCAN_IN;
  assign n39118 = ~P3_STATE2_REG_0__SCAN_IN;
  assign n44838 = ~n26969 | ~n26968;
  assign n23220 = n31037 | n42440;
  assign n23219 = ~n29941 & ~n29942;
  assign n42343 = ~n42373;
  assign n42500 = ~n30327 | ~n42469;
  assign n23954 = ~n31370 & ~n23810;
  assign n42559 = ~n42553;
  assign n42561 = n30348 & n44514;
  assign n30348 = n31424 | n30347;
  assign n30441 = ~n30645;
  assign n26922 = ~n26921 | ~n26920;
  assign n42622 = ~n30615;
  assign n42746 = n44835;
  assign n30729 = ~n23633 ^ n30032;
  assign n23633 = n30117 & n23064;
  assign n30053 = n30117 & n22898;
  assign n30753 = n30074 ^ n30099;
  assign n23837 = ~n42399;
  assign n42915 = ~n43061;
  assign n43061 = n44791 | n30631;
  assign n31032 = ~n23603 | ~n23316;
  assign n23316 = ~n25719 & ~n23317;
  assign n23317 = ~P1_INSTADDRPOINTER_REG_30__SCAN_IN;
  assign n23495 = ~n23440 | ~n23556;
  assign n23556 = ~n23583 | ~n23011;
  assign n31117 = ~n23318 | ~n25713;
  assign n23318 = n23319 & n42963;
  assign n31116 = ~n30673 ^ n23532;
  assign n23532 = ~n30742;
  assign n30775 = ~n23499 ^ P1_INSTADDRPOINTER_REG_21__SCAN_IN;
  assign n43054 = n43050 | n43049;
  assign n44757 = ~n31430 | ~n31429;
  assign n43207 = ~n43976 | ~n43092;
  assign n43312 = ~n43311 & ~n43310;
  assign n43544 = ~n44327 | ~n43480;
  assign n43713 = ~n43641 | ~n43640;
  assign n43876 = ~n43976 | ~n43812;
  assign n44047 = ~n43976 | ~n43975;
  assign n44215 = ~n44138;
  assign n44405 = ~n43098 | ~n43097;
  assign n44214 = ~n44327 | ~n44160;
  assign n44220 = ~n44145 | ~n44144;
  assign n44406 = ~n43064 | ~n43063;
  assign n44326 = ~n44325 & ~n44324;
  assign n44514 = ~n31573 & ~n44851;
  assign n23454 = ~n44517 | ~n22991;
  assign n40117 = ~n39141 | ~n39139;
  assign n31745 = ~n32232;
  assign n23249 = ~n23253 | ~n23252;
  assign n32169 = ~n23863 | ~n28967;
  assign n39653 = ~n42095 | ~n39647;
  assign n32406 = ~n32441 | ~n23902;
  assign n32421 = n32441 & n32440;
  assign n32472 = ~n23887 | ~n23888;
  assign n32493 = ~n32537 & ~n23890;
  assign n32550 = ~n32564 | ~n32563;
  assign n42170 = ~n42112;
  assign n39782 = n31948 & n39805;
  assign n32057 = ~n23513 ^ n31881;
  assign n31886 = ~n23827 | ~n23264;
  assign n39964 = n39888 & n31970;
  assign n39970 = ~n39888;
  assign n40022 = ~P2_STATE2_REG_0__SCAN_IN & ~n39976;
  assign n40077 = ~n40111;
  assign n40114 = ~n40076;
  assign n40273 = ~n40120 | ~n40456;
  assign n32369 = n23294 & n32782;
  assign n23294 = ~n22887 & ~n40323;
  assign n23281 = ~n32403 ^ P2_INSTADDRPOINTER_REG_16__SCAN_IN;
  assign n29905 = ~n29881 & ~n29880;
  assign n23188 = ~n32212 | ~n32638;
  assign n23146 = ~n22924 & ~n32645;
  assign n32230 = ~n28237 ^ P2_INSTADDRPOINTER_REG_27__SCAN_IN;
  assign n32781 = ~n23616 ^ n23615;
  assign n23615 = ~n32360;
  assign n32845 = n32404 & n23296;
  assign n23296 = n32403 & n40356;
  assign n32876 = ~n32433 ^ n23051;
  assign n32989 = ~n23170 ^ n32524;
  assign n33086 = ~n40397;
  assign n42133 = ~n42132;
  assign n40467 = ~P2_INSTQUEUE_REG_0__2__SCAN_IN;
  assign n40482 = ~P2_INSTQUEUE_REG_0__3__SCAN_IN;
  assign n40530 = ~P2_INSTQUEUE_REG_0__6__SCAN_IN;
  assign n40566 = ~n40434 | ~n40433;
  assign n40546 = ~n40427 & ~n40426;
  assign n40637 = n40580 | n42177;
  assign n40740 = n40755 & n41491;
  assign n40808 = ~n40739 & ~n40738;
  assign n40894 = ~n40820;
  assign n41063 = ~n40994 & ~n40993;
  assign n41832 = ~n41624;
  assign n41237 = ~n41176 | ~n41175;
  assign n41311 = ~n41245 & ~n41244;
  assign n41675 = ~n40439 | ~n40438;
  assign n41856 = n27656 | n40551;
  assign n41819 = ~n41710;
  assign n41838 = ~n41720;
  assign n41855 = ~n41740;
  assign n41867 = ~n41756;
  assign n41653 = ~n41590 | ~n41491;
  assign n41672 = ~n41773;
  assign n41690 = ~n40465 | ~n41686;
  assign n41700 = ~n40480 | ~n41686;
  assign n41745 = ~n40543 | ~n41686;
  assign n41796 = ~n41597;
  assign n41762 = ~n41687 | ~n41686;
  assign n41873 = ~n41792 | ~n23972;
  assign n41765 = ~n41675;
  assign n41868 = ~n40448;
  assign n42123 = ~P2_STATE2_REG_1__SCAN_IN;
  assign n33879 = ~n33905 & ~n34376;
  assign n33796 = ~n33795 & ~n38818;
  assign n35487 = n35391;
  assign n35623 = n35970 | n35634;
  assign n35677 = n35493 | n23070;
  assign n23365 = ~n23366 | ~n23069;
  assign n24218 = n24217 & n24216;
  assign n24180 = n24179 & n24178;
  assign n35784 = ~n38756 | ~n35504;
  assign n27595 = ~n24048 | ~n24047;
  assign n24047 = ~n24046 & ~n23948;
  assign n35752 = ~n35784;
  assign n36099 = ~n35966 | ~n35948;
  assign n35944 = n38804 | n35943;
  assign n33338 = ~n33428 & ~n33399;
  assign n37331 = ~n36726 ^ n23537;
  assign n36731 = ~n36691;
  assign n36152 = ~n23763 | ~n23762;
  assign n37383 = ~n37349 | ~n37197;
  assign n37382 = ~P3_INSTADDRPOINTER_REG_0__SCAN_IN;
  assign n39077 = ~n39032 | ~n39031;
  assign n39078 = ~n39077;
  assign n33585 = ~n33487;
  assign n23610 = ~n23798 | ~n31034;
  assign n23169 = n39228 & n23039;
  assign n32765 = ~n32750 | ~n40356;
  assign n23361 = ~n35514 & ~n22931;
  assign n33304 = n33297 & n23658;
  assign n23658 = n33298 & n23659;
  assign P3_U2833 = ~n23644 | ~n23173;
  assign n23173 = ~n33403 & ~n23033;
  assign U212 = ~n33460 | ~U214;
  assign n22865 = ~n28062 | ~n28061;
  assign n22866 = n23459 & P1_STATE2_REG_0__SCAN_IN;
  assign n22867 = n23190 & n22900;
  assign n32482 = ~n23190 | ~n23178;
  assign n34872 = ~n34525;
  assign n23504 = ~n22903;
  assign n22868 = n23504 & P2_INSTADDRPOINTER_REG_18__SCAN_IN;
  assign n29824 = ~n28552;
  assign n27389 = ~n33146;
  assign n22869 = n31788 | n23020;
  assign n43066 = ~n25858 ^ n25860;
  assign n27757 = ~n23473;
  assign n23914 = ~n28072;
  assign n24191 = ~n24297;
  assign n24297 = ~n24009 | ~n38725;
  assign n22870 = n23384 & n22983;
  assign n22871 = ~n28145 | ~n22927;
  assign n22872 = n23914 | n23913;
  assign n22873 = n23190 & n23082;
  assign n27119 = ~n27433;
  assign n22874 = ~n29618 ^ n29617;
  assign n31928 = ~n23251 | ~n23250;
  assign n22875 = ~n32441 | ~n22929;
  assign n30821 = ~n23271 | ~n25551;
  assign n23475 = ~n32198;
  assign n22876 = n29339 & n29340;
  assign n22877 = n25555 & n23166;
  assign n22878 = n28303 & P2_INSTADDRPOINTER_REG_7__SCAN_IN;
  assign n22879 = n25006 & n23726;
  assign n22880 = n28967 & n23862;
  assign n22881 = n23678 & n23041;
  assign n22882 = n23178 & n23076;
  assign n22883 = n23473 | n29855;
  assign n22884 = n23178 & n28313;
  assign n22885 = n22971 & n32527;
  assign n28149 = n28552 & P2_EBX_REG_17__SCAN_IN;
  assign n22886 = ~n23551 | ~P3_PHYADDRPOINTER_REG_21__SCAN_IN;
  assign n22887 = n23005 & n23190;
  assign n22888 = n22928 & n27104;
  assign n22889 = n25446 & n23927;
  assign n22890 = n23849 | n29949;
  assign n22891 = n27646 & P2_REIP_REG_0__SCAN_IN;
  assign n22892 = n34532 & P3_INSTQUEUE_REG_9__5__SCAN_IN;
  assign n22893 = ~n23748 | ~n23080;
  assign n22894 = n25565 & n22920;
  assign n22895 = n22876 & n23974;
  assign n22896 = n23691 & P2_INSTQUEUE_REG_3__1__SCAN_IN;
  assign n22897 = n23693 & P2_INSTQUEUE_REG_1__1__SCAN_IN;
  assign n40734 = ~n23692 | ~n23691;
  assign n34425 = ~n34320;
  assign n22898 = ~n30074 & ~n23632;
  assign n34394 = ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n23642 = ~n34394;
  assign n22899 = n23649 | n37085;
  assign n27569 = ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign n22900 = n23082 & P2_INSTADDRPOINTER_REG_21__SCAN_IN;
  assign n22901 = n22868 & P2_INSTADDRPOINTER_REG_19__SCAN_IN;
  assign n22902 = n22900 & P2_INSTADDRPOINTER_REG_22__SCAN_IN;
  assign n22903 = ~n28313 | ~n29054;
  assign n22904 = n23362 & P3_EAX_REG_26__SCAN_IN;
  assign n25838 = ~n25837 & ~n25836;
  assign n43569 = ~n43568 & ~n44230;
  assign n28366 = n28317;
  assign n25741 = ~n42385;
  assign n26192 = ~n30216;
  assign n22906 = n25390 & n25389;
  assign n40356 = ~n23239;
  assign n23239 = ~n29013 | ~n33220;
  assign n34564 = ~n34585;
  assign n30237 = ~n23841 | ~n23839;
  assign n28580 = ~n31974 & ~n28553;
  assign n30215 = ~n23841 | ~n23628;
  assign n22907 = n23397 & n22876;
  assign n22908 = ~n22830 | ~n23362;
  assign n22909 = ~n23221 & ~n30285;
  assign n22910 = ~n23166 | ~n30674;
  assign n22911 = n28215 | n28216;
  assign n22912 = ~n23777 & ~P1_STATE2_REG_0__SCAN_IN;
  assign n22913 = n23388 & n32574;
  assign n22914 = n28347 & P2_REIP_REG_3__SCAN_IN;
  assign n22915 = ~n31031 & ~P1_INSTADDRPOINTER_REG_30__SCAN_IN;
  assign n22916 = n23905 & n28132;
  assign n22917 = n28204 & n32306;
  assign n22918 = n24203 & n24202;
  assign n22919 = n32527 & n23385;
  assign n22920 = n23166 & n31035;
  assign n22921 = n28174 | n23910;
  assign n27622 = ~n28499;
  assign n22922 = n29302 | n23825;
  assign n22923 = n25660 | n43101;
  assign n22924 = n32633 & n40408;
  assign n22925 = n31928 | n31929;
  assign n22926 = ~n23544 & ~n34376;
  assign n22927 = n23916 & n23915;
  assign n22928 = n25789 & n23804;
  assign n22929 = n23902 & n23901;
  assign n22930 = n36610 | n37210;
  assign n22931 = n35789 | n36018;
  assign n22932 = n23178 & n23504;
  assign n22933 = n35514 | n35789;
  assign n22934 = n24663 | n24662;
  assign n22935 = n29836 | n29835;
  assign n22936 = n23884 | n29780;
  assign n22937 = n30632 | n42373;
  assign n22938 = n29086 | n23878;
  assign n29836 = ~n29828 ^ n29797;
  assign n23575 = ~n29836;
  assign n30152 = n26193 & n23843;
  assign n22939 = n32184 & n32617;
  assign n30171 = n26193 & n23846;
  assign n27103 = n25790 & n22928;
  assign n22940 = n23271 ^ n25454;
  assign n29864 = ~n29851 ^ n29850;
  assign n22941 = n28668 & n28714;
  assign n22942 = n29633 & P2_INSTQUEUE_REG_0__1__SCAN_IN;
  assign n28114 = ~n28080 | ~n28081;
  assign n22943 = n23745 & n28304;
  assign n28178 = ~n23909 | ~n28172;
  assign n22944 = n28835 & n28879;
  assign n28137 = ~n28080 | ~n23573;
  assign n22945 = n23863 & n22880;
  assign n22946 = n23717 & n23716;
  assign n22947 = n23756 | n24185;
  assign n22948 = n29860 & n29859;
  assign n22949 = n36652 & n24185;
  assign n22950 = n25615 & n25643;
  assign n22951 = n25641 & n25640;
  assign n30877 = ~n23730;
  assign n22952 = n30821 | n31078;
  assign n22953 = n23266 & n40348;
  assign n30994 = ~n22906 | ~n25449;
  assign n22954 = n40284 & P2_INSTADDRPOINTER_REG_3__SCAN_IN;
  assign n22955 = n25555 & n23956;
  assign n22956 = n27615 & n31598;
  assign n31033 = ~n29915 ^ n29914;
  assign n22957 = n32816 & n32815;
  assign n22958 = n23289 & n30662;
  assign n22959 = n27726 & n27725;
  assign n22960 = n25848 & n23951;
  assign n22961 = n24308 & P3_INSTQUEUE_REG_0__5__SCAN_IN;
  assign n22962 = n31142 & n31141;
  assign n22963 = P2_STATE2_REG_1__SCAN_IN | n33254;
  assign n28955 = ~n28553 & ~n28552;
  assign n22965 = n39223 & n39222;
  assign n22966 = n23268 & n23696;
  assign n22967 = n24762 & n23953;
  assign n22968 = P1_STATE2_REG_0__SCAN_IN | n44513;
  assign n32549 = n28365 & n28364;
  assign n22969 = n31423 & n31422;
  assign n22970 = n24737 & n24736;
  assign n22971 = n23385 & n23819;
  assign n22972 = n40479 & n40478;
  assign n22973 = n40494 & n40493;
  assign n22974 = n40527 & n40526;
  assign n22975 = n40542 & n40541;
  assign n22976 = n40564 & n40563;
  assign n22977 = n41892 & n41891;
  assign n22978 = n23342 & n23341;
  assign n23775 = ~n24257;
  assign n23218 = n30182 | n30181;
  assign n25790 = ~n23213;
  assign n23213 = n30182 | n23216;
  assign n22979 = n43031 & n30674;
  assign n22980 = n23285 & n26610;
  assign n23894 = ~n23895;
  assign n22981 = n22888 & n30083;
  assign n27570 = ~n29099;
  assign n22982 = n25232 | n23780;
  assign n27433 = ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN;
  assign n36290 = ~P3_PHYADDRPOINTER_REG_21__SCAN_IN;
  assign n22983 = n32390 & n32374;
  assign n22984 = n23830 & n23829;
  assign n22985 = n32454 & n32469;
  assign n22986 = n23132 & n32488;
  assign n22987 = n32634 | n40399;
  assign n22988 = ~n25312 | ~n25311;
  assign n22989 = ~n23546 & ~n23543;
  assign n22990 = n23680 & n22874;
  assign n23784 = ~n25570;
  assign n22991 = n23455 & n31579;
  assign n22992 = n28086 & n39559;
  assign n22993 = n25347 & n25346;
  assign n22994 = n23841 & n23285;
  assign n22995 = ~n23460 & ~n31424;
  assign n22996 = n23888 & n23886;
  assign n34309 = ~P3_PHYADDRPOINTER_REG_7__SCAN_IN;
  assign n22997 = n23482 | n23475;
  assign n22998 = n23121 & n23269;
  assign n22999 = n28073 & n28066;
  assign n23000 = n23252 & n31936;
  assign n23001 = n23626 & n25383;
  assign n23002 = n23912 & n22999;
  assign n23003 = n25464 & n25601;
  assign n23004 = n22927 & n28138;
  assign n23005 = n23178 & n22868;
  assign n23006 = n23178 & n22901;
  assign n23007 = n30898 & n30908;
  assign n23008 = n27348 & P2_INSTQUEUE_REG_9__6__SCAN_IN;
  assign n23009 = n27110 & n27109;
  assign n23010 = n23476 | n23475;
  assign n30010 = ~n23841 | ~n22980;
  assign n23011 = n23784 & n25566;
  assign n23012 = n22929 & n28427;
  assign n23013 = n22988 & n44851;
  assign n23014 = n22984 & n22895;
  assign n23015 = n33398 & n33397;
  assign n23016 = n23843 & n26317;
  assign n28044 = ~P2_INSTQUEUE_REG_12__7__SCAN_IN;
  assign n23017 = n32253 & n32252;
  assign n23018 = n23330 & n25448;
  assign n23019 = n23898 | n23897;
  assign n27644 = ~n42209;
  assign n23020 = n22936 | n23883;
  assign n23021 = n22890 | n23848;
  assign n23022 = ~n25568 & ~n22920;
  assign n23023 = n32832 | n23238;
  assign n23024 = n23665 & n32436;
  assign n23025 = n23789 | n36209;
  assign n23026 = n22941 & n23882;
  assign n23027 = n22944 & n23865;
  assign n28164 = n28552 & P2_EBX_REG_13__SCAN_IN;
  assign n23742 = ~n30821;
  assign n23166 = n30821;
  assign n29278 = ~P2_INSTQUEUE_REG_4__3__SCAN_IN;
  assign n29365 = ~P2_INSTQUEUE_REG_4__5__SCAN_IN;
  assign n29537 = ~P2_INSTQUEUE_REG_12__0__SCAN_IN;
  assign n29501 = ~P2_INSTQUEUE_REG_4__2__SCAN_IN;
  assign n23028 = n25570 | n25566;
  assign n29527 = ~P2_INSTQUEUE_REG_10__0__SCAN_IN;
  assign n23029 = n23421 & n33003;
  assign n28027 = ~P2_INSTQUEUE_REG_4__7__SCAN_IN;
  assign n35319 = n34532;
  assign n42949 = ~n42932;
  assign n23829 = ~n22874;
  assign n28089 = ~n28091 & ~n28090;
  assign n30849 = ~n23732;
  assign n29530 = n29355;
  assign n23030 = n26109 | n26108;
  assign n36554 = ~n36556 | ~n36497;
  assign n26391 = ~n43190 | ~P1_STATE2_REG_2__SCAN_IN;
  assign n23031 = ~n26030 | ~n26029;
  assign n40342 = n39163 | n42208;
  assign n32597 = ~n40342;
  assign n23917 = ~n28146;
  assign n23032 = n31370 | n31352;
  assign n23818 = ~n32454;
  assign n23033 = n33401 | n33400;
  assign n23034 = n28552 & P2_EBX_REG_22__SCAN_IN;
  assign n32511 = ~n32537 & ~n32536;
  assign n23035 = n29728 ^ n29727;
  assign n23036 = ~n28079 | ~n28078;
  assign n23037 = ~n33830 & ~n34376;
  assign n23038 = n23786 & n23789;
  assign n23039 = n39213 | n39495;
  assign n23040 = n28552 & P2_EBX_REG_10__SCAN_IN;
  assign n23041 = P1_STATE_REG_1__SCAN_IN ^ P1_STATE_REG_2__SCAN_IN;
  assign n23042 = n33137 | n23698;
  assign n23043 = n31814 | n28218;
  assign n23044 = n33143 | n23698;
  assign n23045 = n28552 & P2_EBX_REG_27__SCAN_IN;
  assign n23046 = n28552 & P2_EBX_REG_26__SCAN_IN;
  assign n23047 = n32469 & n32468;
  assign n23048 = n29303 & n29633;
  assign n32458 = ~n23887 | ~n22996;
  assign n23251 = ~n32458;
  assign n25549 = ~n25601;
  assign n44142 = n25242 & n25241;
  assign n23621 = ~n44142;
  assign n23049 = n29323 & n29322;
  assign n40323 = n39163 | n40456;
  assign n40348 = ~n40323;
  assign n23050 = n33880 | n33907;
  assign n23051 = n32432 & n32431;
  assign n23052 = n30292 | n30291;
  assign n30054 = ~n26398 & ~n26397;
  assign n23913 = ~n28073;
  assign n23053 = ~n34425 & ~n33880;
  assign n23054 = n32402 & n32401;
  assign n23055 = n32345 & n32344;
  assign n25988 = ~n25042 | ~P1_STATE2_REG_2__SCAN_IN;
  assign n23056 = n23397 & n39780;
  assign n23057 = n28295 & n28294;
  assign n23058 = n29629 & n29633;
  assign n23791 = ~n36234;
  assign n31677 = ~n27404 | ~n27536;
  assign n23059 = n23655 & n23657;
  assign n23060 = n29831 & n23429;
  assign n23061 = n22838 & n31416;
  assign n23062 = n28602 & n27878;
  assign n23063 = ~n30292 & ~n23210;
  assign n23064 = n22898 & n30054;
  assign n35405 = n34575;
  assign n34782 = ~n24318;
  assign n35328 = n34660;
  assign n34717 = ~n24297;
  assign n23066 = ~n36166 ^ n36111;
  assign n23393 = ~n43379;
  assign n23067 = n25747 ^ n27579;
  assign n33186 = ~n42134;
  assign n23648 = ~n23649;
  assign n23649 = ~n37087 | ~P3_INSTADDRPOINTER_REG_8__SCAN_IN;
  assign n23927 = ~P1_INSTADDRPOINTER_REG_5__SCAN_IN;
  assign n23068 = n28552 & n31682;
  assign n23069 = P3_EAX_REG_11__SCAN_IN & P3_EAX_REG_9__SCAN_IN;
  assign n37235 = ~P3_INSTADDRPOINTER_REG_7__SCAN_IN;
  assign n23279 = ~n33176;
  assign n29855 = ~n42214 | ~P2_STATE2_REG_2__SCAN_IN;
  assign n23278 = ~n29855;
  assign n23070 = n35498 | n23365;
  assign n23071 = P3_INSTADDRPOINTER_REG_7__SCAN_IN & P3_INSTADDRPOINTER_REG_6__SCAN_IN;
  assign n23766 = ~n23767;
  assign n23767 = ~n24274 | ~n23768;
  assign n23072 = ~n26911 & ~n23557;
  assign n23643 = ~n34396;
  assign n33023 = ~P2_INSTADDRPOINTER_REG_7__SCAN_IN;
  assign n23768 = ~n24596;
  assign n23581 = ~P1_INSTQUEUE_REG_9__6__SCAN_IN;
  assign n29869 = n28314 & P2_INSTADDRPOINTER_REG_24__SCAN_IN;
  assign n33073 = ~P2_INSTADDRPOINTER_REG_5__SCAN_IN;
  assign n23073 = ~n23937 | ~P2_INSTADDRPOINTER_REG_30__SCAN_IN;
  assign n44851 = ~P1_STATE2_REG_0__SCAN_IN;
  assign n23074 = ~n29773 | ~n29772;
  assign n29053 = ~n32851;
  assign n23075 = n23796 & n23797;
  assign n23640 = ~n23641;
  assign n23641 = ~n23753 & ~n22903;
  assign n23562 = ~n23563;
  assign n23563 = ~n23640 & ~n28533;
  assign n23076 = n28313 & P2_INSTADDRPOINTER_REG_15__SCAN_IN;
  assign n23077 = n22904 & P3_EAX_REG_27__SCAN_IN;
  assign n23078 = ~n23562 & ~n32222;
  assign n31580 = ~P1_STATE2_REG_1__SCAN_IN;
  assign n32362 = ~P2_INSTADDRPOINTER_REG_18__SCAN_IN;
  assign n23364 = ~P3_EAX_REG_26__SCAN_IN;
  assign n32222 = ~P2_INSTADDRPOINTER_REG_27__SCAN_IN;
  assign n23751 = ~P2_INSTADDRPOINTER_REG_25__SCAN_IN;
  assign n23079 = n32818 | n32831;
  assign n23080 = P2_INSTADDRPOINTER_REG_24__SCAN_IN | P2_INSTADDRPOINTER_REG_25__SCAN_IN;
  assign n23081 = ~n32653 & ~n32222;
  assign n32752 = ~P2_INSTADDRPOINTER_REG_22__SCAN_IN;
  assign n23082 = P2_INSTADDRPOINTER_REG_18__SCAN_IN & n28518;
  assign n33003 = ~P2_INSTADDRPOINTER_REG_6__SCAN_IN;
  assign n28542 = ~n22840 | ~n27610;
  assign n27761 = n23194 & n27757;
  assign n36652 = ~n24219 ^ P3_INSTADDRPOINTER_REG_6__SCAN_IN;
  assign n23198 = n36652 & n24184;
  assign n24220 = n24219 | n37257;
  assign n24219 = ~n24221 ^ n35753;
  assign n23083 = n42899;
  assign n42899 = ~n25440 | ~n25439;
  assign n29094 = ~n23276 | ~n27348;
  assign n23084 = n27155 & P2_INSTQUEUE_REG_2__6__SCAN_IN;
  assign n23085 = ~n28250 | ~n27609;
  assign n28258 = ~n28250 | ~n27609;
  assign n23303 = n23141 & n30828;
  assign n30828 = ~n30845 | ~n23184;
  assign n44843 = ~n31568;
  assign n25014 = n24961 & n24960;
  assign n23852 = ~n23480 | ~n23479;
  assign n23698 = n27624 & n31598;
  assign n23950 = n28283 & n27446;
  assign n23697 = n31598 & P2_STATE2_REG_0__SCAN_IN;
  assign n27758 = n23207 & n23086;
  assign n23086 = ~n23473 & ~n40343;
  assign n23087 = n27744 | n27745;
  assign n27722 = n27744 | n27745;
  assign n27863 = n27897 | n28763;
  assign n27749 = n27897 | n28678;
  assign n36706 = ~n24116 ^ P3_INSTADDRPOINTER_REG_3__SCAN_IN;
  assign n36750 = ~n27595 & ~P3_INSTADDRPOINTER_REG_0__SCAN_IN;
  assign n23088 = ~n27156 | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n23089 = ~n33146 & ~n27157;
  assign n39726 = ~n23414 | ~n23413;
  assign n23597 = ~n23090 | ~n23091;
  assign n23414 = n23416 & n22895;
  assign n23416 = ~n23417 | ~n29335;
  assign n27118 = n27116 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n23092 = n24806 & n24805;
  assign n36260 = ~n36347 & ~n22886;
  assign n24186 = ~n24184 | ~n24185;
  assign n26962 = ~n22838 | ~n23678;
  assign n42372 = n43057 & n43101;
  assign n42112 = n31959 & n31958;
  assign n23093 = n23178 & P2_INSTADDRPOINTER_REG_12__SCAN_IN;
  assign n25936 = ~n25498 | ~n23971;
  assign n30926 = ~n30928;
  assign n30928 = ~n25498 | ~n23624;
  assign n23744 = n43161 & n43101;
  assign n23094 = n26964 & n23674;
  assign n23596 = ~n27893 | ~n27899;
  assign n23360 = ~n24627;
  assign n32632 = ~n32200 ^ n23095;
  assign n23095 = n32199 & n32198;
  assign n41378 = n41375 & n23096;
  assign n23096 = ~n23097 & ~n41376;
  assign n23097 = n41400 & n41720;
  assign n23099 = n23697 & n27624;
  assign n23100 = ~n41002 & ~n41332;
  assign n27724 = n23697 & n27624;
  assign n23305 = ~n30663 ^ n23306;
  assign n38723 = ~n38725;
  assign n30995 = n23101 & n23102;
  assign n23102 = n25449 | n25389;
  assign n23103 = n25601 & P1_INSTADDRPOINTER_REG_6__SCAN_IN;
  assign n29103 = ~n27219;
  assign n27219 = ~n27433 & ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n24150 = n24134 & n24133;
  assign n23609 = ~n23611 & ~n23610;
  assign n23603 = ~n31059 & ~n25718;
  assign n31230 = ~n42960 & ~n43026;
  assign n23444 = ~n43051 | ~n23061;
  assign n42227 = ~n43051 | ~n44514;
  assign n31517 = n43051 & n30633;
  assign n23314 = ~n22950 & ~n25624;
  assign n24869 = ~n24947 | ~P1_INSTQUEUE_REG_9__4__SCAN_IN;
  assign n24986 = ~n24947 | ~P1_INSTQUEUE_REG_9__1__SCAN_IN;
  assign n43450 = ~n43397 & ~n44801;
  assign n23104 = ~n28955;
  assign n23105 = ~n23104;
  assign n23106 = ~n28088 | ~n23057;
  assign n28306 = n23189 & n22846;
  assign n30305 = ~n30257 ^ n30258;
  assign n28299 = n28298 & n28297;
  assign n23437 = ~n23301 | ~n23303;
  assign n23301 = ~n30946 | ~n23302;
  assign n41624 = n40501 & n40518;
  assign n23203 = ~n24253 | ~P3_INSTADDRPOINTER_REG_7__SCAN_IN;
  assign n27251 = n27249 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n27905 = ~n27768 | ~n23279;
  assign n27847 = n27904 | n27845;
  assign n27400 = ~n27399 & ~n23133;
  assign n27269 = ~n27380 | ~P2_INSTQUEUE_REG_0__4__SCAN_IN;
  assign n26869 = n24898;
  assign n23674 = ~n22838 | ~n31415;
  assign n24752 = n24905 | n24750;
  assign n39849 = n27632;
  assign n34610 = ~n24289;
  assign n30261 = n23221 | n23030;
  assign n23107 = ~n27881;
  assign n27881 = n27773 & n23279;
  assign n36333 = ~n24271 | ~n36497;
  assign n39729 = ~n39726 & ~n39725;
  assign n23402 = n39726 & n22874;
  assign n23709 = n23401 | n23261;
  assign n30946 = ~n30992 | ~n23392;
  assign n28543 = ~n27404;
  assign n42208 = n27404;
  assign n23441 = ~n23723 | ~n32307;
  assign n23108 = ~n40279 | ~P2_INSTADDRPOINTER_REG_4__SCAN_IN;
  assign n23109 = ~n27344 & ~n40501;
  assign n27603 = ~n27344 & ~n40501;
  assign n23110 = ~n23493 | ~n23112;
  assign n23114 = ~n23110 | ~n23111;
  assign n23111 = n31048 | n23742;
  assign n23112 = n25559 & n25563;
  assign n44391 = ~n44327 | ~n44326;
  assign n44499 = ~n44317 & ~n44801;
  assign n36213 = ~n23764 | ~n36333;
  assign n36215 = n36213 | P3_INSTADDRPOINTER_REG_24__SCAN_IN;
  assign n34777 = ~n35422;
  assign n24535 = ~n34777;
  assign n23405 = ~n23407 | ~n23406;
  assign n27768 = n23207 & n23483;
  assign n23171 = n32837;
  assign n23863 = ~n23171;
  assign n23113 = ~n23592 | ~n27604;
  assign n27606 = ~n23592 | ~n27604;
  assign n31074 = ~n31091 | ~P1_INSTADDRPOINTER_REG_26__SCAN_IN;
  assign n43013 = ~n25837 & ~n25706;
  assign n43031 = ~n25837 & ~n31535;
  assign n23310 = ~n25650 | ~n23308;
  assign n25650 = ~n25646 | ~n25645;
  assign n23605 = n25641 | n25638;
  assign n25637 = ~n25612 | ~n25645;
  assign n31727 = n31701;
  assign n31843 = ~n29086 & ~n23880;
  assign n32090 = ~n29086 & ~n29087;
  assign n27605 = n27643;
  assign n31964 = n27627;
  assign n23403 = ~n39726 | ~n22990;
  assign n27743 = n23140 & n23139;
  assign n23207 = ~n27743 | ~n27742;
  assign n23116 = ~n23903 | ~n23119;
  assign n23682 = ~n23116 | ~n23117;
  assign n23118 = ~n27621;
  assign n23119 = n27617 & n27621;
  assign n23243 = ~n27618 | ~P2_STATE2_REG_0__SCAN_IN;
  assign n23268 = ~n28305 | ~n33073;
  assign n31536 = ~n31474;
  assign n23120 = n23175 & n27880;
  assign n23121 = ~n32562 | ~P2_INSTADDRPOINTER_REG_6__SCAN_IN;
  assign n39106 = n35936;
  assign n23815 = ~n29936 | ~n29994;
  assign n23813 = ~n29994;
  assign n31961 = ~n39817 & ~n23279;
  assign n23131 = n23161 | n27764;
  assign n27279 = ~n29094;
  assign n27270 = ~n23122 & ~n23123;
  assign n23122 = ~n27266 | ~n27269;
  assign n23123 = ~n27267 | ~n27268;
  assign n27192 = ~n27185 & ~n23124;
  assign n23124 = ~n27184 | ~n27183;
  assign n23125 = ~n23129 | ~n23126;
  assign n23127 = n27772 | n27755;
  assign n23129 = ~n23131 & ~n23130;
  assign n23130 = n27756 | n23153;
  assign n23353 = ~n23132 | ~n23565;
  assign n23132 = ~n22919 | ~n32526;
  assign n23372 = ~n23132 | ~n23699;
  assign n23162 = ~n23132 | ~n28122;
  assign n23337 = ~n23340 | ~n23132;
  assign n27418 = ~n27158;
  assign n27135 = ~n27158 | ~P2_INSTQUEUE_REG_4__5__SCAN_IN;
  assign n27268 = ~n27158 | ~P2_INSTQUEUE_REG_4__4__SCAN_IN;
  assign n27374 = ~n27158 | ~P2_INSTQUEUE_REG_12__1__SCAN_IN;
  assign n27196 = ~n27158 | ~P2_INSTQUEUE_REG_4__3__SCAN_IN;
  assign n27335 = ~n27158 | ~P2_INSTQUEUE_REG_4__0__SCAN_IN;
  assign n27246 = ~n27158 | ~P2_INSTQUEUE_REG_12__4__SCAN_IN;
  assign n27314 = ~n27158 | ~P2_INSTQUEUE_REG_12__0__SCAN_IN;
  assign n27230 = ~n27158 | ~P2_INSTQUEUE_REG_4__7__SCAN_IN;
  assign n27289 = ~n27158 | ~P2_INSTQUEUE_REG_12__2__SCAN_IN;
  assign n27301 = ~n27158 | ~P2_INSTQUEUE_REG_4__2__SCAN_IN;
  assign n27158 = n27428 & P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n23526 = ~n23028 & ~n22894;
  assign n23133 = ~n27397 | ~n27398;
  assign n28493 = ~n28507 | ~n27657;
  assign n27171 = ~n23084 & ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n27689 = ~n27729 | ~n42120;
  assign n23160 = ~n23197 | ~n23134;
  assign n23134 = ~n22949 | ~n23199;
  assign n24179 = ~n23135 & ~n22961;
  assign n23135 = n22892 | n24171;
  assign n23136 = ~n23736 | ~n25859;
  assign n23137 = ~n27633 | ~n27634;
  assign n27661 = n23265 & n27278;
  assign n29694 = n27219;
  assign n25547 = ~n30879 & ~n25546;
  assign n27385 = ~n27384 & ~n27383;
  assign n28062 = ~n23138 | ~n29824;
  assign n23138 = ~n28060;
  assign n23820 = ~n28125;
  assign n27344 = ~n40486 | ~n27619;
  assign n23139 = ~n27737 | ~n27736;
  assign n23140 = ~n23149 | ~n23150;
  assign n23398 = ~n27647 | ~n22891;
  assign n42920 = ~n25422 | ~n25421;
  assign n23157 = ~n32210 & ~n32209;
  assign n23496 = ~n23304;
  assign n27176 = ~n27175 & ~n23142;
  assign n23142 = ~n27173 | ~n27174;
  assign n27145 = ~n27137 & ~n23143;
  assign n23143 = ~n27135 | ~n27136;
  assign n27668 = n27654 & n23293;
  assign n25397 = ~n25099 | ~n25098;
  assign n27756 = ~n27749 | ~n27750;
  assign n27720 = ~n27719 & ~n27718;
  assign n23145 = n29694;
  assign n27191 = ~n27190 & ~n23144;
  assign n23144 = ~n27188 | ~n27189;
  assign n27115 = ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN & ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN;
  assign n23265 = n27275 & n27276;
  assign n27265 = ~n27155 | ~P2_INSTQUEUE_REG_2__4__SCAN_IN;
  assign n27267 = n27265 & n29098;
  assign n23601 = ~n27895 & ~n23594;
  assign n23442 = ~n40577;
  assign n27890 = ~n40577 | ~P2_INSTQUEUE_REG_1__5__SCAN_IN;
  assign n27876 = n27875 & n27874;
  assign n23622 = ~n23437 | ~n22877;
  assign n32646 = ~n22987 | ~n23146;
  assign n28573 = ~n33112 | ~n33113;
  assign n23313 = ~n23312 | ~n23311;
  assign n25617 = ~n25610 | ~n23450;
  assign n31062 = ~n31078 & ~n31079;
  assign n25850 = n25412 & n23496;
  assign n23193 = ~n27668 | ~n27667;
  assign n23619 = n44767;
  assign n23718 = ~n23274 | ~n23275;
  assign n28015 = ~n23120 | ~n27947;
  assign n32223 = ~n28236 | ~n28235;
  assign n27889 = n27761 & n33176;
  assign n24832 = ~n23148 | ~n24831;
  assign n23148 = n24829 & n24830;
  assign n23639 = ~n23207 | ~n23473;
  assign n23149 = ~n28327;
  assign n27727 = ~n28317 | ~P2_INSTADDRPOINTER_REG_3__SCAN_IN;
  assign n28317 = ~n27666 | ~n27665;
  assign n32272 = ~n32257 | ~n32256;
  assign n27774 = n22827 & n27743;
  assign n32562 = ~n23151 | ~n23177;
  assign n23151 = n23165 & n28310;
  assign n27177 = ~n27169 & ~n23152;
  assign n23152 = ~n27167 | ~n27168;
  assign n27608 = ~n27599 | ~n22836;
  assign n27897 = ~n27758 | ~n27748;
  assign n23420 = ~n32226 ^ n32227;
  assign n27635 = ~n27627 & ~n27626;
  assign n23825 = ~n27656;
  assign n23153 = ~n27760 | ~n27759;
  assign n27685 = ~n27645 | ~n27644;
  assign n27345 = ~n23825 & ~n28542;
  assign n23473 = ~n23154 | ~n27717;
  assign n23154 = n27721 & n27716;
  assign n23298 = ~n23438 | ~n23078;
  assign n23291 = ~n40734;
  assign n23564 = ~n23163;
  assign n23163 = ~n27879 | ~n27878;
  assign n23387 = ~n23405 | ~n23029;
  assign n23599 = ~n23596 & ~n23595;
  assign n23978 = n28327 & n27738;
  assign n23408 = ~n32260 ^ n32259;
  assign n28507 = ~n28499 & ~n27655;
  assign n27206 = ~n27205 & ~n23155;
  assign n23155 = ~n27203 | ~n27204;
  assign n28328 = n27703 & n27702;
  assign n23688 = ~n23690;
  assign n27859 = ~n27858 & ~n23156;
  assign n23156 = ~n27853 | ~n27854;
  assign n27740 = n27739;
  assign n23274 = ~n22885 | ~n32526;
  assign P2_U2985 = ~n23157 | ~n32211;
  assign n27224 = ~n27222 & ~n27223;
  assign n23423 = ~n23158 | ~n32806;
  assign n23158 = ~n23159 | ~n40356;
  assign n23159 = ~n23292;
  assign n32703 = ~n23192 & ~n22893;
  assign n32271 = ~n23191 & ~n22893;
  assign n42432 = ~n42446 | ~n25884;
  assign n23755 = ~n23160 | ~n23196;
  assign n23668 = ~n23817;
  assign n23589 = ~n23590 | ~n23664;
  assign n23380 = ~n23820 | ~n32469;
  assign n23161 = ~n27780 | ~n27781;
  assign n28131 = ~n32470 | ~n32469;
  assign n32604 = n28088 | n23057;
  assign n28088 = ~n23175 ^ n23163;
  assign n23485 = ~n23431 | ~n23484;
  assign n28236 = ~n23485 | ~n29813;
  assign n27607 = ~n27178 | ~n23164;
  assign n23164 = ~n27176 | ~n27177;
  assign n27638 = ~n23683 | ~n27625;
  assign n23489 = ~n23584 | ~n23586;
  assign n23165 = ~n28308 | ~n28307;
  assign n23431 = ~n23718 | ~n23719;
  assign n23176 = ~n23298 | ~n32653;
  assign n31441 = ~n22839 | ~n23744;
  assign n23525 = ~n23527 | ~n25565;
  assign n28013 = ~n28014;
  assign P2_U3030 = ~n23351 | ~n23167;
  assign n23167 = n32828 & n32826;
  assign n27342 = ~n27325 | ~n27324;
  assign n23325 = ~n30948 | ~n25503;
  assign n31639 = ~n31662 | ~P2_PHYADDRPOINTER_REG_14__SCAN_IN;
  assign n31627 = ~n31668 | ~P2_PHYADDRPOINTER_REG_26__SCAN_IN;
  assign n31635 = ~n31664 | ~P2_PHYADDRPOINTER_REG_18__SCAN_IN;
  assign n31631 = ~n31666 | ~P2_PHYADDRPOINTER_REG_22__SCAN_IN;
  assign n39219 = ~n23168 | ~n39647;
  assign n23168 = ~n39216 ^ n39217;
  assign n29854 = ~n31670 | ~P2_PHYADDRPOINTER_REG_30__SCAN_IN;
  assign P2_U2833 = ~n22965 | ~n23169;
  assign n23170 = ~n28311 | ~n23267;
  assign n32221 = ~n23241 & ~n23240;
  assign n28301 = n32583 & n23189;
  assign n23389 = ~n23390 | ~n33003;
  assign n23593 = ~n23701 | ~n32362;
  assign n23590 = ~n23666;
  assign n23821 = ~n32348 ^ n23055;
  assign n23235 = ~n28595 | ~n31598;
  assign n23941 = ~n32468;
  assign n23391 = n23178 & n23563;
  assign n32687 = n32247 & n23471;
  assign n23679 = ~n23737 | ~n23742;
  assign n23440 = ~n23525 | ~n23526;
  assign n23527 = ~n30663;
  assign n24577 = ~n36704 | ~n36705;
  assign n23172 = ~n36677 | ~n36678;
  assign n24588 = ~n23657 | ~n24584;
  assign n28311 = ~n23694 | ~n23121;
  assign n23190 = ~n23443 | ~n23174;
  assign n23175 = ~n27844 | ~n28290;
  assign n28296 = ~n23564 | ~n23175;
  assign n23241 = ~n23176 | ~n40348;
  assign n23242 = ~n23176 | ~n32212;
  assign n23177 = ~n23687 | ~n28306;
  assign n32211 = ~n23179 | ~n40348;
  assign n32649 = ~n23179 | ~n40356;
  assign n32583 = ~n22964 | ~n23108;
  assign n32573 = ~n23180 | ~n39559;
  assign n30655 = ~n23182 | ~n42949;
  assign n23612 = ~n23182 | ~n43042;
  assign n23185 = ~n23186 | ~n25508;
  assign n23187 = ~n30826 & ~n30823;
  assign n28307 = ~n23189 | ~n23268;
  assign n23266 = ~n23190 | ~n23391;
  assign n32452 = n23190 & n23093;
  assign n32403 = ~n22882 | ~n23190;
  assign n23292 = ~n22884 | ~n23190;
  assign n29028 = ~n23006 | ~n23190;
  assign n32361 = ~n22932 | ~n23190;
  assign n23191 = ~n23746 | ~n40348;
  assign n23192 = ~n23746 | ~n40356;
  assign n27718 = ~n23193 | ~n23851;
  assign n27669 = ~n23851 ^ n23193;
  assign n23197 = ~n23198 | ~n22947;
  assign n23199 = ~n24184;
  assign n24183 = ~n24184 ^ n23756;
  assign n33305 = ~n23200 | ~n33280;
  assign n33381 = ~n23201 | ~n33280;
  assign n23201 = n33281 & n37201;
  assign n36612 = ~n23203 | ~n24256;
  assign n23205 = ~n24281 | ~n36193;
  assign n23542 = ~n24281 | ~n23204;
  assign n36800 = ~n23205 ^ P3_INSTADDRPOINTER_REG_26__SCAN_IN;
  assign n33144 = ~n23207;
  assign n23206 = ~n40343;
  assign n39618 = n33144 & n39639;
  assign n39810 = ~n39817 & ~n23207;
  assign n23521 = ~n23438 | ~n22901;
  assign n30180 = ~n23218;
  assign n29946 = ~n23220 | ~n23219;
  assign n31037 = ~n29952 ^ n29936;
  assign n23221 = ~n30284 & ~n30283;
  assign n28304 = ~n23428 | ~n22878;
  assign n32559 = ~n23222 ^ P2_INSTADDRPOINTER_REG_7__SCAN_IN;
  assign n30970 = n23223 & n23630;
  assign n23223 = n23629 & n23286;
  assign n23224 = ~n23838 | ~n25908;
  assign n23836 = ~n23225 | ~n25849;
  assign n23528 = ~n23225 | ~n25601;
  assign n23225 = ~n23627 ^ n22993;
  assign n27442 = ~n27441 & ~n23226;
  assign n23228 = ~n27509 | ~P2_INSTQUEUE_REG_11__3__SCAN_IN;
  assign n23229 = ~n27510 | ~P2_INSTQUEUE_REG_3__3__SCAN_IN;
  assign n27554 = ~n23233 | ~n23231;
  assign n27486 = ~n23235 | ~n27445;
  assign n27449 = ~n23234 | ~n23235;
  assign n23237 = ~n33228 | ~n23236;
  assign n28276 = ~n23237 | ~n28275;
  assign n29798 = ~n23266 & ~n23073;
  assign n23471 = n23266 & n40356;
  assign n23240 = ~n32212;
  assign n32665 = ~n23242 & ~n23239;
  assign n39579 = ~n23244 | ~n28336;
  assign n39582 = ~n23894 | ~n23244;
  assign n31900 = ~n23896;
  assign n23247 = ~n31901;
  assign n31935 = ~n32458 & ~n23249;
  assign n27748 = ~n27751;
  assign n29318 = ~n33176 | ~n23278;
  assign n33176 = ~n27751 ^ n23255;
  assign n23255 = ~n27718;
  assign n27751 = ~n23256 ^ n27747;
  assign n29682 = ~n31859 & ~n31860;
  assign n23260 = ~n31860;
  assign n23261 = ~n39726 & ~n23262;
  assign n31908 = ~n39726 & ~n23710;
  assign n27601 = ~n27600 | ~n23265;
  assign n28315 = ~n23266 | ~n32222;
  assign n23578 = ~n23159 | ~n23579;
  assign n30953 = ~n23271 | ~n23003;
  assign n23732 = ~n23271 | ~n23733;
  assign n30695 = ~n23679 | ~n23272;
  assign n23272 = ~n25562 | ~n23738;
  assign n23638 = n23860 & n23722;
  assign n27409 = n23276 & P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n23277 = ~n27570 | ~n22858;
  assign n27151 = ~n23008 | ~n22858;
  assign n27413 = ~n29094;
  assign n39667 = n33176 & n39639;
  assign n27882 = ~n27779 | ~n23279;
  assign n32799 = ~n23292 & ~n23079;
  assign n27428 = ~P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN & ~P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN;
  assign n23750 = ~n23280 | ~n32712;
  assign n32398 = n23281 & n40348;
  assign n25858 = ~n23736 | ~n23282;
  assign n23282 = ~n23284 | ~n23283;
  assign n23283 = ~n25138;
  assign n23284 = ~n25397;
  assign n30981 = ~n23629 | ~n23630;
  assign n23286 = ~n30982;
  assign n23288 = ~n23496 | ~n23287;
  assign P1_U2970 = ~n23290 | ~n22958;
  assign n23289 = ~n30657 | ~n42915;
  assign n23290 = ~n23305 | ~n42949;
  assign n27763 = ~n23692 | ~n22896;
  assign n27867 = ~n23291 | ~P2_INSTQUEUE_REG_3__3__SCAN_IN;
  assign n23683 = ~n23682 | ~n23293;
  assign n23293 = n23714 & n23715;
  assign n32356 = ~n23295 & ~n40323;
  assign n32778 = ~n23295 & ~n23239;
  assign n32415 = n32404 & n23297;
  assign n23297 = n32403 & n40348;
  assign n32231 = ~n23298 | ~n28315;
  assign n43210 = ~n25062 | ~n23299;
  assign n23394 = ~n23299;
  assign n32404 = ~n23292 | ~n32831;
  assign n32848 = ~n32419 | ~n23292;
  assign n25003 = ~n23675 | ~n23094;
  assign n25040 = ~n23300 | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN;
  assign n25033 = ~n23300 | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign n25242 = ~n23300 | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n25195 = ~n23300 | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n23300 = ~n25030 | ~n25034;
  assign n25435 = ~n23304 | ~n25424;
  assign n23704 = ~n25425 | ~n23304;
  assign n31045 = ~n23305 | ~n43042;
  assign n23306 = ~n30664;
  assign n23307 = ~n23114 | ~n23272;
  assign n23312 = ~n25617;
  assign n23449 = ~n23314 | ~n23313;
  assign n31380 = ~n42963;
  assign n23319 = ~n42961 | ~n23320;
  assign n25504 = ~n30950;
  assign n30824 = ~n23324 | ~n25508;
  assign n23324 = ~n23325 | ~n25507;
  assign n23327 = n30995 & n25448;
  assign n23330 = ~n23529 | ~n23928;
  assign n28308 = ~n23696 | ~n22846;
  assign n23332 = n43379 | P1_STATE2_REG_0__SCAN_IN;
  assign P2_U2988 = ~n32261 | ~n23333;
  assign n23333 = n23334 & n23017;
  assign n23334 = ~n32247 | ~n22953;
  assign n32332 = ~n23335 | ~n32597;
  assign n29093 = ~n23335 | ~n33086;
  assign n29063 = ~n23336 | ~n23939;
  assign n29026 = ~n23336 | ~n29023;
  assign n23336 = ~n23701 | ~n23700;
  assign n23584 = ~n23372 | ~n23588;
  assign n32346 = ~n23338 | ~n23337;
  assign n23339 = ~n22978 | ~n22870;
  assign n32418 = ~n32452 | ~P2_INSTADDRPOINTER_REG_13__SCAN_IN;
  assign n23344 = ~n23345 | ~n23819;
  assign n23419 = ~n23353 | ~n23819;
  assign n23347 = n28222 | n23348;
  assign n28223 = ~n23346 | ~n23347;
  assign n23346 = n29831 & n29825;
  assign n31768 = n29825 & n23347;
  assign n28226 = ~n28222;
  assign n23348 = ~n23046;
  assign n28166 = ~n23350 | ~n23573;
  assign n23351 = ~n23352 | ~n32820;
  assign n23352 = ~n32819 | ~n32818;
  assign n23436 = ~n23353 | ~n23432;
  assign n23354 = ~n38694 & ~n27589;
  assign n23355 = ~n27583;
  assign n35810 = ~n23359 | ~n38797;
  assign n38710 = ~n23359 | ~n23356;
  assign n23357 = ~n35943;
  assign n23358 = ~n23360 | ~n38797;
  assign n35519 = ~n23361 & ~n35517;
  assign n35558 = ~n22830 | ~n22904;
  assign n35574 = ~n22830 | ~P3_EAX_REG_24__SCAN_IN;
  assign n23363 = ~P3_EAX_REG_24__SCAN_IN;
  assign n24600 = ~n37494 & ~n23367;
  assign n24673 = ~n24625 | ~n23367;
  assign n38725 = P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN & P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign n27275 = ~n27626 | ~n23369;
  assign P2_U3029 = ~n23370 | ~n22957;
  assign n23370 = ~n23371 | ~n32810;
  assign n23371 = ~n32809 | ~n32808;
  assign n32438 = ~n23372 | ~n23817;
  assign n23375 = ~n28575 | ~n31598;
  assign n27808 = ~n23376 & ~n27807;
  assign n23376 = ~n23378 | ~n23377;
  assign n23377 = ~n27509 | ~P2_INSTQUEUE_REG_11__2__SCAN_IN;
  assign n23379 = ~n23667 | ~n23024;
  assign n23384 = ~n23588 | ~n23587;
  assign n23586 = n23384 & n32390;
  assign n32574 = ~n28110 | ~n28109;
  assign n23390 = ~n28087;
  assign n43716 = ~n23394 | ~n23393;
  assign n39772 = ~n23397 | ~n29339;
  assign n39926 = ~n23397 ^ n39780;
  assign n27653 = ~n23398 | ~n23977;
  assign n23399 = ~P2_REIP_REG_0__SCAN_IN;
  assign n23401 = ~n23400 | ~n23403;
  assign n31999 = ~n23404 | ~n39964;
  assign n31858 = ~n23404 | ~n39782;
  assign n23404 = ~n31854 ^ n23035;
  assign n32577 = ~n28087 ^ P2_INSTADDRPOINTER_REG_6__SCAN_IN;
  assign n32261 = ~n23408 | ~n32597;
  assign n32688 = ~n23408 | ~n33086;
  assign n29683 = ~n23409 & ~n29678;
  assign n32014 = ~n23409 ^ n31865;
  assign n23409 = ~n29679 ^ n23048;
  assign n23513 = ~n23709 ^ n23412;
  assign n23417 = ~n23705;
  assign n23415 = ~n39620 | ~n23705;
  assign n32481 = ~n23935 | ~n23745;
  assign n23745 = ~n28312 | ~P2_INSTADDRPOINTER_REG_8__SCAN_IN;
  assign n23859 = ~n23419 | ~n23860;
  assign n23467 = ~n23419 | ~n23468;
  assign n32228 = ~n23420 | ~n32597;
  assign n32666 = ~n23420 | ~n33086;
  assign n23421 = n39559 | n33073;
  assign n32575 = ~n32573 | ~P2_INSTADDRPOINTER_REG_5__SCAN_IN;
  assign n32809 = ~n23423 | ~n32807;
  assign n32819 = ~n23423 | ~P2_INSTADDRPOINTER_REG_15__SCAN_IN;
  assign n28312 = ~n23428;
  assign n23428 = ~n23500 | ~n29831;
  assign n23424 = ~n23500 | ~n23060;
  assign n23427 = ~n23501 | ~P2_INSTADDRPOINTER_REG_8__SCAN_IN;
  assign n23429 = ~P2_INSTADDRPOINTER_REG_8__SCAN_IN;
  assign n23430 = n39559 & n33073;
  assign n32257 = n23431 & n32277;
  assign n23434 = ~n23435 | ~n22917;
  assign n23723 = ~n23859 | ~n22917;
  assign n23494 = ~n30994;
  assign n23623 = ~n23437 | ~n22955;
  assign n30805 = ~n23437 | ~n25555;
  assign P1_U2968 = ~n23439 | ~n30644;
  assign n23439 = ~n23495 | ~n42949;
  assign n27754 = ~n23692 | ~n22897;
  assign n27861 = ~n40577 | ~P2_INSTQUEUE_REG_1__3__SCAN_IN;
  assign n27950 = ~n40577 | ~P2_INSTQUEUE_REG_1__6__SCAN_IN;
  assign n40568 = ~n23442 | ~n40636;
  assign n31419 = ~n23444 | ~n31418;
  assign n25634 = ~n23447 | ~n25631;
  assign n23447 = ~n23448 | ~n25626;
  assign n23448 = ~n23449 | ~n25625;
  assign n25608 = ~n25639;
  assign n23451 = ~n25611;
  assign P1_U3161 = ~n23453 | ~n44516;
  assign n23453 = ~n22968 | ~n23454;
  assign n44510 = ~n44517 | ~n31579;
  assign n23455 = ~n44806;
  assign n23457 = ~n31564 | ~n23456;
  assign n44512 = ~n23457 | ~n23458;
  assign n44515 = ~n31564 | ~n31565;
  assign n23568 = ~n23465 | ~n29840;
  assign n23463 = ~n23464 | ~n23465;
  assign n23464 = n29840 & n32597;
  assign n29931 = ~n23847;
  assign n23466 = ~n29910;
  assign n26964 = ~n25673 | ~n43101;
  assign n25673 = n24966 & n25021;
  assign n26193 = ~n30215;
  assign n40281 = ~n40280 | ~n23472;
  assign n23472 = ~n23934 | ~n28299;
  assign n23483 = ~n23473 & ~n23206;
  assign n27765 = ~n23473 & ~n27748;
  assign n27896 = n23614 & n23473;
  assign n40316 = ~n40344 & ~n23473;
  assign n23474 = n23719 | n22997;
  assign n23480 = ~n23481 | ~n23718;
  assign n32372 = ~n23489 | ~n29020;
  assign n23487 = ~n32374 | ~n23488;
  assign n23488 = ~n29020;
  assign n23490 = ~n23491 | ~n25432;
  assign n23492 = ~n42920 | ~n25423;
  assign n30673 = ~n22855;
  assign n23737 = ~n23493 | ~n25559;
  assign n25562 = ~n23505 | ~n25561;
  assign n23497 = n30992 & n30994;
  assign n23555 = ~n23495 | ~n43042;
  assign n31375 = ~n23497 ^ n23929;
  assign P1_U3010 = ~n23498 | ~n23009;
  assign n23498 = ~n30775 | ~n43042;
  assign n23499 = ~n27095 | ~n27094;
  assign n23500 = ~n23501;
  assign n28303 = ~n23501 | ~n28071;
  assign n28069 = ~n23695 | ~n23501;
  assign n23501 = ~n22849 | ~n28013;
  assign n25461 = ~n25460 | ~n25459;
  assign n23738 = ~n23506 | ~n25559;
  assign n23510 = ~n44767 | ~n23013;
  assign n23511 = ~n23513 | ~n23512;
  assign n23512 = ~n31881;
  assign n23514 = ~n29638;
  assign n23516 = ~n23709 | ~n23058;
  assign n23827 = ~n39726;
  assign n23519 = ~n29683 | ~n23035;
  assign n31854 = ~n29683 & ~n29682;
  assign n23524 = ~n32482 | ~n32771;
  assign n23523 = n22868 | P2_INSTADDRPOINTER_REG_19__SCAN_IN;
  assign n29731 = ~n27155;
  assign n27286 = ~n27155 | ~P2_INSTQUEUE_REG_10__2__SCAN_IN;
  assign n27249 = ~n27155 | ~P2_INSTQUEUE_REG_10__4__SCAN_IN;
  assign n27116 = ~n27155 | ~P2_INSTQUEUE_REG_10__5__SCAN_IN;
  assign n27317 = ~n27155 | ~P2_INSTQUEUE_REG_10__0__SCAN_IN;
  assign n27226 = ~n27155 | ~P2_INSTQUEUE_REG_2__7__SCAN_IN;
  assign n27216 = ~n27155 | ~P2_INSTQUEUE_REG_10__7__SCAN_IN;
  assign n27155 = n27115 & P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign n23529 = ~n23530 | ~n23927;
  assign n23530 = ~n42899 | ~P1_INSTADDRPOINTER_REG_4__SCAN_IN;
  assign n25440 = ~n23531 | ~n25601;
  assign n25907 = ~n23531 | ~n25849;
  assign n23531 = ~n25435 ^ n22988;
  assign n36651 = ~n23533 | ~n24186;
  assign n23533 = ~n24183 | ~P3_INSTADDRPOINTER_REG_5__SCAN_IN;
  assign n36726 = ~n23535;
  assign n24082 = ~n23537 | ~n23535;
  assign n23536 = ~n36749 | ~n36732;
  assign n24080 = ~n24552 ^ n24569;
  assign n36419 = ~n23538 | ~n24265;
  assign n36399 = ~n24268 | ~n23538;
  assign n23538 = ~n24264 | ~n36497;
  assign n24733 = ~n23539 | ~n24731;
  assign n23539 = ~n23540 | ~n22934;
  assign n23540 = ~n23541 | ~n33407;
  assign n23541 = ~n33306;
  assign n24284 = ~n23763 | ~n24283;
  assign n23544 = ~n33956 & ~n33832;
  assign n23545 = n34376 & n23066;
  assign n36312 = ~n36347 & ~n33811;
  assign n23552 = ~P3_PHYADDRPOINTER_REG_20__SCAN_IN;
  assign n33996 = ~n23554 ^ n23553;
  assign n23554 = n33829 | n34376;
  assign P1_U3000 = ~n23555 | ~n22960;
  assign n25013 = ~n25011;
  assign n23731 = ~n25548;
  assign n23561 = ~n25548 | ~n30883;
  assign n27879 = ~n27876 | ~n27877;
  assign n27660 = ~n27659 & ~n23707;
  assign n29907 = ~n23568 & ~n40397;
  assign n23572 = ~n23002 | ~n28089;
  assign n28072 = ~n22865 & ~n23574;
  assign n23574 = ~n28089;
  assign n29820 = ~n29801;
  assign n29827 = ~n23577 | ~n23068;
  assign n23577 = ~n29823;
  assign n29823 = ~n29801 | ~n29818;
  assign n32581 = ~n28309 | ~n23407;
  assign n23582 = ~n24804 | ~n23092;
  assign n23583 = ~n30663 | ~n23022;
  assign n32389 = ~n23585 | ~n23588;
  assign n23585 = ~n23591 | ~n23664;
  assign n23587 = ~n23664;
  assign n28248 = ~n23592;
  assign n23592 = ~n27602 | ~n27603;
  assign n28316 = ~n28248 | ~n28252;
  assign n33218 = ~n31598 | ~n28248;
  assign n23616 = ~n23593 | ~n32359;
  assign n32348 = ~n32347 | ~n23593;
  assign n27913 = ~n23598 & ~n23597;
  assign n23598 = ~n23599 | ~n23600;
  assign n24976 = n24753 & n23602;
  assign n31043 = ~n23603 & ~n31035;
  assign n23604 = ~n23605 | ~n25639;
  assign n23606 = ~n22951 & ~n25642;
  assign P1_U3001 = ~n23612 | ~n23609;
  assign n23614 = n27774 & n27748;
  assign n23936 = ~n23617;
  assign n43969 = ~n31479 | ~n23619;
  assign n26241 = ~n24947 | ~P1_INSTQUEUE_REG_12__1__SCAN_IN;
  assign n25559 = ~n23623 | ~n23742;
  assign n25997 = ~n23625 | ~n25849;
  assign n25382 = ~n23627 | ~n23626;
  assign n31000 = n23630 & n42432;
  assign n23629 = n30999 & n42432;
  assign n42399 = ~n42432 | ~n42431;
  assign n23631 = ~n42431;
  assign n30099 = ~n30117 | ~n30097;
  assign n30115 = ~n22994 | ~n30031;
  assign n30789 = ~n22994 ^ n30131;
  assign n28108 = ~n28093 | ~n23634;
  assign n29839 = ~n32200 | ~n23853;
  assign n23636 = ~n32200 | ~n23637;
  assign n36556 = ~n36612;
  assign n23644 = ~n23645 | ~n24731;
  assign n23645 = ~n23646 | ~n23015;
  assign n23646 = n33391 | n33399;
  assign n36463 = ~n36554 | ~n23647;
  assign n24579 = ~n23651 | ~n36690;
  assign n37293 = ~n23651 ^ n23650;
  assign n23650 = ~n36690;
  assign n23651 = ~n24577 | ~n24578;
  assign n23652 = ~n36662 | ~n23071;
  assign n23657 = ~n36662 | ~P3_INSTADDRPOINTER_REG_6__SCAN_IN;
  assign n23654 = ~n23655;
  assign n24574 = ~n23661 | ~n36750;
  assign n23661 = ~n36732;
  assign n29061 = ~n23662 | ~n33086;
  assign n32343 = ~n23662 | ~n32597;
  assign n23663 = ~n23591 | ~n32437;
  assign n23667 = ~n23668 | ~n32437;
  assign n23670 = ~n31478;
  assign n23671 = n23672 & n23778;
  assign n23672 = ~n31478 | ~n23781;
  assign n31478 = ~n25235 ^ n25234;
  assign n30993 = n23673 & n23018;
  assign n23677 = ~n31441;
  assign n23676 = ~n22881 | ~n22838;
  assign n25652 = ~n25001 | ~n31502;
  assign n31887 = ~n31896 | ~n31897;
  assign n23680 = ~n29626 & ~n23681;
  assign n29679 = ~n31870 | ~n29639;
  assign n31870 = ~n31872 | ~n31871;
  assign n23687 = ~n28309;
  assign n27716 = ~n23689 | ~n23688;
  assign n23689 = ~n27723;
  assign n27721 = ~n27720 | ~n23690;
  assign n28499 = ~n27631 | ~n27619;
  assign n33164 = n33145 | n23698;
  assign n23701 = ~n32346;
  assign n23703 = ~n25434 | ~n25433;
  assign n25885 = ~n23704 | ~n43065;
  assign n39621 = ~n39620 ^ n23705;
  assign n23705 = ~n23826 | ~n29327;
  assign n27598 = ~n23707;
  assign n27343 = n27598 & n39593;
  assign n23715 = ~n23711 | ~n27605;
  assign n23714 = ~n23717 | ~n23712;
  assign n23712 = n27601 & n23713;
  assign n27678 = ~n27605 | ~n23113;
  assign n23713 = n39593 & P2_STATE2_REG_0__SCAN_IN;
  assign n23717 = ~n27598 | ~n27661;
  assign n25046 = ~n23727 | ~n23728;
  assign n25016 = ~n23725 | ~n23724;
  assign n25664 = ~n25007 | ~n25006;
  assign n23726 = ~n25053 | ~n25832;
  assign n30846 = ~n25548 | ~n30883;
  assign n23730 = ~n23007 | ~n30899;
  assign n23734 = ~n24909 & ~n23735;
  assign n24764 = ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN & ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN;
  assign n24919 = ~n24973 | ~P1_INSTQUEUE_REG_8__5__SCAN_IN;
  assign n23736 = ~n25397 | ~n25138;
  assign n25558 = ~n23740 | ~n23166;
  assign n23740 = ~n30805 | ~n23931;
  assign n25233 = ~n23743;
  assign n25412 = ~n22852 | ~n23743;
  assign n23752 = ~n22837 | ~P2_INSTADDRPOINTER_REG_24__SCAN_IN;
  assign n23746 = ~n22837 | ~n23747;
  assign n32246 = ~n22837 | ~n23749;
  assign n32707 = n23750 & n23752;
  assign n36632 = ~n24253;
  assign n23754 = ~n24254;
  assign n24255 = ~n23755 | ~n24220;
  assign n36672 = ~n24183;
  assign n23756 = ~n24185;
  assign n24184 = ~n23757 | ~n24153;
  assign n23757 = ~n36681 | ~n36682;
  assign n33331 = n23763 & n23760;
  assign n23771 = ~n33275 | ~n36610;
  assign n33279 = ~n23771 | ~n23769;
  assign n23770 = ~n36610 | ~n24287;
  assign n36498 = ~n23774 | ~n24257;
  assign n23782 = ~n25229;
  assign n23783 = ~n25041 & ~n25043;
  assign n31476 = ~n31459 | ~n23783;
  assign n25062 = ~n23785 | ~n25139;
  assign n23785 = ~n25040 | ~n25039;
  assign n23786 = ~n33830 | ~n23791;
  assign n33831 = ~n23787 | ~n23025;
  assign n23787 = ~n33830 | ~n23788;
  assign n23788 = ~n36209 & ~n36234;
  assign n23792 = n33906 | n23050;
  assign n36408 = ~n23794 | ~n23796;
  assign n23795 = ~n36639;
  assign n31474 = ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN;
  assign n24759 = ~n31474;
  assign n23798 = ~n23799 | ~n25838;
  assign n23799 = ~n31033;
  assign n23801 = ~n42384;
  assign n31388 = ~n23802;
  assign n23803 = ~n30267;
  assign n23805 = ~n31370;
  assign n30292 = ~n23806 | ~n23805;
  assign n29952 = n29993 & n23812;
  assign n25823 = ~n29993 | ~n23814;
  assign n29975 = ~n29993 | ~n23811;
  assign n29973 = ~n29993 | ~n29994;
  assign n32358 = ~n23821 | ~n32597;
  assign n32780 = ~n23821 | ~n33086;
  assign n31461 = ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN & ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n42931 = ~n23824;
  assign n25406 = ~n42948 | ~P1_INSTADDRPOINTER_REG_0__SCAN_IN;
  assign n31009 = n23823 & n25408;
  assign n23823 = ~n23824 | ~P1_INSTADDRPOINTER_REG_1__SCAN_IN;
  assign n31981 = ~n39850 | ~n23825;
  assign n23826 = ~n39637 | ~n39636;
  assign n31488 = ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n44781 = ~n25850;
  assign n25422 = ~n25850 | ~n25601;
  assign n31534 = n23835 & n43880;
  assign n25099 = ~n23926 | ~n23835;
  assign n31022 = ~n23838;
  assign n31021 = ~n23837 | ~n25908;
  assign n30958 = ~n30957 & ~n30956;
  assign n23842 = ~n30956;
  assign n30195 = ~n26193 | ~n26192;
  assign n29967 = n29991 | n23849;
  assign n29932 = ~n29991 & ~n22890;
  assign n29969 = ~n29991 & ~n29992;
  assign n23850 = ~n29992;
  assign n23851 = ~n27638 | ~n27637;
  assign n27299 = ~n27295 | ~n23858;
  assign n23858 = ~n27409 | ~P2_INSTQUEUE_REG_5__2__SCAN_IN;
  assign n32862 = n32935 & n23027;
  assign n32885 = ~n28836 | ~n22944;
  assign n33046 = ~n23866 | ~n28617;
  assign n23866 = ~n23872 | ~n23873;
  assign n28623 = ~n23871 | ~n23867;
  assign n23870 = ~n28617;
  assign n23871 = ~n39588 | ~n28617;
  assign n32973 = ~n28669 | ~n22941;
  assign n32970 = ~n28669 | ~n28668;
  assign n31722 = ~n31788 & ~n22936;
  assign n31784 = ~n31788 & ~n31789;
  assign n23885 = ~n31789;
  assign n23893 = ~n32585;
  assign n23895 = ~n28344 | ~n28336;
  assign n29071 = ~n31928 & ~n23898;
  assign n23899 = ~n31929;
  assign n23900 = ~n29031;
  assign n27639 = ~n27616 | ~n27615;
  assign n27618 = ~n23903 | ~n27617;
  assign n28208 = ~n23909 | ~n23908;
  assign n28076 = ~n28072 | ~n22999;
  assign n27796 = n27787 | n23919;
  assign n31728 = ~n29820 | ~n29804;
  assign n29811 = ~n23921 | ~n29820;
  assign n23921 = n29804 & n29831;
  assign n28222 = ~n28215 & ~n23924;
  assign n28232 = ~n28215 & ~n23923;
  assign n31019 = ~n23928 ^ P1_INSTADDRPOINTER_REG_5__SCAN_IN;
  assign n23929 = ~n30980;
  assign n30754 = n25559 & n25558;
  assign n25027 = ~n25025 | ~n23930;
  assign n25052 = n25025 & n25024;
  assign n23934 = ~n23106 | ~n28295;
  assign n40279 = ~n23932 | ~n23106;
  assign n23935 = ~n28311 | ~n23936;
  assign n27132 = ~n27155 | ~P2_INSTQUEUE_REG_2__5__SCAN_IN;
  assign n27180 = ~n27155 | ~P2_INSTQUEUE_REG_10__3__SCAN_IN;
  assign n27377 = ~n27155 | ~P2_INSTQUEUE_REG_10__1__SCAN_IN;
  assign n27332 = ~n27155 | ~P2_INSTQUEUE_REG_2__0__SCAN_IN;
  assign n23946 = ~n32433 | ~n32431;
  assign n23943 = ~n23945 | ~n23944;
  assign n25722 = n31415 | n25405;
  assign n31509 = ~n26910 | ~n31415;
  assign n42216 = ~n27531 | ~n28543;
  assign n33112 = ~n28559 | ~n28558;
  assign n30644 = ~n30643 & ~n30642;
  assign n30632 = ~n26908 ^ n26907;
  assign n26923 = n30632 | n31515;
  assign n25183 = ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign n27134 = n27132 & n29098;
  assign n27242 = ~n27225 | ~n27224;
  assign n41808 = n40471 | n40551;
  assign n27904 = ~n27768 | ~n33176;
  assign n27241 = ~n27240 | ~n27239;
  assign n24917 = n22832 | n26748;
  assign n24886 = n22833 | n24885;
  assign n24830 = n26806 | n24822;
  assign n24776 = n22833 | n24775;
  assign n23947 = n26958 & n26957;
  assign n26894 = ~n25877;
  assign n23948 = n24045 | n24044;
  assign n23949 = n40443 & n40442;
  assign n23951 = n25847 & n23955;
  assign n42855 = ~n42761 | ~n43101;
  assign n23952 = n42599 | P1_EAX_REG_31__SCAN_IN;
  assign n23953 = n24761 & n24760;
  assign n23955 = ~n25846 & ~n25845;
  assign n23956 = n25557 & n25556;
  assign n23957 = n31134 & P1_INSTADDRPOINTER_REG_21__SCAN_IN;
  assign n23958 = n25065 | n24969;
  assign n23959 = n25065 | n24739;
  assign n23960 = n29902 | n29901;
  assign n38768 = ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN;
  assign n23961 = n24767 & n24766;
  assign n33722 = n33700;
  assign n23962 = n27429 | n27119;
  assign n23963 = n28811 & n28810;
  assign n40515 = ~BUF2_REG_29__SCAN_IN;
  assign n23964 = ~n28616 | ~n29824;
  assign n42755 = ~n42752 & ~n42746;
  assign n23965 = n40464 & n40463;
  assign n23966 = ~n26049 | ~n26048;
  assign n23967 = n25543 | n25542;
  assign n28476 = ~n28347;
  assign n23968 = n24732 & n33319;
  assign n24287 = ~P3_INSTADDRPOINTER_REG_30__SCAN_IN;
  assign n23969 = n28733 & n28732;
  assign n23970 = n28646 & n28645;
  assign n39945 = ~n39888 | ~n40552;
  assign n31948 = n23042 & n39160;
  assign n25147 = ~n25065;
  assign n23971 = n25497 | n25496;
  assign n23972 = n41791 | n41790;
  assign n23973 = n42096 | n40322;
  assign n23974 = n29342 & n39736;
  assign n23975 = n25869 & P1_STATE2_REG_2__SCAN_IN;
  assign n23976 = n27004 & n27003;
  assign n39520 = ~n42200 & ~n31599;
  assign n40390 = ~n32996;
  assign n32996 = n29013 & n28527;
  assign n33062 = n29013 & n23044;
  assign n23977 = ~n27642 | ~n27641;
  assign n24731 = ~n37349;
  assign n26818 = ~n26349;
  assign n23979 = n24968 & n24967;
  assign n27611 = n28258 & n40486;
  assign n25006 = ~n25015;
  assign n27494 = ~P2_INSTQUEUE_REG_2__0__SCAN_IN;
  assign n26622 = ~n24803;
  assign n24739 = ~P1_INSTQUEUE_REG_5__0__SCAN_IN;
  assign n26759 = ~n26326;
  assign n25199 = ~P1_INSTQUEUE_REG_6__2__SCAN_IN;
  assign n24885 = ~P1_INSTQUEUE_REG_6__4__SCAN_IN;
  assign n27347 = n41324 & P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n24681 = ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n25580 = n25573 & n25572;
  assign n26748 = ~P1_INSTQUEUE_REG_6__5__SCAN_IN;
  assign n25668 = n25015 | n25832;
  assign n24892 = n24891 & n24890;
  assign n27426 = n27425 | n27424;
  assign n27599 = ~n27612;
  assign n27396 = n27394 & n29098;
  assign n25577 = n25584 & n25576;
  assign n25066 = ~P1_INSTQUEUE_REG_6__1__SCAN_IN;
  assign n25399 = n25097 & n25096;
  assign n25023 = n25022 & n25832;
  assign n29283 = ~P2_INSTQUEUE_REG_8__3__SCAN_IN;
  assign n28670 = ~P2_INSTQUEUE_REG_8__1__SCAN_IN;
  assign n29717 = ~P2_INSTQUEUE_REG_4__6__SCAN_IN;
  assign n27836 = ~P2_INSTQUEUE_REG_12__1__SCAN_IN;
  assign n29540 = ~P2_INSTQUEUE_REG_4__0__SCAN_IN;
  assign n28045 = n29581 | n28044;
  assign n27202 = n27199 & n29098;
  assign n27182 = n27180 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n25587 = n44308 & P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN;
  assign n25584 = ~n44306 | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n25103 = ~P1_INSTQUEUE_REG_6__7__SCAN_IN;
  assign n25278 = n25277 & n25276;
  assign n27483 = n33213 & P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN;
  assign n29670 = ~P2_INSTQUEUE_REG_12__5__SCAN_IN;
  assign n29767 = n29100 & n29099;
  assign n29098 = ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n29394 = ~P2_INSTQUEUE_REG_12__3__SCAN_IN;
  assign n27321 = n27412 | n29536;
  assign n28032 = n28031 | n28030;
  assign n27547 = n27546 & P2_STATE2_REG_0__SCAN_IN;
  assign n34545 = ~n34777;
  assign n42328 = ~P1_PHYADDRPOINTER_REG_7__SCAN_IN;
  assign n24748 = ~n24747 & ~n24746;
  assign n44845 = ~n44841;
  assign n26912 = n25685;
  assign n31459 = ~n25660;
  assign n25194 = n25193 & n25192;
  assign n43799 = ~P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN;
  assign n27363 = ~n27483;
  assign n28240 = n27360 & n27522;
  assign n29713 = ~n29767;
  assign n29656 = ~P2_INSTQUEUE_REG_10__5__SCAN_IN;
  assign n28668 = ~n33006;
  assign n31634 = ~P2_PHYADDRPOINTER_REG_21__SCAN_IN;
  assign n28518 = P2_INSTADDRPOINTER_REG_20__SCAN_IN & P2_INSTADDRPOINTER_REG_19__SCAN_IN;
  assign n33145 = n28494;
  assign n27643 = ~n27345 | ~n23109;
  assign n26272 = n26391 | n26266;
  assign n25980 = ~n25938 & ~n42328;
  assign n26151 = ~n30238;
  assign n25946 = ~n30971;
  assign n26904 = n43082 & P1_STATEBS16_REG_SCAN_IN;
  assign n26702 = n26656 & P1_PHYADDRPOINTER_REG_24__SCAN_IN;
  assign n25877 = ~P1_STATE2_REG_2__SCAN_IN & ~P1_STATEBS16_REG_SCAN_IN;
  assign n26275 = ~n26267 | ~P1_PHYADDRPOINTER_REG_16__SCAN_IN;
  assign n25908 = ~n42400;
  assign n25436 = n25310 | n25309;
  assign n25241 = n25240 & n25239;
  assign n43880 = n43210;
  assign n31439 = n25652;
  assign n33237 = n31964 | n41895;
  assign n28179 = n28552 & P2_EBX_REG_21__SCAN_IN;
  assign n31607 = ~n40325 & ~n31606;
  assign n29636 = n29631 & n29301;
  assign n32883 = n28878 & n28877;
  assign n33141 = n28268 | n28267;
  assign n29306 = ~P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN;
  assign n38688 = ~n38681 | ~n39114;
  assign n36109 = ~P3_PHYADDRPOINTER_REG_28__SCAN_IN;
  assign n24595 = P3_INSTADDRPOINTER_REG_14__SCAN_IN & P3_INSTADDRPOINTER_REG_15__SCAN_IN;
  assign n24594 = ~n36554;
  assign n36760 = n33416 | n36808;
  assign n37147 = ~n37184;
  assign n25596 = n25591 | n25613;
  assign n25678 = ~n25002;
  assign n26439 = ~n26318 | ~P1_PHYADDRPOINTER_REG_18__SCAN_IN;
  assign n26972 = ~n44838;
  assign n26900 = ~n26894;
  assign n25803 = ~n30055;
  assign n31424 = ~n43051 & ~n31509;
  assign n30666 = ~P1_PHYADDRPOINTER_REG_28__SCAN_IN;
  assign n30743 = ~P1_PHYADDRPOINTER_REG_23__SCAN_IN;
  assign n30216 = n26191 & n26190;
  assign n30307 = ~P1_PHYADDRPOINTER_REG_11__SCAN_IN;
  assign n25902 = ~P1_PHYADDRPOINTER_REG_3__SCAN_IN;
  assign n25551 = ~n25550 & ~n25549;
  assign n25449 = ~P1_INSTADDRPOINTER_REG_6__SCAN_IN;
  assign n31535 = ~n25052 | ~n25709;
  assign n43717 = ~n43548;
  assign n44311 = ~n31534;
  assign n44792 = ~n43066;
  assign n43191 = ~n43056 | ~P1_STATE2_REG_3__SCAN_IN;
  assign n27560 = n27366 & n27551;
  assign n31632 = ~P2_PHYADDRPOINTER_REG_23__SCAN_IN;
  assign n29032 = n28984 & n28983;
  assign n31638 = ~P2_PHYADDRPOINTER_REG_17__SCAN_IN;
  assign n31642 = ~P2_PHYADDRPOINTER_REG_13__SCAN_IN;
  assign n39516 = ~n42200 | ~n31607;
  assign n28427 = ~n32391;
  assign n31811 = n29001 & n29000;
  assign n32950 = n32932;
  assign n29335 = n29334 & n29333;
  assign n33140 = n31967 & n31966;
  assign n32291 = n31833 | n28214;
  assign n32436 = n39402 | n28192;
  assign n41789 = ~P2_STATEBS16_REG_SCAN_IN;
  assign n41769 = ~P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN;
  assign n40922 = n40991 & n41769;
  assign n40991 = n29306 & P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign n41255 = n41154 & P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN;
  assign n27619 = ~n27310 | ~n27309;
  assign n40547 = ~n40556;
  assign n24720 = ~n24704 & ~n24703;
  assign n36538 = ~P3_PHYADDRPOINTER_REG_11__SCAN_IN;
  assign n33848 = ~n39110 & ~n39132;
  assign n38796 = ~n33789 & ~n33847;
  assign n27587 = ~n27586 & ~n27585;
  assign n38689 = ~n38675 & ~n27584;
  assign n36166 = ~P3_PHYADDRPOINTER_REG_26__SCAN_IN;
  assign n36320 = ~n37008;
  assign n36327 = ~P3_INSTADDRPOINTER_REG_18__SCAN_IN;
  assign n34481 = ~n37453 & ~n39110;
  assign n38788 = ~n38694 & ~n38693;
  assign n37667 = ~n37674;
  assign n26949 = n26936 | n26935;
  assign n42494 = ~n42470;
  assign n30287 = ~n42500;
  assign n42488 = ~n42440;
  assign n30097 = n26438 & n26437;
  assign n42907 = ~n42937 & ~n42944;
  assign n43001 = ~n25838;
  assign n44745 = ~n31535;
  assign n43388 = n43382 & n43381;
  assign n43867 = ~n43898 & ~P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n31582 = ~READY11_REG_SCAN_IN | ~READY1;
  assign n44546 = ~P1_STATE_REG_2__SCAN_IN;
  assign n39138 = n27605 | n39593;
  assign n33240 = n27367 & n27560;
  assign n32823 = n28966 & n28965;
  assign n31648 = ~P2_PHYADDRPOINTER_REG_7__SCAN_IN;
  assign n39678 = n27370 & n31614;
  assign n39656 = n39672;
  assign n39677 = ~n39516;
  assign n31946 = n28434 & n28433;
  assign n39725 = ~n29343;
  assign n39850 = ~n39970 & ~n40552;
  assign n32712 = ~P2_INSTADDRPOINTER_REG_24__SCAN_IN;
  assign n32373 = n39313 | n28196;
  assign n33115 = n29013 & n29012;
  assign n33125 = ~n29013 | ~n28497;
  assign n42154 = ~n41002 & ~n41789;
  assign n40452 = ~P2_INSTQUEUE_REG_0__1__SCAN_IN;
  assign n40513 = ~P2_INSTQUEUE_REG_0__5__SCAN_IN;
  assign n40582 = n40648 & n41769;
  assign n40741 = n40746 & P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n40982 = ~n41071;
  assign n40556 = ~n40435 & ~n40436;
  assign n41422 = ~n41411;
  assign n41606 = ~n41808;
  assign n41642 = ~n41856;
  assign n41693 = ~n40460 | ~n40459;
  assign n41720 = ~n40505 | ~n40504;
  assign n41740 = ~n40538 | ~n40537;
  assign n42204 = ~READY21_REG_SCAN_IN | ~READY12_REG_SCAN_IN;
  assign n41895 = ~n42204;
  assign n38681 = ~n24705 | ~n24710;
  assign n38674 = ~n24632 | ~n24593;
  assign n34405 = ~n33848 | ~n38796;
  assign n34448 = ~n33850 & ~n33849;
  assign n34492 = ~P3_EBX_REG_18__SCAN_IN;
  assign n35447 = ~P3_EBX_REG_6__SCAN_IN;
  assign n35726 = n35687 & n35800;
  assign n36881 = ~n36249;
  assign n36683 = n36681;
  assign n36666 = ~n36751 & ~n33289;
  assign n36745 = ~n36478;
  assign n38678 = n24593 & n34481;
  assign n37292 = ~n38674;
  assign n24730 = n24729 | n24728;
  assign n38483 = ~n36112 & ~n33729;
  assign n39068 = ~n39038;
  assign n39069 = ~P3_STATE2_REG_1__SCAN_IN;
  assign n37805 = ~n37813 & ~n37667;
  assign n37878 = ~n37595 & ~n37667;
  assign n38025 = ~n38776 & ~n37968;
  assign n38248 = ~n38240;
  assign n38468 = ~n38455;
  assign n38537 = ~n38568 & ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n38831 = ~P3_STATE_REG_1__SCAN_IN;
  assign n33659 = ~P3_DATAO_REG_30__SCAN_IN;
  assign n44800 = ~n44418;
  assign n26977 = n30639 & P1_STATE2_REG_1__SCAN_IN;
  assign n42440 = n42461 | n26979;
  assign n42493 = ~n42413;
  assign n31515 = n25022;
  assign n42553 = ~n42561 | ~n43190;
  assign n30984 = ~n30970;
  assign n42599 = ~n42625;
  assign n43070 = ~n42620;
  assign n42758 = ~n44843 | ~n44850;
  assign n42326 = n30984 & n30983;
  assign n42936 = ~n42907;
  assign n43053 = ~n44750 | ~n43052;
  assign n43152 = ~n42598;
  assign n43122 = ~n42610;
  assign n43137 = ~n42604;
  assign n43976 = ~n43471 & ~n43636;
  assign n43113 = ~n42615;
  assign n44327 = ~n43471 & ~n43470;
  assign n44508 = ~P1_STATE2_REG_2__SCAN_IN | ~P1_STATE2_REG_1__SCAN_IN;
  assign n44815 = ~P1_REIP_REG_1__SCAN_IN;
  assign n39160 = ~n42075;
  assign n29031 = n28454 & n28453;
  assign n39628 = n42200 | n33135;
  assign n39495 = ~n39678;
  assign n32471 = n28393 & n28392;
  assign n39898 = ~n31972 & ~n39964;
  assign n40429 = n39837 & n39836;
  assign n40249 = n40117 | n40456;
  assign n40200 = ~n40249;
  assign n29797 = ~P2_INSTADDRPOINTER_REG_31__SCAN_IN;
  assign n40294 = ~n40325;
  assign n40403 = ~n33064;
  assign n27563 = ~P2_STATE2_REG_0__SCAN_IN & ~n42111;
  assign n39140 = ~n27661 | ~n27343;
  assign n40722 = ~n40662 & ~n40654;
  assign n40806 = ~n40741;
  assign n40985 = ~n40910 & ~n40909;
  assign n41071 = n40913 | n41491;
  assign n41143 = ~n41078 & ~n41077;
  assign n41227 = ~n41172;
  assign n41477 = ~n41410 & ~n41409;
  assign n41569 = ~n41422 | ~n42177;
  assign n41562 = ~n41496 & ~n41495;
  assign n41651 = ~n41578 & ~n41577;
  assign n41715 = ~n40495 | ~n41686;
  assign n41814 = ~n41703;
  assign n41850 = ~n41733;
  assign n41870 = n40552 | n40551;
  assign n39976 = ~P2_STATE2_REG_1__SCAN_IN | ~P2_STATE2_REG_2__SCAN_IN;
  assign n39120 = ~P3_STATE2_REG_1__SCAN_IN & ~P3_STATE2_REG_2__SCAN_IN;
  assign n36183 = ~P3_PHYADDRPOINTER_REG_25__SCAN_IN;
  assign n34468 = ~n34371 & ~n34430;
  assign n34469 = ~n34445;
  assign n34459 = ~n34478 | ~P3_STATE2_REG_3__SCAN_IN;
  assign n35006 = ~n34492 & ~n34491;
  assign n35273 = ~P3_EBX_REG_12__SCAN_IN;
  assign n35353 = ~P3_EBX_REG_10__SCAN_IN;
  assign n35394 = ~n34483 & ~n34482;
  assign n35554 = ~n35661;
  assign n35789 = ~n35671;
  assign n37212 = ~n33284;
  assign n35799 = ~n35504;
  assign n35937 = ~n35812 & ~n38687;
  assign n36062 = ~P3_EAX_REG_8__SCAN_IN;
  assign n35966 = ~n36103;
  assign n36400 = n36399;
  assign n37066 = ~P3_INSTADDRPOINTER_REG_13__SCAN_IN;
  assign n36613 = ~n36490;
  assign n36743 = ~n36666;
  assign n37080 = ~P3_INSTADDRPOINTER_REG_14__SCAN_IN;
  assign n37210 = ~P3_INSTADDRPOINTER_REG_8__SCAN_IN;
  assign n37257 = ~P3_INSTADDRPOINTER_REG_6__SCAN_IN;
  assign n37349 = ~n24730 | ~n39105;
  assign n38781 = ~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN;
  assign n38570 = ~n38115;
  assign n37797 = ~n37805;
  assign n37870 = ~n37878;
  assign n37501 = ~n39029 | ~n37436;
  assign n37941 = ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN | ~n37814;
  assign n38017 = ~n38025;
  assign n38087 = ~n38099;
  assign n38240 = ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN | ~n38114;
  assign n38308 = ~n38320;
  assign n38340 = ~n38489;
  assign n38545 = ~n38537;
  assign n38534 = ~n38548;
  assign n38654 = ~n38458;
  assign n38814 = ~n38803 | ~P3_STATE2_REG_3__SCAN_IN;
  assign n38811 = ~n39120;
  assign n39114 = ~READY22_REG_SCAN_IN | ~READY2;
  assign n38890 = ~P3_REIP_REG_7__SCAN_IN;
  assign n38854 = ~P3_STATE_REG_0__SCAN_IN;
  assign n33487 = n33538 | n33460;
  assign n33660 = ~P3_DATAO_REG_31__SCAN_IN & ~n33659;
  assign n42759 = ~n42227 & ~n26962;
  assign n42234 = n44800 & n31580;
  assign n42373 = ~n42469 | ~n26977;
  assign n42389 = ~n42367;
  assign n42481 = n26998 & n26997;
  assign n42562 = ~n42540;
  assign n42540 = n42561 & n31515;
  assign n42556 = ~n42561;
  assign n30536 = ~n30765;
  assign n42592 = ~n42625 & ~n30603;
  assign n42749 = n42755;
  assign n42891 = ~n42759 | ~n42758;
  assign n43018 = ~n25684 | ~n25683;
  assign n44809 = ~n44808;
  assign n44741 = ~n44757;
  assign n43198 = ~n43080 | ~n43079;
  assign n43290 = ~n43224 | ~n43223;
  assign n43458 = ~n43386 | ~n43385;
  assign n43629 = ~n43563 | ~n43562;
  assign n43708 = ~n43654 | ~n43653;
  assign n43796 = ~n43736 | ~n43735;
  assign n43960 = ~n43900 | ~n43899;
  assign n44129 = ~n44064 | ~n44063;
  assign n44303 = ~n44243 | ~n44242;
  assign n44505 = ~n44421 | ~n44420;
  assign n42243 = n42232 | n44522;
  assign n42200 = ~n33223 | ~n39141;
  assign n42075 = ~n27368 | ~P2_STATE2_REG_2__SCAN_IN;
  assign n39681 = n42200 | n31594;
  assign n39686 = ~n39628;
  assign n39639 = ~n39681;
  assign n39647 = ~n41893;
  assign n39817 = ~n31948;
  assign n39954 = ~n39962;
  assign n40037 = ~n40077 & ~n42209;
  assign n42199 = n40022;
  assign n40108 = ~n40111 & ~n42199;
  assign n40324 = ~n40344;
  assign n40337 = n39163 & n29852;
  assign n41786 = ~n27564 & ~n27563;
  assign n40645 = ~n40585 | ~n41686;
  assign n40904 = ~n40843 | ~n40842;
  assign n40981 = ~n40926 | ~n40925;
  assign n41068 = n42139 & n41491;
  assign n41151 = ~n41092 | ~n41091;
  assign n41318 = ~n41259 | ~n41258;
  assign n41486 = ~n41426 | ~n41425;
  assign n41563 = ~n41511 | ~n41510;
  assign n41660 = ~n41594 | ~n41593;
  assign n42181 = ~n39976;
  assign n41926 = ~P2_STATE_REG_2__SCAN_IN;
  assign n42065 = ~n41920 | ~P2_STATE_REG_1__SCAN_IN;
  assign n38799 = ~P3_STATE2_REG_2__SCAN_IN | ~n38815;
  assign n34291 = n34371 | n34286;
  assign n34478 = ~n33796 | ~n38808;
  assign n34843 = n34805 | n34851;
  assign n35391 = ~n35477;
  assign n35477 = ~n35490 & ~n34971;
  assign n35490 = ~n35394;
  assign n35661 = ~n35671 & ~n37502;
  assign n35807 = ~n27590 & ~n35799;
  assign n35872 = n35815 & n35937;
  assign n35909 = ~n39106 & ~n35937;
  assign n36580 = ~n36629;
  assign n36629 = n36727 & n33284;
  assign n36727 = ~n33749 & ~n37453;
  assign n37201 = ~n37349 & ~n33406;
  assign n37352 = ~n37383;
  assign n38489 = ~n39118 | ~n37436;
  assign n38476 = ~n38814;
  assign n37396 = ~P3_STATE2_REG_1__SCAN_IN | ~P3_STATE2_REG_2__SCAN_IN;
  assign n39097 = ~n38854 | ~P3_STATE_REG_1__SCAN_IN;
  assign n39126 = ~n39097;
  assign n33588 = ~U212;
  assign n44859 = n44522 & P1_STATE_REG_1__SCAN_IN;
  assign n43055 = ~P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN;
  assign n44521 = ~n44828 | ~n42243;
  assign n39163 = n33245 | n42075;
  assign n39977 = ~P2_DATAO_REG_31__SCAN_IN;
  assign n40076 = ~n40108;
  assign n33749 = n38668 | n38799;
  assign n35940 = n35909;
  assign n38686 = ~P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN;
  assign n43060 = ~n43062;
  assign U214 = ~n43060 | ~n27017;
  assign n23981 = ~n23065 | ~P3_INSTQUEUE_REG_3__1__SCAN_IN;
  assign n24289 = n24000 & n38725;
  assign n23980 = ~n24289 | ~P3_INSTQUEUE_REG_4__1__SCAN_IN;
  assign n23983 = n23981 & n23980;
  assign n24373 = ~n23999 & ~n24010;
  assign n23982 = ~n24373 | ~P3_INSTQUEUE_REG_14__1__SCAN_IN;
  assign n23986 = ~n23983 | ~n23982;
  assign n23984 = ~P3_INSTQUEUE_REG_7__1__SCAN_IN;
  assign n23985 = ~n24522 & ~n23984;
  assign n23989 = ~n24315 | ~P3_INSTQUEUE_REG_15__1__SCAN_IN;
  assign n23987 = ~n24010;
  assign n23988 = ~n24318 | ~P3_INSTQUEUE_REG_13__1__SCAN_IN;
  assign n23993 = ~n23989 | ~n23988;
  assign n34516 = n24005 & n34451;
  assign n23991 = ~n34516 | ~P3_INSTQUEUE_REG_5__1__SCAN_IN;
  assign n34575 = n24000 & n34451;
  assign n23990 = ~n34575 | ~P3_INSTQUEUE_REG_1__1__SCAN_IN;
  assign n23992 = ~n23991 | ~n23990;
  assign n23994 = ~n23993 & ~n23992;
  assign n24018 = ~n23995 | ~n23994;
  assign n23998 = ~n24191 | ~P3_INSTQUEUE_REG_12__1__SCAN_IN;
  assign n23996 = ~n38719 | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign n34578 = ~n34396 & ~n23996;
  assign n23997 = ~n34578 | ~P3_INSTQUEUE_REG_11__1__SCAN_IN;
  assign n24004 = ~n23998 | ~n23997;
  assign n24002 = ~n24292 | ~P3_INSTQUEUE_REG_10__1__SCAN_IN;
  assign n34660 = n24006 & n24000;
  assign n24001 = ~n34660 | ~P3_INSTQUEUE_REG_2__1__SCAN_IN;
  assign n24003 = ~n24002 | ~n24001;
  assign n24016 = ~n24004 & ~n24003;
  assign n24008 = ~n24300 | ~P3_INSTQUEUE_REG_6__1__SCAN_IN;
  assign n24301 = ~n38728 & ~n38723;
  assign n24007 = ~n24301 | ~P3_INSTQUEUE_REG_8__1__SCAN_IN;
  assign n24014 = ~n24008 | ~n24007;
  assign n34532 = n24009 & n34451;
  assign n24012 = ~n34532 | ~P3_INSTQUEUE_REG_9__1__SCAN_IN;
  assign n24308 = ~n38723 & ~n24010;
  assign n24011 = ~n24308 | ~P3_INSTQUEUE_REG_0__1__SCAN_IN;
  assign n24013 = ~n24012 | ~n24011;
  assign n24015 = ~n24014 & ~n24013;
  assign n24017 = ~n24016 | ~n24015;
  assign n36732 = ~n24569 ^ P3_INSTADDRPOINTER_REG_1__SCAN_IN;
  assign n24020 = ~n24301 | ~P3_INSTQUEUE_REG_8__0__SCAN_IN;
  assign n24019 = ~n24191 | ~P3_INSTQUEUE_REG_12__0__SCAN_IN;
  assign n24022 = ~n24020 | ~n24019;
  assign n24025 = n24022 | n24021;
  assign n24023 = ~P3_INSTQUEUE_REG_7__0__SCAN_IN;
  assign n24024 = ~n24522 & ~n24023;
  assign n24048 = ~n24025 & ~n24024;
  assign n24027 = ~n24300 | ~P3_INSTQUEUE_REG_6__0__SCAN_IN;
  assign n24026 = ~n24318 | ~P3_INSTQUEUE_REG_13__0__SCAN_IN;
  assign n24031 = ~n24027 | ~n24026;
  assign n24029 = ~n24292 | ~P3_INSTQUEUE_REG_10__0__SCAN_IN;
  assign n24028 = ~n23065 | ~P3_INSTQUEUE_REG_3__0__SCAN_IN;
  assign n24030 = ~n24029 | ~n24028;
  assign n24039 = ~n24031 & ~n24030;
  assign n24033 = ~n34578 | ~P3_INSTQUEUE_REG_11__0__SCAN_IN;
  assign n24032 = ~n34660 | ~P3_INSTQUEUE_REG_2__0__SCAN_IN;
  assign n24037 = ~n24033 | ~n24032;
  assign n24035 = ~n24289 | ~P3_INSTQUEUE_REG_4__0__SCAN_IN;
  assign n24034 = ~n24308 | ~P3_INSTQUEUE_REG_0__0__SCAN_IN;
  assign n24036 = ~n24035 | ~n24034;
  assign n24038 = ~n24037 & ~n24036;
  assign n24046 = ~n24039 | ~n24038;
  assign n24041 = ~n34516 | ~P3_INSTQUEUE_REG_5__0__SCAN_IN;
  assign n24040 = ~n34532 | ~P3_INSTQUEUE_REG_9__0__SCAN_IN;
  assign n24045 = ~n24041 | ~n24040;
  assign n24043 = ~n24373 | ~P3_INSTQUEUE_REG_14__0__SCAN_IN;
  assign n24042 = ~n34575 | ~P3_INSTQUEUE_REG_1__0__SCAN_IN;
  assign n24044 = ~n24043 | ~n24042;
  assign n36749 = n27595 & P3_INSTADDRPOINTER_REG_0__SCAN_IN;
  assign n35804 = ~n24569;
  assign n24572 = ~n35804 | ~P3_INSTADDRPOINTER_REG_1__SCAN_IN;
  assign n24050 = ~n23065 | ~P3_INSTQUEUE_REG_3__2__SCAN_IN;
  assign n24049 = ~n24289 | ~P3_INSTQUEUE_REG_4__2__SCAN_IN;
  assign n24052 = n24050 & n24049;
  assign n24051 = ~n24373 | ~P3_INSTQUEUE_REG_14__2__SCAN_IN;
  assign n24055 = ~n24052 | ~n24051;
  assign n24053 = ~P3_INSTQUEUE_REG_7__2__SCAN_IN;
  assign n24054 = ~n24522 & ~n24053;
  assign n24063 = ~n24055 & ~n24054;
  assign n24057 = ~n24315 | ~P3_INSTQUEUE_REG_15__2__SCAN_IN;
  assign n24107 = ~n24318;
  assign n35415 = ~n24107;
  assign n24056 = ~n35415 | ~P3_INSTQUEUE_REG_13__2__SCAN_IN;
  assign n24061 = ~n24057 | ~n24056;
  assign n24059 = ~n34516 | ~P3_INSTQUEUE_REG_5__2__SCAN_IN;
  assign n24058 = ~n34575 | ~P3_INSTQUEUE_REG_1__2__SCAN_IN;
  assign n24060 = ~n24059 | ~n24058;
  assign n24062 = ~n24061 & ~n24060;
  assign n24079 = ~n24063 | ~n24062;
  assign n24065 = ~n24191 | ~P3_INSTQUEUE_REG_12__2__SCAN_IN;
  assign n24064 = ~n34578 | ~P3_INSTQUEUE_REG_11__2__SCAN_IN;
  assign n24069 = ~n24065 | ~n24064;
  assign n24067 = ~n24292 | ~P3_INSTQUEUE_REG_10__2__SCAN_IN;
  assign n24066 = ~n34660 | ~P3_INSTQUEUE_REG_2__2__SCAN_IN;
  assign n24068 = ~n24067 | ~n24066;
  assign n24077 = ~n24069 & ~n24068;
  assign n24098 = ~n24300;
  assign n35422 = ~n24098;
  assign n24071 = ~n24300 | ~P3_INSTQUEUE_REG_6__2__SCAN_IN;
  assign n24070 = ~n24301 | ~P3_INSTQUEUE_REG_8__2__SCAN_IN;
  assign n24075 = ~n24071 | ~n24070;
  assign n24073 = ~n34532 | ~P3_INSTQUEUE_REG_9__2__SCAN_IN;
  assign n24072 = ~n24308 | ~P3_INSTQUEUE_REG_0__2__SCAN_IN;
  assign n24074 = ~n24073 | ~n24072;
  assign n24076 = ~n24075 & ~n24074;
  assign n24078 = ~n24077 | ~n24076;
  assign n24552 = n24079 | n24078;
  assign n24567 = ~P3_INSTADDRPOINTER_REG_2__SCAN_IN;
  assign n24081 = n24080 | n24567;
  assign n36707 = ~n24082 | ~n24081;
  assign n24564 = n24552 & n24569;
  assign n24084 = ~n23065 | ~P3_INSTQUEUE_REG_3__3__SCAN_IN;
  assign n24083 = ~n24308 | ~P3_INSTQUEUE_REG_0__3__SCAN_IN;
  assign n24086 = n24084 & n24083;
  assign n24085 = ~n24540 | ~P3_INSTQUEUE_REG_8__3__SCAN_IN;
  assign n24089 = ~n24086 | ~n24085;
  assign n24087 = ~P3_INSTQUEUE_REG_7__3__SCAN_IN;
  assign n24088 = ~n24522 & ~n24087;
  assign n24097 = ~n24089 & ~n24088;
  assign n24091 = ~n34578 | ~P3_INSTQUEUE_REG_11__3__SCAN_IN;
  assign n24090 = ~n34532 | ~P3_INSTQUEUE_REG_9__3__SCAN_IN;
  assign n24095 = ~n24091 | ~n24090;
  assign n24093 = ~n34575 | ~P3_INSTQUEUE_REG_1__3__SCAN_IN;
  assign n24092 = ~n24289 | ~P3_INSTQUEUE_REG_4__3__SCAN_IN;
  assign n24094 = ~n24093 | ~n24092;
  assign n24096 = ~n24095 & ~n24094;
  assign n24115 = ~n24097 | ~n24096;
  assign n24100 = ~n24300 | ~P3_INSTQUEUE_REG_6__3__SCAN_IN;
  assign n24099 = ~n24292 | ~P3_INSTQUEUE_REG_10__3__SCAN_IN;
  assign n24104 = ~n24100 | ~n24099;
  assign n24102 = ~n24373 | ~P3_INSTQUEUE_REG_14__3__SCAN_IN;
  assign n24101 = ~n34516 | ~P3_INSTQUEUE_REG_5__3__SCAN_IN;
  assign n24103 = ~n24102 | ~n24101;
  assign n24113 = ~n24104 & ~n24103;
  assign n24106 = ~n24315 | ~P3_INSTQUEUE_REG_15__3__SCAN_IN;
  assign n24105 = ~n24191 | ~P3_INSTQUEUE_REG_12__3__SCAN_IN;
  assign n24111 = ~n24106 | ~n24105;
  assign n24109 = ~n34660 | ~P3_INSTQUEUE_REG_2__3__SCAN_IN;
  assign n24108 = ~n24318 | ~P3_INSTQUEUE_REG_13__3__SCAN_IN;
  assign n24110 = ~n24109 | ~n24108;
  assign n24112 = ~n24111 & ~n24110;
  assign n24114 = ~n24113 | ~n24112;
  assign n35782 = n24115 | n24114;
  assign n24119 = ~n36707 | ~n36706;
  assign n24117 = ~n24116;
  assign n24118 = ~n24117 | ~P3_INSTADDRPOINTER_REG_3__SCAN_IN;
  assign n36681 = ~n24119 | ~n24118;
  assign n24121 = ~n23065 | ~P3_INSTQUEUE_REG_3__4__SCAN_IN;
  assign n24120 = ~n24289 | ~P3_INSTQUEUE_REG_4__4__SCAN_IN;
  assign n24123 = n24121 & n24120;
  assign n24122 = ~n24373 | ~P3_INSTQUEUE_REG_14__4__SCAN_IN;
  assign n24126 = ~n24123 | ~n24122;
  assign n24124 = ~P3_INSTQUEUE_REG_7__4__SCAN_IN;
  assign n24125 = ~n24522 & ~n24124;
  assign n24134 = ~n24126 & ~n24125;
  assign n24128 = ~n24315 | ~P3_INSTQUEUE_REG_15__4__SCAN_IN;
  assign n24127 = ~n35415 | ~P3_INSTQUEUE_REG_13__4__SCAN_IN;
  assign n24132 = ~n24128 | ~n24127;
  assign n24130 = ~n34516 | ~P3_INSTQUEUE_REG_5__4__SCAN_IN;
  assign n24129 = ~n34575 | ~P3_INSTQUEUE_REG_1__4__SCAN_IN;
  assign n24131 = ~n24130 | ~n24129;
  assign n24133 = ~n24132 & ~n24131;
  assign n24136 = ~n24191 | ~P3_INSTQUEUE_REG_12__4__SCAN_IN;
  assign n24135 = ~n34578 | ~P3_INSTQUEUE_REG_11__4__SCAN_IN;
  assign n24140 = ~n24136 | ~n24135;
  assign n24138 = ~n24292 | ~P3_INSTQUEUE_REG_10__4__SCAN_IN;
  assign n24137 = ~n34660 | ~P3_INSTQUEUE_REG_2__4__SCAN_IN;
  assign n24139 = ~n24138 | ~n24137;
  assign n24148 = ~n24140 & ~n24139;
  assign n24142 = ~n35422 | ~P3_INSTQUEUE_REG_6__4__SCAN_IN;
  assign n35396 = ~n22844;
  assign n24141 = ~n35396 | ~P3_INSTQUEUE_REG_8__4__SCAN_IN;
  assign n24146 = ~n24142 | ~n24141;
  assign n24144 = ~n34532 | ~P3_INSTQUEUE_REG_9__4__SCAN_IN;
  assign n24143 = ~n24308 | ~P3_INSTQUEUE_REG_0__4__SCAN_IN;
  assign n24145 = ~n24144 | ~n24143;
  assign n24147 = ~n24146 & ~n24145;
  assign n24151 = ~n24188 ^ n35773;
  assign n36682 = ~n24151 ^ P3_INSTADDRPOINTER_REG_4__SCAN_IN;
  assign n24152 = ~n24151;
  assign n24153 = ~n24152 | ~P3_INSTADDRPOINTER_REG_4__SCAN_IN;
  assign n24182 = ~n24188 & ~n35773;
  assign n24155 = ~n34660 | ~P3_INSTQUEUE_REG_2__5__SCAN_IN;
  assign n24154 = ~n24289 | ~P3_INSTQUEUE_REG_4__5__SCAN_IN;
  assign n24157 = ~n24155 | ~n24154;
  assign n24156 = n24315 & P3_INSTQUEUE_REG_15__5__SCAN_IN;
  assign n24160 = ~n24157 & ~n24156;
  assign n24158 = ~P3_INSTQUEUE_REG_7__5__SCAN_IN;
  assign n24159 = n24522 | n24158;
  assign n24168 = ~n24160 | ~n24159;
  assign n24162 = ~n24292 | ~P3_INSTQUEUE_REG_10__5__SCAN_IN;
  assign n24161 = ~n24373 | ~P3_INSTQUEUE_REG_14__5__SCAN_IN;
  assign n24166 = n24162 & n24161;
  assign n24164 = ~n35422 | ~P3_INSTQUEUE_REG_6__5__SCAN_IN;
  assign n24163 = ~n23065 | ~P3_INSTQUEUE_REG_3__5__SCAN_IN;
  assign n24165 = n24164 & n24163;
  assign n24167 = ~n24166 | ~n24165;
  assign n24181 = ~n24168 & ~n24167;
  assign n24170 = ~n24191 | ~P3_INSTQUEUE_REG_12__5__SCAN_IN;
  assign n24169 = ~n34578 | ~P3_INSTQUEUE_REG_11__5__SCAN_IN;
  assign n24171 = ~n24170 | ~n24169;
  assign n24173 = ~n35396 | ~P3_INSTQUEUE_REG_8__5__SCAN_IN;
  assign n24172 = ~n35415 | ~P3_INSTQUEUE_REG_13__5__SCAN_IN;
  assign n24177 = ~n24173 | ~n24172;
  assign n24175 = ~n34516 | ~P3_INSTQUEUE_REG_5__5__SCAN_IN;
  assign n24174 = ~n34575 | ~P3_INSTQUEUE_REG_1__5__SCAN_IN;
  assign n24176 = ~n24175 | ~n24174;
  assign n24178 = ~n24177 & ~n24176;
  assign n35761 = n24181 & n24180;
  assign n24185 = ~n24182 ^ n35761;
  assign n24221 = ~n24188 & ~n24187;
  assign n24190 = ~n35396 | ~P3_INSTQUEUE_REG_8__6__SCAN_IN;
  assign n24189 = ~n34575 | ~P3_INSTQUEUE_REG_1__6__SCAN_IN;
  assign n24195 = ~n24190 | ~n24189;
  assign n24193 = ~n24513 | ~P3_INSTQUEUE_REG_11__6__SCAN_IN;
  assign n24192 = ~n34717 | ~P3_INSTQUEUE_REG_12__6__SCAN_IN;
  assign n24194 = ~n24193 | ~n24192;
  assign n24203 = ~n24195 & ~n24194;
  assign n24197 = ~n24470 | ~P3_INSTQUEUE_REG_3__6__SCAN_IN;
  assign n24196 = ~n24289 | ~P3_INSTQUEUE_REG_4__6__SCAN_IN;
  assign n24201 = ~n24197 | ~n24196;
  assign n24199 = ~n35412 | ~P3_INSTQUEUE_REG_7__6__SCAN_IN;
  assign n24198 = ~n34872 | ~P3_INSTQUEUE_REG_15__6__SCAN_IN;
  assign n24200 = ~n24199 | ~n24198;
  assign n24202 = ~n24201 & ~n24200;
  assign n24205 = ~n35422 | ~P3_INSTQUEUE_REG_6__6__SCAN_IN;
  assign n24204 = ~n35328 | ~P3_INSTQUEUE_REG_2__6__SCAN_IN;
  assign n24209 = ~n24205 | ~n24204;
  assign n24207 = ~n24292 | ~P3_INSTQUEUE_REG_10__6__SCAN_IN;
  assign n24206 = ~n34532 | ~P3_INSTQUEUE_REG_9__6__SCAN_IN;
  assign n24208 = ~n24207 | ~n24206;
  assign n24217 = ~n24209 & ~n24208;
  assign n24211 = ~n35252 | ~P3_INSTQUEUE_REG_14__6__SCAN_IN;
  assign n24210 = ~n35415 | ~P3_INSTQUEUE_REG_13__6__SCAN_IN;
  assign n24215 = ~n24211 | ~n24210;
  assign n24213 = ~n24543 | ~P3_INSTQUEUE_REG_5__6__SCAN_IN;
  assign n24212 = ~n34564 | ~P3_INSTQUEUE_REG_0__6__SCAN_IN;
  assign n24214 = ~n24213 | ~n24212;
  assign n24216 = ~n24215 & ~n24214;
  assign n24223 = ~n24470 | ~P3_INSTQUEUE_REG_3__7__SCAN_IN;
  assign n24222 = ~n24289 | ~P3_INSTQUEUE_REG_4__7__SCAN_IN;
  assign n24225 = n24223 & n24222;
  assign n24224 = ~n35252 | ~P3_INSTQUEUE_REG_14__7__SCAN_IN;
  assign n24228 = ~n24225 | ~n24224;
  assign n24226 = ~P3_INSTQUEUE_REG_7__7__SCAN_IN;
  assign n24227 = ~n24522 & ~n24226;
  assign n24236 = ~n24228 & ~n24227;
  assign n24230 = ~n35396 | ~P3_INSTQUEUE_REG_8__7__SCAN_IN;
  assign n24229 = ~n35319 | ~P3_INSTQUEUE_REG_9__7__SCAN_IN;
  assign n24234 = ~n24230 | ~n24229;
  assign n24232 = ~n34872 | ~P3_INSTQUEUE_REG_15__7__SCAN_IN;
  assign n24231 = ~n35415 | ~P3_INSTQUEUE_REG_13__7__SCAN_IN;
  assign n24233 = ~n24232 | ~n24231;
  assign n24235 = ~n24234 & ~n24233;
  assign n24252 = ~n24236 | ~n24235;
  assign n24238 = ~n24292 | ~P3_INSTQUEUE_REG_10__7__SCAN_IN;
  assign n24237 = ~n24513 | ~P3_INSTQUEUE_REG_11__7__SCAN_IN;
  assign n24242 = ~n24238 | ~n24237;
  assign n24240 = ~n34717 | ~P3_INSTQUEUE_REG_12__7__SCAN_IN;
  assign n24239 = ~n35359 | ~P3_INSTQUEUE_REG_0__7__SCAN_IN;
  assign n24241 = ~n24240 | ~n24239;
  assign n24250 = ~n24242 & ~n24241;
  assign n24244 = ~n35422 | ~P3_INSTQUEUE_REG_6__7__SCAN_IN;
  assign n24243 = ~n35328 | ~P3_INSTQUEUE_REG_2__7__SCAN_IN;
  assign n24248 = ~n24244 | ~n24243;
  assign n24246 = ~n24543 | ~P3_INSTQUEUE_REG_5__7__SCAN_IN;
  assign n24245 = ~n35405 | ~P3_INSTQUEUE_REG_1__7__SCAN_IN;
  assign n24247 = ~n24246 | ~n24245;
  assign n24249 = ~n24248 & ~n24247;
  assign n24251 = ~n24250 | ~n24249;
  assign n24254 = ~n33408 ^ n37212;
  assign n24256 = ~n24255 | ~n24254;
  assign n24257 = ~n36610 | ~n37210;
  assign n37121 = ~P3_INSTADDRPOINTER_REG_9__SCAN_IN | ~P3_INSTADDRPOINTER_REG_10__SCAN_IN;
  assign n37154 = ~P3_INSTADDRPOINTER_REG_11__SCAN_IN;
  assign n37065 = ~n37121 & ~n37154;
  assign n24258 = ~n37065;
  assign n36437 = P3_INSTADDRPOINTER_REG_13__SCAN_IN & P3_INSTADDRPOINTER_REG_12__SCAN_IN;
  assign n24259 = n24595 & n36437;
  assign n24265 = ~n36515 | ~n24259;
  assign n36574 = ~P3_INSTADDRPOINTER_REG_10__SCAN_IN & ~P3_INSTADDRPOINTER_REG_9__SCAN_IN;
  assign n36432 = ~P3_INSTADDRPOINTER_REG_12__SCAN_IN & ~P3_INSTADDRPOINTER_REG_11__SCAN_IN;
  assign n24262 = ~n36574 | ~n36432;
  assign n24260 = ~P3_INSTADDRPOINTER_REG_13__SCAN_IN & ~P3_INSTADDRPOINTER_REG_15__SCAN_IN;
  assign n24261 = ~n24260 | ~n37080;
  assign n24263 = ~n24262 & ~n24261;
  assign n24264 = ~n36498 | ~n24263;
  assign n24267 = ~n36419 | ~P3_INSTADDRPOINTER_REG_16__SCAN_IN;
  assign n24266 = n36610 | P3_INSTADDRPOINTER_REG_16__SCAN_IN;
  assign n24268 = ~n24267 | ~n24266;
  assign n24270 = ~n36399;
  assign n24269 = ~P3_INSTADDRPOINTER_REG_17__SCAN_IN;
  assign n24271 = ~n24270 | ~n24269;
  assign n24272 = P3_INSTADDRPOINTER_REG_16__SCAN_IN & P3_INSTADDRPOINTER_REG_17__SCAN_IN;
  assign n24273 = ~n36419 | ~n24272;
  assign n36322 = P3_INSTADDRPOINTER_REG_19__SCAN_IN & P3_INSTADDRPOINTER_REG_18__SCAN_IN;
  assign n24629 = P3_INSTADDRPOINTER_REG_20__SCAN_IN & P3_INSTADDRPOINTER_REG_21__SCAN_IN;
  assign n36874 = ~n36322 | ~n24629;
  assign n24274 = ~n36874;
  assign n24596 = ~P3_INSTADDRPOINTER_REG_23__SCAN_IN | ~P3_INSTADDRPOINTER_REG_22__SCAN_IN;
  assign n36298 = ~P3_INSTADDRPOINTER_REG_19__SCAN_IN & ~P3_INSTADDRPOINTER_REG_20__SCAN_IN;
  assign n24275 = ~n36298 | ~n36327;
  assign n24276 = P3_INSTADDRPOINTER_REG_21__SCAN_IN | n24275;
  assign n36276 = ~n36610 & ~n24276;
  assign n24277 = ~P3_INSTADDRPOINTER_REG_22__SCAN_IN & ~P3_INSTADDRPOINTER_REG_23__SCAN_IN;
  assign n24278 = ~n36276 | ~n24277;
  assign n24280 = ~n36191 | ~P3_INSTADDRPOINTER_REG_25__SCAN_IN;
  assign n24279 = n36610 | P3_INSTADDRPOINTER_REG_25__SCAN_IN;
  assign n24281 = ~n24280 | ~n24279;
  assign n36193 = ~n36215 | ~n36497;
  assign n24282 = ~P3_INSTADDRPOINTER_REG_26__SCAN_IN;
  assign n36781 = ~P3_INSTADDRPOINTER_REG_26__SCAN_IN | ~P3_INSTADDRPOINTER_REG_25__SCAN_IN;
  assign n24641 = ~n36781;
  assign n36764 = ~P3_INSTADDRPOINTER_REG_27__SCAN_IN;
  assign n24285 = ~n33331 & ~n36610;
  assign n36134 = ~n24285 & ~n36151;
  assign n33399 = ~P3_INSTADDRPOINTER_REG_29__SCAN_IN;
  assign n33267 = ~n36134 | ~n33399;
  assign n33276 = ~n33267 & ~n36610;
  assign n33426 = ~n36151 | ~n36610;
  assign n24286 = ~P3_INSTADDRPOINTER_REG_29__SCAN_IN | ~P3_INSTADDRPOINTER_REG_28__SCAN_IN;
  assign n33268 = ~n33426 & ~n24286;
  assign n24288 = ~n33276 & ~n33268;
  assign n33306 = ~n24288 ^ n24287;
  assign n24470 = ~n34779;
  assign n24291 = ~n24470 | ~P3_INSTQUEUE_REG_2__2__SCAN_IN;
  assign n24290 = ~n34993 | ~P3_INSTQUEUE_REG_3__2__SCAN_IN;
  assign n24296 = ~n24291 | ~n24290;
  assign n24451 = ~n34631;
  assign n24294 = ~n24451 | ~P3_INSTQUEUE_REG_9__2__SCAN_IN;
  assign n24293 = ~n35328 | ~P3_INSTQUEUE_REG_1__2__SCAN_IN;
  assign n24295 = ~n24294 | ~n24293;
  assign n24307 = ~n24296 & ~n24295;
  assign n24299 = ~n24513 | ~P3_INSTQUEUE_REG_10__2__SCAN_IN;
  assign n24298 = ~n34717 | ~P3_INSTQUEUE_REG_11__2__SCAN_IN;
  assign n24305 = ~n24299 | ~n24298;
  assign n24303 = ~n24535 | ~P3_INSTQUEUE_REG_5__2__SCAN_IN;
  assign n24540 = ~n22844;
  assign n24302 = ~n24540 | ~P3_INSTQUEUE_REG_7__2__SCAN_IN;
  assign n24304 = ~n24303 | ~n24302;
  assign n24306 = ~n24305 & ~n24304;
  assign n24326 = ~n24307 | ~n24306;
  assign n24310 = ~n35319 | ~P3_INSTQUEUE_REG_8__2__SCAN_IN;
  assign n24309 = ~n34564 | ~P3_INSTQUEUE_REG_15__2__SCAN_IN;
  assign n24314 = ~n24310 | ~n24309;
  assign n24543 = n34516;
  assign n24312 = ~n24543 | ~P3_INSTQUEUE_REG_4__2__SCAN_IN;
  assign n24311 = ~n35405 | ~P3_INSTQUEUE_REG_0__2__SCAN_IN;
  assign n24313 = ~n24312 | ~n24311;
  assign n24324 = ~n24314 & ~n24313;
  assign n24317 = ~n35412 | ~P3_INSTQUEUE_REG_6__2__SCAN_IN;
  assign n24316 = ~n24315 | ~P3_INSTQUEUE_REG_14__2__SCAN_IN;
  assign n24322 = ~n24317 | ~n24316;
  assign n24320 = ~n35252 | ~P3_INSTQUEUE_REG_13__2__SCAN_IN;
  assign n24516 = ~n34782;
  assign n24319 = ~n24516 | ~P3_INSTQUEUE_REG_12__2__SCAN_IN;
  assign n24321 = ~n24320 | ~n24319;
  assign n24323 = ~n24322 & ~n24321;
  assign n24325 = ~n24324 | ~n24323;
  assign n24328 = ~n24451 | ~P3_INSTQUEUE_REG_9__4__SCAN_IN;
  assign n24327 = ~n34717 | ~P3_INSTQUEUE_REG_11__4__SCAN_IN;
  assign n24332 = ~n24328 | ~n24327;
  assign n24330 = ~n24535 | ~P3_INSTQUEUE_REG_5__4__SCAN_IN;
  assign n24329 = ~n24470 | ~P3_INSTQUEUE_REG_2__4__SCAN_IN;
  assign n24331 = ~n24330 | ~n24329;
  assign n24340 = ~n24332 & ~n24331;
  assign n24334 = ~n35412 | ~P3_INSTQUEUE_REG_6__4__SCAN_IN;
  assign n24333 = ~n34872 | ~P3_INSTQUEUE_REG_14__4__SCAN_IN;
  assign n24338 = ~n24334 | ~n24333;
  assign n24336 = ~n35319 | ~P3_INSTQUEUE_REG_8__4__SCAN_IN;
  assign n24335 = ~n24516 | ~P3_INSTQUEUE_REG_12__4__SCAN_IN;
  assign n24337 = ~n24336 | ~n24335;
  assign n24339 = ~n24338 & ~n24337;
  assign n24356 = ~n24340 | ~n24339;
  assign n24342 = ~n24540 | ~P3_INSTQUEUE_REG_7__4__SCAN_IN;
  assign n24341 = ~n24513 | ~P3_INSTQUEUE_REG_10__4__SCAN_IN;
  assign n24346 = ~n24342 | ~n24341;
  assign n24344 = ~n35328 | ~P3_INSTQUEUE_REG_1__4__SCAN_IN;
  assign n24343 = ~n34993 | ~P3_INSTQUEUE_REG_3__4__SCAN_IN;
  assign n24345 = ~n24344 | ~n24343;
  assign n24354 = ~n24346 & ~n24345;
  assign n24348 = ~n35252 | ~P3_INSTQUEUE_REG_13__4__SCAN_IN;
  assign n24347 = ~n34575 | ~P3_INSTQUEUE_REG_0__4__SCAN_IN;
  assign n24352 = ~n24348 | ~n24347;
  assign n24350 = ~n24543 | ~P3_INSTQUEUE_REG_4__4__SCAN_IN;
  assign n24349 = ~n34564 | ~P3_INSTQUEUE_REG_15__4__SCAN_IN;
  assign n24351 = ~n24350 | ~n24349;
  assign n24353 = ~n24352 & ~n24351;
  assign n24355 = ~n24354 | ~n24353;
  assign n24482 = ~n37463 | ~n37482;
  assign n24358 = ~n24516 | ~P3_INSTQUEUE_REG_12__5__SCAN_IN;
  assign n24357 = ~n34564 | ~P3_INSTQUEUE_REG_15__5__SCAN_IN;
  assign n24362 = ~n24358 | ~n24357;
  assign n24360 = ~n24513 | ~P3_INSTQUEUE_REG_10__5__SCAN_IN;
  assign n24359 = ~n34717 | ~P3_INSTQUEUE_REG_11__5__SCAN_IN;
  assign n24361 = ~n24360 | ~n24359;
  assign n24370 = ~n24362 & ~n24361;
  assign n24364 = ~n34872 | ~P3_INSTQUEUE_REG_14__5__SCAN_IN;
  assign n24363 = ~n34575 | ~P3_INSTQUEUE_REG_0__5__SCAN_IN;
  assign n24368 = ~n24364 | ~n24363;
  assign n24366 = ~n35412 | ~P3_INSTQUEUE_REG_6__5__SCAN_IN;
  assign n24365 = ~n34545 | ~P3_INSTQUEUE_REG_5__5__SCAN_IN;
  assign n24367 = ~n24366 | ~n24365;
  assign n24369 = ~n24368 & ~n24367;
  assign n24387 = ~n24370 | ~n24369;
  assign n24372 = ~n24540 | ~P3_INSTQUEUE_REG_7__5__SCAN_IN;
  assign n24371 = ~n35319 | ~P3_INSTQUEUE_REG_8__5__SCAN_IN;
  assign n24377 = ~n24372 | ~n24371;
  assign n24375 = ~n35252 | ~P3_INSTQUEUE_REG_13__5__SCAN_IN;
  assign n24374 = ~n24543 | ~P3_INSTQUEUE_REG_4__5__SCAN_IN;
  assign n24376 = ~n24375 | ~n24374;
  assign n24385 = ~n24377 & ~n24376;
  assign n24379 = ~n24451 | ~P3_INSTQUEUE_REG_9__5__SCAN_IN;
  assign n24378 = ~n35328 | ~P3_INSTQUEUE_REG_1__5__SCAN_IN;
  assign n24383 = ~n24379 | ~n24378;
  assign n24381 = ~n24470 | ~P3_INSTQUEUE_REG_2__5__SCAN_IN;
  assign n24380 = ~n34993 | ~P3_INSTQUEUE_REG_3__5__SCAN_IN;
  assign n24382 = ~n24381 | ~n24380;
  assign n24384 = ~n24383 & ~n24382;
  assign n24386 = ~n24385 | ~n24384;
  assign n24388 = ~P3_INSTQUEUE_REG_7__6__SCAN_IN;
  assign n24390 = ~n22844 & ~n24388;
  assign n34783 = ~P3_INSTQUEUE_REG_3__6__SCAN_IN;
  assign n24389 = ~n34610 & ~n34783;
  assign n24392 = ~n24390 & ~n24389;
  assign n24391 = ~n34872 | ~P3_INSTQUEUE_REG_14__6__SCAN_IN;
  assign n24394 = ~n24392 | ~n24391;
  assign n34778 = ~P3_INSTQUEUE_REG_6__6__SCAN_IN;
  assign n24393 = ~n24522 & ~n34778;
  assign n24402 = ~n24394 & ~n24393;
  assign n24396 = ~n35319 | ~P3_INSTQUEUE_REG_8__6__SCAN_IN;
  assign n24395 = ~n34564 | ~P3_INSTQUEUE_REG_15__6__SCAN_IN;
  assign n24400 = ~n24396 | ~n24395;
  assign n24398 = ~n34575 | ~P3_INSTQUEUE_REG_0__6__SCAN_IN;
  assign n24397 = ~n24516 | ~P3_INSTQUEUE_REG_12__6__SCAN_IN;
  assign n24399 = ~n24398 | ~n24397;
  assign n24401 = ~n24400 & ~n24399;
  assign n24418 = ~n24402 | ~n24401;
  assign n24404 = ~n34545 | ~P3_INSTQUEUE_REG_5__6__SCAN_IN;
  assign n24403 = ~n34717 | ~P3_INSTQUEUE_REG_11__6__SCAN_IN;
  assign n24408 = ~n24404 | ~n24403;
  assign n24406 = ~n35252 | ~P3_INSTQUEUE_REG_13__6__SCAN_IN;
  assign n24405 = ~n24543 | ~P3_INSTQUEUE_REG_4__6__SCAN_IN;
  assign n24407 = ~n24406 | ~n24405;
  assign n24416 = ~n24408 & ~n24407;
  assign n24410 = ~n24451 | ~P3_INSTQUEUE_REG_9__6__SCAN_IN;
  assign n24409 = ~n24513 | ~P3_INSTQUEUE_REG_10__6__SCAN_IN;
  assign n24414 = ~n24410 | ~n24409;
  assign n24412 = ~n35328 | ~P3_INSTQUEUE_REG_1__6__SCAN_IN;
  assign n24411 = ~n24470 | ~P3_INSTQUEUE_REG_2__6__SCAN_IN;
  assign n24413 = ~n24412 | ~n24411;
  assign n24415 = ~n24414 & ~n24413;
  assign n24417 = ~n24416 | ~n24415;
  assign n24616 = ~n24721;
  assign n24420 = ~n35412 | ~P3_INSTQUEUE_REG_6__3__SCAN_IN;
  assign n24419 = ~n34872 | ~P3_INSTQUEUE_REG_14__3__SCAN_IN;
  assign n24424 = ~n24420 | ~n24419;
  assign n24422 = ~n24451 | ~P3_INSTQUEUE_REG_9__3__SCAN_IN;
  assign n24421 = ~n35252 | ~P3_INSTQUEUE_REG_13__3__SCAN_IN;
  assign n24423 = ~n24422 | ~n24421;
  assign n24432 = ~n24424 & ~n24423;
  assign n24426 = ~n34717 | ~P3_INSTQUEUE_REG_11__3__SCAN_IN;
  assign n24425 = ~n24543 | ~P3_INSTQUEUE_REG_4__3__SCAN_IN;
  assign n24430 = ~n24426 | ~n24425;
  assign n24428 = ~n24513 | ~P3_INSTQUEUE_REG_10__3__SCAN_IN;
  assign n24427 = ~n35319 | ~P3_INSTQUEUE_REG_8__3__SCAN_IN;
  assign n24429 = ~n24428 | ~n24427;
  assign n24431 = ~n24430 & ~n24429;
  assign n24448 = ~n24432 | ~n24431;
  assign n24434 = ~n34575 | ~P3_INSTQUEUE_REG_0__3__SCAN_IN;
  assign n24433 = ~n24470 | ~P3_INSTQUEUE_REG_2__3__SCAN_IN;
  assign n24438 = ~n24434 | ~n24433;
  assign n24436 = ~n24535 | ~P3_INSTQUEUE_REG_5__3__SCAN_IN;
  assign n24435 = ~n35328 | ~P3_INSTQUEUE_REG_1__3__SCAN_IN;
  assign n24437 = ~n24436 | ~n24435;
  assign n24446 = ~n24438 & ~n24437;
  assign n24440 = ~n24540 | ~P3_INSTQUEUE_REG_7__3__SCAN_IN;
  assign n24439 = ~n34564 | ~P3_INSTQUEUE_REG_15__3__SCAN_IN;
  assign n24444 = ~n24440 | ~n24439;
  assign n24442 = ~n34993 | ~P3_INSTQUEUE_REG_3__3__SCAN_IN;
  assign n24441 = ~n24516 | ~P3_INSTQUEUE_REG_12__3__SCAN_IN;
  assign n24443 = ~n24442 | ~n24441;
  assign n24445 = ~n24444 & ~n24443;
  assign n24447 = ~n24446 | ~n24445;
  assign n24450 = ~n34717 | ~P3_INSTQUEUE_REG_11__7__SCAN_IN;
  assign n24449 = ~n24540 | ~P3_INSTQUEUE_REG_7__7__SCAN_IN;
  assign n24455 = ~n24450 | ~n24449;
  assign n24453 = ~n24451 | ~P3_INSTQUEUE_REG_9__7__SCAN_IN;
  assign n24452 = ~n35252 | ~P3_INSTQUEUE_REG_13__7__SCAN_IN;
  assign n24454 = ~n24453 | ~n24452;
  assign n24463 = ~n24455 & ~n24454;
  assign n24457 = ~n24535 | ~P3_INSTQUEUE_REG_5__7__SCAN_IN;
  assign n24456 = ~n35328 | ~P3_INSTQUEUE_REG_1__7__SCAN_IN;
  assign n24461 = ~n24457 | ~n24456;
  assign n24459 = ~n35412 | ~P3_INSTQUEUE_REG_6__7__SCAN_IN;
  assign n24458 = ~n34872 | ~P3_INSTQUEUE_REG_14__7__SCAN_IN;
  assign n24460 = ~n24459 | ~n24458;
  assign n24462 = ~n24461 & ~n24460;
  assign n24480 = ~n24463 | ~n24462;
  assign n24465 = ~n24513 | ~P3_INSTQUEUE_REG_10__7__SCAN_IN;
  assign n24464 = ~n24543 | ~P3_INSTQUEUE_REG_4__7__SCAN_IN;
  assign n24469 = ~n24465 | ~n24464;
  assign n24467 = ~n34575 | ~P3_INSTQUEUE_REG_0__7__SCAN_IN;
  assign n24466 = ~n24516 | ~P3_INSTQUEUE_REG_12__7__SCAN_IN;
  assign n24468 = ~n24467 | ~n24466;
  assign n24478 = ~n24469 & ~n24468;
  assign n24472 = ~n24470 | ~P3_INSTQUEUE_REG_2__7__SCAN_IN;
  assign n24471 = ~n34564 | ~P3_INSTQUEUE_REG_15__7__SCAN_IN;
  assign n24476 = ~n24472 | ~n24471;
  assign n24474 = ~n35319 | ~P3_INSTQUEUE_REG_8__7__SCAN_IN;
  assign n24473 = ~n34993 | ~P3_INSTQUEUE_REG_3__7__SCAN_IN;
  assign n24475 = ~n24474 | ~n24473;
  assign n24477 = ~n24476 & ~n24475;
  assign n24479 = ~n24478 | ~n24477;
  assign n24481 = ~n24616 | ~n24668;
  assign n24484 = ~n35412 | ~P3_INSTQUEUE_REG_6__1__SCAN_IN;
  assign n24483 = ~n35319 | ~P3_INSTQUEUE_REG_8__1__SCAN_IN;
  assign n24488 = ~n24484 | ~n24483;
  assign n24486 = ~n34872 | ~P3_INSTQUEUE_REG_14__1__SCAN_IN;
  assign n24485 = ~n24516 | ~P3_INSTQUEUE_REG_12__1__SCAN_IN;
  assign n24487 = ~n24486 | ~n24485;
  assign n24496 = ~n24488 & ~n24487;
  assign n24490 = ~n24513 | ~P3_INSTQUEUE_REG_10__1__SCAN_IN;
  assign n24489 = ~n24543 | ~P3_INSTQUEUE_REG_4__1__SCAN_IN;
  assign n24494 = ~n24490 | ~n24489;
  assign n24492 = ~n35252 | ~P3_INSTQUEUE_REG_13__1__SCAN_IN;
  assign n24491 = ~n34564 | ~P3_INSTQUEUE_REG_15__1__SCAN_IN;
  assign n24493 = ~n24492 | ~n24491;
  assign n24495 = ~n24494 & ~n24493;
  assign n24512 = ~n24496 | ~n24495;
  assign n24498 = ~n35328 | ~P3_INSTQUEUE_REG_1__1__SCAN_IN;
  assign n24497 = ~n34993 | ~P3_INSTQUEUE_REG_3__1__SCAN_IN;
  assign n24502 = ~n24498 | ~n24497;
  assign n24500 = ~n34717 | ~P3_INSTQUEUE_REG_11__1__SCAN_IN;
  assign n24499 = ~n24540 | ~P3_INSTQUEUE_REG_7__1__SCAN_IN;
  assign n24501 = ~n24500 | ~n24499;
  assign n24510 = ~n24502 & ~n24501;
  assign n24504 = ~n24451 | ~P3_INSTQUEUE_REG_9__1__SCAN_IN;
  assign n24503 = ~n35405 | ~P3_INSTQUEUE_REG_0__1__SCAN_IN;
  assign n24508 = ~n24504 | ~n24503;
  assign n24506 = ~n34545 | ~P3_INSTQUEUE_REG_5__1__SCAN_IN;
  assign n24505 = ~n24470 | ~P3_INSTQUEUE_REG_2__1__SCAN_IN;
  assign n24507 = ~n24506 | ~n24505;
  assign n24509 = ~n24508 & ~n24507;
  assign n24511 = ~n24510 | ~n24509;
  assign n24515 = ~n34564 | ~P3_INSTQUEUE_REG_15__0__SCAN_IN;
  assign n24514 = ~n24513 | ~P3_INSTQUEUE_REG_10__0__SCAN_IN;
  assign n24520 = ~n24515 | ~n24514;
  assign n24518 = ~n34872 | ~P3_INSTQUEUE_REG_14__0__SCAN_IN;
  assign n24517 = ~n24516 | ~P3_INSTQUEUE_REG_12__0__SCAN_IN;
  assign n24519 = ~n24518 | ~n24517;
  assign n24532 = ~n24520 & ~n24519;
  assign n24521 = ~P3_INSTQUEUE_REG_6__0__SCAN_IN;
  assign n24530 = ~n24522 & ~n24521;
  assign n24523 = ~P3_INSTQUEUE_REG_9__0__SCAN_IN;
  assign n24526 = ~n34631 & ~n24523;
  assign n24524 = ~P3_INSTQUEUE_REG_2__0__SCAN_IN;
  assign n24525 = ~n34779 & ~n24524;
  assign n24528 = ~n24526 & ~n24525;
  assign n24527 = ~n35252 | ~P3_INSTQUEUE_REG_13__0__SCAN_IN;
  assign n24529 = ~n24528 | ~n24527;
  assign n24531 = ~n24530 & ~n24529;
  assign n24551 = ~n24532 | ~n24531;
  assign n24534 = ~n35328 | ~P3_INSTQUEUE_REG_1__0__SCAN_IN;
  assign n24533 = ~n34993 | ~P3_INSTQUEUE_REG_3__0__SCAN_IN;
  assign n24539 = ~n24534 | ~n24533;
  assign n24537 = ~n24535 | ~P3_INSTQUEUE_REG_5__0__SCAN_IN;
  assign n24536 = ~n34717 | ~P3_INSTQUEUE_REG_11__0__SCAN_IN;
  assign n24538 = ~n24537 | ~n24536;
  assign n24549 = ~n24539 & ~n24538;
  assign n24542 = ~n35319 | ~P3_INSTQUEUE_REG_8__0__SCAN_IN;
  assign n24541 = ~n24540 | ~P3_INSTQUEUE_REG_7__0__SCAN_IN;
  assign n24547 = ~n24542 | ~n24541;
  assign n24545 = ~n34575 | ~P3_INSTQUEUE_REG_0__0__SCAN_IN;
  assign n24544 = ~n24543 | ~P3_INSTQUEUE_REG_4__0__SCAN_IN;
  assign n24546 = ~n24545 | ~n24544;
  assign n24548 = ~n24547 & ~n24546;
  assign n24550 = ~n24549 | ~n24548;
  assign n33406 = ~n38678 | ~n33284;
  assign n24631 = ~P3_INSTADDRPOINTER_REG_27__SCAN_IN | ~P3_INSTADDRPOINTER_REG_28__SCAN_IN;
  assign n24646 = ~n24631;
  assign n36380 = ~P3_INSTADDRPOINTER_REG_16__SCAN_IN | ~P3_INSTADDRPOINTER_REG_17__SCAN_IN;
  assign n36258 = ~n36380 & ~n36874;
  assign n33412 = ~n36258;
  assign n37059 = ~P3_INSTADDRPOINTER_REG_12__SCAN_IN | ~n37065;
  assign n37056 = ~n37066 & ~n37059;
  assign n35794 = ~n24552;
  assign n24553 = ~n27595 | ~n24569;
  assign n24565 = ~n35794 | ~n24553;
  assign n24559 = ~n24565 | ~n35782;
  assign n24557 = ~n24559 & ~n35773;
  assign n24554 = ~n24557;
  assign n24556 = ~n24554 & ~n35761;
  assign n24555 = ~n24556 | ~n35753;
  assign n24586 = ~n37212 & ~n24555;
  assign n24587 = ~n33284 ^ n24555;
  assign n24583 = n35753 ^ n24556;
  assign n24558 = ~n24557 ^ n35761;
  assign n24581 = ~P3_INSTADDRPOINTER_REG_5__SCAN_IN | ~n24558;
  assign n36678 = P3_INSTADDRPOINTER_REG_5__SCAN_IN ^ n24558;
  assign n24561 = ~n24559 ^ n35773;
  assign n24560 = ~n24561;
  assign n24580 = ~n24560 | ~P3_INSTADDRPOINTER_REG_4__SCAN_IN;
  assign n36690 = ~n24561 ^ P3_INSTADDRPOINTER_REG_4__SCAN_IN;
  assign n24563 = ~n24565 ^ n35782;
  assign n24562 = ~n24563;
  assign n24578 = ~n24562 | ~P3_INSTADDRPOINTER_REG_3__SCAN_IN;
  assign n36705 = ~n24563 ^ P3_INSTADDRPOINTER_REG_3__SCAN_IN;
  assign n24566 = ~n24564 | ~n27595;
  assign n24568 = ~n24566 | ~n24565;
  assign n24576 = ~n24568 | ~P3_INSTADDRPOINTER_REG_2__SCAN_IN;
  assign n36716 = ~n24568 ^ n24567;
  assign n24570 = ~n27595;
  assign n24571 = ~n24570 | ~n24569;
  assign n24573 = ~n24572 | ~n24571;
  assign n36715 = n24574 & n24573;
  assign n24575 = ~n36716 | ~n36715;
  assign n36677 = ~n24580 | ~n24579;
  assign n24584 = ~n24583 | ~n24582;
  assign n24592 = ~n24586 | ~n24585;
  assign n24590 = ~n24586 ^ n24585;
  assign n36645 = n24588 & n24587;
  assign n24589 = ~n36645;
  assign n36619 = ~n24590 | ~n24589;
  assign n24591 = ~P3_INSTADDRPOINTER_REG_8__SCAN_IN | ~n36619;
  assign n36462 = n37056 & n37185;
  assign n36201 = ~P3_INSTADDRPOINTER_REG_24__SCAN_IN | ~n36833;
  assign n24597 = ~n33338 & ~n38674;
  assign n37087 = ~n37121;
  assign n37085 = ~P3_INSTADDRPOINTER_REG_11__SCAN_IN | ~P3_INSTADDRPOINTER_REG_12__SCAN_IN;
  assign n24628 = ~n24595;
  assign n37184 = ~n37212 | ~n38678;
  assign n33393 = ~n33307 & ~n37184;
  assign n24649 = ~P3_INSTADDRPOINTER_REG_30__SCAN_IN | ~n33388;
  assign n24605 = ~n35948 | ~n39110;
  assign n24667 = ~n24605;
  assign n24599 = ~n37473 | ~n37514;
  assign n24665 = ~n39110 | ~n37482;
  assign n38745 = ~n24599 & ~n24598;
  assign n24678 = ~n37463 & ~n38745;
  assign n33740 = ~n37463;
  assign n24601 = ~n24668 | ~n24600;
  assign n24602 = ~n39110 & ~n24601;
  assign n24603 = ~n33740 & ~n24602;
  assign n35943 = ~n34481 | ~n24604;
  assign n24606 = ~n37473 | ~n24605;
  assign n27588 = ~n37453 | ~n39110;
  assign n24623 = ~n34971 & ~n27588;
  assign n24614 = ~n24606 & ~n24623;
  assign n38756 = ~n24634 & ~n24625;
  assign n24664 = ~n37482 | ~n38756;
  assign n24607 = ~n37463 | ~n39110;
  assign n24611 = ~n24608 & ~n24607;
  assign n24609 = ~n34971 & ~n24616;
  assign n24610 = ~n37482 & ~n24609;
  assign n24612 = ~n24611 & ~n24610;
  assign n24613 = ~n24664 | ~n24612;
  assign n24622 = ~n24614 & ~n24613;
  assign n24615 = ~n24667 & ~n33740;
  assign n24620 = ~n24616 & ~n24615;
  assign n27590 = n34971 | n38756;
  assign n24675 = ~n24632 | ~n27590;
  assign n24618 = n24675 & n24617;
  assign n24619 = ~n37473 & ~n24618;
  assign n24621 = ~n24620 & ~n24619;
  assign n38732 = ~n24622 | ~n24621;
  assign n24626 = ~n24623;
  assign n24642 = ~n37463 | ~n37473;
  assign n24624 = ~n37502 & ~n24642;
  assign n27586 = ~n24625 | ~n24624;
  assign n24627 = ~n24626 & ~n27586;
  assign n38703 = ~n38732 & ~n38710;
  assign n27583 = ~n35943 | ~n38763;
  assign n36962 = ~P3_INSTADDRPOINTER_REG_19__SCAN_IN;
  assign n37295 = ~P3_INSTADDRPOINTER_REG_2__SCAN_IN | ~P3_INSTADDRPOINTER_REG_1__SCAN_IN;
  assign n37302 = ~P3_INSTADDRPOINTER_REG_4__SCAN_IN;
  assign n37317 = ~P3_INSTADDRPOINTER_REG_3__SCAN_IN;
  assign n37278 = ~n37302 & ~n37317;
  assign n37256 = ~P3_INSTADDRPOINTER_REG_5__SCAN_IN | ~n37278;
  assign n37259 = ~n37295 & ~n37256;
  assign n37188 = ~P3_INSTADDRPOINTER_REG_6__SCAN_IN | ~n37259;
  assign n37058 = ~n37210 & ~n37235;
  assign n24638 = ~n37058;
  assign n37140 = ~n37188 & ~n24638;
  assign n37062 = ~n37056 | ~n37140;
  assign n36968 = ~n24628 & ~n37062;
  assign n36863 = ~n36380 & ~n36327;
  assign n36916 = ~n36968 | ~n36863;
  assign n36884 = ~n36962 & ~n36916;
  assign n33413 = n24629 & n36884;
  assign n36869 = ~P3_INSTADDRPOINTER_REG_23__SCAN_IN;
  assign n36849 = ~P3_INSTADDRPOINTER_REG_24__SCAN_IN;
  assign n36811 = ~n36869 & ~n36849;
  assign n24630 = ~P3_INSTADDRPOINTER_REG_22__SCAN_IN | ~n36811;
  assign n33417 = ~n24630 & ~n36781;
  assign n33433 = ~n33413 | ~n33417;
  assign n24652 = ~n24631 & ~n33433;
  assign n33386 = ~n22828 & ~n24652;
  assign n39129 = ~n24632 & ~n24667;
  assign n24636 = ~n39129;
  assign n24635 = ~n24633;
  assign n38706 = ~n24634 & ~n37482;
  assign n27584 = ~n24635 | ~n38706;
  assign n38730 = ~n24636 & ~n27584;
  assign n36774 = ~n36811;
  assign n37369 = ~P3_INSTADDRPOINTER_REG_1__SCAN_IN;
  assign n24637 = ~n37369 & ~n37382;
  assign n37294 = ~P3_INSTADDRPOINTER_REG_2__SCAN_IN & ~n24637;
  assign n37260 = ~n37294 & ~n37256;
  assign n37218 = ~P3_INSTADDRPOINTER_REG_6__SCAN_IN | ~n37260;
  assign n37064 = ~n24638 & ~n37218;
  assign n36990 = P3_INSTADDRPOINTER_REG_14__SCAN_IN & n37056;
  assign n37012 = ~n37064 | ~n36990;
  assign n24639 = ~n36380 & ~n37012;
  assign n36975 = ~P3_INSTADDRPOINTER_REG_15__SCAN_IN | ~n24639;
  assign n36919 = ~n36327 & ~n36975;
  assign n36893 = ~P3_INSTADDRPOINTER_REG_21__SCAN_IN;
  assign n36951 = ~P3_INSTADDRPOINTER_REG_20__SCAN_IN;
  assign n36909 = ~n36962 & ~n36951;
  assign n24640 = ~P3_INSTADDRPOINTER_REG_22__SCAN_IN | ~n36909;
  assign n36864 = ~n36893 & ~n24640;
  assign n36842 = ~n36919 | ~n36864;
  assign n36792 = ~n36774 & ~n36842;
  assign n24654 = n36792 & n24641;
  assign n33382 = n38673 | n24654;
  assign n38744 = ~n38703;
  assign n38704 = ~n37453 & ~n24668;
  assign n38705 = ~n24642;
  assign n24643 = ~n38704 & ~n38705;
  assign n24644 = ~n38744 & ~n24643;
  assign n37010 = ~P3_INSTADDRPOINTER_REG_0__SCAN_IN | ~n36968;
  assign n36879 = ~n33412 & ~n37010;
  assign n36836 = ~P3_INSTADDRPOINTER_REG_22__SCAN_IN | ~n36879;
  assign n36770 = ~n36774 & ~n36836;
  assign n24645 = ~n36781 & ~n36764;
  assign n24653 = ~n36770 | ~n24645;
  assign n33384 = ~n38757 | ~n24653;
  assign n33432 = ~n33382 | ~n33384;
  assign n24648 = ~n33386 & ~n33432;
  assign n33313 = ~n24646 | ~P3_INSTADDRPOINTER_REG_29__SCAN_IN;
  assign n36932 = ~n38757 & ~n38730;
  assign n37356 = ~n22828 | ~n36932;
  assign n24647 = ~n33313 | ~n37356;
  assign n33365 = ~n24648 | ~n24647;
  assign n24663 = ~n24649 & ~n33365;
  assign n24651 = ~n37292 | ~n33338;
  assign n24650 = ~n33307 | ~n37147;
  assign n24661 = ~n24651 | ~n24650;
  assign n24659 = ~n24652 | ~n38758;
  assign n24656 = n22834 | n24653;
  assign n24655 = n24654 & P3_INSTADDRPOINTER_REG_27__SCAN_IN;
  assign n33419 = ~n38730 | ~n24655;
  assign n24657 = ~n24656 | ~n33419;
  assign n24658 = ~n24657 | ~P3_INSTADDRPOINTER_REG_28__SCAN_IN;
  assign n33395 = ~n24659 | ~n24658;
  assign n33362 = ~P3_INSTADDRPOINTER_REG_29__SCAN_IN | ~n33395;
  assign n24660 = ~n33362 | ~n24287;
  assign n24662 = ~n24661 & ~n24660;
  assign n24671 = ~n24665 | ~n24664;
  assign n24666 = ~n37482 & ~n37502;
  assign n24669 = ~n24667 & ~n24666;
  assign n24670 = ~n24669 | ~n24668;
  assign n24672 = ~n24671 & ~n24670;
  assign n24674 = ~n24673 | ~n24672;
  assign n24676 = ~n24674 | ~n37463;
  assign n24677 = ~n24676 | ~n24675;
  assign n38692 = ~n24678 & ~n24677;
  assign n24716 = ~n23759 ^ n38768;
  assign n24679 = ~n38695 & ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n24692 = ~n24716 ^ n24679;
  assign n24690 = ~P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN | ~n38686;
  assign n24693 = ~P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN & ~n38686;
  assign n37428 = ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign n24685 = ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~n37428;
  assign n24680 = ~n38768 | ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN;
  assign n24682 = ~n38723 | ~n24680;
  assign n24684 = ~n24682 | ~n24681;
  assign n24683 = ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN | ~n38768;
  assign n24699 = ~n24684 | ~n24683;
  assign n24698 = ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN ^ P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign n24701 = ~n24699 | ~n24698;
  assign n24687 = ~n24685 | ~n24701;
  assign n24686 = ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN & ~n24687;
  assign n24697 = ~n24693 & ~n24686;
  assign n24694 = ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~n24687;
  assign n24688 = ~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | ~n24694;
  assign n24689 = ~n24697 | ~n24688;
  assign n24691 = ~n24704;
  assign n24705 = ~n24692 | ~n24691;
  assign n24695 = n24694 & n24693;
  assign n24696 = ~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & ~n24695;
  assign n24718 = ~n24697 & ~n24696;
  assign n24700 = n24699 | n24698;
  assign n24702 = ~n24701 | ~n24700;
  assign n24703 = ~n24718 & ~n24702;
  assign n33737 = ~P3_STATE_REG_1__SCAN_IN & ~P3_STATE_REG_2__SCAN_IN;
  assign n24706 = ~P3_STATE_REG_0__SCAN_IN & ~n33737;
  assign n39005 = ~n39126 | ~P3_STATE_REG_2__SCAN_IN;
  assign n39112 = ~n24706 | ~n39005;
  assign n24707 = ~n37453 & ~n35811;
  assign n33742 = ~n37463 & ~n24707;
  assign n24708 = ~n39112 & ~n37494;
  assign n24709 = ~n33742 & ~n24708;
  assign n24726 = ~n38688 & ~n24709;
  assign n24713 = ~n37494 & ~n38688;
  assign n24715 = ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN ^ P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n24711 = ~n24710 | ~n24715;
  assign n38677 = ~n38681 | ~n24711;
  assign n24712 = ~n37502 & ~n38677;
  assign n24714 = ~n24713 & ~n24712;
  assign n24723 = ~n37453 & ~n24714;
  assign n24717 = ~n24716 | ~n24715;
  assign n24719 = n24718 | n24717;
  assign n24722 = ~n24721 & ~n38675;
  assign n24724 = ~n24723 & ~n24722;
  assign n24725 = ~n24724 & ~n33740;
  assign n24727 = ~n24726 & ~n24725;
  assign n24729 = ~n38692 | ~n24727;
  assign n24728 = ~n38675 & ~n37482;
  assign n39056 = ~n39069 | ~n38487;
  assign n38803 = ~P3_STATE2_REG_2__SCAN_IN;
  assign n38810 = ~n38803 | ~n39118;
  assign n24732 = ~n37352 | ~P3_INSTADDRPOINTER_REG_30__SCAN_IN;
  assign n33319 = ~n22843 | ~P3_REIP_REG_30__SCAN_IN;
  assign P3_U2832 = ~n24733 | ~n23968;
  assign n25574 = ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n24741 = ~n22832 & ~n24735;
  assign n24737 = ~n24911 | ~P1_INSTQUEUE_REG_13__0__SCAN_IN;
  assign n24736 = ~n25196 | ~P1_INSTQUEUE_REG_0__0__SCAN_IN;
  assign n24740 = ~n22970 | ~n23959;
  assign n24749 = ~n24741 & ~n24740;
  assign n24743 = ~n26851 | ~P1_INSTQUEUE_REG_7__0__SCAN_IN;
  assign n24742 = ~n26630 | ~P1_INSTQUEUE_REG_8__0__SCAN_IN;
  assign n24747 = ~n24743 | ~n24742;
  assign n26629 = n31445 & n24753;
  assign n24745 = ~n26629 | ~P1_INSTQUEUE_REG_10__0__SCAN_IN;
  assign n24744 = ~n24976 | ~P1_INSTQUEUE_REG_14__0__SCAN_IN;
  assign n24746 = ~n24745 | ~n24744;
  assign n24769 = ~n24749 | ~n24748;
  assign n24905 = ~n31536 | ~n31445;
  assign n24750 = ~P1_INSTQUEUE_REG_11__0__SCAN_IN;
  assign n24751 = ~n25085 | ~P1_INSTQUEUE_REG_3__0__SCAN_IN;
  assign n24758 = ~n24752 | ~n24751;
  assign n25088 = n24753 & n31461;
  assign n24756 = ~n25088 | ~P1_INSTQUEUE_REG_2__0__SCAN_IN;
  assign n24755 = ~n25089 | ~P1_INSTQUEUE_REG_12__0__SCAN_IN;
  assign n24757 = ~n24756 | ~n24755;
  assign n24947 = n24763 & n31445;
  assign n24761 = ~n24947 | ~P1_INSTQUEUE_REG_9__0__SCAN_IN;
  assign n24760 = ~n22826 | ~P1_INSTQUEUE_REG_15__0__SCAN_IN;
  assign n24767 = ~n24898 | ~P1_INSTQUEUE_REG_1__0__SCAN_IN;
  assign n24766 = ~n25118 | ~P1_INSTQUEUE_REG_4__0__SCAN_IN;
  assign n24768 = ~n22967 | ~n23961;
  assign n24771 = ~n25100 | ~P1_INSTQUEUE_REG_13__3__SCAN_IN;
  assign n24770 = ~n25196 | ~P1_INSTQUEUE_REG_0__3__SCAN_IN;
  assign n24774 = ~n24771 | ~n24770;
  assign n24772 = ~P1_INSTQUEUE_REG_5__3__SCAN_IN;
  assign n24773 = ~n25065 & ~n24772;
  assign n24777 = ~n24774 & ~n24773;
  assign n24775 = ~P1_INSTQUEUE_REG_6__3__SCAN_IN;
  assign n24785 = ~n24777 | ~n24776;
  assign n24779 = ~n24972 | ~P1_INSTQUEUE_REG_7__3__SCAN_IN;
  assign n24778 = ~n24973 | ~P1_INSTQUEUE_REG_8__3__SCAN_IN;
  assign n24781 = ~n26629 | ~P1_INSTQUEUE_REG_10__3__SCAN_IN;
  assign n24780 = ~n24976 | ~P1_INSTQUEUE_REG_14__3__SCAN_IN;
  assign n24782 = n24781 & n24780;
  assign n24784 = ~n24783 | ~n24782;
  assign n24786 = ~P1_INSTQUEUE_REG_11__3__SCAN_IN;
  assign n24788 = n24905 | n24786;
  assign n24787 = ~n22829 | ~P1_INSTQUEUE_REG_3__3__SCAN_IN;
  assign n24792 = ~n24788 | ~n24787;
  assign n24790 = ~n25088 | ~P1_INSTQUEUE_REG_2__3__SCAN_IN;
  assign n24789 = ~n25089 | ~P1_INSTQUEUE_REG_12__3__SCAN_IN;
  assign n24791 = ~n24790 | ~n24789;
  assign n24800 = ~n24792 & ~n24791;
  assign n24794 = ~n24898 | ~P1_INSTQUEUE_REG_1__3__SCAN_IN;
  assign n24793 = ~n25118 | ~P1_INSTQUEUE_REG_4__3__SCAN_IN;
  assign n24798 = ~n24794 | ~n24793;
  assign n24796 = ~n24947 | ~P1_INSTQUEUE_REG_9__3__SCAN_IN;
  assign n24795 = ~n22826 | ~P1_INSTQUEUE_REG_15__3__SCAN_IN;
  assign n24797 = ~n24796 | ~n24795;
  assign n24799 = ~n24798 & ~n24797;
  assign n24803 = ~n24947;
  assign n24804 = ~n24898 | ~P1_INSTQUEUE_REG_1__6__SCAN_IN;
  assign n25123 = ~n24905;
  assign n24806 = ~n25123 | ~P1_INSTQUEUE_REG_11__6__SCAN_IN;
  assign n24805 = ~n25088 | ~P1_INSTQUEUE_REG_2__6__SCAN_IN;
  assign n24808 = ~n22862 | ~P1_INSTQUEUE_REG_5__6__SCAN_IN;
  assign n24807 = ~n24976 | ~P1_INSTQUEUE_REG_14__6__SCAN_IN;
  assign n24812 = ~n24808 | ~n24807;
  assign n26851 = n24936;
  assign n24810 = ~n26851 | ~P1_INSTQUEUE_REG_7__6__SCAN_IN;
  assign n24809 = ~n22826 | ~P1_INSTQUEUE_REG_15__6__SCAN_IN;
  assign n24811 = ~n24810 | ~n24809;
  assign n24833 = ~n24814 | ~n24813;
  assign n25100 = ~n26482;
  assign n24817 = ~n25100 | ~P1_INSTQUEUE_REG_13__6__SCAN_IN;
  assign n24816 = ~n24973 | ~P1_INSTQUEUE_REG_8__6__SCAN_IN;
  assign n24821 = ~n24817 | ~n24816;
  assign n24819 = ~n26629 | ~P1_INSTQUEUE_REG_10__6__SCAN_IN;
  assign n24818 = ~n25118 | ~P1_INSTQUEUE_REG_4__6__SCAN_IN;
  assign n24820 = ~n24819 | ~n24818;
  assign n24831 = ~n24821 & ~n24820;
  assign n24822 = ~P1_INSTQUEUE_REG_6__6__SCAN_IN;
  assign n24824 = ~n25196 | ~P1_INSTQUEUE_REG_0__6__SCAN_IN;
  assign n24823 = ~n25085 | ~P1_INSTQUEUE_REG_3__6__SCAN_IN;
  assign n24828 = ~n24823 | ~n24824;
  assign n24826 = ~n25089;
  assign n24825 = ~P1_INSTQUEUE_REG_12__6__SCAN_IN;
  assign n24827 = ~n24826 & ~n24825;
  assign n24829 = ~n24828 & ~n24827;
  assign n24835 = ~n24947 | ~P1_INSTQUEUE_REG_9__7__SCAN_IN;
  assign n24834 = ~n24898 | ~P1_INSTQUEUE_REG_1__7__SCAN_IN;
  assign n24839 = ~n24835 | ~n24834;
  assign n24837 = ~n24989 | ~P1_INSTQUEUE_REG_11__7__SCAN_IN;
  assign n24836 = ~n25089 | ~P1_INSTQUEUE_REG_12__7__SCAN_IN;
  assign n24838 = ~n24837 | ~n24836;
  assign n24847 = ~n24839 & ~n24838;
  assign n24841 = ~n22862 | ~P1_INSTQUEUE_REG_5__7__SCAN_IN;
  assign n24840 = ~n26629 | ~P1_INSTQUEUE_REG_10__7__SCAN_IN;
  assign n24845 = ~n24841 | ~n24840;
  assign n24843 = ~n25088 | ~P1_INSTQUEUE_REG_2__7__SCAN_IN;
  assign n24842 = ~n25196 | ~P1_INSTQUEUE_REG_0__7__SCAN_IN;
  assign n24844 = ~n24843 | ~n24842;
  assign n24846 = ~n24845 & ~n24844;
  assign n24863 = ~n24847 | ~n24846;
  assign n24853 = ~n22832 & ~n25103;
  assign n24911 = ~n26482;
  assign n24849 = ~n24911 | ~P1_INSTQUEUE_REG_13__7__SCAN_IN;
  assign n24848 = ~n22829 | ~P1_INSTQUEUE_REG_3__7__SCAN_IN;
  assign n24850 = ~n26851 | ~P1_INSTQUEUE_REG_7__7__SCAN_IN;
  assign n24852 = ~n24851 | ~n24850;
  assign n24855 = ~n26630 | ~P1_INSTQUEUE_REG_8__7__SCAN_IN;
  assign n24854 = ~n24976 | ~P1_INSTQUEUE_REG_14__7__SCAN_IN;
  assign n24859 = ~n24855 | ~n24854;
  assign n24857 = ~n25118 | ~P1_INSTQUEUE_REG_4__7__SCAN_IN;
  assign n24856 = ~n22826 | ~P1_INSTQUEUE_REG_15__7__SCAN_IN;
  assign n24858 = ~n24857 | ~n24856;
  assign n24860 = ~n24859 & ~n24858;
  assign n24862 = ~n24861 | ~n24860;
  assign n25002 = ~n25685 | ~n25022;
  assign n24864 = ~n25002;
  assign n24929 = ~n24865 | ~n24864;
  assign n24867 = ~n24898 | ~P1_INSTQUEUE_REG_1__4__SCAN_IN;
  assign n24866 = ~n25118 | ~P1_INSTQUEUE_REG_4__4__SCAN_IN;
  assign n24871 = ~n24867 | ~n24866;
  assign n24868 = ~n22826 | ~P1_INSTQUEUE_REG_15__4__SCAN_IN;
  assign n24870 = ~n24869 | ~n24868;
  assign n24879 = ~n24871 & ~n24870;
  assign n24873 = ~n24989 | ~P1_INSTQUEUE_REG_11__4__SCAN_IN;
  assign n24872 = ~n22829 | ~P1_INSTQUEUE_REG_3__4__SCAN_IN;
  assign n24877 = ~n24873 | ~n24872;
  assign n24875 = ~n25088 | ~P1_INSTQUEUE_REG_2__4__SCAN_IN;
  assign n24874 = ~n25089 | ~P1_INSTQUEUE_REG_12__4__SCAN_IN;
  assign n24876 = ~n24875 | ~n24874;
  assign n24881 = ~n25100 | ~P1_INSTQUEUE_REG_13__4__SCAN_IN;
  assign n24880 = ~n25196 | ~P1_INSTQUEUE_REG_0__4__SCAN_IN;
  assign n24884 = ~n24881 | ~n24880;
  assign n24883 = ~n25065 & ~n24882;
  assign n24887 = ~n24884 & ~n24883;
  assign n24895 = ~n24887 | ~n24886;
  assign n24889 = ~n24972 | ~P1_INSTQUEUE_REG_7__4__SCAN_IN;
  assign n24888 = ~n24973 | ~P1_INSTQUEUE_REG_8__4__SCAN_IN;
  assign n24891 = ~n26629 | ~P1_INSTQUEUE_REG_10__4__SCAN_IN;
  assign n24890 = ~n24976 | ~P1_INSTQUEUE_REG_14__4__SCAN_IN;
  assign n24894 = ~n24893 | ~n24892;
  assign n24900 = ~n24898 | ~P1_INSTQUEUE_REG_1__5__SCAN_IN;
  assign n24899 = ~n25118 | ~P1_INSTQUEUE_REG_4__5__SCAN_IN;
  assign n24904 = ~n24900 | ~n24899;
  assign n24902 = ~n24947 | ~P1_INSTQUEUE_REG_9__5__SCAN_IN;
  assign n24901 = ~n22826 | ~P1_INSTQUEUE_REG_15__5__SCAN_IN;
  assign n24903 = ~n24902 | ~n24901;
  assign n24910 = ~n24904 & ~n24903;
  assign n24906 = ~n25123 | ~P1_INSTQUEUE_REG_11__5__SCAN_IN;
  assign n24908 = ~n25088 | ~P1_INSTQUEUE_REG_2__5__SCAN_IN;
  assign n24907 = ~n25089 | ~P1_INSTQUEUE_REG_12__5__SCAN_IN;
  assign n24909 = ~n24908 | ~n24907;
  assign n24913 = ~n24911 | ~P1_INSTQUEUE_REG_13__5__SCAN_IN;
  assign n24912 = ~n25196 | ~P1_INSTQUEUE_REG_0__5__SCAN_IN;
  assign n24916 = ~n24913 | ~n24912;
  assign n24914 = ~P1_INSTQUEUE_REG_5__5__SCAN_IN;
  assign n24915 = ~n25065 & ~n24914;
  assign n24918 = ~n24916 & ~n24915;
  assign n24926 = ~n24918 | ~n24917;
  assign n24920 = ~n24972 | ~P1_INSTQUEUE_REG_7__5__SCAN_IN;
  assign n24922 = ~n26629 | ~P1_INSTQUEUE_REG_10__5__SCAN_IN;
  assign n24921 = ~n24976 | ~P1_INSTQUEUE_REG_14__5__SCAN_IN;
  assign n24966 = ~n24929 & ~n25011;
  assign n24931 = ~n25100 | ~P1_INSTQUEUE_REG_13__2__SCAN_IN;
  assign n24930 = ~n25196 | ~P1_INSTQUEUE_REG_0__2__SCAN_IN;
  assign n24933 = ~n24931 | ~n24930;
  assign n25513 = ~P1_INSTQUEUE_REG_5__2__SCAN_IN;
  assign n24932 = ~n25065 & ~n25513;
  assign n24935 = ~n24933 & ~n24932;
  assign n24934 = n22832 | n25199;
  assign n24944 = ~n24935 | ~n24934;
  assign n24938 = ~n26851 | ~P1_INSTQUEUE_REG_7__2__SCAN_IN;
  assign n24937 = ~n24973 | ~P1_INSTQUEUE_REG_8__2__SCAN_IN;
  assign n24942 = n24938 & n24937;
  assign n24940 = ~n26629 | ~P1_INSTQUEUE_REG_10__2__SCAN_IN;
  assign n24939 = ~n24976 | ~P1_INSTQUEUE_REG_14__2__SCAN_IN;
  assign n24941 = n24940 & n24939;
  assign n24943 = ~n24942 | ~n24941;
  assign n24946 = ~n24898 | ~P1_INSTQUEUE_REG_1__2__SCAN_IN;
  assign n24945 = ~n25118 | ~P1_INSTQUEUE_REG_4__2__SCAN_IN;
  assign n24951 = ~n24946 | ~n24945;
  assign n24949 = ~n24947 | ~P1_INSTQUEUE_REG_9__2__SCAN_IN;
  assign n24948 = ~n22826 | ~P1_INSTQUEUE_REG_15__2__SCAN_IN;
  assign n24950 = ~n24949 | ~n24948;
  assign n24959 = ~n24951 & ~n24950;
  assign n24953 = ~n24989 | ~P1_INSTQUEUE_REG_11__2__SCAN_IN;
  assign n24952 = ~n25085 | ~P1_INSTQUEUE_REG_3__2__SCAN_IN;
  assign n24957 = ~n24953 | ~n24952;
  assign n24955 = ~n25088 | ~P1_INSTQUEUE_REG_2__2__SCAN_IN;
  assign n24954 = ~n25089 | ~P1_INSTQUEUE_REG_12__2__SCAN_IN;
  assign n24956 = ~n24955 | ~n24954;
  assign n24958 = ~n24957 & ~n24956;
  assign n24960 = n24959 & n24958;
  assign n24963 = ~n25609 | ~n25685;
  assign n24964 = ~n24963 | ~n25014;
  assign n25021 = ~n44864 | ~n24964;
  assign n24971 = ~n22833 & ~n25066;
  assign n24968 = ~n24911 | ~P1_INSTQUEUE_REG_13__1__SCAN_IN;
  assign n24967 = ~n25196 | ~P1_INSTQUEUE_REG_0__1__SCAN_IN;
  assign n24970 = ~n23979 | ~n23958;
  assign n24982 = ~n24971 & ~n24970;
  assign n24975 = ~n26851 | ~P1_INSTQUEUE_REG_7__1__SCAN_IN;
  assign n24974 = ~n26630 | ~P1_INSTQUEUE_REG_8__1__SCAN_IN;
  assign n24980 = ~n24975 | ~n24974;
  assign n24978 = ~n26629 | ~P1_INSTQUEUE_REG_10__1__SCAN_IN;
  assign n24977 = ~n24976 | ~P1_INSTQUEUE_REG_14__1__SCAN_IN;
  assign n24979 = ~n24978 | ~n24977;
  assign n24981 = ~n24980 & ~n24979;
  assign n24999 = ~n24982 | ~n24981;
  assign n24984 = ~n24898 | ~P1_INSTQUEUE_REG_1__1__SCAN_IN;
  assign n24983 = ~n25118 | ~P1_INSTQUEUE_REG_4__1__SCAN_IN;
  assign n24988 = ~n24984 | ~n24983;
  assign n24985 = ~n22826 | ~P1_INSTQUEUE_REG_15__1__SCAN_IN;
  assign n24987 = ~n24986 | ~n24985;
  assign n24997 = ~n24988 & ~n24987;
  assign n24991 = ~n24989 | ~P1_INSTQUEUE_REG_11__1__SCAN_IN;
  assign n24990 = ~n25085 | ~P1_INSTQUEUE_REG_3__1__SCAN_IN;
  assign n24995 = ~n24991 | ~n24990;
  assign n24993 = ~n25088 | ~P1_INSTQUEUE_REG_2__1__SCAN_IN;
  assign n24992 = ~n25089 | ~P1_INSTQUEUE_REG_12__1__SCAN_IN;
  assign n24994 = ~n24993 | ~n24992;
  assign n24996 = ~n24995 & ~n24994;
  assign n24998 = ~n24997 | ~n24996;
  assign n25018 = ~n25685;
  assign n25000 = ~n25018 | ~n25022;
  assign n25041 = n26914 | n26986;
  assign n25034 = ~n25003 | ~P1_STATE2_REG_0__SCAN_IN;
  assign n25053 = ~n25018 | ~n25609;
  assign n25832 = ~n25017;
  assign n25007 = n25053 | n25832;
  assign n25005 = ~n25004 | ~n25685;
  assign n25015 = ~n25005 | ~n25022;
  assign n25010 = ~n43131 | ~n26986;
  assign n25731 = ~n25010 | ~n25055;
  assign n25693 = ~n25731 | ~n25661;
  assign n25012 = ~n25055;
  assign n31438 = ~n25013 | ~n25012;
  assign n25599 = ~n43116;
  assign n25691 = ~n26986 | ~n25599;
  assign n31568 = n43101 & n26986;
  assign n25029 = ~n25016 | ~P1_STATE2_REG_0__SCAN_IN;
  assign n25019 = ~n43146 | ~n25042;
  assign n25020 = n25019 & n31515;
  assign n25025 = n25021 & n25020;
  assign n25024 = ~n25660 | ~n25054;
  assign n25026 = n26914 & n43101;
  assign n25028 = ~n25027 | ~n25134;
  assign n30634 = ~n44744 | ~n44851;
  assign n25031 = n44152 | n30634;
  assign n25185 = ~n31573 | ~P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN;
  assign n25032 = n25031 & n25185;
  assign n25035 = ~n25033 | ~n25032;
  assign n25187 = ~n25034;
  assign n25038 = ~n30634 | ~n44308;
  assign n25036 = ~n31573;
  assign n25037 = ~n25036 | ~P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n25039 = ~n25038 | ~n25037;
  assign n25703 = ~n22839 | ~n25042;
  assign n42393 = ~n43057 | ~n42760;
  assign n44748 = ~n44744;
  assign n25044 = ~n44748 & ~n44851;
  assign n25045 = n42393 & n25044;
  assign n25047 = ~n25703 | ~n25045;
  assign n25051 = ~n25047 & ~n25046;
  assign n25049 = ~n25048;
  assign n25050 = ~n25049 | ~n42760;
  assign n25061 = n25051 & n25050;
  assign n25059 = ~n25052 | ~n42372;
  assign n25056 = ~n30440 | ~n25054;
  assign n25057 = ~n25056 | ~n27579;
  assign n31497 = ~n42372;
  assign n25058 = ~n25057 | ~n31497;
  assign n25060 = ~n25059 | ~n25058;
  assign n25064 = ~n26875 | ~P1_INSTQUEUE_REG_14__1__SCAN_IN;
  assign n25063 = ~n26876 | ~P1_INSTQUEUE_REG_1__1__SCAN_IN;
  assign n25068 = ~n25064 | ~n25063;
  assign n25067 = ~n26360 & ~n25066;
  assign n25070 = ~n25068 & ~n25067;
  assign n26483 = ~P1_INSTQUEUE_REG_7__1__SCAN_IN;
  assign n25069 = n22832 | n26483;
  assign n25078 = ~n25070 | ~n25069;
  assign n25072 = ~n26851 | ~P1_INSTQUEUE_REG_8__1__SCAN_IN;
  assign n26035 = ~n26630;
  assign n25071 = ~n26866 | ~P1_INSTQUEUE_REG_9__1__SCAN_IN;
  assign n25076 = n25072 & n25071;
  assign n25074 = ~n26707 | ~P1_INSTQUEUE_REG_11__1__SCAN_IN;
  assign n26326 = ~n24976;
  assign n25073 = ~n26759 | ~P1_INSTQUEUE_REG_15__1__SCAN_IN;
  assign n25075 = n25074 & n25073;
  assign n25077 = ~n25076 | ~n25075;
  assign n25097 = ~n25078 & ~n25077;
  assign n25080 = ~n22841 | ~P1_INSTQUEUE_REG_2__1__SCAN_IN;
  assign n25079 = ~n25118 | ~P1_INSTQUEUE_REG_5__1__SCAN_IN;
  assign n25084 = ~n25080 | ~n25079;
  assign n25082 = ~n24947 | ~P1_INSTQUEUE_REG_10__1__SCAN_IN;
  assign n31463 = ~n22826;
  assign n25081 = ~n22842 | ~P1_INSTQUEUE_REG_0__1__SCAN_IN;
  assign n25083 = ~n25082 | ~n25081;
  assign n25095 = ~n25084 & ~n25083;
  assign n25294 = ~n24989;
  assign n25087 = ~n26879 | ~P1_INSTQUEUE_REG_12__1__SCAN_IN;
  assign n25267 = ~n25085;
  assign n25086 = ~n26859 | ~P1_INSTQUEUE_REG_4__1__SCAN_IN;
  assign n25093 = ~n25087 | ~n25086;
  assign n25091 = ~n25220 | ~P1_INSTQUEUE_REG_3__1__SCAN_IN;
  assign n26349 = ~n25089;
  assign n25090 = ~n25337 | ~P1_INSTQUEUE_REG_13__1__SCAN_IN;
  assign n25092 = ~n25091 | ~n25090;
  assign n25094 = ~n25093 & ~n25092;
  assign n25096 = n25095 & n25094;
  assign n25098 = n25243 | n25399;
  assign n25102 = ~n25100 | ~P1_INSTQUEUE_REG_14__7__SCAN_IN;
  assign n25101 = ~n26759 | ~P1_INSTQUEUE_REG_15__7__SCAN_IN;
  assign n25105 = ~n25102 | ~n25101;
  assign n25104 = ~n26360 & ~n25103;
  assign n26154 = ~P1_INSTQUEUE_REG_7__7__SCAN_IN;
  assign n25106 = ~n22833 & ~n26154;
  assign n25115 = ~n25107 & ~n25106;
  assign n25109 = ~n26851 | ~P1_INSTQUEUE_REG_8__7__SCAN_IN;
  assign n25108 = ~n26866 | ~P1_INSTQUEUE_REG_9__7__SCAN_IN;
  assign n25113 = ~n25109 | ~n25108;
  assign n25111 = ~n26707 | ~P1_INSTQUEUE_REG_11__7__SCAN_IN;
  assign n25110 = ~n22842 | ~P1_INSTQUEUE_REG_0__7__SCAN_IN;
  assign n25112 = ~n25111 | ~n25110;
  assign n25114 = ~n25113 & ~n25112;
  assign n25133 = ~n25115 | ~n25114;
  assign n25117 = ~n26622 | ~P1_INSTQUEUE_REG_10__7__SCAN_IN;
  assign n25116 = ~n26869 | ~P1_INSTQUEUE_REG_2__7__SCAN_IN;
  assign n25122 = ~n25117 | ~n25116;
  assign n25465 = ~n25118;
  assign n25120 = ~n26686 | ~P1_INSTQUEUE_REG_5__7__SCAN_IN;
  assign n25119 = ~n25337 | ~P1_INSTQUEUE_REG_13__7__SCAN_IN;
  assign n25121 = ~n25120 | ~n25119;
  assign n25131 = ~n25122 & ~n25121;
  assign n25125 = ~n24989 | ~P1_INSTQUEUE_REG_12__7__SCAN_IN;
  assign n25124 = ~n26876 | ~P1_INSTQUEUE_REG_1__7__SCAN_IN;
  assign n25129 = ~n25125 | ~n25124;
  assign n25127 = ~n25088 | ~P1_INSTQUEUE_REG_3__7__SCAN_IN;
  assign n25126 = ~n26859 | ~P1_INSTQUEUE_REG_4__7__SCAN_IN;
  assign n25128 = ~n25127 | ~n25126;
  assign n25130 = ~n25129 & ~n25128;
  assign n25132 = ~n25131 | ~n25130;
  assign n25172 = n25243 | n25499;
  assign n25135 = n25462 | n25399;
  assign n25137 = n25172 & n25135;
  assign n25136 = ~n25639 | ~P1_INSTQUEUE_REG_0__1__SCAN_IN;
  assign n25138 = ~n25137 | ~n25136;
  assign n25141 = ~n26875 | ~P1_INSTQUEUE_REG_14__0__SCAN_IN;
  assign n25140 = ~n26859 | ~P1_INSTQUEUE_REG_4__0__SCAN_IN;
  assign n25143 = ~n25141 | ~n25140;
  assign n25142 = ~n26320 & ~n24750;
  assign n25146 = ~n25143 & ~n25142;
  assign n25144 = ~P1_INSTQUEUE_REG_7__0__SCAN_IN;
  assign n25145 = n22833 | n25144;
  assign n25155 = ~n25146 | ~n25145;
  assign n25149 = ~n25147 | ~P1_INSTQUEUE_REG_6__0__SCAN_IN;
  assign n25148 = ~n22842 | ~P1_INSTQUEUE_REG_0__0__SCAN_IN;
  assign n25153 = n25149 & n25148;
  assign n25151 = ~n26851 | ~P1_INSTQUEUE_REG_8__0__SCAN_IN;
  assign n25150 = ~n25337 | ~P1_INSTQUEUE_REG_13__0__SCAN_IN;
  assign n25152 = n25151 & n25150;
  assign n25154 = ~n25153 | ~n25152;
  assign n25171 = ~n25155 & ~n25154;
  assign n25157 = ~n26622 | ~P1_INSTQUEUE_REG_10__0__SCAN_IN;
  assign n25156 = ~n22841 | ~P1_INSTQUEUE_REG_2__0__SCAN_IN;
  assign n25161 = ~n25157 | ~n25156;
  assign n25159 = ~n26686 | ~P1_INSTQUEUE_REG_5__0__SCAN_IN;
  assign n25158 = ~n25220 | ~P1_INSTQUEUE_REG_3__0__SCAN_IN;
  assign n25160 = ~n25159 | ~n25158;
  assign n25169 = ~n25161 & ~n25160;
  assign n25163 = ~n26866 | ~P1_INSTQUEUE_REG_9__0__SCAN_IN;
  assign n25162 = ~n26759 | ~P1_INSTQUEUE_REG_15__0__SCAN_IN;
  assign n25167 = ~n25163 | ~n25162;
  assign n25165 = ~n24989 | ~P1_INSTQUEUE_REG_12__0__SCAN_IN;
  assign n25164 = ~n26876 | ~P1_INSTQUEUE_REG_1__0__SCAN_IN;
  assign n25166 = ~n25165 | ~n25164;
  assign n25168 = ~n25167 & ~n25166;
  assign n25170 = n25169 & n25168;
  assign n25174 = ~n25550 | ~n25398;
  assign n25177 = ~n25398;
  assign n25173 = ~n25172 | ~n25177;
  assign n25175 = ~n25174 | ~n25173;
  assign n25181 = ~n25639 | ~P1_INSTQUEUE_REG_0__0__SCAN_IN;
  assign n25176 = ~n43146 | ~n25499;
  assign n25179 = ~n25176 | ~P1_STATE2_REG_0__SCAN_IN;
  assign n25178 = n43057 & n25177;
  assign n25180 = ~n25179 & ~n25178;
  assign n25391 = ~n25181 | ~n25180;
  assign n25184 = n25183;
  assign n25186 = ~n25185 | ~n25184;
  assign n25188 = ~n25187 | ~n25186;
  assign n25236 = ~n25189 | ~P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign n25190 = ~n25189;
  assign n25191 = ~n25190 | ~n44132;
  assign n25238 = ~n30634;
  assign n25193 = ~n43081 | ~n25238;
  assign n25192 = ~n31573 | ~P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign n25198 = ~n26875 | ~P1_INSTQUEUE_REG_14__2__SCAN_IN;
  assign n26750 = ~n25196;
  assign n26876 = ~n26750;
  assign n25197 = ~n26876 | ~P1_INSTQUEUE_REG_1__2__SCAN_IN;
  assign n25201 = ~n25198 | ~n25197;
  assign n25200 = ~n26360 & ~n25199;
  assign n25203 = ~n25201 & ~n25200;
  assign n26612 = ~P1_INSTQUEUE_REG_7__2__SCAN_IN;
  assign n25202 = n22833 | n26612;
  assign n25211 = ~n25203 | ~n25202;
  assign n25205 = ~n26851 | ~P1_INSTQUEUE_REG_8__2__SCAN_IN;
  assign n25204 = ~n26866 | ~P1_INSTQUEUE_REG_9__2__SCAN_IN;
  assign n25209 = n25205 & n25204;
  assign n25207 = ~n26707 | ~P1_INSTQUEUE_REG_11__2__SCAN_IN;
  assign n25206 = ~n26759 | ~P1_INSTQUEUE_REG_15__2__SCAN_IN;
  assign n25208 = n25207 & n25206;
  assign n25210 = ~n25209 | ~n25208;
  assign n25228 = ~n25211 & ~n25210;
  assign n25213 = ~n22841 | ~P1_INSTQUEUE_REG_2__2__SCAN_IN;
  assign n25212 = ~n26858 | ~P1_INSTQUEUE_REG_5__2__SCAN_IN;
  assign n25217 = ~n25213 | ~n25212;
  assign n25215 = ~n24947 | ~P1_INSTQUEUE_REG_10__2__SCAN_IN;
  assign n25214 = ~n22842 | ~P1_INSTQUEUE_REG_0__2__SCAN_IN;
  assign n25216 = ~n25215 | ~n25214;
  assign n25226 = ~n25217 & ~n25216;
  assign n25219 = ~n26879 | ~P1_INSTQUEUE_REG_12__2__SCAN_IN;
  assign n25218 = ~n26859 | ~P1_INSTQUEUE_REG_4__2__SCAN_IN;
  assign n25224 = ~n25219 | ~n25218;
  assign n25481 = ~n25088;
  assign n25220 = ~n25481;
  assign n25222 = ~n25220 | ~P1_INSTQUEUE_REG_3__2__SCAN_IN;
  assign n25337 = ~n26349;
  assign n25221 = ~n25337 | ~P1_INSTQUEUE_REG_13__2__SCAN_IN;
  assign n25223 = ~n25222 | ~n25221;
  assign n25225 = ~n25224 & ~n25223;
  assign n25227 = n25226 & n25225;
  assign n25229 = n25243 | n25414;
  assign n25231 = ~n25639 | ~P1_INSTQUEUE_REG_0__2__SCAN_IN;
  assign n25230 = n25462 | n25414;
  assign n44307 = ~P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign n43729 = ~n44307 & ~P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN;
  assign n43718 = ~n43729 | ~P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n25237 = ~n25236 | ~P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN;
  assign n44153 = ~n43718 | ~n25237;
  assign n25240 = ~n44153 | ~n25238;
  assign n25239 = ~n31573 | ~P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN;
  assign n25277 = ~n25639 | ~P1_INSTQUEUE_REG_0__3__SCAN_IN;
  assign n25245 = ~n26851 | ~P1_INSTQUEUE_REG_8__3__SCAN_IN;
  assign n25244 = ~n22842 | ~P1_INSTQUEUE_REG_0__3__SCAN_IN;
  assign n25247 = n25245 & n25244;
  assign n25246 = ~n25147 | ~P1_INSTQUEUE_REG_6__3__SCAN_IN;
  assign n25250 = ~n25247 | ~n25246;
  assign n25248 = ~P1_INSTQUEUE_REG_7__3__SCAN_IN;
  assign n25249 = ~n22833 & ~n25248;
  assign n25258 = ~n25250 & ~n25249;
  assign n25252 = ~n26866 | ~P1_INSTQUEUE_REG_9__3__SCAN_IN;
  assign n25251 = ~n26759 | ~P1_INSTQUEUE_REG_15__3__SCAN_IN;
  assign n25256 = ~n25252 | ~n25251;
  assign n25254 = ~n26707 | ~P1_INSTQUEUE_REG_11__3__SCAN_IN;
  assign n25253 = ~n25337 | ~P1_INSTQUEUE_REG_13__3__SCAN_IN;
  assign n25255 = ~n25254 | ~n25253;
  assign n25257 = ~n25256 & ~n25255;
  assign n25275 = ~n25258 | ~n25257;
  assign n25260 = ~n26879 | ~P1_INSTQUEUE_REG_12__3__SCAN_IN;
  assign n25259 = ~n25220 | ~P1_INSTQUEUE_REG_3__3__SCAN_IN;
  assign n25264 = ~n25260 | ~n25259;
  assign n25262 = ~n24947 | ~P1_INSTQUEUE_REG_10__3__SCAN_IN;
  assign n26577 = ~n26750;
  assign n25261 = ~n26577 | ~P1_INSTQUEUE_REG_1__3__SCAN_IN;
  assign n25263 = ~n25262 | ~n25261;
  assign n25273 = ~n25264 & ~n25263;
  assign n25266 = ~n26875 | ~P1_INSTQUEUE_REG_14__3__SCAN_IN;
  assign n25265 = ~n26686 | ~P1_INSTQUEUE_REG_5__3__SCAN_IN;
  assign n25271 = ~n25266 | ~n25265;
  assign n25269 = ~n22841 | ~P1_INSTQUEUE_REG_2__3__SCAN_IN;
  assign n25268 = ~n26859 | ~P1_INSTQUEUE_REG_4__3__SCAN_IN;
  assign n25270 = ~n25269 | ~n25268;
  assign n25272 = ~n25271 & ~n25270;
  assign n25274 = ~n25273 | ~n25272;
  assign n25276 = ~n25629 | ~n25426;
  assign n25312 = ~n25639 | ~P1_INSTQUEUE_REG_0__4__SCAN_IN;
  assign n25280 = ~n26622 | ~P1_INSTQUEUE_REG_10__4__SCAN_IN;
  assign n25279 = ~n22841 | ~P1_INSTQUEUE_REG_2__4__SCAN_IN;
  assign n25282 = n25280 & n25279;
  assign n25281 = ~n26686 | ~P1_INSTQUEUE_REG_5__4__SCAN_IN;
  assign n25285 = ~n25282 | ~n25281;
  assign n25283 = ~P1_INSTQUEUE_REG_7__4__SCAN_IN;
  assign n25284 = ~n22832 & ~n25283;
  assign n25293 = ~n25285 & ~n25284;
  assign n25287 = ~n25147 | ~P1_INSTQUEUE_REG_6__4__SCAN_IN;
  assign n25286 = ~n26859 | ~P1_INSTQUEUE_REG_4__4__SCAN_IN;
  assign n25291 = ~n25287 | ~n25286;
  assign n25289 = ~n24972 | ~P1_INSTQUEUE_REG_8__4__SCAN_IN;
  assign n25288 = ~n22842 | ~P1_INSTQUEUE_REG_0__4__SCAN_IN;
  assign n25290 = ~n25289 | ~n25288;
  assign n25292 = ~n25291 & ~n25290;
  assign n25310 = ~n25293 | ~n25292;
  assign n26879 = ~n25294;
  assign n25296 = ~n26879 | ~P1_INSTQUEUE_REG_12__4__SCAN_IN;
  assign n25295 = ~n26759 | ~P1_INSTQUEUE_REG_15__4__SCAN_IN;
  assign n25300 = ~n25296 | ~n25295;
  assign n25298 = ~n26707 | ~P1_INSTQUEUE_REG_11__4__SCAN_IN;
  assign n25297 = ~n26817 | ~P1_INSTQUEUE_REG_3__4__SCAN_IN;
  assign n25299 = ~n25298 | ~n25297;
  assign n25308 = ~n25300 & ~n25299;
  assign n25302 = ~n26875 | ~P1_INSTQUEUE_REG_14__4__SCAN_IN;
  assign n25301 = ~n25337 | ~P1_INSTQUEUE_REG_13__4__SCAN_IN;
  assign n25306 = ~n25302 | ~n25301;
  assign n25304 = ~n26866 | ~P1_INSTQUEUE_REG_9__4__SCAN_IN;
  assign n25303 = ~n26876 | ~P1_INSTQUEUE_REG_1__4__SCAN_IN;
  assign n25305 = ~n25304 | ~n25303;
  assign n25307 = ~n25306 & ~n25305;
  assign n25309 = ~n25308 | ~n25307;
  assign n25311 = ~n25629 | ~n25436;
  assign n25347 = ~n25639 | ~P1_INSTQUEUE_REG_0__5__SCAN_IN;
  assign n25313 = ~P1_INSTQUEUE_REG_7__5__SCAN_IN;
  assign n25320 = ~n22832 & ~n25313;
  assign n25316 = ~n26875 | ~P1_INSTQUEUE_REG_14__5__SCAN_IN;
  assign n25315 = ~n26577 | ~P1_INSTQUEUE_REG_1__5__SCAN_IN;
  assign n25318 = ~n25316 | ~n25315;
  assign n25317 = ~n26360 & ~n26748;
  assign n25319 = n25318 | n25317;
  assign n25328 = ~n25320 & ~n25319;
  assign n25322 = ~n26851 | ~P1_INSTQUEUE_REG_8__5__SCAN_IN;
  assign n25321 = ~n26866 | ~P1_INSTQUEUE_REG_9__5__SCAN_IN;
  assign n25326 = ~n25322 | ~n25321;
  assign n25324 = ~n26707 | ~P1_INSTQUEUE_REG_11__5__SCAN_IN;
  assign n25323 = ~n26759 | ~P1_INSTQUEUE_REG_15__5__SCAN_IN;
  assign n25325 = ~n25324 | ~n25323;
  assign n25327 = ~n25326 & ~n25325;
  assign n25345 = ~n25328 | ~n25327;
  assign n25330 = ~n22841 | ~P1_INSTQUEUE_REG_2__5__SCAN_IN;
  assign n26686 = ~n25465;
  assign n25329 = ~n26686 | ~P1_INSTQUEUE_REG_5__5__SCAN_IN;
  assign n25334 = ~n25330 | ~n25329;
  assign n25332 = ~n26622 | ~P1_INSTQUEUE_REG_10__5__SCAN_IN;
  assign n25331 = ~n22842 | ~P1_INSTQUEUE_REG_0__5__SCAN_IN;
  assign n25333 = ~n25332 | ~n25331;
  assign n25343 = ~n25334 & ~n25333;
  assign n25336 = ~n26879 | ~P1_INSTQUEUE_REG_12__5__SCAN_IN;
  assign n25335 = ~n26859 | ~P1_INSTQUEUE_REG_4__5__SCAN_IN;
  assign n25341 = ~n25336 | ~n25335;
  assign n25339 = ~n26817 | ~P1_INSTQUEUE_REG_3__5__SCAN_IN;
  assign n25338 = ~n25337 | ~P1_INSTQUEUE_REG_13__5__SCAN_IN;
  assign n25340 = ~n25339 | ~n25338;
  assign n25342 = ~n25341 & ~n25340;
  assign n25344 = ~n25343 | ~n25342;
  assign n25346 = ~n25629 | ~n25443;
  assign n25380 = ~n25639 | ~P1_INSTQUEUE_REG_0__6__SCAN_IN;
  assign n25349 = ~n26622 | ~P1_INSTQUEUE_REG_10__6__SCAN_IN;
  assign n25348 = ~n26866 | ~P1_INSTQUEUE_REG_9__6__SCAN_IN;
  assign n25351 = n25349 & n25348;
  assign n25350 = ~n26818 | ~P1_INSTQUEUE_REG_13__6__SCAN_IN;
  assign n25353 = ~n25351 | ~n25350;
  assign n26800 = ~P1_INSTQUEUE_REG_7__6__SCAN_IN;
  assign n25352 = ~n22833 & ~n26800;
  assign n25361 = ~n25353 & ~n25352;
  assign n25355 = ~n22841 | ~P1_INSTQUEUE_REG_2__6__SCAN_IN;
  assign n25354 = ~n26577 | ~P1_INSTQUEUE_REG_1__6__SCAN_IN;
  assign n25359 = ~n25355 | ~n25354;
  assign n26870 = ~n26326;
  assign n25357 = ~n26870 | ~P1_INSTQUEUE_REG_15__6__SCAN_IN;
  assign n25356 = ~n22842 | ~P1_INSTQUEUE_REG_0__6__SCAN_IN;
  assign n25358 = ~n25357 | ~n25356;
  assign n25360 = ~n25359 & ~n25358;
  assign n25378 = ~n25361 | ~n25360;
  assign n25364 = ~n25147 | ~P1_INSTQUEUE_REG_6__6__SCAN_IN;
  assign n25363 = ~n26851 | ~P1_INSTQUEUE_REG_8__6__SCAN_IN;
  assign n25368 = ~n25364 | ~n25363;
  assign n25366 = ~n26707 | ~P1_INSTQUEUE_REG_11__6__SCAN_IN;
  assign n26817 = ~n25481;
  assign n25365 = ~n26817 | ~P1_INSTQUEUE_REG_3__6__SCAN_IN;
  assign n25367 = ~n25366 | ~n25365;
  assign n25376 = ~n25368 & ~n25367;
  assign n25370 = ~n26875 | ~P1_INSTQUEUE_REG_14__6__SCAN_IN;
  assign n26858 = ~n25465;
  assign n25369 = ~n26858 | ~P1_INSTQUEUE_REG_5__6__SCAN_IN;
  assign n25374 = ~n25370 | ~n25369;
  assign n25372 = ~n26879 | ~P1_INSTQUEUE_REG_12__6__SCAN_IN;
  assign n25371 = ~n26859 | ~P1_INSTQUEUE_REG_4__6__SCAN_IN;
  assign n25373 = ~n25372 | ~n25371;
  assign n25375 = ~n25374 & ~n25373;
  assign n25377 = ~n25376 | ~n25375;
  assign n25379 = ~n25629 | ~n25455;
  assign n25383 = ~n25380 | ~n25379;
  assign n25381 = ~n25383;
  assign n25384 = ~n25382 | ~n25381;
  assign n25390 = ~n25916 | ~n25601;
  assign n25413 = n25399 | n25398;
  assign n25428 = ~n25413 | ~n25414;
  assign n25437 = ~n25428 | ~n25426;
  assign n25385 = ~n25436;
  assign n25444 = n25437 | n25385;
  assign n25386 = ~n25443;
  assign n25456 = ~n25444 & ~n25386;
  assign n25387 = ~n25456;
  assign n25388 = ~n25387 ^ n25455;
  assign n25389 = ~n25388 | ~n31568;
  assign n25396 = ~n25868 | ~n25601;
  assign n25394 = ~n31568 | ~n25398;
  assign n25419 = n26986 | n43131;
  assign n25395 = n25394 & n25419;
  assign n42948 = ~n25396 | ~n25395;
  assign n25404 = n25397 | n25549;
  assign n25400 = ~n25399 ^ n25398;
  assign n25402 = n44843 | n25400;
  assign n25401 = ~n25661 & ~n43161;
  assign n25403 = n25402 & n25401;
  assign n25407 = n25404 & n25403;
  assign n25405 = ~P1_INSTADDRPOINTER_REG_1__SCAN_IN;
  assign n25408 = n25407 | n25406;
  assign n25409 = ~n31009;
  assign n31010 = ~n25409 | ~P1_INSTADDRPOINTER_REG_2__SCAN_IN;
  assign n25410 = ~P1_INSTADDRPOINTER_REG_2__SCAN_IN;
  assign n25423 = ~n31009 | ~n25410;
  assign n25416 = ~n25413;
  assign n25415 = ~n25414;
  assign n25417 = ~n25416 | ~n25415;
  assign n25418 = ~n25417 | ~n25428;
  assign n25420 = ~n25418 | ~n31568;
  assign n25421 = n25420 & n25419;
  assign n25425 = ~n25424;
  assign n25431 = ~n25885 | ~n25601;
  assign n25427 = ~n25426;
  assign n25429 = ~n25428 ^ n25427;
  assign n25430 = ~n25429 | ~n31568;
  assign n25432 = ~n31012 | ~P1_INSTADDRPOINTER_REG_3__SCAN_IN;
  assign n25434 = ~n31012;
  assign n25433 = ~P1_INSTADDRPOINTER_REG_3__SCAN_IN;
  assign n25438 = ~n25437 ^ n25436;
  assign n25439 = ~n25438 | ~n31568;
  assign n25442 = ~n42899;
  assign n25441 = ~P1_INSTADDRPOINTER_REG_4__SCAN_IN;
  assign n25445 = ~n25444 ^ n25443;
  assign n25446 = ~n25445 | ~n31568;
  assign n25447 = P1_INSTADDRPOINTER_REG_4__SCAN_IN & P1_INSTADDRPOINTER_REG_5__SCAN_IN;
  assign n25448 = ~n42899 | ~n25447;
  assign n25450 = ~P1_INSTQUEUE_REG_0__7__SCAN_IN;
  assign n25453 = ~n25608 & ~n25450;
  assign n25451 = n25462 | n25457;
  assign n25452 = ~n25550 | ~n25451;
  assign n25454 = ~n25453 & ~n25452;
  assign n25460 = ~n22940 | ~n25601;
  assign n25501 = ~n25456 | ~n25455;
  assign n25458 = ~n25501 ^ n25457;
  assign n25459 = n25458 | n44843;
  assign n30947 = ~n25461 | ~P1_INSTADDRPOINTER_REG_7__SCAN_IN;
  assign n25463 = ~n25608 | ~n25462;
  assign n25542 = ~n25550;
  assign n25467 = ~n26622 | ~P1_INSTQUEUE_REG_11__0__SCAN_IN;
  assign n25466 = ~n26858 | ~P1_INSTQUEUE_REG_6__0__SCAN_IN;
  assign n25471 = ~n25467 | ~n25466;
  assign n26707 = ~n26320;
  assign n25469 = ~n26707 | ~P1_INSTQUEUE_REG_12__0__SCAN_IN;
  assign n25468 = ~n26870 | ~P1_INSTQUEUE_REG_0__0__SCAN_IN;
  assign n25470 = ~n25469 | ~n25468;
  assign n25479 = ~n25471 & ~n25470;
  assign n25473 = ~n26875 | ~P1_INSTQUEUE_REG_15__0__SCAN_IN;
  assign n25472 = ~n22841 | ~P1_INSTQUEUE_REG_3__0__SCAN_IN;
  assign n25477 = ~n25473 | ~n25472;
  assign n25475 = ~n26577 | ~P1_INSTQUEUE_REG_2__0__SCAN_IN;
  assign n25474 = ~n26818 | ~P1_INSTQUEUE_REG_14__0__SCAN_IN;
  assign n25476 = ~n25475 | ~n25474;
  assign n25478 = ~n25477 & ~n25476;
  assign n25480 = n25479 & n25478;
  assign n25497 = ~n25550 | ~n25480;
  assign n25483 = ~n26879 | ~P1_INSTQUEUE_REG_13__0__SCAN_IN;
  assign n25482 = ~n26817 | ~P1_INSTQUEUE_REG_4__0__SCAN_IN;
  assign n25487 = ~n25483 | ~n25482;
  assign n25485 = ~n25147 | ~P1_INSTQUEUE_REG_7__0__SCAN_IN;
  assign n25484 = ~n26859 | ~P1_INSTQUEUE_REG_5__0__SCAN_IN;
  assign n25486 = ~n25485 | ~n25484;
  assign n25495 = ~n25487 & ~n25486;
  assign n25489 = ~n26630 | ~P1_INSTQUEUE_REG_10__0__SCAN_IN;
  assign n25488 = ~n22842 | ~P1_INSTQUEUE_REG_1__0__SCAN_IN;
  assign n25493 = ~n25489 | ~n25488;
  assign n26847 = ~n22833;
  assign n25491 = ~n26847 | ~P1_INSTQUEUE_REG_8__0__SCAN_IN;
  assign n25490 = ~n26753 | ~P1_INSTQUEUE_REG_9__0__SCAN_IN;
  assign n25492 = ~n25491 | ~n25490;
  assign n25494 = ~n25493 & ~n25492;
  assign n25496 = ~n25495 | ~n25494;
  assign n25500 = ~n31568 | ~n25499;
  assign n25502 = n25501 | n25500;
  assign n30951 = ~n30950 | ~P1_INSTADDRPOINTER_REG_8__SCAN_IN;
  assign n25503 = n30947 & n30951;
  assign n30949 = ~P1_INSTADDRPOINTER_REG_8__SCAN_IN;
  assign n25506 = ~n25504 | ~n30949;
  assign n31332 = ~P1_INSTADDRPOINTER_REG_9__SCAN_IN;
  assign n25505 = ~n30953 | ~n31332;
  assign n25508 = n30953 | n31332;
  assign n25509 = ~P1_INSTQUEUE_REG_0__2__SCAN_IN;
  assign n25511 = ~n26326 & ~n25509;
  assign n26617 = ~P1_INSTQUEUE_REG_10__2__SCAN_IN;
  assign n25510 = ~n26035 & ~n26617;
  assign n25517 = ~n25511 & ~n25510;
  assign n25512 = ~P1_INSTQUEUE_REG_14__2__SCAN_IN;
  assign n25515 = ~n26349 & ~n25512;
  assign n25514 = ~n25267 & ~n25513;
  assign n25516 = ~n25515 & ~n25514;
  assign n25521 = ~n25517 | ~n25516;
  assign n26875 = ~n26482;
  assign n25519 = ~n26875 | ~P1_INSTQUEUE_REG_15__2__SCAN_IN;
  assign n25518 = ~n26869 | ~P1_INSTQUEUE_REG_3__2__SCAN_IN;
  assign n25520 = ~n25519 | ~n25518;
  assign n25541 = ~n25521 & ~n25520;
  assign n25523 = ~n26879 | ~P1_INSTQUEUE_REG_13__2__SCAN_IN;
  assign n25522 = ~n26817 | ~P1_INSTQUEUE_REG_4__2__SCAN_IN;
  assign n25539 = ~n25523 | ~n25522;
  assign n25525 = ~n26858 | ~P1_INSTQUEUE_REG_6__2__SCAN_IN;
  assign n25524 = ~n26577 | ~P1_INSTQUEUE_REG_2__2__SCAN_IN;
  assign n25529 = ~n25525 | ~n25524;
  assign n25527 = ~n26622 | ~P1_INSTQUEUE_REG_11__2__SCAN_IN;
  assign n25526 = ~n26707 | ~P1_INSTQUEUE_REG_12__2__SCAN_IN;
  assign n25528 = ~n25527 | ~n25526;
  assign n25537 = ~n25529 & ~n25528;
  assign n25531 = ~n25147 | ~P1_INSTQUEUE_REG_7__2__SCAN_IN;
  assign n25530 = ~n26753 | ~P1_INSTQUEUE_REG_9__2__SCAN_IN;
  assign n25535 = ~n25531 | ~n25530;
  assign n25533 = ~n26847 | ~P1_INSTQUEUE_REG_8__2__SCAN_IN;
  assign n25532 = ~n22842 | ~P1_INSTQUEUE_REG_1__2__SCAN_IN;
  assign n25534 = ~n25533 | ~n25532;
  assign n25536 = ~n25535 & ~n25534;
  assign n25538 = ~n25537 | ~n25536;
  assign n25540 = ~n25539 & ~n25538;
  assign n25543 = ~n25541 | ~n25540;
  assign n30927 = ~P1_INSTADDRPOINTER_REG_10__SCAN_IN;
  assign n25545 = ~n30928 | ~n30927;
  assign n31287 = ~P1_INSTADDRPOINTER_REG_11__SCAN_IN;
  assign n25544 = ~n30953 | ~n31287;
  assign n30879 = ~n25545 | ~n25544;
  assign n31233 = ~P1_INSTADDRPOINTER_REG_14__SCAN_IN;
  assign n25546 = n30953 & n31233;
  assign n30903 = ~n30953 ^ P1_INSTADDRPOINTER_REG_13__SCAN_IN;
  assign n31286 = ~P1_INSTADDRPOINTER_REG_12__SCAN_IN;
  assign n30907 = ~n30953 | ~n31286;
  assign n31261 = ~P1_INSTADDRPOINTER_REG_13__SCAN_IN;
  assign n25548 = n30953 | n31233;
  assign n31216 = ~P1_INSTADDRPOINTER_REG_15__SCAN_IN;
  assign n25552 = ~P1_INSTADDRPOINTER_REG_16__SCAN_IN;
  assign n30844 = ~n30821 ^ n25552;
  assign n30864 = n30821 & n31216;
  assign n31189 = ~P1_INSTADDRPOINTER_REG_17__SCAN_IN;
  assign n30823 = n30821 & n31189;
  assign n30898 = n30953 | n31287;
  assign n25553 = ~P1_INSTADDRPOINTER_REG_17__SCAN_IN & ~P1_INSTADDRPOINTER_REG_16__SCAN_IN;
  assign n25554 = ~n30821 & ~n25553;
  assign n30804 = ~n30821 ^ P1_INSTADDRPOINTER_REG_18__SCAN_IN;
  assign n31134 = P1_INSTADDRPOINTER_REG_19__SCAN_IN & P1_INSTADDRPOINTER_REG_20__SCAN_IN;
  assign n25557 = ~P1_INSTADDRPOINTER_REG_21__SCAN_IN & ~P1_INSTADDRPOINTER_REG_20__SCAN_IN;
  assign n25556 = ~P1_INSTADDRPOINTER_REG_19__SCAN_IN & ~P1_INSTADDRPOINTER_REG_18__SCAN_IN;
  assign n25560 = ~P1_INSTADDRPOINTER_REG_25__SCAN_IN & ~P1_INSTADDRPOINTER_REG_23__SCAN_IN;
  assign n31105 = ~P1_INSTADDRPOINTER_REG_24__SCAN_IN;
  assign n30706 = n25560 & n31105;
  assign n31078 = ~P1_INSTADDRPOINTER_REG_26__SCAN_IN;
  assign n31075 = P1_INSTADDRPOINTER_REG_23__SCAN_IN & P1_INSTADDRPOINTER_REG_24__SCAN_IN;
  assign n30674 = ~n31075 | ~P1_INSTADDRPOINTER_REG_25__SCAN_IN;
  assign n25842 = ~n30674;
  assign n25561 = ~n25842 | ~P1_INSTADDRPOINTER_REG_26__SCAN_IN;
  assign n31063 = ~P1_INSTADDRPOINTER_REG_27__SCAN_IN;
  assign n30683 = ~P1_INSTADDRPOINTER_REG_28__SCAN_IN;
  assign n31048 = ~n31063 | ~n30683;
  assign n25563 = ~n31048;
  assign n31049 = P1_INSTADDRPOINTER_REG_27__SCAN_IN & P1_INSTADDRPOINTER_REG_28__SCAN_IN;
  assign n31035 = ~P1_INSTADDRPOINTER_REG_29__SCAN_IN;
  assign n25564 = ~P1_INSTADDRPOINTER_REG_29__SCAN_IN & ~P1_INSTADDRPOINTER_REG_30__SCAN_IN;
  assign n25567 = ~n23166 & ~n25564;
  assign n25565 = ~n25567;
  assign n25566 = ~n23166 ^ P1_INSTADDRPOINTER_REG_31__SCAN_IN;
  assign n25568 = ~n23742 & ~P1_INSTADDRPOINTER_REG_30__SCAN_IN;
  assign n25569 = ~n25568 & ~n25567;
  assign n25570 = ~n25569 & ~P1_INSTADDRPOINTER_REG_31__SCAN_IN;
  assign n44522 = ~P1_STATE_REG_0__SCAN_IN;
  assign n44841 = ~n23041 | ~n44522;
  assign n25598 = ~n44841 | ~n42760;
  assign n25588 = ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN ^ P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN;
  assign n25590 = ~n25588 | ~n25587;
  assign n25571 = ~n43799 | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign n25581 = ~n25590 | ~n25571;
  assign n25573 = ~n44132 | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n25572 = ~n31488 | ~P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign n25583 = ~n25581 | ~n25580;
  assign n25578 = ~n25583 | ~n25573;
  assign n25575 = n25574;
  assign n25576 = ~n25575 | ~P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN;
  assign n25585 = ~n25578 | ~n25577;
  assign n25579 = n25578 | n25577;
  assign n25632 = ~n25585 | ~n25579;
  assign n25582 = n25581 | n25580;
  assign n25627 = ~n25583 | ~n25582;
  assign n25586 = ~n25632 & ~n25627;
  assign n25640 = ~n25592 | ~n25593;
  assign n25591 = ~n25586 | ~n25640;
  assign n25589 = n25588 | n25587;
  assign n25613 = ~n25590 | ~n25589;
  assign n31512 = ~n25596 | ~n25647;
  assign n26911 = ~n31417 | ~n31582;
  assign n25597 = ~n26911;
  assign n25600 = ~n25598 | ~n25597;
  assign n25659 = ~n25600 | ~n25599;
  assign n25643 = ~n25639 | ~n25601;
  assign n25602 = ~n25643;
  assign n25636 = ~n25602 | ~n25632;
  assign n25605 = ~n25608 | ~n25627;
  assign n25603 = ~n25627;
  assign n25604 = ~n25645 | ~n25603;
  assign n25607 = ~n25605 | ~n25604;
  assign n25606 = ~n43161 & ~n42760;
  assign n25628 = ~n42372 & ~n25606;
  assign n25626 = ~n25607 | ~n25628;
  assign n25611 = ~n25609 & ~n44851;
  assign n25610 = ~n25629 | ~n42760;
  assign n25612 = ~n25611 & ~n43101;
  assign n25625 = ~n25617 | ~n25616;
  assign n25618 = ~n25614 ^ P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n25620 = ~n43146 & ~n25618;
  assign n25622 = ~n25620 & ~n25619;
  assign n25621 = ~n31502;
  assign n25623 = ~n25622 | ~n25621;
  assign n25624 = n25628 & n25623;
  assign n25630 = ~n25628 & ~n25627;
  assign n25631 = ~n25630 | ~n25629;
  assign n25633 = ~n25608 | ~n25632;
  assign n25635 = ~n25634 | ~n25633;
  assign n25641 = ~n25636 | ~n25635;
  assign n25638 = ~n25637 & ~n25640;
  assign n25644 = ~n25647 & ~n25643;
  assign n25649 = ~n25648 | ~n25647;
  assign n25651 = ~n43101 | ~n44841;
  assign n26985 = n25651 & n31582;
  assign n25653 = ~n26985;
  assign n25655 = n25653 | n31439;
  assign n25654 = n25002 & n26986;
  assign n25656 = ~n25655 | ~n25654;
  assign n25657 = ~n43051 | ~n25656;
  assign n25658 = ~n25657 | ~n43116;
  assign n25676 = ~n25659 | ~n25658;
  assign n31503 = n25661 | n43057;
  assign n25663 = ~n31503;
  assign n25662 = ~n25661;
  assign n25666 = n25663 | n26910;
  assign n25665 = ~n25664;
  assign n25672 = n25666 & n25665;
  assign n25667 = n30440 & n26986;
  assign n25671 = ~n25668 | ~n25667;
  assign n25670 = ~n25669 | ~n31568;
  assign n25697 = n25671 & n25670;
  assign n25674 = ~n25672 | ~n25697;
  assign n31493 = ~n25673;
  assign n31423 = ~n25674 | ~n31493;
  assign n25684 = ~n25837;
  assign n25681 = ~n25833 & ~n43146;
  assign n25680 = ~n30633;
  assign n31451 = ~n26910 | ~n42372;
  assign n31506 = ~n25680 | ~n31451;
  assign n25682 = ~n25681 & ~n31506;
  assign n25683 = ~n25682 | ~n23094;
  assign n25690 = ~n25664 | ~n25822;
  assign n25686 = n26912 | n43116;
  assign n25687 = n25686 & n31515;
  assign n25688 = ~n25041 | ~n25687;
  assign n25689 = ~n25688 | ~n42760;
  assign n25696 = ~n25690 | ~n25689;
  assign n44842 = ~n42393;
  assign n25694 = n25692 & n25691;
  assign n25695 = ~n25694 | ~n25693;
  assign n25698 = ~n25696 & ~n25695;
  assign n25701 = n25698 & n25697;
  assign n25699 = ~n25052;
  assign n25700 = ~n25699 | ~n42372;
  assign n31444 = ~n25701 | ~n25700;
  assign n25702 = ~n31438;
  assign n25704 = ~n25702 | ~n43057;
  assign n25705 = ~n25704 | ~n25703;
  assign n25706 = ~n31444 & ~n25705;
  assign n27066 = ~n43013;
  assign n25714 = ~n31075 & ~n27066;
  assign n25712 = ~P1_INSTADDRPOINTER_REG_21__SCAN_IN | ~P1_INSTADDRPOINTER_REG_22__SCAN_IN;
  assign n27064 = ~P1_INSTADDRPOINTER_REG_12__SCAN_IN | ~P1_INSTADDRPOINTER_REG_11__SCAN_IN;
  assign n31232 = ~n27064;
  assign n25710 = ~P1_INSTADDRPOINTER_REG_9__SCAN_IN | ~P1_INSTADDRPOINTER_REG_10__SCAN_IN;
  assign n31315 = P1_INSTADDRPOINTER_REG_8__SCAN_IN & P1_INSTADDRPOINTER_REG_7__SCAN_IN;
  assign n44753 = ~P1_INSTADDRPOINTER_REG_0__SCAN_IN;
  assign n42993 = ~n44753 & ~n25405;
  assign n42965 = ~P1_INSTADDRPOINTER_REG_2__SCAN_IN & ~n42993;
  assign n42972 = ~P1_INSTADDRPOINTER_REG_4__SCAN_IN | ~P1_INSTADDRPOINTER_REG_3__SCAN_IN;
  assign n31395 = ~n42965 & ~n42972;
  assign n31381 = ~P1_INSTADDRPOINTER_REG_5__SCAN_IN | ~n31395;
  assign n31348 = ~n25449 & ~n31381;
  assign n31318 = ~n31315 | ~n31348;
  assign n31277 = ~n25710 & ~n31318;
  assign n31243 = ~n31232 | ~n31277;
  assign n31187 = ~P1_INSTADDRPOINTER_REG_16__SCAN_IN | ~P1_INSTADDRPOINTER_REG_15__SCAN_IN;
  assign n31173 = ~n31189 & ~n31187;
  assign n25711 = ~P1_INSTADDRPOINTER_REG_18__SCAN_IN | ~n31173;
  assign n31167 = ~P1_INSTADDRPOINTER_REG_14__SCAN_IN | ~P1_INSTADDRPOINTER_REG_13__SCAN_IN;
  assign n27068 = n25711 | n31167;
  assign n27072 = ~n31243 & ~n27068;
  assign n27097 = ~n31134 | ~n27072;
  assign n25840 = ~n25712 & ~n27097;
  assign n25707 = ~n25840 | ~P1_INSTADDRPOINTER_REG_23__SCAN_IN;
  assign n43014 = ~n25837 & ~n31509;
  assign n25713 = ~n25707 | ~n43014;
  assign n25708 = ~n43013 | ~n44753;
  assign n43032 = n25837 & n42947;
  assign n31248 = ~n43032;
  assign n42968 = ~P1_INSTADDRPOINTER_REG_2__SCAN_IN | ~P1_INSTADDRPOINTER_REG_1__SCAN_IN;
  assign n31404 = ~n42968 & ~n42972;
  assign n31312 = ~P1_INSTADDRPOINTER_REG_5__SCAN_IN | ~n31404;
  assign n31347 = ~n25449 & ~n31312;
  assign n31317 = ~n31347 | ~n31315;
  assign n31279 = ~n31317 & ~n25710;
  assign n27065 = ~n31279 | ~n31232;
  assign n31241 = ~n31261 & ~n27065;
  assign n31170 = ~P1_INSTADDRPOINTER_REG_14__SCAN_IN | ~n31241;
  assign n27069 = ~n31170 & ~n25711;
  assign n27096 = ~n31134 | ~n27069;
  assign n25839 = ~n27096 & ~n25712;
  assign n25715 = n43014 & n31105;
  assign n43027 = ~n43014 & ~n42961;
  assign n25720 = ~n31091 | ~n43027;
  assign n25717 = ~n25720;
  assign n31090 = ~P1_INSTADDRPOINTER_REG_25__SCAN_IN;
  assign n25716 = ~n31090 & ~n31074;
  assign n31059 = ~n25717 & ~n25716;
  assign n25718 = ~n31049 & ~n25717;
  assign n25719 = ~P1_INSTADDRPOINTER_REG_29__SCAN_IN & ~n43027;
  assign n25721 = P1_INSTADDRPOINTER_REG_31__SCAN_IN & n25720;
  assign n25848 = ~n31032 | ~n25721;
  assign n25723 = ~n25731 | ~P1_EBX_REG_1__SCAN_IN;
  assign n25724 = ~n25723 | ~n25722;
  assign n25728 = ~n25724 ^ n27579;
  assign n25727 = n27579 | P1_EBX_REG_0__SCAN_IN;
  assign n25725 = n26986 & P1_EBX_REG_0__SCAN_IN;
  assign n25726 = ~n25725 | ~n43131;
  assign n42486 = ~n25727 | ~n25726;
  assign n25729 = ~n25728 | ~n42486;
  assign n42439 = ~n42464 | ~n25730;
  assign n42485 = n25731;
  assign n25733 = ~n42485 | ~P1_EBX_REG_2__SCAN_IN;
  assign n25732 = ~n42461 | ~P1_INSTADDRPOINTER_REG_2__SCAN_IN;
  assign n25734 = ~n25733 | ~n25732;
  assign n42438 = ~n25734 ^ n25822;
  assign n25736 = ~n42485 | ~P1_EBX_REG_3__SCAN_IN;
  assign n25735 = ~n42461 | ~P1_INSTADDRPOINTER_REG_3__SCAN_IN;
  assign n25737 = ~n25736 | ~n25735;
  assign n42420 = ~n25737 ^ n27579;
  assign n42384 = ~n42421 | ~n42420;
  assign n25739 = ~n42485 | ~P1_EBX_REG_4__SCAN_IN;
  assign n25738 = ~n42461 | ~P1_INSTADDRPOINTER_REG_4__SCAN_IN;
  assign n25740 = ~n25739 | ~n25738;
  assign n42385 = ~n25740 ^ n25822;
  assign n25743 = ~n42485 | ~P1_EBX_REG_5__SCAN_IN;
  assign n25742 = ~n42461 | ~P1_INSTADDRPOINTER_REG_5__SCAN_IN;
  assign n25744 = ~n25743 | ~n25742;
  assign n31401 = ~n25744 ^ n25822;
  assign n25746 = ~n42485 | ~P1_EBX_REG_6__SCAN_IN;
  assign n25745 = ~n42461 | ~P1_INSTADDRPOINTER_REG_6__SCAN_IN;
  assign n25747 = ~n25746 | ~n25745;
  assign n25749 = ~n42485 | ~P1_EBX_REG_7__SCAN_IN;
  assign n25748 = ~n42461 | ~P1_INSTADDRPOINTER_REG_7__SCAN_IN;
  assign n25750 = ~n25749 | ~n25748;
  assign n31367 = ~n25750 ^ n27579;
  assign n25752 = ~n42485 | ~P1_EBX_REG_8__SCAN_IN;
  assign n25751 = ~n42461 | ~P1_INSTADDRPOINTER_REG_8__SCAN_IN;
  assign n25753 = ~n25752 | ~n25751;
  assign n31352 = ~n25753 ^ n25822;
  assign n25755 = ~n42485 | ~P1_EBX_REG_9__SCAN_IN;
  assign n25754 = ~n42461 | ~P1_INSTADDRPOINTER_REG_9__SCAN_IN;
  assign n25756 = ~n25755 | ~n25754;
  assign n31338 = ~n25756 ^ n25822;
  assign n25758 = ~n42485 | ~P1_EBX_REG_10__SCAN_IN;
  assign n25757 = ~n42461 | ~P1_INSTADDRPOINTER_REG_10__SCAN_IN;
  assign n25759 = ~n25758 | ~n25757;
  assign n30330 = ~n25759 ^ n27579;
  assign n25761 = ~n42485 | ~P1_EBX_REG_11__SCAN_IN;
  assign n25760 = ~n42461 | ~P1_INSTADDRPOINTER_REG_11__SCAN_IN;
  assign n25762 = ~n25761 | ~n25760;
  assign n30314 = ~n25762 ^ n27579;
  assign n25764 = ~n42485 | ~P1_EBX_REG_12__SCAN_IN;
  assign n25763 = ~n42461 | ~P1_INSTADDRPOINTER_REG_12__SCAN_IN;
  assign n25765 = ~n25764 | ~n25763;
  assign n30291 = ~n25765 ^ n25822;
  assign n25767 = ~n42485 | ~P1_EBX_REG_13__SCAN_IN;
  assign n25766 = ~n42461 | ~P1_INSTADDRPOINTER_REG_13__SCAN_IN;
  assign n25768 = ~n25767 | ~n25766;
  assign n30267 = ~n25768 ^ n25822;
  assign n25770 = ~n42485 | ~P1_EBX_REG_14__SCAN_IN;
  assign n25769 = ~n42461 | ~P1_INSTADDRPOINTER_REG_14__SCAN_IN;
  assign n25771 = ~n25770 | ~n25769;
  assign n30243 = ~n25771 ^ n25822;
  assign n25773 = ~n42485 | ~P1_EBX_REG_15__SCAN_IN;
  assign n25772 = ~n42461 | ~P1_INSTADDRPOINTER_REG_15__SCAN_IN;
  assign n25774 = ~n25773 | ~n25772;
  assign n30226 = ~n25774 ^ n27579;
  assign n25779 = ~n30228;
  assign n25776 = ~n42485 | ~P1_EBX_REG_16__SCAN_IN;
  assign n25775 = ~n42461 | ~P1_INSTADDRPOINTER_REG_16__SCAN_IN;
  assign n25777 = ~n25776 | ~n25775;
  assign n30199 = ~n25777 ^ n25822;
  assign n30182 = ~n25779 | ~n25778;
  assign n25781 = ~n42485 | ~P1_EBX_REG_17__SCAN_IN;
  assign n25780 = ~n42461 | ~P1_INSTADDRPOINTER_REG_17__SCAN_IN;
  assign n25782 = ~n25781 | ~n25780;
  assign n30181 = ~n25782 ^ n25822;
  assign n25784 = ~n42485 | ~P1_EBX_REG_18__SCAN_IN;
  assign n25783 = ~n42461 | ~P1_INSTADDRPOINTER_REG_18__SCAN_IN;
  assign n25785 = ~n25784 | ~n25783;
  assign n30156 = ~n25785 ^ n27579;
  assign n25787 = ~n42485 | ~P1_EBX_REG_19__SCAN_IN;
  assign n25786 = ~n42461 | ~P1_INSTADDRPOINTER_REG_19__SCAN_IN;
  assign n25788 = ~n25787 | ~n25786;
  assign n30138 = ~n25788 ^ n25822;
  assign n25792 = ~n42485 | ~P1_EBX_REG_20__SCAN_IN;
  assign n25791 = ~n42461 | ~P1_INSTADDRPOINTER_REG_20__SCAN_IN;
  assign n25793 = ~n25792 | ~n25791;
  assign n27082 = ~n25793 ^ n25822;
  assign n25795 = ~n42485 | ~P1_EBX_REG_21__SCAN_IN;
  assign n25794 = ~n42461 | ~P1_INSTADDRPOINTER_REG_21__SCAN_IN;
  assign n25796 = ~n25795 | ~n25794;
  assign n27104 = ~n25796 ^ n27579;
  assign n25798 = ~n42485 | ~P1_EBX_REG_22__SCAN_IN;
  assign n25797 = ~n42461 | ~P1_INSTADDRPOINTER_REG_22__SCAN_IN;
  assign n25799 = ~n25798 | ~n25797;
  assign n30083 = ~n25799 ^ n27579;
  assign n25801 = ~n42485 | ~P1_EBX_REG_23__SCAN_IN;
  assign n25800 = ~n42461 | ~P1_INSTADDRPOINTER_REG_23__SCAN_IN;
  assign n25802 = ~n25801 | ~n25800;
  assign n30055 = ~n25802 ^ n25822;
  assign n25806 = ~n42485 | ~P1_EBX_REG_24__SCAN_IN;
  assign n25805 = ~n42461 | ~P1_INSTADDRPOINTER_REG_24__SCAN_IN;
  assign n25807 = ~n25806 | ~n25805;
  assign n30033 = ~n25807 ^ n25822;
  assign n25809 = ~n42485 | ~P1_EBX_REG_25__SCAN_IN;
  assign n25808 = ~n42461 | ~P1_INSTADDRPOINTER_REG_25__SCAN_IN;
  assign n25810 = ~n25809 | ~n25808;
  assign n30014 = ~n25810 ^ n27579;
  assign n25812 = ~n42485 | ~P1_EBX_REG_26__SCAN_IN;
  assign n25811 = ~n42461 | ~P1_INSTADDRPOINTER_REG_26__SCAN_IN;
  assign n25813 = ~n25812 | ~n25811;
  assign n29994 = ~n25813 ^ n27579;
  assign n25815 = ~n42485 | ~P1_EBX_REG_27__SCAN_IN;
  assign n25814 = ~n42461 | ~P1_INSTADDRPOINTER_REG_27__SCAN_IN;
  assign n25816 = ~n25815 | ~n25814;
  assign n29972 = ~n25816 ^ n25822;
  assign n25818 = ~n42485 | ~P1_EBX_REG_28__SCAN_IN;
  assign n25817 = ~n42461 | ~P1_INSTADDRPOINTER_REG_28__SCAN_IN;
  assign n25819 = ~n25818 | ~n25817;
  assign n29950 = ~n25819 ^ n25822;
  assign n25821 = ~n42485 | ~P1_EBX_REG_29__SCAN_IN;
  assign n25820 = ~n42461 | ~P1_INSTADDRPOINTER_REG_29__SCAN_IN;
  assign n29911 = ~n25821 | ~n25820;
  assign n29936 = ~n29911 ^ n27579;
  assign n29913 = ~n25823 | ~n25822;
  assign n25825 = ~n42485 | ~P1_EBX_REG_30__SCAN_IN;
  assign n25824 = ~n42461 | ~P1_INSTADDRPOINTER_REG_30__SCAN_IN;
  assign n29914 = ~n25825 | ~n25824;
  assign n25826 = n29936 & n29914;
  assign n25827 = ~n29952 | ~n25826;
  assign n25831 = ~n29913 | ~n25827;
  assign n25829 = ~n42485 | ~P1_EBX_REG_31__SCAN_IN;
  assign n25828 = ~n42461 | ~P1_INSTADDRPOINTER_REG_31__SCAN_IN;
  assign n25830 = n25829 & n25828;
  assign n42503 = ~n25831 ^ n25830;
  assign n25835 = ~n25833 & ~n25832;
  assign n25834 = ~n31439 & ~n44843;
  assign n25836 = ~n25835 & ~n25834;
  assign n25847 = ~n42503 | ~n25838;
  assign n43026 = ~P1_INSTADDRPOINTER_REG_0__SCAN_IN & ~n43031;
  assign n31102 = ~n25839 | ~n31230;
  assign n25841 = ~n43014 | ~n25840;
  assign n31119 = ~n31102 | ~n25841;
  assign n31079 = ~n31119 | ~n25842;
  assign n31036 = ~n31049 | ~n31062;
  assign n31031 = ~n31035 & ~n31036;
  assign n25843 = ~P1_INSTADDRPOINTER_REG_31__SCAN_IN;
  assign n25844 = n25843 & P1_INSTADDRPOINTER_REG_30__SCAN_IN;
  assign n25846 = n31031 & n25844;
  assign n30637 = ~n42929 | ~P1_REIP_REG_31__SCAN_IN;
  assign n25845 = ~n30637;
  assign n25849 = ~n25988;
  assign n25920 = ~n26904;
  assign n25895 = ~n25002 & ~n43082;
  assign n25857 = ~n25895 | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n25851 = ~P1_EAX_REG_2__SCAN_IN;
  assign n25855 = n26391 | n25851;
  assign n25853 = ~n26904 | ~P1_PHYADDRPOINTER_REG_2__SCAN_IN;
  assign n42919 = ~P1_PHYADDRPOINTER_REG_1__SCAN_IN ^ P1_PHYADDRPOINTER_REG_2__SCAN_IN;
  assign n25852 = ~n25877 | ~n42919;
  assign n25854 = n25853 & n25852;
  assign n25856 = n25855 & n25854;
  assign n25881 = n25857 & n25856;
  assign n25860 = ~n25859;
  assign n25867 = ~n43066 | ~n25849;
  assign n25865 = ~n25895 | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign n25861 = ~P1_EAX_REG_1__SCAN_IN;
  assign n25863 = n26391 | n25861;
  assign n25862 = ~n43082 | ~P1_PHYADDRPOINTER_REG_1__SCAN_IN;
  assign n25864 = n25863 & n25862;
  assign n25866 = n25865 & n25864;
  assign n42459 = ~n25867 | ~n25866;
  assign n44801 = n25868;
  assign n25869 = n44801 | n26912;
  assign n25876 = n43379 | n25988;
  assign n25874 = ~n25895 | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN;
  assign n25870 = ~P1_EAX_REG_0__SCAN_IN;
  assign n25872 = n26391 | n25870;
  assign n25871 = ~n43082 | ~P1_PHYADDRPOINTER_REG_0__SCAN_IN;
  assign n25873 = n25872 & n25871;
  assign n25875 = n25874 & n25873;
  assign n42482 = ~n25876 | ~n25875;
  assign n25880 = ~n23975 | ~n42482;
  assign n25878 = ~n42482;
  assign n25879 = ~n25878 | ~n26900;
  assign n42458 = ~n25880 | ~n25879;
  assign n25882 = ~n25881;
  assign n25884 = ~n25883 | ~n25882;
  assign n43072 = n25885;
  assign n25894 = ~n43072 | ~n25849;
  assign n25890 = ~n25895 | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n25886 = ~P1_EAX_REG_3__SCAN_IN;
  assign n25888 = n26391 | n25886;
  assign n25887 = ~n26904 | ~P1_PHYADDRPOINTER_REG_3__SCAN_IN;
  assign n25889 = n25888 & n25887;
  assign n25892 = ~n25890 | ~n25889;
  assign n25903 = ~P1_PHYADDRPOINTER_REG_1__SCAN_IN | ~P1_PHYADDRPOINTER_REG_2__SCAN_IN;
  assign n42906 = n25902 ^ n25903;
  assign n25891 = ~n42906 & ~n26894;
  assign n25893 = ~n25892 & ~n25891;
  assign n42431 = ~n25894 | ~n25893;
  assign n25901 = ~n25895 | ~P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN;
  assign n25896 = ~P1_EAX_REG_4__SCAN_IN;
  assign n25899 = n26391 | n25896;
  assign n25897 = ~n43082 | ~P1_PHYADDRPOINTER_REG_4__SCAN_IN;
  assign n25898 = n26894 & n25897;
  assign n25900 = n25899 & n25898;
  assign n25905 = ~n25901 | ~n25900;
  assign n42894 = P1_PHYADDRPOINTER_REG_4__SCAN_IN ^ n25912;
  assign n25904 = ~n42894 | ~n26900;
  assign n25906 = ~n25905 | ~n25904;
  assign n25909 = ~P1_EAX_REG_5__SCAN_IN;
  assign n25911 = n26391 | n25909;
  assign n25910 = n25920 | n31023;
  assign n25914 = ~n25911 | ~n25910;
  assign n25918 = ~n25912 | ~P1_PHYADDRPOINTER_REG_4__SCAN_IN;
  assign n42363 = ~n25918 ^ P1_PHYADDRPOINTER_REG_5__SCAN_IN;
  assign n25913 = ~n42363 & ~n26894;
  assign n25915 = ~n25914 & ~n25913;
  assign n25926 = ~n25916 | ~n25849;
  assign n25917 = ~P1_EAX_REG_6__SCAN_IN;
  assign n25924 = n26391 | n25917;
  assign n25928 = ~n25918 & ~n31023;
  assign n25919 = ~n25928;
  assign n42350 = ~P1_PHYADDRPOINTER_REG_6__SCAN_IN ^ n25919;
  assign n25922 = n42350 | n26894;
  assign n25921 = ~n26904 | ~P1_PHYADDRPOINTER_REG_6__SCAN_IN;
  assign n25923 = n25922 & n25921;
  assign n25925 = n25924 & n25923;
  assign n30999 = ~n25926 | ~n25925;
  assign n25935 = ~n22940 | ~n25849;
  assign n25927 = ~P1_EAX_REG_7__SCAN_IN;
  assign n25933 = n26391 | n25927;
  assign n25938 = ~n25928 | ~P1_PHYADDRPOINTER_REG_6__SCAN_IN;
  assign n25929 = ~n25938;
  assign n42327 = ~P1_PHYADDRPOINTER_REG_7__SCAN_IN ^ n25929;
  assign n25931 = ~n42327 | ~n25877;
  assign n25930 = ~n26904 | ~P1_PHYADDRPOINTER_REG_7__SCAN_IN;
  assign n25932 = n25931 & n25930;
  assign n25934 = n25933 & n25932;
  assign n25945 = n25936 | n25988;
  assign n25937 = ~P1_EAX_REG_8__SCAN_IN;
  assign n25943 = n26391 | n25937;
  assign n25939 = ~n25980;
  assign n42306 = ~P1_PHYADDRPOINTER_REG_8__SCAN_IN ^ n25939;
  assign n25941 = n42306 | n26894;
  assign n25940 = ~n26904 | ~P1_PHYADDRPOINTER_REG_8__SCAN_IN;
  assign n25942 = n25941 & n25940;
  assign n25944 = n25943 & n25942;
  assign n25948 = ~n26707 | ~P1_INSTQUEUE_REG_12__1__SCAN_IN;
  assign n25947 = ~n26630 | ~P1_INSTQUEUE_REG_10__1__SCAN_IN;
  assign n25952 = ~n25948 | ~n25947;
  assign n25950 = ~n26875 | ~P1_INSTQUEUE_REG_15__1__SCAN_IN;
  assign n25949 = ~n26879 | ~P1_INSTQUEUE_REG_13__1__SCAN_IN;
  assign n25951 = ~n25950 | ~n25949;
  assign n25960 = ~n25952 & ~n25951;
  assign n25954 = ~n26858 | ~P1_INSTQUEUE_REG_6__1__SCAN_IN;
  assign n25953 = ~n26817 | ~P1_INSTQUEUE_REG_4__1__SCAN_IN;
  assign n25958 = ~n25954 | ~n25953;
  assign n25956 = ~n25147 | ~P1_INSTQUEUE_REG_7__1__SCAN_IN;
  assign n25955 = ~n26869 | ~P1_INSTQUEUE_REG_3__1__SCAN_IN;
  assign n25957 = ~n25956 | ~n25955;
  assign n25959 = ~n25958 & ~n25957;
  assign n25977 = ~n25960 | ~n25959;
  assign n25962 = ~n26577 | ~P1_INSTQUEUE_REG_2__1__SCAN_IN;
  assign n25961 = ~n26818 | ~P1_INSTQUEUE_REG_14__1__SCAN_IN;
  assign n25964 = ~n25962 | ~n25961;
  assign n26481 = ~P1_INSTQUEUE_REG_1__1__SCAN_IN;
  assign n25963 = ~n31463 & ~n26481;
  assign n25967 = ~n25964 & ~n25963;
  assign n25965 = ~P1_INSTQUEUE_REG_8__1__SCAN_IN;
  assign n25966 = n22833 | n25965;
  assign n25975 = n25967 & n25966;
  assign n25969 = ~n26753 | ~P1_INSTQUEUE_REG_9__1__SCAN_IN;
  assign n25968 = ~n26870 | ~P1_INSTQUEUE_REG_0__1__SCAN_IN;
  assign n25973 = ~n25969 | ~n25968;
  assign n25971 = ~n26622 | ~P1_INSTQUEUE_REG_11__1__SCAN_IN;
  assign n25970 = ~n26859 | ~P1_INSTQUEUE_REG_5__1__SCAN_IN;
  assign n25972 = ~n25971 | ~n25970;
  assign n25974 = ~n25973 & ~n25972;
  assign n25976 = ~n25975 | ~n25974;
  assign n25978 = ~n25977 & ~n25976;
  assign n25987 = n25988 | n25978;
  assign n25979 = ~P1_EAX_REG_9__SCAN_IN;
  assign n25985 = n26391 | n25979;
  assign n25991 = ~n25980 | ~P1_PHYADDRPOINTER_REG_8__SCAN_IN;
  assign n25981 = ~n25991;
  assign n42290 = ~P1_PHYADDRPOINTER_REG_9__SCAN_IN ^ n25981;
  assign n25983 = ~n42290 | ~n25877;
  assign n25982 = ~n26904 | ~P1_PHYADDRPOINTER_REG_9__SCAN_IN;
  assign n25984 = n25983 & n25982;
  assign n25986 = n25985 & n25984;
  assign n30956 = n25987 & n25986;
  assign n25989 = ~P1_EAX_REG_10__SCAN_IN;
  assign n25995 = n26391 | n25989;
  assign n25993 = ~n26904 | ~P1_PHYADDRPOINTER_REG_10__SCAN_IN;
  assign n30937 = ~P1_PHYADDRPOINTER_REG_10__SCAN_IN ^ n26031;
  assign n25992 = ~n30937 | ~n25877;
  assign n25994 = n25993 & n25992;
  assign n25996 = n25995 & n25994;
  assign n30323 = ~n25997 | ~n25996;
  assign n25999 = ~n26847 | ~P1_INSTQUEUE_REG_8__4__SCAN_IN;
  assign n25998 = ~n26870 | ~P1_INSTQUEUE_REG_0__4__SCAN_IN;
  assign n26003 = ~n25999 | ~n25998;
  assign n26001 = ~n26753 | ~P1_INSTQUEUE_REG_9__4__SCAN_IN;
  assign n26000 = ~n22842 | ~P1_INSTQUEUE_REG_1__4__SCAN_IN;
  assign n26002 = ~n26001 | ~n26000;
  assign n26011 = ~n26003 & ~n26002;
  assign n26005 = ~n26858 | ~P1_INSTQUEUE_REG_6__4__SCAN_IN;
  assign n26004 = ~n26818 | ~P1_INSTQUEUE_REG_14__4__SCAN_IN;
  assign n26009 = ~n26005 | ~n26004;
  assign n26007 = ~n25147 | ~P1_INSTQUEUE_REG_7__4__SCAN_IN;
  assign n26006 = ~n26630 | ~P1_INSTQUEUE_REG_10__4__SCAN_IN;
  assign n26008 = ~n26007 | ~n26006;
  assign n26010 = ~n26009 & ~n26008;
  assign n26027 = ~n26011 | ~n26010;
  assign n26013 = ~n26875 | ~P1_INSTQUEUE_REG_15__4__SCAN_IN;
  assign n26012 = ~n26859 | ~P1_INSTQUEUE_REG_5__4__SCAN_IN;
  assign n26017 = ~n26013 | ~n26012;
  assign n26015 = ~n26622 | ~P1_INSTQUEUE_REG_11__4__SCAN_IN;
  assign n26014 = ~n26869 | ~P1_INSTQUEUE_REG_3__4__SCAN_IN;
  assign n26016 = ~n26015 | ~n26014;
  assign n26025 = ~n26017 & ~n26016;
  assign n26019 = ~n26707 | ~P1_INSTQUEUE_REG_12__4__SCAN_IN;
  assign n26018 = ~n26817 | ~P1_INSTQUEUE_REG_4__4__SCAN_IN;
  assign n26023 = ~n26019 | ~n26018;
  assign n26021 = ~n26879 | ~P1_INSTQUEUE_REG_13__4__SCAN_IN;
  assign n26020 = ~n26577 | ~P1_INSTQUEUE_REG_2__4__SCAN_IN;
  assign n26022 = ~n26021 | ~n26020;
  assign n26024 = ~n26023 & ~n26022;
  assign n26026 = ~n26025 | ~n26024;
  assign n26028 = ~n26027 & ~n26026;
  assign n26030 = n25988 | n26028;
  assign n26029 = ~n26904 | ~P1_PHYADDRPOINTER_REG_12__SCAN_IN;
  assign n26066 = ~n26031 | ~P1_PHYADDRPOINTER_REG_10__SCAN_IN;
  assign n30911 = ~n26072 ^ P1_PHYADDRPOINTER_REG_12__SCAN_IN;
  assign n26033 = ~n30911 | ~n25877;
  assign n42872 = ~P1_EAX_REG_12__SCAN_IN;
  assign n26032 = n26391 | n42872;
  assign n26034 = ~n26033 | ~n26032;
  assign n26037 = ~n25147 | ~P1_INSTQUEUE_REG_7__3__SCAN_IN;
  assign n26036 = ~n26866 | ~P1_INSTQUEUE_REG_10__3__SCAN_IN;
  assign n26041 = ~n26037 | ~n26036;
  assign n26039 = ~n22841 | ~P1_INSTQUEUE_REG_3__3__SCAN_IN;
  assign n26038 = ~n26870 | ~P1_INSTQUEUE_REG_0__3__SCAN_IN;
  assign n26040 = ~n26039 | ~n26038;
  assign n26049 = ~n26041 & ~n26040;
  assign n26043 = ~n26875 | ~P1_INSTQUEUE_REG_15__3__SCAN_IN;
  assign n26042 = ~n26859 | ~P1_INSTQUEUE_REG_5__3__SCAN_IN;
  assign n26047 = ~n26043 | ~n26042;
  assign n26045 = ~n26817 | ~P1_INSTQUEUE_REG_4__3__SCAN_IN;
  assign n26044 = ~n26818 | ~P1_INSTQUEUE_REG_14__3__SCAN_IN;
  assign n26046 = ~n26045 | ~n26044;
  assign n26048 = ~n26047 & ~n26046;
  assign n26051 = ~n26622 | ~P1_INSTQUEUE_REG_11__3__SCAN_IN;
  assign n26050 = ~n26879 | ~P1_INSTQUEUE_REG_13__3__SCAN_IN;
  assign n26055 = ~n26051 | ~n26050;
  assign n26053 = ~n26858 | ~P1_INSTQUEUE_REG_6__3__SCAN_IN;
  assign n26052 = ~n26577 | ~P1_INSTQUEUE_REG_2__3__SCAN_IN;
  assign n26054 = ~n26053 | ~n26052;
  assign n26063 = ~n26055 & ~n26054;
  assign n26057 = ~n26847 | ~P1_INSTQUEUE_REG_8__3__SCAN_IN;
  assign n26056 = ~n26707 | ~P1_INSTQUEUE_REG_12__3__SCAN_IN;
  assign n26061 = ~n26057 | ~n26056;
  assign n26059 = ~n26753 | ~P1_INSTQUEUE_REG_9__3__SCAN_IN;
  assign n26058 = ~n22842 | ~P1_INSTQUEUE_REG_1__3__SCAN_IN;
  assign n26060 = ~n26059 | ~n26058;
  assign n26062 = ~n26061 & ~n26060;
  assign n26064 = ~n26063 | ~n26062;
  assign n26065 = n23966 | n26064;
  assign n30304 = ~n26065 | ~n25849;
  assign n30921 = n30307 ^ n26066;
  assign n26071 = ~n30921 & ~n26894;
  assign n26067 = ~P1_EAX_REG_11__SCAN_IN;
  assign n26069 = n26391 | n26067;
  assign n26068 = ~n26904 | ~P1_PHYADDRPOINTER_REG_11__SCAN_IN;
  assign n26070 = ~n26069 | ~n26068;
  assign n30258 = ~n26071 & ~n26070;
  assign n26110 = ~n30304 | ~n30258;
  assign n26113 = ~n26072 | ~P1_PHYADDRPOINTER_REG_12__SCAN_IN;
  assign n30893 = n30891 ^ n26113;
  assign n26109 = ~n30893 & ~n26894;
  assign n26074 = ~n26707 | ~P1_INSTQUEUE_REG_12__5__SCAN_IN;
  assign n26073 = ~n26869 | ~P1_INSTQUEUE_REG_3__5__SCAN_IN;
  assign n26078 = ~n26074 | ~n26073;
  assign n26076 = ~n26870 | ~P1_INSTQUEUE_REG_0__5__SCAN_IN;
  assign n26075 = ~n26817 | ~P1_INSTQUEUE_REG_4__5__SCAN_IN;
  assign n26077 = ~n26076 | ~n26075;
  assign n26086 = ~n26078 & ~n26077;
  assign n26080 = ~n26622 | ~P1_INSTQUEUE_REG_11__5__SCAN_IN;
  assign n26079 = ~n26630 | ~P1_INSTQUEUE_REG_10__5__SCAN_IN;
  assign n26084 = ~n26080 | ~n26079;
  assign n26082 = ~n25147 | ~P1_INSTQUEUE_REG_7__5__SCAN_IN;
  assign n26081 = ~n26859 | ~P1_INSTQUEUE_REG_5__5__SCAN_IN;
  assign n26083 = ~n26082 | ~n26081;
  assign n26085 = ~n26084 & ~n26083;
  assign n26102 = ~n26086 | ~n26085;
  assign n26088 = ~n26847 | ~P1_INSTQUEUE_REG_8__5__SCAN_IN;
  assign n26087 = ~n22842 | ~P1_INSTQUEUE_REG_1__5__SCAN_IN;
  assign n26092 = ~n26088 | ~n26087;
  assign n26090 = ~n26875 | ~P1_INSTQUEUE_REG_15__5__SCAN_IN;
  assign n26089 = ~n26753 | ~P1_INSTQUEUE_REG_9__5__SCAN_IN;
  assign n26091 = ~n26090 | ~n26089;
  assign n26100 = ~n26092 & ~n26091;
  assign n26094 = ~n26879 | ~P1_INSTQUEUE_REG_13__5__SCAN_IN;
  assign n26093 = ~n26818 | ~P1_INSTQUEUE_REG_14__5__SCAN_IN;
  assign n26098 = ~n26094 | ~n26093;
  assign n26096 = ~n26858 | ~P1_INSTQUEUE_REG_6__5__SCAN_IN;
  assign n26095 = ~n26577 | ~P1_INSTQUEUE_REG_2__5__SCAN_IN;
  assign n26097 = ~n26096 | ~n26095;
  assign n26099 = ~n26098 & ~n26097;
  assign n26101 = ~n26100 | ~n26099;
  assign n26103 = ~n26102 & ~n26101;
  assign n26107 = n25988 | n26103;
  assign n42877 = ~P1_EAX_REG_13__SCAN_IN;
  assign n26105 = n26391 | n42877;
  assign n26104 = ~n26904 | ~P1_PHYADDRPOINTER_REG_13__SCAN_IN;
  assign n26106 = n26105 & n26104;
  assign n26108 = ~n26107 | ~n26106;
  assign n26111 = ~n26110 | ~n23030;
  assign n26112 = ~n30283 & ~n26111;
  assign n30871 = ~n26184 ^ P1_PHYADDRPOINTER_REG_14__SCAN_IN;
  assign n26150 = ~n30871 | ~n25877;
  assign n26115 = ~n26622 | ~P1_INSTQUEUE_REG_11__6__SCAN_IN;
  assign n26114 = ~n26870 | ~P1_INSTQUEUE_REG_0__6__SCAN_IN;
  assign n26119 = ~n26115 | ~n26114;
  assign n26117 = ~n26875 | ~P1_INSTQUEUE_REG_15__6__SCAN_IN;
  assign n26116 = ~n26818 | ~P1_INSTQUEUE_REG_14__6__SCAN_IN;
  assign n26118 = ~n26117 | ~n26116;
  assign n26127 = ~n26119 & ~n26118;
  assign n26121 = ~n25147 | ~P1_INSTQUEUE_REG_7__6__SCAN_IN;
  assign n26120 = ~n26859 | ~P1_INSTQUEUE_REG_5__6__SCAN_IN;
  assign n26125 = ~n26121 | ~n26120;
  assign n26123 = ~n26879 | ~P1_INSTQUEUE_REG_13__6__SCAN_IN;
  assign n26122 = ~n26817 | ~P1_INSTQUEUE_REG_4__6__SCAN_IN;
  assign n26124 = ~n26123 | ~n26122;
  assign n26126 = ~n26125 & ~n26124;
  assign n26143 = ~n26127 | ~n26126;
  assign n26129 = ~n22841 | ~P1_INSTQUEUE_REG_3__6__SCAN_IN;
  assign n26128 = ~n26577 | ~P1_INSTQUEUE_REG_2__6__SCAN_IN;
  assign n26131 = n26129 & n26128;
  assign n26130 = ~n26707 | ~P1_INSTQUEUE_REG_12__6__SCAN_IN;
  assign n26133 = ~n26131 | ~n26130;
  assign n26799 = ~P1_INSTQUEUE_REG_8__6__SCAN_IN;
  assign n26132 = ~n22832 & ~n26799;
  assign n26141 = ~n26133 & ~n26132;
  assign n26135 = ~n26753 | ~P1_INSTQUEUE_REG_9__6__SCAN_IN;
  assign n26134 = ~n26866 | ~P1_INSTQUEUE_REG_10__6__SCAN_IN;
  assign n26139 = ~n26135 | ~n26134;
  assign n26137 = ~n26858 | ~P1_INSTQUEUE_REG_6__6__SCAN_IN;
  assign n26136 = ~n22842 | ~P1_INSTQUEUE_REG_1__6__SCAN_IN;
  assign n26138 = ~n26137 | ~n26136;
  assign n26140 = ~n26139 & ~n26138;
  assign n26142 = ~n26141 | ~n26140;
  assign n26144 = ~n26143 & ~n26142;
  assign n26148 = n25988 | n26144;
  assign n42882 = ~P1_EAX_REG_14__SCAN_IN;
  assign n26146 = n26391 | n42882;
  assign n26145 = ~n26904 | ~P1_PHYADDRPOINTER_REG_14__SCAN_IN;
  assign n26147 = n26146 & n26145;
  assign n26149 = n26148 & n26147;
  assign n30238 = n26150 & n26149;
  assign n26327 = ~P1_INSTQUEUE_REG_8__7__SCAN_IN;
  assign n26158 = ~n22832 & ~n26327;
  assign n26153 = ~n26875 | ~P1_INSTQUEUE_REG_15__7__SCAN_IN;
  assign n26152 = ~n26577 | ~P1_INSTQUEUE_REG_2__7__SCAN_IN;
  assign n26156 = ~n26153 | ~n26152;
  assign n26155 = ~n26360 & ~n26154;
  assign n26157 = n26156 | n26155;
  assign n26166 = ~n26158 & ~n26157;
  assign n26160 = ~n26753 | ~P1_INSTQUEUE_REG_9__7__SCAN_IN;
  assign n26159 = ~n26866 | ~P1_INSTQUEUE_REG_10__7__SCAN_IN;
  assign n26164 = ~n26160 | ~n26159;
  assign n26162 = ~n26707 | ~P1_INSTQUEUE_REG_12__7__SCAN_IN;
  assign n26161 = ~n26870 | ~P1_INSTQUEUE_REG_0__7__SCAN_IN;
  assign n26163 = ~n26162 | ~n26161;
  assign n26165 = ~n26164 & ~n26163;
  assign n26182 = ~n26166 | ~n26165;
  assign n26168 = ~n26869 | ~P1_INSTQUEUE_REG_3__7__SCAN_IN;
  assign n26167 = ~n26858 | ~P1_INSTQUEUE_REG_6__7__SCAN_IN;
  assign n26172 = ~n26168 | ~n26167;
  assign n26170 = ~n24947 | ~P1_INSTQUEUE_REG_11__7__SCAN_IN;
  assign n26169 = ~n22842 | ~P1_INSTQUEUE_REG_1__7__SCAN_IN;
  assign n26171 = ~n26170 | ~n26169;
  assign n26180 = ~n26172 & ~n26171;
  assign n26174 = ~n26879 | ~P1_INSTQUEUE_REG_13__7__SCAN_IN;
  assign n26173 = ~n26859 | ~P1_INSTQUEUE_REG_5__7__SCAN_IN;
  assign n26178 = ~n26174 | ~n26173;
  assign n26176 = ~n26817 | ~P1_INSTQUEUE_REG_4__7__SCAN_IN;
  assign n26175 = ~n26818 | ~P1_INSTQUEUE_REG_14__7__SCAN_IN;
  assign n26177 = ~n26176 | ~n26175;
  assign n26179 = ~n26178 & ~n26177;
  assign n26181 = ~n26180 | ~n26179;
  assign n26183 = ~n26182 & ~n26181;
  assign n26191 = n25988 | n26183;
  assign n30606 = ~P1_EAX_REG_15__SCAN_IN;
  assign n26189 = n26391 | n30606;
  assign n26231 = ~n26184 | ~P1_PHYADDRPOINTER_REG_14__SCAN_IN;
  assign n26185 = ~n26231;
  assign n30858 = ~P1_PHYADDRPOINTER_REG_15__SCAN_IN ^ n26185;
  assign n26187 = ~n30858 | ~n26900;
  assign n26186 = ~n26904 | ~P1_PHYADDRPOINTER_REG_15__SCAN_IN;
  assign n26188 = n26187 & n26186;
  assign n26190 = n26189 & n26188;
  assign n26195 = ~n25147 | ~P1_INSTQUEUE_REG_8__0__SCAN_IN;
  assign n26194 = ~n26859 | ~P1_INSTQUEUE_REG_6__0__SCAN_IN;
  assign n26199 = ~n26195 | ~n26194;
  assign n26197 = ~n26707 | ~P1_INSTQUEUE_REG_13__0__SCAN_IN;
  assign n26196 = ~n26817 | ~P1_INSTQUEUE_REG_5__0__SCAN_IN;
  assign n26198 = ~n26197 | ~n26196;
  assign n26207 = ~n26199 & ~n26198;
  assign n26201 = ~n26753 | ~P1_INSTQUEUE_REG_10__0__SCAN_IN;
  assign n26200 = ~n26818 | ~P1_INSTQUEUE_REG_15__0__SCAN_IN;
  assign n26205 = ~n26201 | ~n26200;
  assign n26203 = ~n26847 | ~P1_INSTQUEUE_REG_9__0__SCAN_IN;
  assign n26202 = ~n22842 | ~P1_INSTQUEUE_REG_2__0__SCAN_IN;
  assign n26204 = ~n26203 | ~n26202;
  assign n26206 = ~n26205 & ~n26204;
  assign n26223 = ~n26207 | ~n26206;
  assign n26209 = ~n26622 | ~P1_INSTQUEUE_REG_12__0__SCAN_IN;
  assign n26208 = ~n26858 | ~P1_INSTQUEUE_REG_7__0__SCAN_IN;
  assign n26213 = ~n26209 | ~n26208;
  assign n26211 = ~n26866 | ~P1_INSTQUEUE_REG_11__0__SCAN_IN;
  assign n26210 = ~n26870 | ~P1_INSTQUEUE_REG_1__0__SCAN_IN;
  assign n26212 = ~n26211 | ~n26210;
  assign n26221 = ~n26213 & ~n26212;
  assign n26215 = ~n26875 | ~P1_INSTQUEUE_REG_0__0__SCAN_IN;
  assign n26214 = ~n26879 | ~P1_INSTQUEUE_REG_14__0__SCAN_IN;
  assign n26219 = ~n26215 | ~n26214;
  assign n26217 = ~n26869 | ~P1_INSTQUEUE_REG_4__0__SCAN_IN;
  assign n26216 = ~n26577 | ~P1_INSTQUEUE_REG_3__0__SCAN_IN;
  assign n26218 = ~n26217 | ~n26216;
  assign n26220 = ~n26219 & ~n26218;
  assign n26222 = ~n26221 | ~n26220;
  assign n26224 = n26223 | n26222;
  assign n26230 = ~n26890 | ~n26224;
  assign n26225 = ~P1_EAX_REG_16__SCAN_IN;
  assign n26228 = n26391 | n26225;
  assign n26226 = ~n43082 | ~P1_PHYADDRPOINTER_REG_16__SCAN_IN;
  assign n26227 = n26894 & n26226;
  assign n26229 = n26228 & n26227;
  assign n26234 = ~n26230 | ~n26229;
  assign n26232 = ~n26267;
  assign n30839 = ~P1_PHYADDRPOINTER_REG_16__SCAN_IN ^ n26232;
  assign n26233 = ~n30839 | ~n26900;
  assign n30196 = ~n26234 | ~n26233;
  assign n26236 = ~n26859 | ~P1_INSTQUEUE_REG_6__1__SCAN_IN;
  assign n26235 = ~n26818 | ~P1_INSTQUEUE_REG_15__1__SCAN_IN;
  assign n26240 = ~n26236 | ~n26235;
  assign n26238 = ~n26707 | ~P1_INSTQUEUE_REG_13__1__SCAN_IN;
  assign n26237 = ~n26630 | ~P1_INSTQUEUE_REG_11__1__SCAN_IN;
  assign n26239 = ~n26238 | ~n26237;
  assign n26248 = ~n26240 & ~n26239;
  assign n26242 = ~n26847 | ~P1_INSTQUEUE_REG_9__1__SCAN_IN;
  assign n26246 = ~n26242 | ~n26241;
  assign n26244 = ~n26753 | ~P1_INSTQUEUE_REG_10__1__SCAN_IN;
  assign n26243 = ~n22842 | ~P1_INSTQUEUE_REG_2__1__SCAN_IN;
  assign n26245 = ~n26244 | ~n26243;
  assign n26247 = ~n26246 & ~n26245;
  assign n26264 = ~n26248 | ~n26247;
  assign n26250 = ~n25147 | ~P1_INSTQUEUE_REG_8__1__SCAN_IN;
  assign n26249 = ~n26870 | ~P1_INSTQUEUE_REG_1__1__SCAN_IN;
  assign n26254 = ~n26250 | ~n26249;
  assign n26252 = ~n26869 | ~P1_INSTQUEUE_REG_4__1__SCAN_IN;
  assign n26251 = ~n26817 | ~P1_INSTQUEUE_REG_5__1__SCAN_IN;
  assign n26253 = ~n26252 | ~n26251;
  assign n26262 = ~n26254 & ~n26253;
  assign n26256 = ~n26875 | ~P1_INSTQUEUE_REG_0__1__SCAN_IN;
  assign n26255 = ~n26879 | ~P1_INSTQUEUE_REG_14__1__SCAN_IN;
  assign n26260 = ~n26256 | ~n26255;
  assign n26258 = ~n26858 | ~P1_INSTQUEUE_REG_7__1__SCAN_IN;
  assign n26257 = ~n26577 | ~P1_INSTQUEUE_REG_3__1__SCAN_IN;
  assign n26259 = ~n26258 | ~n26257;
  assign n26261 = ~n26260 & ~n26259;
  assign n26263 = ~n26262 | ~n26261;
  assign n26265 = n26264 | n26263;
  assign n26274 = ~n26890 | ~n26265;
  assign n26266 = ~P1_EAX_REG_17__SCAN_IN;
  assign n26268 = ~n26275;
  assign n30815 = ~P1_PHYADDRPOINTER_REG_17__SCAN_IN ^ n26268;
  assign n26270 = ~n30815 | ~n26900;
  assign n26269 = ~n26904 | ~P1_PHYADDRPOINTER_REG_17__SCAN_IN;
  assign n26271 = n26270 & n26269;
  assign n30172 = ~n26274 | ~n26273;
  assign n30807 = P1_PHYADDRPOINTER_REG_18__SCAN_IN ^ n26318;
  assign n26316 = ~n30807 | ~n25877;
  assign n26277 = ~n26707 | ~P1_INSTQUEUE_REG_13__2__SCAN_IN;
  assign n26276 = ~n26817 | ~P1_INSTQUEUE_REG_5__2__SCAN_IN;
  assign n26281 = ~n26277 | ~n26276;
  assign n26279 = ~n26622 | ~P1_INSTQUEUE_REG_12__2__SCAN_IN;
  assign n26278 = ~n26875 | ~P1_INSTQUEUE_REG_0__2__SCAN_IN;
  assign n26280 = ~n26279 | ~n26278;
  assign n26289 = ~n26281 & ~n26280;
  assign n26283 = ~n25147 | ~P1_INSTQUEUE_REG_8__2__SCAN_IN;
  assign n26282 = ~n26630 | ~P1_INSTQUEUE_REG_11__2__SCAN_IN;
  assign n26287 = ~n26283 | ~n26282;
  assign n26285 = ~n26858 | ~P1_INSTQUEUE_REG_7__2__SCAN_IN;
  assign n26284 = ~n26876 | ~P1_INSTQUEUE_REG_3__2__SCAN_IN;
  assign n26286 = ~n26285 | ~n26284;
  assign n26288 = ~n26287 & ~n26286;
  assign n26307 = n26289 & n26288;
  assign n26291 = ~n26859 | ~P1_INSTQUEUE_REG_6__2__SCAN_IN;
  assign n26290 = ~n26818 | ~P1_INSTQUEUE_REG_15__2__SCAN_IN;
  assign n26294 = ~n26291 | ~n26290;
  assign n26292 = ~P1_INSTQUEUE_REG_2__2__SCAN_IN;
  assign n26293 = ~n31463 & ~n26292;
  assign n26297 = ~n26294 & ~n26293;
  assign n26295 = ~P1_INSTQUEUE_REG_9__2__SCAN_IN;
  assign n26296 = n22833 | n26295;
  assign n26305 = ~n26297 | ~n26296;
  assign n26299 = ~n26879 | ~P1_INSTQUEUE_REG_14__2__SCAN_IN;
  assign n26298 = ~n26869 | ~P1_INSTQUEUE_REG_4__2__SCAN_IN;
  assign n26303 = ~n26299 | ~n26298;
  assign n26301 = ~n26753 | ~P1_INSTQUEUE_REG_10__2__SCAN_IN;
  assign n26300 = ~n26870 | ~P1_INSTQUEUE_REG_1__2__SCAN_IN;
  assign n26302 = ~n26301 | ~n26300;
  assign n26304 = n26303 | n26302;
  assign n26306 = ~n26305 & ~n26304;
  assign n26308 = ~n26307 | ~n26306;
  assign n26314 = ~n26890 | ~n26308;
  assign n26309 = ~P1_EAX_REG_18__SCAN_IN;
  assign n26312 = n26391 | n26309;
  assign n26310 = ~n43082 | ~P1_PHYADDRPOINTER_REG_18__SCAN_IN;
  assign n26311 = n26894 & n26310;
  assign n26313 = n26312 & n26311;
  assign n26315 = ~n26314 | ~n26313;
  assign n30153 = ~n26316 | ~n26315;
  assign n26317 = ~n30153;
  assign n30059 = P1_PHYADDRPOINTER_REG_23__SCAN_IN ^ n26522;
  assign n26398 = ~n30059 & ~n26894;
  assign n26319 = ~P1_INSTQUEUE_REG_13__7__SCAN_IN;
  assign n26324 = ~n26320 & ~n26319;
  assign n26322 = ~n26622 | ~P1_INSTQUEUE_REG_12__7__SCAN_IN;
  assign n26321 = ~n26858 | ~P1_INSTQUEUE_REG_7__7__SCAN_IN;
  assign n26323 = ~n26322 | ~n26321;
  assign n26331 = ~n26324 & ~n26323;
  assign n26325 = ~P1_INSTQUEUE_REG_1__7__SCAN_IN;
  assign n26329 = ~n26326 & ~n26325;
  assign n26328 = ~n26360 & ~n26327;
  assign n26330 = ~n26329 & ~n26328;
  assign n26347 = ~n26331 | ~n26330;
  assign n26333 = ~n26879 | ~P1_INSTQUEUE_REG_14__7__SCAN_IN;
  assign n26332 = ~n26817 | ~P1_INSTQUEUE_REG_5__7__SCAN_IN;
  assign n26337 = ~n26333 | ~n26332;
  assign n26335 = ~n26577 | ~P1_INSTQUEUE_REG_3__7__SCAN_IN;
  assign n26334 = ~n26859 | ~P1_INSTQUEUE_REG_6__7__SCAN_IN;
  assign n26336 = ~n26335 | ~n26334;
  assign n26345 = ~n26337 & ~n26336;
  assign n26339 = ~n26630 | ~P1_INSTQUEUE_REG_11__7__SCAN_IN;
  assign n26338 = ~n22842 | ~P1_INSTQUEUE_REG_2__7__SCAN_IN;
  assign n26343 = ~n26339 | ~n26338;
  assign n26341 = ~n26847 | ~P1_INSTQUEUE_REG_9__7__SCAN_IN;
  assign n26340 = ~n26753 | ~P1_INSTQUEUE_REG_10__7__SCAN_IN;
  assign n26342 = ~n26341 | ~n26340;
  assign n26344 = ~n26343 & ~n26342;
  assign n26346 = ~n26345 | ~n26344;
  assign n26355 = ~n26347 & ~n26346;
  assign n26348 = ~P1_INSTQUEUE_REG_15__7__SCAN_IN;
  assign n26353 = ~n26349 & ~n26348;
  assign n26351 = ~n26875 | ~P1_INSTQUEUE_REG_0__7__SCAN_IN;
  assign n26350 = ~n26869 | ~P1_INSTQUEUE_REG_4__7__SCAN_IN;
  assign n26352 = ~n26351 | ~n26350;
  assign n26354 = ~n26353 & ~n26352;
  assign n26480 = ~n26355 | ~n26354;
  assign n26356 = ~P1_INSTQUEUE_REG_10__0__SCAN_IN;
  assign n26364 = ~n22832 & ~n26356;
  assign n26358 = ~n26875 | ~P1_INSTQUEUE_REG_1__0__SCAN_IN;
  assign n26357 = ~n26577 | ~P1_INSTQUEUE_REG_4__0__SCAN_IN;
  assign n26362 = ~n26358 | ~n26357;
  assign n26359 = ~P1_INSTQUEUE_REG_9__0__SCAN_IN;
  assign n26361 = ~n26360 & ~n26359;
  assign n26363 = n26362 | n26361;
  assign n26372 = ~n26364 & ~n26363;
  assign n26366 = ~n26753 | ~P1_INSTQUEUE_REG_11__0__SCAN_IN;
  assign n26365 = ~n26630 | ~P1_INSTQUEUE_REG_12__0__SCAN_IN;
  assign n26370 = ~n26366 | ~n26365;
  assign n26368 = ~n26707 | ~P1_INSTQUEUE_REG_14__0__SCAN_IN;
  assign n26367 = ~n26870 | ~P1_INSTQUEUE_REG_2__0__SCAN_IN;
  assign n26369 = ~n26368 | ~n26367;
  assign n26371 = ~n26370 & ~n26369;
  assign n26388 = ~n26372 | ~n26371;
  assign n26374 = ~n26869 | ~P1_INSTQUEUE_REG_5__0__SCAN_IN;
  assign n26373 = ~n26858 | ~P1_INSTQUEUE_REG_8__0__SCAN_IN;
  assign n26378 = ~n26374 | ~n26373;
  assign n26376 = ~n26622 | ~P1_INSTQUEUE_REG_13__0__SCAN_IN;
  assign n26375 = ~n22842 | ~P1_INSTQUEUE_REG_3__0__SCAN_IN;
  assign n26377 = ~n26376 | ~n26375;
  assign n26386 = ~n26378 & ~n26377;
  assign n26380 = ~n26879 | ~P1_INSTQUEUE_REG_15__0__SCAN_IN;
  assign n26379 = ~n26859 | ~P1_INSTQUEUE_REG_7__0__SCAN_IN;
  assign n26384 = ~n26380 | ~n26379;
  assign n26382 = ~n26817 | ~P1_INSTQUEUE_REG_6__0__SCAN_IN;
  assign n26381 = ~n26818 | ~P1_INSTQUEUE_REG_0__0__SCAN_IN;
  assign n26383 = ~n26382 | ~n26381;
  assign n26385 = ~n26384 & ~n26383;
  assign n26387 = ~n26386 | ~n26385;
  assign n26479 = n26388 | n26387;
  assign n26390 = ~n26480 ^ n26479;
  assign n26389 = ~n26890;
  assign n26396 = ~n26390 & ~n26389;
  assign n26903 = ~n26391;
  assign n26394 = ~n26903 | ~P1_EAX_REG_23__SCAN_IN;
  assign n26392 = ~n30743 & ~P1_STATE2_REG_2__SCAN_IN;
  assign n26393 = ~n26392 & ~n26900;
  assign n26395 = ~n26394 | ~n26393;
  assign n26397 = ~n26396 & ~n26395;
  assign n30770 = ~n26399 ^ P1_PHYADDRPOINTER_REG_21__SCAN_IN;
  assign n26438 = ~n30770 | ~n25877;
  assign n26401 = ~n26858 | ~P1_INSTQUEUE_REG_7__5__SCAN_IN;
  assign n26400 = ~n26577 | ~P1_INSTQUEUE_REG_3__5__SCAN_IN;
  assign n26405 = ~n26401 | ~n26400;
  assign n26403 = ~n26879 | ~P1_INSTQUEUE_REG_14__5__SCAN_IN;
  assign n26402 = ~n26818 | ~P1_INSTQUEUE_REG_15__5__SCAN_IN;
  assign n26404 = ~n26403 | ~n26402;
  assign n26429 = ~n26405 & ~n26404;
  assign n26407 = ~n25147 | ~P1_INSTQUEUE_REG_8__5__SCAN_IN;
  assign n26406 = ~n26622 | ~P1_INSTQUEUE_REG_12__5__SCAN_IN;
  assign n26411 = ~n26407 | ~n26406;
  assign n26409 = ~n26875 | ~P1_INSTQUEUE_REG_0__5__SCAN_IN;
  assign n26408 = ~n26817 | ~P1_INSTQUEUE_REG_5__5__SCAN_IN;
  assign n26410 = ~n26409 | ~n26408;
  assign n26427 = n26411 | n26410;
  assign n26413 = ~n26707 | ~P1_INSTQUEUE_REG_13__5__SCAN_IN;
  assign n26412 = ~n26870 | ~P1_INSTQUEUE_REG_1__5__SCAN_IN;
  assign n26417 = ~n26413 | ~n26412;
  assign n26415 = ~n26869 | ~P1_INSTQUEUE_REG_4__5__SCAN_IN;
  assign n26414 = ~n26859 | ~P1_INSTQUEUE_REG_6__5__SCAN_IN;
  assign n26416 = ~n26415 | ~n26414;
  assign n26425 = ~n26417 & ~n26416;
  assign n26419 = ~n26753 | ~P1_INSTQUEUE_REG_10__5__SCAN_IN;
  assign n26418 = ~n26866 | ~P1_INSTQUEUE_REG_11__5__SCAN_IN;
  assign n26423 = ~n26419 | ~n26418;
  assign n26421 = ~n26847 | ~P1_INSTQUEUE_REG_9__5__SCAN_IN;
  assign n26420 = ~n22842 | ~P1_INSTQUEUE_REG_2__5__SCAN_IN;
  assign n26422 = ~n26421 | ~n26420;
  assign n26424 = ~n26423 & ~n26422;
  assign n26426 = ~n26425 | ~n26424;
  assign n26428 = ~n26427 & ~n26426;
  assign n26430 = ~n26429 | ~n26428;
  assign n26436 = ~n26890 | ~n26430;
  assign n26431 = ~P1_EAX_REG_21__SCAN_IN;
  assign n26434 = n26391 | n26431;
  assign n26432 = ~P1_PHYADDRPOINTER_REG_21__SCAN_IN & ~n44765;
  assign n26433 = P1_STATE2_REG_2__SCAN_IN | n26432;
  assign n26435 = n26434 & n26433;
  assign n26437 = ~n26436 | ~n26435;
  assign n30795 = ~n26439 ^ n30792;
  assign n26478 = n30795 | n26894;
  assign n26441 = ~n26869 | ~P1_INSTQUEUE_REG_4__3__SCAN_IN;
  assign n26440 = ~n26817 | ~P1_INSTQUEUE_REG_5__3__SCAN_IN;
  assign n26445 = ~n26441 | ~n26440;
  assign n26443 = ~n26875 | ~P1_INSTQUEUE_REG_0__3__SCAN_IN;
  assign n26442 = ~n26577 | ~P1_INSTQUEUE_REG_3__3__SCAN_IN;
  assign n26444 = ~n26443 | ~n26442;
  assign n26449 = n26445 | n26444;
  assign n26447 = ~n26879 | ~P1_INSTQUEUE_REG_14__3__SCAN_IN;
  assign n26446 = ~n26859 | ~P1_INSTQUEUE_REG_6__3__SCAN_IN;
  assign n26448 = ~n26447 | ~n26446;
  assign n26469 = ~n26449 & ~n26448;
  assign n26451 = ~n26707 | ~P1_INSTQUEUE_REG_13__3__SCAN_IN;
  assign n26450 = ~n26866 | ~P1_INSTQUEUE_REG_11__3__SCAN_IN;
  assign n26467 = ~n26451 | ~n26450;
  assign n26453 = ~n25147 | ~P1_INSTQUEUE_REG_8__3__SCAN_IN;
  assign n26452 = ~n26818 | ~P1_INSTQUEUE_REG_15__3__SCAN_IN;
  assign n26457 = ~n26453 | ~n26452;
  assign n26455 = ~n26622 | ~P1_INSTQUEUE_REG_12__3__SCAN_IN;
  assign n26454 = ~n26870 | ~P1_INSTQUEUE_REG_1__3__SCAN_IN;
  assign n26456 = ~n26455 | ~n26454;
  assign n26465 = ~n26457 & ~n26456;
  assign n26459 = ~n26847 | ~P1_INSTQUEUE_REG_9__3__SCAN_IN;
  assign n26458 = ~n22842 | ~P1_INSTQUEUE_REG_2__3__SCAN_IN;
  assign n26463 = ~n26459 | ~n26458;
  assign n26461 = ~n26753 | ~P1_INSTQUEUE_REG_10__3__SCAN_IN;
  assign n26460 = ~n26858 | ~P1_INSTQUEUE_REG_7__3__SCAN_IN;
  assign n26462 = ~n26461 | ~n26460;
  assign n26464 = ~n26463 & ~n26462;
  assign n26466 = ~n26465 | ~n26464;
  assign n26468 = ~n26467 & ~n26466;
  assign n26470 = ~n26469 | ~n26468;
  assign n26476 = ~n26890 | ~n26470;
  assign n26471 = ~P1_EAX_REG_19__SCAN_IN;
  assign n26474 = n26391 | n26471;
  assign n26472 = ~P1_PHYADDRPOINTER_REG_19__SCAN_IN & ~n44765;
  assign n26473 = P1_STATE2_REG_2__SCAN_IN | n26472;
  assign n26475 = n26474 & n26473;
  assign n26477 = ~n26476 | ~n26475;
  assign n30131 = ~n26478 | ~n26477;
  assign n26647 = ~n26480 | ~n26479;
  assign n26485 = ~n26482 & ~n26481;
  assign n26484 = ~n25267 & ~n26483;
  assign n26487 = ~n26485 & ~n26484;
  assign n26486 = ~n25147 | ~P1_INSTQUEUE_REG_9__1__SCAN_IN;
  assign n26490 = ~n26487 | ~n26486;
  assign n26488 = ~P1_INSTQUEUE_REG_10__1__SCAN_IN;
  assign n26489 = ~n22833 & ~n26488;
  assign n26498 = ~n26490 & ~n26489;
  assign n26492 = ~n26753 | ~P1_INSTQUEUE_REG_11__1__SCAN_IN;
  assign n26491 = ~n26818 | ~P1_INSTQUEUE_REG_0__1__SCAN_IN;
  assign n26496 = ~n26492 | ~n26491;
  assign n26494 = ~n26630 | ~P1_INSTQUEUE_REG_12__1__SCAN_IN;
  assign n26493 = ~n22842 | ~P1_INSTQUEUE_REG_3__1__SCAN_IN;
  assign n26495 = ~n26494 | ~n26493;
  assign n26497 = ~n26496 & ~n26495;
  assign n26514 = ~n26498 | ~n26497;
  assign n26500 = ~n26879 | ~P1_INSTQUEUE_REG_15__1__SCAN_IN;
  assign n26499 = ~n26869 | ~P1_INSTQUEUE_REG_5__1__SCAN_IN;
  assign n26504 = ~n26500 | ~n26499;
  assign n26502 = ~n26870 | ~P1_INSTQUEUE_REG_2__1__SCAN_IN;
  assign n26501 = ~n26817 | ~P1_INSTQUEUE_REG_6__1__SCAN_IN;
  assign n26503 = ~n26502 | ~n26501;
  assign n26512 = ~n26504 & ~n26503;
  assign n26506 = ~n26622 | ~P1_INSTQUEUE_REG_13__1__SCAN_IN;
  assign n26505 = ~n26629 | ~P1_INSTQUEUE_REG_14__1__SCAN_IN;
  assign n26510 = ~n26506 | ~n26505;
  assign n26508 = ~n26858 | ~P1_INSTQUEUE_REG_8__1__SCAN_IN;
  assign n26507 = ~n26577 | ~P1_INSTQUEUE_REG_4__1__SCAN_IN;
  assign n26509 = ~n26508 | ~n26507;
  assign n26511 = ~n26510 & ~n26509;
  assign n26513 = ~n26512 | ~n26511;
  assign n26648 = ~n26514 & ~n26513;
  assign n26515 = n26647 ^ n26648;
  assign n26521 = ~n26515 | ~n26890;
  assign n26516 = ~P1_EAX_REG_24__SCAN_IN;
  assign n26519 = ~n26391 & ~n26516;
  assign n26517 = ~n43082 | ~P1_PHYADDRPOINTER_REG_24__SCAN_IN;
  assign n26518 = ~n26894 | ~n26517;
  assign n26520 = ~n26519 & ~n26518;
  assign n26524 = ~n26521 | ~n26520;
  assign n30734 = n26656 ^ P1_PHYADDRPOINTER_REG_24__SCAN_IN;
  assign n26523 = ~n30734 | ~n25877;
  assign n30032 = ~n26524 | ~n26523;
  assign n26525 = ~n30131 & ~n30032;
  assign n26566 = ~n30097 | ~n26525;
  assign n30781 = P1_PHYADDRPOINTER_REG_20__SCAN_IN ^ n26526;
  assign n26565 = ~n30781 | ~n25877;
  assign n26528 = ~n25147 | ~P1_INSTQUEUE_REG_8__4__SCAN_IN;
  assign n26527 = ~n26630 | ~P1_INSTQUEUE_REG_11__4__SCAN_IN;
  assign n26532 = ~n26528 | ~n26527;
  assign n26530 = ~n26869 | ~P1_INSTQUEUE_REG_4__4__SCAN_IN;
  assign n26529 = ~n26817 | ~P1_INSTQUEUE_REG_5__4__SCAN_IN;
  assign n26531 = ~n26530 | ~n26529;
  assign n26540 = ~n26532 & ~n26531;
  assign n26534 = ~n26707 | ~P1_INSTQUEUE_REG_13__4__SCAN_IN;
  assign n26533 = ~n26818 | ~P1_INSTQUEUE_REG_15__4__SCAN_IN;
  assign n26538 = ~n26534 | ~n26533;
  assign n26536 = ~n26577 | ~P1_INSTQUEUE_REG_3__4__SCAN_IN;
  assign n26535 = ~n26859 | ~P1_INSTQUEUE_REG_6__4__SCAN_IN;
  assign n26537 = ~n26536 | ~n26535;
  assign n26539 = ~n26538 & ~n26537;
  assign n26556 = ~n26540 | ~n26539;
  assign n26542 = ~n26879 | ~P1_INSTQUEUE_REG_14__4__SCAN_IN;
  assign n26541 = ~n26870 | ~P1_INSTQUEUE_REG_1__4__SCAN_IN;
  assign n26546 = ~n26542 | ~n26541;
  assign n26544 = ~n26875 | ~P1_INSTQUEUE_REG_0__4__SCAN_IN;
  assign n26543 = ~n26858 | ~P1_INSTQUEUE_REG_7__4__SCAN_IN;
  assign n26545 = ~n26544 | ~n26543;
  assign n26554 = ~n26546 & ~n26545;
  assign n26548 = ~n26753 | ~P1_INSTQUEUE_REG_10__4__SCAN_IN;
  assign n26547 = ~n22842 | ~P1_INSTQUEUE_REG_2__4__SCAN_IN;
  assign n26552 = ~n26548 | ~n26547;
  assign n26550 = ~n26847 | ~P1_INSTQUEUE_REG_9__4__SCAN_IN;
  assign n26549 = ~n24947 | ~P1_INSTQUEUE_REG_12__4__SCAN_IN;
  assign n26551 = ~n26550 | ~n26549;
  assign n26553 = ~n26552 & ~n26551;
  assign n26555 = ~n26554 | ~n26553;
  assign n26557 = n26556 | n26555;
  assign n26563 = ~n26557 | ~n26890;
  assign n26558 = ~P1_EAX_REG_20__SCAN_IN;
  assign n26561 = n26391 | n26558;
  assign n26559 = ~n43082 | ~P1_PHYADDRPOINTER_REG_20__SCAN_IN;
  assign n26560 = n26894 & n26559;
  assign n26562 = n26561 & n26560;
  assign n26564 = ~n26563 | ~n26562;
  assign n30114 = ~n26565 | ~n26564;
  assign n26567 = ~n26566 & ~n30114;
  assign n26609 = ~n30054 | ~n26567;
  assign n30758 = P1_PHYADDRPOINTER_REG_22__SCAN_IN ^ n26568;
  assign n26608 = ~n30758 | ~n26900;
  assign n26570 = ~n26875 | ~P1_INSTQUEUE_REG_0__6__SCAN_IN;
  assign n26569 = ~n26817 | ~P1_INSTQUEUE_REG_5__6__SCAN_IN;
  assign n26574 = ~n26570 | ~n26569;
  assign n26572 = ~n26707 | ~P1_INSTQUEUE_REG_13__6__SCAN_IN;
  assign n26571 = ~n26866 | ~P1_INSTQUEUE_REG_11__6__SCAN_IN;
  assign n26573 = ~n26572 | ~n26571;
  assign n26583 = ~n26574 & ~n26573;
  assign n26576 = ~n26686 | ~P1_INSTQUEUE_REG_7__6__SCAN_IN;
  assign n26575 = ~n26870 | ~P1_INSTQUEUE_REG_1__6__SCAN_IN;
  assign n26581 = ~n26576 | ~n26575;
  assign n26579 = ~n26577 | ~P1_INSTQUEUE_REG_3__6__SCAN_IN;
  assign n26578 = ~n26859 | ~P1_INSTQUEUE_REG_6__6__SCAN_IN;
  assign n26580 = ~n26579 | ~n26578;
  assign n26582 = ~n26581 & ~n26580;
  assign n26599 = ~n26583 | ~n26582;
  assign n26585 = ~n26879 | ~P1_INSTQUEUE_REG_14__6__SCAN_IN;
  assign n26584 = ~n26869 | ~P1_INSTQUEUE_REG_4__6__SCAN_IN;
  assign n26587 = n26585 & n26584;
  assign n26586 = ~n26753 | ~P1_INSTQUEUE_REG_10__6__SCAN_IN;
  assign n26589 = ~n26587 | ~n26586;
  assign n26588 = ~n22832 & ~n23581;
  assign n26597 = ~n26589 & ~n26588;
  assign n26591 = ~n26622 | ~P1_INSTQUEUE_REG_12__6__SCAN_IN;
  assign n26590 = ~n26818 | ~P1_INSTQUEUE_REG_15__6__SCAN_IN;
  assign n26595 = ~n26591 | ~n26590;
  assign n26593 = ~n25147 | ~P1_INSTQUEUE_REG_8__6__SCAN_IN;
  assign n26592 = ~n22842 | ~P1_INSTQUEUE_REG_2__6__SCAN_IN;
  assign n26594 = ~n26593 | ~n26592;
  assign n26596 = ~n26595 & ~n26594;
  assign n26598 = ~n26597 | ~n26596;
  assign n26600 = n26599 | n26598;
  assign n26606 = ~n26890 | ~n26600;
  assign n26601 = ~P1_EAX_REG_22__SCAN_IN;
  assign n26604 = n26391 | n26601;
  assign n26602 = ~n43082 | ~P1_PHYADDRPOINTER_REG_22__SCAN_IN;
  assign n26603 = n26894 & n26602;
  assign n26605 = n26604 & n26603;
  assign n26607 = ~n26606 | ~n26605;
  assign n30074 = ~n26608 | ~n26607;
  assign n26610 = ~n26609 & ~n30074;
  assign n26611 = ~P1_INSTQUEUE_REG_15__2__SCAN_IN;
  assign n26614 = ~n25294 & ~n26611;
  assign n26613 = ~n25267 & ~n26612;
  assign n26616 = ~n26614 & ~n26613;
  assign n26615 = ~n26753 | ~P1_INSTQUEUE_REG_11__2__SCAN_IN;
  assign n26619 = ~n26616 | ~n26615;
  assign n26618 = ~n22832 & ~n26617;
  assign n26628 = ~n26619 & ~n26618;
  assign n26621 = ~n25147 | ~P1_INSTQUEUE_REG_9__2__SCAN_IN;
  assign n26620 = ~n22842 | ~P1_INSTQUEUE_REG_3__2__SCAN_IN;
  assign n26626 = ~n26621 | ~n26620;
  assign n26624 = ~n26622 | ~P1_INSTQUEUE_REG_13__2__SCAN_IN;
  assign n26623 = ~n26858 | ~P1_INSTQUEUE_REG_8__2__SCAN_IN;
  assign n26625 = ~n26624 | ~n26623;
  assign n26627 = ~n26626 & ~n26625;
  assign n26646 = ~n26628 | ~n26627;
  assign n26632 = ~n26629 | ~P1_INSTQUEUE_REG_14__2__SCAN_IN;
  assign n26631 = ~n26630 | ~P1_INSTQUEUE_REG_12__2__SCAN_IN;
  assign n26636 = ~n26632 | ~n26631;
  assign n26634 = ~n26869 | ~P1_INSTQUEUE_REG_5__2__SCAN_IN;
  assign n26633 = ~n26870 | ~P1_INSTQUEUE_REG_2__2__SCAN_IN;
  assign n26635 = ~n26634 | ~n26633;
  assign n26644 = ~n26636 & ~n26635;
  assign n26638 = ~n26875 | ~P1_INSTQUEUE_REG_1__2__SCAN_IN;
  assign n26637 = ~n26577 | ~P1_INSTQUEUE_REG_4__2__SCAN_IN;
  assign n26642 = ~n26638 | ~n26637;
  assign n26640 = ~n26817 | ~P1_INSTQUEUE_REG_6__2__SCAN_IN;
  assign n26639 = ~n26818 | ~P1_INSTQUEUE_REG_0__2__SCAN_IN;
  assign n26641 = ~n26640 | ~n26639;
  assign n26643 = ~n26642 & ~n26641;
  assign n26645 = ~n26644 | ~n26643;
  assign n26663 = ~n26646 & ~n26645;
  assign n26662 = n26648 | n26647;
  assign n26649 = n26663 ^ n26662;
  assign n26655 = ~n26649 | ~n26890;
  assign n26650 = ~P1_EAX_REG_25__SCAN_IN;
  assign n26653 = n26391 | n26650;
  assign n26651 = ~P1_PHYADDRPOINTER_REG_25__SCAN_IN & ~n44765;
  assign n26652 = P1_STATE2_REG_2__SCAN_IN | n26651;
  assign n26654 = n26653 & n26652;
  assign n26659 = ~n26655 | ~n26654;
  assign n26657 = ~n26702;
  assign n30716 = ~P1_PHYADDRPOINTER_REG_25__SCAN_IN ^ n26657;
  assign n26658 = ~n30716 | ~n26900;
  assign n30011 = ~n26659 | ~n26658;
  assign n26705 = n26663 | n26662;
  assign n26665 = ~n26817 | ~P1_INSTQUEUE_REG_6__3__SCAN_IN;
  assign n26664 = ~n26859 | ~P1_INSTQUEUE_REG_7__3__SCAN_IN;
  assign n26669 = ~n26665 | ~n26664;
  assign n26667 = ~n26707 | ~P1_INSTQUEUE_REG_14__3__SCAN_IN;
  assign n26666 = ~n26870 | ~P1_INSTQUEUE_REG_2__3__SCAN_IN;
  assign n26668 = ~n26667 | ~n26666;
  assign n26677 = ~n26669 & ~n26668;
  assign n26671 = ~n26847 | ~P1_INSTQUEUE_REG_10__3__SCAN_IN;
  assign n26670 = ~n26875 | ~P1_INSTQUEUE_REG_1__3__SCAN_IN;
  assign n26675 = ~n26671 | ~n26670;
  assign n26673 = ~n26753 | ~P1_INSTQUEUE_REG_11__3__SCAN_IN;
  assign n26672 = ~n22842 | ~P1_INSTQUEUE_REG_3__3__SCAN_IN;
  assign n26674 = ~n26673 | ~n26672;
  assign n26676 = ~n26675 & ~n26674;
  assign n26694 = ~n26677 | ~n26676;
  assign n26679 = ~n25147 | ~P1_INSTQUEUE_REG_9__3__SCAN_IN;
  assign n26678 = ~n26866 | ~P1_INSTQUEUE_REG_12__3__SCAN_IN;
  assign n26683 = ~n26679 | ~n26678;
  assign n26681 = ~n26622 | ~P1_INSTQUEUE_REG_13__3__SCAN_IN;
  assign n26680 = ~n26869 | ~P1_INSTQUEUE_REG_5__3__SCAN_IN;
  assign n26682 = ~n26681 | ~n26680;
  assign n26692 = ~n26683 & ~n26682;
  assign n26685 = ~n26879 | ~P1_INSTQUEUE_REG_15__3__SCAN_IN;
  assign n26684 = ~n26876 | ~P1_INSTQUEUE_REG_4__3__SCAN_IN;
  assign n26690 = ~n26685 | ~n26684;
  assign n26688 = ~n26686 | ~P1_INSTQUEUE_REG_8__3__SCAN_IN;
  assign n26687 = ~n26818 | ~P1_INSTQUEUE_REG_0__3__SCAN_IN;
  assign n26689 = ~n26688 | ~n26687;
  assign n26691 = ~n26690 & ~n26689;
  assign n26693 = ~n26692 | ~n26691;
  assign n26706 = ~n26694 & ~n26693;
  assign n26695 = n26705 ^ n26706;
  assign n26701 = ~n26695 | ~n26890;
  assign n26696 = ~P1_EAX_REG_26__SCAN_IN;
  assign n26699 = ~n26391 & ~n26696;
  assign n26697 = ~n43082 | ~P1_PHYADDRPOINTER_REG_26__SCAN_IN;
  assign n26698 = ~n26894 | ~n26697;
  assign n26700 = ~n26699 & ~n26698;
  assign n26704 = ~n26701 | ~n26700;
  assign n30700 = n26745 ^ P1_PHYADDRPOINTER_REG_26__SCAN_IN;
  assign n26703 = ~n30700 | ~n26900;
  assign n29992 = ~n26704 | ~n26703;
  assign n26786 = ~n26706 & ~n26705;
  assign n26709 = ~n26707 | ~P1_INSTQUEUE_REG_14__4__SCAN_IN;
  assign n26708 = ~n26870 | ~P1_INSTQUEUE_REG_2__4__SCAN_IN;
  assign n26713 = ~n26709 | ~n26708;
  assign n26711 = ~n26875 | ~P1_INSTQUEUE_REG_1__4__SCAN_IN;
  assign n26710 = ~n26686 | ~P1_INSTQUEUE_REG_8__4__SCAN_IN;
  assign n26712 = ~n26711 | ~n26710;
  assign n26721 = ~n26713 & ~n26712;
  assign n26715 = ~n26847 | ~P1_INSTQUEUE_REG_10__4__SCAN_IN;
  assign n26714 = ~n24947 | ~P1_INSTQUEUE_REG_13__4__SCAN_IN;
  assign n26719 = ~n26715 | ~n26714;
  assign n26717 = ~n26753 | ~P1_INSTQUEUE_REG_11__4__SCAN_IN;
  assign n26716 = ~n22842 | ~P1_INSTQUEUE_REG_3__4__SCAN_IN;
  assign n26718 = ~n26717 | ~n26716;
  assign n26720 = ~n26719 & ~n26718;
  assign n26737 = ~n26721 | ~n26720;
  assign n26723 = ~n25147 | ~P1_INSTQUEUE_REG_9__4__SCAN_IN;
  assign n26722 = ~n26577 | ~P1_INSTQUEUE_REG_4__4__SCAN_IN;
  assign n26727 = ~n26723 | ~n26722;
  assign n26725 = ~n26869 | ~P1_INSTQUEUE_REG_5__4__SCAN_IN;
  assign n26724 = ~n26866 | ~P1_INSTQUEUE_REG_12__4__SCAN_IN;
  assign n26726 = ~n26725 | ~n26724;
  assign n26735 = ~n26727 & ~n26726;
  assign n26729 = ~n26879 | ~P1_INSTQUEUE_REG_15__4__SCAN_IN;
  assign n26728 = ~n26818 | ~P1_INSTQUEUE_REG_0__4__SCAN_IN;
  assign n26733 = ~n26729 | ~n26728;
  assign n26731 = ~n26817 | ~P1_INSTQUEUE_REG_6__4__SCAN_IN;
  assign n26730 = ~n26859 | ~P1_INSTQUEUE_REG_7__4__SCAN_IN;
  assign n26732 = ~n26731 | ~n26730;
  assign n26734 = ~n26733 & ~n26732;
  assign n26736 = ~n26735 | ~n26734;
  assign n26784 = ~n26737 & ~n26736;
  assign n26738 = ~n26786 ^ n26784;
  assign n26744 = ~n26890 | ~n26738;
  assign n26739 = ~P1_EAX_REG_27__SCAN_IN;
  assign n26742 = ~n26391 & ~n26739;
  assign n26740 = ~n43082 | ~P1_PHYADDRPOINTER_REG_27__SCAN_IN;
  assign n26741 = ~n26894 | ~n26740;
  assign n26743 = ~n26742 & ~n26741;
  assign n26747 = n26744 & n26743;
  assign n30688 = ~P1_PHYADDRPOINTER_REG_27__SCAN_IN ^ n26794;
  assign n26746 = ~n30688 & ~n26894;
  assign n29968 = ~n26747 & ~n26746;
  assign n26752 = ~n25481 & ~n26748;
  assign n26749 = ~P1_INSTQUEUE_REG_4__5__SCAN_IN;
  assign n26751 = ~n26750 & ~n26749;
  assign n26755 = ~n26752 & ~n26751;
  assign n26754 = ~n26753 | ~P1_INSTQUEUE_REG_11__5__SCAN_IN;
  assign n26758 = ~n26755 | ~n26754;
  assign n26756 = ~P1_INSTQUEUE_REG_10__5__SCAN_IN;
  assign n26757 = ~n22833 & ~n26756;
  assign n26767 = ~n26758 & ~n26757;
  assign n26761 = ~n26866 | ~P1_INSTQUEUE_REG_12__5__SCAN_IN;
  assign n26760 = ~n26759 | ~P1_INSTQUEUE_REG_2__5__SCAN_IN;
  assign n26765 = ~n26761 | ~n26760;
  assign n26763 = ~n26818 | ~P1_INSTQUEUE_REG_0__5__SCAN_IN;
  assign n26762 = ~n22842 | ~P1_INSTQUEUE_REG_3__5__SCAN_IN;
  assign n26764 = ~n26763 | ~n26762;
  assign n26766 = ~n26765 & ~n26764;
  assign n26783 = ~n26767 | ~n26766;
  assign n26769 = ~n26879 | ~P1_INSTQUEUE_REG_15__5__SCAN_IN;
  assign n26768 = ~n26869 | ~P1_INSTQUEUE_REG_5__5__SCAN_IN;
  assign n26773 = ~n26769 | ~n26768;
  assign n26771 = ~n25147 | ~P1_INSTQUEUE_REG_9__5__SCAN_IN;
  assign n26770 = ~n26707 | ~P1_INSTQUEUE_REG_14__5__SCAN_IN;
  assign n26772 = ~n26771 | ~n26770;
  assign n26781 = ~n26773 & ~n26772;
  assign n26775 = ~n26622 | ~P1_INSTQUEUE_REG_13__5__SCAN_IN;
  assign n26774 = ~n26875 | ~P1_INSTQUEUE_REG_1__5__SCAN_IN;
  assign n26779 = ~n26775 | ~n26774;
  assign n26777 = ~n26686 | ~P1_INSTQUEUE_REG_8__5__SCAN_IN;
  assign n26776 = ~n26859 | ~P1_INSTQUEUE_REG_7__5__SCAN_IN;
  assign n26778 = ~n26777 | ~n26776;
  assign n26780 = ~n26779 & ~n26778;
  assign n26782 = ~n26781 | ~n26780;
  assign n26798 = ~n26783 & ~n26782;
  assign n26785 = ~n26784;
  assign n26797 = ~n26786 | ~n26785;
  assign n26787 = n26798 ^ n26797;
  assign n26793 = ~n26787 | ~n26890;
  assign n26788 = ~P1_EAX_REG_28__SCAN_IN;
  assign n26791 = n26391 | n26788;
  assign n26789 = ~n43082 | ~P1_PHYADDRPOINTER_REG_28__SCAN_IN;
  assign n26790 = n26894 & n26789;
  assign n26792 = n26791 & n26790;
  assign n26796 = ~n26793 | ~n26792;
  assign n30668 = ~P1_PHYADDRPOINTER_REG_28__SCAN_IN ^ n26842;
  assign n26795 = ~n30668 | ~n26900;
  assign n29949 = ~n26796 | ~n26795;
  assign n26845 = n26798 | n26797;
  assign n26802 = ~n25465 & ~n26799;
  assign n26801 = ~n25267 & ~n26800;
  assign n26804 = ~n26802 & ~n26801;
  assign n26803 = ~n26851 | ~P1_INSTQUEUE_REG_11__6__SCAN_IN;
  assign n26808 = ~n26804 | ~n26803;
  assign n26805 = ~P1_INSTQUEUE_REG_10__6__SCAN_IN;
  assign n26807 = ~n22833 & ~n26805;
  assign n26816 = ~n26808 & ~n26807;
  assign n26810 = ~n25147 | ~P1_INSTQUEUE_REG_9__6__SCAN_IN;
  assign n26809 = ~n22842 | ~P1_INSTQUEUE_REG_3__6__SCAN_IN;
  assign n26814 = ~n26810 | ~n26809;
  assign n26812 = ~n26622 | ~P1_INSTQUEUE_REG_13__6__SCAN_IN;
  assign n26811 = ~n26869 | ~P1_INSTQUEUE_REG_5__6__SCAN_IN;
  assign n26813 = ~n26812 | ~n26811;
  assign n26815 = ~n26814 & ~n26813;
  assign n26834 = ~n26816 | ~n26815;
  assign n26820 = ~n26817 | ~P1_INSTQUEUE_REG_6__6__SCAN_IN;
  assign n26819 = ~n26818 | ~P1_INSTQUEUE_REG_0__6__SCAN_IN;
  assign n26824 = ~n26820 | ~n26819;
  assign n26822 = ~n26707 | ~P1_INSTQUEUE_REG_14__6__SCAN_IN;
  assign n26821 = ~n26870 | ~P1_INSTQUEUE_REG_2__6__SCAN_IN;
  assign n26823 = ~n26822 | ~n26821;
  assign n26832 = ~n26824 & ~n26823;
  assign n26826 = ~n26879 | ~P1_INSTQUEUE_REG_15__6__SCAN_IN;
  assign n26825 = ~n26866 | ~P1_INSTQUEUE_REG_12__6__SCAN_IN;
  assign n26830 = ~n26826 | ~n26825;
  assign n26828 = ~n26875 | ~P1_INSTQUEUE_REG_1__6__SCAN_IN;
  assign n26827 = ~n26577 | ~P1_INSTQUEUE_REG_4__6__SCAN_IN;
  assign n26829 = ~n26828 | ~n26827;
  assign n26831 = ~n26830 & ~n26829;
  assign n26833 = ~n26832 | ~n26831;
  assign n26846 = ~n26834 & ~n26833;
  assign n26835 = n26845 ^ n26846;
  assign n26841 = ~n26835 | ~n26890;
  assign n26836 = ~P1_EAX_REG_29__SCAN_IN;
  assign n26839 = ~n26391 & ~n26836;
  assign n26837 = ~n43082 | ~P1_PHYADDRPOINTER_REG_29__SCAN_IN;
  assign n26838 = ~n26894 | ~n26837;
  assign n26840 = ~n26839 & ~n26838;
  assign n26844 = n26841 & n26840;
  assign n30658 = ~P1_PHYADDRPOINTER_REG_29__SCAN_IN ^ n26899;
  assign n26843 = ~n30658 & ~n26894;
  assign n29933 = ~n26844 & ~n26843;
  assign n26889 = ~n26846 & ~n26845;
  assign n26850 = ~n26847 | ~P1_INSTQUEUE_REG_10__7__SCAN_IN;
  assign n26849 = ~n25147 | ~P1_INSTQUEUE_REG_9__7__SCAN_IN;
  assign n26855 = ~n26850 | ~n26849;
  assign n26853 = ~n26851 | ~P1_INSTQUEUE_REG_11__7__SCAN_IN;
  assign n26852 = ~n22842 | ~P1_INSTQUEUE_REG_3__7__SCAN_IN;
  assign n26854 = ~n26853 | ~n26852;
  assign n26865 = ~n26855 & ~n26854;
  assign n26857 = ~n26622 | ~P1_INSTQUEUE_REG_13__7__SCAN_IN;
  assign n26856 = ~n25220 | ~P1_INSTQUEUE_REG_6__7__SCAN_IN;
  assign n26863 = ~n26857 | ~n26856;
  assign n26861 = ~n26858 | ~P1_INSTQUEUE_REG_8__7__SCAN_IN;
  assign n26860 = ~n26859 | ~P1_INSTQUEUE_REG_7__7__SCAN_IN;
  assign n26862 = ~n26861 | ~n26860;
  assign n26864 = ~n26863 & ~n26862;
  assign n26887 = ~n26865 | ~n26864;
  assign n26868 = ~n26707 | ~P1_INSTQUEUE_REG_14__7__SCAN_IN;
  assign n26867 = ~n26866 | ~P1_INSTQUEUE_REG_12__7__SCAN_IN;
  assign n26874 = ~n26868 | ~n26867;
  assign n26872 = ~n26869 | ~P1_INSTQUEUE_REG_5__7__SCAN_IN;
  assign n26871 = ~n26870 | ~P1_INSTQUEUE_REG_2__7__SCAN_IN;
  assign n26873 = ~n26872 | ~n26871;
  assign n26885 = ~n26874 & ~n26873;
  assign n26878 = ~n26875 | ~P1_INSTQUEUE_REG_1__7__SCAN_IN;
  assign n26877 = ~n26876 | ~P1_INSTQUEUE_REG_4__7__SCAN_IN;
  assign n26883 = ~n26878 | ~n26877;
  assign n26881 = ~n26879 | ~P1_INSTQUEUE_REG_15__7__SCAN_IN;
  assign n26880 = ~n26818 | ~P1_INSTQUEUE_REG_0__7__SCAN_IN;
  assign n26882 = ~n26881 | ~n26880;
  assign n26884 = ~n26883 & ~n26882;
  assign n26886 = ~n26885 | ~n26884;
  assign n26888 = ~n26887 & ~n26886;
  assign n26891 = ~n26889 ^ n26888;
  assign n26898 = ~n26891 | ~n26890;
  assign n26892 = ~P1_EAX_REG_30__SCAN_IN;
  assign n26896 = ~n26391 & ~n26892;
  assign n26893 = ~n43082 | ~P1_PHYADDRPOINTER_REG_30__SCAN_IN;
  assign n26895 = ~n26894 | ~n26893;
  assign n26897 = ~n26896 & ~n26895;
  assign n26902 = ~n26898 | ~n26897;
  assign n30647 = n26975 ^ P1_PHYADDRPOINTER_REG_30__SCAN_IN;
  assign n26901 = ~n30647 | ~n26900;
  assign n29910 = ~n26902 | ~n26901;
  assign n26906 = ~n26903 | ~P1_EAX_REG_31__SCAN_IN;
  assign n26905 = ~n26904 | ~P1_PHYADDRPOINTER_REG_31__SCAN_IN;
  assign n26907 = ~n26906 | ~n26905;
  assign n26909 = ~n42461 & ~n44850;
  assign n26921 = ~n31570 | ~n26909;
  assign n26918 = ~n23147 | ~n26910;
  assign n26916 = ~n25052 | ~n23072;
  assign n26913 = ~n43190 | ~n26912;
  assign n26915 = ~n26914 & ~n26913;
  assign n30346 = ~n26915 | ~n31502;
  assign n26917 = n26916 & n30346;
  assign n26919 = ~n26918 | ~n26917;
  assign n26920 = ~n26919 | ~n42372;
  assign n26924 = ~n26923 | ~n42599;
  assign n26959 = ~n26924 | ~n23952;
  assign n26926 = ~P1_ADDRESS_REG_22__SCAN_IN & ~P1_ADDRESS_REG_21__SCAN_IN;
  assign n26925 = ~P1_ADDRESS_REG_20__SCAN_IN & ~P1_ADDRESS_REG_19__SCAN_IN;
  assign n26930 = ~n26926 | ~n26925;
  assign n26928 = ~P1_ADDRESS_REG_26__SCAN_IN & ~P1_ADDRESS_REG_25__SCAN_IN;
  assign n26927 = ~P1_ADDRESS_REG_24__SCAN_IN & ~P1_ADDRESS_REG_23__SCAN_IN;
  assign n26929 = ~n26928 | ~n26927;
  assign n26951 = ~n26930 & ~n26929;
  assign n26932 = ~P1_ADDRESS_REG_14__SCAN_IN & ~P1_ADDRESS_REG_13__SCAN_IN;
  assign n26931 = ~P1_ADDRESS_REG_12__SCAN_IN & ~P1_ADDRESS_REG_11__SCAN_IN;
  assign n26936 = ~n26932 | ~n26931;
  assign n26934 = ~P1_ADDRESS_REG_18__SCAN_IN & ~P1_ADDRESS_REG_17__SCAN_IN;
  assign n26933 = ~P1_ADDRESS_REG_16__SCAN_IN & ~P1_ADDRESS_REG_15__SCAN_IN;
  assign n26935 = ~n26934 | ~n26933;
  assign n26938 = ~P1_ADDRESS_REG_6__SCAN_IN & ~P1_ADDRESS_REG_5__SCAN_IN;
  assign n26937 = ~P1_ADDRESS_REG_4__SCAN_IN & ~P1_ADDRESS_REG_3__SCAN_IN;
  assign n26942 = ~n26938 | ~n26937;
  assign n26940 = ~P1_ADDRESS_REG_1__SCAN_IN & ~P1_ADDRESS_REG_0__SCAN_IN;
  assign n26939 = ~P1_ADDRESS_REG_28__SCAN_IN & ~P1_ADDRESS_REG_27__SCAN_IN;
  assign n26941 = ~n26940 | ~n26939;
  assign n26947 = ~n26942 & ~n26941;
  assign n26944 = ~P1_ADDRESS_REG_10__SCAN_IN & ~P1_ADDRESS_REG_9__SCAN_IN;
  assign n26943 = ~P1_ADDRESS_REG_8__SCAN_IN & ~P1_ADDRESS_REG_7__SCAN_IN;
  assign n26945 = ~n26944 | ~n26943;
  assign n26946 = ~n26945 & ~P1_ADDRESS_REG_2__SCAN_IN;
  assign n26948 = ~n26947 | ~n26946;
  assign n26950 = ~n26949 & ~n26948;
  assign n26952 = ~n26951 | ~n26950;
  assign n26953 = ~n25678 | ~n43062;
  assign n26958 = ~n26954 | ~DATAI_31_;
  assign n26955 = ~n25678 | ~n43060;
  assign n26957 = ~n26956 | ~BUF1_REG_31__SCAN_IN;
  assign P1_U2873 = ~n26959 | ~n23947;
  assign n26960 = n25877 & P1_STATE2_REG_1__SCAN_IN;
  assign n26961 = n42234 | n26960;
  assign n26974 = ~n26961 | ~n44851;
  assign n27056 = ~n42227;
  assign n26963 = ~n31535 | ~n26962;
  assign n26969 = ~n27056 | ~n26963;
  assign n26965 = n26964;
  assign n26966 = ~n44514;
  assign n26967 = ~n26965 & ~n26966;
  assign n26968 = ~n31417 | ~n26967;
  assign n26970 = ~n44851 & ~n44853;
  assign n26971 = ~P1_STATE2_REG_3__SCAN_IN | ~n26970;
  assign n42469 = ~n26974 | ~n26973;
  assign n26976 = ~n26975 | ~P1_PHYADDRPOINTER_REG_30__SCAN_IN;
  assign n30639 = ~P1_PHYADDRPOINTER_REG_31__SCAN_IN ^ n26976;
  assign n31566 = ~n31582 | ~n44765;
  assign n26978 = n31566 & P1_EBX_REG_31__SCAN_IN;
  assign n26979 = ~n42391 | ~n26978;
  assign n26990 = ~n42503 | ~n42488;
  assign n44676 = ~P1_REIP_REG_27__SCAN_IN;
  assign n44671 = ~P1_REIP_REG_26__SCAN_IN;
  assign n26992 = ~n44676 & ~n44671;
  assign n26984 = n26992 & P1_REIP_REG_28__SCAN_IN;
  assign n30263 = ~n42469;
  assign n44661 = ~P1_REIP_REG_24__SCAN_IN;
  assign n30080 = ~P1_REIP_REG_21__SCAN_IN | ~P1_REIP_REG_20__SCAN_IN;
  assign n30079 = ~P1_REIP_REG_18__SCAN_IN | ~P1_REIP_REG_17__SCAN_IN;
  assign n44621 = ~P1_REIP_REG_16__SCAN_IN;
  assign n44611 = ~P1_REIP_REG_14__SCAN_IN;
  assign n44586 = ~P1_REIP_REG_9__SCAN_IN;
  assign n44576 = ~P1_REIP_REG_7__SCAN_IN;
  assign n44566 = ~P1_REIP_REG_5__SCAN_IN;
  assign n26980 = ~P1_REIP_REG_3__SCAN_IN | ~P1_REIP_REG_2__SCAN_IN;
  assign n42404 = ~n44815 & ~n26980;
  assign n42379 = ~P1_REIP_REG_4__SCAN_IN | ~n42404;
  assign n42355 = ~n44566 & ~n42379;
  assign n42334 = ~P1_REIP_REG_6__SCAN_IN | ~n42355;
  assign n42313 = ~n44576 & ~n42334;
  assign n42296 = ~P1_REIP_REG_8__SCAN_IN | ~n42313;
  assign n30328 = ~n44586 & ~n42296;
  assign n30264 = ~P1_REIP_REG_10__SCAN_IN | ~n30328;
  assign n30265 = ~P1_REIP_REG_12__SCAN_IN | ~P1_REIP_REG_11__SCAN_IN;
  assign n26981 = ~n30264 & ~n30265;
  assign n30245 = ~P1_REIP_REG_13__SCAN_IN | ~n26981;
  assign n30218 = ~n44611 & ~n30245;
  assign n30202 = ~P1_REIP_REG_15__SCAN_IN | ~n30218;
  assign n30141 = ~n44621 & ~n30202;
  assign n26982 = ~P1_REIP_REG_19__SCAN_IN | ~n30141;
  assign n30075 = ~n30079 & ~n26982;
  assign n26983 = ~P1_REIP_REG_22__SCAN_IN | ~n30075;
  assign n30060 = ~n30080 & ~n26983;
  assign n30015 = ~P1_REIP_REG_23__SCAN_IN | ~n30060;
  assign n30017 = ~n44661 & ~n30015;
  assign n26991 = ~P1_REIP_REG_25__SCAN_IN | ~n30017;
  assign n29976 = ~n30263 & ~n26991;
  assign n26987 = ~n26984 | ~n29976;
  assign n26998 = ~n26985 | ~n44765;
  assign n26995 = ~n23678 | ~n42391;
  assign n29959 = ~n26987 | ~n42500;
  assign n44692 = ~P1_REIP_REG_30__SCAN_IN;
  assign n44686 = ~P1_REIP_REG_29__SCAN_IN;
  assign n26993 = ~n44692 & ~n44686;
  assign n26988 = n26993 | n30287;
  assign n29924 = ~n29959 | ~n26988;
  assign n26989 = ~P1_REIP_REG_31__SCAN_IN | ~n29924;
  assign n27004 = n26990 & n26989;
  assign n44681 = ~P1_REIP_REG_28__SCAN_IN;
  assign n30005 = ~n30327 & ~n26991;
  assign n29960 = ~n30005 | ~n26992;
  assign n29943 = ~n44681 & ~n29960;
  assign n26994 = ~n29943 | ~n26993;
  assign n27002 = ~P1_REIP_REG_31__SCAN_IN & ~n26994;
  assign n26996 = n42760 & P1_EBX_REG_31__SCAN_IN;
  assign n26997 = ~n26996 & ~n26995;
  assign n27000 = ~n42481 | ~P1_EBX_REG_31__SCAN_IN;
  assign n42470 = n42469 & P1_STATE2_REG_3__SCAN_IN;
  assign n26999 = ~n42470 | ~P1_PHYADDRPOINTER_REG_31__SCAN_IN;
  assign n27001 = ~n27000 | ~n26999;
  assign n27003 = ~n27002 & ~n27001;
  assign P1_U2809 = ~n22937 | ~n23976;
  assign n27010 = ~P2_BE_N_REG_0__SCAN_IN & ~P2_BE_N_REG_1__SCAN_IN;
  assign n27006 = ~P2_BE_N_REG_2__SCAN_IN & ~P2_BE_N_REG_3__SCAN_IN;
  assign n27005 = ~P2_D_C_N_REG_SCAN_IN & ~P2_ADS_N_REG_SCAN_IN;
  assign n27008 = ~n27006 | ~n27005;
  assign n27007 = ~P2_W_R_N_REG_SCAN_IN | ~P2_M_IO_N_REG_SCAN_IN;
  assign n27009 = ~n27008 & ~n27007;
  assign n27046 = ~n27010 | ~n27009;
  assign U215 = P2_ADDRESS_REG_29__SCAN_IN | n27046;
  assign n27016 = ~P1_W_R_N_REG_SCAN_IN | ~P1_M_IO_N_REG_SCAN_IN;
  assign n27012 = ~P1_D_C_N_REG_SCAN_IN & ~P1_ADS_N_REG_SCAN_IN;
  assign n27011 = ~P1_BE_N_REG_2__SCAN_IN & ~P1_BE_N_REG_3__SCAN_IN;
  assign n27014 = n27012 & n27011;
  assign n27013 = ~P1_BE_N_REG_0__SCAN_IN & ~P1_BE_N_REG_1__SCAN_IN;
  assign n27015 = ~n27014 | ~n27013;
  assign n27017 = ~n27016 & ~n27015;
  assign n27019 = ~P2_ADDRESS_REG_6__SCAN_IN & ~P2_ADDRESS_REG_5__SCAN_IN;
  assign n27018 = ~P2_ADDRESS_REG_4__SCAN_IN & ~P2_ADDRESS_REG_3__SCAN_IN;
  assign n27023 = ~n27019 | ~n27018;
  assign n27021 = ~P2_ADDRESS_REG_1__SCAN_IN & ~P2_ADDRESS_REG_0__SCAN_IN;
  assign n27020 = ~P2_ADDRESS_REG_28__SCAN_IN & ~P2_ADDRESS_REG_27__SCAN_IN;
  assign n27022 = ~n27021 | ~n27020;
  assign n27028 = ~n27023 & ~n27022;
  assign n27025 = ~P2_ADDRESS_REG_10__SCAN_IN & ~P2_ADDRESS_REG_9__SCAN_IN;
  assign n27024 = ~P2_ADDRESS_REG_8__SCAN_IN & ~P2_ADDRESS_REG_7__SCAN_IN;
  assign n27026 = ~n27025 | ~n27024;
  assign n27027 = ~n27026 & ~P2_ADDRESS_REG_2__SCAN_IN;
  assign n27044 = ~n27028 | ~n27027;
  assign n27030 = ~P2_ADDRESS_REG_22__SCAN_IN & ~P2_ADDRESS_REG_21__SCAN_IN;
  assign n27029 = ~P2_ADDRESS_REG_20__SCAN_IN & ~P2_ADDRESS_REG_19__SCAN_IN;
  assign n27034 = ~n27030 | ~n27029;
  assign n27032 = ~P2_ADDRESS_REG_26__SCAN_IN & ~P2_ADDRESS_REG_25__SCAN_IN;
  assign n27031 = ~P2_ADDRESS_REG_24__SCAN_IN & ~P2_ADDRESS_REG_23__SCAN_IN;
  assign n27033 = ~n27032 | ~n27031;
  assign n27042 = ~n27034 & ~n27033;
  assign n27036 = ~P2_ADDRESS_REG_14__SCAN_IN & ~P2_ADDRESS_REG_13__SCAN_IN;
  assign n27035 = ~P2_ADDRESS_REG_12__SCAN_IN & ~P2_ADDRESS_REG_11__SCAN_IN;
  assign n27040 = ~n27036 | ~n27035;
  assign n27038 = ~P2_ADDRESS_REG_18__SCAN_IN & ~P2_ADDRESS_REG_17__SCAN_IN;
  assign n27037 = ~P2_ADDRESS_REG_16__SCAN_IN & ~P2_ADDRESS_REG_15__SCAN_IN;
  assign n27039 = ~n27038 | ~n27037;
  assign n27041 = ~n27040 & ~n27039;
  assign n27043 = ~n27042 | ~n27041;
  assign n33460 = ~n40437 & ~n27046;
  assign n42232 = ~P1_STATE_REG_2__SCAN_IN & ~n42244;
  assign n27047 = ~HOLD | ~n42232;
  assign n44530 = ~P1_STATE_REG_1__SCAN_IN | ~n44850;
  assign n27052 = ~n27047 | ~n44530;
  assign n41918 = ~HOLD;
  assign n27049 = ~n44546 & ~n41918;
  assign n27048 = ~P1_STATE_REG_0__SCAN_IN | ~P1_REQUESTPENDING_REG_SCAN_IN;
  assign n27050 = n27049 | n27048;
  assign n27051 = ~n44841 | ~n27050;
  assign P1_U3195 = n27052 | n27051;
  assign n27053 = ~n44745 | ~n44845;
  assign n27058 = ~n31420 | ~n44514;
  assign n27054 = ~n31568 | ~n44845;
  assign n27055 = ~n31439 & ~n27054;
  assign n27057 = ~n27056 | ~n27055;
  assign P1_U2905 = n42755 & P1_DATAO_REG_31__SCAN_IN;
  assign n27059 = ~n23742 | ~P1_INSTADDRPOINTER_REG_18__SCAN_IN;
  assign n30790 = P1_INSTADDRPOINTER_REG_19__SCAN_IN ^ n23166;
  assign n27062 = ~n30791 & ~n30790;
  assign n31151 = ~P1_INSTADDRPOINTER_REG_19__SCAN_IN;
  assign n27061 = ~n23166 & ~n31151;
  assign n27090 = ~n27062 & ~n27061;
  assign n27063 = ~n23166 ^ P1_INSTADDRPOINTER_REG_20__SCAN_IN;
  assign n30786 = ~n27090 ^ n27063;
  assign n27089 = n30786 & n43042;
  assign n31231 = ~n43014 | ~n31277;
  assign n31162 = ~n27064 & ~n31231;
  assign n31268 = ~n27065;
  assign n31244 = ~P1_INSTADDRPOINTER_REG_0__SCAN_IN | ~n31268;
  assign n27067 = ~n27066 & ~n31244;
  assign n31259 = ~n31162 & ~n27067;
  assign n27079 = ~n31259 & ~n27068;
  assign n27075 = ~n27069;
  assign n31242 = ~n43031;
  assign n27070 = ~n27075 & ~n31242;
  assign n31150 = ~n27079 & ~n27070;
  assign n27071 = P1_INSTADDRPOINTER_REG_20__SCAN_IN | n31151;
  assign n27087 = n31150 | n27071;
  assign n27074 = ~n31242 & ~P1_INSTADDRPOINTER_REG_19__SCAN_IN;
  assign n42966 = ~n43014;
  assign n27073 = ~n42966 & ~n27072;
  assign n27077 = ~n27074 & ~n27073;
  assign n27076 = ~n42961 | ~n27075;
  assign n27078 = ~n27077 | ~n27076;
  assign n31147 = ~n31380 & ~n27078;
  assign n27080 = ~n27079 | ~n31151;
  assign n27081 = ~n31147 | ~n27080;
  assign n27085 = ~n27081 | ~P1_INSTADDRPOINTER_REG_20__SCAN_IN;
  assign n30396 = ~n30140 ^ n27082;
  assign n27083 = n30396 | n43001;
  assign n30780 = ~n42929 | ~P1_REIP_REG_20__SCAN_IN;
  assign n27084 = n27083 & n30780;
  assign n27086 = n27085 & n27084;
  assign n27088 = ~n27087 | ~n27086;
  assign P1_U3011 = n27089 | n27088;
  assign n27095 = ~n27090 | ~P1_INSTADDRPOINTER_REG_20__SCAN_IN;
  assign n27091 = ~n23166 & ~P1_INSTADDRPOINTER_REG_19__SCAN_IN;
  assign n27093 = ~n30791 | ~n27091;
  assign n27092 = ~n23166 | ~P1_INSTADDRPOINTER_REG_20__SCAN_IN;
  assign n27094 = ~n27093 | ~n27092;
  assign n27099 = ~n27096 | ~n42961;
  assign n27098 = ~n43014 | ~n27097;
  assign n27100 = ~n27099 | ~n27098;
  assign n31137 = ~n31380 & ~n27100;
  assign n27101 = ~P1_INSTADDRPOINTER_REG_21__SCAN_IN;
  assign n27110 = n31137 | n27101;
  assign n27105 = ~n27103 & ~n27104;
  assign n30390 = n27102 | n27105;
  assign n27108 = ~n30390 & ~n43001;
  assign n30766 = ~n42929 | ~P1_REIP_REG_21__SCAN_IN;
  assign n31131 = ~P1_INSTADDRPOINTER_REG_21__SCAN_IN & ~n31150;
  assign n27106 = ~n31134 | ~n31131;
  assign n27107 = ~n30766 | ~n27106;
  assign n27109 = ~n27108 & ~n27107;
  assign n29853 = ~P2_STATE2_REG_1__SCAN_IN | ~P2_STATEBS16_REG_SCAN_IN;
  assign n27111 = ~n29853 | ~n41664;
  assign n33131 = ~P2_STATE2_REG_0__SCAN_IN | ~n41664;
  assign n27113 = n27111 & n33131;
  assign n41887 = ~P2_STATE2_REG_0__SCAN_IN | ~n42204;
  assign n27112 = ~n42123 & ~n41887;
  assign n27114 = ~n27113 & ~n27112;
  assign n33265 = ~P2_STATE2_REG_0__SCAN_IN | ~n42181;
  assign n42079 = ~n33265;
  assign P2_U3178 = ~n27114 & ~n42079;
  assign n27117 = ~n29694 | ~P2_INSTQUEUE_REG_11__5__SCAN_IN;
  assign n27123 = ~n27118 | ~n27117;
  assign n27120 = ~n22864 | ~P2_INSTQUEUE_REG_15__5__SCAN_IN;
  assign n27122 = ~n27121 | ~n27120;
  assign n27131 = ~n27122 & ~n27123;
  assign n29688 = n42134 | n33165;
  assign n27200 = ~n29688;
  assign n27124 = ~n27200 | ~P2_INSTQUEUE_REG_14__5__SCAN_IN;
  assign n27129 = ~n27125 | ~n27124;
  assign n27127 = ~n27409 | ~P2_INSTQUEUE_REG_13__5__SCAN_IN;
  assign n27126 = ~n27279 | ~P2_INSTQUEUE_REG_9__5__SCAN_IN;
  assign n27128 = ~n27126 | ~n27127;
  assign n27130 = ~n27129 & ~n27128;
  assign n27147 = ~n27131 | ~n27130;
  assign n27133 = ~n29694 | ~P2_INSTQUEUE_REG_3__5__SCAN_IN;
  assign n27137 = ~n27134 | ~n27133;
  assign n27139 = ~n27409 | ~P2_INSTQUEUE_REG_5__5__SCAN_IN;
  assign n27138 = ~n27279 | ~P2_INSTQUEUE_REG_1__5__SCAN_IN;
  assign n27143 = ~n27139 | ~n27138;
  assign n27141 = ~n22864 | ~P2_INSTQUEUE_REG_7__5__SCAN_IN;
  assign n27140 = ~n27200 | ~P2_INSTQUEUE_REG_6__5__SCAN_IN;
  assign n27142 = ~n27141 | ~n27140;
  assign n27144 = ~n27142 & ~n27143;
  assign n27146 = ~n27145 | ~n27144;
  assign n27612 = ~n27146 | ~n27147;
  assign n27179 = ~n27612;
  assign n27148 = ~n29694 | ~P2_INSTQUEUE_REG_11__6__SCAN_IN;
  assign n27154 = ~n27149 | ~n27148;
  assign n27150 = ~P2_INSTQUEUE_REG_13__6__SCAN_IN;
  assign n27152 = ~n27409 | ~P2_INSTQUEUE_REG_13__6__SCAN_IN;
  assign n27153 = ~n27152 | ~n27151;
  assign n27164 = ~n27154 & ~n27153;
  assign n27156 = ~n27155 | ~P2_INSTQUEUE_REG_10__6__SCAN_IN;
  assign n27157 = ~P2_INSTQUEUE_REG_15__6__SCAN_IN;
  assign n27160 = ~n27158 | ~P2_INSTQUEUE_REG_12__6__SCAN_IN;
  assign n27159 = ~n27200 | ~P2_INSTQUEUE_REG_14__6__SCAN_IN;
  assign n27161 = ~n27160 | ~n27159;
  assign n27178 = ~n27164 | ~n27163;
  assign n27166 = ~n22863 | ~P2_INSTQUEUE_REG_7__6__SCAN_IN;
  assign n27165 = ~n27200 | ~P2_INSTQUEUE_REG_6__6__SCAN_IN;
  assign n27169 = ~n27166 | ~n27165;
  assign n27168 = ~n27279 | ~P2_INSTQUEUE_REG_1__6__SCAN_IN;
  assign n27167 = ~n27409 | ~P2_INSTQUEUE_REG_5__6__SCAN_IN;
  assign n27170 = ~n27219 | ~P2_INSTQUEUE_REG_3__6__SCAN_IN;
  assign n27175 = ~n27171 | ~n27170;
  assign n27172 = ~n27412 & ~n40530;
  assign n27174 = ~n27172;
  assign n27173 = ~n27158 | ~P2_INSTQUEUE_REG_4__6__SCAN_IN;
  assign n27181 = ~n29694 | ~P2_INSTQUEUE_REG_11__3__SCAN_IN;
  assign n27185 = ~n27182 | ~n27181;
  assign n27187 = ~n27409 | ~P2_INSTQUEUE_REG_13__3__SCAN_IN;
  assign n27186 = ~n27279 | ~P2_INSTQUEUE_REG_9__3__SCAN_IN;
  assign n27190 = ~n27187 | ~n27186;
  assign n27189 = ~n22864 | ~P2_INSTQUEUE_REG_15__3__SCAN_IN;
  assign n27260 = ~n29688;
  assign n27188 = ~n27260 | ~P2_INSTQUEUE_REG_14__3__SCAN_IN;
  assign n27194 = ~n27413 | ~P2_INSTQUEUE_REG_1__3__SCAN_IN;
  assign n27193 = ~n27409 | ~P2_INSTQUEUE_REG_5__3__SCAN_IN;
  assign n27198 = ~n27194 | ~n27193;
  assign n27197 = ~n27196 | ~n27195;
  assign n27207 = ~n27198 & ~n27197;
  assign n27199 = ~n27155 | ~P2_INSTQUEUE_REG_2__3__SCAN_IN;
  assign n27201 = ~n27421 | ~P2_INSTQUEUE_REG_6__3__SCAN_IN;
  assign n27205 = ~n27202 | ~n27201;
  assign n27204 = ~n27389 | ~P2_INSTQUEUE_REG_7__3__SCAN_IN;
  assign n27203 = ~n29694 | ~P2_INSTQUEUE_REG_3__3__SCAN_IN;
  assign n40486 = ~n27631;
  assign n27276 = ~n27632 | ~n40486;
  assign n27211 = ~n27409 | ~P2_INSTQUEUE_REG_13__7__SCAN_IN;
  assign n27210 = ~n27413 | ~P2_INSTQUEUE_REG_9__7__SCAN_IN;
  assign n27215 = ~n27211 | ~n27210;
  assign n27212 = ~n27260 | ~P2_INSTQUEUE_REG_14__7__SCAN_IN;
  assign n27214 = ~n27213 | ~n27212;
  assign n27225 = ~n27215 & ~n27214;
  assign n28017 = ~P2_INSTQUEUE_REG_10__7__SCAN_IN;
  assign n27217 = ~n27389 | ~P2_INSTQUEUE_REG_15__7__SCAN_IN;
  assign n27223 = ~n27218 | ~n27217;
  assign n27220 = ~n29694 | ~P2_INSTQUEUE_REG_11__7__SCAN_IN;
  assign n27222 = ~n27221 | ~n27220;
  assign n28020 = ~P2_INSTQUEUE_REG_2__7__SCAN_IN;
  assign n27227 = ~n29694 | ~P2_INSTQUEUE_REG_3__7__SCAN_IN;
  assign n27232 = ~n27228 | ~n27227;
  assign n27229 = ~n27260 | ~P2_INSTQUEUE_REG_6__7__SCAN_IN;
  assign n27231 = ~n27230 | ~n27229;
  assign n27240 = ~n27232 & ~n27231;
  assign n27234 = ~n27409 | ~P2_INSTQUEUE_REG_5__7__SCAN_IN;
  assign n27233 = ~n27413 | ~P2_INSTQUEUE_REG_1__7__SCAN_IN;
  assign n27238 = ~n27234 | ~n27233;
  assign n40545 = ~P2_INSTQUEUE_REG_0__7__SCAN_IN;
  assign n27236 = n27412 | n40545;
  assign n27235 = ~n27389 | ~P2_INSTQUEUE_REG_7__7__SCAN_IN;
  assign n27237 = ~n27236 | ~n27235;
  assign n27239 = ~n27238 & ~n27237;
  assign n27244 = ~n27413 | ~P2_INSTQUEUE_REG_9__4__SCAN_IN;
  assign n27243 = ~n27409 | ~P2_INSTQUEUE_REG_13__4__SCAN_IN;
  assign n27248 = ~n27244 | ~n27243;
  assign n27476 = ~P2_INSTQUEUE_REG_12__4__SCAN_IN;
  assign n29116 = ~P2_INSTQUEUE_REG_8__4__SCAN_IN;
  assign n27247 = ~n27246 | ~n27245;
  assign n27257 = ~n27248 & ~n27247;
  assign n29126 = ~P2_INSTQUEUE_REG_10__4__SCAN_IN;
  assign n27250 = ~n27260 | ~P2_INSTQUEUE_REG_14__4__SCAN_IN;
  assign n27255 = ~n27251 | ~n27250;
  assign n27253 = ~n29694 | ~P2_INSTQUEUE_REG_11__4__SCAN_IN;
  assign n27252 = ~n27389 | ~P2_INSTQUEUE_REG_15__4__SCAN_IN;
  assign n27254 = ~n27253 | ~n27252;
  assign n27256 = ~n27255 & ~n27254;
  assign n27273 = ~n27257 | ~n27256;
  assign n27259 = ~n27409 | ~P2_INSTQUEUE_REG_5__4__SCAN_IN;
  assign n27258 = ~n27413 | ~P2_INSTQUEUE_REG_1__4__SCAN_IN;
  assign n27264 = ~n27259 | ~n27258;
  assign n27262 = ~n22863 | ~P2_INSTQUEUE_REG_7__4__SCAN_IN;
  assign n27261 = ~n27260 | ~P2_INSTQUEUE_REG_6__4__SCAN_IN;
  assign n27263 = ~n27261 | ~n27262;
  assign n27271 = ~n27264 & ~n27263;
  assign n27453 = ~P2_INSTQUEUE_REG_2__4__SCAN_IN;
  assign n27266 = ~n29694 | ~P2_INSTQUEUE_REG_3__4__SCAN_IN;
  assign n29111 = ~P2_INSTQUEUE_REG_4__4__SCAN_IN;
  assign n27272 = ~n27270 | ~n27271;
  assign n27277 = n27273 & n27272;
  assign n27626 = ~n27610 | ~n27277;
  assign n27274 = ~n27277;
  assign n40552 = n27613;
  assign n27278 = ~n40501 & ~n40552;
  assign n40519 = ~n27612;
  assign n27281 = ~n27409 | ~P2_INSTQUEUE_REG_13__2__SCAN_IN;
  assign n27280 = ~n27413 | ~P2_INSTQUEUE_REG_9__2__SCAN_IN;
  assign n27285 = ~n27281 | ~n27280;
  assign n27283 = ~n27389 | ~P2_INSTQUEUE_REG_15__2__SCAN_IN;
  assign n27282 = ~n27200 | ~P2_INSTQUEUE_REG_14__2__SCAN_IN;
  assign n27284 = ~n27283 | ~n27282;
  assign n27294 = ~n27285 & ~n27284;
  assign n29502 = ~P2_INSTQUEUE_REG_10__2__SCAN_IN;
  assign n27288 = n27286 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n27287 = ~n29694 | ~P2_INSTQUEUE_REG_11__2__SCAN_IN;
  assign n27292 = ~n27288 | ~n27287;
  assign n27290 = n27412 | n29497;
  assign n29498 = ~P2_INSTQUEUE_REG_12__2__SCAN_IN;
  assign n27291 = ~n27290 | ~n27289;
  assign n27293 = ~n27292 & ~n27291;
  assign n27310 = ~n27294 | ~n27293;
  assign n27295 = ~n27413 | ~P2_INSTQUEUE_REG_1__2__SCAN_IN;
  assign n27297 = ~n22863 | ~P2_INSTQUEUE_REG_7__2__SCAN_IN;
  assign n27296 = ~n29694 | ~P2_INSTQUEUE_REG_3__2__SCAN_IN;
  assign n27298 = ~n27297 | ~n27296;
  assign n27308 = ~n27299 & ~n27298;
  assign n27300 = ~n27155 | ~P2_INSTQUEUE_REG_2__2__SCAN_IN;
  assign n27302 = n27300 & n29098;
  assign n27306 = ~n27302 | ~n27301;
  assign n27304 = n27412 | n40467;
  assign n27303 = ~n27260 | ~P2_INSTQUEUE_REG_6__2__SCAN_IN;
  assign n27305 = ~n27304 | ~n27303;
  assign n27307 = ~n27306 & ~n27305;
  assign n27309 = ~n27308 | ~n27307;
  assign n27312 = ~n27413 | ~P2_INSTQUEUE_REG_9__0__SCAN_IN;
  assign n27311 = ~n27409 | ~P2_INSTQUEUE_REG_13__0__SCAN_IN;
  assign n27316 = ~n27312 | ~n27311;
  assign n27313 = ~n29694 | ~P2_INSTQUEUE_REG_11__0__SCAN_IN;
  assign n27315 = ~n27314 | ~n27313;
  assign n27325 = ~n27316 & ~n27315;
  assign n27318 = ~n27389 | ~P2_INSTQUEUE_REG_15__0__SCAN_IN;
  assign n27323 = ~n27319 | ~n27318;
  assign n27421 = ~n29688;
  assign n27320 = ~n27421 | ~P2_INSTQUEUE_REG_14__0__SCAN_IN;
  assign n27322 = ~n27321 | ~n27320;
  assign n27324 = ~n27323 & ~n27322;
  assign n27327 = ~n27409 | ~P2_INSTQUEUE_REG_5__0__SCAN_IN;
  assign n27326 = ~n27413 | ~P2_INSTQUEUE_REG_1__0__SCAN_IN;
  assign n27331 = ~n27327 | ~n27326;
  assign n27329 = ~n22863 | ~P2_INSTQUEUE_REG_7__0__SCAN_IN;
  assign n27328 = ~n27421 | ~P2_INSTQUEUE_REG_6__0__SCAN_IN;
  assign n27330 = ~n27329 | ~n27328;
  assign n27340 = ~n27331 & ~n27330;
  assign n27333 = ~n29694 | ~P2_INSTQUEUE_REG_3__0__SCAN_IN;
  assign n27338 = ~n27334 | ~n27333;
  assign n27337 = ~n27336 | ~n27335;
  assign n27339 = ~n27338 & ~n27337;
  assign n27341 = ~n27340 | ~n27339;
  assign n27358 = ~n42120 ^ P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN;
  assign n27357 = ~n27358 | ~n27359;
  assign n27346 = ~n41769 | ~n42120;
  assign n27354 = ~n27357 | ~n27346;
  assign n27349 = ~n27348 | ~P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign n27444 = ~n29098 ^ P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN;
  assign n27355 = ~n27444;
  assign n27352 = ~n27446 | ~n27355;
  assign n27351 = ~n27447;
  assign n27364 = ~n27352 | ~n27351;
  assign n27353 = ~n27348 ^ P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign n27539 = ~n27354 ^ n27353;
  assign n27356 = ~n27552 | ~n27539;
  assign n27543 = ~n27446 ^ n27355;
  assign n27362 = ~n27566;
  assign n27361 = ~n27357;
  assign n27360 = ~n27358;
  assign n27522 = ~n27359;
  assign n27525 = ~n27361 & ~n28240;
  assign n27367 = ~n27362 | ~n27525;
  assign n27366 = ~n27364 | ~n27363;
  assign n27365 = ~P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN;
  assign n27551 = ~n27365 | ~P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN;
  assign n27370 = ~n42200;
  assign n39150 = ~n41002 & ~P2_STATE2_REG_1__SCAN_IN;
  assign n27369 = ~n39150 & ~P2_READREQUEST_REG_SCAN_IN;
  assign n27406 = ~n27370 & ~n27369;
  assign n27372 = ~n27413 | ~P2_INSTQUEUE_REG_9__1__SCAN_IN;
  assign n27371 = ~n27409 | ~P2_INSTQUEUE_REG_13__1__SCAN_IN;
  assign n27376 = ~n27372 | ~n27371;
  assign n27373 = ~n27421 | ~P2_INSTQUEUE_REG_14__1__SCAN_IN;
  assign n27375 = ~n27374 | ~n27373;
  assign n27386 = ~n27376 & ~n27375;
  assign n27378 = ~n27389 | ~P2_INSTQUEUE_REG_15__1__SCAN_IN;
  assign n27384 = ~n27379 | ~n27378;
  assign n27380 = ~n27412;
  assign n27382 = ~n27380 | ~P2_INSTQUEUE_REG_8__1__SCAN_IN;
  assign n27381 = ~n29694 | ~P2_INSTQUEUE_REG_11__1__SCAN_IN;
  assign n27383 = ~n27382 | ~n27381;
  assign n27403 = ~n27386 | ~n27385;
  assign n27388 = ~n27409 | ~P2_INSTQUEUE_REG_5__1__SCAN_IN;
  assign n27387 = ~n27413 | ~P2_INSTQUEUE_REG_1__1__SCAN_IN;
  assign n27393 = ~n27388 | ~n27387;
  assign n27391 = ~n22863 | ~P2_INSTQUEUE_REG_7__1__SCAN_IN;
  assign n27390 = ~n27421 | ~P2_INSTQUEUE_REG_6__1__SCAN_IN;
  assign n27392 = ~n27391 | ~n27390;
  assign n27401 = ~n27393 & ~n27392;
  assign n27394 = ~n27155 | ~P2_INSTQUEUE_REG_2__1__SCAN_IN;
  assign n27395 = ~n29694 | ~P2_INSTQUEUE_REG_3__1__SCAN_IN;
  assign n27399 = ~n27396 | ~n27395;
  assign n27398 = ~n27380 | ~P2_INSTQUEUE_REG_0__1__SCAN_IN;
  assign n27397 = ~n27158 | ~P2_INSTQUEUE_REG_4__1__SCAN_IN;
  assign n27402 = ~n27401 | ~n27400;
  assign n27404 = ~n27402 | ~n27403;
  assign n27627 = ~n42216 | ~n31677;
  assign n27405 = ~n42200 & ~n31964;
  assign P2_U3612 = n27406 | n27405;
  assign n27407 = ~n42123 & ~P2_STATE2_REG_0__SCAN_IN;
  assign n42206 = ~n23278 & ~n27407;
  assign n27564 = ~n42206 & ~n42181;
  assign n27408 = ~P2_INSTQUEUE_REG_10__3__SCAN_IN;
  assign n27411 = n29575 | n27408;
  assign n27845 = ~P2_INSTQUEUE_REG_6__3__SCAN_IN;
  assign n27417 = ~n27411 | ~n27410;
  assign n29718 = n27412;
  assign n29355 = n29752 & n29098;
  assign n27415 = ~n29530 | ~P2_INSTQUEUE_REG_1__3__SCAN_IN;
  assign n29660 = n27413;
  assign n27852 = ~P2_INSTQUEUE_REG_2__3__SCAN_IN;
  assign n27414 = n29580 | n27852;
  assign n27416 = ~n27415 | ~n27414;
  assign n27427 = n27417 | n27416;
  assign n27420 = ~n27817 | ~P2_INSTQUEUE_REG_5__3__SCAN_IN;
  assign n27419 = n33147 | n29283;
  assign n27425 = ~n27420 | ~n27419;
  assign n29602 = ~n23145 | ~n29098;
  assign n27423 = n29602 | n29278;
  assign n29569 = ~n27421 | ~n29098;
  assign n28763 = ~P2_INSTQUEUE_REG_7__3__SCAN_IN;
  assign n27422 = n29569 | n28763;
  assign n27424 = ~n27423 | ~n27422;
  assign n27443 = ~n27427 & ~n27426;
  assign n29099 = ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n27431 = ~n28734 | ~P2_INSTQUEUE_REG_14__3__SCAN_IN;
  assign n27429 = n27428;
  assign n29591 = n27429 & n27570;
  assign n27430 = ~n29591 | ~P2_INSTQUEUE_REG_13__3__SCAN_IN;
  assign n27437 = ~n27431 | ~n27430;
  assign n27432 = n33186 & n42120;
  assign n29592 = n27432 & n27570;
  assign n27435 = ~n29592 | ~P2_INSTQUEUE_REG_15__3__SCAN_IN;
  assign n27434 = ~n29588 | ~P2_INSTQUEUE_REG_0__3__SCAN_IN;
  assign n27436 = ~n27435 | ~n27434;
  assign n27438 = ~n27437 & ~n27436;
  assign n29436 = n29752 & P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n27440 = ~n29436 | ~P2_INSTQUEUE_REG_9__3__SCAN_IN;
  assign n27439 = n29581 | n29394;
  assign n27441 = ~n27440 | ~n27439;
  assign n31598 = n28543 & n27536;
  assign n27445 = ~n28283 | ~n27444;
  assign n27448 = ~n28283 | ~n27447;
  assign n27452 = n29575 | n29126;
  assign n27450 = ~P2_INSTQUEUE_REG_6__4__SCAN_IN;
  assign n27451 = n29577 | n27450;
  assign n27457 = ~n27452 | ~n27451;
  assign n29519 = n29355;
  assign n27455 = ~n29519 | ~P2_INSTQUEUE_REG_1__4__SCAN_IN;
  assign n27454 = n29580 | n27453;
  assign n27456 = ~n27455 | ~n27454;
  assign n27465 = n27457 | n27456;
  assign n27459 = ~n27817 | ~P2_INSTQUEUE_REG_5__4__SCAN_IN;
  assign n27458 = n33147 | n29116;
  assign n27463 = ~n27459 | ~n27458;
  assign n27461 = n29602 | n29111;
  assign n29447 = ~P2_INSTQUEUE_REG_7__4__SCAN_IN;
  assign n27460 = n29569 | n29447;
  assign n27462 = ~n27461 | ~n27460;
  assign n27464 = n27463 | n27462;
  assign n27482 = ~n27465 & ~n27464;
  assign n27467 = ~n28734 | ~P2_INSTQUEUE_REG_14__4__SCAN_IN;
  assign n27466 = ~n29591 | ~P2_INSTQUEUE_REG_13__4__SCAN_IN;
  assign n27471 = ~n27467 | ~n27466;
  assign n27469 = ~n29592 | ~P2_INSTQUEUE_REG_15__4__SCAN_IN;
  assign n27468 = ~n29588 | ~P2_INSTQUEUE_REG_0__4__SCAN_IN;
  assign n27470 = ~n27469 | ~n27468;
  assign n27475 = ~n27471 & ~n27470;
  assign n27473 = ~n27509 | ~P2_INSTQUEUE_REG_11__4__SCAN_IN;
  assign n29597 = n27510;
  assign n27472 = ~n29597 | ~P2_INSTQUEUE_REG_3__4__SCAN_IN;
  assign n27474 = n27473 & n27472;
  assign n27480 = ~n27475 | ~n27474;
  assign n27478 = ~n29436 | ~P2_INSTQUEUE_REG_9__4__SCAN_IN;
  assign n27477 = n29581 | n27476;
  assign n27479 = ~n27478 | ~n27477;
  assign n27481 = ~n27480 & ~n27479;
  assign n27484 = ~n31598 | ~n28601;
  assign n27550 = ~n28283 | ~n27483;
  assign n27485 = ~n27484 | ~n27550;
  assign n28060 = ~n27549 | ~n27485;
  assign n28051 = ~n27486 ^ n23950;
  assign n28245 = n28051 & n28060;
  assign n27487 = ~n28245;
  assign n27548 = ~n27487 | ~n28283;
  assign n27489 = ~n29519 | ~P2_INSTQUEUE_REG_1__0__SCAN_IN;
  assign n27488 = n29581 | n29537;
  assign n27493 = ~n27489 | ~n27488;
  assign n27491 = ~n29436 | ~P2_INSTQUEUE_REG_9__0__SCAN_IN;
  assign n27490 = n33147 | n29536;
  assign n27492 = ~n27491 | ~n27490;
  assign n27502 = n27493 | n27492;
  assign n27496 = n29580 | n27494;
  assign n27495 = n29575 | n29527;
  assign n27500 = ~n27496 | ~n27495;
  assign n29558 = ~P2_INSTQUEUE_REG_6__0__SCAN_IN;
  assign n27497 = n29602 | n29540;
  assign n27499 = ~n27498 | ~n27497;
  assign n27520 = ~n27502 & ~n27501;
  assign n27504 = ~n28734 | ~P2_INSTQUEUE_REG_14__0__SCAN_IN;
  assign n27503 = ~n29588 | ~P2_INSTQUEUE_REG_0__0__SCAN_IN;
  assign n27508 = ~n27504 | ~n27503;
  assign n27506 = ~n29591 | ~P2_INSTQUEUE_REG_13__0__SCAN_IN;
  assign n27505 = ~n29592 | ~P2_INSTQUEUE_REG_15__0__SCAN_IN;
  assign n27507 = ~n27506 | ~n27505;
  assign n27514 = ~n27508 & ~n27507;
  assign n27512 = ~n27509 | ~P2_INSTQUEUE_REG_11__0__SCAN_IN;
  assign n27511 = ~n27510 | ~P2_INSTQUEUE_REG_3__0__SCAN_IN;
  assign n27513 = n27512 & n27511;
  assign n27518 = ~n27514 | ~n27513;
  assign n27516 = ~n27817 | ~P2_INSTQUEUE_REG_5__0__SCAN_IN;
  assign n28647 = ~P2_INSTQUEUE_REG_7__0__SCAN_IN;
  assign n27515 = n29569 | n28647;
  assign n27517 = ~n27516 | ~n27515;
  assign n27519 = ~n27518 & ~n27517;
  assign n28554 = ~n27520 | ~n27519;
  assign n28285 = ~n28554;
  assign n27524 = ~n31598 | ~n28285;
  assign n27521 = ~n33186 | ~P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n27565 = ~n27522 | ~n27521;
  assign n27523 = ~n28283 | ~n27565;
  assign n28241 = ~n27524 | ~n27523;
  assign n27527 = ~n28241 | ~n42208;
  assign n27528 = ~n27525;
  assign n27526 = ~n40444 & ~n27528;
  assign n27535 = ~n27527 | ~n27526;
  assign n27530 = ~n31598 | ~n27528;
  assign n27529 = ~n31598 | ~n27565;
  assign n27533 = ~n27530 | ~n27529;
  assign n27655 = ~n27531 | ~n27404;
  assign n27537 = ~n27539;
  assign n27532 = ~n27655 & ~n27537;
  assign n27534 = ~n27533 & ~n27532;
  assign n27542 = ~n27535 | ~n27534;
  assign n40456 = n28543;
  assign n27538 = ~n42209 | ~n40456;
  assign n27540 = ~n27538 | ~n27537;
  assign n28054 = ~n28283 | ~n27539;
  assign n27541 = ~n27540 | ~n28054;
  assign n27545 = ~n27542 | ~n27541;
  assign n27544 = ~n27543;
  assign n27546 = ~n27545 | ~n27544;
  assign n27559 = ~n27548 | ~n27547;
  assign n27553 = ~n31598 | ~n27552;
  assign n27555 = ~n27554 | ~n27553;
  assign n27557 = ~n27555 | ~P2_STATE2_REG_0__SCAN_IN;
  assign n27556 = ~n42214 | ~n33213;
  assign n27558 = ~n27557 | ~n27556;
  assign n27567 = n27565 | n27566;
  assign n27568 = ~n33240 | ~n27567;
  assign n27575 = ~n27568 | ~n42123;
  assign n27571 = ~n33186 | ~n22856;
  assign n27572 = ~n27571 | ~n27570;
  assign n27574 = ~n27572 | ~n33213;
  assign n27573 = ~n42123 & ~P2_FLUSH_REG_SCAN_IN;
  assign n42180 = ~n27574 | ~n27573;
  assign n27576 = n33217 | P2_FLUSH_REG_SCAN_IN;
  assign n27577 = ~n27576 | ~n42079;
  assign n42186 = n41786 & n27577;
  assign P2_U3047 = n42186 & P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN;
  assign n27578 = ~n42234 & ~P1_READREQUEST_REG_SCAN_IN;
  assign n27582 = n44838 | n27578;
  assign n27580 = ~n31497 | ~n27579;
  assign n27581 = ~n44838 | ~n27580;
  assign P1_U3487 = ~n27582 | ~n27581;
  assign n27585 = ~n37482 | ~n34971;
  assign n27589 = ~n34483 & ~n27588;
  assign n35745 = ~n34971 | ~n35504;
  assign n27594 = ~P3_EAX_REG_0__SCAN_IN & ~n35745;
  assign n27592 = ~BUF2_REG_0__SCAN_IN | ~n35807;
  assign n27591 = ~P3_EAX_REG_0__SCAN_IN | ~n35799;
  assign n27593 = ~n27592 | ~n27591;
  assign n27597 = ~n27594 & ~n27593;
  assign n27596 = ~n35752 | ~n27595;
  assign P3_U2735 = ~n27597 | ~n27596;
  assign n27600 = n27608 & n40471;
  assign n27602 = ~n27608 & ~n40552;
  assign n27604 = n28543 & n40471;
  assign n27628 = ~n27607 | ~n27612;
  assign n28250 = n27608 & n27628;
  assign n27609 = ~n40501;
  assign n28261 = ~n27632 | ~n40501;
  assign n27616 = ~n27611 | ~n28512;
  assign n27614 = ~n22840 | ~n27613;
  assign n27615 = ~n28498 | ~n27631;
  assign n27623 = ~n28498;
  assign n27640 = ~n27623 | ~n28500;
  assign n27617 = ~n27640 | ~n39593;
  assign n27620 = n31598 & P2_STATE2_REG_0__SCAN_IN;
  assign n27621 = ~n27620 | ~n27622;
  assign n27624 = ~n27623 & ~n28499;
  assign n28318 = ~n23099;
  assign n27625 = ~n28318 | ~n33186;
  assign n27630 = ~n28543 & ~n40486;
  assign n27629 = ~n27628;
  assign n27634 = ~n27630 | ~n27629;
  assign n27633 = n27632 | n27631;
  assign n27636 = ~n42197 | ~P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n27642 = ~n27639 | ~n40444;
  assign n27641 = n27640 & P2_STATE2_REG_0__SCAN_IN;
  assign n27645 = ~n27643;
  assign n27647 = ~n27685;
  assign n27646 = ~n42208;
  assign n27651 = ~n27724 | ~P2_EBX_REG_0__SCAN_IN;
  assign n27649 = ~n42197;
  assign n27648 = ~P2_STATE2_REG_1__SCAN_IN | ~P2_PHYADDRPOINTER_REG_0__SCAN_IN;
  assign n27650 = n27649 & n27648;
  assign n27652 = ~n27651 | ~n27650;
  assign n27654 = ~n27653 & ~n27652;
  assign n27657 = ~n28542 & ~n27656;
  assign n27658 = ~n28493;
  assign n27663 = ~n27658 | ~P2_STATE2_REG_0__SCAN_IN;
  assign n27659 = n40444 | n42214;
  assign n27662 = ~n27661 | ~n27660;
  assign n27683 = ~n27662 | ~n27663;
  assign n27664 = ~n27685 & ~n40456;
  assign n27666 = ~n27683 & ~n27664;
  assign n27667 = ~n28317 | ~P2_INSTADDRPOINTER_REG_0__SCAN_IN;
  assign n40343 = n27669;
  assign n27671 = ~n29320 | ~n42134;
  assign n27670 = n41002 | P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n27673 = ~n42214 & ~P2_STATE2_REG_3__SCAN_IN;
  assign n27675 = n27656 & n27673;
  assign n27674 = ~n40456 | ~P2_INSTQUEUE_REG_0__0__SCAN_IN;
  assign n27676 = ~n27675 | ~n27674;
  assign n33230 = ~n27677 | ~n27678;
  assign n27682 = ~n42177 | ~n39782;
  assign n28057 = ~P2_EBX_REG_0__SCAN_IN;
  assign n27680 = ~n39817 | ~n28057;
  assign n27679 = ~n40343 | ~n31948;
  assign n27681 = ~n27680 | ~n27679;
  assign P2_U2887 = ~n27682 | ~n27681;
  assign n27687 = ~n27683;
  assign n27684 = ~n42197 | ~P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN;
  assign n27686 = n27685 & n27684;
  assign n27744 = ~n27689 | ~n27688;
  assign n27696 = ~n28317 | ~P2_INSTADDRPOINTER_REG_1__SCAN_IN;
  assign n27691 = ~n23098 | ~P2_EBX_REG_1__SCAN_IN;
  assign n27690 = ~P2_STATE2_REG_1__SCAN_IN | ~P2_PHYADDRPOINTER_REG_1__SCAN_IN;
  assign n27694 = ~n27691 | ~n27690;
  assign n27692 = ~P2_REIP_REG_1__SCAN_IN;
  assign n27745 = ~n27696 | ~n27695;
  assign n27698 = ~n23099 | ~P2_EBX_REG_2__SCAN_IN;
  assign n27697 = ~P2_STATE2_REG_1__SCAN_IN | ~P2_PHYADDRPOINTER_REG_2__SCAN_IN;
  assign n27701 = ~n27698 | ~n27697;
  assign n27699 = ~P2_REIP_REG_2__SCAN_IN;
  assign n27703 = ~n27701 & ~n27700;
  assign n27702 = ~n28317 | ~P2_INSTADDRPOINTER_REG_2__SCAN_IN;
  assign n27734 = ~n27703 | ~n27702;
  assign n27705 = ~n23087 | ~n27734;
  assign n27704 = ~n27715 | ~n28328;
  assign n27709 = ~n27705 | ~n27704;
  assign n27708 = ~n27729 | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n27706 = ~n42214 | ~P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign n27707 = n27706 & n42123;
  assign n27735 = ~n27708 | ~n27707;
  assign n27714 = ~n27709 | ~n27735;
  assign n27711 = ~n27722 | ~n28328;
  assign n27710 = ~n27715 | ~n27734;
  assign n27712 = ~n27711 | ~n27710;
  assign n28325 = ~n27735;
  assign n27713 = ~n27712 | ~n28325;
  assign n27717 = ~n27714 | ~n27713;
  assign n27719 = ~n27722;
  assign n28327 = ~n27723 | ~n23087;
  assign n27726 = ~n23098 | ~P2_EBX_REG_3__SCAN_IN;
  assign n27725 = ~P2_STATE2_REG_1__SCAN_IN | ~P2_PHYADDRPOINTER_REG_3__SCAN_IN;
  assign n27728 = ~n27727 | ~n22959;
  assign n28332 = ~n27728 & ~n22914;
  assign n27731 = ~n27729 | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n27730 = ~n42197 | ~P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN;
  assign n28335 = ~n27731 | ~n27730;
  assign n27739 = ~n28332 ^ n28335;
  assign n27733 = ~n27739;
  assign n27737 = ~n27733 | ~n27732;
  assign n27738 = ~n27735 | ~n27734;
  assign n27736 = ~n27739 | ~n27738;
  assign n27741 = ~n27740;
  assign n27746 = ~n27745;
  assign n27750 = ~n41503 | ~P2_INSTQUEUE_REG_12__1__SCAN_IN;
  assign n28678 = ~P2_INSTQUEUE_REG_7__1__SCAN_IN;
  assign n27752 = n27751;
  assign n29424 = ~P2_INSTQUEUE_REG_1__1__SCAN_IN;
  assign n27753 = ~n27896 | ~P2_INSTQUEUE_REG_11__1__SCAN_IN;
  assign n27755 = ~n27754 | ~n27753;
  assign n27760 = ~n27908 | ~P2_INSTQUEUE_REG_15__1__SCAN_IN;
  assign n27892 = ~n27758 | ~n27752;
  assign n28700 = ~P2_INSTQUEUE_REG_5__1__SCAN_IN;
  assign n28681 = ~P2_INSTQUEUE_REG_3__1__SCAN_IN;
  assign n27762 = ~n27889 | ~P2_INSTQUEUE_REG_14__1__SCAN_IN;
  assign n27764 = ~n27763 | ~n27762;
  assign n29222 = ~P2_INSTQUEUE_REG_6__1__SCAN_IN;
  assign n41574 = ~n27774 | ~n27765;
  assign n28682 = ~P2_INSTQUEUE_REG_13__1__SCAN_IN;
  assign n27766 = n41574 | n28682;
  assign n27772 = ~n27767 | ~n27766;
  assign n27770 = n27905 | n29226;
  assign n27769 = ~n27881 | ~P2_INSTQUEUE_REG_8__1__SCAN_IN;
  assign n27771 = ~n27769 | ~n27770;
  assign n27778 = ~n41336 | ~P2_INSTQUEUE_REG_10__1__SCAN_IN;
  assign n27776 = ~n27900 | ~P2_INSTQUEUE_REG_9__1__SCAN_IN;
  assign n27782 = ~n27778 | ~n27777;
  assign n27783 = n29575 | n29502;
  assign n29520 = ~P2_INSTQUEUE_REG_6__2__SCAN_IN;
  assign n27786 = ~n29530 | ~P2_INSTQUEUE_REG_1__2__SCAN_IN;
  assign n27784 = ~P2_INSTQUEUE_REG_2__2__SCAN_IN;
  assign n27785 = n29580 | n27784;
  assign n27787 = ~n27786 | ~n27785;
  assign n27789 = ~n27817 | ~P2_INSTQUEUE_REG_5__2__SCAN_IN;
  assign n27788 = n33147 | n29497;
  assign n27794 = ~n27789 | ~n27788;
  assign n27792 = n29602 | n29501;
  assign n27790 = ~P2_INSTQUEUE_REG_7__2__SCAN_IN;
  assign n27791 = n29569 | n27790;
  assign n27793 = ~n27792 | ~n27791;
  assign n27809 = ~n27796 & ~n27795;
  assign n27798 = ~n28734 | ~P2_INSTQUEUE_REG_14__2__SCAN_IN;
  assign n27797 = ~n29591 | ~P2_INSTQUEUE_REG_13__2__SCAN_IN;
  assign n27802 = ~n27798 | ~n27797;
  assign n27800 = ~n29592 | ~P2_INSTQUEUE_REG_15__2__SCAN_IN;
  assign n27799 = ~n29588 | ~P2_INSTQUEUE_REG_0__2__SCAN_IN;
  assign n27801 = ~n27800 | ~n27799;
  assign n27804 = ~n27802 & ~n27801;
  assign n27803 = ~n27510 | ~P2_INSTQUEUE_REG_3__2__SCAN_IN;
  assign n27806 = ~n29436 | ~P2_INSTQUEUE_REG_9__2__SCAN_IN;
  assign n27805 = n29581 | n29498;
  assign n27807 = ~n27806 | ~n27805;
  assign n33116 = n28285 | n40456;
  assign n27843 = ~n33116;
  assign n27812 = n29575 | n27810;
  assign n27811 = n29577 | n29222;
  assign n27816 = ~n27812 | ~n27811;
  assign n27814 = ~n29519 | ~P2_INSTQUEUE_REG_1__1__SCAN_IN;
  assign n27813 = n29580 | n29426;
  assign n27815 = ~n27814 | ~n27813;
  assign n27825 = n27816 | n27815;
  assign n29491 = n27817;
  assign n27819 = ~n29491 | ~P2_INSTQUEUE_REG_5__1__SCAN_IN;
  assign n27818 = n33147 | n28670;
  assign n27823 = ~n27819 | ~n27818;
  assign n27821 = n29602 | n29226;
  assign n27820 = n29569 | n28678;
  assign n27822 = ~n27821 | ~n27820;
  assign n27824 = n27823 | n27822;
  assign n27842 = ~n27825 & ~n27824;
  assign n27827 = ~n28734 | ~P2_INSTQUEUE_REG_14__1__SCAN_IN;
  assign n27826 = ~n29591 | ~P2_INSTQUEUE_REG_13__1__SCAN_IN;
  assign n27831 = ~n27827 | ~n27826;
  assign n27829 = ~n29592 | ~P2_INSTQUEUE_REG_15__1__SCAN_IN;
  assign n27828 = ~n29588 | ~P2_INSTQUEUE_REG_0__1__SCAN_IN;
  assign n27830 = ~n27829 | ~n27828;
  assign n27835 = ~n27831 & ~n27830;
  assign n27833 = ~n27509 | ~P2_INSTQUEUE_REG_11__1__SCAN_IN;
  assign n27832 = ~n27510 | ~P2_INSTQUEUE_REG_3__1__SCAN_IN;
  assign n27834 = n27833 & n27832;
  assign n27840 = ~n27835 | ~n27834;
  assign n27838 = ~n29436 | ~P2_INSTQUEUE_REG_9__1__SCAN_IN;
  assign n27837 = n29581 | n27836;
  assign n27839 = ~n27838 | ~n27837;
  assign n27841 = ~n27840 & ~n27839;
  assign n28565 = ~n27842 | ~n27841;
  assign n28767 = ~P2_INSTQUEUE_REG_13__3__SCAN_IN;
  assign n27846 = n41574 | n28767;
  assign n27851 = ~n27847 | ~n27846;
  assign n27848 = ~n27881 | ~P2_INSTQUEUE_REG_8__3__SCAN_IN;
  assign n27850 = ~n27849 | ~n27848;
  assign n27860 = ~n27851 & ~n27850;
  assign n40421 = ~n27882;
  assign n27854 = ~n40421 | ~P2_INSTQUEUE_REG_0__3__SCAN_IN;
  assign n27857 = ~n41336 | ~P2_INSTQUEUE_REG_10__3__SCAN_IN;
  assign n27855 = ~n27900 | ~P2_INSTQUEUE_REG_9__3__SCAN_IN;
  assign n27856 = n27855 & n40456;
  assign n27858 = ~n27857 | ~n27856;
  assign n27862 = ~n41418 | ~P2_INSTQUEUE_REG_11__3__SCAN_IN;
  assign n27866 = ~n27862 | ~n27861;
  assign n27864 = ~n41503 | ~P2_INSTQUEUE_REG_12__3__SCAN_IN;
  assign n27865 = ~n27864 | ~n27863;
  assign n27875 = ~n27866 & ~n27865;
  assign n27868 = ~n27889 | ~P2_INSTQUEUE_REG_14__3__SCAN_IN;
  assign n28766 = ~P2_INSTQUEUE_REG_3__3__SCAN_IN;
  assign n27873 = ~n27868 | ~n27867;
  assign n27869 = ~n27892;
  assign n27871 = ~n27869 | ~P2_INSTQUEUE_REG_5__3__SCAN_IN;
  assign n27870 = ~n27908 | ~P2_INSTQUEUE_REG_15__3__SCAN_IN;
  assign n27872 = ~n27870 | ~n27871;
  assign n27874 = ~n27873 & ~n27872;
  assign n27878 = ~n28595 | ~n42208;
  assign n27885 = ~n27881 | ~P2_INSTQUEUE_REG_8__5__SCAN_IN;
  assign n27888 = ~n41336 | ~P2_INSTQUEUE_REG_10__5__SCAN_IN;
  assign n27891 = ~n27889 | ~P2_INSTQUEUE_REG_14__5__SCAN_IN;
  assign n29350 = ~P2_INSTQUEUE_REG_1__5__SCAN_IN;
  assign n27895 = ~n27891 | ~n27890;
  assign n29356 = ~P2_INSTQUEUE_REG_3__5__SCAN_IN;
  assign n27894 = n40734 | n29356;
  assign n28840 = ~P2_INSTQUEUE_REG_5__5__SCAN_IN;
  assign n27899 = ~n41418 | ~P2_INSTQUEUE_REG_11__5__SCAN_IN;
  assign n28845 = ~P2_INSTQUEUE_REG_7__5__SCAN_IN;
  assign n27902 = ~n27956 | ~P2_INSTQUEUE_REG_9__5__SCAN_IN;
  assign n28865 = ~P2_INSTQUEUE_REG_13__5__SCAN_IN;
  assign n27901 = n41574 | n28865;
  assign n27903 = n27902 & n27901;
  assign n29651 = ~P2_INSTQUEUE_REG_6__5__SCAN_IN;
  assign n27907 = n27904 | n29651;
  assign n27906 = n27905 | n29365;
  assign n27911 = ~n27907 | ~n27906;
  assign n41766 = ~n41782;
  assign n27909 = ~P2_INSTQUEUE_REG_15__5__SCAN_IN;
  assign n27910 = ~n41766 & ~n27909;
  assign n27912 = ~n27911 & ~n27910;
  assign n27946 = ~n27913 | ~n27912;
  assign n27915 = n29575 | n29656;
  assign n27914 = n29577 | n29651;
  assign n27920 = ~n27915 | ~n27914;
  assign n27918 = ~n29530 | ~P2_INSTQUEUE_REG_1__5__SCAN_IN;
  assign n27917 = n29580 | n27916;
  assign n27919 = ~n27918 | ~n27917;
  assign n27928 = n27920 | n27919;
  assign n27922 = ~n27817 | ~P2_INSTQUEUE_REG_5__5__SCAN_IN;
  assign n27921 = n33147 | n29669;
  assign n27926 = ~n27922 | ~n27921;
  assign n27924 = n29602 | n29365;
  assign n27923 = n29569 | n28845;
  assign n27925 = ~n27924 | ~n27923;
  assign n27927 = n27926 | n27925;
  assign n27944 = ~n27928 & ~n27927;
  assign n27930 = ~n28734 | ~P2_INSTQUEUE_REG_14__5__SCAN_IN;
  assign n27929 = ~n29591 | ~P2_INSTQUEUE_REG_13__5__SCAN_IN;
  assign n27934 = ~n27930 | ~n27929;
  assign n27932 = ~n29592 | ~P2_INSTQUEUE_REG_15__5__SCAN_IN;
  assign n27931 = ~n29588 | ~P2_INSTQUEUE_REG_0__5__SCAN_IN;
  assign n27933 = ~n27932 | ~n27931;
  assign n27938 = ~n27934 & ~n27933;
  assign n27936 = ~n27509 | ~P2_INSTQUEUE_REG_11__5__SCAN_IN;
  assign n27935 = ~n27510 | ~P2_INSTQUEUE_REG_3__5__SCAN_IN;
  assign n27937 = n27936 & n27935;
  assign n27942 = ~n27938 | ~n27937;
  assign n27940 = ~n29436 | ~P2_INSTQUEUE_REG_9__5__SCAN_IN;
  assign n27939 = n29581 | n29670;
  assign n27941 = ~n27940 | ~n27939;
  assign n27943 = ~n27942 & ~n27941;
  assign n28609 = ~n27944 | ~n27943;
  assign n27945 = n28609 | n40456;
  assign n27947 = ~n28070;
  assign n27949 = ~n41782 | ~P2_INSTQUEUE_REG_15__6__SCAN_IN;
  assign n28905 = ~P2_INSTQUEUE_REG_5__6__SCAN_IN;
  assign n27948 = n27892 | n28905;
  assign n27953 = ~n27949 | ~n27948;
  assign n27951 = ~n27889 | ~P2_INSTQUEUE_REG_14__6__SCAN_IN;
  assign n27952 = ~n27951 | ~n27950;
  assign n27964 = ~n27953 & ~n27952;
  assign n27955 = ~n41418 | ~P2_INSTQUEUE_REG_11__6__SCAN_IN;
  assign n27954 = ~n41503 | ~P2_INSTQUEUE_REG_12__6__SCAN_IN;
  assign n27962 = ~n27955 | ~n27954;
  assign n27958 = ~n27956 | ~P2_INSTQUEUE_REG_9__6__SCAN_IN;
  assign n27957 = n41574 | n27150;
  assign n27960 = n27958 & n27957;
  assign n27988 = ~P2_INSTQUEUE_REG_7__6__SCAN_IN;
  assign n27959 = n27897 | n27988;
  assign n27961 = ~n27960 | ~n27959;
  assign n27963 = ~n27962 & ~n27961;
  assign n27978 = ~n27964 | ~n27963;
  assign n27966 = ~n41336 | ~P2_INSTQUEUE_REG_10__6__SCAN_IN;
  assign n27965 = n27883 | n40530;
  assign n27970 = ~n27966 | ~n27965;
  assign n27968 = ~n27881 | ~P2_INSTQUEUE_REG_8__6__SCAN_IN;
  assign n27967 = n40657 | n27981;
  assign n27969 = ~n27968 | ~n27967;
  assign n27976 = ~n27970 & ~n27969;
  assign n29712 = ~P2_INSTQUEUE_REG_6__6__SCAN_IN;
  assign n27972 = n27904 | n29712;
  assign n27971 = n27905 | n29717;
  assign n27974 = ~n27972 | ~n27971;
  assign n28904 = ~P2_INSTQUEUE_REG_3__6__SCAN_IN;
  assign n27973 = ~n40734 & ~n28904;
  assign n27975 = ~n27974 & ~n27973;
  assign n27977 = ~n27976 | ~n27975;
  assign n27980 = n29575 | n29687;
  assign n27979 = n29577 | n29712;
  assign n27985 = ~n27980 | ~n27979;
  assign n27983 = ~n29519 | ~P2_INSTQUEUE_REG_1__6__SCAN_IN;
  assign n27982 = n29580 | n27981;
  assign n27984 = ~n27983 | ~n27982;
  assign n27994 = n27985 | n27984;
  assign n27987 = ~n27817 | ~P2_INSTQUEUE_REG_5__6__SCAN_IN;
  assign n27986 = n33147 | n29576;
  assign n27992 = ~n27987 | ~n27986;
  assign n27990 = n29602 | n29717;
  assign n27989 = n29569 | n27988;
  assign n27991 = ~n27990 | ~n27989;
  assign n27993 = n27992 | n27991;
  assign n28010 = ~n27994 & ~n27993;
  assign n27996 = ~n28734 | ~P2_INSTQUEUE_REG_14__6__SCAN_IN;
  assign n27995 = ~n29591 | ~P2_INSTQUEUE_REG_13__6__SCAN_IN;
  assign n28000 = ~n27996 | ~n27995;
  assign n27998 = ~n29592 | ~P2_INSTQUEUE_REG_15__6__SCAN_IN;
  assign n27997 = ~n29588 | ~P2_INSTQUEUE_REG_0__6__SCAN_IN;
  assign n27999 = ~n27998 | ~n27997;
  assign n28004 = ~n28000 & ~n27999;
  assign n28002 = ~n27509 | ~P2_INSTQUEUE_REG_11__6__SCAN_IN;
  assign n28001 = ~n29597 | ~P2_INSTQUEUE_REG_3__6__SCAN_IN;
  assign n28003 = n28002 & n28001;
  assign n28008 = ~n28004 | ~n28003;
  assign n28006 = ~n29436 | ~P2_INSTQUEUE_REG_9__6__SCAN_IN;
  assign n28005 = n29581 | n29574;
  assign n28007 = ~n28006 | ~n28005;
  assign n28009 = ~n28008 & ~n28007;
  assign n28616 = ~n28010 | ~n28009;
  assign n28011 = n28616 | n40456;
  assign n28014 = ~n28012 | ~n28011;
  assign n28016 = ~n28015 | ~n28014;
  assign n28019 = n29575 | n28017;
  assign n29730 = ~P2_INSTQUEUE_REG_6__7__SCAN_IN;
  assign n28018 = n29577 | n29730;
  assign n28024 = ~n28019 | ~n28018;
  assign n28022 = ~n29530 | ~P2_INSTQUEUE_REG_1__7__SCAN_IN;
  assign n28021 = n29580 | n28020;
  assign n28023 = ~n28022 | ~n28021;
  assign n28026 = ~n29491 | ~P2_INSTQUEUE_REG_5__7__SCAN_IN;
  assign n28025 = n33147 | n29749;
  assign n28031 = ~n28026 | ~n28025;
  assign n28029 = n29602 | n28027;
  assign n28928 = ~P2_INSTQUEUE_REG_7__7__SCAN_IN;
  assign n28028 = n29569 | n28928;
  assign n28030 = ~n28029 | ~n28028;
  assign n28050 = ~n28033 & ~n28032;
  assign n28035 = ~n28734 | ~P2_INSTQUEUE_REG_14__7__SCAN_IN;
  assign n28034 = ~n29591 | ~P2_INSTQUEUE_REG_13__7__SCAN_IN;
  assign n28039 = ~n28035 | ~n28034;
  assign n28037 = ~n29592 | ~P2_INSTQUEUE_REG_15__7__SCAN_IN;
  assign n28036 = ~n29588 | ~P2_INSTQUEUE_REG_0__7__SCAN_IN;
  assign n28038 = ~n28037 | ~n28036;
  assign n28043 = ~n28039 & ~n28038;
  assign n28041 = ~n27509 | ~P2_INSTQUEUE_REG_11__7__SCAN_IN;
  assign n28040 = ~n29597 | ~P2_INSTQUEUE_REG_3__7__SCAN_IN;
  assign n28042 = n28041 & n28040;
  assign n28048 = ~n28043 | ~n28042;
  assign n28046 = ~n29436 | ~P2_INSTQUEUE_REG_9__7__SCAN_IN;
  assign n28047 = ~n28046 | ~n28045;
  assign n28049 = ~n28048 & ~n28047;
  assign n28077 = ~n28050 | ~n28049;
  assign n28053 = n28051 | n28552;
  assign n28052 = ~n28552 | ~P2_EBX_REG_3__SCAN_IN;
  assign n28091 = ~n28053 | ~n28052;
  assign n28055 = ~P2_EBX_REG_2__SCAN_IN;
  assign n28056 = ~n28552 | ~n28055;
  assign n28059 = ~n28565 | ~n40519;
  assign n28095 = ~n28552 | ~n28057;
  assign n28058 = n28095 | P2_EBX_REG_1__SCAN_IN;
  assign n28099 = ~n28059 | ~n28058;
  assign n28061 = ~n28552 | ~P2_EBX_REG_4__SCAN_IN;
  assign n28063 = ~n28552 | ~P2_EBX_REG_5__SCAN_IN;
  assign n39790 = ~P2_EBX_REG_6__SCAN_IN;
  assign n28065 = ~n28552 | ~n39790;
  assign n28066 = ~n23964 | ~n28065;
  assign n28067 = ~n28066;
  assign n28068 = ~n22872 | ~n28067;
  assign n39544 = ~n28076 | ~n28068;
  assign n28074 = ~n23914 | ~n23913;
  assign n39559 = ~n22872 | ~n28074;
  assign n28075 = P2_INSTADDRPOINTER_REG_6__SCAN_IN & P2_INSTADDRPOINTER_REG_5__SCAN_IN;
  assign n28079 = n28077 | n28552;
  assign n28078 = ~n28552 | ~P2_EBX_REG_7__SCAN_IN;
  assign n28081 = ~n28552 | ~P2_EBX_REG_8__SCAN_IN;
  assign n28083 = ~n28080;
  assign n28082 = ~n28081;
  assign n28084 = ~n28083 | ~n28082;
  assign n39498 = ~n28114 | ~n28084;
  assign n28085 = ~n29831 | ~P2_INSTADDRPOINTER_REG_8__SCAN_IN;
  assign n32533 = n39498 | n28085;
  assign n32529 = ~n28076 ^ n23036;
  assign n32530 = n32529 | n33023;
  assign n28086 = n32533 & n32530;
  assign n28093 = ~n28088 | ~n28071;
  assign n28092 = ~n28091 | ~n28090;
  assign n39605 = ~n23574 | ~n28092;
  assign n39629 = ~n28094 ^ n28099;
  assign n40302 = ~n39629 ^ P2_INSTADDRPOINTER_REG_2__SCAN_IN;
  assign n28096 = ~n28241 | ~n29824;
  assign n39682 = ~n28096 | ~n28095;
  assign n33123 = ~P2_INSTADDRPOINTER_REG_0__SCAN_IN;
  assign n28100 = ~n39682 & ~n33123;
  assign n28097 = P2_EBX_REG_0__SCAN_IN & P2_EBX_REG_1__SCAN_IN;
  assign n28098 = n28552 & n28097;
  assign n28101 = ~n28099 & ~n28098;
  assign n40320 = ~n28100 | ~n28101;
  assign n42096 = ~P2_INSTADDRPOINTER_REG_1__SCAN_IN;
  assign n28102 = ~n40320 | ~n42096;
  assign n33111 = ~n28100;
  assign n39665 = ~n28101;
  assign n40319 = ~n33111 | ~n39665;
  assign n40301 = n28102 & n40319;
  assign n28105 = ~n40302 | ~n40301;
  assign n28103 = ~n39629;
  assign n28104 = ~n28103 | ~P2_INSTADDRPOINTER_REG_2__SCAN_IN;
  assign n40284 = ~n28105 | ~n28104;
  assign n39583 = ~n23574 ^ n22865;
  assign n40289 = ~n39583 ^ P2_INSTADDRPOINTER_REG_4__SCAN_IN;
  assign n28106 = n40284 | P2_INSTADDRPOINTER_REG_3__SCAN_IN;
  assign n28107 = n40289 & n28106;
  assign n28110 = ~n28108 | ~n28107;
  assign n40368 = ~P2_INSTADDRPOINTER_REG_4__SCAN_IN;
  assign n28109 = n39583 | n40368;
  assign n28111 = ~n39498;
  assign n28112 = ~n28111 | ~n29831;
  assign n32532 = ~n28112 | ~n23429;
  assign n39521 = ~n32529;
  assign n28113 = n39521 | P2_INSTADDRPOINTER_REG_7__SCAN_IN;
  assign n32488 = n32532 & n28113;
  assign n28115 = n28552 & P2_EBX_REG_9__SCAN_IN;
  assign n28116 = ~n28114 | ~n28115;
  assign n39479 = n28118 & n28116;
  assign n28117 = ~n39479 | ~n29831;
  assign n32975 = ~P2_INSTADDRPOINTER_REG_9__SCAN_IN;
  assign n32509 = ~n28117 | ~n32975;
  assign n28121 = n32488 & n32509;
  assign n28119 = ~n28118 | ~n23040;
  assign n39458 = ~n28126 | ~n28119;
  assign n28120 = n39458 | n28071;
  assign n32502 = ~P2_INSTADDRPOINTER_REG_10__SCAN_IN;
  assign n32487 = ~n28120 | ~n32502;
  assign n28122 = n28121 & n32487;
  assign n28123 = ~n29831 | ~P2_INSTADDRPOINTER_REG_10__SCAN_IN;
  assign n32486 = n39458 | n28123;
  assign n28124 = n29831 & P2_INSTADDRPOINTER_REG_9__SCAN_IN;
  assign n32508 = ~n39479 | ~n28124;
  assign n28125 = n32486 & n32508;
  assign n28128 = ~n28126 | ~n28127;
  assign n39439 = n23904 & n28128;
  assign n28129 = ~n39439 | ~n29831;
  assign n32927 = ~P2_INSTADDRPOINTER_REG_11__SCAN_IN;
  assign n32469 = ~n28129 | ~n32927;
  assign n28130 = n29831 & P2_INSTADDRPOINTER_REG_11__SCAN_IN;
  assign n32468 = ~n39439 | ~n28130;
  assign n28132 = ~n28552 | ~P2_EBX_REG_12__SCAN_IN;
  assign n28133 = ~n28132;
  assign n28134 = ~n23904 | ~n28133;
  assign n39416 = ~n28137 | ~n28134;
  assign n28135 = ~n29831 | ~P2_INSTADDRPOINTER_REG_12__SCAN_IN;
  assign n32455 = ~n39416 & ~n28135;
  assign n28136 = n39416 | n28071;
  assign n32899 = ~P2_INSTADDRPOINTER_REG_12__SCAN_IN;
  assign n32454 = ~n28136 | ~n32899;
  assign n28155 = ~n28552 | ~P2_EBX_REG_15__SCAN_IN;
  assign n28146 = ~n28552 | ~P2_EBX_REG_16__SCAN_IN;
  assign n28138 = ~n28552 | ~P2_EBX_REG_19__SCAN_IN;
  assign n28139 = ~n28138;
  assign n28140 = ~n22871 | ~n28139;
  assign n28184 = n28174 & n28140;
  assign n28141 = ~n28184 | ~n29831;
  assign n32771 = ~P2_INSTADDRPOINTER_REG_19__SCAN_IN;
  assign n32345 = ~n28141 | ~n32771;
  assign n28143 = ~n28152 | ~n28142;
  assign n39296 = ~n22871 | ~n28143;
  assign n28187 = ~n39296;
  assign n32360 = ~n28187 | ~n29831;
  assign n28144 = ~n32360 | ~n32362;
  assign n29022 = ~n32345 | ~n28144;
  assign n28158 = ~n28145;
  assign n28147 = ~n28158 | ~n23917;
  assign n39340 = ~n28150 | ~n28147;
  assign n28148 = n39340 | n28071;
  assign n32390 = ~n28148 ^ P2_INSTADDRPOINTER_REG_16__SCAN_IN;
  assign n28151 = ~n28150 | ~n28149;
  assign n39313 = ~n28152 | ~n28151;
  assign n28153 = n39313 | n28071;
  assign n32808 = ~P2_INSTADDRPOINTER_REG_17__SCAN_IN;
  assign n32374 = ~n28153 | ~n32808;
  assign n28162 = ~n28154;
  assign n28156 = ~n28155;
  assign n28157 = ~n28162 | ~n28156;
  assign n28159 = ~n39356 | ~n29831;
  assign n32831 = ~P2_INSTADDRPOINTER_REG_15__SCAN_IN;
  assign n32402 = ~n28159 | ~n32831;
  assign n28161 = ~n28166 | ~n28160;
  assign n39376 = ~n28162 | ~n28161;
  assign n28163 = n39376 | n28071;
  assign n32858 = ~P2_INSTADDRPOINTER_REG_14__SCAN_IN;
  assign n32432 = ~n28163 | ~n32858;
  assign n28165 = ~n28137 | ~n28164;
  assign n28191 = n28166 & n28165;
  assign n28167 = ~n28191 | ~n29831;
  assign n32849 = ~P2_INSTADDRPOINTER_REG_13__SCAN_IN;
  assign n32437 = ~n28167 | ~n32849;
  assign n28168 = n32432 & n32437;
  assign n28169 = n32402 & n28168;
  assign n28170 = n32374 & n28169;
  assign n28171 = ~n32390 | ~n28170;
  assign n28177 = ~n29022 & ~n28171;
  assign n28172 = ~n28552 | ~P2_EBX_REG_20__SCAN_IN;
  assign n28173 = ~n28172;
  assign n28175 = ~n28174 | ~n28173;
  assign n39255 = ~n28178 | ~n28175;
  assign n29062 = ~P2_INSTADDRPOINTER_REG_20__SCAN_IN;
  assign n28176 = ~n29025 | ~n29062;
  assign n28182 = ~n28177 | ~n28176;
  assign n28180 = ~n28178 | ~n28179;
  assign n28201 = n22921 & n28180;
  assign n28181 = ~n28201 | ~n29831;
  assign n29075 = ~P2_INSTADDRPOINTER_REG_21__SCAN_IN;
  assign n29067 = n28181 & n29075;
  assign n28183 = ~n28182 & ~n29067;
  assign n29024 = ~n29025;
  assign n28200 = ~n29024 | ~P2_INSTADDRPOINTER_REG_20__SCAN_IN;
  assign n39280 = ~n28184;
  assign n28185 = ~n29831 | ~P2_INSTADDRPOINTER_REG_19__SCAN_IN;
  assign n28186 = n29831 & P2_INSTADDRPOINTER_REG_18__SCAN_IN;
  assign n28188 = ~n28187 | ~n28186;
  assign n29021 = ~n32344 | ~n28188;
  assign n28189 = n29831 & P2_INSTADDRPOINTER_REG_15__SCAN_IN;
  assign n32401 = ~n39356 | ~n28189;
  assign n28190 = ~n29831 | ~P2_INSTADDRPOINTER_REG_14__SCAN_IN;
  assign n32431 = n39376 | n28190;
  assign n39402 = ~n28191;
  assign n28192 = ~n29831 | ~P2_INSTADDRPOINTER_REG_13__SCAN_IN;
  assign n28193 = n32431 & n32436;
  assign n28195 = n32401 & n28193;
  assign n28194 = ~n29831 | ~P2_INSTADDRPOINTER_REG_16__SCAN_IN;
  assign n29020 = n39340 | n28194;
  assign n28197 = n28195 & n29020;
  assign n28196 = ~n29831 | ~P2_INSTADDRPOINTER_REG_17__SCAN_IN;
  assign n28198 = ~n28197 | ~n32373;
  assign n28199 = ~n29021 & ~n28198;
  assign n28203 = ~n28200 | ~n28199;
  assign n39243 = ~n28201;
  assign n28202 = ~n29831 | ~P2_INSTADDRPOINTER_REG_21__SCAN_IN;
  assign n29066 = ~n39243 & ~n28202;
  assign n28204 = ~n28203 & ~n29066;
  assign n28205 = ~n22921 | ~n23034;
  assign n39225 = ~n28208 | ~n28205;
  assign n28206 = ~n29831 | ~P2_INSTADDRPOINTER_REG_22__SCAN_IN;
  assign n32306 = n39225 | n28206;
  assign n28207 = n39225 | n28071;
  assign n32307 = ~n28207 | ~n32752;
  assign n28209 = ~n28208;
  assign n28210 = ~n28552 | ~P2_EBX_REG_23__SCAN_IN;
  assign n28215 = ~n28209 | ~n28210;
  assign n28211 = ~n28210;
  assign n28212 = ~n28208 | ~n28211;
  assign n31833 = ~n28215 | ~n28212;
  assign n28213 = n31833 | n28071;
  assign n28993 = ~P2_INSTADDRPOINTER_REG_23__SCAN_IN;
  assign n32292 = ~n28213 | ~n28993;
  assign n28214 = ~n29831 | ~P2_INSTADDRPOINTER_REG_23__SCAN_IN;
  assign n28216 = n28552 & P2_EBX_REG_24__SCAN_IN;
  assign n28217 = ~n28215 | ~n28216;
  assign n31814 = ~n22911 | ~n28217;
  assign n28218 = ~n29831 | ~P2_INSTADDRPOINTER_REG_24__SCAN_IN;
  assign n28219 = ~n31814;
  assign n28220 = ~n28219 | ~n29831;
  assign n32277 = ~n28220 | ~n32712;
  assign n28224 = n28552 & P2_EBX_REG_25__SCAN_IN;
  assign n28221 = ~n28224;
  assign n29825 = ~n28232;
  assign n32259 = ~n28223 ^ P2_INSTADDRPOINTER_REG_26__SCAN_IN;
  assign n28225 = ~n22911 | ~n28224;
  assign n31790 = ~n28226 | ~n28225;
  assign n28227 = ~n32254 | ~n23751;
  assign n29808 = ~n32259 | ~n28227;
  assign n28228 = ~n29808;
  assign n32256 = ~n32254;
  assign n28231 = ~n32256 | ~P2_INSTADDRPOINTER_REG_25__SCAN_IN;
  assign n28229 = n29831 & P2_INSTADDRPOINTER_REG_26__SCAN_IN;
  assign n28230 = ~n31768 | ~n28229;
  assign n28234 = ~n28236;
  assign n28233 = ~n29825 | ~n23045;
  assign n31746 = ~n29803 | ~n28233;
  assign n32224 = ~n28234 | ~n29805;
  assign n28235 = ~n29805;
  assign n28237 = ~n32224 | ~n32223;
  assign n28238 = n33228 | n40444;
  assign n28239 = n28238 & n40501;
  assign n28281 = ~n28239 | ~n33136;
  assign n28243 = n28241 | n28240;
  assign n28244 = ~n28243 | ~n28242;
  assign n28247 = ~n28245 | ~n28244;
  assign n33221 = ~n28247 | ~n28246;
  assign n28249 = ~n40456 | ~n28248;
  assign n28269 = ~n33217 & ~n28249;
  assign n28251 = ~n28250;
  assign n28253 = ~n28251 | ~n39805;
  assign n28252 = ~n31677;
  assign n28514 = n28253 & n28252;
  assign n28254 = ~n42208 | ~n40501;
  assign n28255 = ~n28254 | ~n39593;
  assign n28256 = ~n28255 | ~n39805;
  assign n28257 = n28256 & n40471;
  assign n28260 = ~n28514 & ~n28257;
  assign n28259 = n28499 & n23085;
  assign n28264 = n28260 & n28259;
  assign n28262 = ~n28261 | ~n40471;
  assign n28263 = ~n39140 | ~n28262;
  assign n28268 = ~n28264 | ~n28263;
  assign n41920 = ~P2_STATE_REG_0__SCAN_IN;
  assign n39153 = ~P2_STATE_REG_1__SCAN_IN;
  assign n28265 = ~n39153 ^ P2_STATE_REG_2__SCAN_IN;
  assign n41909 = ~n41920 | ~n28265;
  assign n31608 = ~n41909 & ~n41895;
  assign n33236 = ~n31608;
  assign n28266 = ~n27605 & ~n33236;
  assign n28267 = n33240 & n28266;
  assign n28278 = ~n28269 & ~n33141;
  assign n28270 = ~n41909 & ~n40471;
  assign n28271 = ~n27605;
  assign n28273 = ~n40456 | ~n28271;
  assign n28272 = ~n23706 | ~n42208;
  assign n28274 = ~n28273 | ~n28272;
  assign n28275 = ~n33240 | ~n28274;
  assign n28277 = ~n42204 | ~n28276;
  assign n28279 = ~n28278 | ~n28277;
  assign n28280 = ~n29800 & ~n28279;
  assign n28282 = ~n28281 | ~n28280;
  assign n28284 = ~n33218;
  assign n29019 = ~n32230 | ~n33086;
  assign n28287 = ~n28285 ^ n28565;
  assign n28286 = n33116 & P2_INSTADDRPOINTER_REG_0__SCAN_IN;
  assign n28288 = ~n28287 | ~n28286;
  assign n40322 = ~n28287 ^ n28286;
  assign n28289 = ~n28291;
  assign n28292 = ~n28289 | ~P2_INSTADDRPOINTER_REG_2__SCAN_IN;
  assign n40306 = ~n28290 ^ n28575;
  assign n40305 = P2_INSTADDRPOINTER_REG_2__SCAN_IN ^ n28291;
  assign n40308 = n40306 | n40305;
  assign n28293 = ~n28292 | ~n40308;
  assign n28294 = n28293 | P2_INSTADDRPOINTER_REG_3__SCAN_IN;
  assign n28297 = ~n28296 | ~n28601;
  assign n28302 = ~n32581 | ~n33073;
  assign n28310 = ~n22966 | ~n28309;
  assign n32925 = P2_INSTADDRPOINTER_REG_10__SCAN_IN & P2_INSTADDRPOINTER_REG_9__SCAN_IN;
  assign n32851 = ~n32925 | ~P2_INSTADDRPOINTER_REG_11__SCAN_IN;
  assign n32859 = P2_INSTADDRPOINTER_REG_13__SCAN_IN & P2_INSTADDRPOINTER_REG_12__SCAN_IN;
  assign n32376 = ~n32859 | ~P2_INSTADDRPOINTER_REG_14__SCAN_IN;
  assign n28313 = ~n32376;
  assign n32807 = P2_INSTADDRPOINTER_REG_16__SCAN_IN & P2_INSTADDRPOINTER_REG_15__SCAN_IN;
  assign n29054 = n32807 & P2_INSTADDRPOINTER_REG_17__SCAN_IN;
  assign n28314 = P2_INSTADDRPOINTER_REG_26__SCAN_IN & P2_INSTADDRPOINTER_REG_25__SCAN_IN;
  assign n33220 = ~n28316;
  assign n29017 = ~n32231 & ~n23239;
  assign n28324 = ~n28366 | ~P2_INSTADDRPOINTER_REG_27__SCAN_IN;
  assign n28320 = ~n29843 | ~P2_EBX_REG_27__SCAN_IN;
  assign n28319 = ~P2_PHYADDRPOINTER_REG_27__SCAN_IN | ~P2_STATE2_REG_1__SCAN_IN;
  assign n28322 = ~n28320 | ~n28319;
  assign n42040 = ~P2_REIP_REG_27__SCAN_IN;
  assign n28321 = ~n28476 & ~n42040;
  assign n28323 = ~n28322 & ~n28321;
  assign n28326 = ~n23149 | ~n27734;
  assign n28330 = ~n28326 | ~n28325;
  assign n28329 = ~n28327 | ~n28328;
  assign n28331 = ~n28330 | ~n28329;
  assign n28333 = n28332;
  assign n28334 = ~n28333;
  assign n28336 = n28335 | n28334;
  assign n28343 = ~n28366 | ~P2_INSTADDRPOINTER_REG_4__SCAN_IN;
  assign n28338 = ~n29843 | ~P2_EBX_REG_4__SCAN_IN;
  assign n28337 = ~P2_PHYADDRPOINTER_REG_4__SCAN_IN | ~P2_STATE2_REG_1__SCAN_IN;
  assign n28341 = ~n28338 | ~n28337;
  assign n28339 = ~P2_REIP_REG_4__SCAN_IN;
  assign n28340 = ~n28476 & ~n28339;
  assign n28342 = ~n28341 & ~n28340;
  assign n39580 = n28343 & n28342;
  assign n28351 = ~n28366 | ~P2_INSTADDRPOINTER_REG_5__SCAN_IN;
  assign n28346 = ~n29843 | ~P2_EBX_REG_5__SCAN_IN;
  assign n28345 = ~P2_PHYADDRPOINTER_REG_5__SCAN_IN | ~P2_STATE2_REG_1__SCAN_IN;
  assign n28349 = ~n28346 | ~n28345;
  assign n32586 = ~P2_REIP_REG_5__SCAN_IN;
  assign n28348 = ~n28476 & ~n32586;
  assign n28350 = ~n28349 & ~n28348;
  assign n28358 = ~n28366 | ~P2_INSTADDRPOINTER_REG_6__SCAN_IN;
  assign n28353 = ~n29843 | ~P2_EBX_REG_6__SCAN_IN;
  assign n28352 = ~P2_PHYADDRPOINTER_REG_6__SCAN_IN | ~P2_STATE2_REG_1__SCAN_IN;
  assign n28356 = ~n28353 | ~n28352;
  assign n28354 = ~P2_REIP_REG_6__SCAN_IN;
  assign n28355 = ~n28476 & ~n28354;
  assign n28357 = ~n28356 & ~n28355;
  assign n32563 = ~n28358 | ~n28357;
  assign n28365 = ~n28366 | ~P2_INSTADDRPOINTER_REG_7__SCAN_IN;
  assign n28360 = ~n29843 | ~P2_EBX_REG_7__SCAN_IN;
  assign n28359 = ~P2_PHYADDRPOINTER_REG_7__SCAN_IN | ~P2_STATE2_REG_1__SCAN_IN;
  assign n28363 = ~n28360 | ~n28359;
  assign n28361 = ~P2_REIP_REG_7__SCAN_IN;
  assign n28362 = ~n28476 & ~n28361;
  assign n28364 = ~n28363 & ~n28362;
  assign n28373 = ~n28366 | ~P2_INSTADDRPOINTER_REG_8__SCAN_IN;
  assign n28368 = ~n29843 | ~P2_EBX_REG_8__SCAN_IN;
  assign n28367 = ~P2_PHYADDRPOINTER_REG_8__SCAN_IN | ~P2_STATE2_REG_1__SCAN_IN;
  assign n28371 = ~n28368 | ~n28367;
  assign n28369 = ~P2_REIP_REG_8__SCAN_IN;
  assign n28370 = ~n28476 & ~n28369;
  assign n28372 = ~n28371 & ~n28370;
  assign n28379 = ~n28366 | ~P2_INSTADDRPOINTER_REG_9__SCAN_IN;
  assign n28375 = ~n29843 | ~P2_EBX_REG_9__SCAN_IN;
  assign n28374 = ~P2_PHYADDRPOINTER_REG_9__SCAN_IN | ~P2_STATE2_REG_1__SCAN_IN;
  assign n28377 = ~n28375 | ~n28374;
  assign n32974 = ~P2_REIP_REG_9__SCAN_IN;
  assign n28376 = ~n28476 & ~n32974;
  assign n28378 = ~n28377 & ~n28376;
  assign n32512 = ~n28379 | ~n28378;
  assign n28386 = ~n28366 | ~P2_INSTADDRPOINTER_REG_10__SCAN_IN;
  assign n28381 = ~n29843 | ~P2_EBX_REG_10__SCAN_IN;
  assign n28380 = ~P2_PHYADDRPOINTER_REG_10__SCAN_IN | ~P2_STATE2_REG_1__SCAN_IN;
  assign n28384 = ~n28381 | ~n28380;
  assign n28382 = ~P2_REIP_REG_10__SCAN_IN;
  assign n28383 = ~n28476 & ~n28382;
  assign n28385 = ~n28384 & ~n28383;
  assign n32492 = ~n28386 | ~n28385;
  assign n28393 = ~n28366 | ~P2_INSTADDRPOINTER_REG_11__SCAN_IN;
  assign n28388 = ~n29843 | ~P2_EBX_REG_11__SCAN_IN;
  assign n28387 = ~P2_PHYADDRPOINTER_REG_11__SCAN_IN | ~P2_STATE2_REG_1__SCAN_IN;
  assign n28391 = ~n28388 | ~n28387;
  assign n28389 = ~P2_REIP_REG_11__SCAN_IN;
  assign n28390 = ~n28476 & ~n28389;
  assign n28392 = ~n28391 & ~n28390;
  assign n28400 = ~n28366 | ~P2_INSTADDRPOINTER_REG_12__SCAN_IN;
  assign n28395 = ~n29843 | ~P2_EBX_REG_12__SCAN_IN;
  assign n28394 = ~P2_PHYADDRPOINTER_REG_12__SCAN_IN | ~P2_STATE2_REG_1__SCAN_IN;
  assign n28398 = ~n28395 | ~n28394;
  assign n28396 = ~P2_REIP_REG_12__SCAN_IN;
  assign n28397 = ~n28476 & ~n28396;
  assign n28399 = ~n28398 & ~n28397;
  assign n28407 = ~n28366 | ~P2_INSTADDRPOINTER_REG_13__SCAN_IN;
  assign n28402 = ~n29843 | ~P2_EBX_REG_13__SCAN_IN;
  assign n28401 = ~P2_PHYADDRPOINTER_REG_13__SCAN_IN | ~P2_STATE2_REG_1__SCAN_IN;
  assign n28405 = ~n28402 | ~n28401;
  assign n28403 = ~P2_REIP_REG_13__SCAN_IN;
  assign n28404 = ~n28476 & ~n28403;
  assign n28406 = ~n28405 & ~n28404;
  assign n32440 = ~n28407 | ~n28406;
  assign n28413 = ~n28366 | ~P2_INSTADDRPOINTER_REG_14__SCAN_IN;
  assign n28409 = ~n29843 | ~P2_EBX_REG_14__SCAN_IN;
  assign n28408 = ~P2_PHYADDRPOINTER_REG_14__SCAN_IN | ~P2_STATE2_REG_1__SCAN_IN;
  assign n28411 = ~n28409 | ~n28408;
  assign n32422 = ~P2_REIP_REG_14__SCAN_IN;
  assign n28410 = ~n28476 & ~n32422;
  assign n28412 = ~n28411 & ~n28410;
  assign n32420 = ~n28413 | ~n28412;
  assign n28419 = ~n28366 | ~P2_INSTADDRPOINTER_REG_15__SCAN_IN;
  assign n28415 = ~n29843 | ~P2_EBX_REG_15__SCAN_IN;
  assign n28414 = ~P2_PHYADDRPOINTER_REG_15__SCAN_IN | ~P2_STATE2_REG_1__SCAN_IN;
  assign n28417 = ~n28415 | ~n28414;
  assign n41984 = ~P2_REIP_REG_15__SCAN_IN;
  assign n28416 = ~n28476 & ~n41984;
  assign n28418 = ~n28417 & ~n28416;
  assign n28426 = ~n28366 | ~P2_INSTADDRPOINTER_REG_16__SCAN_IN;
  assign n28421 = ~n29843 | ~P2_EBX_REG_16__SCAN_IN;
  assign n28420 = ~P2_PHYADDRPOINTER_REG_16__SCAN_IN | ~P2_STATE2_REG_1__SCAN_IN;
  assign n28424 = ~n28421 | ~n28420;
  assign n28422 = ~P2_REIP_REG_16__SCAN_IN;
  assign n28423 = ~n28476 & ~n28422;
  assign n28425 = ~n28424 & ~n28423;
  assign n28434 = ~n28366 | ~P2_INSTADDRPOINTER_REG_17__SCAN_IN;
  assign n28429 = ~n29843 | ~P2_EBX_REG_17__SCAN_IN;
  assign n28428 = ~P2_PHYADDRPOINTER_REG_17__SCAN_IN | ~P2_STATE2_REG_1__SCAN_IN;
  assign n28432 = ~n28429 | ~n28428;
  assign n28430 = ~P2_REIP_REG_17__SCAN_IN;
  assign n28431 = ~n28476 & ~n28430;
  assign n28433 = ~n28432 & ~n28431;
  assign n28440 = ~n28366 | ~P2_INSTADDRPOINTER_REG_18__SCAN_IN;
  assign n28436 = ~n29843 | ~P2_EBX_REG_18__SCAN_IN;
  assign n28435 = ~P2_PHYADDRPOINTER_REG_18__SCAN_IN | ~P2_STATE2_REG_1__SCAN_IN;
  assign n28438 = ~n28436 | ~n28435;
  assign n41997 = ~P2_REIP_REG_18__SCAN_IN;
  assign n28437 = ~n28476 & ~n41997;
  assign n28439 = ~n28438 & ~n28437;
  assign n31936 = ~n28440 | ~n28439;
  assign n28447 = ~n28366 | ~P2_INSTADDRPOINTER_REG_19__SCAN_IN;
  assign n28442 = ~n29843 | ~P2_EBX_REG_19__SCAN_IN;
  assign n28441 = ~P2_PHYADDRPOINTER_REG_19__SCAN_IN | ~P2_STATE2_REG_1__SCAN_IN;
  assign n28445 = ~n28442 | ~n28441;
  assign n28443 = ~P2_REIP_REG_19__SCAN_IN;
  assign n28444 = ~n28476 & ~n28443;
  assign n28446 = ~n28445 & ~n28444;
  assign n28454 = ~n28366 | ~P2_INSTADDRPOINTER_REG_20__SCAN_IN;
  assign n28449 = ~n29843 | ~P2_EBX_REG_20__SCAN_IN;
  assign n28448 = ~P2_PHYADDRPOINTER_REG_20__SCAN_IN | ~P2_STATE2_REG_1__SCAN_IN;
  assign n28452 = ~n28449 | ~n28448;
  assign n28450 = ~P2_REIP_REG_20__SCAN_IN;
  assign n28451 = ~n28476 & ~n28450;
  assign n28453 = ~n28452 & ~n28451;
  assign n28461 = ~n28366 | ~P2_INSTADDRPOINTER_REG_21__SCAN_IN;
  assign n28456 = ~n29843 | ~P2_EBX_REG_21__SCAN_IN;
  assign n28455 = ~P2_PHYADDRPOINTER_REG_21__SCAN_IN | ~P2_STATE2_REG_1__SCAN_IN;
  assign n28459 = ~n28456 | ~n28455;
  assign n28457 = ~P2_REIP_REG_21__SCAN_IN;
  assign n28458 = ~n28476 & ~n28457;
  assign n28460 = ~n28459 & ~n28458;
  assign n29072 = ~n28461 | ~n28460;
  assign n28467 = ~n28366 | ~P2_INSTADDRPOINTER_REG_22__SCAN_IN;
  assign n28463 = ~n29843 | ~P2_EBX_REG_22__SCAN_IN;
  assign n28462 = ~P2_PHYADDRPOINTER_REG_22__SCAN_IN | ~P2_STATE2_REG_1__SCAN_IN;
  assign n28465 = ~n28463 | ~n28462;
  assign n32310 = ~P2_REIP_REG_22__SCAN_IN;
  assign n28464 = ~n28476 & ~n32310;
  assign n28466 = ~n28465 & ~n28464;
  assign n28473 = ~n28366 | ~P2_INSTADDRPOINTER_REG_23__SCAN_IN;
  assign n28469 = ~n29843 | ~P2_EBX_REG_23__SCAN_IN;
  assign n28468 = ~P2_PHYADDRPOINTER_REG_23__SCAN_IN | ~P2_STATE2_REG_1__SCAN_IN;
  assign n28471 = ~n28469 | ~n28468;
  assign n42018 = ~P2_REIP_REG_23__SCAN_IN;
  assign n28470 = ~n28476 & ~n42018;
  assign n28472 = ~n28471 & ~n28470;
  assign n28480 = ~n28366 | ~P2_INSTADDRPOINTER_REG_24__SCAN_IN;
  assign n28475 = ~n29843 | ~P2_EBX_REG_24__SCAN_IN;
  assign n28474 = ~P2_PHYADDRPOINTER_REG_24__SCAN_IN | ~P2_STATE2_REG_1__SCAN_IN;
  assign n28478 = ~n28475 | ~n28474;
  assign n42025 = ~P2_REIP_REG_24__SCAN_IN;
  assign n28477 = ~n28476 & ~n42025;
  assign n28479 = ~n28478 & ~n28477;
  assign n31809 = ~n28480 | ~n28479;
  assign n31788 = ~n31810 | ~n31809;
  assign n28486 = ~n28366 | ~P2_INSTADDRPOINTER_REG_25__SCAN_IN;
  assign n28482 = ~n29843 | ~P2_EBX_REG_25__SCAN_IN;
  assign n28481 = ~P2_PHYADDRPOINTER_REG_25__SCAN_IN | ~P2_STATE2_REG_1__SCAN_IN;
  assign n28484 = ~n28482 | ~n28481;
  assign n42030 = ~P2_REIP_REG_25__SCAN_IN;
  assign n28483 = ~n28476 & ~n42030;
  assign n28485 = ~n28484 & ~n28483;
  assign n28492 = ~n28366 | ~P2_INSTADDRPOINTER_REG_26__SCAN_IN;
  assign n28488 = ~n29843 | ~P2_EBX_REG_26__SCAN_IN;
  assign n28487 = ~P2_PHYADDRPOINTER_REG_26__SCAN_IN | ~P2_STATE2_REG_1__SCAN_IN;
  assign n28490 = ~n28488 | ~n28487;
  assign n42035 = ~P2_REIP_REG_26__SCAN_IN;
  assign n28489 = ~n28476 & ~n42035;
  assign n28491 = ~n28490 & ~n28489;
  assign n31785 = ~n28492 | ~n28491;
  assign n33184 = ~n33239 | ~n28493;
  assign n28496 = ~n33184 | ~n42208;
  assign n28495 = ~n33145;
  assign n28497 = ~n28496 | ~n28495;
  assign n28541 = ~n31745 & ~n33125;
  assign n28502 = ~n28499 & ~n28498;
  assign n28501 = ~n28500;
  assign n28504 = ~n28502 | ~n28501;
  assign n28503 = ~n31964;
  assign n28506 = ~n28504 | ~n28503;
  assign n28505 = n27622 | n40501;
  assign n28510 = ~n28506 | ~n28505;
  assign n31968 = ~n28507 | ~n28498;
  assign n28508 = ~n23706 | ~n40444;
  assign n28509 = n31968 & n28508;
  assign n28511 = ~n28510 | ~n28509;
  assign n28517 = ~n28511 & ~n22946;
  assign n28513 = ~n28512 | ~n23085;
  assign n28524 = n28513 & n40456;
  assign n28515 = n28524 | n28514;
  assign n28516 = ~n28515 | ~n40486;
  assign n33143 = ~n28517 | ~n28516;
  assign n32736 = ~n29075 & ~n32752;
  assign n28523 = ~P2_INSTADDRPOINTER_REG_23__SCAN_IN | ~n32736;
  assign n29038 = ~n29054 | ~P2_INSTADDRPOINTER_REG_18__SCAN_IN;
  assign n29043 = ~n32851 & ~n32376;
  assign n28519 = ~n28518 | ~n29043;
  assign n29073 = ~n29038 & ~n28519;
  assign n33015 = ~n33023 & ~n33003;
  assign n28522 = ~P2_INSTADDRPOINTER_REG_8__SCAN_IN | ~n33015;
  assign n33061 = ~P2_INSTADDRPOINTER_REG_1__SCAN_IN | ~P2_INSTADDRPOINTER_REG_0__SCAN_IN;
  assign n40377 = ~n33061;
  assign n33074 = ~P2_INSTADDRPOINTER_REG_3__SCAN_IN | ~P2_INSTADDRPOINTER_REG_4__SCAN_IN;
  assign n33002 = ~n33073 & ~n33074;
  assign n28520 = n40377 & n33002;
  assign n32991 = ~P2_INSTADDRPOINTER_REG_2__SCAN_IN | ~n28520;
  assign n32852 = ~n28522 & ~n32991;
  assign n29074 = ~n29073 | ~n32852;
  assign n32671 = ~n28523 & ~n29074;
  assign n28521 = ~n29869 | ~n32671;
  assign n28531 = ~n33062 | ~n28521;
  assign n28581 = ~P2_INSTADDRPOINTER_REG_2__SCAN_IN;
  assign n33065 = ~n28581 | ~n33061;
  assign n32995 = ~n33065 | ~n33002;
  assign n29050 = ~n32995 & ~n28522;
  assign n29078 = ~n29050 | ~n29073;
  assign n29866 = ~n29078 & ~n28523;
  assign n32673 = ~n29866;
  assign n28533 = ~n29869;
  assign n28536 = ~n32673 & ~n28533;
  assign n33185 = n28524 | n27677;
  assign n28525 = n40456 | n28552;
  assign n28526 = ~n28525 & ~n23706;
  assign n33229 = ~n33185 | ~n28526;
  assign n28527 = ~n33229;
  assign n28529 = ~n28536 & ~n40390;
  assign n28528 = ~n29013;
  assign n40325 = n41785 & n42197;
  assign n33064 = ~n28528 | ~n40294;
  assign n28530 = ~n28529 & ~n40403;
  assign n29873 = ~n28531 | ~n28530;
  assign n32993 = ~n33062;
  assign n28532 = ~P2_INSTADDRPOINTER_REG_27__SCAN_IN & ~n32993;
  assign n32637 = ~n29873 & ~n28532;
  assign n29867 = ~n33062 | ~n32671;
  assign n28534 = ~n28533 & ~n29867;
  assign n28535 = ~P2_INSTADDRPOINTER_REG_27__SCAN_IN & ~n28534;
  assign n28539 = ~n32637 & ~n28535;
  assign n32635 = n32996 & n32222;
  assign n28537 = ~n32635 | ~n28536;
  assign n32236 = ~n40325 | ~P2_REIP_REG_27__SCAN_IN;
  assign n28538 = ~n28537 | ~n32236;
  assign n28540 = n28539 | n28538;
  assign n29015 = ~n28541 & ~n28540;
  assign n28547 = ~n29896 & ~n42040;
  assign n28555 = ~n28543 | ~n42196;
  assign n29897 = ~n29891;
  assign n28545 = ~n29897 | ~P2_INSTADDRPOINTER_REG_27__SCAN_IN;
  assign n29898 = ~n28596;
  assign n28544 = ~n29898 | ~P2_EAX_REG_27__SCAN_IN;
  assign n28546 = ~n28545 | ~n28544;
  assign n29882 = ~n28547 & ~n28546;
  assign n28551 = ~n28580 | ~P2_REIP_REG_1__SCAN_IN;
  assign n28549 = n28555 | n42096;
  assign n40205 = ~P2_EAX_REG_1__SCAN_IN;
  assign n28548 = n22860 | n40205;
  assign n28550 = n28549 & n28548;
  assign n28559 = ~n28955 | ~n28554;
  assign n28566 = n40552 | P2_STATE2_REG_3__SCAN_IN;
  assign n42179 = ~P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & ~n42196;
  assign n28556 = ~n42179;
  assign n28557 = ~n28566 | ~n28556;
  assign n28558 = n28577 & n28557;
  assign n28564 = ~n28580 | ~P2_REIP_REG_0__SCAN_IN;
  assign n28562 = n28555 | n33123;
  assign n28560 = ~n40552 | ~P2_EAX_REG_0__SCAN_IN;
  assign n28561 = n28560 & n42196;
  assign n28563 = n28562 & n28561;
  assign n33113 = ~n28564 | ~n28563;
  assign n28571 = ~n23105 | ~n28565;
  assign n28567 = ~n28566;
  assign n28569 = ~n28567 | ~n39849;
  assign n28568 = ~P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~P2_STATE2_REG_3__SCAN_IN;
  assign n28570 = n28569 & n28568;
  assign n39659 = ~n28571 | ~n28570;
  assign n28574 = ~n28573 | ~n28572;
  assign n28579 = ~n23105 | ~n28575;
  assign n28576 = ~P2_STATE2_REG_3__SCAN_IN | ~P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign n28578 = n28577 & n28576;
  assign n28587 = ~n28579 | ~n28578;
  assign n28585 = ~n28980 | ~P2_REIP_REG_2__SCAN_IN;
  assign n28583 = n29891 | n28581;
  assign n40210 = ~P2_EAX_REG_2__SCAN_IN;
  assign n28582 = n28596 | n40210;
  assign n28584 = n28583 & n28582;
  assign n39626 = n28585 & n28584;
  assign n28590 = ~n39627 | ~n39626;
  assign n28588 = ~n28587;
  assign n28589 = ~n28586 | ~n28588;
  assign n33094 = ~n28590 | ~n28589;
  assign n28594 = ~n28980 | ~P2_REIP_REG_3__SCAN_IN;
  assign n33104 = ~P2_INSTADDRPOINTER_REG_3__SCAN_IN;
  assign n28592 = n29891 | n33104;
  assign n28591 = ~P2_STATE2_REG_3__SCAN_IN | ~P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN;
  assign n28593 = n28592 & n28591;
  assign n28600 = ~n28594 | ~n28593;
  assign n28598 = n23104 | n28595;
  assign n40215 = ~P2_EAX_REG_3__SCAN_IN;
  assign n28597 = n28596 | n40215;
  assign n28599 = ~n28598 | ~n28597;
  assign n33093 = ~n28600 & ~n28599;
  assign n28602 = ~n28601;
  assign n28606 = ~n23105 | ~n28602;
  assign n28604 = n29891 | n40368;
  assign n40220 = ~P2_EAX_REG_4__SCAN_IN;
  assign n28603 = n28596 | n40220;
  assign n28605 = n28604 & n28603;
  assign n28608 = n28606 & n28605;
  assign n28607 = ~n28980 | ~P2_REIP_REG_4__SCAN_IN;
  assign n39587 = n28608 & n28607;
  assign n28613 = ~n23105 | ~n28609;
  assign n28611 = n29891 | n33073;
  assign n40225 = ~P2_EAX_REG_5__SCAN_IN;
  assign n28610 = n28596 | n40225;
  assign n28612 = n28611 & n28610;
  assign n28615 = n28613 & n28612;
  assign n28614 = ~n28980 | ~P2_REIP_REG_5__SCAN_IN;
  assign n33072 = ~n28615 | ~n28614;
  assign n28617 = ~n23105 | ~n28616;
  assign n28621 = n29896 | n28354;
  assign n28619 = n29891 | n33003;
  assign n40231 = ~P2_EAX_REG_6__SCAN_IN;
  assign n28618 = n28596 | n40231;
  assign n28620 = n28619 & n28618;
  assign n33045 = ~n28621 | ~n28620;
  assign n28622 = ~n23105 | ~n29831;
  assign n33026 = ~n28623 | ~n28622;
  assign n28627 = n29896 | n28361;
  assign n28625 = n29891 | n33023;
  assign n40236 = ~P2_EAX_REG_7__SCAN_IN;
  assign n28624 = n28596 | n40236;
  assign n28626 = n28625 & n28624;
  assign n33025 = ~n28627 | ~n28626;
  assign n33027 = ~n33026 | ~n33025;
  assign n28629 = ~n29436 | ~P2_INSTQUEUE_REG_10__0__SCAN_IN;
  assign n28628 = ~n27509 | ~P2_INSTQUEUE_REG_12__0__SCAN_IN;
  assign n28633 = ~n28629 | ~n28628;
  assign n29474 = ~n33147;
  assign n28631 = ~n29474 | ~P2_INSTQUEUE_REG_9__0__SCAN_IN;
  assign n28630 = ~n29597 | ~P2_INSTQUEUE_REG_4__0__SCAN_IN;
  assign n28632 = ~n28631 | ~n28630;
  assign n28646 = ~n28633 & ~n28632;
  assign n28634 = ~P2_INSTQUEUE_REG_15__0__SCAN_IN;
  assign n28638 = ~n23277 & ~n28634;
  assign n28636 = ~n29591 | ~P2_INSTQUEUE_REG_14__0__SCAN_IN;
  assign n28635 = ~n29592 | ~P2_INSTQUEUE_REG_0__0__SCAN_IN;
  assign n28637 = ~n28636 | ~n28635;
  assign n28640 = ~n28638 & ~n28637;
  assign n29469 = ~n29580;
  assign n28639 = ~n29469 | ~P2_INSTQUEUE_REG_3__0__SCAN_IN;
  assign n28644 = ~n28640 | ~n28639;
  assign n29478 = ~n29569;
  assign n28642 = ~n29478 | ~P2_INSTQUEUE_REG_8__0__SCAN_IN;
  assign n29475 = ~n29581;
  assign n28641 = ~n29475 | ~P2_INSTQUEUE_REG_13__0__SCAN_IN;
  assign n28643 = ~n28642 | ~n28641;
  assign n28645 = ~n28644 & ~n28643;
  assign n28649 = ~n29519 | ~P2_INSTQUEUE_REG_2__0__SCAN_IN;
  assign n28648 = n29577 | n28647;
  assign n28654 = ~n28649 | ~n28648;
  assign n28650 = ~P2_INSTQUEUE_REG_11__0__SCAN_IN;
  assign n28652 = n29575 | n28650;
  assign n28651 = ~n29588 | ~P2_INSTQUEUE_REG_1__0__SCAN_IN;
  assign n28653 = ~n28652 | ~n28651;
  assign n28659 = n28654 | n28653;
  assign n28657 = ~n29491 | ~P2_INSTQUEUE_REG_6__0__SCAN_IN;
  assign n28655 = ~P2_INSTQUEUE_REG_5__0__SCAN_IN;
  assign n28656 = n29602 | n28655;
  assign n28658 = ~n28657 | ~n28656;
  assign n28660 = ~n28659 & ~n28658;
  assign n29340 = ~n23970 | ~n28660;
  assign n28667 = ~n29340 | ~n23105;
  assign n28665 = ~n28980 | ~P2_REIP_REG_8__SCAN_IN;
  assign n28663 = n29891 | n23429;
  assign n28661 = ~P2_EAX_REG_8__SCAN_IN;
  assign n28662 = n28596 | n28661;
  assign n28664 = n28663 & n28662;
  assign n28666 = n28665 & n28664;
  assign n33006 = n28667 & n28666;
  assign n28672 = ~n29436 | ~P2_INSTQUEUE_REG_10__1__SCAN_IN;
  assign n28671 = n29569 | n28670;
  assign n28677 = ~n28672 | ~n28671;
  assign n28675 = ~n27817 | ~P2_INSTQUEUE_REG_6__1__SCAN_IN;
  assign n28673 = ~P2_INSTQUEUE_REG_9__1__SCAN_IN;
  assign n28674 = n33147 | n28673;
  assign n28676 = ~n28675 | ~n28674;
  assign n28688 = n28677 | n28676;
  assign n28680 = n29577 | n28678;
  assign n29437 = ~P2_INSTQUEUE_REG_11__1__SCAN_IN;
  assign n28679 = n29575 | n29437;
  assign n28686 = ~n28680 | ~n28679;
  assign n28684 = n29580 | n28681;
  assign n28683 = n29581 | n28682;
  assign n28685 = ~n28684 | ~n28683;
  assign n28687 = n28686 | n28685;
  assign n28706 = ~n28688 & ~n28687;
  assign n28691 = ~n28734 | ~P2_INSTQUEUE_REG_15__1__SCAN_IN;
  assign n28690 = ~n29592 | ~P2_INSTQUEUE_REG_0__1__SCAN_IN;
  assign n28695 = ~n28691 | ~n28690;
  assign n28693 = ~n29591 | ~P2_INSTQUEUE_REG_14__1__SCAN_IN;
  assign n28692 = ~n29588 | ~P2_INSTQUEUE_REG_1__1__SCAN_IN;
  assign n28694 = ~n28693 | ~n28692;
  assign n28699 = ~n28695 & ~n28694;
  assign n28697 = ~n29597 | ~P2_INSTQUEUE_REG_4__1__SCAN_IN;
  assign n28696 = ~n27509 | ~P2_INSTQUEUE_REG_12__1__SCAN_IN;
  assign n28698 = n28697 & n28696;
  assign n28704 = ~n28699 | ~n28698;
  assign n28702 = ~n29519 | ~P2_INSTQUEUE_REG_2__1__SCAN_IN;
  assign n28701 = n29602 | n28700;
  assign n28703 = ~n28702 | ~n28701;
  assign n28705 = ~n28704 & ~n28703;
  assign n39762 = ~n28706 | ~n28705;
  assign n28711 = ~n23105 | ~n39762;
  assign n28709 = n29891 | n32975;
  assign n28707 = ~P2_EAX_REG_9__SCAN_IN;
  assign n28708 = n28596 | n28707;
  assign n28710 = n28709 & n28708;
  assign n28713 = n28711 & n28710;
  assign n28712 = ~n28980 | ~P2_REIP_REG_9__SCAN_IN;
  assign n32971 = n28713 & n28712;
  assign n28716 = ~n27817 | ~P2_INSTQUEUE_REG_6__2__SCAN_IN;
  assign n28715 = ~n29597 | ~P2_INSTQUEUE_REG_4__2__SCAN_IN;
  assign n28720 = ~n28716 | ~n28715;
  assign n28718 = ~n29436 | ~P2_INSTQUEUE_REG_10__2__SCAN_IN;
  assign n28717 = ~n29474 | ~P2_INSTQUEUE_REG_9__2__SCAN_IN;
  assign n28719 = ~n28718 | ~n28717;
  assign n28733 = ~n28720 & ~n28719;
  assign n28721 = ~P2_INSTQUEUE_REG_5__2__SCAN_IN;
  assign n28725 = ~n29602 & ~n28721;
  assign n28723 = ~n29591 | ~P2_INSTQUEUE_REG_14__2__SCAN_IN;
  assign n28722 = ~n29592 | ~P2_INSTQUEUE_REG_0__2__SCAN_IN;
  assign n28724 = ~n28723 | ~n28722;
  assign n28727 = ~n28725 & ~n28724;
  assign n28726 = ~n29519 | ~P2_INSTQUEUE_REG_2__2__SCAN_IN;
  assign n28731 = ~n28727 | ~n28726;
  assign n29466 = ~n29575;
  assign n28729 = ~n29466 | ~P2_INSTQUEUE_REG_11__2__SCAN_IN;
  assign n29465 = ~n29577;
  assign n28728 = ~n29465 | ~P2_INSTQUEUE_REG_7__2__SCAN_IN;
  assign n28730 = ~n28729 | ~n28728;
  assign n28732 = ~n28731 & ~n28730;
  assign n28736 = ~n28734 | ~P2_INSTQUEUE_REG_15__2__SCAN_IN;
  assign n28735 = ~n29588 | ~P2_INSTQUEUE_REG_1__2__SCAN_IN;
  assign n28738 = n28736 & n28735;
  assign n28737 = ~n27509 | ~P2_INSTQUEUE_REG_12__2__SCAN_IN;
  assign n28740 = ~n28738 | ~n28737;
  assign n28739 = ~n29569 & ~n29497;
  assign n28746 = ~n28740 & ~n28739;
  assign n28741 = ~P2_INSTQUEUE_REG_3__2__SCAN_IN;
  assign n28744 = n29580 | n28741;
  assign n28742 = ~P2_INSTQUEUE_REG_13__2__SCAN_IN;
  assign n28743 = n29581 | n28742;
  assign n28745 = n28744 & n28743;
  assign n28747 = n28746 & n28745;
  assign n39736 = ~n23969 | ~n28747;
  assign n28754 = ~n39736 | ~n23105;
  assign n28752 = ~n28980 | ~P2_REIP_REG_10__SCAN_IN;
  assign n28750 = n29891 | n32502;
  assign n28748 = ~P2_EAX_REG_10__SCAN_IN;
  assign n28749 = n28596 | n28748;
  assign n28751 = n28750 & n28749;
  assign n28753 = n28752 & n28751;
  assign n32951 = n28754 & n28753;
  assign n28757 = ~n27817 | ~P2_INSTQUEUE_REG_6__3__SCAN_IN;
  assign n28755 = ~P2_INSTQUEUE_REG_9__3__SCAN_IN;
  assign n28756 = n33147 | n28755;
  assign n28761 = ~n28757 | ~n28756;
  assign n28759 = ~n29355 | ~P2_INSTQUEUE_REG_2__3__SCAN_IN;
  assign n28758 = n29569 | n29283;
  assign n28760 = ~n28759 | ~n28758;
  assign n28773 = n28761 | n28760;
  assign n28762 = ~P2_INSTQUEUE_REG_11__3__SCAN_IN;
  assign n28765 = n29575 | n28762;
  assign n28764 = n29577 | n28763;
  assign n28771 = ~n28765 | ~n28764;
  assign n28769 = n29580 | n28766;
  assign n28768 = n29581 | n28767;
  assign n28770 = ~n28769 | ~n28768;
  assign n28772 = n28771 | n28770;
  assign n28790 = ~n28773 & ~n28772;
  assign n28775 = ~n28734 | ~P2_INSTQUEUE_REG_15__3__SCAN_IN;
  assign n28774 = ~n29588 | ~P2_INSTQUEUE_REG_1__3__SCAN_IN;
  assign n28779 = ~n28775 | ~n28774;
  assign n28777 = ~n29591 | ~P2_INSTQUEUE_REG_14__3__SCAN_IN;
  assign n28776 = ~n29592 | ~P2_INSTQUEUE_REG_0__3__SCAN_IN;
  assign n28778 = ~n28777 | ~n28776;
  assign n28783 = ~n28779 & ~n28778;
  assign n28781 = ~n27509 | ~P2_INSTQUEUE_REG_12__3__SCAN_IN;
  assign n28780 = ~n29597 | ~P2_INSTQUEUE_REG_4__3__SCAN_IN;
  assign n28782 = n28781 & n28780;
  assign n28788 = ~n28783 | ~n28782;
  assign n28786 = ~n29436 | ~P2_INSTQUEUE_REG_10__3__SCAN_IN;
  assign n28784 = ~P2_INSTQUEUE_REG_5__3__SCAN_IN;
  assign n28785 = n29602 | n28784;
  assign n28787 = ~n28786 | ~n28785;
  assign n28789 = ~n28788 & ~n28787;
  assign n39744 = ~n28790 | ~n28789;
  assign n28795 = ~n23105 | ~n39744;
  assign n28793 = n29891 | n32927;
  assign n28791 = ~P2_EAX_REG_11__SCAN_IN;
  assign n28792 = n28596 | n28791;
  assign n28794 = n28793 & n28792;
  assign n28797 = n28795 & n28794;
  assign n28796 = ~n28980 | ~P2_REIP_REG_11__SCAN_IN;
  assign n32933 = ~n28797 | ~n28796;
  assign n28836 = ~n32931;
  assign n28799 = ~n29519 | ~P2_INSTQUEUE_REG_2__4__SCAN_IN;
  assign n28798 = ~n29591 | ~P2_INSTQUEUE_REG_14__4__SCAN_IN;
  assign n28803 = ~n28799 | ~n28798;
  assign n28801 = ~n29474 | ~P2_INSTQUEUE_REG_9__4__SCAN_IN;
  assign n28800 = ~n29588 | ~P2_INSTQUEUE_REG_1__4__SCAN_IN;
  assign n28802 = ~n28801 | ~n28800;
  assign n28811 = ~n28803 & ~n28802;
  assign n28805 = ~n27817 | ~P2_INSTQUEUE_REG_6__4__SCAN_IN;
  assign n28804 = ~n27510 | ~P2_INSTQUEUE_REG_4__4__SCAN_IN;
  assign n28809 = ~n28805 | ~n28804;
  assign n28807 = ~n29478 | ~P2_INSTQUEUE_REG_8__4__SCAN_IN;
  assign n28806 = ~n29475 | ~P2_INSTQUEUE_REG_13__4__SCAN_IN;
  assign n28808 = ~n28807 | ~n28806;
  assign n28810 = ~n28809 & ~n28808;
  assign n28815 = n27509 & P2_INSTQUEUE_REG_12__4__SCAN_IN;
  assign n28813 = ~n28734 | ~P2_INSTQUEUE_REG_15__4__SCAN_IN;
  assign n28812 = ~n29592 | ~P2_INSTQUEUE_REG_0__4__SCAN_IN;
  assign n28814 = ~n28813 | ~n28812;
  assign n28817 = ~n28815 & ~n28814;
  assign n28816 = ~n29436 | ~P2_INSTQUEUE_REG_10__4__SCAN_IN;
  assign n28826 = ~n28817 | ~n28816;
  assign n29125 = ~P2_INSTQUEUE_REG_11__4__SCAN_IN;
  assign n28819 = n29575 | n29125;
  assign n28818 = n29577 | n29447;
  assign n28824 = ~n28819 | ~n28818;
  assign n29449 = ~P2_INSTQUEUE_REG_3__4__SCAN_IN;
  assign n28822 = n29580 | n29449;
  assign n28820 = ~P2_INSTQUEUE_REG_5__4__SCAN_IN;
  assign n28821 = n29602 | n28820;
  assign n28823 = ~n28822 | ~n28821;
  assign n28825 = n28824 | n28823;
  assign n28827 = ~n28826 & ~n28825;
  assign n39737 = ~n23963 | ~n28827;
  assign n28834 = ~n39737 | ~n23105;
  assign n28832 = ~n28980 | ~P2_REIP_REG_12__SCAN_IN;
  assign n28830 = n29891 | n32899;
  assign n28828 = ~P2_EAX_REG_12__SCAN_IN;
  assign n28829 = n28596 | n28828;
  assign n28831 = n28830 & n28829;
  assign n28833 = n28832 & n28831;
  assign n32902 = n28834 & n28833;
  assign n28838 = ~n29491 | ~P2_INSTQUEUE_REG_6__5__SCAN_IN;
  assign n28837 = ~n29436 | ~P2_INSTQUEUE_REG_10__5__SCAN_IN;
  assign n28844 = ~n28838 | ~n28837;
  assign n28839 = ~P2_INSTQUEUE_REG_9__5__SCAN_IN;
  assign n28842 = n33147 | n28839;
  assign n28841 = n29602 | n28840;
  assign n28843 = ~n28842 | ~n28841;
  assign n28854 = n28844 | n28843;
  assign n28848 = n29577 | n28845;
  assign n28846 = ~P2_INSTQUEUE_REG_11__5__SCAN_IN;
  assign n28847 = n29575 | n28846;
  assign n28852 = ~n28848 | ~n28847;
  assign n28850 = n29580 | n29356;
  assign n28849 = n29569 | n29669;
  assign n28851 = ~n28850 | ~n28849;
  assign n28853 = n28852 | n28851;
  assign n28871 = ~n28854 & ~n28853;
  assign n28856 = ~n28734 | ~P2_INSTQUEUE_REG_15__5__SCAN_IN;
  assign n28855 = ~n29592 | ~P2_INSTQUEUE_REG_0__5__SCAN_IN;
  assign n28860 = ~n28856 | ~n28855;
  assign n28858 = ~n29591 | ~P2_INSTQUEUE_REG_14__5__SCAN_IN;
  assign n28857 = ~n29588 | ~P2_INSTQUEUE_REG_1__5__SCAN_IN;
  assign n28859 = ~n28858 | ~n28857;
  assign n28864 = ~n28860 & ~n28859;
  assign n28862 = ~n29597 | ~P2_INSTQUEUE_REG_4__5__SCAN_IN;
  assign n28861 = ~n27509 | ~P2_INSTQUEUE_REG_12__5__SCAN_IN;
  assign n28863 = n28862 & n28861;
  assign n28869 = ~n28864 | ~n28863;
  assign n28867 = ~n29519 | ~P2_INSTQUEUE_REG_2__5__SCAN_IN;
  assign n28866 = n29581 | n28865;
  assign n28868 = ~n28867 | ~n28866;
  assign n28870 = ~n28869 & ~n28868;
  assign n29343 = ~n28871 | ~n28870;
  assign n28876 = ~n23105 | ~n29343;
  assign n28874 = n29891 | n32849;
  assign n28872 = ~P2_EAX_REG_13__SCAN_IN;
  assign n28873 = n28596 | n28872;
  assign n28875 = n28874 & n28873;
  assign n28878 = n28876 & n28875;
  assign n28877 = ~n28980 | ~P2_REIP_REG_13__SCAN_IN;
  assign n28881 = ~n29475 | ~P2_INSTQUEUE_REG_13__6__SCAN_IN;
  assign n28880 = ~n27509 | ~P2_INSTQUEUE_REG_12__6__SCAN_IN;
  assign n28885 = ~n28881 | ~n28880;
  assign n28883 = ~n29466 | ~P2_INSTQUEUE_REG_11__6__SCAN_IN;
  assign n28882 = ~n27817 | ~P2_INSTQUEUE_REG_6__6__SCAN_IN;
  assign n28884 = ~n28883 | ~n28882;
  assign n28897 = ~n28885 & ~n28884;
  assign n29568 = ~P2_INSTQUEUE_REG_9__6__SCAN_IN;
  assign n28889 = ~n33147 & ~n29568;
  assign n28887 = ~n29591 | ~P2_INSTQUEUE_REG_14__6__SCAN_IN;
  assign n28886 = ~n29588 | ~P2_INSTQUEUE_REG_1__6__SCAN_IN;
  assign n28888 = ~n28887 | ~n28886;
  assign n28891 = ~n28889 & ~n28888;
  assign n28890 = ~n29519 | ~P2_INSTQUEUE_REG_2__6__SCAN_IN;
  assign n28895 = ~n28891 | ~n28890;
  assign n28893 = ~n29465 | ~P2_INSTQUEUE_REG_7__6__SCAN_IN;
  assign n28892 = ~n29478 | ~P2_INSTQUEUE_REG_8__6__SCAN_IN;
  assign n28894 = ~n28893 | ~n28892;
  assign n28896 = ~n28895 & ~n28894;
  assign n28911 = n28897 & n28896;
  assign n28901 = n29597 & P2_INSTQUEUE_REG_4__6__SCAN_IN;
  assign n28899 = ~n28734 | ~P2_INSTQUEUE_REG_15__6__SCAN_IN;
  assign n28898 = ~n29592 | ~P2_INSTQUEUE_REG_0__6__SCAN_IN;
  assign n28900 = ~n28899 | ~n28898;
  assign n28903 = ~n28901 & ~n28900;
  assign n28902 = ~n29436 | ~P2_INSTQUEUE_REG_10__6__SCAN_IN;
  assign n28909 = ~n28903 | ~n28902;
  assign n28907 = n29580 | n28904;
  assign n28906 = n29602 | n28905;
  assign n28908 = ~n28907 | ~n28906;
  assign n28910 = ~n28909 & ~n28908;
  assign n39717 = ~n28911 | ~n28910;
  assign n28918 = ~n39717 | ~n23105;
  assign n28916 = ~n28980 | ~P2_REIP_REG_14__SCAN_IN;
  assign n28914 = n29891 | n32858;
  assign n28912 = ~P2_EAX_REG_14__SCAN_IN;
  assign n28913 = n28596 | n28912;
  assign n28915 = n28914 & n28913;
  assign n28917 = n28916 & n28915;
  assign n32863 = n28918 & n28917;
  assign n28920 = ~n27817 | ~P2_INSTQUEUE_REG_6__7__SCAN_IN;
  assign n28919 = ~n29519 | ~P2_INSTQUEUE_REG_2__7__SCAN_IN;
  assign n28926 = ~n28920 | ~n28919;
  assign n28921 = ~P2_INSTQUEUE_REG_9__7__SCAN_IN;
  assign n28924 = n33147 | n28921;
  assign n28922 = ~P2_INSTQUEUE_REG_13__7__SCAN_IN;
  assign n28923 = n29581 | n28922;
  assign n28925 = ~n28924 | ~n28923;
  assign n28937 = n28926 | n28925;
  assign n28927 = ~P2_INSTQUEUE_REG_11__7__SCAN_IN;
  assign n28930 = n29575 | n28927;
  assign n28929 = n29577 | n28928;
  assign n28935 = ~n28930 | ~n28929;
  assign n28933 = ~n29436 | ~P2_INSTQUEUE_REG_10__7__SCAN_IN;
  assign n28931 = ~P2_INSTQUEUE_REG_3__7__SCAN_IN;
  assign n28932 = n29580 | n28931;
  assign n28934 = ~n28933 | ~n28932;
  assign n28936 = n28935 | n28934;
  assign n28954 = ~n28937 & ~n28936;
  assign n28939 = ~n28734 | ~P2_INSTQUEUE_REG_15__7__SCAN_IN;
  assign n28938 = ~n29588 | ~P2_INSTQUEUE_REG_1__7__SCAN_IN;
  assign n28943 = ~n28939 | ~n28938;
  assign n28941 = ~n29591 | ~P2_INSTQUEUE_REG_14__7__SCAN_IN;
  assign n28940 = ~n29592 | ~P2_INSTQUEUE_REG_0__7__SCAN_IN;
  assign n28942 = ~n28941 | ~n28940;
  assign n28947 = ~n28943 & ~n28942;
  assign n28945 = ~n29597 | ~P2_INSTQUEUE_REG_4__7__SCAN_IN;
  assign n28944 = ~n27509 | ~P2_INSTQUEUE_REG_12__7__SCAN_IN;
  assign n28946 = n28945 & n28944;
  assign n28952 = ~n28947 | ~n28946;
  assign n28948 = ~P2_INSTQUEUE_REG_5__7__SCAN_IN;
  assign n28950 = n29602 | n28948;
  assign n28949 = n29569 | n29749;
  assign n28951 = ~n28950 | ~n28949;
  assign n28953 = ~n28952 & ~n28951;
  assign n29609 = ~n28954 | ~n28953;
  assign n28960 = ~n23105 | ~n29609;
  assign n28958 = n29891 | n32831;
  assign n28956 = ~P2_EAX_REG_15__SCAN_IN;
  assign n28957 = n28596 | n28956;
  assign n28959 = n28958 & n28957;
  assign n28962 = n28960 & n28959;
  assign n28961 = ~n28980 | ~P2_REIP_REG_15__SCAN_IN;
  assign n32835 = ~n28962 | ~n28961;
  assign n28966 = ~n28980 | ~P2_REIP_REG_16__SCAN_IN;
  assign n32818 = ~P2_INSTADDRPOINTER_REG_16__SCAN_IN;
  assign n28964 = n29891 | n32818;
  assign n40118 = ~P2_EAX_REG_16__SCAN_IN;
  assign n28963 = n28596 | n40118;
  assign n28965 = n28964 & n28963;
  assign n28971 = n29896 | n28430;
  assign n28969 = n29891 | n32808;
  assign n40123 = ~P2_EAX_REG_17__SCAN_IN;
  assign n28968 = n28596 | n40123;
  assign n28970 = n28969 & n28968;
  assign n28975 = n29896 | n41997;
  assign n28973 = n29891 | n32362;
  assign n40128 = ~P2_EAX_REG_18__SCAN_IN;
  assign n28972 = n28596 | n40128;
  assign n28974 = n28973 & n28972;
  assign n32151 = ~n28975 | ~n28974;
  assign n28979 = n29896 | n28443;
  assign n28977 = n29891 | n32771;
  assign n40133 = ~P2_EAX_REG_19__SCAN_IN;
  assign n28976 = n28596 | n40133;
  assign n28978 = n28977 & n28976;
  assign n32136 = ~n28979 | ~n28978;
  assign n29033 = ~n32153 | ~n32136;
  assign n28984 = ~n28980 | ~P2_REIP_REG_20__SCAN_IN;
  assign n28982 = n29891 | n29062;
  assign n40138 = ~P2_EAX_REG_20__SCAN_IN;
  assign n28981 = n28596 | n40138;
  assign n28983 = n28982 & n28981;
  assign n28988 = n29896 | n28457;
  assign n28986 = n29891 | n29075;
  assign n40143 = ~P2_EAX_REG_21__SCAN_IN;
  assign n28985 = n28596 | n40143;
  assign n28987 = n28986 & n28985;
  assign n28992 = n29896 | n32310;
  assign n28990 = n29891 | n32752;
  assign n40148 = ~P2_EAX_REG_22__SCAN_IN;
  assign n28989 = n28596 | n40148;
  assign n28991 = n28990 & n28989;
  assign n32089 = ~n28992 | ~n28991;
  assign n28997 = ~n28980 | ~P2_REIP_REG_23__SCAN_IN;
  assign n28995 = n29891 | n28993;
  assign n40153 = ~P2_EAX_REG_23__SCAN_IN;
  assign n28994 = n28596 | n40153;
  assign n28996 = n28995 & n28994;
  assign n31844 = ~n28997 | ~n28996;
  assign n29001 = ~n28980 | ~P2_REIP_REG_24__SCAN_IN;
  assign n28999 = n29891 | n32712;
  assign n40158 = ~P2_EAX_REG_24__SCAN_IN;
  assign n28998 = n28596 | n40158;
  assign n29000 = n28999 & n28998;
  assign n31805 = ~n29002;
  assign n29006 = n29896 | n42030;
  assign n29004 = n29891 | n23751;
  assign n40164 = ~P2_EAX_REG_25__SCAN_IN;
  assign n29003 = n28596 | n40164;
  assign n29005 = n29004 & n29003;
  assign n31765 = ~n31805 & ~n31806;
  assign n29010 = ~n28980 | ~P2_REIP_REG_26__SCAN_IN;
  assign n32245 = ~P2_INSTADDRPOINTER_REG_26__SCAN_IN;
  assign n29008 = ~n29891 & ~n32245;
  assign n40170 = ~P2_EAX_REG_26__SCAN_IN;
  assign n29007 = ~n28596 & ~n40170;
  assign n29009 = ~n29008 & ~n29007;
  assign n31764 = ~n29010 | ~n29009;
  assign n31763 = ~n31765 | ~n31764;
  assign n32015 = n29882 ^ n31763;
  assign n29011 = ~n33223 | ~n40456;
  assign n29012 = ~n29011 | ~n33230;
  assign n29014 = ~n32015 | ~n33115;
  assign n29016 = ~n29015 | ~n29014;
  assign n29018 = ~n29017 & ~n29016;
  assign P2_U3019 = ~n29019 | ~n29018;
  assign n29023 = ~n29022;
  assign n29064 = ~n29026 | ~n29025;
  assign n29027 = ~n29063 | ~n29064;
  assign n29030 = ~n29028 | ~n29062;
  assign n32333 = ~n29030 | ~n29029;
  assign n29059 = ~n32333 & ~n23239;
  assign n39267 = n29031 ^ n22925;
  assign n31917 = ~n39267;
  assign n29037 = ~n31917 & ~n33125;
  assign n29034 = ~n29033 | ~n29032;
  assign n39248 = n29086 & n29034;
  assign n29035 = ~n39248 | ~n33115;
  assign n32335 = ~n40325 | ~P2_REIP_REG_20__SCAN_IN;
  assign n29036 = ~n29035 | ~n32335;
  assign n29049 = ~n29037 & ~n29036;
  assign n29041 = ~n29054 & ~n40390;
  assign n32800 = ~n29043 | ~n32852;
  assign n29039 = ~n29038 & ~n32800;
  assign n29040 = ~n32993 & ~n29039;
  assign n29046 = ~n29041 & ~n29040;
  assign n29042 = n40390 | n29050;
  assign n32921 = ~n29042 | ~n33064;
  assign n29044 = ~n29043;
  assign n29045 = n32996 & n29044;
  assign n32803 = ~n32921 & ~n29045;
  assign n32784 = ~n29046 | ~n32803;
  assign n29047 = n32996 & n32362;
  assign n32772 = n32784 | n29047;
  assign n29048 = ~n32772 | ~P2_INSTADDRPOINTER_REG_20__SCAN_IN;
  assign n29057 = n29049 & n29048;
  assign n29055 = P2_INSTADDRPOINTER_REG_19__SCAN_IN ^ P2_INSTADDRPOINTER_REG_20__SCAN_IN;
  assign n29052 = ~n32852 | ~n33062;
  assign n29051 = ~n29050 | ~n32996;
  assign n32969 = ~n29052 | ~n29051;
  assign n32861 = ~n32969 | ~n29053;
  assign n32830 = ~n32861 & ~n32376;
  assign n32791 = ~n29054 | ~n32830;
  assign n32770 = ~n32362 & ~n32791;
  assign n29056 = ~n29055 | ~n32770;
  assign n29058 = ~n29057 | ~n29056;
  assign n29060 = ~n29059 & ~n29058;
  assign P2_U3026 = ~n29061 | ~n29060;
  assign n29065 = ~n29063 | ~n29062;
  assign n29069 = ~n29065 | ~n29064;
  assign n29068 = ~n29067 & ~n29066;
  assign n29091 = ~n32321 & ~n23239;
  assign n39230 = n29072 ^ n29071;
  assign n29085 = ~n39230 | ~n40408;
  assign n32734 = ~n29073 | ~n32969;
  assign n29083 = ~P2_INSTADDRPOINTER_REG_21__SCAN_IN & ~n32734;
  assign n29076 = ~n29075 & ~n29074;
  assign n29077 = ~n32993 & ~n29076;
  assign n29080 = ~n40403 & ~n29077;
  assign n29079 = ~n32996 | ~n29078;
  assign n32732 = ~n29080 | ~n29079;
  assign n29081 = ~n32732 | ~P2_INSTADDRPOINTER_REG_21__SCAN_IN;
  assign n32324 = ~n40325 | ~P2_REIP_REG_21__SCAN_IN;
  assign n29082 = ~n29081 | ~n32324;
  assign n29084 = ~n29083 & ~n29082;
  assign n29089 = n29085 & n29084;
  assign n32105 = n29087 ^ n29086;
  assign n29088 = ~n32105 | ~n33115;
  assign n29090 = ~n29089 | ~n29088;
  assign n29092 = ~n29091 & ~n29090;
  assign P2_U3025 = ~n29093 | ~n29092;
  assign n29095 = n29094;
  assign n29757 = ~n29095;
  assign n29097 = ~n29757 | ~P2_INSTQUEUE_REG_5__4__SCAN_IN;
  assign n29756 = ~n23571;
  assign n29096 = ~n29756 | ~P2_INSTQUEUE_REG_3__4__SCAN_IN;
  assign n29110 = ~n29097 | ~n29096;
  assign n29100 = ~n27348 | ~n29098;
  assign n29102 = ~n29753 | ~P2_INSTQUEUE_REG_1__4__SCAN_IN;
  assign n29101 = ~n29760 | ~P2_INSTQUEUE_REG_2__4__SCAN_IN;
  assign n29107 = ~n29102 | ~n29101;
  assign n29105 = ~n29761 | ~P2_INSTQUEUE_REG_6__4__SCAN_IN;
  assign n29104 = ~n23145 | ~P2_INSTQUEUE_REG_7__4__SCAN_IN;
  assign n29106 = ~n29105 | ~n29104;
  assign n29108 = ~n29107 & ~n29106;
  assign n29109 = ~n29713 | ~n29108;
  assign n29115 = n29110 | n29109;
  assign n29113 = n29718 | n29111;
  assign n29112 = n27418 | n40497;
  assign n29114 = ~n29113 | ~n29112;
  assign n29137 = n29115 | n29114;
  assign n29119 = n27418 | n29116;
  assign n29117 = ~P2_INSTQUEUE_REG_14__4__SCAN_IN;
  assign n29118 = n29731 | n29117;
  assign n29135 = n29119 & n29118;
  assign n29121 = ~n29752 | ~P2_INSTQUEUE_REG_12__4__SCAN_IN;
  assign n29120 = ~n23145 | ~P2_INSTQUEUE_REG_15__4__SCAN_IN;
  assign n29132 = ~n29121 | ~n29120;
  assign n29122 = ~P2_INSTQUEUE_REG_13__4__SCAN_IN;
  assign n29123 = ~n29095 & ~n29122;
  assign n29130 = ~n29124 & ~n29123;
  assign n29128 = ~n23571 & ~n29125;
  assign n29127 = ~n29688 & ~n29126;
  assign n29129 = ~n29128 & ~n29127;
  assign n29131 = ~n29130 | ~n29129;
  assign n29133 = n29132 | n29131;
  assign n29134 = ~n29713 & ~n29133;
  assign n29136 = ~n29135 | ~n29134;
  assign n29680 = ~n29137 | ~n29136;
  assign n29139 = ~n29591 | ~P2_INSTQUEUE_REG_15__7__SCAN_IN;
  assign n29138 = ~n29588 | ~P2_INSTQUEUE_REG_2__7__SCAN_IN;
  assign n29143 = ~n29139 | ~n29138;
  assign n29141 = ~n29469 | ~P2_INSTQUEUE_REG_4__7__SCAN_IN;
  assign n29140 = ~n29597 | ~P2_INSTQUEUE_REG_5__7__SCAN_IN;
  assign n29142 = ~n29141 | ~n29140;
  assign n29151 = ~n29143 & ~n29142;
  assign n29145 = ~n28734 | ~P2_INSTQUEUE_REG_0__7__SCAN_IN;
  assign n29144 = ~n29592 | ~P2_INSTQUEUE_REG_1__7__SCAN_IN;
  assign n29149 = ~n29145 | ~n29144;
  assign n29147 = ~n29519 | ~P2_INSTQUEUE_REG_3__7__SCAN_IN;
  assign n29479 = ~n29602;
  assign n29146 = ~n29479 | ~P2_INSTQUEUE_REG_6__7__SCAN_IN;
  assign n29148 = ~n29147 | ~n29146;
  assign n29150 = ~n29149 & ~n29148;
  assign n29167 = n29151 & n29150;
  assign n29153 = ~n29465 | ~P2_INSTQUEUE_REG_8__7__SCAN_IN;
  assign n29152 = ~n29475 | ~P2_INSTQUEUE_REG_14__7__SCAN_IN;
  assign n29157 = ~n29153 | ~n29152;
  assign n29155 = ~n29436 | ~P2_INSTQUEUE_REG_11__7__SCAN_IN;
  assign n29154 = ~n27509 | ~P2_INSTQUEUE_REG_13__7__SCAN_IN;
  assign n29156 = ~n29155 | ~n29154;
  assign n29165 = ~n29157 & ~n29156;
  assign n29159 = ~n27817 | ~P2_INSTQUEUE_REG_7__7__SCAN_IN;
  assign n29158 = ~n29474 | ~P2_INSTQUEUE_REG_10__7__SCAN_IN;
  assign n29163 = ~n29159 | ~n29158;
  assign n29161 = ~n29466 | ~P2_INSTQUEUE_REG_12__7__SCAN_IN;
  assign n29160 = ~n29478 | ~P2_INSTQUEUE_REG_9__7__SCAN_IN;
  assign n29162 = ~n29161 | ~n29160;
  assign n29164 = ~n29163 & ~n29162;
  assign n29166 = n29165 & n29164;
  assign n29618 = ~n29167 | ~n29166;
  assign n29169 = ~n29753 | ~P2_INSTQUEUE_REG_9__0__SCAN_IN;
  assign n29168 = ~n29757 | ~P2_INSTQUEUE_REG_13__0__SCAN_IN;
  assign n29178 = ~n29169 | ~n29168;
  assign n29170 = ~n29761 | ~P2_INSTQUEUE_REG_14__0__SCAN_IN;
  assign n29175 = ~n29171 | ~n29170;
  assign n29173 = ~n29739 | ~P2_INSTQUEUE_REG_8__0__SCAN_IN;
  assign n29172 = ~n23145 | ~P2_INSTQUEUE_REG_15__0__SCAN_IN;
  assign n29174 = ~n29173 | ~n29172;
  assign n29176 = ~n29175 & ~n29174;
  assign n29177 = ~n29767 | ~n29176;
  assign n29182 = ~n29178 & ~n29177;
  assign n29180 = n29718 | n29537;
  assign n29760 = ~n29688;
  assign n29179 = ~n29760 | ~P2_INSTQUEUE_REG_10__0__SCAN_IN;
  assign n29181 = n29180 & n29179;
  assign n29199 = ~n29182 | ~n29181;
  assign n29184 = ~n29753 | ~P2_INSTQUEUE_REG_1__0__SCAN_IN;
  assign n29183 = n29718 | n29540;
  assign n29193 = ~n29184 | ~n29183;
  assign n29186 = ~n29660 | ~P2_INSTQUEUE_REG_5__0__SCAN_IN;
  assign n29185 = ~n23145 | ~P2_INSTQUEUE_REG_7__0__SCAN_IN;
  assign n29190 = ~n29186 | ~n29185;
  assign n29187 = ~n29761 | ~P2_INSTQUEUE_REG_6__0__SCAN_IN;
  assign n29189 = ~n29188 | ~n29187;
  assign n29191 = ~n29190 & ~n29189;
  assign n29192 = ~n29713 | ~n29191;
  assign n29197 = ~n29193 & ~n29192;
  assign n29195 = n27418 | n40428;
  assign n29194 = ~n29760 | ~P2_INSTQUEUE_REG_2__0__SCAN_IN;
  assign n29196 = n29195 & n29194;
  assign n29198 = ~n29197 | ~n29196;
  assign n29619 = n29199 & n29198;
  assign n29621 = ~n29618 | ~n29619;
  assign n29200 = ~P2_INSTQUEUE_REG_15__1__SCAN_IN;
  assign n29203 = ~n29103 & ~n29200;
  assign n29201 = ~n29739 | ~P2_INSTQUEUE_REG_8__1__SCAN_IN;
  assign n29202 = ~n29201 | ~n29767;
  assign n29211 = ~n29203 & ~n29202;
  assign n29205 = ~n29660 | ~P2_INSTQUEUE_REG_13__1__SCAN_IN;
  assign n29204 = ~n29760 | ~P2_INSTQUEUE_REG_10__1__SCAN_IN;
  assign n29209 = ~n29205 | ~n29204;
  assign n29207 = ~n29752 | ~P2_INSTQUEUE_REG_12__1__SCAN_IN;
  assign n29206 = ~n29761 | ~P2_INSTQUEUE_REG_14__1__SCAN_IN;
  assign n29208 = ~n29207 | ~n29206;
  assign n29210 = ~n29209 & ~n29208;
  assign n29215 = ~n29211 | ~n29210;
  assign n29213 = ~n29753 | ~P2_INSTQUEUE_REG_9__1__SCAN_IN;
  assign n29212 = ~n29756 | ~P2_INSTQUEUE_REG_11__1__SCAN_IN;
  assign n29214 = ~n29213 | ~n29212;
  assign n29234 = n29215 | n29214;
  assign n29217 = ~n29753 | ~P2_INSTQUEUE_REG_1__1__SCAN_IN;
  assign n29216 = ~n29757 | ~P2_INSTQUEUE_REG_5__1__SCAN_IN;
  assign n29221 = ~n29217 | ~n29216;
  assign n29219 = ~n29756 | ~P2_INSTQUEUE_REG_3__1__SCAN_IN;
  assign n29218 = ~n29760 | ~P2_INSTQUEUE_REG_2__1__SCAN_IN;
  assign n29220 = ~n29219 | ~n29218;
  assign n29232 = ~n29221 & ~n29220;
  assign n29223 = n29731 | n29222;
  assign n29225 = n29223 & n29713;
  assign n29224 = ~n23145 | ~P2_INSTQUEUE_REG_7__1__SCAN_IN;
  assign n29230 = ~n29225 | ~n29224;
  assign n29228 = n29718 | n29226;
  assign n29227 = n27418 | n40452;
  assign n29229 = ~n29228 | ~n29227;
  assign n29231 = ~n29230 & ~n29229;
  assign n29233 = ~n29232 | ~n29231;
  assign n29625 = ~n29234 | ~n29233;
  assign n29624 = ~n29621 & ~n29625;
  assign n29628 = ~n29624;
  assign n29236 = ~n29753 | ~P2_INSTQUEUE_REG_9__2__SCAN_IN;
  assign n29235 = ~n29757 | ~P2_INSTQUEUE_REG_13__2__SCAN_IN;
  assign n29245 = ~n29236 | ~n29235;
  assign n29238 = ~n29761 | ~P2_INSTQUEUE_REG_14__2__SCAN_IN;
  assign n29237 = ~n23145 | ~P2_INSTQUEUE_REG_15__2__SCAN_IN;
  assign n29242 = ~n29238 | ~n29237;
  assign n29240 = ~n29752 | ~P2_INSTQUEUE_REG_12__2__SCAN_IN;
  assign n29239 = ~n29739 | ~P2_INSTQUEUE_REG_8__2__SCAN_IN;
  assign n29241 = ~n29240 | ~n29239;
  assign n29243 = ~n29242 & ~n29241;
  assign n29244 = ~n29767 | ~n29243;
  assign n29249 = ~n29245 & ~n29244;
  assign n29247 = ~n29756 | ~P2_INSTQUEUE_REG_11__2__SCAN_IN;
  assign n29246 = ~n29760 | ~P2_INSTQUEUE_REG_10__2__SCAN_IN;
  assign n29248 = n29247 & n29246;
  assign n29266 = ~n29249 | ~n29248;
  assign n29251 = n29718 | n29501;
  assign n29250 = ~n29756 | ~P2_INSTQUEUE_REG_3__2__SCAN_IN;
  assign n29260 = ~n29251 | ~n29250;
  assign n29253 = ~n29660 | ~P2_INSTQUEUE_REG_5__2__SCAN_IN;
  assign n29252 = ~n29761 | ~P2_INSTQUEUE_REG_6__2__SCAN_IN;
  assign n29257 = ~n29253 | ~n29252;
  assign n29255 = ~n29753 | ~P2_INSTQUEUE_REG_1__2__SCAN_IN;
  assign n29254 = ~n23145 | ~P2_INSTQUEUE_REG_7__2__SCAN_IN;
  assign n29256 = ~n29255 | ~n29254;
  assign n29258 = ~n29257 & ~n29256;
  assign n29259 = ~n29713 | ~n29258;
  assign n29264 = ~n29260 & ~n29259;
  assign n29262 = n27418 | n40467;
  assign n29261 = ~n29760 | ~P2_INSTQUEUE_REG_2__2__SCAN_IN;
  assign n29263 = n29262 & n29261;
  assign n29265 = ~n29264 | ~n29263;
  assign n29627 = n29266 & n29265;
  assign n29630 = ~n29627;
  assign n29631 = ~n29628 & ~n29630;
  assign n29267 = ~n29761 | ~P2_INSTQUEUE_REG_6__3__SCAN_IN;
  assign n29269 = ~n29267 | ~n29713;
  assign n29268 = ~n27418 & ~n40482;
  assign n29277 = ~n29269 & ~n29268;
  assign n29271 = ~n29753 | ~P2_INSTQUEUE_REG_1__3__SCAN_IN;
  assign n29270 = ~n29660 | ~P2_INSTQUEUE_REG_5__3__SCAN_IN;
  assign n29275 = ~n29271 | ~n29270;
  assign n29273 = ~n29756 | ~P2_INSTQUEUE_REG_3__3__SCAN_IN;
  assign n29272 = ~n23145 | ~P2_INSTQUEUE_REG_7__3__SCAN_IN;
  assign n29274 = ~n29273 | ~n29272;
  assign n29276 = ~n29275 & ~n29274;
  assign n29282 = ~n29277 | ~n29276;
  assign n29280 = n29718 | n29278;
  assign n29279 = ~n29760 | ~P2_INSTQUEUE_REG_2__3__SCAN_IN;
  assign n29281 = ~n29280 | ~n29279;
  assign n29300 = n29282 | n29281;
  assign n29286 = ~n27418 & ~n29283;
  assign n29284 = ~n29760 | ~P2_INSTQUEUE_REG_10__3__SCAN_IN;
  assign n29285 = ~n29284 | ~n29767;
  assign n29294 = ~n29286 & ~n29285;
  assign n29288 = ~n29752 | ~P2_INSTQUEUE_REG_12__3__SCAN_IN;
  assign n29287 = ~n23145 | ~P2_INSTQUEUE_REG_15__3__SCAN_IN;
  assign n29292 = ~n29288 | ~n29287;
  assign n29290 = ~n29753 | ~P2_INSTQUEUE_REG_9__3__SCAN_IN;
  assign n29289 = ~n29756 | ~P2_INSTQUEUE_REG_11__3__SCAN_IN;
  assign n29291 = ~n29290 | ~n29289;
  assign n29293 = ~n29292 & ~n29291;
  assign n29298 = ~n29294 | ~n29293;
  assign n29296 = ~n29757 | ~P2_INSTQUEUE_REG_13__3__SCAN_IN;
  assign n29403 = ~P2_INSTQUEUE_REG_14__3__SCAN_IN;
  assign n29295 = n29731 | n29403;
  assign n29297 = ~n29296 | ~n29295;
  assign n29299 = n29298 | n29297;
  assign n29637 = ~n29300 | ~n29299;
  assign n29301 = ~n29637;
  assign n29681 = ~n29636;
  assign n29303 = n29680 ^ n29681;
  assign n29302 = ~n40456 | ~P2_STATE2_REG_0__SCAN_IN;
  assign n29312 = ~n33144 | ~n23278;
  assign n29310 = ~n29320 | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n41089 = ~n40991 | ~P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN;
  assign n29308 = ~n41158;
  assign n40648 = ~P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & ~P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN;
  assign n40553 = ~n40582 | ~n41575;
  assign n41768 = ~P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN | ~P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN;
  assign n29304 = ~n41768;
  assign n29305 = P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & n29304;
  assign n41869 = ~n29305 | ~P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN;
  assign n40432 = ~n40553 | ~n41869;
  assign n29307 = n40432 | n29306;
  assign n41493 = ~n29308 | ~n29307;
  assign n29309 = ~n41493 | ~n41785;
  assign n29328 = ~n29633 | ~P2_INSTQUEUE_REG_0__3__SCAN_IN;
  assign n29316 = ~n29320 | ~n42120;
  assign n40992 = ~n41575 ^ P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN;
  assign n29315 = ~n40992 | ~n41785;
  assign n29317 = n29316 & n29315;
  assign n29323 = ~n29320 | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n29321 = ~P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n40823 = ~P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ^ n29321;
  assign n29322 = ~n40823 | ~n41785;
  assign n29324 = ~n29633 | ~P2_INSTQUEUE_REG_0__2__SCAN_IN;
  assign n29325 = ~n29324;
  assign n29327 = ~n29326 | ~n29325;
  assign n29329 = ~n29328;
  assign n29334 = ~n29330 | ~n29329;
  assign n29332 = ~n29331;
  assign n29333 = ~n29332 | ~P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN;
  assign n29337 = P2_INSTQUEUE_REG_0__7__SCAN_IN & P2_INSTQUEUE_REG_0__5__SCAN_IN;
  assign n29336 = P2_INSTQUEUE_REG_0__6__SCAN_IN & P2_INSTQUEUE_REG_0__4__SCAN_IN;
  assign n29338 = ~n29337 | ~n29336;
  assign n29339 = ~n22922 & ~n29338;
  assign n39773 = ~n29340;
  assign n29341 = n39744 & n39762;
  assign n29342 = n39737 & n29341;
  assign n29345 = ~n29436 | ~P2_INSTQUEUE_REG_11__5__SCAN_IN;
  assign n29344 = ~n29475 | ~P2_INSTQUEUE_REG_14__5__SCAN_IN;
  assign n29349 = ~n29345 | ~n29344;
  assign n29347 = ~n29465 | ~P2_INSTQUEUE_REG_8__5__SCAN_IN;
  assign n29346 = ~n29491 | ~P2_INSTQUEUE_REG_7__5__SCAN_IN;
  assign n29348 = ~n29347 | ~n29346;
  assign n29364 = ~n29349 & ~n29348;
  assign n29352 = ~n23277 & ~n40513;
  assign n29425 = ~n29592;
  assign n29351 = ~n29425 & ~n29350;
  assign n29354 = ~n29352 & ~n29351;
  assign n29353 = ~n29588 | ~P2_INSTQUEUE_REG_2__5__SCAN_IN;
  assign n29358 = ~n29354 | ~n29353;
  assign n29450 = ~n29355;
  assign n29357 = ~n29450 & ~n29356;
  assign n29362 = n29358 | n29357;
  assign n29360 = ~n29466 | ~P2_INSTQUEUE_REG_12__5__SCAN_IN;
  assign n29359 = ~n29478 | ~P2_INSTQUEUE_REG_9__5__SCAN_IN;
  assign n29361 = ~n29360 | ~n29359;
  assign n29363 = ~n29362 & ~n29361;
  assign n29377 = ~n29364 | ~n29363;
  assign n29367 = n29580 | n29365;
  assign n29366 = ~n29597 | ~P2_INSTQUEUE_REG_5__5__SCAN_IN;
  assign n29371 = ~n29367 | ~n29366;
  assign n29369 = ~n27509 | ~P2_INSTQUEUE_REG_13__5__SCAN_IN;
  assign n29368 = ~n29591 | ~P2_INSTQUEUE_REG_15__5__SCAN_IN;
  assign n29370 = ~n29369 | ~n29368;
  assign n29375 = ~n29371 & ~n29370;
  assign n29373 = n29602 | n29651;
  assign n29372 = n33147 | n29656;
  assign n29374 = n29373 & n29372;
  assign n29376 = ~n29375 | ~n29374;
  assign n31914 = ~n29377 & ~n29376;
  assign n29379 = ~n29479 | ~P2_INSTQUEUE_REG_6__3__SCAN_IN;
  assign n29378 = ~n28734 | ~P2_INSTQUEUE_REG_0__3__SCAN_IN;
  assign n29383 = ~n29379 | ~n29378;
  assign n29381 = ~n29469 | ~P2_INSTQUEUE_REG_4__3__SCAN_IN;
  assign n29380 = ~n29474 | ~P2_INSTQUEUE_REG_10__3__SCAN_IN;
  assign n29382 = ~n29381 | ~n29380;
  assign n29391 = ~n29383 & ~n29382;
  assign n29385 = ~n29436 | ~P2_INSTQUEUE_REG_11__3__SCAN_IN;
  assign n29384 = ~n27509 | ~P2_INSTQUEUE_REG_13__3__SCAN_IN;
  assign n29389 = ~n29385 | ~n29384;
  assign n29387 = ~n29465 | ~P2_INSTQUEUE_REG_8__3__SCAN_IN;
  assign n29386 = ~n29478 | ~P2_INSTQUEUE_REG_9__3__SCAN_IN;
  assign n29388 = ~n29387 | ~n29386;
  assign n29390 = ~n29389 & ~n29388;
  assign n29409 = ~n29391 | ~n29390;
  assign n29393 = ~n29519 | ~P2_INSTQUEUE_REG_3__3__SCAN_IN;
  assign n29392 = ~n27817 | ~P2_INSTQUEUE_REG_7__3__SCAN_IN;
  assign n29400 = ~n29393 | ~n29392;
  assign n29398 = n29575 | n29394;
  assign n29396 = ~n29592 | ~P2_INSTQUEUE_REG_1__3__SCAN_IN;
  assign n29395 = ~n29588 | ~P2_INSTQUEUE_REG_2__3__SCAN_IN;
  assign n29397 = n29396 & n29395;
  assign n29399 = ~n29398 | ~n29397;
  assign n29407 = ~n29400 & ~n29399;
  assign n29402 = ~n29597 | ~P2_INSTQUEUE_REG_5__3__SCAN_IN;
  assign n29401 = ~n29591 | ~P2_INSTQUEUE_REG_15__3__SCAN_IN;
  assign n29405 = ~n29402 | ~n29401;
  assign n29404 = ~n29581 & ~n29403;
  assign n29406 = ~n29405 & ~n29404;
  assign n29408 = ~n29407 | ~n29406;
  assign n31932 = ~n29409 & ~n29408;
  assign n29615 = ~n31914 & ~n31932;
  assign n29411 = ~n29479 | ~P2_INSTQUEUE_REG_6__1__SCAN_IN;
  assign n29410 = ~n29591 | ~P2_INSTQUEUE_REG_15__1__SCAN_IN;
  assign n29415 = ~n29411 | ~n29410;
  assign n29413 = ~n29519 | ~P2_INSTQUEUE_REG_3__1__SCAN_IN;
  assign n29412 = ~n27509 | ~P2_INSTQUEUE_REG_13__1__SCAN_IN;
  assign n29414 = ~n29413 | ~n29412;
  assign n29423 = ~n29415 & ~n29414;
  assign n29417 = ~n29474 | ~P2_INSTQUEUE_REG_10__1__SCAN_IN;
  assign n29416 = ~n29478 | ~P2_INSTQUEUE_REG_9__1__SCAN_IN;
  assign n29421 = ~n29417 | ~n29416;
  assign n29419 = ~n27817 | ~P2_INSTQUEUE_REG_7__1__SCAN_IN;
  assign n29418 = ~n29475 | ~P2_INSTQUEUE_REG_14__1__SCAN_IN;
  assign n29420 = ~n29419 | ~n29418;
  assign n29422 = ~n29421 & ~n29420;
  assign n29446 = ~n29423 | ~n29422;
  assign n29429 = ~n29425 & ~n29424;
  assign n29427 = ~n29588;
  assign n29428 = ~n29427 & ~n29426;
  assign n29431 = ~n29429 & ~n29428;
  assign n29430 = ~n29466 | ~P2_INSTQUEUE_REG_12__1__SCAN_IN;
  assign n29435 = ~n29431 | ~n29430;
  assign n29433 = ~n29465 | ~P2_INSTQUEUE_REG_8__1__SCAN_IN;
  assign n29432 = ~n29469 | ~P2_INSTQUEUE_REG_4__1__SCAN_IN;
  assign n29434 = ~n29433 | ~n29432;
  assign n29444 = ~n29435 & ~n29434;
  assign n29438 = ~n29436;
  assign n29442 = ~n29438 & ~n29437;
  assign n29440 = ~n29597 | ~P2_INSTQUEUE_REG_5__1__SCAN_IN;
  assign n29439 = ~n28734 | ~P2_INSTQUEUE_REG_0__1__SCAN_IN;
  assign n29441 = ~n29440 | ~n29439;
  assign n29443 = ~n29442 & ~n29441;
  assign n29445 = ~n29444 | ~n29443;
  assign n31951 = ~n29446 & ~n29445;
  assign n29448 = ~n29491;
  assign n29452 = ~n29448 & ~n29447;
  assign n29451 = ~n29450 & ~n29449;
  assign n29464 = ~n29452 & ~n29451;
  assign n29454 = ~n28734 | ~P2_INSTQUEUE_REG_0__4__SCAN_IN;
  assign n29453 = ~n29591 | ~P2_INSTQUEUE_REG_15__4__SCAN_IN;
  assign n29458 = ~n29454 | ~n29453;
  assign n29456 = ~n29592 | ~P2_INSTQUEUE_REG_1__4__SCAN_IN;
  assign n29455 = ~n29588 | ~P2_INSTQUEUE_REG_2__4__SCAN_IN;
  assign n29457 = ~n29456 | ~n29455;
  assign n29462 = n29458 | n29457;
  assign n29460 = ~n27509 | ~P2_INSTQUEUE_REG_13__4__SCAN_IN;
  assign n29459 = ~n29597 | ~P2_INSTQUEUE_REG_5__4__SCAN_IN;
  assign n29461 = ~n29460 | ~n29459;
  assign n29463 = ~n29462 & ~n29461;
  assign n29487 = ~n29464 | ~n29463;
  assign n29468 = ~n29465 | ~P2_INSTQUEUE_REG_8__4__SCAN_IN;
  assign n29467 = ~n29466 | ~P2_INSTQUEUE_REG_12__4__SCAN_IN;
  assign n29473 = ~n29468 | ~n29467;
  assign n29471 = ~n29469 | ~P2_INSTQUEUE_REG_4__4__SCAN_IN;
  assign n29470 = ~n29436 | ~P2_INSTQUEUE_REG_11__4__SCAN_IN;
  assign n29472 = ~n29471 | ~n29470;
  assign n29485 = ~n29473 & ~n29472;
  assign n29477 = ~n29474 | ~P2_INSTQUEUE_REG_10__4__SCAN_IN;
  assign n29476 = ~n29475 | ~P2_INSTQUEUE_REG_14__4__SCAN_IN;
  assign n29483 = ~n29477 | ~n29476;
  assign n29481 = ~n29478 | ~P2_INSTQUEUE_REG_9__4__SCAN_IN;
  assign n29480 = ~n29479 | ~P2_INSTQUEUE_REG_6__4__SCAN_IN;
  assign n29482 = ~n29481 | ~n29480;
  assign n29484 = ~n29483 & ~n29482;
  assign n29486 = ~n29485 | ~n29484;
  assign n31905 = ~n29487 & ~n29486;
  assign n29490 = ~n29436 | ~P2_INSTQUEUE_REG_11__2__SCAN_IN;
  assign n29488 = ~P2_INSTQUEUE_REG_14__2__SCAN_IN;
  assign n29489 = n29581 | n29488;
  assign n29496 = ~n29490 | ~n29489;
  assign n29494 = ~n29491 | ~P2_INSTQUEUE_REG_7__2__SCAN_IN;
  assign n29492 = ~P2_INSTQUEUE_REG_9__2__SCAN_IN;
  assign n29493 = n29569 | n29492;
  assign n29495 = ~n29494 | ~n29493;
  assign n29508 = n29496 | n29495;
  assign n29500 = n29577 | n29497;
  assign n29499 = n29575 | n29498;
  assign n29506 = ~n29500 | ~n29499;
  assign n29504 = n29580 | n29501;
  assign n29503 = n33147 | n29502;
  assign n29505 = ~n29504 | ~n29503;
  assign n29507 = n29506 | n29505;
  assign n29526 = ~n29508 & ~n29507;
  assign n29510 = ~n28734 | ~P2_INSTQUEUE_REG_0__2__SCAN_IN;
  assign n29509 = ~n29592 | ~P2_INSTQUEUE_REG_1__2__SCAN_IN;
  assign n29514 = ~n29510 | ~n29509;
  assign n29512 = ~n29591 | ~P2_INSTQUEUE_REG_15__2__SCAN_IN;
  assign n29511 = ~n29588 | ~P2_INSTQUEUE_REG_2__2__SCAN_IN;
  assign n29513 = ~n29512 | ~n29511;
  assign n29518 = ~n29514 & ~n29513;
  assign n29516 = ~n29597 | ~P2_INSTQUEUE_REG_5__2__SCAN_IN;
  assign n29515 = ~n27509 | ~P2_INSTQUEUE_REG_13__2__SCAN_IN;
  assign n29517 = n29516 & n29515;
  assign n29524 = ~n29518 | ~n29517;
  assign n29522 = ~n29519 | ~P2_INSTQUEUE_REG_3__2__SCAN_IN;
  assign n29521 = n29602 | n29520;
  assign n29523 = ~n29522 | ~n29521;
  assign n29525 = ~n29524 & ~n29523;
  assign n31904 = n29526 & n29525;
  assign n29612 = ~n31905 & ~n31904;
  assign n29529 = ~n29436 | ~P2_INSTQUEUE_REG_11__0__SCAN_IN;
  assign n29528 = n33147 | n29527;
  assign n29535 = ~n29529 | ~n29528;
  assign n29533 = ~n29530 | ~P2_INSTQUEUE_REG_3__0__SCAN_IN;
  assign n29531 = ~P2_INSTQUEUE_REG_9__0__SCAN_IN;
  assign n29532 = n29569 | n29531;
  assign n29534 = ~n29533 | ~n29532;
  assign n29547 = n29535 | n29534;
  assign n29539 = n29577 | n29536;
  assign n29538 = n29575 | n29537;
  assign n29545 = ~n29539 | ~n29538;
  assign n29543 = n29580 | n29540;
  assign n29541 = ~P2_INSTQUEUE_REG_14__0__SCAN_IN;
  assign n29542 = n29581 | n29541;
  assign n29544 = ~n29543 | ~n29542;
  assign n29546 = n29545 | n29544;
  assign n29564 = ~n29547 & ~n29546;
  assign n29549 = ~n28734 | ~P2_INSTQUEUE_REG_0__0__SCAN_IN;
  assign n29548 = ~n29588 | ~P2_INSTQUEUE_REG_2__0__SCAN_IN;
  assign n29553 = ~n29549 | ~n29548;
  assign n29551 = ~n29591 | ~P2_INSTQUEUE_REG_15__0__SCAN_IN;
  assign n29550 = ~n29592 | ~P2_INSTQUEUE_REG_1__0__SCAN_IN;
  assign n29552 = ~n29551 | ~n29550;
  assign n29557 = ~n29553 & ~n29552;
  assign n29555 = ~n27509 | ~P2_INSTQUEUE_REG_13__0__SCAN_IN;
  assign n29554 = ~n27510 | ~P2_INSTQUEUE_REG_5__0__SCAN_IN;
  assign n29556 = n29555 & n29554;
  assign n29562 = ~n29557 | ~n29556;
  assign n29560 = ~n27817 | ~P2_INSTQUEUE_REG_7__0__SCAN_IN;
  assign n29559 = n29602 | n29558;
  assign n29561 = ~n29560 | ~n29559;
  assign n29563 = ~n29562 & ~n29561;
  assign n39698 = ~n29564 | ~n29563;
  assign n29567 = ~n27817 | ~P2_INSTQUEUE_REG_7__6__SCAN_IN;
  assign n29566 = ~n29436 | ~P2_INSTQUEUE_REG_11__6__SCAN_IN;
  assign n29573 = ~n29567 | ~n29566;
  assign n29571 = n33147 | n29687;
  assign n29570 = n29569 | n29568;
  assign n29572 = ~n29571 | ~n29570;
  assign n29587 = n29573 | n29572;
  assign n29579 = n29575 | n29574;
  assign n29578 = n29577 | n29576;
  assign n29585 = ~n29579 | ~n29578;
  assign n29583 = n29580 | n29717;
  assign n29701 = ~P2_INSTQUEUE_REG_14__6__SCAN_IN;
  assign n29582 = n29581 | n29701;
  assign n29584 = ~n29583 | ~n29582;
  assign n29586 = n29585 | n29584;
  assign n29608 = ~n29587 & ~n29586;
  assign n29590 = ~n28734 | ~P2_INSTQUEUE_REG_0__6__SCAN_IN;
  assign n29589 = ~n29588 | ~P2_INSTQUEUE_REG_2__6__SCAN_IN;
  assign n29596 = ~n29590 | ~n29589;
  assign n29594 = ~n29591 | ~P2_INSTQUEUE_REG_15__6__SCAN_IN;
  assign n29593 = ~n29592 | ~P2_INSTQUEUE_REG_1__6__SCAN_IN;
  assign n29595 = ~n29594 | ~n29593;
  assign n29601 = ~n29596 & ~n29595;
  assign n29599 = ~n27509 | ~P2_INSTQUEUE_REG_13__6__SCAN_IN;
  assign n29598 = ~n29597 | ~P2_INSTQUEUE_REG_5__6__SCAN_IN;
  assign n29600 = n29599 & n29598;
  assign n29606 = ~n29601 | ~n29600;
  assign n29604 = ~n29355 | ~P2_INSTQUEUE_REG_3__6__SCAN_IN;
  assign n29603 = n29602 | n29712;
  assign n29605 = ~n29604 | ~n29603;
  assign n29607 = ~n29606 & ~n29605;
  assign n31906 = ~n29608 | ~n29607;
  assign n29610 = ~n39698 | ~n31906;
  assign n39708 = ~n29609;
  assign n29611 = ~n29610 & ~n39708;
  assign n29613 = ~n29612 | ~n29611;
  assign n29614 = ~n31951 & ~n29613;
  assign n29616 = ~n29615 | ~n29614;
  assign n29617 = ~n40456 | ~n29619;
  assign n29620 = ~n29619;
  assign n31897 = ~n40456 & ~n29620;
  assign n29622 = ~n29621 | ~n29625;
  assign n29623 = ~n29622 | ~n29633;
  assign n31889 = ~n29624 & ~n29623;
  assign n31888 = ~n29625 & ~n40456;
  assign n29626 = ~n31889 & ~n31888;
  assign n29629 = ~n29628 ^ n29627;
  assign n31881 = n40456 | n29630;
  assign n29632 = ~n29631;
  assign n29634 = ~n29632 | ~n29637;
  assign n29635 = ~n29634 | ~n29633;
  assign n29638 = ~n29636 & ~n29635;
  assign n31871 = ~n29637 & ~n40456;
  assign n29639 = ~n23515 | ~n29638;
  assign n29640 = ~n29660 | ~P2_INSTQUEUE_REG_5__5__SCAN_IN;
  assign n29642 = ~n29640 | ~n29713;
  assign n29641 = ~n27418 & ~n40513;
  assign n29650 = ~n29642 & ~n29641;
  assign n29644 = ~n29760 | ~P2_INSTQUEUE_REG_2__5__SCAN_IN;
  assign n29643 = ~n23145 | ~P2_INSTQUEUE_REG_7__5__SCAN_IN;
  assign n29648 = ~n29644 | ~n29643;
  assign n29646 = ~n29752 | ~P2_INSTQUEUE_REG_4__5__SCAN_IN;
  assign n29645 = ~n29756 | ~P2_INSTQUEUE_REG_3__5__SCAN_IN;
  assign n29647 = ~n29646 | ~n29645;
  assign n29649 = ~n29648 & ~n29647;
  assign n29655 = ~n29650 | ~n29649;
  assign n29653 = ~n29753 | ~P2_INSTQUEUE_REG_1__5__SCAN_IN;
  assign n29652 = n29731 | n29651;
  assign n29654 = ~n29653 | ~n29652;
  assign n29676 = n29655 | n29654;
  assign n29659 = ~n29688 & ~n29656;
  assign n29657 = ~n29756 | ~P2_INSTQUEUE_REG_11__5__SCAN_IN;
  assign n29658 = ~n29657 | ~n29767;
  assign n29668 = ~n29659 & ~n29658;
  assign n29662 = ~n29660 | ~P2_INSTQUEUE_REG_13__5__SCAN_IN;
  assign n29661 = ~n23145 | ~P2_INSTQUEUE_REG_15__5__SCAN_IN;
  assign n29666 = ~n29662 | ~n29661;
  assign n29664 = ~n29753 | ~P2_INSTQUEUE_REG_9__5__SCAN_IN;
  assign n29663 = ~n29761 | ~P2_INSTQUEUE_REG_14__5__SCAN_IN;
  assign n29665 = ~n29664 | ~n29663;
  assign n29667 = ~n29666 & ~n29665;
  assign n29674 = ~n29668 | ~n29667;
  assign n29672 = n27418 | n29669;
  assign n29671 = n29718 | n29670;
  assign n29673 = ~n29672 | ~n29671;
  assign n29675 = n29674 | n29673;
  assign n29684 = ~n29676 | ~n29675;
  assign n29677 = ~n29684;
  assign n31865 = ~n40456 & ~n29680;
  assign n29678 = ~n29677 | ~n31865;
  assign n31859 = ~n29679 | ~n23048;
  assign n29686 = ~n29681 & ~n29680;
  assign n31860 = n29684 ^ n29686;
  assign n29685 = ~n29684 & ~n42208;
  assign n29728 = ~n29686 | ~n29685;
  assign n29691 = ~n29688 & ~n29687;
  assign n29689 = ~n29753 | ~P2_INSTQUEUE_REG_9__6__SCAN_IN;
  assign n29690 = ~n29689 | ~n29767;
  assign n29700 = ~n29691 & ~n29690;
  assign n29693 = ~n29752 | ~P2_INSTQUEUE_REG_12__6__SCAN_IN;
  assign n29692 = ~n29739 | ~P2_INSTQUEUE_REG_8__6__SCAN_IN;
  assign n29698 = ~n29693 | ~n29692;
  assign n29695 = ~n23145 | ~P2_INSTQUEUE_REG_15__6__SCAN_IN;
  assign n29697 = ~n29696 | ~n29695;
  assign n29699 = ~n29698 & ~n29697;
  assign n29705 = ~n29700 | ~n29699;
  assign n29703 = ~n29757 | ~P2_INSTQUEUE_REG_13__6__SCAN_IN;
  assign n29702 = n29731 | n29701;
  assign n29704 = ~n29703 | ~n29702;
  assign n29726 = n29705 | n29704;
  assign n29707 = ~n29753 | ~P2_INSTQUEUE_REG_1__6__SCAN_IN;
  assign n29706 = ~n29757 | ~P2_INSTQUEUE_REG_5__6__SCAN_IN;
  assign n29711 = ~n29707 | ~n29706;
  assign n29708 = ~n29760 | ~P2_INSTQUEUE_REG_2__6__SCAN_IN;
  assign n29710 = ~n29709 | ~n29708;
  assign n29724 = ~n29711 & ~n29710;
  assign n29714 = n29731 | n29712;
  assign n29716 = n29714 & n29713;
  assign n29715 = ~n23145 | ~P2_INSTQUEUE_REG_7__6__SCAN_IN;
  assign n29722 = ~n29716 | ~n29715;
  assign n29720 = n29718 | n29717;
  assign n29719 = n27418 | n40530;
  assign n29721 = ~n29720 | ~n29719;
  assign n29723 = ~n29722 & ~n29721;
  assign n29725 = ~n29724 | ~n29723;
  assign n29727 = ~n29726 | ~n29725;
  assign n29729 = ~n29728 & ~n29727;
  assign n29732 = ~n29731 & ~n29730;
  assign n29734 = ~n29732 & ~n29767;
  assign n29733 = ~n23145 | ~P2_INSTQUEUE_REG_7__7__SCAN_IN;
  assign n29738 = ~n29734 | ~n29733;
  assign n29736 = ~n29752 | ~P2_INSTQUEUE_REG_4__7__SCAN_IN;
  assign n29735 = ~n29760 | ~P2_INSTQUEUE_REG_2__7__SCAN_IN;
  assign n29737 = ~n29736 | ~n29735;
  assign n29747 = ~n29738 & ~n29737;
  assign n29741 = ~n29739 | ~P2_INSTQUEUE_REG_0__7__SCAN_IN;
  assign n29740 = ~n29756 | ~P2_INSTQUEUE_REG_3__7__SCAN_IN;
  assign n29745 = ~n29741 | ~n29740;
  assign n29743 = ~n29753 | ~P2_INSTQUEUE_REG_1__7__SCAN_IN;
  assign n29742 = ~n29757 | ~P2_INSTQUEUE_REG_5__7__SCAN_IN;
  assign n29744 = ~n29743 | ~n29742;
  assign n29746 = ~n29745 & ~n29744;
  assign n29773 = ~n29747 | ~n29746;
  assign n29748 = ~P2_INSTQUEUE_REG_15__7__SCAN_IN;
  assign n29751 = ~n29103 & ~n29748;
  assign n29750 = ~n27418 & ~n29749;
  assign n29771 = ~n29751 & ~n29750;
  assign n29755 = ~n29752 | ~P2_INSTQUEUE_REG_12__7__SCAN_IN;
  assign n29754 = ~n29753 | ~P2_INSTQUEUE_REG_9__7__SCAN_IN;
  assign n29769 = ~n29755 | ~n29754;
  assign n29759 = ~n29756 | ~P2_INSTQUEUE_REG_11__7__SCAN_IN;
  assign n29758 = ~n29757 | ~P2_INSTQUEUE_REG_13__7__SCAN_IN;
  assign n29765 = ~n29759 | ~n29758;
  assign n29763 = ~n29760 | ~P2_INSTQUEUE_REG_10__7__SCAN_IN;
  assign n29762 = ~n29761 | ~P2_INSTQUEUE_REG_14__7__SCAN_IN;
  assign n29764 = ~n29763 | ~n29762;
  assign n29766 = ~n29765 & ~n29764;
  assign n29768 = ~n29767 | ~n29766;
  assign n29770 = ~n29769 & ~n29768;
  assign n29772 = ~n29771 | ~n29770;
  assign n29796 = ~n31971 | ~n39782;
  assign n29779 = ~n28366 | ~P2_INSTADDRPOINTER_REG_30__SCAN_IN;
  assign n29775 = ~n29843 | ~P2_EBX_REG_30__SCAN_IN;
  assign n29774 = ~P2_PHYADDRPOINTER_REG_30__SCAN_IN | ~P2_STATE2_REG_1__SCAN_IN;
  assign n29777 = ~n29775 | ~n29774;
  assign n42056 = ~P2_REIP_REG_30__SCAN_IN;
  assign n29776 = ~n28476 & ~n42056;
  assign n29778 = ~n29777 & ~n29776;
  assign n29841 = ~n29779 | ~n29778;
  assign n29786 = ~n28366 | ~P2_INSTADDRPOINTER_REG_28__SCAN_IN;
  assign n29782 = ~n29843 | ~P2_EBX_REG_28__SCAN_IN;
  assign n29781 = ~P2_PHYADDRPOINTER_REG_28__SCAN_IN | ~P2_STATE2_REG_1__SCAN_IN;
  assign n29784 = ~n29782 | ~n29781;
  assign n42045 = ~P2_REIP_REG_28__SCAN_IN;
  assign n29783 = ~n28476 & ~n42045;
  assign n29785 = ~n29784 & ~n29783;
  assign n31723 = ~n29786 | ~n29785;
  assign n29792 = ~n28366 | ~P2_INSTADDRPOINTER_REG_29__SCAN_IN;
  assign n29788 = ~n29843 | ~P2_EBX_REG_29__SCAN_IN;
  assign n29787 = ~P2_PHYADDRPOINTER_REG_29__SCAN_IN | ~P2_STATE2_REG_1__SCAN_IN;
  assign n29790 = ~n29788 | ~n29787;
  assign n42050 = ~P2_REIP_REG_29__SCAN_IN;
  assign n29789 = ~n28476 & ~n42050;
  assign n29791 = ~n29790 & ~n29789;
  assign n31680 = ~n32615;
  assign n29794 = ~n31680 | ~n31948;
  assign n31682 = ~P2_EBX_REG_30__SCAN_IN;
  assign n29793 = ~n39817 | ~n31682;
  assign n29795 = ~n29794 | ~n29793;
  assign P2_U2857 = ~n29796 | ~n29795;
  assign n32617 = ~P2_INSTADDRPOINTER_REG_30__SCAN_IN;
  assign n29863 = ~n29798 ^ n29797;
  assign n29862 = ~n29863 | ~n40348;
  assign n29802 = n28552 & P2_EBX_REG_28__SCAN_IN;
  assign n29804 = ~n29803 | ~n29802;
  assign n32227 = ~n29811 ^ P2_INSTADDRPOINTER_REG_28__SCAN_IN;
  assign n29806 = ~n29805 | ~n32222;
  assign n29807 = ~n29806 | ~n32277;
  assign n29809 = ~n29808 & ~n29807;
  assign n29816 = ~n29811 & ~n32222;
  assign n29812 = ~n29831 | ~P2_INSTADDRPOINTER_REG_28__SCAN_IN;
  assign n29814 = n31728 | n29812;
  assign n29815 = ~n29814 | ~n29813;
  assign n29817 = ~n29816 & ~n29815;
  assign n29818 = ~n28552 | ~P2_EBX_REG_29__SCAN_IN;
  assign n29819 = ~n29818;
  assign n29821 = ~n29820 | ~n29819;
  assign n31705 = ~n29823 | ~n29821;
  assign n32638 = ~P2_INSTADDRPOINTER_REG_29__SCAN_IN;
  assign n32198 = ~n29829 | ~n32638;
  assign n29822 = n28552 & P2_EBX_REG_30__SCAN_IN;
  assign n31681 = ~n29823 ^ n29822;
  assign n32184 = n31681 | n28071;
  assign n29826 = ~n29825 | ~n29824;
  assign n31596 = ~n29827 | ~n29826;
  assign n29828 = ~n31596 | ~n29831;
  assign n29830 = ~n29829;
  assign n32199 = ~n29830 | ~P2_INSTADDRPOINTER_REG_29__SCAN_IN;
  assign n29832 = ~n29831 | ~P2_INSTADDRPOINTER_REG_30__SCAN_IN;
  assign n29834 = ~n32199 | ~n29832;
  assign n29833 = ~n31681;
  assign n29835 = ~n29834 | ~n29833;
  assign n29837 = ~n29835;
  assign n29838 = ~n29837 & ~n23575;
  assign n29840 = ~n29839 | ~n29838;
  assign n29851 = ~n29842 | ~n29841;
  assign n29849 = ~n28366 | ~P2_INSTADDRPOINTER_REG_31__SCAN_IN;
  assign n29845 = ~n29843 | ~P2_EBX_REG_31__SCAN_IN;
  assign n29844 = ~P2_PHYADDRPOINTER_REG_31__SCAN_IN | ~P2_STATE2_REG_1__SCAN_IN;
  assign n29847 = ~n29845 | ~n29844;
  assign n42055 = ~P2_REIP_REG_31__SCAN_IN;
  assign n29846 = ~n28476 & ~n42055;
  assign n29848 = ~n29847 & ~n29846;
  assign n29850 = ~n29849 | ~n29848;
  assign n42137 = ~n42123 | ~n42196;
  assign n42176 = ~n41002 | ~n42137;
  assign n29852 = ~n42176 | ~n42214;
  assign n29860 = ~n29864 | ~n40324;
  assign n31626 = ~P2_PHYADDRPOINTER_REG_29__SCAN_IN;
  assign n31628 = ~P2_PHYADDRPOINTER_REG_27__SCAN_IN;
  assign n31630 = ~P2_PHYADDRPOINTER_REG_25__SCAN_IN;
  assign n31636 = ~P2_PHYADDRPOINTER_REG_19__SCAN_IN;
  assign n31640 = ~P2_PHYADDRPOINTER_REG_15__SCAN_IN;
  assign n31644 = ~P2_PHYADDRPOINTER_REG_11__SCAN_IN;
  assign n31650 = ~P2_PHYADDRPOINTER_REG_5__SCAN_IN;
  assign n31652 = ~P2_PHYADDRPOINTER_REG_3__SCAN_IN;
  assign n31649 = ~P2_PHYADDRPOINTER_REG_4__SCAN_IN | ~n31657;
  assign n31647 = ~P2_PHYADDRPOINTER_REG_6__SCAN_IN | ~n31658;
  assign n31645 = ~P2_PHYADDRPOINTER_REG_8__SCAN_IN | ~n31659;
  assign n31643 = ~P2_PHYADDRPOINTER_REG_10__SCAN_IN | ~n31660;
  assign n31641 = ~P2_PHYADDRPOINTER_REG_12__SCAN_IN | ~n31661;
  assign n31637 = ~P2_PHYADDRPOINTER_REG_16__SCAN_IN | ~n31663;
  assign n31633 = ~P2_PHYADDRPOINTER_REG_20__SCAN_IN | ~n31665;
  assign n31629 = ~P2_PHYADDRPOINTER_REG_24__SCAN_IN | ~n31667;
  assign n31625 = ~P2_PHYADDRPOINTER_REG_28__SCAN_IN | ~n31669;
  assign n31622 = ~P2_PHYADDRPOINTER_REG_31__SCAN_IN ^ n29854;
  assign n31601 = ~n41789 | ~P2_STATE2_REG_1__SCAN_IN;
  assign n40338 = n29855 & n31601;
  assign n40304 = n40337 | n40338;
  assign n40330 = ~n40304;
  assign n29858 = n31622 & n40330;
  assign n29878 = ~n40325 | ~P2_REIP_REG_31__SCAN_IN;
  assign n29856 = ~n40337 | ~P2_PHYADDRPOINTER_REG_31__SCAN_IN;
  assign n29857 = ~n29878 | ~n29856;
  assign n29859 = ~n29858 & ~n29857;
  assign P2_U2983 = ~n29862 | ~n29861;
  assign n29909 = ~n29863 | ~n40356;
  assign n29881 = ~n31595 & ~n33125;
  assign n29865 = ~n32222 & ~n32638;
  assign n29871 = ~P2_INSTADDRPOINTER_REG_28__SCAN_IN | ~n29865;
  assign n29868 = ~n32996 | ~n29866;
  assign n32713 = ~n29868 | ~n29867;
  assign n32655 = ~n32713 | ~n29869;
  assign n32618 = ~n29871 & ~n32655;
  assign n29870 = ~n32618 | ~P2_INSTADDRPOINTER_REG_30__SCAN_IN;
  assign n29877 = ~n29870 | ~n29797;
  assign n33124 = ~n40390 | ~n32993;
  assign n29874 = ~n33124 | ~n32617;
  assign n29872 = n33124 & n29871;
  assign n32616 = ~n29873 & ~n29872;
  assign n29875 = ~n29874 | ~n32616;
  assign n29876 = n29875 | n29797;
  assign n29879 = ~n29877 | ~n29876;
  assign n29880 = ~n29879 | ~n29878;
  assign n31725 = ~n31763 & ~n29882;
  assign n29886 = ~n28980 | ~P2_REIP_REG_28__SCAN_IN;
  assign n29884 = ~n29891 & ~n32653;
  assign n40182 = ~P2_EAX_REG_28__SCAN_IN;
  assign n29883 = ~n28596 & ~n40182;
  assign n29885 = ~n29884 & ~n29883;
  assign n31724 = ~n29886 | ~n29885;
  assign n31701 = ~n31725 | ~n31724;
  assign n29890 = ~n29896 & ~n42050;
  assign n29888 = ~n29897 | ~P2_INSTADDRPOINTER_REG_29__SCAN_IN;
  assign n29887 = ~n29898 | ~P2_EAX_REG_29__SCAN_IN;
  assign n29889 = ~n29888 | ~n29887;
  assign n31702 = ~n29890 & ~n29889;
  assign n29895 = n29896 | n42056;
  assign n29893 = n29891 | n32617;
  assign n40194 = ~P2_EAX_REG_30__SCAN_IN;
  assign n29892 = n28596 | n40194;
  assign n29894 = n29893 & n29892;
  assign n31696 = ~n29895 | ~n29894;
  assign n29903 = ~n31700 | ~n31696;
  assign n29902 = ~n29896 & ~n42055;
  assign n29900 = ~n29897 | ~P2_INSTADDRPOINTER_REG_31__SCAN_IN;
  assign n29899 = ~n29898 | ~P2_EAX_REG_31__SCAN_IN;
  assign n29901 = ~n29900 | ~n29899;
  assign n29904 = ~n39820 | ~n33115;
  assign n29906 = ~n29905 | ~n29904;
  assign n29908 = ~n29907 & ~n29906;
  assign P2_U3015 = ~n29909 | ~n29908;
  assign n29930 = ~n30441 | ~n42343;
  assign n29912 = ~n29952 | ~n29911;
  assign n29915 = ~n29913 | ~n29912;
  assign n29922 = ~n23799 | ~n42488;
  assign n30036 = ~n42481;
  assign n30349 = ~P1_EBX_REG_30__SCAN_IN;
  assign n29920 = ~n30036 & ~n30349;
  assign n29918 = ~n42470 | ~P1_PHYADDRPOINTER_REG_30__SCAN_IN;
  assign n29916 = ~n30639 & ~n31580;
  assign n29917 = ~n42413 | ~n30647;
  assign n29919 = ~n29918 | ~n29917;
  assign n29921 = ~n29920 & ~n29919;
  assign n29928 = ~n29922 | ~n29921;
  assign n29923 = n29943 & P1_REIP_REG_29__SCAN_IN;
  assign n29926 = ~n29923 & ~P1_REIP_REG_30__SCAN_IN;
  assign n29925 = ~n29924;
  assign n29927 = ~n29926 & ~n29925;
  assign n29929 = ~n29928 & ~n29927;
  assign P1_U2810 = ~n29930 | ~n29929;
  assign n29935 = ~n29931;
  assign n29934 = ~n29932 & ~n29933;
  assign n29948 = ~n30657 | ~n42343;
  assign n29940 = ~P1_EBX_REG_29__SCAN_IN | ~n42481;
  assign n29938 = P1_PHYADDRPOINTER_REG_29__SCAN_IN & n42470;
  assign n29937 = ~n30658 & ~n42493;
  assign n29939 = ~n29938 & ~n29937;
  assign n29941 = ~n29940 | ~n29939;
  assign n29942 = ~n29959 & ~n44686;
  assign n29944 = ~n29943;
  assign n29945 = ~n29944 & ~P1_REIP_REG_29__SCAN_IN;
  assign n29947 = ~n29946 & ~n29945;
  assign P1_U2811 = ~n29948 | ~n29947;
  assign n29966 = ~n30665 & ~n42373;
  assign n29951 = n29975 & n29950;
  assign n31047 = ~n29952 & ~n29951;
  assign n29958 = ~n31047 | ~n42488;
  assign n29954 = ~n42481 | ~P1_EBX_REG_28__SCAN_IN;
  assign n29953 = ~n42413 | ~n30668;
  assign n29956 = ~n29954 | ~n29953;
  assign n29955 = ~n30666 & ~n42494;
  assign n29957 = ~n29956 & ~n29955;
  assign n29964 = n29958 & n29957;
  assign n29962 = ~n29959 & ~n44681;
  assign n29961 = ~P1_REIP_REG_28__SCAN_IN & ~n29960;
  assign n29963 = ~n29962 & ~n29961;
  assign n29965 = ~n29964 | ~n29963;
  assign P1_U2812 = n29966 | n29965;
  assign n29971 = ~n29967;
  assign n29970 = ~n29969 & ~n29968;
  assign n29990 = ~n30687 | ~n42343;
  assign n29974 = ~n29973 | ~n29972;
  assign n31061 = ~n29975 | ~n29974;
  assign n29979 = ~n31061 & ~n42440;
  assign n29996 = P1_REIP_REG_26__SCAN_IN & n29976;
  assign n29977 = ~n42500 | ~P1_REIP_REG_27__SCAN_IN;
  assign n29978 = ~n29996 & ~n29977;
  assign n29982 = ~n29979 & ~n29978;
  assign n29980 = ~n44671 & ~P1_REIP_REG_27__SCAN_IN;
  assign n29981 = ~n29980 | ~n30005;
  assign n29988 = n29982 & n29981;
  assign n29984 = ~n42481 | ~P1_EBX_REG_27__SCAN_IN;
  assign n29983 = ~n42470 | ~P1_PHYADDRPOINTER_REG_27__SCAN_IN;
  assign n29986 = ~n29984 | ~n29983;
  assign n29985 = ~n30688 & ~n22835;
  assign n29987 = ~n29986 & ~n29985;
  assign n29989 = n29988 & n29987;
  assign P1_U2813 = ~n29990 | ~n29989;
  assign n30698 = ~n29991 ^ n29992;
  assign n30009 = ~n30698 & ~n42373;
  assign n31082 = n29994 ^ n29993;
  assign n30004 = ~n31082 | ~n42488;
  assign n29995 = ~n42500 | ~P1_REIP_REG_26__SCAN_IN;
  assign n30002 = ~n29996 & ~n29995;
  assign n30000 = ~n42481 | ~P1_EBX_REG_26__SCAN_IN;
  assign n29998 = ~n42413 | ~n30700;
  assign n29997 = ~P1_PHYADDRPOINTER_REG_26__SCAN_IN | ~n42470;
  assign n29999 = n29998 & n29997;
  assign n30001 = ~n30000 | ~n29999;
  assign n30003 = ~n30002 & ~n30001;
  assign n30007 = n30004 & n30003;
  assign n30006 = ~n30005 | ~n44671;
  assign n30008 = ~n30007 | ~n30006;
  assign P1_U2814 = n30009 | n30008;
  assign n30012 = ~n30010 | ~n30011;
  assign n30713 = ~n29991 | ~n30012;
  assign n30495 = ~n30713;
  assign n30030 = ~n30495 | ~n42343;
  assign n31092 = ~n30013 ^ n30014;
  assign n30028 = ~n31092 & ~n42440;
  assign n30048 = ~n30327 & ~P1_REIP_REG_24__SCAN_IN;
  assign n44666 = ~P1_REIP_REG_25__SCAN_IN;
  assign n30016 = ~n30048 & ~n44666;
  assign n30047 = ~n30015;
  assign n30041 = ~n42469 | ~n30047;
  assign n30062 = ~n42500 | ~n30041;
  assign n30020 = ~n30016 | ~n30062;
  assign n30018 = ~n42411 | ~n30017;
  assign n30019 = ~n30018 | ~n44666;
  assign n30026 = ~n30020 | ~n30019;
  assign n30371 = ~P1_EBX_REG_25__SCAN_IN;
  assign n30024 = ~n30036 & ~n30371;
  assign n30022 = ~n42413 | ~n30716;
  assign n30021 = ~n42470 | ~P1_PHYADDRPOINTER_REG_25__SCAN_IN;
  assign n30023 = ~n30022 | ~n30021;
  assign n30025 = ~n30024 & ~n30023;
  assign n30027 = ~n30026 | ~n30025;
  assign n30029 = ~n30028 & ~n30027;
  assign P1_U2815 = ~n30030 | ~n30029;
  assign n30031 = ~n30131;
  assign n30117 = ~n30115 & ~n30114;
  assign n30052 = ~n30729 | ~n42343;
  assign n30035 = ~n30013;
  assign n30034 = ~n30058 | ~n30033;
  assign n31109 = ~n30035 | ~n30034;
  assign n30046 = ~n31109 & ~n42440;
  assign n30376 = ~P1_EBX_REG_24__SCAN_IN;
  assign n30040 = ~n30036 & ~n30376;
  assign n30038 = ~n42413 | ~n30734;
  assign n30037 = ~n42470 | ~P1_PHYADDRPOINTER_REG_24__SCAN_IN;
  assign n30039 = ~n30038 | ~n30037;
  assign n30044 = ~n30040 & ~n30039;
  assign n30042 = n30041 & P1_REIP_REG_24__SCAN_IN;
  assign n30043 = ~n42500 | ~n30042;
  assign n30045 = ~n30044 | ~n30043;
  assign n30050 = ~n30046 & ~n30045;
  assign n30049 = ~n30048 | ~n30047;
  assign n30051 = n30050 & n30049;
  assign P1_U2816 = ~n30052 | ~n30051;
  assign n30073 = ~n30741 | ~n42343;
  assign n30057 = ~n30056 | ~n30055;
  assign n31118 = ~n30058 | ~n30057;
  assign n30071 = ~n31118 & ~n42440;
  assign n30746 = ~n30059;
  assign n30069 = ~n30746 | ~n42413;
  assign n30061 = n30060 & n42411;
  assign n30063 = ~n30061 & ~P1_REIP_REG_23__SCAN_IN;
  assign n30067 = ~n30063 & ~n30062;
  assign n30065 = ~n42481 | ~P1_EBX_REG_23__SCAN_IN;
  assign n30064 = ~n42470 | ~P1_PHYADDRPOINTER_REG_23__SCAN_IN;
  assign n30066 = ~n30065 | ~n30064;
  assign n30068 = ~n30067 & ~n30066;
  assign n30070 = ~n30069 | ~n30068;
  assign n30072 = ~n30071 & ~n30070;
  assign P1_U2817 = ~n30073 | ~n30072;
  assign n30096 = ~n30753 | ~n42343;
  assign n44651 = ~P1_REIP_REG_22__SCAN_IN;
  assign n30101 = ~P1_REIP_REG_20__SCAN_IN | ~n30075;
  assign n30076 = ~n30101 & ~n30263;
  assign n30119 = ~n30076 & ~n30287;
  assign n44646 = ~P1_REIP_REG_21__SCAN_IN;
  assign n30100 = ~n42411 | ~n44646;
  assign n30077 = ~n30100;
  assign n30078 = ~n30119 & ~n30077;
  assign n30094 = ~n44651 & ~n30078;
  assign n30185 = ~n42411 | ~n30141;
  assign n30137 = ~n30079 & ~n30185;
  assign n30118 = ~P1_REIP_REG_19__SCAN_IN | ~n30137;
  assign n30082 = ~n30118;
  assign n30081 = ~P1_REIP_REG_22__SCAN_IN & ~n30080;
  assign n30092 = ~n30082 | ~n30081;
  assign n30084 = ~n30083;
  assign n31138 = ~n27102 ^ n30084;
  assign n30086 = ~n31138 | ~n42488;
  assign n30085 = ~n42470 | ~P1_PHYADDRPOINTER_REG_22__SCAN_IN;
  assign n30090 = ~n30086 | ~n30085;
  assign n30088 = ~n42481 | ~P1_EBX_REG_22__SCAN_IN;
  assign n30087 = ~n42413 | ~n30758;
  assign n30089 = ~n30088 | ~n30087;
  assign n30091 = ~n30090 & ~n30089;
  assign n30093 = ~n30092 | ~n30091;
  assign n30095 = ~n30094 & ~n30093;
  assign P1_U2818 = ~n30096 | ~n30095;
  assign n30098 = n30117 | n30097;
  assign n30765 = ~n30099 | ~n30098;
  assign n30113 = ~n30536 | ~n42343;
  assign n30111 = ~n30390 & ~n42440;
  assign n30107 = ~n30119 | ~P1_REIP_REG_21__SCAN_IN;
  assign n30105 = ~n30101 & ~n30100;
  assign n30103 = ~n42481 | ~P1_EBX_REG_21__SCAN_IN;
  assign n30102 = ~n42470 | ~P1_PHYADDRPOINTER_REG_21__SCAN_IN;
  assign n30104 = ~n30103 | ~n30102;
  assign n30106 = ~n30105 & ~n30104;
  assign n30109 = n30107 & n30106;
  assign n30108 = ~n30770 | ~n42413;
  assign n30110 = ~n30109 | ~n30108;
  assign n30112 = ~n30111 & ~n30110;
  assign P1_U2819 = ~n30113 | ~n30112;
  assign n30116 = n30115 & n30114;
  assign n30778 = n30117 | n30116;
  assign n30130 = ~n30778 & ~n42373;
  assign n44641 = ~P1_REIP_REG_20__SCAN_IN;
  assign n30120 = ~n30118 | ~n44641;
  assign n30128 = ~n30120 | ~n30119;
  assign n30122 = ~n42481 | ~P1_EBX_REG_20__SCAN_IN;
  assign n30121 = ~n42413 | ~n30781;
  assign n30126 = ~n30122 | ~n30121;
  assign n30124 = ~n30396 & ~n42440;
  assign n30123 = P1_PHYADDRPOINTER_REG_20__SCAN_IN & n42470;
  assign n30125 = n30124 | n30123;
  assign n30127 = ~n30126 & ~n30125;
  assign n30129 = ~n30128 | ~n30127;
  assign P1_U2820 = n30130 | n30129;
  assign n30151 = ~n30789 | ~n42343;
  assign n30136 = ~n30795 & ~n22835;
  assign n30134 = ~P1_EBX_REG_19__SCAN_IN | ~n42481;
  assign n42367 = ~n42469 | ~n42234;
  assign n30132 = ~n42494 & ~n30792;
  assign n30133 = ~n42389 & ~n30132;
  assign n30135 = ~n30134 | ~n30133;
  assign n30149 = ~n30136 & ~n30135;
  assign n44636 = ~P1_REIP_REG_19__SCAN_IN;
  assign n30147 = ~n44636 | ~n30137;
  assign n30139 = ~n23213 | ~n30138;
  assign n31148 = ~n30140 | ~n30139;
  assign n30145 = ~n31148 & ~n42440;
  assign n30158 = ~P1_REIP_REG_17__SCAN_IN | ~n30141;
  assign n30142 = ~n30263 & ~n30158;
  assign n30184 = ~n30287 & ~n30142;
  assign n30157 = ~n30327 & ~P1_REIP_REG_18__SCAN_IN;
  assign n30143 = ~n30184 & ~n30157;
  assign n30144 = ~n30143 & ~n44636;
  assign n30146 = ~n30145 & ~n30144;
  assign n30148 = n30147 & n30146;
  assign n30150 = n30149 & n30148;
  assign P1_U2821 = ~n30151 | ~n30150;
  assign n30803 = ~n30152 ^ n30153;
  assign n30170 = ~n30803 | ~n42343;
  assign n30155 = ~n42481 | ~P1_EBX_REG_18__SCAN_IN;
  assign n30154 = ~n42413 | ~n30807;
  assign n30168 = ~n30155 | ~n30154;
  assign n31177 = ~n30180 ^ n30156;
  assign n30166 = ~n31177 & ~n42440;
  assign n30159 = ~n30157;
  assign n30162 = ~n30159 & ~n30158;
  assign n30160 = ~n42470 | ~P1_PHYADDRPOINTER_REG_18__SCAN_IN;
  assign n30161 = ~n42367 | ~n30160;
  assign n30164 = ~n30162 & ~n30161;
  assign n30163 = ~n30184 | ~P1_REIP_REG_18__SCAN_IN;
  assign n30165 = ~n30164 | ~n30163;
  assign n30167 = n30166 | n30165;
  assign n30169 = ~n30168 & ~n30167;
  assign P1_U2822 = ~n30170 | ~n30169;
  assign n30173 = ~n30171 & ~n30172;
  assign n30814 = n30152 | n30173;
  assign n30194 = ~n30814 & ~n42373;
  assign n30175 = ~n30174 & ~n42494;
  assign n30177 = ~n30175 & ~n42389;
  assign n30176 = ~n42481 | ~P1_EBX_REG_17__SCAN_IN;
  assign n30179 = ~n30177 | ~n30176;
  assign n30178 = ~n30815 & ~n42493;
  assign n30192 = ~n30179 & ~n30178;
  assign n30183 = ~n30182 | ~n30181;
  assign n31194 = ~n23218 | ~n30183;
  assign n30190 = ~n31194 & ~n42440;
  assign n30188 = ~n30184;
  assign n30186 = ~n30185;
  assign n30187 = ~n30186 & ~P1_REIP_REG_17__SCAN_IN;
  assign n30189 = ~n30188 & ~n30187;
  assign n30191 = ~n30190 & ~n30189;
  assign n30193 = ~n30192 | ~n30191;
  assign P1_U2823 = n30194 | n30193;
  assign n30837 = ~n30195 ^ n30196;
  assign n30589 = ~n30837;
  assign n30214 = ~n30589 | ~n42343;
  assign n30198 = ~n42481 | ~P1_EBX_REG_16__SCAN_IN;
  assign n30197 = ~n42413 | ~n30839;
  assign n30212 = ~n30198 | ~n30197;
  assign n31204 = n30199 ^ n30228;
  assign n30210 = ~n31204 | ~n42488;
  assign n44616 = ~P1_REIP_REG_15__SCAN_IN;
  assign n30219 = ~n42411 | ~n44616;
  assign n30201 = ~n30219 | ~P1_REIP_REG_16__SCAN_IN;
  assign n30200 = ~n42469 | ~n30218;
  assign n30247 = n42500 & n30200;
  assign n30205 = ~n30201 & ~n30247;
  assign n30203 = ~n30327 & ~n30202;
  assign n30204 = ~n30203 & ~P1_REIP_REG_16__SCAN_IN;
  assign n30208 = ~n30205 & ~n30204;
  assign n30206 = ~P1_PHYADDRPOINTER_REG_16__SCAN_IN | ~n42470;
  assign n30207 = ~n42367 | ~n30206;
  assign n30209 = ~n30208 & ~n30207;
  assign n30211 = ~n30210 | ~n30209;
  assign n30213 = ~n30212 & ~n30211;
  assign P1_U2824 = ~n30214 | ~n30213;
  assign n30217 = ~n30215 | ~n30216;
  assign n30854 = ~n30195 | ~n30217;
  assign n30601 = ~n30854;
  assign n30236 = ~n30601 | ~n42343;
  assign n30225 = ~n30855 & ~n42494;
  assign n30220 = ~n30218;
  assign n30222 = ~n30220 & ~n30219;
  assign n30221 = ~n30858 & ~n22835;
  assign n30223 = ~n30222 & ~n30221;
  assign n30224 = ~n42367 | ~n30223;
  assign n30234 = ~n30225 & ~n30224;
  assign n30227 = n23063 | n30226;
  assign n31222 = ~n30228 | ~n30227;
  assign n30232 = ~n31222 & ~n42440;
  assign n30230 = ~n30247 | ~P1_REIP_REG_15__SCAN_IN;
  assign n30229 = ~n42481 | ~P1_EBX_REG_15__SCAN_IN;
  assign n30231 = ~n30230 | ~n30229;
  assign n30233 = ~n30232 & ~n30231;
  assign n30235 = n30234 & n30233;
  assign P1_U2825 = ~n30236 | ~n30235;
  assign n30239 = ~n30237 | ~n30238;
  assign n30869 = ~n30215 | ~n30239;
  assign n30256 = ~n30869 & ~n42373;
  assign n30242 = ~n30871 & ~n22835;
  assign n30240 = ~P1_PHYADDRPOINTER_REG_14__SCAN_IN | ~n42470;
  assign n30241 = ~n42367 | ~n30240;
  assign n30254 = ~n30242 & ~n30241;
  assign n31236 = n30243 ^ n30269;
  assign n30244 = ~n31236;
  assign n30252 = ~n30244 & ~n42440;
  assign n30246 = ~n30245 & ~n30327;
  assign n30248 = n30246 | P1_REIP_REG_14__SCAN_IN;
  assign n30250 = ~n30248 | ~n30247;
  assign n30249 = ~n42481 | ~P1_EBX_REG_14__SCAN_IN;
  assign n30251 = ~n30250 | ~n30249;
  assign n30253 = ~n30252 & ~n30251;
  assign n30255 = ~n30254 | ~n30253;
  assign P1_U2826 = n30256 | n30255;
  assign n30260 = ~n30305 & ~n30304;
  assign n30259 = ~n30257 & ~n30258;
  assign n30284 = ~n30260 & ~n30259;
  assign n30616 = ~n30889;
  assign n30282 = ~n30616 | ~n42343;
  assign n30262 = ~P1_REIP_REG_13__SCAN_IN & ~n30265;
  assign n30313 = ~n30327 & ~n30264;
  assign n30280 = n30262 & n30313;
  assign n30306 = n30264 | n30263;
  assign n30288 = ~n30265 & ~n30306;
  assign n30266 = ~n42500 | ~P1_REIP_REG_13__SCAN_IN;
  assign n30278 = n30288 | n30266;
  assign n30268 = ~n23052 | ~n30267;
  assign n31265 = ~n30269 | ~n30268;
  assign n30276 = ~n31265 & ~n42440;
  assign n30274 = ~n30893 | ~n42413;
  assign n30272 = ~n42481 | ~P1_EBX_REG_13__SCAN_IN;
  assign n30270 = ~n42470 | ~P1_PHYADDRPOINTER_REG_13__SCAN_IN;
  assign n30271 = n30270 & n42367;
  assign n30273 = n30272 & n30271;
  assign n30275 = ~n30274 | ~n30273;
  assign n30277 = ~n30276 & ~n30275;
  assign n30279 = ~n30278 | ~n30277;
  assign n30281 = ~n30280 & ~n30279;
  assign P1_U2827 = ~n30282 | ~n30281;
  assign n30285 = n30284 & n30283;
  assign n30303 = ~n22909 | ~n42343;
  assign n30286 = ~P1_REIP_REG_11__SCAN_IN | ~n30313;
  assign n44602 = ~P1_REIP_REG_12__SCAN_IN;
  assign n30290 = n30286 & n44602;
  assign n30289 = n30288 | n30287;
  assign n30301 = ~n30290 & ~n30289;
  assign n31290 = ~n30292 ^ n30291;
  assign n30299 = ~n31290 & ~n42440;
  assign n30297 = n30911 | n22835;
  assign n30295 = ~n42481 | ~P1_EBX_REG_12__SCAN_IN;
  assign n30293 = ~n42470 | ~P1_PHYADDRPOINTER_REG_12__SCAN_IN;
  assign n30294 = n30293 & n42367;
  assign n30296 = n30295 & n30294;
  assign n30298 = ~n30297 | ~n30296;
  assign n30300 = n30299 | n30298;
  assign n30302 = ~n30301 & ~n30300;
  assign P1_U2828 = ~n30303 | ~n30302;
  assign n30919 = ~n30305 ^ n30304;
  assign n30322 = ~n30919 & ~n42373;
  assign n30326 = ~n42500 | ~n30306;
  assign n44596 = ~P1_REIP_REG_11__SCAN_IN;
  assign n30312 = ~n30326 & ~n44596;
  assign n30308 = ~n30307 & ~n42494;
  assign n30310 = ~n30308 & ~n42389;
  assign n30309 = ~n42413 | ~n30921;
  assign n30311 = ~n30310 | ~n30309;
  assign n30320 = ~n30312 & ~n30311;
  assign n30318 = ~n30313 | ~n44596;
  assign n31303 = n30314 ^ n30332;
  assign n30316 = ~n31303 | ~n42488;
  assign n30315 = ~n42481 | ~P1_EBX_REG_11__SCAN_IN;
  assign n30317 = n30316 & n30315;
  assign n30319 = n30318 & n30317;
  assign n30321 = ~n30320 | ~n30319;
  assign P1_U2829 = n30322 | n30321;
  assign n30325 = ~n30257;
  assign n30324 = ~n30958 & ~n30323;
  assign n42506 = ~n30325 & ~n30324;
  assign n30345 = ~n42506 | ~n42343;
  assign n44591 = ~P1_REIP_REG_10__SCAN_IN;
  assign n30343 = ~n30326 & ~n44591;
  assign n30329 = ~P1_REIP_REG_10__SCAN_IN & ~n30327;
  assign n30341 = ~n30329 | ~n30328;
  assign n30331 = ~n23954 & ~n30330;
  assign n42507 = n30332 | n30331;
  assign n30339 = ~n42507 & ~n42440;
  assign n30337 = ~n42481 | ~P1_EBX_REG_10__SCAN_IN;
  assign n30335 = ~n42493 & ~n30937;
  assign n30333 = ~n42470 | ~P1_PHYADDRPOINTER_REG_10__SCAN_IN;
  assign n30334 = ~n42367 | ~n30333;
  assign n30336 = ~n30335 & ~n30334;
  assign n30338 = ~n30337 | ~n30336;
  assign n30340 = ~n30339 & ~n30338;
  assign n30342 = ~n30341 | ~n30340;
  assign n30344 = ~n30343 & ~n30342;
  assign P1_U2830 = ~n30345 | ~n30344;
  assign n30347 = ~n30346 & ~n42461;
  assign n30353 = ~n30441 | ~n42540;
  assign n30351 = ~n31033 & ~n42553;
  assign n30350 = ~n42561 & ~n30349;
  assign n30352 = ~n30351 & ~n30350;
  assign P1_U2842 = ~n30353 | ~n30352;
  assign n30357 = ~n30657 | ~n42540;
  assign n30355 = ~n31037 & ~n42553;
  assign n30354 = n42556 & P1_EBX_REG_29__SCAN_IN;
  assign n30356 = ~n30355 & ~n30354;
  assign P1_U2843 = ~n30357 | ~n30356;
  assign n30361 = ~n30665 & ~n42562;
  assign n30359 = ~n31047 | ~n42559;
  assign n30358 = ~n42556 | ~P1_EBX_REG_28__SCAN_IN;
  assign n30360 = ~n30359 | ~n30358;
  assign P1_U2844 = n30361 | n30360;
  assign n30362 = ~n30687;
  assign n30366 = ~n30362 & ~n42562;
  assign n30364 = n31061 | n42553;
  assign n30363 = ~n42556 | ~P1_EBX_REG_27__SCAN_IN;
  assign n30365 = ~n30364 | ~n30363;
  assign P1_U2845 = n30366 | n30365;
  assign n30370 = ~n30698 & ~n42562;
  assign n30368 = ~n31082 | ~n42559;
  assign n30367 = ~n42556 | ~P1_EBX_REG_26__SCAN_IN;
  assign n30369 = ~n30368 | ~n30367;
  assign P1_U2846 = n30370 | n30369;
  assign n30375 = ~n30495 | ~n42540;
  assign n30373 = ~n31092 & ~n42553;
  assign n30372 = ~n42561 & ~n30371;
  assign n30374 = ~n30373 & ~n30372;
  assign P1_U2847 = ~n30375 | ~n30374;
  assign n30380 = ~n30729 | ~n42540;
  assign n30378 = ~n31109 & ~n42553;
  assign n30377 = ~n42561 & ~n30376;
  assign n30379 = ~n30378 & ~n30377;
  assign P1_U2848 = ~n30380 | ~n30379;
  assign n30385 = ~n30741 | ~n42540;
  assign n30383 = ~n31118 & ~n42553;
  assign n30381 = ~P1_EBX_REG_23__SCAN_IN;
  assign n30382 = ~n42561 & ~n30381;
  assign n30384 = ~n30383 & ~n30382;
  assign P1_U2849 = ~n30385 | ~n30384;
  assign n30389 = ~n30753 | ~n42540;
  assign n30387 = ~n31138 | ~n42559;
  assign n30386 = ~n42556 | ~P1_EBX_REG_22__SCAN_IN;
  assign n30388 = n30387 & n30386;
  assign P1_U2850 = ~n30389 | ~n30388;
  assign n30395 = ~n30536 | ~n42540;
  assign n30393 = ~n30390 & ~n42553;
  assign n30391 = ~P1_EBX_REG_21__SCAN_IN;
  assign n30392 = ~n42561 & ~n30391;
  assign n30394 = ~n30393 & ~n30392;
  assign P1_U2851 = ~n30395 | ~n30394;
  assign n30547 = ~n30778;
  assign n30400 = ~n30547 | ~n42540;
  assign n30398 = ~n30396 & ~n42553;
  assign n30397 = n42556 & P1_EBX_REG_20__SCAN_IN;
  assign n30399 = ~n30398 & ~n30397;
  assign P1_U2852 = ~n30400 | ~n30399;
  assign n30404 = ~n30789 | ~n42540;
  assign n30402 = ~n31148 & ~n42553;
  assign n30401 = n42556 & P1_EBX_REG_19__SCAN_IN;
  assign n30403 = ~n30402 & ~n30401;
  assign P1_U2853 = ~n30404 | ~n30403;
  assign n30408 = ~n30803 | ~n42540;
  assign n30406 = ~n31177 & ~n42553;
  assign n30405 = n42556 & P1_EBX_REG_18__SCAN_IN;
  assign n30407 = ~n30406 & ~n30405;
  assign P1_U2854 = ~n30408 | ~n30407;
  assign n30578 = ~n30814;
  assign n30412 = ~n30578 | ~n42540;
  assign n30410 = ~n31194 & ~n42553;
  assign n30409 = n42556 & P1_EBX_REG_17__SCAN_IN;
  assign n30411 = ~n30410 & ~n30409;
  assign P1_U2855 = ~n30412 | ~n30411;
  assign n30416 = ~n30837 & ~n42562;
  assign n30414 = ~n42559 | ~n31204;
  assign n30413 = ~n42556 | ~P1_EBX_REG_16__SCAN_IN;
  assign n30415 = ~n30414 | ~n30413;
  assign P1_U2856 = n30416 | n30415;
  assign n30421 = ~n30601 | ~n42540;
  assign n30419 = ~n42553 & ~n31222;
  assign n30417 = ~P1_EBX_REG_15__SCAN_IN;
  assign n30418 = ~n42561 & ~n30417;
  assign n30420 = ~n30419 & ~n30418;
  assign P1_U2857 = ~n30421 | ~n30420;
  assign n30425 = ~n30869 & ~n42562;
  assign n30423 = ~n42559 | ~n31236;
  assign n30422 = ~n42556 | ~P1_EBX_REG_14__SCAN_IN;
  assign n30424 = ~n30423 | ~n30422;
  assign P1_U2858 = n30425 | n30424;
  assign n30430 = ~n30616 | ~n42540;
  assign n30428 = ~n42553 & ~n31265;
  assign n30426 = ~P1_EBX_REG_13__SCAN_IN;
  assign n30427 = ~n42561 & ~n30426;
  assign n30429 = ~n30428 & ~n30427;
  assign P1_U2859 = ~n30430 | ~n30429;
  assign n30435 = ~n22909 | ~n42540;
  assign n30433 = ~n42553 & ~n31290;
  assign n30431 = ~P1_EBX_REG_12__SCAN_IN;
  assign n30432 = ~n42561 & ~n30431;
  assign n30434 = ~n30433 & ~n30432;
  assign P1_U2860 = ~n30435 | ~n30434;
  assign n30439 = ~n30919 & ~n42562;
  assign n30437 = ~n42559 | ~n31303;
  assign n30436 = ~n42556 | ~P1_EBX_REG_11__SCAN_IN;
  assign n30438 = ~n30437 | ~n30436;
  assign P1_U2861 = n30439 | n30438;
  assign n30452 = ~n30441 | ~n44865;
  assign n30442 = ~n43161 | ~n31515;
  assign n30592 = ~n42625 & ~n30442;
  assign n30444 = ~n43060 | ~BUF1_REG_14__SCAN_IN;
  assign n30443 = ~n43062 | ~DATAI_14_;
  assign n42818 = ~n30444 | ~n30443;
  assign n30446 = ~n30592 | ~n42818;
  assign n30445 = ~n26954 | ~DATAI_30_;
  assign n30450 = ~n30446 | ~n30445;
  assign n30448 = ~n26956 | ~BUF1_REG_30__SCAN_IN;
  assign n30447 = ~n42625 | ~P1_EAX_REG_30__SCAN_IN;
  assign n30449 = ~n30448 | ~n30447;
  assign n30451 = ~n30450 & ~n30449;
  assign P1_U2874 = ~n30452 | ~n30451;
  assign n30462 = ~n30657 | ~n30615;
  assign n30454 = ~n43060 | ~BUF1_REG_13__SCAN_IN;
  assign n30453 = ~n43062 | ~DATAI_13_;
  assign n30617 = ~n30454 | ~n30453;
  assign n30456 = ~n30592 | ~n30617;
  assign n30455 = ~n26954 | ~DATAI_29_;
  assign n30460 = ~n30456 | ~n30455;
  assign n30458 = ~n26956 | ~BUF1_REG_29__SCAN_IN;
  assign n30457 = ~n42625 | ~P1_EAX_REG_29__SCAN_IN;
  assign n30459 = ~n30458 | ~n30457;
  assign n30461 = ~n30460 & ~n30459;
  assign P1_U2875 = ~n30462 | ~n30461;
  assign n30463 = ~n30665;
  assign n30473 = ~n30463 | ~n30615;
  assign n30465 = ~n43060 | ~BUF1_REG_12__SCAN_IN;
  assign n30464 = ~n43062 | ~DATAI_12_;
  assign n30622 = ~n30465 | ~n30464;
  assign n30467 = ~n30592 | ~n30622;
  assign n30466 = ~n26954 | ~DATAI_28_;
  assign n30471 = ~n30467 | ~n30466;
  assign n30469 = ~n26956 | ~BUF1_REG_28__SCAN_IN;
  assign n30468 = ~n42625 | ~P1_EAX_REG_28__SCAN_IN;
  assign n30470 = ~n30469 | ~n30468;
  assign n30472 = ~n30471 & ~n30470;
  assign P1_U2876 = ~n30473 | ~n30472;
  assign n30483 = ~n30687 | ~n44865;
  assign n30475 = ~n43062 | ~DATAI_11_;
  assign n30474 = ~n43060 | ~BUF1_REG_11__SCAN_IN;
  assign n42805 = ~n30475 | ~n30474;
  assign n30477 = ~n30592 | ~n42805;
  assign n30476 = ~n26954 | ~DATAI_27_;
  assign n30481 = ~n30477 | ~n30476;
  assign n30479 = ~n26956 | ~BUF1_REG_27__SCAN_IN;
  assign n30478 = ~n42625 | ~P1_EAX_REG_27__SCAN_IN;
  assign n30480 = ~n30479 | ~n30478;
  assign n30482 = ~n30481 & ~n30480;
  assign P1_U2877 = ~n30483 | ~n30482;
  assign n30484 = ~n30698;
  assign n30494 = ~n30484 | ~n44865;
  assign n30486 = ~n43062 | ~DATAI_10_;
  assign n30485 = ~n43060 | ~BUF1_REG_10__SCAN_IN;
  assign n42800 = ~n30486 | ~n30485;
  assign n30488 = ~n30592 | ~n42800;
  assign n30487 = ~n26954 | ~DATAI_26_;
  assign n30492 = ~n30488 | ~n30487;
  assign n30490 = ~n26956 | ~BUF1_REG_26__SCAN_IN;
  assign n30489 = ~n42625 | ~P1_EAX_REG_26__SCAN_IN;
  assign n30491 = ~n30490 | ~n30489;
  assign n30493 = ~n30492 & ~n30491;
  assign P1_U2878 = ~n30494 | ~n30493;
  assign n30505 = ~n30495 | ~n30615;
  assign n30497 = ~n43062 | ~DATAI_9_;
  assign n30496 = ~n43060 | ~BUF1_REG_9__SCAN_IN;
  assign n42795 = ~n30497 | ~n30496;
  assign n30499 = ~n30592 | ~n42795;
  assign n30498 = ~n26954 | ~DATAI_25_;
  assign n30503 = ~n30499 | ~n30498;
  assign n30501 = ~n26956 | ~BUF1_REG_25__SCAN_IN;
  assign n30500 = ~n42625 | ~P1_EAX_REG_25__SCAN_IN;
  assign n30502 = ~n30501 | ~n30500;
  assign n30504 = ~n30503 & ~n30502;
  assign P1_U2879 = ~n30505 | ~n30504;
  assign n30515 = ~n30729 | ~n30615;
  assign n30507 = ~n43062 | ~DATAI_8_;
  assign n30506 = ~n43060 | ~BUF1_REG_8__SCAN_IN;
  assign n42790 = ~n30507 | ~n30506;
  assign n30509 = ~n30592 | ~n42790;
  assign n30508 = ~n26954 | ~DATAI_24_;
  assign n30513 = ~n30509 | ~n30508;
  assign n30511 = ~n26956 | ~BUF1_REG_24__SCAN_IN;
  assign n30510 = ~n42625 | ~P1_EAX_REG_24__SCAN_IN;
  assign n30512 = ~n30511 | ~n30510;
  assign n30514 = ~n30513 & ~n30512;
  assign P1_U2880 = ~n30515 | ~n30514;
  assign n30525 = ~n30741 | ~n44865;
  assign n30517 = ~n43062 | ~DATAI_7_;
  assign n30516 = ~n43060 | ~BUF1_REG_7__SCAN_IN;
  assign n42785 = ~n30517 | ~n30516;
  assign n30519 = ~n30592 | ~n42785;
  assign n30518 = ~n26954 | ~DATAI_23_;
  assign n30523 = ~n30519 | ~n30518;
  assign n30521 = ~n26956 | ~BUF1_REG_23__SCAN_IN;
  assign n30520 = ~n42625 | ~P1_EAX_REG_23__SCAN_IN;
  assign n30522 = ~n30521 | ~n30520;
  assign n30524 = ~n30523 & ~n30522;
  assign P1_U2881 = ~n30525 | ~n30524;
  assign n30535 = ~n30753 | ~n44865;
  assign n30527 = ~n43062 | ~DATAI_6_;
  assign n30526 = ~n43060 | ~BUF1_REG_6__SCAN_IN;
  assign n42781 = ~n30527 | ~n30526;
  assign n30529 = ~n30592 | ~n42781;
  assign n30528 = ~n26954 | ~DATAI_22_;
  assign n30533 = ~n30529 | ~n30528;
  assign n30531 = ~n26956 | ~BUF1_REG_22__SCAN_IN;
  assign n30530 = ~n42625 | ~P1_EAX_REG_22__SCAN_IN;
  assign n30532 = ~n30531 | ~n30530;
  assign n30534 = ~n30533 & ~n30532;
  assign P1_U2882 = ~n30535 | ~n30534;
  assign n30546 = ~n30536 | ~n30615;
  assign n30538 = ~n43062 | ~DATAI_5_;
  assign n30537 = ~n43060 | ~BUF1_REG_5__SCAN_IN;
  assign n42777 = ~n30538 | ~n30537;
  assign n30540 = ~n30592 | ~n42777;
  assign n30539 = ~n26954 | ~DATAI_21_;
  assign n30544 = ~n30540 | ~n30539;
  assign n30542 = ~n26956 | ~BUF1_REG_21__SCAN_IN;
  assign n30541 = ~n42625 | ~P1_EAX_REG_21__SCAN_IN;
  assign n30543 = ~n30542 | ~n30541;
  assign n30545 = ~n30544 & ~n30543;
  assign P1_U2883 = ~n30546 | ~n30545;
  assign n30557 = ~n30547 | ~n30615;
  assign n30549 = ~n43062 | ~DATAI_4_;
  assign n30548 = ~n43060 | ~BUF1_REG_4__SCAN_IN;
  assign n42598 = ~n30549 | ~n30548;
  assign n30551 = ~n30592 | ~n42598;
  assign n30550 = ~n26954 | ~DATAI_20_;
  assign n30555 = ~n30551 | ~n30550;
  assign n30553 = ~n26956 | ~BUF1_REG_20__SCAN_IN;
  assign n30552 = ~n42625 | ~P1_EAX_REG_20__SCAN_IN;
  assign n30554 = ~n30553 | ~n30552;
  assign n30556 = ~n30555 & ~n30554;
  assign P1_U2884 = ~n30557 | ~n30556;
  assign n30567 = ~n30789 | ~n44865;
  assign n30559 = ~n43062 | ~DATAI_3_;
  assign n30558 = ~n43060 | ~BUF1_REG_3__SCAN_IN;
  assign n42604 = ~n30559 | ~n30558;
  assign n30561 = ~n30592 | ~n42604;
  assign n30560 = ~n26954 | ~DATAI_19_;
  assign n30565 = ~n30561 | ~n30560;
  assign n30563 = ~n26956 | ~BUF1_REG_19__SCAN_IN;
  assign n30562 = ~n42625 | ~P1_EAX_REG_19__SCAN_IN;
  assign n30564 = ~n30563 | ~n30562;
  assign n30566 = ~n30565 & ~n30564;
  assign P1_U2885 = ~n30567 | ~n30566;
  assign n30577 = ~n30803 | ~n44865;
  assign n30569 = ~n43062 | ~DATAI_2_;
  assign n30568 = ~n43060 | ~BUF1_REG_2__SCAN_IN;
  assign n42610 = ~n30569 | ~n30568;
  assign n30571 = ~n30592 | ~n42610;
  assign n30570 = ~n26954 | ~DATAI_18_;
  assign n30575 = ~n30571 | ~n30570;
  assign n30573 = ~n26956 | ~BUF1_REG_18__SCAN_IN;
  assign n30572 = ~n42625 | ~P1_EAX_REG_18__SCAN_IN;
  assign n30574 = ~n30573 | ~n30572;
  assign n30576 = ~n30575 & ~n30574;
  assign P1_U2886 = ~n30577 | ~n30576;
  assign n30588 = ~n30578 | ~n30615;
  assign n30580 = ~n43062 | ~DATAI_1_;
  assign n30579 = ~n43060 | ~BUF1_REG_1__SCAN_IN;
  assign n42615 = ~n30580 | ~n30579;
  assign n30582 = ~n30592 | ~n42615;
  assign n30581 = ~n26954 | ~DATAI_17_;
  assign n30586 = ~n30582 | ~n30581;
  assign n30584 = ~n26956 | ~BUF1_REG_17__SCAN_IN;
  assign n30583 = ~n42625 | ~P1_EAX_REG_17__SCAN_IN;
  assign n30585 = ~n30584 | ~n30583;
  assign n30587 = ~n30586 & ~n30585;
  assign P1_U2887 = ~n30588 | ~n30587;
  assign n30600 = ~n30589 | ~n44865;
  assign n30591 = ~n43062 | ~DATAI_0_;
  assign n30590 = ~n43060 | ~BUF1_REG_0__SCAN_IN;
  assign n42620 = ~n30591 | ~n30590;
  assign n30594 = ~n30592 | ~n42620;
  assign n30593 = ~n26954 | ~DATAI_16_;
  assign n30598 = ~n30594 | ~n30593;
  assign n30596 = ~n26956 | ~BUF1_REG_16__SCAN_IN;
  assign n30595 = ~n42625 | ~P1_EAX_REG_16__SCAN_IN;
  assign n30597 = ~n30596 | ~n30595;
  assign n30599 = ~n30598 & ~n30597;
  assign P1_U2888 = ~n30600 | ~n30599;
  assign n30610 = ~n30601 | ~n44865;
  assign n30603 = ~n30602;
  assign n30605 = ~n43060 | ~BUF1_REG_15__SCAN_IN;
  assign n30604 = ~n43062 | ~DATAI_15_;
  assign n42887 = n30605 & n30604;
  assign n30608 = ~n42621 & ~n42887;
  assign n30607 = ~n42599 & ~n30606;
  assign n30609 = ~n30608 & ~n30607;
  assign P1_U2889 = ~n30610 | ~n30609;
  assign n30614 = ~n30869 & ~n42622;
  assign n30612 = ~n42592 | ~n42818;
  assign n30611 = ~n42625 | ~P1_EAX_REG_14__SCAN_IN;
  assign n30613 = ~n30612 | ~n30611;
  assign P1_U2890 = n30614 | n30613;
  assign n30621 = ~n30616 | ~n44865;
  assign n42814 = ~n30617;
  assign n30619 = ~n42621 & ~n42814;
  assign n30618 = ~n42599 & ~n42877;
  assign n30620 = ~n30619 & ~n30618;
  assign P1_U2891 = ~n30621 | ~n30620;
  assign n30626 = ~n22909 | ~n44865;
  assign n42810 = ~n30622;
  assign n30624 = ~n42621 & ~n42810;
  assign n30623 = ~n42599 & ~n42872;
  assign n30625 = ~n30624 & ~n30623;
  assign P1_U2892 = ~n30626 | ~n30625;
  assign n30630 = ~n30919 & ~n42622;
  assign n30628 = ~n42592 | ~n42805;
  assign n30627 = ~n42625 | ~P1_EAX_REG_11__SCAN_IN;
  assign n30629 = ~n30628 | ~n30627;
  assign P1_U2893 = n30630 | n30629;
  assign n44791 = ~n44800 | ~P1_STATEBS16_REG_SCAN_IN;
  assign n30631 = ~n44851 | ~P1_STATE2_REG_1__SCAN_IN;
  assign n30643 = ~n30632 & ~n43061;
  assign n44837 = ~n30634 | ~n44418;
  assign n30635 = ~n44837 | ~n44851;
  assign n30636 = ~n42937 | ~P1_PHYADDRPOINTER_REG_31__SCAN_IN;
  assign n30641 = n30637 & n30636;
  assign n31571 = ~n44851 | ~P1_STATE2_REG_2__SCAN_IN;
  assign n30638 = ~n44765 | ~P1_STATE2_REG_1__SCAN_IN;
  assign n42944 = n31571 & n30638;
  assign n30640 = ~n42895 | ~n30639;
  assign n30642 = ~n30641 | ~n30640;
  assign n30651 = ~n30645 & ~n43061;
  assign n31034 = ~n42929 | ~P1_REIP_REG_30__SCAN_IN;
  assign n30646 = ~n42937 | ~P1_PHYADDRPOINTER_REG_30__SCAN_IN;
  assign n30649 = n31034 & n30646;
  assign n30648 = ~n42895 | ~n30647;
  assign n30650 = ~n30649 | ~n30648;
  assign n30656 = ~n30651 & ~n30650;
  assign n30664 = ~n23166 ^ P1_INSTADDRPOINTER_REG_29__SCAN_IN;
  assign n30653 = ~n30652 | ~n23166;
  assign P1_U2969 = ~n30656 | ~n30655;
  assign n30661 = ~n42936 & ~n30658;
  assign n31038 = ~n42929 | ~P1_REIP_REG_29__SCAN_IN;
  assign n30659 = ~n42937 | ~P1_PHYADDRPOINTER_REG_29__SCAN_IN;
  assign n30660 = ~n31038 | ~n30659;
  assign n30662 = ~n30661 & ~n30660;
  assign n30672 = ~n30665 & ~n43061;
  assign n31052 = ~n42947 & ~n44681;
  assign n30667 = ~n42945 & ~n30666;
  assign n30670 = ~n31052 & ~n30667;
  assign n30669 = ~n42907 | ~n30668;
  assign n30671 = ~n30670 | ~n30669;
  assign n30686 = ~n30672 & ~n30671;
  assign n30675 = ~n30706 | ~n31078;
  assign n30678 = ~n30676 & ~n30675;
  assign n30705 = ~n30676;
  assign n30677 = ~n30705 & ~n31063;
  assign n30682 = ~n30678 & ~n30677;
  assign n30680 = ~n23742 & ~n31078;
  assign n30679 = ~n23166 & ~P1_INSTADDRPOINTER_REG_27__SCAN_IN;
  assign n30681 = ~n30680 & ~n30679;
  assign n31046 = ~n30684 ^ n30683;
  assign n30685 = ~n31046 | ~n42949;
  assign P1_U2971 = ~n30686 | ~n30685;
  assign n30693 = ~n30687 | ~n42915;
  assign n30691 = ~n42936 & ~n30688;
  assign n31065 = ~n42929 | ~P1_REIP_REG_27__SCAN_IN;
  assign n30689 = ~n42937 | ~P1_PHYADDRPOINTER_REG_27__SCAN_IN;
  assign n30690 = ~n31065 | ~n30689;
  assign n30692 = ~n30691 & ~n30690;
  assign n30697 = ~n30693 | ~n30692;
  assign n30694 = ~n23166 ^ P1_INSTADDRPOINTER_REG_27__SCAN_IN;
  assign n31070 = ~n22854 ^ n30694;
  assign n30696 = ~n31070 & ~n42932;
  assign P1_U2972 = n30697 | n30696;
  assign n30704 = ~n30698 & ~n43061;
  assign n31083 = ~n42929 | ~P1_REIP_REG_26__SCAN_IN;
  assign n30699 = ~n42937 | ~P1_PHYADDRPOINTER_REG_26__SCAN_IN;
  assign n30702 = n31083 & n30699;
  assign n30701 = ~n42907 | ~n30700;
  assign n30703 = ~n30702 | ~n30701;
  assign n30712 = ~n30704 & ~n30703;
  assign n30709 = ~n30705 & ~n23742;
  assign n30707 = ~n23742 | ~n30706;
  assign n30708 = ~n22855 & ~n30707;
  assign n30710 = ~n30709 & ~n30708;
  assign n31073 = ~n30710 ^ P1_INSTADDRPOINTER_REG_26__SCAN_IN;
  assign n30711 = ~n31073 | ~n42949;
  assign P1_U2973 = ~n30712 | ~n30711;
  assign n30720 = ~n30713 & ~n43061;
  assign n31093 = ~n42947 & ~n44666;
  assign n30714 = ~P1_PHYADDRPOINTER_REG_25__SCAN_IN;
  assign n30715 = ~n42945 & ~n30714;
  assign n30718 = ~n31093 & ~n30715;
  assign n30717 = ~n42895 | ~n30716;
  assign n30719 = ~n30718 | ~n30717;
  assign n30728 = ~n30720 & ~n30719;
  assign n30742 = ~n23166 ^ P1_INSTADDRPOINTER_REG_23__SCAN_IN;
  assign n30722 = ~n22855 | ~n30742;
  assign n30721 = ~n23742 | ~P1_INSTADDRPOINTER_REG_23__SCAN_IN;
  assign n30731 = ~n30722 | ~n30721;
  assign n30730 = ~n23166 ^ P1_INSTADDRPOINTER_REG_24__SCAN_IN;
  assign n30724 = ~n30731 | ~n30730;
  assign n30723 = ~n23742 | ~P1_INSTADDRPOINTER_REG_24__SCAN_IN;
  assign n30726 = ~n30724 | ~n30723;
  assign n30725 = P1_INSTADDRPOINTER_REG_25__SCAN_IN ^ n23166;
  assign n31089 = ~n30726 ^ n30725;
  assign n30727 = ~n31089 | ~n42949;
  assign P1_U2974 = ~n30728 | ~n30727;
  assign n30740 = ~n30729 | ~n42915;
  assign n31101 = ~n30731 ^ n30730;
  assign n30738 = ~n31101 & ~n42932;
  assign n31110 = ~n42947 & ~n44661;
  assign n30733 = ~n31110;
  assign n30732 = ~n42937 | ~P1_PHYADDRPOINTER_REG_24__SCAN_IN;
  assign n30736 = n30733 & n30732;
  assign n30735 = ~n42895 | ~n30734;
  assign n30737 = ~n30736 | ~n30735;
  assign n30739 = ~n30738 & ~n30737;
  assign P1_U2975 = ~n30740 | ~n30739;
  assign n30752 = ~n30741 | ~n42915;
  assign n30750 = ~n31116 & ~n42932;
  assign n31122 = ~n42929 | ~P1_REIP_REG_23__SCAN_IN;
  assign n30745 = ~n31122;
  assign n30744 = ~n42945 & ~n30743;
  assign n30748 = ~n30745 & ~n30744;
  assign n30747 = ~n42907 | ~n30746;
  assign n30749 = ~n30748 | ~n30747;
  assign n30751 = ~n30750 & ~n30749;
  assign P1_U2976 = ~n30752 | ~n30751;
  assign n30764 = ~n30753 | ~n42915;
  assign n31129 = ~n30754 ^ P1_INSTADDRPOINTER_REG_22__SCAN_IN;
  assign n30762 = ~n31129 & ~n42932;
  assign n31139 = ~n42929 | ~P1_REIP_REG_22__SCAN_IN;
  assign n30757 = ~n31139;
  assign n30755 = ~P1_PHYADDRPOINTER_REG_22__SCAN_IN;
  assign n30756 = ~n42945 & ~n30755;
  assign n30760 = ~n30757 & ~n30756;
  assign n30759 = ~n42895 | ~n30758;
  assign n30761 = ~n30760 | ~n30759;
  assign n30763 = ~n30762 & ~n30761;
  assign P1_U2977 = ~n30764 | ~n30763;
  assign n30774 = ~n30765 & ~n43061;
  assign n30769 = ~n30766;
  assign n30768 = ~n42945 & ~n30767;
  assign n30772 = ~n30769 & ~n30768;
  assign n30771 = ~n42895 | ~n30770;
  assign n30773 = ~n30772 | ~n30771;
  assign n30777 = ~n30774 & ~n30773;
  assign n30776 = ~n30775 | ~n42949;
  assign P1_U2978 = ~n30777 | ~n30776;
  assign n30785 = ~n30778 & ~n43061;
  assign n30779 = ~n42937 | ~P1_PHYADDRPOINTER_REG_20__SCAN_IN;
  assign n30783 = n30780 & n30779;
  assign n30782 = ~n42895 | ~n30781;
  assign n30784 = ~n30783 | ~n30782;
  assign n30788 = ~n30785 & ~n30784;
  assign n30787 = ~n30786 | ~n42949;
  assign P1_U2979 = ~n30788 | ~n30787;
  assign n30802 = ~n30789 | ~n42915;
  assign n31146 = ~n30791 ^ n30790;
  assign n30800 = ~n31146 & ~n42932;
  assign n31154 = ~n42929 | ~P1_REIP_REG_19__SCAN_IN;
  assign n30794 = ~n31154;
  assign n30793 = ~n42945 & ~n30792;
  assign n30798 = ~n30794 & ~n30793;
  assign n30796 = ~n30795;
  assign n30797 = ~n42907 | ~n30796;
  assign n30799 = ~n30798 | ~n30797;
  assign n30801 = ~n30800 & ~n30799;
  assign P1_U2980 = ~n30802 | ~n30801;
  assign n30813 = ~n30803 | ~n42915;
  assign n31183 = ~n30805 ^ n30804;
  assign n30811 = ~n31183 & ~n42932;
  assign n31179 = ~n42929 | ~P1_REIP_REG_18__SCAN_IN;
  assign n30806 = ~n42937 | ~P1_PHYADDRPOINTER_REG_18__SCAN_IN;
  assign n30809 = n31179 & n30806;
  assign n30808 = ~n42907 | ~n30807;
  assign n30810 = ~n30809 | ~n30808;
  assign n30812 = ~n30811 & ~n30810;
  assign P1_U2981 = ~n30813 | ~n30812;
  assign n30820 = ~n30814 & ~n43061;
  assign n30818 = ~n42936 & ~n30815;
  assign n31196 = ~n42929 | ~P1_REIP_REG_17__SCAN_IN;
  assign n30816 = ~n42937 | ~P1_PHYADDRPOINTER_REG_17__SCAN_IN;
  assign n30817 = ~n31196 | ~n30816;
  assign n30819 = n30818 | n30817;
  assign n30836 = ~n30820 & ~n30819;
  assign n30822 = ~n23166 & ~n31189;
  assign n30834 = ~n30823 & ~n30822;
  assign n30830 = ~n30824 & ~n30825;
  assign n30827 = ~n30826;
  assign n30829 = ~n30828 | ~n30827;
  assign n30832 = n30830 | n30829;
  assign n30831 = ~n23742 | ~P1_INSTADDRPOINTER_REG_16__SCAN_IN;
  assign n30833 = ~n30832 | ~n30831;
  assign n31186 = n30834 ^ n30833;
  assign n30835 = ~n31186 | ~n42949;
  assign P1_U2982 = ~n30836 | ~n30835;
  assign n30843 = ~n30837 & ~n43061;
  assign n31207 = ~n42929 | ~P1_REIP_REG_16__SCAN_IN;
  assign n30838 = ~n42937 | ~P1_PHYADDRPOINTER_REG_16__SCAN_IN;
  assign n30841 = n31207 & n30838;
  assign n30840 = ~n42895 | ~n30839;
  assign n30842 = ~n30841 | ~n30840;
  assign n30853 = ~n30843 & ~n30842;
  assign n30929 = ~n30824;
  assign n30848 = n30929 | n30845;
  assign n30847 = ~n23730 & ~n30846;
  assign n30866 = ~n30848 | ~n30847;
  assign n30850 = ~n30866 & ~n30849;
  assign n31202 = ~n30844 ^ n30851;
  assign n30852 = ~n31202 | ~n42949;
  assign P1_U2983 = ~n30853 | ~n30852;
  assign n30863 = ~n30854 & ~n43061;
  assign n31224 = ~n42929 | ~P1_REIP_REG_15__SCAN_IN;
  assign n30857 = ~n31224;
  assign n30856 = ~n42945 & ~n30855;
  assign n30861 = ~n30857 & ~n30856;
  assign n30859 = ~n30858;
  assign n30860 = ~n42895 | ~n30859;
  assign n30862 = ~n30861 | ~n30860;
  assign n30868 = ~n30863 & ~n30862;
  assign n30865 = ~n30849 & ~n30864;
  assign n31214 = n30866 ^ n30865;
  assign n30867 = ~n31214 | ~n42949;
  assign P1_U2984 = ~n30868 | ~n30867;
  assign n30876 = n30869 | n43061;
  assign n31237 = ~n42929 | ~P1_REIP_REG_14__SCAN_IN;
  assign n30870 = ~n42937 | ~P1_PHYADDRPOINTER_REG_14__SCAN_IN;
  assign n30874 = ~n31237 | ~n30870;
  assign n30872 = ~n30871;
  assign n30873 = n42895 & n30872;
  assign n30875 = ~n30874 & ~n30873;
  assign n30888 = ~n30876 | ~n30875;
  assign n30882 = ~n30929 | ~n30877;
  assign n30880 = ~n30878;
  assign n30881 = ~n30880 & ~n30879;
  assign n30884 = ~n30882 | ~n30881;
  assign n30886 = ~n30884 | ~n30883;
  assign n30885 = ~n30953 ^ P1_INSTADDRPOINTER_REG_14__SCAN_IN;
  assign n31255 = ~n30886 ^ n30885;
  assign n30887 = ~n31255 & ~n42932;
  assign P1_U2985 = n30888 | n30887;
  assign n30897 = ~n30889 & ~n43061;
  assign n30890 = ~P1_REIP_REG_13__SCAN_IN;
  assign n31266 = ~n42947 & ~n30890;
  assign n30892 = ~n42945 & ~n30891;
  assign n30895 = ~n31266 & ~n30892;
  assign n30894 = ~n42907 | ~n30893;
  assign n30896 = ~n30895 | ~n30894;
  assign n30906 = ~n30897 & ~n30896;
  assign n30901 = ~n30929 & ~n30879;
  assign n30900 = ~n30899 | ~n30898;
  assign n30909 = ~n30901 & ~n30900;
  assign n30902 = ~n30909 | ~n30908;
  assign n30904 = ~n30902 | ~n30907;
  assign n31258 = ~n30904 ^ n30903;
  assign n30905 = ~n31258 | ~n42949;
  assign P1_U2986 = ~n30906 | ~n30905;
  assign n30918 = ~n22909 | ~n42915;
  assign n30910 = ~n30908 | ~n30907;
  assign n31276 = n30910 ^ n30909;
  assign n30916 = ~n31276 | ~n42949;
  assign n30914 = ~n42936 & ~n30911;
  assign n31292 = ~n42929 | ~P1_REIP_REG_12__SCAN_IN;
  assign n30912 = ~n42937 | ~P1_PHYADDRPOINTER_REG_12__SCAN_IN;
  assign n30913 = ~n31292 | ~n30912;
  assign n30915 = ~n30914 & ~n30913;
  assign n30917 = n30916 & n30915;
  assign P1_U2987 = ~n30918 | ~n30917;
  assign n30925 = ~n30919 & ~n43061;
  assign n31304 = ~n42929 | ~P1_REIP_REG_11__SCAN_IN;
  assign n30920 = ~n42937 | ~P1_PHYADDRPOINTER_REG_11__SCAN_IN;
  assign n30923 = n31304 & n30920;
  assign n30922 = ~n42907 | ~n30921;
  assign n30924 = ~n30923 | ~n30922;
  assign n30935 = ~n30925 & ~n30924;
  assign n30936 = ~n30824 ^ n30926;
  assign n30931 = ~n30936 & ~n30927;
  assign n30930 = ~n30929 & ~n30928;
  assign n30933 = ~n30931 & ~n30930;
  assign n30932 = ~n30953 ^ P1_INSTADDRPOINTER_REG_11__SCAN_IN;
  assign n31300 = ~n30933 ^ n30932;
  assign n30934 = ~n31300 | ~n42949;
  assign P1_U2988 = ~n30935 | ~n30934;
  assign n31329 = ~n30936 ^ P1_INSTADDRPOINTER_REG_10__SCAN_IN;
  assign n30945 = ~n31329 | ~n42949;
  assign n30943 = ~n42506 | ~n42915;
  assign n30941 = ~n42936 & ~n30937;
  assign n31323 = ~n42947 & ~n44591;
  assign n30939 = ~n31323;
  assign n30938 = ~n42937 | ~P1_PHYADDRPOINTER_REG_10__SCAN_IN;
  assign n30940 = ~n30939 | ~n30938;
  assign n30942 = ~n30941 & ~n30940;
  assign n30944 = n30943 & n30942;
  assign P1_U2989 = ~n30945 | ~n30944;
  assign n30948 = n30946;
  assign n30969 = ~n30948 | ~n30947;
  assign n30968 = ~n30950 ^ n30949;
  assign n30952 = ~n30969 | ~n30968;
  assign n30955 = ~n30952 | ~n30951;
  assign n30954 = ~n30953 ^ P1_INSTADDRPOINTER_REG_9__SCAN_IN;
  assign n31337 = ~n30955 ^ n30954;
  assign n30967 = ~n31337 & ~n42932;
  assign n30959 = n30957 & n30956;
  assign n42572 = n30959 | n30958;
  assign n30960 = ~n42572;
  assign n30965 = ~n30960 | ~n42915;
  assign n30963 = ~n42936 & ~n42290;
  assign n31339 = ~n42929 | ~P1_REIP_REG_9__SCAN_IN;
  assign n30961 = ~n42937 | ~P1_PHYADDRPOINTER_REG_9__SCAN_IN;
  assign n30962 = ~n31339 | ~n30961;
  assign n30964 = ~n30963 & ~n30962;
  assign n30966 = ~n30965 | ~n30964;
  assign P1_U2990 = n30967 | n30966;
  assign n31346 = ~n30969 ^ n30968;
  assign n30979 = ~n31346 & ~n42932;
  assign n42579 = n30971 ^ n30984;
  assign n30977 = ~n42579 | ~n42915;
  assign n30972 = ~n42306;
  assign n30975 = ~n42936 & ~n30972;
  assign n31353 = ~n42929 | ~P1_REIP_REG_8__SCAN_IN;
  assign n30973 = ~n42937 | ~P1_PHYADDRPOINTER_REG_8__SCAN_IN;
  assign n30974 = ~n31353 | ~n30973;
  assign n30976 = ~n30975 & ~n30974;
  assign n30978 = ~n30977 | ~n30976;
  assign P1_U2991 = n30979 | n30978;
  assign n30991 = ~n31375 & ~n42932;
  assign n30983 = ~n30981 | ~n30982;
  assign n30989 = ~n42326 | ~n42915;
  assign n30987 = ~n42936 & ~n42327;
  assign n31371 = ~n42929 | ~P1_REIP_REG_7__SCAN_IN;
  assign n30985 = ~n42937 | ~P1_PHYADDRPOINTER_REG_7__SCAN_IN;
  assign n30986 = ~n31371 | ~n30985;
  assign n30988 = ~n30987 & ~n30986;
  assign n30990 = ~n30989 | ~n30988;
  assign P1_U2992 = n30991 | n30990;
  assign n30998 = ~n30992 & ~n23494;
  assign n30996 = n30995 & n30994;
  assign n30997 = ~n30993 & ~n30996;
  assign n31387 = ~n30998 & ~n30997;
  assign n31008 = ~n31387 & ~n42932;
  assign n31001 = n31000 | n30999;
  assign n42587 = ~n30981 | ~n31001;
  assign n31006 = n42587 | n43061;
  assign n31389 = ~n42929 | ~P1_REIP_REG_6__SCAN_IN;
  assign n31002 = ~n42937 | ~P1_PHYADDRPOINTER_REG_6__SCAN_IN;
  assign n31004 = ~n31389 | ~n31002;
  assign n31003 = n42895 & n42350;
  assign n31005 = ~n31004 & ~n31003;
  assign n31007 = ~n31006 | ~n31005;
  assign P1_U2993 = n31008 | n31007;
  assign n42921 = ~n31009 ^ P1_INSTADDRPOINTER_REG_2__SCAN_IN;
  assign n31011 = ~n42921 | ~n42920;
  assign n31013 = ~n31011 | ~n31010;
  assign n42910 = P1_INSTADDRPOINTER_REG_3__SCAN_IN ^ n31013;
  assign n31015 = ~n42910 | ~n31012;
  assign n31014 = ~n31013 | ~P1_INSTADDRPOINTER_REG_3__SCAN_IN;
  assign n31016 = ~n31015 | ~n31014;
  assign n42898 = P1_INSTADDRPOINTER_REG_4__SCAN_IN ^ n31016;
  assign n31018 = ~n42898 | ~n23083;
  assign n31017 = ~n31016 | ~P1_INSTADDRPOINTER_REG_4__SCAN_IN;
  assign n31020 = ~n31018 | ~n31017;
  assign n31411 = ~n31020 ^ n31019;
  assign n31030 = ~n31411 | ~n42949;
  assign n42371 = ~n31021 ^ n31022;
  assign n31028 = ~n42371 & ~n43061;
  assign n31398 = ~n42947 & ~n44566;
  assign n31024 = ~n42945 & ~n31023;
  assign n31026 = ~n31398 & ~n31024;
  assign n31025 = ~n42895 | ~n42363;
  assign n31027 = ~n31026 | ~n31025;
  assign n31029 = ~n31028 & ~n31027;
  assign P1_U2994 = ~n31030 | ~n31029;
  assign n31041 = ~P1_INSTADDRPOINTER_REG_29__SCAN_IN & ~n31036;
  assign n31039 = n31037 | n43001;
  assign n31040 = ~n31039 | ~n31038;
  assign n31042 = n31041 | n31040;
  assign n31044 = ~n31043 & ~n31042;
  assign P1_U3002 = ~n31045 | ~n31044;
  assign n31058 = ~n31046 | ~n43042;
  assign n31056 = n31059 & P1_INSTADDRPOINTER_REG_28__SCAN_IN;
  assign n31054 = ~n31047 | ~n25838;
  assign n31050 = ~n31048 | ~n31062;
  assign n31051 = ~n31050 & ~n31049;
  assign n31053 = ~n31052 & ~n31051;
  assign n31055 = ~n31054 | ~n31053;
  assign n31057 = ~n31056 & ~n31055;
  assign P1_U3003 = ~n31058 | ~n31057;
  assign n31060 = ~n31059;
  assign n31069 = ~n31060 & ~n31063;
  assign n31067 = n31061 | n43001;
  assign n31064 = ~n31063 | ~n31062;
  assign n31066 = n31065 & n31064;
  assign n31068 = ~n31067 | ~n31066;
  assign n31072 = ~n31069 & ~n31068;
  assign n31071 = n31070 | n43018;
  assign P1_U3004 = ~n31072 | ~n31071;
  assign n31088 = ~n31073 | ~n43042;
  assign n31077 = ~n31074;
  assign n31076 = n31075 & n31090;
  assign n31095 = ~n31119 | ~n31076;
  assign n31081 = ~n31077 | ~n31095;
  assign n31080 = ~n31079 | ~n31078;
  assign n31086 = n31081 & n31080;
  assign n31084 = ~n31082 | ~n25838;
  assign n31085 = ~n31084 | ~n31083;
  assign n31087 = ~n31086 & ~n31085;
  assign P1_U3005 = ~n31088 | ~n31087;
  assign n31100 = ~n31089 | ~n43042;
  assign n31098 = ~n31091 & ~n31090;
  assign n31094 = ~n31092 & ~n43001;
  assign n31096 = ~n31094 & ~n31093;
  assign n31097 = ~n31096 | ~n31095;
  assign n31099 = ~n31098 & ~n31097;
  assign P1_U3006 = ~n31100 | ~n31099;
  assign n31115 = ~n31101 & ~n43018;
  assign n31103 = ~P1_INSTADDRPOINTER_REG_23__SCAN_IN & ~n31102;
  assign n31104 = ~n31117 & ~n31103;
  assign n31108 = ~n31104 | ~P1_INSTADDRPOINTER_REG_24__SCAN_IN;
  assign n31106 = ~n31119 | ~P1_INSTADDRPOINTER_REG_23__SCAN_IN;
  assign n31107 = ~n31106 | ~n31105;
  assign n31113 = ~n31108 | ~n31107;
  assign n31111 = ~n31109 & ~n43001;
  assign n31112 = ~n31111 & ~n31110;
  assign n31114 = ~n31113 | ~n31112;
  assign P1_U3007 = n31115 | n31114;
  assign n31128 = ~n31116 & ~n43018;
  assign n31126 = ~P1_INSTADDRPOINTER_REG_23__SCAN_IN | ~n31117;
  assign n31124 = ~n31118 & ~n43001;
  assign n31120 = ~P1_INSTADDRPOINTER_REG_23__SCAN_IN;
  assign n31121 = ~n31120 | ~n31119;
  assign n31123 = ~n31122 | ~n31121;
  assign n31125 = ~n31124 & ~n31123;
  assign n31127 = ~n31126 | ~n31125;
  assign P1_U3008 = n31128 | n31127;
  assign n31145 = ~n31129 & ~n43018;
  assign n31136 = ~P1_INSTADDRPOINTER_REG_22__SCAN_IN;
  assign n31130 = ~n31136 | ~P1_INSTADDRPOINTER_REG_21__SCAN_IN;
  assign n31133 = n31150 | n31130;
  assign n31132 = ~P1_INSTADDRPOINTER_REG_22__SCAN_IN | ~n31131;
  assign n31135 = ~n31133 | ~n31132;
  assign n31143 = ~n31135 | ~n31134;
  assign n31142 = n31137 | n31136;
  assign n31140 = ~n31138 | ~n25838;
  assign n31141 = n31140 & n31139;
  assign n31144 = ~n31143 | ~n22962;
  assign P1_U3009 = n31145 | n31144;
  assign n31160 = ~n31146 & ~n43018;
  assign n31158 = n31147 | n31151;
  assign n31149 = ~n31148;
  assign n31156 = ~n25838 | ~n31149;
  assign n31152 = ~n31150;
  assign n31153 = ~n31152 | ~n31151;
  assign n31155 = n31154 & n31153;
  assign n31157 = n31156 & n31155;
  assign n31159 = ~n31158 | ~n31157;
  assign P1_U3012 = n31160 | n31159;
  assign n42967 = ~n31230;
  assign n31164 = n42967 | n31170;
  assign n31161 = ~n31167;
  assign n31163 = ~n31162 | ~n31161;
  assign n31215 = ~n31164 | ~n31163;
  assign n31166 = ~n31215 | ~n31173;
  assign n31165 = ~P1_INSTADDRPOINTER_REG_18__SCAN_IN;
  assign n31176 = ~n31166 | ~n31165;
  assign n31168 = ~n31243 & ~n31167;
  assign n31169 = ~n42966 & ~n31168;
  assign n31172 = ~n31169 & ~n31380;
  assign n31171 = ~n31170 | ~n42961;
  assign n31218 = ~n31172 | ~n31171;
  assign n31174 = ~n43027 & ~n31173;
  assign n31191 = ~n31218 & ~n31174;
  assign n31175 = ~n31191 | ~P1_INSTADDRPOINTER_REG_18__SCAN_IN;
  assign n31182 = ~n31176 | ~n31175;
  assign n31178 = ~n31177;
  assign n31180 = ~n25838 | ~n31178;
  assign n31181 = n31180 & n31179;
  assign n31185 = ~n31182 | ~n31181;
  assign n31184 = ~n31183 & ~n43018;
  assign P1_U3013 = n31185 | n31184;
  assign n31201 = n31186 & n43042;
  assign n31188 = ~n31187;
  assign n31190 = ~n31215 | ~n31188;
  assign n31193 = ~n31190 | ~n31189;
  assign n31192 = ~n31191;
  assign n31199 = ~n31193 | ~n31192;
  assign n31195 = ~n31194;
  assign n31197 = ~n25838 | ~n31195;
  assign n31198 = n31197 & n31196;
  assign n31200 = ~n31199 | ~n31198;
  assign P1_U3014 = n31201 | n31200;
  assign n31213 = ~n31202 | ~n43042;
  assign n31203 = ~P1_INSTADDRPOINTER_REG_16__SCAN_IN ^ n31216;
  assign n31211 = ~n31215 | ~n31203;
  assign n31205 = ~n31204;
  assign n31209 = ~n43001 & ~n31205;
  assign n31206 = ~P1_INSTADDRPOINTER_REG_16__SCAN_IN | ~n31218;
  assign n31208 = ~n31207 | ~n31206;
  assign n31210 = ~n31209 & ~n31208;
  assign n31212 = n31211 & n31210;
  assign P1_U3015 = ~n31213 | ~n31212;
  assign n31229 = n31214 & n43042;
  assign n31217 = ~n31215;
  assign n31221 = ~n31217 | ~n31216;
  assign n31219 = ~n31218;
  assign n31220 = ~n31219 | ~P1_INSTADDRPOINTER_REG_15__SCAN_IN;
  assign n31227 = ~n31221 | ~n31220;
  assign n31223 = ~n31222;
  assign n31225 = ~n25838 | ~n31223;
  assign n31226 = n31225 & n31224;
  assign n31228 = ~n31227 | ~n31226;
  assign P1_U3016 = n31229 | n31228;
  assign n31283 = ~n31279 | ~n31230;
  assign n31301 = n31283 & n31231;
  assign n31289 = ~n31301;
  assign n31234 = ~n31233 | ~n31232;
  assign n31235 = ~n31234 & ~n31261;
  assign n31240 = n31289 & n31235;
  assign n31238 = ~n25838 | ~n31236;
  assign n31239 = ~n31238 | ~n31237;
  assign n31254 = ~n31240 & ~n31239;
  assign n31251 = n31259 | P1_INSTADDRPOINTER_REG_13__SCAN_IN;
  assign n31269 = ~n31242 & ~n31241;
  assign n31246 = ~n43014 | ~n31243;
  assign n31245 = ~n43013 | ~n31244;
  assign n31247 = ~n31246 | ~n31245;
  assign n31249 = ~n31269 & ~n31247;
  assign n31262 = ~n31249 | ~n31248;
  assign n31250 = ~n31262;
  assign n31252 = ~n31251 | ~n31250;
  assign n31253 = ~n31252 | ~P1_INSTADDRPOINTER_REG_14__SCAN_IN;
  assign n31257 = ~n31254 | ~n31253;
  assign n31256 = ~n31255 & ~n43018;
  assign P1_U3017 = n31257 | n31256;
  assign n31275 = ~n31258 | ~n43042;
  assign n31260 = ~n31259;
  assign n31264 = ~n31260 & ~P1_INSTADDRPOINTER_REG_13__SCAN_IN;
  assign n31263 = ~n31262 & ~n31261;
  assign n31273 = ~n31264 & ~n31263;
  assign n31267 = ~n43001 & ~n31265;
  assign n31271 = ~n31267 & ~n31266;
  assign n31270 = ~n31269 | ~n31268;
  assign n31272 = ~n31271 | ~n31270;
  assign n31274 = ~n31273 & ~n31272;
  assign P1_U3018 = ~n31275 | ~n31274;
  assign n31299 = ~n31276 | ~n43042;
  assign n31278 = ~n31277 | ~P1_INSTADDRPOINTER_REG_11__SCAN_IN;
  assign n31282 = ~n31278 | ~n43014;
  assign n31280 = ~n42960 & ~n31279;
  assign n31281 = ~n31380 & ~n31280;
  assign n31302 = ~n31282 | ~n31281;
  assign n31284 = ~P1_INSTADDRPOINTER_REG_11__SCAN_IN & ~n31283;
  assign n31285 = ~n31302 & ~n31284;
  assign n31297 = ~n31286 & ~n31285;
  assign n31288 = ~n31287 & ~P1_INSTADDRPOINTER_REG_12__SCAN_IN;
  assign n31295 = ~n31289 | ~n31288;
  assign n31291 = ~n31290;
  assign n31293 = ~n25838 | ~n31291;
  assign n31294 = n31293 & n31292;
  assign n31296 = ~n31295 | ~n31294;
  assign n31298 = ~n31297 & ~n31296;
  assign P1_U3019 = ~n31299 | ~n31298;
  assign n31311 = ~n31300 | ~n43042;
  assign n31309 = ~n31301 & ~P1_INSTADDRPOINTER_REG_11__SCAN_IN;
  assign n31307 = ~P1_INSTADDRPOINTER_REG_11__SCAN_IN | ~n31302;
  assign n31305 = ~n25838 | ~n31303;
  assign n31306 = n31305 & n31304;
  assign n31308 = ~n31307 | ~n31306;
  assign n31310 = ~n31309 & ~n31308;
  assign P1_U3020 = ~n31311 | ~n31310;
  assign n31314 = ~n31312 & ~n42967;
  assign n31313 = ~n31381 & ~n42966;
  assign n31378 = ~n31314 & ~n31313;
  assign n31362 = ~n31378 & ~n25449;
  assign n31333 = ~n31315 | ~n31362;
  assign n31316 = ~P1_INSTADDRPOINTER_REG_10__SCAN_IN ^ P1_INSTADDRPOINTER_REG_9__SCAN_IN;
  assign n31328 = ~n31333 & ~n31316;
  assign n31320 = ~n31317 | ~n42961;
  assign n31319 = ~n43014 | ~n31318;
  assign n31321 = ~n31320 | ~n31319;
  assign n31334 = ~n31380 & ~n31321;
  assign n31322 = ~n31334;
  assign n31326 = ~n31322 | ~P1_INSTADDRPOINTER_REG_10__SCAN_IN;
  assign n31324 = ~n43001 & ~n42507;
  assign n31325 = ~n31324 & ~n31323;
  assign n31327 = ~n31326 | ~n31325;
  assign n31331 = ~n31328 & ~n31327;
  assign n31330 = ~n31329 | ~n43042;
  assign P1_U3021 = ~n31331 | ~n31330;
  assign n31336 = ~n31333 | ~n31332;
  assign n31335 = ~n31334 | ~P1_INSTADDRPOINTER_REG_9__SCAN_IN;
  assign n31344 = ~n31336 | ~n31335;
  assign n31342 = ~n31337 & ~n43018;
  assign n42512 = n31338 ^ n23032;
  assign n31340 = ~n25838 | ~n42512;
  assign n31341 = ~n31340 | ~n31339;
  assign n31343 = ~n31342 & ~n31341;
  assign P1_U3022 = ~n31344 | ~n31343;
  assign n31364 = ~P1_INSTADDRPOINTER_REG_7__SCAN_IN;
  assign n31345 = ~P1_INSTADDRPOINTER_REG_8__SCAN_IN ^ n31364;
  assign n31360 = ~n31345 | ~n31362;
  assign n31358 = ~n31346 & ~n43018;
  assign n31350 = ~n31347 & ~n42960;
  assign n31349 = ~n31348 & ~n42966;
  assign n31351 = ~n31350 & ~n31349;
  assign n31361 = ~n31351 | ~n42963;
  assign n31356 = ~n31361 | ~P1_INSTADDRPOINTER_REG_8__SCAN_IN;
  assign n42518 = n31352 ^ n31370;
  assign n31354 = ~n25838 | ~n42518;
  assign n31355 = n31354 & n31353;
  assign n31357 = ~n31356 | ~n31355;
  assign n31359 = ~n31358 & ~n31357;
  assign P1_U3023 = ~n31360 | ~n31359;
  assign n31366 = n31361 | n31364;
  assign n31363 = ~n31362;
  assign n31365 = ~n31364 | ~n31363;
  assign n31374 = ~n31366 | ~n31365;
  assign n31369 = n31368 | n31367;
  assign n42323 = n31370 & n31369;
  assign n31372 = ~n25838 | ~n42323;
  assign n31373 = n31372 & n31371;
  assign n31377 = ~n31374 | ~n31373;
  assign n31376 = ~n31375 & ~n43018;
  assign P1_U3024 = n31377 | n31376;
  assign n31386 = ~n31378 | ~n25449;
  assign n31379 = ~n42960 & ~n31404;
  assign n31382 = ~n31380 & ~n31379;
  assign n31396 = ~n43014 | ~n31381;
  assign n31406 = ~n31382 | ~n31396;
  assign n31383 = ~P1_INSTADDRPOINTER_REG_5__SCAN_IN & ~n42960;
  assign n31384 = ~n31406 & ~n31383;
  assign n31385 = ~n31384 | ~P1_INSTADDRPOINTER_REG_6__SCAN_IN;
  assign n31394 = ~n31386 | ~n31385;
  assign n31392 = ~n31387 & ~n43018;
  assign n42342 = ~n31388 ^ n23067;
  assign n31390 = ~n25838 | ~n42342;
  assign n31391 = ~n31390 | ~n31389;
  assign n31393 = ~n31392 & ~n31391;
  assign P1_U3025 = ~n31394 | ~n31393;
  assign n31397 = ~n31395;
  assign n31399 = ~n31397 & ~n31396;
  assign n31403 = ~n31399 & ~n31398;
  assign n42533 = n31401 ^ n31400;
  assign n31402 = ~n25838 | ~n42533;
  assign n31410 = ~n31403 | ~n31402;
  assign n31405 = ~P1_INSTADDRPOINTER_REG_5__SCAN_IN & ~n42967;
  assign n31408 = ~n31405 | ~n31404;
  assign n31407 = ~P1_INSTADDRPOINTER_REG_5__SCAN_IN | ~n31406;
  assign n31409 = ~n31408 | ~n31407;
  assign n31413 = ~n31410 & ~n31409;
  assign n31412 = ~n31411 | ~n43042;
  assign P1_U3026 = ~n31413 | ~n31412;
  assign n31414 = ~n31451;
  assign n31425 = ~n43051 | ~n31414;
  assign n31498 = ~n31415 & ~n44845;
  assign n31416 = ~n31498;
  assign n31433 = ~n26965;
  assign n31418 = ~n31417 | ~n31433;
  assign n31421 = ~n31420 & ~n31419;
  assign n31422 = ~n43116 | ~n44842;
  assign n31430 = ~n31541 | ~n44514;
  assign n31471 = ~P1_FLUSH_REG_SCAN_IN;
  assign n31426 = n31471 | n44508;
  assign n31428 = ~n31426 | ~P1_STATE2_REG_0__SCAN_IN;
  assign n31427 = ~n44851 | ~n44766;
  assign n31429 = ~n31428 | ~n31427;
  assign n31432 = ~n31431 & ~n44142;
  assign n42390 = n31528 ^ n31432;
  assign n31434 = ~n31433 | ~n44744;
  assign n31435 = ~n42390 & ~n31434;
  assign n31437 = ~n44757 | ~n31435;
  assign n31436 = ~n44741 | ~P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN;
  assign P1_U3468 = ~n31437 | ~n31436;
  assign n31440 = n31439 & n31438;
  assign n31442 = n31441 & n31440;
  assign n31443 = ~n31442 | ~n26965;
  assign n31543 = n31444 | n31443;
  assign n31467 = ~n23619 | ~n31543;
  assign n31448 = ~n31446 | ~n31474;
  assign n31447 = ~n31536 | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n31450 = ~n31448 | ~n31447;
  assign n31452 = ~n31450 | ~n31449;
  assign n31475 = ~n31509 | ~n31451;
  assign n31458 = ~n31452 | ~n31475;
  assign n31455 = n31449 | n25184;
  assign n31453 = ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign n31454 = ~n31453 | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n31456 = ~n31455 | ~n31454;
  assign n31457 = ~n44745 | ~n31456;
  assign n31465 = ~n31458 | ~n31457;
  assign n31460 = n31474 & n25575;
  assign n31462 = ~n31461 & ~n31460;
  assign n44712 = ~n31463 | ~n31462;
  assign n31464 = ~n31476 & ~n44712;
  assign n31466 = ~n31465 & ~n31464;
  assign n44713 = ~n31467 | ~n31466;
  assign n31469 = ~n31541 | ~n44713;
  assign n31468 = ~n31524 | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n31559 = ~n31469 | ~n31468;
  assign n31470 = ~n31559;
  assign n31473 = ~n31470 & ~P1_STATE2_REG_1__SCAN_IN;
  assign n31529 = ~P1_STATE2_REG_1__SCAN_IN | ~n31471;
  assign n31472 = ~n25575 & ~n31529;
  assign n31492 = ~n31473 & ~n31472;
  assign n31487 = ~n31524 | ~n31488;
  assign n44719 = ~n31474 ^ n31488;
  assign n31485 = ~n31475 | ~n44719;
  assign n31483 = ~n31476 & ~n44719;
  assign n31477 = P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN ^ P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign n31481 = ~n44745 | ~n31477;
  assign n31479 = n31478;
  assign n44784 = ~n31479;
  assign n31480 = ~n44784 | ~n31543;
  assign n31482 = ~n31481 | ~n31480;
  assign n31484 = ~n31483 & ~n31482;
  assign n44721 = ~n31485 | ~n31484;
  assign n31486 = n31524 | n44721;
  assign n31490 = n31555 & n31580;
  assign n31489 = ~n31488 & ~n31529;
  assign n31491 = ~n31490 & ~n31489;
  assign n43046 = ~n31492 & ~n31491;
  assign n31522 = ~n43046;
  assign n31496 = ~n23147 & ~n42372;
  assign n42228 = ~n31512 & ~n31493;
  assign n31494 = ~n26962;
  assign n31495 = ~n42228 & ~n31494;
  assign n42235 = ~n31496 & ~n31495;
  assign n31499 = ~n31498 | ~n31497;
  assign n31500 = ~n31499 | ~n31582;
  assign n42248 = ~n42235 | ~n31500;
  assign n31501 = ~P1_FLUSH_REG_SCAN_IN & ~P1_MORE_REG_SCAN_IN;
  assign n31520 = ~n42248 & ~n31501;
  assign n31504 = ~n31502 | ~n25042;
  assign n31505 = ~n31504 & ~n31503;
  assign n31507 = ~n31506 & ~n31505;
  assign n31511 = ~n31508 | ~n31507;
  assign n31510 = ~n23147 | ~n31509;
  assign n31514 = ~n31511 | ~n31510;
  assign n31513 = ~n31512 | ~n25673;
  assign n31516 = ~n31514 | ~n31513;
  assign n44832 = ~n31516 | ~n31515;
  assign n31518 = ~n31517;
  assign n31519 = ~n44832 | ~n31518;
  assign n31521 = ~n31520 & ~n31519;
  assign n31533 = ~n31522 | ~n31521;
  assign n31523 = ~n42390 & ~n26965;
  assign n31527 = ~n31524 & ~n31523;
  assign n31525 = ~P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN & ~n31541;
  assign n31526 = P1_STATE2_REG_1__SCAN_IN | n31525;
  assign n31531 = ~n31527 & ~n31526;
  assign n31530 = ~n31529 & ~n31528;
  assign n43047 = ~n31531 & ~n31530;
  assign n31532 = ~n43047;
  assign n31565 = ~n31533 & ~n31532;
  assign n31540 = ~n31534 | ~n31543;
  assign n31538 = ~n31535 & ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign n44729 = n31536 | n24764;
  assign n31537 = ~n25660 & ~n44729;
  assign n31539 = ~n31538 & ~n31537;
  assign n44732 = ~n31540 | ~n31539;
  assign n31542 = ~n31541 | ~n44732;
  assign n31552 = ~P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~n31542;
  assign n31549 = ~P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & ~n31542;
  assign n31544 = ~n31543;
  assign n31546 = ~n43379 & ~n31544;
  assign n31545 = ~n25660 & ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN;
  assign n44749 = ~n31546 & ~n31545;
  assign n31547 = ~n44745 | ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN;
  assign n31548 = ~n44749 | ~n31547;
  assign n31550 = ~n31549 & ~n31548;
  assign n31551 = ~P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN | ~n31550;
  assign n31553 = ~n31552 | ~n31551;
  assign n31557 = P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN | n31553;
  assign n31554 = ~P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN | ~n31553;
  assign n31556 = ~n31555 | ~n31554;
  assign n31560 = ~n31557 | ~n31556;
  assign n31558 = ~n31560 & ~n31559;
  assign n31563 = ~n31558 & ~P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN;
  assign n31561 = ~n31560 | ~n31559;
  assign n31562 = ~P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | ~n31561;
  assign n31564 = ~n31563 | ~n31562;
  assign n31567 = ~n44841 & ~n31566;
  assign n31569 = n31568 & n31567;
  assign n31576 = ~n31570 | ~n31569;
  assign n31572 = ~n31571;
  assign n31574 = ~n44850 | ~n31572;
  assign n31575 = ~n31574 | ~n31573;
  assign n31587 = ~n31576 | ~n31575;
  assign n44517 = ~n44512 & ~n44851;
  assign n31578 = ~n44766 & ~n44853;
  assign n31577 = ~P1_STATE2_REG_2__SCAN_IN & ~n31582;
  assign n31579 = ~n31578 & ~n31577;
  assign n31589 = ~n44510 | ~n31580;
  assign n31581 = ~n44851 & ~P1_STATE2_REG_2__SCAN_IN;
  assign n31584 = ~n31582 | ~n31581;
  assign n31583 = ~n44851 | ~P1_STATEBS16_REG_SCAN_IN;
  assign n31585 = ~n31584 | ~n31583;
  assign n44519 = ~n31585 | ~P1_STATE2_REG_1__SCAN_IN;
  assign n31586 = ~n44519 | ~n44508;
  assign n31588 = ~n31587 | ~n31586;
  assign P1_U3162 = n31589 & n31588;
  assign n31590 = ~n44517;
  assign n31592 = ~n31590 | ~P1_STATE2_REG_3__SCAN_IN;
  assign n31591 = ~n44508;
  assign n43049 = ~n31591 | ~P1_STATE2_REG_0__SCAN_IN;
  assign P1_U3466 = ~n31592 | ~n43049;
  assign n31610 = ~n42204 | ~n41789;
  assign n31593 = ~n31610;
  assign n31594 = ~n31598 | ~n31593;
  assign n31675 = ~n31595 & ~n39681;
  assign n31600 = ~n31596;
  assign n31597 = n31610 & P2_EBX_REG_31__SCAN_IN;
  assign n31599 = ~n31598 | ~n31597;
  assign n39683 = ~n39520;
  assign n31621 = ~n31600 & ~n39683;
  assign n31603 = ~n31601;
  assign n31602 = ~P2_STATE2_REG_0__SCAN_IN & ~n42181;
  assign n41893 = ~n31603 | ~n31602;
  assign n31604 = ~n42123 | ~n41664;
  assign n31605 = ~n31604 & ~n42196;
  assign n33133 = ~P2_STATE2_REG_0__SCAN_IN | ~n31605;
  assign n31606 = ~n41893 | ~n33133;
  assign n31619 = ~n39656 | ~P2_PHYADDRPOINTER_REG_31__SCAN_IN;
  assign n31676 = ~n41789 | ~n31608;
  assign n31609 = ~n31676;
  assign n31613 = n31677 | n31609;
  assign n31615 = ~P2_EBX_REG_31__SCAN_IN;
  assign n31611 = n31610 & n31615;
  assign n31612 = ~n40444 | ~n31611;
  assign n31614 = ~n31613 | ~n31612;
  assign n31617 = ~n39495 & ~n31615;
  assign n31616 = ~n39516 & ~n42055;
  assign n31618 = ~n31617 & ~n31616;
  assign n31620 = ~n31619 | ~n31618;
  assign n31673 = ~n31621 & ~n31620;
  assign n31624 = ~n31622 | ~n42214;
  assign n31623 = ~P2_STATE2_REG_0__SCAN_IN | ~P2_INSTADDRPOINTER_REG_31__SCAN_IN;
  assign n42095 = ~n31624 | ~n31623;
  assign n32201 = n31626 ^ n31625;
  assign n32233 = n31628 ^ n31627;
  assign n32263 = n31630 ^ n31629;
  assign n32294 = n31632 ^ n31631;
  assign n39231 = n31634 ^ n31633;
  assign n39272 = n31636 ^ n31635;
  assign n39324 = n31638 ^ n31637;
  assign n39367 = n31640 ^ n31639;
  assign n39396 = n31642 ^ n31641;
  assign n39453 = n31644 ^ n31643;
  assign n39485 = n31646 ^ n31645;
  assign n39531 = n31648 ^ n31647;
  assign n39565 = n31650 ^ n31649;
  assign n39613 = n31651 ^ n31652;
  assign n31654 = ~n42214 | ~P2_PHYADDRPOINTER_REG_0__SCAN_IN;
  assign n31653 = ~P2_STATE2_REG_0__SCAN_IN | ~P2_INSTADDRPOINTER_REG_0__SCAN_IN;
  assign n39675 = ~n31654 | ~n31653;
  assign n31656 = ~n42214 | ~n40329;
  assign n31655 = ~P2_STATE2_REG_0__SCAN_IN | ~P2_INSTADDRPOINTER_REG_1__SCAN_IN;
  assign n39652 = ~n31656 | ~n31655;
  assign n39644 = ~n39675 & ~n39652;
  assign n39612 = ~n39644 | ~n40303;
  assign n39598 = ~n39613 & ~n39612;
  assign n40293 = ~P2_PHYADDRPOINTER_REG_4__SCAN_IN ^ n31657;
  assign n39564 = ~n39598 | ~n40293;
  assign n39549 = ~n39565 & ~n39564;
  assign n39550 = ~P2_PHYADDRPOINTER_REG_6__SCAN_IN ^ n31658;
  assign n39530 = ~n39549 | ~n39550;
  assign n39510 = ~n39531 & ~n39530;
  assign n39511 = ~P2_PHYADDRPOINTER_REG_8__SCAN_IN ^ n31659;
  assign n39484 = ~n39510 | ~n39511;
  assign n39462 = ~n39485 & ~n39484;
  assign n39461 = ~P2_PHYADDRPOINTER_REG_10__SCAN_IN ^ n31660;
  assign n39444 = ~n39462 | ~n39461;
  assign n39419 = ~P2_PHYADDRPOINTER_REG_12__SCAN_IN ^ n31661;
  assign n39394 = ~n39443 | ~n39419;
  assign n39379 = ~P2_PHYADDRPOINTER_REG_14__SCAN_IN ^ n31662;
  assign n39360 = ~n39380 | ~n39379;
  assign n39333 = ~n39367 & ~n39360;
  assign n39336 = ~P2_PHYADDRPOINTER_REG_16__SCAN_IN ^ n31663;
  assign n39317 = ~n39333 | ~n39336;
  assign n39297 = ~P2_PHYADDRPOINTER_REG_18__SCAN_IN ^ n31664;
  assign n39271 = ~n39291 | ~n39297;
  assign n39259 = ~n39272 & ~n39271;
  assign n39258 = ~P2_PHYADDRPOINTER_REG_20__SCAN_IN ^ n31665;
  assign n39261 = ~n39259 | ~n39258;
  assign n39215 = ~n39231 & ~n39261;
  assign n39217 = ~P2_PHYADDRPOINTER_REG_22__SCAN_IN ^ n31666;
  assign n31845 = ~n39215 | ~n39217;
  assign n31824 = ~n32294 & ~n31845;
  assign n32280 = ~P2_PHYADDRPOINTER_REG_24__SCAN_IN ^ n31667;
  assign n31798 = ~n31824 | ~n32280;
  assign n31777 = ~n32263 & ~n31798;
  assign n32248 = ~P2_PHYADDRPOINTER_REG_26__SCAN_IN ^ n31668;
  assign n31754 = ~n31777 | ~n32248;
  assign n32213 = ~P2_PHYADDRPOINTER_REG_28__SCAN_IN ^ n31669;
  assign n31713 = ~n31736 | ~n32213;
  assign n32187 = ~P2_PHYADDRPOINTER_REG_30__SCAN_IN ^ n31670;
  assign n31671 = ~n31689 | ~n32187;
  assign n31672 = n39653 | n31671;
  assign n31674 = ~n31673 | ~n31672;
  assign n31679 = ~n31675 & ~n31674;
  assign n33135 = n31677 | n31676;
  assign n31678 = ~n39820 | ~n39686;
  assign P2_U2824 = ~n31679 | ~n31678;
  assign n31695 = ~n31680 & ~n39681;
  assign n31688 = ~n31681 & ~n39683;
  assign n31686 = ~P2_PHYADDRPOINTER_REG_30__SCAN_IN | ~n39656;
  assign n31684 = ~n39495 & ~n31682;
  assign n31683 = ~n39516 & ~n42056;
  assign n31685 = ~n31684 & ~n31683;
  assign n31687 = ~n31686 | ~n31685;
  assign n31693 = ~n31688 & ~n31687;
  assign n42097 = ~n42095;
  assign n31690 = ~n42097 & ~n31689;
  assign n31691 = ~n32187 ^ n31690;
  assign n31692 = ~n39647 | ~n31691;
  assign n31694 = ~n31693 | ~n31692;
  assign n31698 = ~n31695 & ~n31694;
  assign n32625 = n31696 ^ n31700;
  assign n31697 = ~n32625 | ~n39686;
  assign P2_U2825 = ~n31698 | ~n31697;
  assign n32633 = n31699 ^ n22869;
  assign n31721 = ~n32633 | ~n39639;
  assign n31704 = ~n31700;
  assign n31703 = ~n31727 | ~n31702;
  assign n31719 = ~n32634 & ~n39628;
  assign n31712 = ~n31705 & ~n39683;
  assign n31710 = ~P2_PHYADDRPOINTER_REG_29__SCAN_IN | ~n39672;
  assign n31706 = ~P2_EBX_REG_29__SCAN_IN;
  assign n31708 = ~n39495 & ~n31706;
  assign n31707 = ~n39516 & ~n42050;
  assign n31709 = ~n31708 & ~n31707;
  assign n31711 = ~n31710 | ~n31709;
  assign n31717 = ~n31712 & ~n31711;
  assign n31714 = ~n42095 | ~n31713;
  assign n31715 = ~n31714 ^ n32201;
  assign n31716 = ~n31715 | ~n39647;
  assign n31718 = ~n31717 | ~n31716;
  assign n31720 = ~n31719 & ~n31718;
  assign P2_U2826 = ~n31721 | ~n31720;
  assign n32650 = n31723 ^ n31722;
  assign n31744 = ~n32650 | ~n39639;
  assign n31726 = n31725 | n31724;
  assign n32651 = ~n31727 | ~n31726;
  assign n31742 = ~n32651 & ~n39628;
  assign n31735 = ~n31728 & ~n39683;
  assign n31733 = ~P2_PHYADDRPOINTER_REG_28__SCAN_IN | ~n39672;
  assign n31729 = ~P2_EBX_REG_28__SCAN_IN;
  assign n31731 = ~n39495 & ~n31729;
  assign n31730 = ~n39516 & ~n42045;
  assign n31732 = ~n31731 & ~n31730;
  assign n31734 = ~n31733 | ~n31732;
  assign n31740 = ~n31735 & ~n31734;
  assign n31737 = ~n42097 & ~n31736;
  assign n31738 = ~n32213 ^ n31737;
  assign n31739 = ~n39647 | ~n31738;
  assign n31741 = ~n31740 | ~n31739;
  assign n31743 = ~n31742 & ~n31741;
  assign P2_U2827 = ~n31744 | ~n31743;
  assign n31760 = ~n31745 & ~n39681;
  assign n31753 = ~n31746 & ~n39683;
  assign n31751 = ~P2_PHYADDRPOINTER_REG_27__SCAN_IN | ~n39656;
  assign n31747 = ~P2_EBX_REG_27__SCAN_IN;
  assign n31749 = ~n39495 & ~n31747;
  assign n31748 = ~n39516 & ~n42040;
  assign n31750 = ~n31749 & ~n31748;
  assign n31752 = ~n31751 | ~n31750;
  assign n31758 = ~n31753 & ~n31752;
  assign n31755 = ~n42095 | ~n31754;
  assign n31756 = ~n31755 ^ n32233;
  assign n31757 = ~n31756 | ~n39647;
  assign n31759 = ~n31758 | ~n31757;
  assign n31762 = ~n31760 & ~n31759;
  assign n31761 = ~n32015 | ~n39686;
  assign P2_U2828 = ~n31762 | ~n31761;
  assign n31767 = ~n31763;
  assign n31766 = ~n31765 & ~n31764;
  assign n32669 = ~n31767 & ~n31766;
  assign n32031 = ~n32669;
  assign n31783 = ~n32031 & ~n39628;
  assign n31769 = ~n31768;
  assign n31776 = ~n31769 & ~n39683;
  assign n31774 = ~P2_PHYADDRPOINTER_REG_26__SCAN_IN | ~n39656;
  assign n31770 = ~P2_EBX_REG_26__SCAN_IN;
  assign n31772 = ~n39495 & ~n31770;
  assign n31771 = ~n39516 & ~n42035;
  assign n31773 = ~n31772 & ~n31771;
  assign n31775 = ~n31774 | ~n31773;
  assign n31781 = ~n31776 & ~n31775;
  assign n31778 = ~n42097 & ~n31777;
  assign n31779 = ~n32248 ^ n31778;
  assign n31780 = ~n39647 | ~n31779;
  assign n31782 = ~n31781 | ~n31780;
  assign n31787 = ~n31783 & ~n31782;
  assign n32668 = n31785 ^ n31784;
  assign n31786 = ~n32668 | ~n39639;
  assign P2_U2829 = ~n31787 | ~n31786;
  assign n32262 = n31789 ^ n31788;
  assign n32690 = ~n32262;
  assign n31804 = ~n32690 & ~n39681;
  assign n31797 = ~n31790 & ~n39683;
  assign n31795 = ~P2_PHYADDRPOINTER_REG_25__SCAN_IN | ~n39656;
  assign n31791 = ~P2_EBX_REG_25__SCAN_IN;
  assign n31793 = ~n39495 & ~n31791;
  assign n31792 = ~n39516 & ~n42030;
  assign n31794 = ~n31793 & ~n31792;
  assign n31796 = ~n31795 | ~n31794;
  assign n31802 = ~n31797 & ~n31796;
  assign n31799 = ~n42095 | ~n31798;
  assign n31800 = ~n31799 ^ n32263;
  assign n31801 = ~n31800 | ~n39647;
  assign n31803 = ~n31802 | ~n31801;
  assign n31808 = ~n31804 & ~n31803;
  assign n32699 = n31806 ^ n31813;
  assign n31807 = ~n32699 | ~n39686;
  assign P2_U2830 = ~n31808 | ~n31807;
  assign n32709 = ~n31810 ^ n31809;
  assign n31830 = ~n32709 & ~n39681;
  assign n31812 = ~n22938 | ~n31811;
  assign n32710 = ~n31813 | ~n31812;
  assign n31823 = ~n32710 & ~n39628;
  assign n31821 = ~n31814 & ~n39683;
  assign n31819 = ~P2_PHYADDRPOINTER_REG_24__SCAN_IN | ~n39656;
  assign n31815 = ~P2_EBX_REG_24__SCAN_IN;
  assign n31817 = ~n39495 & ~n31815;
  assign n31816 = ~n39516 & ~n42025;
  assign n31818 = ~n31817 & ~n31816;
  assign n31820 = ~n31819 | ~n31818;
  assign n31822 = n31821 | n31820;
  assign n31828 = ~n31823 & ~n31822;
  assign n31825 = ~n42097 & ~n31824;
  assign n31826 = ~n32280 ^ n31825;
  assign n31827 = ~n39647 | ~n31826;
  assign n31829 = ~n31828 | ~n31827;
  assign P2_U2831 = n31830 | n31829;
  assign n32728 = n31832 ^ n31831;
  assign n31842 = ~n32728 | ~n39639;
  assign n31840 = ~n31833 & ~n39683;
  assign n31838 = ~P2_PHYADDRPOINTER_REG_23__SCAN_IN | ~n39656;
  assign n31834 = ~P2_EBX_REG_23__SCAN_IN;
  assign n31836 = ~n39495 & ~n31834;
  assign n31835 = ~n39516 & ~n42018;
  assign n31837 = ~n31836 & ~n31835;
  assign n31839 = ~n31838 | ~n31837;
  assign n31841 = ~n31840 & ~n31839;
  assign n31851 = ~n31842 | ~n31841;
  assign n32743 = n31844 ^ n31843;
  assign n31849 = ~n32743 | ~n39686;
  assign n31846 = ~n42095 | ~n31845;
  assign n31847 = ~n31846 ^ n32294;
  assign n31848 = ~n31847 | ~n39647;
  assign n31850 = ~n31849 | ~n31848;
  assign P2_U2832 = n31851 | n31850;
  assign n31853 = ~n29864 | ~n31948;
  assign n31852 = ~n39817 | ~P2_EBX_REG_31__SCAN_IN;
  assign P2_U2856 = ~n31853 | ~n31852;
  assign n31856 = ~n32633 & ~n39817;
  assign n31855 = ~n31948 & ~P2_EBX_REG_29__SCAN_IN;
  assign n31857 = n31856 | n31855;
  assign P2_U2858 = ~n31858 | ~n31857;
  assign n32000 = n31860 ^ n31859;
  assign n31864 = ~n32000 | ~n39782;
  assign n31862 = ~n32650 & ~n39817;
  assign n31861 = ~n31948 & ~P2_EBX_REG_28__SCAN_IN;
  assign n31863 = n31862 | n31861;
  assign P2_U2859 = ~n31864 | ~n31863;
  assign n31869 = ~n32014 | ~n39782;
  assign n31867 = ~n32232 & ~n39817;
  assign n31866 = ~n31948 & ~P2_EBX_REG_27__SCAN_IN;
  assign n31868 = n31867 | n31866;
  assign P2_U2860 = ~n31869 | ~n31868;
  assign n31874 = ~n31870;
  assign n31873 = ~n31872 & ~n31871;
  assign n32030 = ~n31874 & ~n31873;
  assign n31878 = ~n32030 | ~n39782;
  assign n31876 = ~n32668 & ~n39817;
  assign n31875 = ~n31948 & ~P2_EBX_REG_26__SCAN_IN;
  assign n31877 = n31876 | n31875;
  assign P2_U2861 = ~n31878 | ~n31877;
  assign n31880 = ~n32262 & ~n39817;
  assign n31879 = ~n31948 & ~P2_EBX_REG_25__SCAN_IN;
  assign n31883 = n31880 | n31879;
  assign n31882 = ~n32057 | ~n39782;
  assign P2_U2862 = ~n31883 | ~n31882;
  assign n31885 = ~n32709 | ~n31948;
  assign n31884 = n31948 | P2_EBX_REG_24__SCAN_IN;
  assign n31893 = ~n31885 | ~n31884;
  assign n31891 = ~n31887 | ~n31886;
  assign n31890 = ~n31889 ^ n31888;
  assign n32071 = ~n31891 ^ n31890;
  assign n31892 = ~n32071 | ~n39782;
  assign P2_U2863 = ~n31893 | ~n31892;
  assign n31895 = ~n32728 & ~n39817;
  assign n31894 = ~n31948 & ~P2_EBX_REG_23__SCAN_IN;
  assign n31899 = n31895 | n31894;
  assign n32074 = n31897 ^ n31896;
  assign n31898 = ~n32074 | ~n39782;
  assign P2_U2864 = ~n31899 | ~n31898;
  assign n39214 = n31901 ^ n31900;
  assign n31903 = ~n39214 & ~n39817;
  assign n31902 = ~n31948 & ~P2_EBX_REG_22__SCAN_IN;
  assign n31911 = n31903 | n31902;
  assign n39699 = ~n39709 & ~n39708;
  assign n39701 = ~n39699 | ~n39698;
  assign n31941 = ~n39701 & ~n31951;
  assign n31940 = ~n31904;
  assign n31939 = ~n31941 | ~n31940;
  assign n31923 = ~n31939 & ~n31932;
  assign n31922 = ~n31905;
  assign n31921 = ~n31923 | ~n31922;
  assign n31907 = ~n31921 & ~n31914;
  assign n31909 = ~n31907 & ~n31906;
  assign n32088 = ~n31909 & ~n31908;
  assign n31910 = ~n32088 | ~n39782;
  assign P2_U2865 = ~n31911 | ~n31910;
  assign n31913 = ~n39230 & ~n39817;
  assign n31912 = ~n31948 & ~P2_EBX_REG_21__SCAN_IN;
  assign n31916 = n31913 | n31912;
  assign n32117 = n31914 ^ n31921;
  assign n31915 = ~n32117 | ~n39782;
  assign P2_U2866 = ~n31916 | ~n31915;
  assign n31920 = ~n31917 | ~n31948;
  assign n31918 = ~P2_EBX_REG_20__SCAN_IN;
  assign n31919 = ~n39817 | ~n31918;
  assign n31927 = ~n31920 | ~n31919;
  assign n31925 = ~n31921;
  assign n31924 = ~n31923 & ~n31922;
  assign n32120 = ~n31925 & ~n31924;
  assign n31926 = ~n32120 | ~n39782;
  assign P2_U2867 = ~n31927 | ~n31926;
  assign n39275 = n31929 ^ n31928;
  assign n31931 = ~n39275 & ~n39817;
  assign n31930 = ~n31948 & ~P2_EBX_REG_19__SCAN_IN;
  assign n31934 = n31931 | n31930;
  assign n32135 = n31932 ^ n31939;
  assign n31933 = ~n32135 | ~n39782;
  assign P2_U2868 = ~n31934 | ~n31933;
  assign n39308 = n31936 ^ n31935;
  assign n31938 = ~n39308 & ~n39817;
  assign n31937 = ~n31948 & ~P2_EBX_REG_18__SCAN_IN;
  assign n31945 = n31938 | n31937;
  assign n31943 = ~n31939;
  assign n31942 = ~n31941 & ~n31940;
  assign n32150 = ~n31943 & ~n31942;
  assign n31944 = ~n32150 | ~n39782;
  assign P2_U2869 = ~n31945 | ~n31944;
  assign n39325 = n31947 ^ n31946;
  assign n31950 = ~n39325 & ~n39817;
  assign n31949 = ~n31948 & ~P2_EBX_REG_17__SCAN_IN;
  assign n31953 = n31950 | n31949;
  assign n32167 = n31951 ^ n39701;
  assign n31952 = ~n32167 | ~n39782;
  assign P2_U2870 = ~n31953 | ~n31952;
  assign n31957 = ~n31954;
  assign n31956 = ~n31955;
  assign n31959 = ~n31957 | ~n31956;
  assign n31963 = ~n42170 | ~n39782;
  assign n31960 = n39817 & P2_EBX_REG_1__SCAN_IN;
  assign n31962 = ~n31961 & ~n31960;
  assign P2_U2886 = ~n31963 | ~n31962;
  assign n31965 = ~n33239 & ~n33237;
  assign n31967 = ~n31965 | ~n33240;
  assign n33231 = ~n33228;
  assign n31970 = ~n39849;
  assign n31987 = ~n31971 | ~n39964;
  assign n31972 = ~n39945;
  assign n31985 = n32625 & n31972;
  assign n39828 = ~n31981 & ~n40435;
  assign n31973 = ~BUF2_REG_30__SCAN_IN;
  assign n31980 = ~n32171 & ~n31973;
  assign n39835 = ~n39970 & ~n31974;
  assign n31976 = ~BUF1_REG_14__SCAN_IN | ~n40435;
  assign n31975 = ~n40437 | ~BUF2_REG_14__SCAN_IN;
  assign n40195 = ~n31976 | ~n31975;
  assign n31978 = ~n39835 | ~n40195;
  assign n31977 = ~n39970 | ~P2_EAX_REG_30__SCAN_IN;
  assign n31979 = ~n31978 | ~n31977;
  assign n31983 = ~n31980 & ~n31979;
  assign n39839 = ~n31981 & ~n40437;
  assign n31982 = ~n39839 | ~BUF1_REG_30__SCAN_IN;
  assign n31984 = ~n31983 | ~n31982;
  assign n31986 = ~n31985 & ~n31984;
  assign P2_U2889 = ~n31987 | ~n31986;
  assign n31997 = ~n32634 & ~n39945;
  assign n31993 = ~n32171 & ~n40515;
  assign n31989 = ~n40435 | ~BUF1_REG_13__SCAN_IN;
  assign n31988 = ~n40437 | ~BUF2_REG_13__SCAN_IN;
  assign n40189 = ~n31989 | ~n31988;
  assign n31991 = ~n39835 | ~n40189;
  assign n31990 = ~n39970 | ~P2_EAX_REG_29__SCAN_IN;
  assign n31992 = ~n31991 | ~n31990;
  assign n31995 = ~n31993 & ~n31992;
  assign n31994 = ~n39839 | ~BUF1_REG_29__SCAN_IN;
  assign n31996 = ~n31995 | ~n31994;
  assign n31998 = ~n31997 & ~n31996;
  assign P2_U2890 = ~n31999 | ~n31998;
  assign n32013 = ~n32000 | ~n39964;
  assign n32011 = ~n32651 & ~n39945;
  assign n32001 = ~BUF2_REG_28__SCAN_IN;
  assign n32007 = ~n32171 & ~n32001;
  assign n32003 = ~n40435 | ~BUF1_REG_12__SCAN_IN;
  assign n32002 = ~n40437 | ~BUF2_REG_12__SCAN_IN;
  assign n40183 = ~n32003 | ~n32002;
  assign n32005 = ~n39835 | ~n40183;
  assign n32004 = ~n39970 | ~P2_EAX_REG_28__SCAN_IN;
  assign n32006 = ~n32005 | ~n32004;
  assign n32009 = ~n32007 & ~n32006;
  assign n32008 = ~n39839 | ~BUF1_REG_28__SCAN_IN;
  assign n32010 = ~n32009 | ~n32008;
  assign n32012 = ~n32011 & ~n32010;
  assign P2_U2891 = ~n32013 | ~n32012;
  assign n32029 = ~n32014 | ~n39964;
  assign n32016 = ~n32015;
  assign n32027 = ~n32016 & ~n39945;
  assign n32017 = ~BUF2_REG_27__SCAN_IN;
  assign n32023 = ~n32171 & ~n32017;
  assign n32019 = ~n40435 | ~BUF1_REG_11__SCAN_IN;
  assign n32018 = ~n40437 | ~BUF2_REG_11__SCAN_IN;
  assign n40177 = ~n32019 | ~n32018;
  assign n32021 = ~n39835 | ~n40177;
  assign n32020 = ~n39970 | ~P2_EAX_REG_27__SCAN_IN;
  assign n32022 = ~n32021 | ~n32020;
  assign n32025 = ~n32023 & ~n32022;
  assign n32024 = ~n39839 | ~BUF1_REG_27__SCAN_IN;
  assign n32026 = ~n32025 | ~n32024;
  assign n32028 = ~n32027 & ~n32026;
  assign P2_U2892 = ~n32029 | ~n32028;
  assign n32044 = ~n32030 | ~n39964;
  assign n32042 = ~n32031 & ~n39945;
  assign n32032 = ~BUF2_REG_26__SCAN_IN;
  assign n32038 = ~n32171 & ~n32032;
  assign n32034 = ~n40435 | ~BUF1_REG_10__SCAN_IN;
  assign n32033 = ~n40437 | ~BUF2_REG_10__SCAN_IN;
  assign n40171 = ~n32034 | ~n32033;
  assign n32036 = ~n39835 | ~n40171;
  assign n32035 = ~n39970 | ~P2_EAX_REG_26__SCAN_IN;
  assign n32037 = ~n32036 | ~n32035;
  assign n32040 = ~n32038 & ~n32037;
  assign n32039 = ~n39839 | ~BUF1_REG_26__SCAN_IN;
  assign n32041 = ~n32040 | ~n32039;
  assign n32043 = ~n32042 & ~n32041;
  assign P2_U2893 = ~n32044 | ~n32043;
  assign n32045 = ~n32699;
  assign n32056 = ~n32045 & ~n39945;
  assign n32046 = ~BUF2_REG_25__SCAN_IN;
  assign n32052 = ~n32171 & ~n32046;
  assign n32048 = ~n40435 | ~BUF1_REG_9__SCAN_IN;
  assign n32047 = ~n40437 | ~BUF2_REG_9__SCAN_IN;
  assign n40165 = ~n32048 | ~n32047;
  assign n32050 = ~n39835 | ~n40165;
  assign n32049 = ~n39970 | ~P2_EAX_REG_25__SCAN_IN;
  assign n32051 = ~n32050 | ~n32049;
  assign n32054 = ~n32052 & ~n32051;
  assign n32053 = ~n39839 | ~BUF1_REG_25__SCAN_IN;
  assign n32055 = ~n32054 | ~n32053;
  assign n32059 = ~n32056 & ~n32055;
  assign n32058 = ~n32057 | ~n39964;
  assign P2_U2894 = ~n32059 | ~n32058;
  assign n32070 = ~n32710 & ~n39945;
  assign n32060 = ~BUF2_REG_24__SCAN_IN;
  assign n32066 = ~n32171 & ~n32060;
  assign n32062 = ~n40435 | ~BUF1_REG_8__SCAN_IN;
  assign n32061 = ~n40437 | ~BUF2_REG_8__SCAN_IN;
  assign n40159 = ~n32062 | ~n32061;
  assign n32064 = ~n39835 | ~n40159;
  assign n32063 = ~n39970 | ~P2_EAX_REG_24__SCAN_IN;
  assign n32065 = ~n32064 | ~n32063;
  assign n32068 = ~n32066 & ~n32065;
  assign n32067 = ~n39839 | ~BUF1_REG_24__SCAN_IN;
  assign n32069 = ~n32068 | ~n32067;
  assign n32073 = ~n32070 & ~n32069;
  assign n32072 = ~n32071 | ~n39964;
  assign P2_U2895 = ~n32073 | ~n32072;
  assign n32087 = ~n32743 | ~n31972;
  assign n32085 = n32074 & n39964;
  assign n32075 = ~BUF2_REG_23__SCAN_IN;
  assign n32081 = ~n32171 & ~n32075;
  assign n32077 = ~n40435 | ~BUF1_REG_7__SCAN_IN;
  assign n32076 = ~n40437 | ~BUF2_REG_7__SCAN_IN;
  assign n40565 = ~n32077 | ~n32076;
  assign n32079 = ~n39835 | ~n40565;
  assign n32078 = ~n39970 | ~P2_EAX_REG_23__SCAN_IN;
  assign n32080 = ~n32079 | ~n32078;
  assign n32083 = ~n32081 & ~n32080;
  assign n32082 = ~n39839 | ~BUF1_REG_23__SCAN_IN;
  assign n32084 = ~n32083 | ~n32082;
  assign n32086 = ~n32085 & ~n32084;
  assign P2_U2896 = ~n32087 | ~n32086;
  assign n32104 = ~n32088 | ~n39964;
  assign n32091 = ~n32090 & ~n32089;
  assign n39224 = n31843 | n32091;
  assign n32102 = ~n39224 & ~n39945;
  assign n32092 = ~BUF2_REG_22__SCAN_IN;
  assign n32098 = ~n32171 & ~n32092;
  assign n32094 = ~n40435 | ~BUF1_REG_6__SCAN_IN;
  assign n32093 = ~n40437 | ~BUF2_REG_6__SCAN_IN;
  assign n40543 = ~n32094 | ~n32093;
  assign n32096 = ~n39835 | ~n40543;
  assign n32095 = ~n39970 | ~P2_EAX_REG_22__SCAN_IN;
  assign n32097 = ~n32096 | ~n32095;
  assign n32100 = ~n32098 & ~n32097;
  assign n32099 = ~n39839 | ~BUF1_REG_22__SCAN_IN;
  assign n32101 = ~n32100 | ~n32099;
  assign n32103 = ~n32102 & ~n32101;
  assign P2_U2897 = ~n32104 | ~n32103;
  assign n39242 = ~n32105;
  assign n32116 = ~n39242 & ~n39945;
  assign n32106 = ~BUF2_REG_21__SCAN_IN;
  assign n32112 = ~n32171 & ~n32106;
  assign n32108 = ~n40435 | ~BUF1_REG_5__SCAN_IN;
  assign n32107 = ~n40437 | ~BUF2_REG_5__SCAN_IN;
  assign n40528 = ~n32108 | ~n32107;
  assign n32110 = ~n39835 | ~n40528;
  assign n32109 = ~n39970 | ~P2_EAX_REG_21__SCAN_IN;
  assign n32111 = ~n32110 | ~n32109;
  assign n32114 = ~n32112 & ~n32111;
  assign n32113 = ~n39839 | ~BUF1_REG_21__SCAN_IN;
  assign n32115 = ~n32114 | ~n32113;
  assign n32119 = ~n32116 & ~n32115;
  assign n32118 = ~n32117 | ~n39964;
  assign P2_U2898 = ~n32119 | ~n32118;
  assign n32134 = ~n32120 | ~n39964;
  assign n32121 = ~n39248;
  assign n32132 = ~n32121 & ~n39945;
  assign n32122 = ~BUF2_REG_20__SCAN_IN;
  assign n32128 = ~n32171 & ~n32122;
  assign n32124 = ~n40435 | ~BUF1_REG_4__SCAN_IN;
  assign n32123 = ~n40437 | ~BUF2_REG_4__SCAN_IN;
  assign n40510 = ~n32124 | ~n32123;
  assign n32126 = ~n39835 | ~n40510;
  assign n32125 = ~n39970 | ~P2_EAX_REG_20__SCAN_IN;
  assign n32127 = ~n32126 | ~n32125;
  assign n32130 = ~n32128 & ~n32127;
  assign n32129 = ~n39839 | ~BUF1_REG_20__SCAN_IN;
  assign n32131 = ~n32130 | ~n32129;
  assign n32133 = ~n32132 & ~n32131;
  assign P2_U2899 = ~n32134 | ~n32133;
  assign n32149 = ~n32135 | ~n39964;
  assign n39270 = ~n32153 ^ n32136;
  assign n32147 = ~n39270 & ~n39945;
  assign n32137 = ~BUF2_REG_19__SCAN_IN;
  assign n32143 = ~n32171 & ~n32137;
  assign n32139 = ~n40435 | ~BUF1_REG_3__SCAN_IN;
  assign n32138 = ~n40437 | ~BUF2_REG_3__SCAN_IN;
  assign n40495 = ~n32139 | ~n32138;
  assign n32141 = ~n39835 | ~n40495;
  assign n32140 = ~n39970 | ~P2_EAX_REG_19__SCAN_IN;
  assign n32142 = ~n32141 | ~n32140;
  assign n32145 = ~n32143 & ~n32142;
  assign n32144 = ~n39839 | ~BUF1_REG_19__SCAN_IN;
  assign n32146 = ~n32145 | ~n32144;
  assign n32148 = ~n32147 & ~n32146;
  assign P2_U2900 = ~n32149 | ~n32148;
  assign n32166 = ~n32150 | ~n39964;
  assign n32152 = ~n22945 & ~n32151;
  assign n39290 = n32153 | n32152;
  assign n32164 = ~n39290 & ~n39945;
  assign n32154 = ~BUF2_REG_18__SCAN_IN;
  assign n32160 = ~n32171 & ~n32154;
  assign n32156 = ~n40435 | ~BUF1_REG_2__SCAN_IN;
  assign n32155 = ~n40437 | ~BUF2_REG_2__SCAN_IN;
  assign n40480 = ~n32156 | ~n32155;
  assign n32158 = ~n39835 | ~n40480;
  assign n32157 = ~n39970 | ~P2_EAX_REG_18__SCAN_IN;
  assign n32159 = ~n32158 | ~n32157;
  assign n32162 = ~n32160 & ~n32159;
  assign n32161 = ~n39839 | ~BUF1_REG_18__SCAN_IN;
  assign n32163 = ~n32162 | ~n32161;
  assign n32165 = ~n32164 & ~n32163;
  assign P2_U2901 = ~n32166 | ~n32165;
  assign n32183 = ~n32167 | ~n39964;
  assign n39328 = ~n32169 ^ n32168;
  assign n32181 = ~n39328 & ~n39945;
  assign n32170 = ~BUF2_REG_17__SCAN_IN;
  assign n32177 = ~n32171 & ~n32170;
  assign n32173 = ~n40435 | ~BUF1_REG_1__SCAN_IN;
  assign n32172 = ~n40437 | ~BUF2_REG_1__SCAN_IN;
  assign n40465 = ~n32173 | ~n32172;
  assign n32175 = ~n39835 | ~n40465;
  assign n32174 = ~n39970 | ~P2_EAX_REG_17__SCAN_IN;
  assign n32176 = ~n32175 | ~n32174;
  assign n32179 = ~n32177 & ~n32176;
  assign n32178 = ~n39839 | ~BUF1_REG_17__SCAN_IN;
  assign n32180 = ~n32179 | ~n32178;
  assign n32182 = ~n32181 & ~n32180;
  assign P2_U2902 = ~n32183 | ~n32182;
  assign n32196 = ~n32613 | ~n40348;
  assign n32185 = ~n32184 ^ n32617;
  assign n32614 = ~n32186 ^ n32185;
  assign n32194 = ~n32614 & ~n40342;
  assign n32192 = ~n32615 | ~n40324;
  assign n32190 = ~n32187 & ~n40304;
  assign n32619 = ~n40325 | ~P2_REIP_REG_30__SCAN_IN;
  assign n32188 = ~n40337 | ~P2_PHYADDRPOINTER_REG_30__SCAN_IN;
  assign n32189 = ~n32619 | ~n32188;
  assign n32191 = ~n32190 & ~n32189;
  assign n32193 = ~n32192 | ~n32191;
  assign n32195 = ~n32194 & ~n32193;
  assign P2_U2984 = ~n32196 | ~n32195;
  assign n32210 = ~n32632 & ~n40342;
  assign n32208 = ~n32633 | ~n40324;
  assign n32202 = ~n32201;
  assign n32206 = ~n32202 & ~n40304;
  assign n32641 = ~n40294 & ~n42050;
  assign n32204 = ~n32641;
  assign n32203 = ~n40337 | ~P2_PHYADDRPOINTER_REG_29__SCAN_IN;
  assign n32205 = ~n32204 | ~n32203;
  assign n32207 = ~n32206 & ~n32205;
  assign n32209 = ~n32208 | ~n32207;
  assign n32219 = ~n32650 | ~n40324;
  assign n32217 = ~n32213 & ~n40304;
  assign n32656 = ~n40294 & ~n42045;
  assign n32215 = ~n32656;
  assign n32214 = ~n40337 | ~P2_PHYADDRPOINTER_REG_28__SCAN_IN;
  assign n32216 = ~n32215 | ~n32214;
  assign n32218 = ~n32217 & ~n32216;
  assign n32220 = ~n32219 | ~n32218;
  assign n32229 = ~n32221 & ~n32220;
  assign n32225 = ~n32223 | ~n32222;
  assign n32226 = ~n32225 | ~n32224;
  assign P2_U2986 = ~n32229 | ~n32228;
  assign n32244 = ~n32230 | ~n32597;
  assign n32242 = ~n32231 & ~n40323;
  assign n32240 = ~n32232 | ~n40324;
  assign n32234 = ~n32233;
  assign n32238 = ~n32234 & ~n40304;
  assign n32235 = ~n40337 | ~P2_PHYADDRPOINTER_REG_27__SCAN_IN;
  assign n32237 = ~n32236 | ~n32235;
  assign n32239 = ~n32238 & ~n32237;
  assign n32241 = ~n32240 | ~n32239;
  assign n32243 = ~n32242 & ~n32241;
  assign P2_U2987 = ~n32244 | ~n32243;
  assign n32247 = ~n32246 | ~n32245;
  assign n32253 = ~n32668 | ~n40324;
  assign n32251 = ~n32248 & ~n40304;
  assign n32679 = ~n40325 | ~P2_REIP_REG_26__SCAN_IN;
  assign n32249 = ~n40337 | ~P2_PHYADDRPOINTER_REG_26__SCAN_IN;
  assign n32250 = ~n32679 | ~n32249;
  assign n32252 = ~n32251 & ~n32250;
  assign n32255 = ~n32257;
  assign n32273 = ~n32255 | ~n32254;
  assign n32258 = ~n32272 | ~n23751;
  assign n32260 = ~n32273 | ~n32258;
  assign n32269 = ~n32262 | ~n40324;
  assign n32264 = ~n32263;
  assign n32267 = ~n32264 & ~n40304;
  assign n32695 = ~n40325 | ~P2_REIP_REG_25__SCAN_IN;
  assign n32265 = ~n40337 | ~P2_PHYADDRPOINTER_REG_25__SCAN_IN;
  assign n32266 = ~n32695 | ~n32265;
  assign n32268 = ~n32267 & ~n32266;
  assign n32270 = ~n32269 | ~n32268;
  assign n32276 = ~n32271 & ~n32270;
  assign n32274 = ~n32273 | ~n32272;
  assign n32704 = ~n32274 ^ P2_INSTADDRPOINTER_REG_25__SCAN_IN;
  assign n32275 = ~n32704 | ~n32597;
  assign P2_U2989 = ~n32276 | ~n32275;
  assign n32289 = ~n32707 | ~n40348;
  assign n32278 = n23043 & n32277;
  assign n32708 = ~n32279 ^ n32278;
  assign n32287 = n32708 | n40342;
  assign n32285 = n32709 | n40344;
  assign n32283 = ~n32280 & ~n40304;
  assign n32714 = ~n40325 | ~P2_REIP_REG_24__SCAN_IN;
  assign n32281 = ~n40337 | ~P2_PHYADDRPOINTER_REG_24__SCAN_IN;
  assign n32282 = ~n32714 | ~n32281;
  assign n32284 = ~n32283 & ~n32282;
  assign n32286 = n32285 & n32284;
  assign n32288 = n32287 & n32286;
  assign P2_U2990 = ~n32289 | ~n32288;
  assign n32290 = ~n32305 & ~P2_INSTADDRPOINTER_REG_23__SCAN_IN;
  assign n32304 = ~n32726 | ~n40348;
  assign n32293 = ~n32292 | ~n32291;
  assign n32302 = ~n32727 & ~n40342;
  assign n32300 = ~n32728 | ~n40324;
  assign n32295 = ~n32294;
  assign n32298 = ~n32295 & ~n40304;
  assign n32737 = ~n40325 | ~P2_REIP_REG_23__SCAN_IN;
  assign n32296 = ~n40337 | ~P2_PHYADDRPOINTER_REG_23__SCAN_IN;
  assign n32297 = ~n32737 | ~n32296;
  assign n32299 = ~n32298 & ~n32297;
  assign n32301 = ~n32300 | ~n32299;
  assign n32303 = ~n32302 & ~n32301;
  assign P2_U2991 = ~n32304 | ~n32303;
  assign n32320 = ~n32750 | ~n40348;
  assign n32308 = ~n32307 | ~n32306;
  assign n32751 = ~n32309 ^ n32308;
  assign n32318 = ~n32751 & ~n40342;
  assign n32316 = ~n39214 | ~n40324;
  assign n32314 = ~n39217 & ~n40304;
  assign n32754 = ~n40294 & ~n32310;
  assign n32312 = ~n32754;
  assign n32311 = ~n40337 | ~P2_PHYADDRPOINTER_REG_22__SCAN_IN;
  assign n32313 = ~n32312 | ~n32311;
  assign n32315 = ~n32314 & ~n32313;
  assign n32317 = ~n32316 | ~n32315;
  assign n32319 = ~n32318 & ~n32317;
  assign P2_U2992 = ~n32320 | ~n32319;
  assign n32330 = ~n32321 & ~n40323;
  assign n32328 = ~n39230 | ~n40324;
  assign n32322 = ~n39231;
  assign n32326 = ~n32322 & ~n40304;
  assign n32323 = ~n40337 | ~P2_PHYADDRPOINTER_REG_21__SCAN_IN;
  assign n32325 = ~n32324 | ~n32323;
  assign n32327 = ~n32326 & ~n32325;
  assign n32329 = ~n32328 | ~n32327;
  assign n32331 = ~n32330 & ~n32329;
  assign P2_U2993 = ~n32332 | ~n32331;
  assign n32341 = ~n32333 & ~n40323;
  assign n32339 = ~n39267 | ~n40324;
  assign n32337 = ~n39258 & ~n40304;
  assign n32334 = ~n40337 | ~P2_PHYADDRPOINTER_REG_20__SCAN_IN;
  assign n32336 = ~n32335 | ~n32334;
  assign n32338 = ~n32337 & ~n32336;
  assign n32340 = ~n32339 | ~n32338;
  assign n32342 = ~n32341 & ~n32340;
  assign P2_U2994 = ~n32343 | ~n32342;
  assign n32347 = ~n32359 | ~n32360;
  assign n32354 = ~n39275 | ~n40324;
  assign n32349 = ~n39272;
  assign n32352 = ~n32349 & ~n40304;
  assign n32766 = ~n40325 | ~P2_REIP_REG_19__SCAN_IN;
  assign n32350 = ~n40337 | ~P2_PHYADDRPOINTER_REG_19__SCAN_IN;
  assign n32351 = ~n32766 | ~n32350;
  assign n32353 = ~n32352 & ~n32351;
  assign n32355 = ~n32354 | ~n32353;
  assign n32357 = ~n32356 & ~n32355;
  assign P2_U2995 = ~n32358 | ~n32357;
  assign n32371 = ~n32781 | ~n32597;
  assign n32367 = ~n39308 | ~n40324;
  assign n32365 = ~n39297 & ~n40304;
  assign n32786 = ~n40325 | ~P2_REIP_REG_18__SCAN_IN;
  assign n32363 = ~n40337 | ~P2_PHYADDRPOINTER_REG_18__SCAN_IN;
  assign n32364 = ~n32786 | ~n32363;
  assign n32366 = ~n32365 & ~n32364;
  assign n32368 = ~n32367 | ~n32366;
  assign n32370 = ~n32369 & ~n32368;
  assign P2_U2996 = ~n32371 | ~n32370;
  assign n32375 = ~n32374 | ~n32373;
  assign n32798 = ~n32372 ^ n32375;
  assign n32388 = ~n32798 | ~n32597;
  assign n32378 = ~n32799 & ~P2_INSTADDRPOINTER_REG_17__SCAN_IN;
  assign n32377 = ~n32361 | ~n40348;
  assign n32386 = ~n32378 & ~n32377;
  assign n32384 = ~n39325 | ~n40324;
  assign n32379 = ~n39324;
  assign n32382 = ~n32379 & ~n40304;
  assign n32811 = ~n40325 | ~P2_REIP_REG_17__SCAN_IN;
  assign n32380 = ~n40337 | ~P2_PHYADDRPOINTER_REG_17__SCAN_IN;
  assign n32381 = ~n32811 | ~n32380;
  assign n32383 = ~n32382 & ~n32381;
  assign n32385 = ~n32384 | ~n32383;
  assign n32387 = ~n32386 & ~n32385;
  assign P2_U2997 = ~n32388 | ~n32387;
  assign n32827 = n32389 ^ n32390;
  assign n32400 = ~n32827 | ~n32597;
  assign n39704 = n32391 ^ n22875;
  assign n32396 = ~n39704 | ~n40324;
  assign n32394 = ~n40304 & ~n39336;
  assign n32821 = ~n40325 | ~P2_REIP_REG_16__SCAN_IN;
  assign n32392 = ~n40337 | ~P2_PHYADDRPOINTER_REG_16__SCAN_IN;
  assign n32393 = ~n32821 | ~n32392;
  assign n32395 = ~n32394 & ~n32393;
  assign n32397 = ~n32396 | ~n32395;
  assign n32399 = ~n32398 & ~n32397;
  assign P2_U2998 = ~n32400 | ~n32399;
  assign n32417 = ~n32829 | ~n32597;
  assign n39713 = n32406 ^ n32405;
  assign n32413 = ~n39713 | ~n40324;
  assign n32838 = ~n40294 & ~n41984;
  assign n32408 = ~n32838;
  assign n32407 = ~n40337 | ~P2_PHYADDRPOINTER_REG_15__SCAN_IN;
  assign n32411 = ~n32408 | ~n32407;
  assign n32409 = ~n39367;
  assign n32410 = ~n32409 & ~n40304;
  assign n32412 = ~n32411 & ~n32410;
  assign n32414 = ~n32413 | ~n32412;
  assign n32416 = ~n32415 & ~n32414;
  assign P2_U2999 = ~n32417 | ~n32416;
  assign n32419 = ~n32418 | ~n32858;
  assign n32430 = ~n32848 & ~n40323;
  assign n39721 = n32421 ^ n32420;
  assign n32428 = ~n39721 | ~n40324;
  assign n32866 = ~n40294 & ~n32422;
  assign n32424 = ~n32866;
  assign n32423 = ~n40337 | ~P2_PHYADDRPOINTER_REG_14__SCAN_IN;
  assign n32426 = ~n32424 | ~n32423;
  assign n32425 = ~n40304 & ~n39379;
  assign n32427 = ~n32426 & ~n32425;
  assign n32429 = ~n32428 | ~n32427;
  assign n32435 = ~n32430 & ~n32429;
  assign n32434 = ~n32876 | ~n32597;
  assign P2_U3000 = ~n32435 | ~n32434;
  assign n32439 = ~n32437 | ~n32436;
  assign n32879 = n32439 ^ n32438;
  assign n32449 = ~n32879 & ~n40342;
  assign n39732 = n32441 ^ n32440;
  assign n32447 = ~n39732 | ~n40324;
  assign n32882 = ~n40325 | ~P2_REIP_REG_13__SCAN_IN;
  assign n32442 = ~n40337 | ~P2_PHYADDRPOINTER_REG_13__SCAN_IN;
  assign n32445 = ~n32882 | ~n32442;
  assign n32443 = ~n39396;
  assign n32444 = ~n40304 & ~n32443;
  assign n32446 = ~n32445 & ~n32444;
  assign n32448 = ~n32447 | ~n32446;
  assign n32451 = ~n32449 & ~n32448;
  assign n32894 = ~n32452 ^ n32849;
  assign n32450 = ~n32894 | ~n40348;
  assign P2_U3001 = ~n32451 | ~n32450;
  assign n32453 = ~n23438 & ~P2_INSTADDRPOINTER_REG_12__SCAN_IN;
  assign n32897 = ~n32453 & ~n32452;
  assign n32467 = ~n32897 | ~n40348;
  assign n32456 = ~n23818 & ~n32455;
  assign n32465 = ~n32898 & ~n40342;
  assign n39741 = n32458 ^ n32457;
  assign n32463 = ~n39741 | ~n40324;
  assign n32905 = ~n40325 | ~P2_REIP_REG_12__SCAN_IN;
  assign n32459 = ~n40337 | ~P2_PHYADDRPOINTER_REG_12__SCAN_IN;
  assign n32461 = ~n32905 | ~n32459;
  assign n32460 = ~n40304 & ~n39419;
  assign n32462 = ~n32461 & ~n32460;
  assign n32464 = ~n32463 | ~n32462;
  assign n32466 = ~n32465 & ~n32464;
  assign P2_U3002 = ~n32467 | ~n32466;
  assign n32480 = ~n32917 & ~n40342;
  assign n39751 = n32472 ^ n32471;
  assign n32478 = ~n39751 | ~n40324;
  assign n32936 = ~n40325 | ~P2_REIP_REG_11__SCAN_IN;
  assign n32473 = ~n40337 | ~P2_PHYADDRPOINTER_REG_11__SCAN_IN;
  assign n32476 = ~n32936 | ~n32473;
  assign n32474 = ~n39453;
  assign n32475 = ~n40304 & ~n32474;
  assign n32477 = ~n32476 & ~n32475;
  assign n32479 = ~n32478 | ~n32477;
  assign n32485 = ~n32480 & ~n32479;
  assign n32504 = ~n32481 | ~n32925;
  assign n32483 = ~n32504 | ~n32927;
  assign n32944 = n32482 & n32483;
  assign n32484 = ~n32944 | ~n40348;
  assign P2_U3003 = ~n32485 | ~n32484;
  assign n32491 = ~n32487 | ~n32486;
  assign n32489 = ~n22986 | ~n32509;
  assign n32490 = ~n32489 | ~n32508;
  assign n32947 = n32491 ^ n32490;
  assign n32501 = ~n32947 & ~n40342;
  assign n39759 = n32493 ^ n32492;
  assign n32499 = ~n39759 | ~n40324;
  assign n32954 = ~n40294 & ~n28382;
  assign n32495 = ~n32954;
  assign n32494 = ~n40337 | ~P2_PHYADDRPOINTER_REG_10__SCAN_IN;
  assign n32497 = ~n32495 | ~n32494;
  assign n32496 = ~n40304 & ~n39461;
  assign n32498 = ~n32497 & ~n32496;
  assign n32500 = ~n32499 | ~n32498;
  assign n32507 = ~n32501 & ~n32500;
  assign n32503 = ~n32481 | ~P2_INSTADDRPOINTER_REG_9__SCAN_IN;
  assign n32505 = ~n32503 | ~n32502;
  assign n32964 = n32505 & n32504;
  assign n32506 = ~n32964 | ~n40348;
  assign P2_U3004 = ~n32507 | ~n32506;
  assign n32967 = ~n32481 ^ n32975;
  assign n32523 = ~n32967 | ~n40348;
  assign n32510 = n32509 & n32508;
  assign n32968 = ~n22986 ^ n32510;
  assign n32521 = n32968 | n40342;
  assign n39492 = ~n32511 ^ n32512;
  assign n32519 = n39492 | n40344;
  assign n32514 = n40294 | n32974;
  assign n32513 = ~n40337 | ~P2_PHYADDRPOINTER_REG_9__SCAN_IN;
  assign n32517 = ~n32514 | ~n32513;
  assign n32515 = ~n39485;
  assign n32516 = ~n40304 & ~n32515;
  assign n32518 = ~n32517 & ~n32516;
  assign n32520 = n32519 & n32518;
  assign n32522 = n32521 & n32520;
  assign P2_U3005 = ~n32523 | ~n32522;
  assign n32546 = ~n32989 | ~n40348;
  assign n32528 = n32526 & n32525;
  assign n32548 = ~n32528 | ~n32527;
  assign n32547 = ~n32529 ^ P2_INSTADDRPOINTER_REG_7__SCAN_IN;
  assign n32531 = ~n32548 | ~n32547;
  assign n32535 = ~n32531 | ~n32530;
  assign n32534 = ~n32533 | ~n32532;
  assign n32990 = ~n32535 ^ n32534;
  assign n32544 = ~n32990 | ~n32597;
  assign n39496 = ~n32537 ^ n32536;
  assign n32540 = ~n39496 & ~n40344;
  assign n33008 = ~n40325 | ~P2_REIP_REG_8__SCAN_IN;
  assign n32538 = ~n40337 | ~P2_PHYADDRPOINTER_REG_8__SCAN_IN;
  assign n32539 = ~n33008 | ~n32538;
  assign n32542 = n32540 | n32539;
  assign n32541 = ~n40304 & ~n39511;
  assign n32543 = ~n32542 & ~n32541;
  assign n32545 = n32544 & n32543;
  assign P2_U3006 = ~n32546 | ~n32545;
  assign n33022 = ~n32548 ^ n32547;
  assign n32558 = ~n33022 & ~n40342;
  assign n39787 = n32550 ^ n32549;
  assign n32556 = ~n39787 | ~n40324;
  assign n33030 = ~n40325 | ~P2_REIP_REG_7__SCAN_IN;
  assign n32551 = ~n40337 | ~P2_PHYADDRPOINTER_REG_7__SCAN_IN;
  assign n32554 = ~n33030 | ~n32551;
  assign n32552 = ~n39531;
  assign n32553 = ~n40304 & ~n32552;
  assign n32555 = ~n32554 & ~n32553;
  assign n32557 = ~n32556 | ~n32555;
  assign n32561 = ~n32558 & ~n32557;
  assign n33039 = ~n22998 ^ n32559;
  assign n32560 = ~n33039 | ~n40348;
  assign P2_U3007 = ~n32561 | ~n32560;
  assign n33042 = ~n32562 ^ P2_INSTADDRPOINTER_REG_6__SCAN_IN;
  assign n32572 = ~n33042 & ~n40323;
  assign n39543 = ~n32564 ^ n32563;
  assign n39794 = ~n39543;
  assign n32570 = ~n39794 | ~n40324;
  assign n33048 = ~n28354 & ~n40294;
  assign n32566 = ~n33048;
  assign n32565 = ~n40337 | ~P2_PHYADDRPOINTER_REG_6__SCAN_IN;
  assign n32568 = ~n32566 | ~n32565;
  assign n32567 = ~n40304 & ~n39550;
  assign n32569 = ~n32568 & ~n32567;
  assign n32571 = ~n32570 | ~n32569;
  assign n32580 = ~n32572 & ~n32571;
  assign n32596 = ~n32573 ^ n33073;
  assign n32576 = ~n32596 | ~n32574;
  assign n32578 = ~n32576 | ~n32575;
  assign n33057 = ~n32578 ^ n32577;
  assign n32579 = ~n33057 | ~n32597;
  assign P2_U3008 = ~n32580 | ~n32579;
  assign n32582 = n32581;
  assign n32584 = ~n32583 | ~n32582;
  assign n33060 = ~n32584 ^ n33073;
  assign n32595 = ~n33060 & ~n40323;
  assign n39802 = n32585 ^ n39582;
  assign n32593 = ~n39802 | ~n40324;
  assign n33077 = ~n40294 & ~n32586;
  assign n32588 = ~n33077;
  assign n32587 = ~n40337 | ~P2_PHYADDRPOINTER_REG_5__SCAN_IN;
  assign n32591 = ~n32588 | ~n32587;
  assign n32589 = ~n39565;
  assign n32590 = ~n40304 & ~n32589;
  assign n32592 = ~n32591 & ~n32590;
  assign n32594 = ~n32593 | ~n32592;
  assign n32599 = ~n32595 & ~n32594;
  assign n33087 = n32574 ^ n32596;
  assign n32598 = ~n33087 | ~n32597;
  assign P2_U3009 = ~n32599 | ~n32598;
  assign n32600 = ~n39613 | ~n40330;
  assign n33092 = ~n40325 | ~P2_REIP_REG_3__SCAN_IN;
  assign n32610 = ~n32600 | ~n33092;
  assign n32601 = ~n32602;
  assign n32603 = ~n32601 | ~P2_INSTADDRPOINTER_REG_3__SCAN_IN;
  assign n40286 = ~n32602 | ~n33104;
  assign n40285 = ~n32603 | ~n40286;
  assign n33098 = n40284 ^ n40285;
  assign n32606 = ~n33098 & ~n40342;
  assign n33099 = ~n22845 | ~n32604;
  assign n32605 = ~n33099 & ~n40323;
  assign n32608 = ~n32606 & ~n32605;
  assign n32607 = ~P2_PHYADDRPOINTER_REG_3__SCAN_IN | ~n40337;
  assign n32609 = ~n32608 | ~n32607;
  assign n32612 = ~n32610 & ~n32609;
  assign n32611 = ~n33144 | ~n40324;
  assign P2_U3011 = ~n32612 | ~n32611;
  assign n32631 = ~n32613 | ~n40356;
  assign n32629 = ~n32614 & ~n40397;
  assign n32624 = ~n32615 | ~n40408;
  assign n32622 = ~n32616 & ~n32617;
  assign n32620 = ~n32618 | ~n32617;
  assign n32621 = ~n32620 | ~n32619;
  assign n32623 = ~n32622 & ~n32621;
  assign n32627 = n32624 & n32623;
  assign n32626 = ~n32625 | ~n33115;
  assign n32628 = ~n32627 | ~n32626;
  assign n32630 = ~n32629 & ~n32628;
  assign P2_U3016 = ~n32631 | ~n32630;
  assign n32647 = ~n32632 & ~n40397;
  assign n32636 = ~n32635;
  assign n32652 = ~n32637 | ~n32636;
  assign n32644 = ~P2_INSTADDRPOINTER_REG_29__SCAN_IN | ~n32652;
  assign n32639 = ~n32638 ^ P2_INSTADDRPOINTER_REG_28__SCAN_IN;
  assign n32640 = ~P2_INSTADDRPOINTER_REG_27__SCAN_IN | ~n32639;
  assign n32642 = ~n32655 & ~n32640;
  assign n32643 = ~n32642 & ~n32641;
  assign n32645 = ~n32644 | ~n32643;
  assign n32648 = ~n32647 & ~n32646;
  assign P2_U3017 = ~n32649 | ~n32648;
  assign n32663 = ~n32650 | ~n40408;
  assign n32661 = ~n32651 & ~n40399;
  assign n32659 = ~P2_INSTADDRPOINTER_REG_28__SCAN_IN | ~n32652;
  assign n32654 = ~n32653 | ~P2_INSTADDRPOINTER_REG_27__SCAN_IN;
  assign n32657 = ~n32655 & ~n32654;
  assign n32658 = ~n32657 & ~n32656;
  assign n32660 = ~n32659 | ~n32658;
  assign n32662 = ~n32661 & ~n32660;
  assign n32664 = ~n32663 | ~n32662;
  assign n32667 = ~n32665 & ~n32664;
  assign P2_U3018 = ~n32667 | ~n32666;
  assign n32685 = ~n32668 | ~n40408;
  assign n32683 = ~n32669 | ~n33115;
  assign n32692 = ~n32713 | ~P2_INSTADDRPOINTER_REG_24__SCAN_IN;
  assign n32670 = ~P2_INSTADDRPOINTER_REG_26__SCAN_IN ^ P2_INSTADDRPOINTER_REG_25__SCAN_IN;
  assign n32681 = ~n32692 & ~n32670;
  assign n32672 = ~P2_INSTADDRPOINTER_REG_24__SCAN_IN | ~n32671;
  assign n32675 = ~n32672 | ~n33062;
  assign n32674 = ~n32996 | ~n32673;
  assign n32676 = ~n32675 | ~n32674;
  assign n32711 = ~n40403 & ~n32676;
  assign n32677 = ~n32996 | ~n32712;
  assign n32691 = ~n32711 | ~n32677;
  assign n32678 = ~P2_INSTADDRPOINTER_REG_26__SCAN_IN | ~n32691;
  assign n32680 = ~n32679 | ~n32678;
  assign n32682 = ~n32681 & ~n32680;
  assign n32684 = n32683 & n32682;
  assign n32686 = ~n32685 | ~n32684;
  assign n32689 = ~n32687 & ~n32686;
  assign P2_U3020 = ~n32689 | ~n32688;
  assign n32698 = ~n32690 & ~n33125;
  assign n32694 = n32691 | n23751;
  assign n32693 = ~n32692 | ~n23751;
  assign n32696 = ~n32694 | ~n32693;
  assign n32697 = ~n32696 | ~n32695;
  assign n32701 = ~n32698 & ~n32697;
  assign n32700 = ~n32699 | ~n33115;
  assign n32702 = ~n32701 | ~n32700;
  assign n32706 = ~n32703 & ~n32702;
  assign n32705 = ~n32704 | ~n33086;
  assign P2_U3021 = ~n32706 | ~n32705;
  assign n32725 = ~n32707 | ~n40356;
  assign n32723 = n32708 | n40397;
  assign n32721 = n32709 | n33125;
  assign n32719 = ~n32710 & ~n40399;
  assign n32717 = ~n32711 & ~n32712;
  assign n32715 = ~n32713 | ~n32712;
  assign n32716 = ~n32715 | ~n32714;
  assign n32718 = n32717 | n32716;
  assign n32720 = ~n32719 & ~n32718;
  assign n32722 = n32721 & n32720;
  assign n32724 = n32723 & n32722;
  assign P2_U3022 = ~n32725 | ~n32724;
  assign n32749 = ~n32726 | ~n40356;
  assign n32747 = ~n32727 & ~n40397;
  assign n32729 = ~n32728;
  assign n32742 = ~n32729 & ~n33125;
  assign n32730 = ~P2_INSTADDRPOINTER_REG_22__SCAN_IN & ~n32734;
  assign n32756 = ~P2_INSTADDRPOINTER_REG_21__SCAN_IN | ~n32730;
  assign n32731 = ~n40390 & ~P2_INSTADDRPOINTER_REG_21__SCAN_IN;
  assign n32753 = ~n32732 & ~n32731;
  assign n32733 = ~n32756 | ~n32753;
  assign n32740 = ~n32733 | ~P2_INSTADDRPOINTER_REG_23__SCAN_IN;
  assign n32735 = ~P2_INSTADDRPOINTER_REG_23__SCAN_IN & ~n32734;
  assign n32738 = ~n32736 | ~n32735;
  assign n32739 = n32738 & n32737;
  assign n32741 = ~n32740 | ~n32739;
  assign n32745 = ~n32742 & ~n32741;
  assign n32744 = ~n32743 | ~n33115;
  assign n32746 = ~n32745 | ~n32744;
  assign n32748 = ~n32747 & ~n32746;
  assign P2_U3023 = ~n32749 | ~n32748;
  assign n32763 = ~n32751 & ~n40397;
  assign n32761 = ~n39214 | ~n40408;
  assign n32759 = ~n39224 & ~n40399;
  assign n32755 = ~n32753 & ~n32752;
  assign n32757 = ~n32755 & ~n32754;
  assign n32758 = ~n32757 | ~n32756;
  assign n32760 = ~n32759 & ~n32758;
  assign n32762 = ~n32761 | ~n32760;
  assign n32764 = ~n32763 & ~n32762;
  assign P2_U3024 = ~n32765 | ~n32764;
  assign n32767 = ~n39275 | ~n40408;
  assign n32769 = ~n32767 | ~n32766;
  assign n32768 = ~n39270 & ~n40399;
  assign n32776 = ~n32769 & ~n32768;
  assign n32774 = ~n32770 & ~P2_INSTADDRPOINTER_REG_19__SCAN_IN;
  assign n32773 = ~n32772 & ~n32771;
  assign n32775 = n32774 | n32773;
  assign n32777 = ~n32776 | ~n32775;
  assign n32779 = ~n32778 & ~n32777;
  assign P2_U3027 = ~n32780 | ~n32779;
  assign n32797 = ~n32781 | ~n33086;
  assign n32783 = ~n32782 | ~n40356;
  assign n32795 = ~n22887 & ~n32783;
  assign n32790 = ~n39308 | ~n40408;
  assign n32788 = ~n39290 & ~n40399;
  assign n32785 = ~P2_INSTADDRPOINTER_REG_18__SCAN_IN | ~n32784;
  assign n32787 = ~n32786 | ~n32785;
  assign n32789 = ~n32788 & ~n32787;
  assign n32793 = ~n32790 | ~n32789;
  assign n32792 = ~P2_INSTADDRPOINTER_REG_18__SCAN_IN & ~n32791;
  assign n32794 = n32793 | n32792;
  assign n32796 = ~n32795 & ~n32794;
  assign P2_U3028 = ~n32797 | ~n32796;
  assign n32816 = ~n32798 | ~n33086;
  assign n32801 = n32831 | n32800;
  assign n32802 = ~n33062 | ~n32801;
  assign n32832 = ~n32803 | ~n32802;
  assign n40412 = ~n33124;
  assign n32804 = ~n40412 & ~P2_INSTADDRPOINTER_REG_16__SCAN_IN;
  assign n32805 = ~n32804 & ~n32808;
  assign n32810 = ~n32817 | ~n32805;
  assign n32806 = ~n32830;
  assign n32812 = ~n39325 | ~n40408;
  assign n32814 = ~n32812 | ~n32811;
  assign n32813 = ~n39328 & ~n40399;
  assign n32815 = ~n32814 & ~n32813;
  assign n32820 = ~n32817 | ~P2_INSTADDRPOINTER_REG_16__SCAN_IN;
  assign n32822 = ~n39704 | ~n40408;
  assign n32825 = ~n32822 | ~n32821;
  assign n39351 = ~n23171 ^ n32823;
  assign n32824 = ~n39351 & ~n40399;
  assign n32826 = ~n32825 & ~n32824;
  assign n32828 = ~n32827 | ~n33086;
  assign n32847 = ~n32829 | ~n33086;
  assign n32834 = ~n32830 & ~P2_INSTADDRPOINTER_REG_15__SCAN_IN;
  assign n32833 = ~n32832 & ~n32831;
  assign n32843 = ~n32834 & ~n32833;
  assign n32841 = ~n39713 | ~n40408;
  assign n32836 = n32862 | n32835;
  assign n39846 = ~n23171 | ~n32836;
  assign n32839 = ~n39846 & ~n40399;
  assign n32840 = ~n32839 & ~n32838;
  assign n32842 = ~n32841 | ~n32840;
  assign n32844 = n32843 | n32842;
  assign n32846 = ~n32845 & ~n32844;
  assign P2_U3031 = ~n32847 | ~n32846;
  assign n32875 = ~n32848 & ~n23239;
  assign n32850 = ~P2_INSTADDRPOINTER_REG_12__SCAN_IN | ~n32849;
  assign n32889 = ~n32861 & ~n32850;
  assign n32854 = ~n33124 | ~n32851;
  assign n32918 = ~n32852;
  assign n32853 = ~n33062 | ~n32918;
  assign n32855 = ~n32854 | ~n32853;
  assign n32900 = ~n32855 & ~n32921;
  assign n32856 = ~n32861;
  assign n32909 = ~n32856 | ~n32899;
  assign n32880 = ~n32900 | ~n32909;
  assign n32857 = ~n32889 & ~n32880;
  assign n32873 = ~n32858 & ~n32857;
  assign n32860 = ~n32859 | ~n32858;
  assign n32871 = ~n32861 & ~n32860;
  assign n32869 = ~n39721 | ~n40408;
  assign n32865 = ~n32862;
  assign n32864 = ~n32885 | ~n32863;
  assign n39855 = ~n32865 | ~n32864;
  assign n32867 = ~n39855 & ~n40399;
  assign n32868 = ~n32867 & ~n32866;
  assign n32870 = ~n32869 | ~n32868;
  assign n32872 = n32871 | n32870;
  assign n32874 = n32873 | n32872;
  assign n32878 = ~n32875 & ~n32874;
  assign n32877 = ~n32876 | ~n33086;
  assign P2_U3032 = ~n32878 | ~n32877;
  assign n32893 = ~n32879 & ~n40397;
  assign n32881 = ~P2_INSTADDRPOINTER_REG_13__SCAN_IN | ~n32880;
  assign n32891 = ~n32882 | ~n32881;
  assign n32887 = ~n39732 | ~n40408;
  assign n32884 = ~n32904 | ~n32883;
  assign n39405 = n32885 & n32884;
  assign n32886 = ~n39405 | ~n33115;
  assign n32888 = ~n32887 | ~n32886;
  assign n32890 = n32889 | n32888;
  assign n32892 = n32891 | n32890;
  assign n32896 = ~n32893 & ~n32892;
  assign n32895 = ~n32894 | ~n40356;
  assign P2_U3033 = ~n32896 | ~n32895;
  assign n32916 = ~n32897 | ~n40356;
  assign n32914 = ~n32898 & ~n40397;
  assign n32912 = ~n32900 & ~n32899;
  assign n32901 = ~n39741;
  assign n32908 = ~n32901 & ~n33125;
  assign n32903 = ~n32931 | ~n32902;
  assign n39429 = n32904 & n32903;
  assign n32906 = ~n39429 | ~n33115;
  assign n32907 = ~n32906 | ~n32905;
  assign n32910 = ~n32908 & ~n32907;
  assign n32911 = ~n32910 | ~n32909;
  assign n32913 = n32912 | n32911;
  assign n32915 = ~n32914 & ~n32913;
  assign P2_U3034 = ~n32916 | ~n32915;
  assign n32943 = ~n32917 & ~n40397;
  assign n32919 = ~n32918 & ~n32975;
  assign n32920 = ~n32993 & ~n32919;
  assign n32976 = ~n32921 & ~n32920;
  assign n32922 = ~n32996 | ~n32975;
  assign n32948 = ~n32976 | ~n32922;
  assign n32924 = ~n32927 & ~n32948;
  assign n32923 = ~P2_INSTADDRPOINTER_REG_10__SCAN_IN & ~n32975;
  assign n32949 = ~n32969 | ~n32923;
  assign n32929 = ~n32924 | ~n32949;
  assign n32926 = ~n32925 | ~n32969;
  assign n32928 = ~n32927 | ~n32926;
  assign n32941 = ~n32929 | ~n32928;
  assign n32930 = ~n39751;
  assign n32939 = ~n32930 & ~n33125;
  assign n32935 = ~n32931;
  assign n32934 = ~n32950 & ~n32933;
  assign n39870 = ~n28836 & ~n32934;
  assign n32937 = ~n39870 | ~n33115;
  assign n32938 = ~n32937 | ~n32936;
  assign n32940 = ~n32939 & ~n32938;
  assign n32942 = ~n32941 | ~n32940;
  assign n32946 = ~n32943 & ~n32942;
  assign n32945 = ~n32944 | ~n40356;
  assign P2_U3035 = ~n32946 | ~n32945;
  assign n32963 = ~n32947 & ~n40397;
  assign n32961 = ~n32948 | ~P2_INSTADDRPOINTER_REG_10__SCAN_IN;
  assign n32959 = ~n32949;
  assign n32957 = ~n39759 | ~n40408;
  assign n32953 = ~n32950;
  assign n32952 = ~n32973 | ~n32951;
  assign n39876 = ~n32953 | ~n32952;
  assign n32955 = ~n39876 & ~n40399;
  assign n32956 = ~n32955 & ~n32954;
  assign n32958 = ~n32957 | ~n32956;
  assign n32960 = ~n32959 & ~n32958;
  assign n32962 = ~n32961 | ~n32960;
  assign n32966 = ~n32963 & ~n32962;
  assign n32965 = ~n32964 | ~n40356;
  assign P2_U3036 = ~n32966 | ~n32965;
  assign n32988 = ~n32967 | ~n40356;
  assign n32986 = ~n32968 & ~n40397;
  assign n32984 = ~n32969 | ~n32975;
  assign n32982 = ~n39492 & ~n33125;
  assign n32972 = ~n32970 | ~n32971;
  assign n39881 = n32973 & n32972;
  assign n32980 = ~n39881 | ~n33115;
  assign n32978 = ~n40294 & ~n32974;
  assign n32977 = ~n32976 & ~n32975;
  assign n32979 = ~n32978 & ~n32977;
  assign n32981 = ~n32980 | ~n32979;
  assign n32983 = ~n32982 & ~n32981;
  assign n32985 = ~n32984 | ~n32983;
  assign n32987 = ~n32986 & ~n32985;
  assign P2_U3037 = ~n32988 | ~n32987;
  assign n33021 = ~n32989 | ~n40356;
  assign n33019 = n32990 & n33086;
  assign n32992 = ~n33003 & ~n32991;
  assign n32994 = ~n32993 & ~n32992;
  assign n32998 = ~n40403 & ~n32994;
  assign n32997 = ~n32996 | ~n32995;
  assign n33043 = ~n32998 | ~n32997;
  assign n32999 = ~n40390 & ~P2_INSTADDRPOINTER_REG_6__SCAN_IN;
  assign n33024 = ~n33043 & ~n32999;
  assign n40389 = ~P2_INSTADDRPOINTER_REG_2__SCAN_IN | ~n40377;
  assign n33000 = ~n40390 | ~n40389;
  assign n33001 = ~n33000 | ~n33065;
  assign n33105 = ~n40412 & ~n33001;
  assign n33044 = ~n33002 | ~n33105;
  assign n33004 = ~n33003 & ~n33044;
  assign n33029 = ~n33004 | ~n33023;
  assign n33005 = ~n33024 | ~n33029;
  assign n33013 = ~n33005 | ~P2_INSTADDRPOINTER_REG_8__SCAN_IN;
  assign n33011 = ~n39496 & ~n33125;
  assign n33007 = ~n33027 | ~n33006;
  assign n39497 = n32970 & n33007;
  assign n33009 = ~n39497 | ~n33115;
  assign n33010 = ~n33009 | ~n33008;
  assign n33012 = ~n33011 & ~n33010;
  assign n33017 = n33013 & n33012;
  assign n33014 = ~P2_INSTADDRPOINTER_REG_8__SCAN_IN & ~n33044;
  assign n33016 = ~n33015 | ~n33014;
  assign n33018 = ~n33017 | ~n33016;
  assign n33020 = ~n33019 & ~n33018;
  assign P2_U3038 = ~n33021 | ~n33020;
  assign n33038 = ~n33022 & ~n40397;
  assign n33036 = ~n33024 & ~n33023;
  assign n33034 = ~n39787 | ~n40408;
  assign n33028 = n33026 | n33025;
  assign n39893 = ~n33028 | ~n33027;
  assign n33032 = ~n39893 & ~n40399;
  assign n33031 = ~n33030 | ~n33029;
  assign n33033 = ~n33032 & ~n33031;
  assign n33035 = ~n33034 | ~n33033;
  assign n33037 = n33036 | n33035;
  assign n33041 = ~n33038 & ~n33037;
  assign n33040 = ~n33039 | ~n40356;
  assign P2_U3039 = ~n33041 | ~n33040;
  assign n33056 = ~n33042 & ~n23239;
  assign n33054 = ~n33043 | ~P2_INSTADDRPOINTER_REG_6__SCAN_IN;
  assign n33052 = ~n39543 & ~n33125;
  assign n33050 = P2_INSTADDRPOINTER_REG_6__SCAN_IN | n33044;
  assign n39899 = ~n33046 ^ n33045;
  assign n33047 = ~n40399 & ~n39899;
  assign n33049 = ~n33048 & ~n33047;
  assign n33051 = ~n33050 | ~n33049;
  assign n33053 = ~n33052 & ~n33051;
  assign n33055 = ~n33054 | ~n33053;
  assign n33059 = ~n33056 & ~n33055;
  assign n33058 = ~n33057 | ~n33086;
  assign P2_U3040 = ~n33059 | ~n33058;
  assign n33085 = ~n33060 & ~n23239;
  assign n33063 = ~n33062 | ~n33061;
  assign n40384 = ~n33064 | ~n33063;
  assign n33067 = ~n40384;
  assign n40388 = ~n40390 & ~n33065;
  assign n40378 = ~n32993 & ~P2_INSTADDRPOINTER_REG_2__SCAN_IN;
  assign n33066 = ~n40388 & ~n40378;
  assign n33090 = ~n33067 | ~n33066;
  assign n33068 = ~P2_INSTADDRPOINTER_REG_3__SCAN_IN & ~n40412;
  assign n40367 = ~n33090 & ~n33068;
  assign n33069 = ~n33104 & ~P2_INSTADDRPOINTER_REG_4__SCAN_IN;
  assign n40360 = ~n33105 | ~n33069;
  assign n33070 = ~n40367 | ~n40360;
  assign n33083 = ~n33070 | ~P2_INSTADDRPOINTER_REG_5__SCAN_IN;
  assign n33071 = ~n39802;
  assign n33081 = ~n33071 & ~n33125;
  assign n39558 = n39586 ^ n33072;
  assign n33079 = ~n39558 | ~n33115;
  assign n33075 = ~n33105 | ~n33073;
  assign n33076 = ~n33075 & ~n33074;
  assign n33078 = ~n33077 & ~n33076;
  assign n33080 = ~n33079 | ~n33078;
  assign n33082 = ~n33081 & ~n33080;
  assign n33084 = ~n33083 | ~n33082;
  assign n33089 = ~n33085 & ~n33084;
  assign n33088 = ~n33087 | ~n33086;
  assign P2_U3041 = ~n33089 | ~n33088;
  assign n33091 = ~P2_INSTADDRPOINTER_REG_3__SCAN_IN | ~n33090;
  assign n33097 = ~n33092 | ~n33091;
  assign n33095 = ~n33094 | ~n33093;
  assign n42147 = ~n39588 | ~n33095;
  assign n33096 = ~n40399 & ~n42147;
  assign n33103 = ~n33097 & ~n33096;
  assign n33101 = ~n33098 & ~n40397;
  assign n33100 = ~n33099 & ~n23239;
  assign n33102 = ~n33101 & ~n33100;
  assign n33109 = ~n33103 | ~n33102;
  assign n33107 = ~n33105 | ~n33104;
  assign n33106 = ~n33144 | ~n40408;
  assign n33108 = ~n33107 | ~n33106;
  assign P2_U3043 = n33109 | n33108;
  assign n33110 = ~n39682 | ~n33123;
  assign n40341 = ~n33111 | ~n33110;
  assign n33120 = ~n40397 & ~n40341;
  assign n33114 = ~n33112;
  assign n39963 = ~n33114 ^ n33113;
  assign n33118 = ~n33115 | ~n39963;
  assign n40347 = ~n33116 ^ n33123;
  assign n33117 = ~n40356 | ~n40347;
  assign n33119 = ~n33118 | ~n33117;
  assign n33122 = ~n33120 & ~n33119;
  assign n33121 = ~n40403 | ~P2_INSTADDRPOINTER_REG_0__SCAN_IN;
  assign n33130 = ~n33122 | ~n33121;
  assign n33128 = ~n33124 | ~n33123;
  assign n33126 = ~n33125 & ~n40343;
  assign n40346 = ~n40294 & ~n23399;
  assign n33127 = ~n33126 & ~n40346;
  assign n33129 = ~n33128 | ~n33127;
  assign P2_U3046 = n33130 | n33129;
  assign n41884 = ~n42204 & ~n33131;
  assign n33132 = ~n33217 & ~n33265;
  assign n33134 = ~n41884 & ~n33132;
  assign n33258 = ~n33134 | ~n33133;
  assign n33252 = n27605 | n33135;
  assign n33138 = ~n39973 & ~n33236;
  assign n33139 = ~n33138 & ~n33137;
  assign n33142 = ~n33140 | ~n33139;
  assign n33183 = ~n33143;
  assign n33157 = ~n33144 | ~n33143;
  assign n33148 = ~n23571 | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n33149 = ~n33148 | ~n33147;
  assign n33152 = ~n33164 | ~n33149;
  assign n33160 = n27433 & n27348;
  assign n33150 = ~n33160 ^ P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n33161 = ~n33229 | ~n33230;
  assign n33151 = ~n33150 | ~n33161;
  assign n33155 = ~n33152 | ~n33151;
  assign n33153 = ~n33165 ^ P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n33154 = n33184 & n33153;
  assign n33156 = ~n33155 & ~n33154;
  assign n42086 = n33157 & n33156;
  assign n33159 = n42076 | n42086;
  assign n33158 = ~n42076 | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n33201 = n33159 & n33158;
  assign n33175 = ~n42076 | ~n27348;
  assign n33173 = ~n33161 | ~n33162;
  assign n33163 = ~n33162;
  assign n33171 = n33164 & n33163;
  assign n33169 = ~n27757 | ~n33143;
  assign n33212 = ~n33165;
  assign n33166 = ~n42120 & ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n33167 = ~n33212 & ~n33166;
  assign n33168 = ~n33167 | ~n33184;
  assign n33170 = ~n33169 | ~n33168;
  assign n33172 = ~n33171 & ~n33170;
  assign n42102 = ~n33173 | ~n33172;
  assign n33174 = n42076 | n42102;
  assign n33196 = ~n33175 | ~n33174;
  assign n33211 = ~n33201 & ~n33196;
  assign n33182 = ~n33176 | ~n33143;
  assign n33177 = ~n33184;
  assign n33180 = ~n33177 & ~n42120;
  assign n33178 = ~n33185;
  assign n33179 = ~n33178 & ~n23962;
  assign n33181 = ~n33180 & ~n33179;
  assign n42116 = ~n33182 | ~n33181;
  assign n33190 = n40343 | n33183;
  assign n33188 = n33184 | n33186;
  assign n33187 = ~n33178 | ~n33186;
  assign n33189 = ~n33188 | ~n33187;
  assign n42125 = n33190 & n33189;
  assign n33192 = ~P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN | ~n42125;
  assign n33191 = ~n42116 & ~n33192;
  assign n33195 = ~n33191 & ~n42076;
  assign n33193 = ~n42116 | ~n33192;
  assign n33194 = ~P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~n33193;
  assign n33198 = ~n33195 | ~n33194;
  assign n33197 = n33198 & P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign n33200 = ~n33197 & ~n33196;
  assign n33199 = ~n33198 & ~P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign n33203 = ~n33201;
  assign n33202 = ~n33204 & ~n33203;
  assign n33207 = ~n33202 & ~P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN;
  assign n33205 = ~n33204 | ~n33203;
  assign n33206 = ~P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | ~n33205;
  assign n33209 = ~n33207 | ~n33206;
  assign n33208 = ~P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN | ~n42076;
  assign n33210 = ~n33209 | ~n33208;
  assign n33248 = ~n33211 & ~n33210;
  assign n33214 = ~n33212 | ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n33215 = ~n33214 | ~n33213;
  assign n33216 = ~n42208 | ~n33215;
  assign n42082 = ~n39140 & ~n33216;
  assign n33219 = ~n33217;
  assign n33227 = ~n33219 & ~n33218;
  assign n33225 = ~n33221 | ~n33220;
  assign n33222 = ~n33240;
  assign n33224 = ~n33223 | ~n33222;
  assign n33226 = ~n33225 | ~n33224;
  assign n33235 = ~n33227 & ~n33226;
  assign n33233 = ~n33229 & ~n33228;
  assign n33232 = ~n33231 & ~n33230;
  assign n33234 = ~n33233 & ~n33232;
  assign n42192 = ~n33235 | ~n33234;
  assign n33238 = ~n33237 | ~n33236;
  assign n33241 = ~n33239 & ~n33238;
  assign n39161 = ~n33241 | ~n33240;
  assign n33242 = ~P2_MORE_REG_SCAN_IN & ~P2_FLUSH_REG_SCAN_IN;
  assign n33243 = ~n39161 & ~n33242;
  assign n33244 = ~n42192 & ~n33243;
  assign n33246 = ~n33245 | ~n33244;
  assign n33247 = ~n42082 & ~n33246;
  assign n33254 = ~n33248 | ~n33247;
  assign n33249 = ~P2_STATE2_REG_0__SCAN_IN | ~n22963;
  assign n33250 = ~n33249 | ~P2_STATE2_REG_2__SCAN_IN;
  assign n33251 = ~n42197 & ~n33250;
  assign n41890 = ~n33252 | ~n33251;
  assign n33253 = ~n41890;
  assign n33256 = ~P2_STATE2_REG_0__SCAN_IN | ~n33253;
  assign n33255 = ~n33254 | ~n39160;
  assign n33257 = ~n33256 | ~n33255;
  assign n33263 = ~n33258 & ~n33257;
  assign n33259 = ~n42111 | ~n42214;
  assign n33261 = ~n33259 | ~n42206;
  assign n41885 = ~n42204 & ~n41890;
  assign n33260 = ~n41885;
  assign n33262 = ~n33261 | ~n33260;
  assign P2_U3176 = ~n33263 | ~n33262;
  assign n33264 = ~n41890 | ~P2_STATE2_REG_0__SCAN_IN;
  assign n33266 = ~n33264 | ~P2_STATE2_REG_3__SCAN_IN;
  assign P2_U3593 = ~n33266 | ~n33265;
  assign n33269 = n33267 & n36497;
  assign n33275 = ~n33269 & ~n33268;
  assign n39046 = ~P3_INSTADDRPOINTER_REG_31__SCAN_IN;
  assign n33363 = ~n39046 | ~P3_INSTADDRPOINTER_REG_30__SCAN_IN;
  assign n33274 = ~n33275 | ~n33363;
  assign n33272 = ~n36497 | ~n39046;
  assign n33270 = ~n24287 & ~n39046;
  assign n33271 = ~n36610 | ~n33270;
  assign n33273 = ~n33272 | ~n33271;
  assign n33281 = ~n33274 | ~n33273;
  assign n33277 = ~n33276 | ~n24287;
  assign n33278 = ~n33277 | ~P3_INSTADDRPOINTER_REG_31__SCAN_IN;
  assign n33280 = ~n33279 | ~n33278;
  assign n33283 = ~n38677 & ~n37363;
  assign n33282 = ~n38675 & ~n38674;
  assign n38668 = ~n33283 & ~n33282;
  assign n33348 = ~P3_PHYADDRPOINTER_REG_29__SCAN_IN;
  assign n36229 = ~P3_PHYADDRPOINTER_REG_23__SCAN_IN;
  assign n34343 = ~P3_PHYADDRPOINTER_REG_5__SCAN_IN;
  assign n36686 = ~P3_PHYADDRPOINTER_REG_2__SCAN_IN | ~P3_PHYADDRPOINTER_REG_3__SCAN_IN;
  assign n33285 = ~n36686;
  assign n36639 = ~n36653 | ~P3_PHYADDRPOINTER_REG_6__SCAN_IN;
  assign n33286 = ~n36622 & ~n36590;
  assign n36537 = ~P3_PHYADDRPOINTER_REG_10__SCAN_IN | ~n33286;
  assign n33820 = ~n36537 & ~n36538;
  assign n33822 = ~n36511 & ~n36483;
  assign n33287 = ~n33822;
  assign n36405 = ~P3_PHYADDRPOINTER_REG_15__SCAN_IN | ~P3_PHYADDRPOINTER_REG_16__SCAN_IN;
  assign n33811 = ~P3_PHYADDRPOINTER_REG_18__SCAN_IN | ~P3_PHYADDRPOINTER_REG_19__SCAN_IN;
  assign n36205 = ~P3_PHYADDRPOINTER_REG_24__SCAN_IN;
  assign n33803 = ~n36205 & ~n36183;
  assign n33288 = ~P3_PHYADDRPOINTER_REG_30__SCAN_IN | ~n33322;
  assign n36751 = ~n33749;
  assign n33729 = ~n38803 | ~n38487;
  assign n39104 = n33729 & n39056;
  assign n33289 = ~P3_STATE2_REG_0__SCAN_IN & ~n39104;
  assign n36112 = ~P3_STATEBS16_REG_SCAN_IN;
  assign n33794 = ~P3_STATE2_REG_1__SCAN_IN | ~n36112;
  assign n33303 = ~n34425 | ~n36389;
  assign n33292 = P3_PHYADDRPOINTER_REG_31__SCAN_IN ^ P3_PHYADDRPOINTER_REG_30__SCAN_IN;
  assign n37441 = ~n38483;
  assign n39038 = ~n38487 & ~P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN;
  assign n33290 = ~n38811 | ~n37396;
  assign n37436 = ~n39068 | ~n33290;
  assign n38115 = ~n37441 & ~n38489;
  assign n34460 = ~P3_PHYADDRPOINTER_REG_1__SCAN_IN;
  assign n36478 = ~n39118 | ~P3_STATE2_REG_2__SCAN_IN;
  assign n36262 = ~n36743 | ~n36745;
  assign n33291 = ~n34460 & ~n36262;
  assign n36484 = ~n38115 & ~n33291;
  assign n33299 = ~n33342 | ~P3_PHYADDRPOINTER_REG_29__SCAN_IN;
  assign n33315 = ~n36484 & ~n33299;
  assign n33298 = ~n33292 | ~n33315;
  assign n33376 = ~n22843 | ~P3_REIP_REG_31__SCAN_IN;
  assign n33293 = ~n33307 | ~P3_INSTADDRPOINTER_REG_30__SCAN_IN;
  assign n33369 = ~P3_INSTADDRPOINTER_REG_31__SCAN_IN ^ n33293;
  assign n33296 = n36490 & n33369;
  assign n36691 = ~n33749 & ~n35948;
  assign n33372 = n33294 ^ P3_INSTADDRPOINTER_REG_31__SCAN_IN;
  assign n33295 = ~n36731 & ~n33372;
  assign n33297 = ~n33296 & ~n33295;
  assign n33343 = ~n38115 | ~n33299;
  assign n33300 = ~n36745 | ~n33801;
  assign n33301 = ~n33343 | ~n33300;
  assign n33347 = ~n36666 & ~n33301;
  assign n36390 = ~n36262;
  assign n33349 = ~n36390 | ~n33348;
  assign n33317 = ~n33347 | ~n33349;
  assign n33302 = ~P3_PHYADDRPOINTER_REG_31__SCAN_IN | ~n33317;
  assign P3_U2799 = ~n33305 | ~n33304;
  assign n33330 = ~n33306 & ~n36580;
  assign n33309 = n33338 | n36731;
  assign n33308 = ~n33307;
  assign n33339 = ~n36490 | ~n33308;
  assign n33310 = ~n33309 | ~n33339;
  assign n33328 = ~n33310 | ~P3_INSTADDRPOINTER_REG_30__SCAN_IN;
  assign n33312 = ~n36832 | ~n36490;
  assign n33311 = ~n36833 | ~n36691;
  assign n36220 = ~n33312 | ~n33311;
  assign n36172 = ~P3_INSTADDRPOINTER_REG_24__SCAN_IN | ~n36220;
  assign n36142 = ~n36781 & ~n36172;
  assign n33314 = ~n36142 | ~n24287;
  assign n33326 = ~n33314 & ~n33313;
  assign n33316 = ~n33315;
  assign n33321 = ~P3_PHYADDRPOINTER_REG_30__SCAN_IN & ~n33316;
  assign n33318 = ~P3_PHYADDRPOINTER_REG_30__SCAN_IN | ~n33317;
  assign n33320 = ~n33319 | ~n33318;
  assign n33324 = ~n33321 & ~n33320;
  assign n33863 = P3_PHYADDRPOINTER_REG_30__SCAN_IN ^ n33322;
  assign n33323 = ~n36389 | ~n33863;
  assign n33325 = ~n33324 | ~n33323;
  assign n33327 = ~n33326 & ~n33325;
  assign n33329 = ~n33328 | ~n33327;
  assign P3_U2800 = n33330 | n33329;
  assign n33334 = ~n33331 | ~n36497;
  assign n33332 = ~n33426;
  assign n33333 = ~n33332 | ~P3_INSTADDRPOINTER_REG_28__SCAN_IN;
  assign n33335 = ~n33334 | ~n33333;
  assign n33402 = ~n33335 ^ P3_INSTADDRPOINTER_REG_29__SCAN_IN;
  assign n33361 = ~n33402 & ~n36580;
  assign n33336 = ~n33428 | ~n33399;
  assign n33337 = ~n33336 | ~n36691;
  assign n33359 = n33338 | n33337;
  assign n33341 = ~n33429 | ~n33399;
  assign n33340 = ~n33339;
  assign n33357 = ~n33341 | ~n33340;
  assign n33344 = ~n33342;
  assign n33345 = ~n33344 & ~n33343;
  assign n33346 = ~P3_PHYADDRPOINTER_REG_29__SCAN_IN & ~n33345;
  assign n33355 = ~n33347 & ~n33346;
  assign n33880 = n33348 ^ n33801;
  assign n33350 = ~n33349 | ~n36508;
  assign n33353 = ~n33880 | ~n33350;
  assign n33351 = ~P3_REIP_REG_29__SCAN_IN;
  assign n33400 = ~n37197 & ~n33351;
  assign n33352 = ~n33400;
  assign n33354 = ~n33353 | ~n33352;
  assign n33356 = ~n33355 & ~n33354;
  assign n33358 = n33357 & n33356;
  assign n33360 = ~n33359 | ~n33358;
  assign P3_U2801 = n33361 | n33360;
  assign n33368 = ~n33363 & ~n33362;
  assign n37300 = ~n37356;
  assign n33364 = ~n37300 & ~P3_INSTADDRPOINTER_REG_30__SCAN_IN;
  assign n33366 = ~n33365 & ~n33364;
  assign n33367 = ~n39046 & ~n33366;
  assign n33371 = ~n33368 & ~n33367;
  assign n33370 = ~n33369 | ~n37147;
  assign n33374 = ~n33371 | ~n33370;
  assign n33373 = ~n38674 & ~n33372;
  assign n33375 = ~n33374 & ~n33373;
  assign n33379 = ~n33375 & ~n37349;
  assign n33377 = ~n37352 | ~P3_INSTADDRPOINTER_REG_31__SCAN_IN;
  assign n33378 = ~n33377 | ~n33376;
  assign n33380 = ~n33379 & ~n33378;
  assign P3_U2831 = ~n33381 | ~n33380;
  assign n33390 = ~P3_INSTADDRPOINTER_REG_28__SCAN_IN & ~n36932;
  assign n36780 = ~P3_INSTADDRPOINTER_REG_27__SCAN_IN | ~n33382;
  assign n33383 = ~n38730 | ~n36780;
  assign n33385 = ~n33384 | ~n33383;
  assign n33387 = ~n33386 & ~n33385;
  assign n33389 = ~n33388 | ~n33387;
  assign n33391 = ~n33390 & ~n33389;
  assign n33392 = ~n33429;
  assign n33398 = ~n33393 | ~n33392;
  assign n33394 = ~n33428 & ~n38674;
  assign n33396 = ~n33395 & ~n33394;
  assign n33397 = P3_INSTADDRPOINTER_REG_29__SCAN_IN | n33396;
  assign n33401 = ~n37383 & ~n33399;
  assign n37165 = ~n37201;
  assign n33403 = ~n33402 & ~n37165;
  assign n36132 = ~n36610 ^ P3_INSTADDRPOINTER_REG_28__SCAN_IN;
  assign n33405 = ~n36151 & ~n36132;
  assign n33404 = ~n36152 | ~n36497;
  assign n36135 = ~n33405 | ~n33404;
  assign n33407 = ~n33406;
  assign n33425 = ~n36135 | ~n33407;
  assign n33409 = ~n33408;
  assign n33422 = ~n33425 & ~n33409;
  assign n33411 = ~n38674 & ~n36321;
  assign n33410 = ~n37184 & ~n36320;
  assign n36987 = ~n33411 & ~n33410;
  assign n33416 = ~n36987 & ~n33412;
  assign n33415 = ~n36879 | ~n38757;
  assign n33414 = ~n33413 | ~n38758;
  assign n36808 = ~n33415 | ~n33414;
  assign n33418 = n33417 & P3_INSTADDRPOINTER_REG_27__SCAN_IN;
  assign n33420 = ~n36760 | ~n33418;
  assign n33421 = ~n33420 | ~n33419;
  assign n33423 = ~n33422 & ~n33421;
  assign n33424 = ~n33423 & ~n37349;
  assign n33445 = n33424 | P3_INSTADDRPOINTER_REG_28__SCAN_IN;
  assign n33427 = ~n33425;
  assign n33441 = ~n33427 | ~n33426;
  assign n33431 = ~n37292 | ~n33428;
  assign n33430 = ~n37147 | ~n33429;
  assign n33439 = ~n33431 | ~n33430;
  assign n36892 = ~n22828 | ~n38673;
  assign n33437 = n36892 & n36764;
  assign n33435 = ~n37352 & ~n33432;
  assign n33434 = ~n33433 | ~n38758;
  assign n33436 = ~n33435 | ~n33434;
  assign n33438 = n33437 | n33436;
  assign n33440 = ~n33439 & ~n33438;
  assign n33442 = ~n33441 | ~n33440;
  assign n33443 = ~n33442 | ~n37197;
  assign n33444 = ~n33443 | ~P3_INSTADDRPOINTER_REG_28__SCAN_IN;
  assign n33450 = ~n33445 | ~n33444;
  assign n33446 = ~n37201 | ~n36132;
  assign n33448 = ~n36152 & ~n33446;
  assign n33447 = ~P3_REIP_REG_28__SCAN_IN;
  assign n36122 = ~n37197 & ~n33447;
  assign n33449 = ~n33448 & ~n36122;
  assign P3_U2834 = ~n33450 | ~n33449;
  assign n33457 = ~P3_BE_N_REG_2__SCAN_IN & ~P3_BE_N_REG_3__SCAN_IN;
  assign n33651 = ~U215;
  assign n33451 = ~P3_W_R_N_REG_SCAN_IN & ~P3_BE_N_REG_1__SCAN_IN;
  assign n33452 = ~P3_M_IO_N_REG_SCAN_IN | ~n33451;
  assign n33454 = ~P3_BE_N_REG_0__SCAN_IN & ~n33452;
  assign n33453 = ~P3_D_C_N_REG_SCAN_IN & ~P3_ADS_N_REG_SCAN_IN;
  assign n33455 = ~n33454 | ~n33453;
  assign n33456 = ~n33651 & ~n33455;
  assign U213 = ~n33457 | ~n33456;
  assign n33459 = ~n39977 & ~U212;
  assign n33656 = ~P1_DATAO_REG_31__SCAN_IN;
  assign n33458 = ~n33656 & ~U214;
  assign n33462 = ~n33459 & ~n33458;
  assign n33461 = ~BUF1_REG_31__SCAN_IN | ~n33585;
  assign U216 = ~n33462 | ~n33461;
  assign n33464 = P2_DATAO_REG_30__SCAN_IN & n33588;
  assign n40532 = ~BUF1_REG_30__SCAN_IN;
  assign n33463 = ~n40532 & ~n33487;
  assign n33466 = ~n33464 & ~n33463;
  assign n33465 = ~P1_DATAO_REG_30__SCAN_IN | ~n33538;
  assign U217 = ~n33466 | ~n33465;
  assign n33468 = P2_DATAO_REG_29__SCAN_IN & n33588;
  assign n40514 = ~BUF1_REG_29__SCAN_IN;
  assign n33467 = ~n40514 & ~n33487;
  assign n33470 = ~n33468 & ~n33467;
  assign n33469 = ~P1_DATAO_REG_29__SCAN_IN | ~n33538;
  assign U218 = ~n33470 | ~n33469;
  assign n33472 = P2_DATAO_REG_28__SCAN_IN & n33588;
  assign n40498 = ~BUF1_REG_28__SCAN_IN;
  assign n33471 = ~n40498 & ~n33487;
  assign n33474 = ~n33472 & ~n33471;
  assign n33473 = ~P1_DATAO_REG_28__SCAN_IN | ~n33538;
  assign U219 = ~n33474 | ~n33473;
  assign n33476 = P2_DATAO_REG_27__SCAN_IN & n33588;
  assign n40483 = ~BUF1_REG_27__SCAN_IN;
  assign n33475 = ~n40483 & ~n33487;
  assign n33478 = ~n33476 & ~n33475;
  assign n33477 = ~P1_DATAO_REG_27__SCAN_IN | ~n33538;
  assign U220 = ~n33478 | ~n33477;
  assign n33480 = P2_DATAO_REG_26__SCAN_IN & n33588;
  assign n40468 = ~BUF1_REG_26__SCAN_IN;
  assign n33479 = ~n40468 & ~n33487;
  assign n33482 = ~n33480 & ~n33479;
  assign n33481 = ~P1_DATAO_REG_26__SCAN_IN | ~n33538;
  assign U221 = ~n33482 | ~n33481;
  assign n33484 = P2_DATAO_REG_25__SCAN_IN & n33588;
  assign n40453 = ~BUF1_REG_25__SCAN_IN;
  assign n33483 = ~n40453 & ~n33487;
  assign n33486 = ~n33484 & ~n33483;
  assign n33485 = ~P1_DATAO_REG_25__SCAN_IN | ~n33538;
  assign U222 = ~n33486 | ~n33485;
  assign n33489 = P2_DATAO_REG_24__SCAN_IN & n33588;
  assign n40445 = ~BUF1_REG_24__SCAN_IN;
  assign n33488 = ~n40445 & ~n33487;
  assign n33491 = ~n33489 & ~n33488;
  assign n33490 = ~P1_DATAO_REG_24__SCAN_IN | ~n33538;
  assign U223 = ~n33491 | ~n33490;
  assign n33493 = ~P1_DATAO_REG_23__SCAN_IN | ~n33538;
  assign n33492 = ~n33585 | ~BUF1_REG_23__SCAN_IN;
  assign n33495 = n33493 & n33492;
  assign n33494 = ~P2_DATAO_REG_23__SCAN_IN | ~n33588;
  assign U224 = ~n33495 | ~n33494;
  assign n33497 = ~P1_DATAO_REG_22__SCAN_IN | ~n33538;
  assign n33496 = ~n33585 | ~BUF1_REG_22__SCAN_IN;
  assign n33499 = n33497 & n33496;
  assign n33498 = ~P2_DATAO_REG_22__SCAN_IN | ~n33588;
  assign U225 = ~n33499 | ~n33498;
  assign n33501 = ~P1_DATAO_REG_21__SCAN_IN | ~n33538;
  assign n33500 = ~n33585 | ~BUF1_REG_21__SCAN_IN;
  assign n33503 = n33501 & n33500;
  assign n33502 = ~P2_DATAO_REG_21__SCAN_IN | ~n33588;
  assign U226 = ~n33503 | ~n33502;
  assign n33505 = ~P1_DATAO_REG_20__SCAN_IN | ~n33538;
  assign n33504 = ~n33585 | ~BUF1_REG_20__SCAN_IN;
  assign n33507 = n33505 & n33504;
  assign n33506 = ~P2_DATAO_REG_20__SCAN_IN | ~n33588;
  assign U227 = ~n33507 | ~n33506;
  assign n33509 = ~P1_DATAO_REG_19__SCAN_IN | ~n33538;
  assign n33508 = ~n33585 | ~BUF1_REG_19__SCAN_IN;
  assign n33511 = n33509 & n33508;
  assign n33510 = ~P2_DATAO_REG_19__SCAN_IN | ~n33588;
  assign U228 = ~n33511 | ~n33510;
  assign n33513 = ~P1_DATAO_REG_18__SCAN_IN | ~n33538;
  assign n33512 = ~n33585 | ~BUF1_REG_18__SCAN_IN;
  assign n33515 = n33513 & n33512;
  assign n33514 = ~P2_DATAO_REG_18__SCAN_IN | ~n33588;
  assign U229 = ~n33515 | ~n33514;
  assign n33517 = ~P1_DATAO_REG_17__SCAN_IN | ~n33538;
  assign n33516 = ~n33585 | ~BUF1_REG_17__SCAN_IN;
  assign n33519 = n33517 & n33516;
  assign n33518 = ~P2_DATAO_REG_17__SCAN_IN | ~n33588;
  assign U230 = ~n33519 | ~n33518;
  assign n33521 = ~P1_DATAO_REG_16__SCAN_IN | ~n33538;
  assign n33520 = ~n33585 | ~BUF1_REG_16__SCAN_IN;
  assign n33523 = n33521 & n33520;
  assign n33522 = ~P2_DATAO_REG_16__SCAN_IN | ~n33588;
  assign U231 = ~n33523 | ~n33522;
  assign n40040 = ~P2_DATAO_REG_15__SCAN_IN;
  assign n33525 = ~n40040 & ~U212;
  assign n33524 = BUF1_REG_15__SCAN_IN & n33585;
  assign n33527 = ~n33525 & ~n33524;
  assign n33526 = ~P1_DATAO_REG_15__SCAN_IN | ~n33538;
  assign U232 = ~n33527 | ~n33526;
  assign n40045 = ~P2_DATAO_REG_14__SCAN_IN;
  assign n33529 = ~n40045 & ~U212;
  assign n33528 = BUF1_REG_14__SCAN_IN & n33585;
  assign n33531 = ~n33529 & ~n33528;
  assign n33530 = ~P1_DATAO_REG_14__SCAN_IN | ~n33538;
  assign U233 = ~n33531 | ~n33530;
  assign n40050 = ~P2_DATAO_REG_13__SCAN_IN;
  assign n33533 = ~n40050 & ~U212;
  assign n33532 = BUF1_REG_13__SCAN_IN & n33585;
  assign n33535 = ~n33533 & ~n33532;
  assign n33534 = ~P1_DATAO_REG_13__SCAN_IN | ~n33538;
  assign U234 = ~n33535 | ~n33534;
  assign n40055 = ~P2_DATAO_REG_12__SCAN_IN;
  assign n33537 = ~n40055 & ~U212;
  assign n33536 = BUF1_REG_12__SCAN_IN & n33585;
  assign n33540 = ~n33537 & ~n33536;
  assign n33539 = ~P1_DATAO_REG_12__SCAN_IN | ~n33538;
  assign U235 = ~n33540 | ~n33539;
  assign n40060 = ~P2_DATAO_REG_11__SCAN_IN;
  assign n33542 = ~n40060 & ~U212;
  assign n33541 = BUF1_REG_11__SCAN_IN & n33585;
  assign n33544 = ~n33542 & ~n33541;
  assign n33543 = ~P1_DATAO_REG_11__SCAN_IN | ~n33538;
  assign U236 = ~n33544 | ~n33543;
  assign n40065 = ~P2_DATAO_REG_10__SCAN_IN;
  assign n33546 = ~n40065 & ~U212;
  assign n33545 = BUF1_REG_10__SCAN_IN & n33585;
  assign n33548 = ~n33546 & ~n33545;
  assign n33547 = ~P1_DATAO_REG_10__SCAN_IN | ~n33538;
  assign U237 = ~n33548 | ~n33547;
  assign n40070 = ~P2_DATAO_REG_9__SCAN_IN;
  assign n33550 = ~n40070 & ~U212;
  assign n33549 = BUF1_REG_9__SCAN_IN & n33585;
  assign n33552 = ~n33550 & ~n33549;
  assign n33551 = ~P1_DATAO_REG_9__SCAN_IN | ~n33538;
  assign U238 = ~n33552 | ~n33551;
  assign n40075 = ~P2_DATAO_REG_8__SCAN_IN;
  assign n33554 = ~n40075 & ~U212;
  assign n33553 = BUF1_REG_8__SCAN_IN & n33585;
  assign n33556 = ~n33554 & ~n33553;
  assign n33555 = ~P1_DATAO_REG_8__SCAN_IN | ~n33538;
  assign U239 = ~n33556 | ~n33555;
  assign n33558 = ~P1_DATAO_REG_7__SCAN_IN | ~n33538;
  assign n33557 = ~n33585 | ~BUF1_REG_7__SCAN_IN;
  assign n33560 = n33558 & n33557;
  assign n33559 = ~P2_DATAO_REG_7__SCAN_IN | ~n33588;
  assign U240 = ~n33560 | ~n33559;
  assign n33562 = ~P1_DATAO_REG_6__SCAN_IN | ~n33538;
  assign n33561 = ~n33585 | ~BUF1_REG_6__SCAN_IN;
  assign n33564 = n33562 & n33561;
  assign n33563 = ~P2_DATAO_REG_6__SCAN_IN | ~n33588;
  assign U241 = ~n33564 | ~n33563;
  assign n33566 = ~P1_DATAO_REG_5__SCAN_IN | ~n33538;
  assign n33565 = ~n33585 | ~BUF1_REG_5__SCAN_IN;
  assign n33568 = n33566 & n33565;
  assign n33567 = ~P2_DATAO_REG_5__SCAN_IN | ~n33588;
  assign U242 = ~n33568 | ~n33567;
  assign n33570 = ~P1_DATAO_REG_4__SCAN_IN | ~n33538;
  assign n33569 = ~n33585 | ~BUF1_REG_4__SCAN_IN;
  assign n33572 = n33570 & n33569;
  assign n33571 = ~P2_DATAO_REG_4__SCAN_IN | ~n33588;
  assign U243 = ~n33572 | ~n33571;
  assign n33574 = ~P1_DATAO_REG_3__SCAN_IN | ~n33538;
  assign n33573 = ~n33585 | ~BUF1_REG_3__SCAN_IN;
  assign n33576 = n33574 & n33573;
  assign n33575 = ~P2_DATAO_REG_3__SCAN_IN | ~n33588;
  assign U244 = ~n33576 | ~n33575;
  assign n33578 = ~P1_DATAO_REG_2__SCAN_IN | ~n33538;
  assign n33577 = ~n33585 | ~BUF1_REG_2__SCAN_IN;
  assign n33580 = n33578 & n33577;
  assign n33579 = ~P2_DATAO_REG_2__SCAN_IN | ~n33588;
  assign U245 = ~n33580 | ~n33579;
  assign n33582 = ~P1_DATAO_REG_1__SCAN_IN | ~n33538;
  assign n33581 = ~n33585 | ~BUF1_REG_1__SCAN_IN;
  assign n33584 = n33582 & n33581;
  assign n33583 = ~P2_DATAO_REG_1__SCAN_IN | ~n33588;
  assign U246 = ~n33584 | ~n33583;
  assign n33587 = ~P1_DATAO_REG_0__SCAN_IN | ~n33538;
  assign n33586 = ~n33585 | ~BUF1_REG_0__SCAN_IN;
  assign n33590 = n33587 & n33586;
  assign n33589 = ~P2_DATAO_REG_0__SCAN_IN | ~n33588;
  assign U247 = ~n33590 | ~n33589;
  assign n33592 = ~BUF2_REG_0__SCAN_IN | ~U215;
  assign n33591 = ~P2_DATAO_REG_0__SCAN_IN | ~n33651;
  assign U251 = ~n33592 | ~n33591;
  assign n33594 = ~U215 | ~BUF2_REG_1__SCAN_IN;
  assign n33593 = ~n33651 | ~P2_DATAO_REG_1__SCAN_IN;
  assign U252 = ~n33594 | ~n33593;
  assign n33596 = ~U215 | ~BUF2_REG_2__SCAN_IN;
  assign n33595 = ~n33651 | ~P2_DATAO_REG_2__SCAN_IN;
  assign U253 = ~n33596 | ~n33595;
  assign n33598 = ~U215 | ~BUF2_REG_3__SCAN_IN;
  assign n33597 = ~n33651 | ~P2_DATAO_REG_3__SCAN_IN;
  assign U254 = ~n33598 | ~n33597;
  assign n33600 = ~U215 | ~BUF2_REG_4__SCAN_IN;
  assign n33599 = ~n33651 | ~P2_DATAO_REG_4__SCAN_IN;
  assign U255 = ~n33600 | ~n33599;
  assign n33602 = ~U215 | ~BUF2_REG_5__SCAN_IN;
  assign n33601 = ~n33651 | ~P2_DATAO_REG_5__SCAN_IN;
  assign U256 = ~n33602 | ~n33601;
  assign n33604 = ~U215 | ~BUF2_REG_6__SCAN_IN;
  assign n33603 = ~n33651 | ~P2_DATAO_REG_6__SCAN_IN;
  assign U257 = ~n33604 | ~n33603;
  assign n33606 = ~U215 | ~BUF2_REG_7__SCAN_IN;
  assign n33605 = ~n33651 | ~P2_DATAO_REG_7__SCAN_IN;
  assign U258 = ~n33606 | ~n33605;
  assign n33608 = ~U215 | ~BUF2_REG_8__SCAN_IN;
  assign n33607 = ~n33651 | ~P2_DATAO_REG_8__SCAN_IN;
  assign U259 = ~n33608 | ~n33607;
  assign n33610 = ~U215 | ~BUF2_REG_9__SCAN_IN;
  assign n33609 = ~n33651 | ~P2_DATAO_REG_9__SCAN_IN;
  assign U260 = ~n33610 | ~n33609;
  assign n33612 = ~U215 | ~BUF2_REG_10__SCAN_IN;
  assign n33611 = ~n33651 | ~P2_DATAO_REG_10__SCAN_IN;
  assign U261 = ~n33612 | ~n33611;
  assign n33614 = ~U215 | ~BUF2_REG_11__SCAN_IN;
  assign n33613 = ~n33651 | ~P2_DATAO_REG_11__SCAN_IN;
  assign U262 = ~n33614 | ~n33613;
  assign n33616 = ~U215 | ~BUF2_REG_12__SCAN_IN;
  assign n33615 = ~n33651 | ~P2_DATAO_REG_12__SCAN_IN;
  assign U263 = ~n33616 | ~n33615;
  assign n33618 = ~U215 | ~BUF2_REG_13__SCAN_IN;
  assign n33617 = ~n33651 | ~P2_DATAO_REG_13__SCAN_IN;
  assign U264 = ~n33618 | ~n33617;
  assign n33620 = ~U215 | ~BUF2_REG_14__SCAN_IN;
  assign n33619 = ~n33651 | ~P2_DATAO_REG_14__SCAN_IN;
  assign U265 = ~n33620 | ~n33619;
  assign n33622 = ~U215 | ~BUF2_REG_15__SCAN_IN;
  assign n33621 = ~n33651 | ~P2_DATAO_REG_15__SCAN_IN;
  assign U266 = ~n33622 | ~n33621;
  assign n33624 = ~U215 | ~BUF2_REG_16__SCAN_IN;
  assign n33623 = ~n33651 | ~P2_DATAO_REG_16__SCAN_IN;
  assign U267 = ~n33624 | ~n33623;
  assign n33626 = ~U215 | ~BUF2_REG_17__SCAN_IN;
  assign n33625 = ~n33651 | ~P2_DATAO_REG_17__SCAN_IN;
  assign U268 = ~n33626 | ~n33625;
  assign n33628 = ~U215 | ~BUF2_REG_18__SCAN_IN;
  assign n33627 = ~n33651 | ~P2_DATAO_REG_18__SCAN_IN;
  assign U269 = ~n33628 | ~n33627;
  assign n33630 = ~U215 | ~BUF2_REG_19__SCAN_IN;
  assign n33629 = ~n33651 | ~P2_DATAO_REG_19__SCAN_IN;
  assign U270 = ~n33630 | ~n33629;
  assign n33632 = ~U215 | ~BUF2_REG_20__SCAN_IN;
  assign n33631 = ~n33651 | ~P2_DATAO_REG_20__SCAN_IN;
  assign U271 = ~n33632 | ~n33631;
  assign n33634 = ~U215 | ~BUF2_REG_21__SCAN_IN;
  assign n33633 = ~n33651 | ~P2_DATAO_REG_21__SCAN_IN;
  assign U272 = ~n33634 | ~n33633;
  assign n33636 = ~U215 | ~BUF2_REG_22__SCAN_IN;
  assign n33635 = ~n33651 | ~P2_DATAO_REG_22__SCAN_IN;
  assign U273 = ~n33636 | ~n33635;
  assign n33638 = ~U215 | ~BUF2_REG_23__SCAN_IN;
  assign n33637 = ~n33651 | ~P2_DATAO_REG_23__SCAN_IN;
  assign U274 = ~n33638 | ~n33637;
  assign n33640 = ~U215 | ~BUF2_REG_24__SCAN_IN;
  assign n33639 = ~n33651 | ~P2_DATAO_REG_24__SCAN_IN;
  assign U275 = ~n33640 | ~n33639;
  assign n33642 = ~U215 | ~BUF2_REG_25__SCAN_IN;
  assign n33641 = ~n33651 | ~P2_DATAO_REG_25__SCAN_IN;
  assign U276 = ~n33642 | ~n33641;
  assign n33644 = ~U215 | ~BUF2_REG_26__SCAN_IN;
  assign n33643 = ~n33651 | ~P2_DATAO_REG_26__SCAN_IN;
  assign U277 = ~n33644 | ~n33643;
  assign n33646 = ~U215 | ~BUF2_REG_27__SCAN_IN;
  assign n33645 = ~n33651 | ~P2_DATAO_REG_27__SCAN_IN;
  assign U278 = ~n33646 | ~n33645;
  assign n33648 = ~U215 | ~BUF2_REG_28__SCAN_IN;
  assign n33647 = ~n33651 | ~P2_DATAO_REG_28__SCAN_IN;
  assign U279 = ~n33648 | ~n33647;
  assign n33650 = ~U215 | ~BUF2_REG_29__SCAN_IN;
  assign n33649 = ~n33651 | ~P2_DATAO_REG_29__SCAN_IN;
  assign U280 = ~n33650 | ~n33649;
  assign n33653 = ~U215 | ~BUF2_REG_30__SCAN_IN;
  assign n33652 = ~n33651 | ~P2_DATAO_REG_30__SCAN_IN;
  assign U281 = ~n33653 | ~n33652;
  assign n33655 = ~U215 | ~BUF2_REG_31__SCAN_IN;
  assign n33654 = ~n33651 | ~P2_DATAO_REG_31__SCAN_IN;
  assign U282 = ~n33655 | ~n33654;
  assign n33658 = ~P1_DATAO_REG_30__SCAN_IN | ~n33656;
  assign n33657 = ~P2_DATAO_REG_30__SCAN_IN | ~n39977;
  assign n33661 = ~n33658 | ~n33657;
  assign n33700 = ~n33661 & ~n33660;
  assign n33719 = ~n33722;
  assign n33663 = ~n33719 | ~P2_ADDRESS_REG_9__SCAN_IN;
  assign n33662 = ~n33722 | ~P3_ADDRESS_REG_9__SCAN_IN;
  assign U347 = ~n33663 | ~n33662;
  assign n33665 = ~n33719 | ~P2_ADDRESS_REG_8__SCAN_IN;
  assign n33664 = ~n33722 | ~P3_ADDRESS_REG_8__SCAN_IN;
  assign U348 = ~n33665 | ~n33664;
  assign n33667 = ~n33719 | ~P2_ADDRESS_REG_7__SCAN_IN;
  assign n33666 = ~n33722 | ~P3_ADDRESS_REG_7__SCAN_IN;
  assign U349 = ~n33667 | ~n33666;
  assign n33669 = ~n33719 | ~P2_ADDRESS_REG_6__SCAN_IN;
  assign n33668 = ~n33722 | ~P3_ADDRESS_REG_6__SCAN_IN;
  assign U350 = ~n33669 | ~n33668;
  assign n33671 = ~n33719 | ~P2_ADDRESS_REG_5__SCAN_IN;
  assign n33670 = ~n33722 | ~P3_ADDRESS_REG_5__SCAN_IN;
  assign U351 = ~n33671 | ~n33670;
  assign n33673 = ~n33719 | ~P2_ADDRESS_REG_4__SCAN_IN;
  assign n33672 = ~n33722 | ~P3_ADDRESS_REG_4__SCAN_IN;
  assign U352 = ~n33673 | ~n33672;
  assign n33675 = ~n33719 | ~P2_ADDRESS_REG_3__SCAN_IN;
  assign n33674 = ~n33722 | ~P3_ADDRESS_REG_3__SCAN_IN;
  assign U353 = ~n33675 | ~n33674;
  assign n33677 = ~n33719 | ~P2_ADDRESS_REG_2__SCAN_IN;
  assign n33676 = ~n33722 | ~P3_ADDRESS_REG_2__SCAN_IN;
  assign U354 = ~n33677 | ~n33676;
  assign n33679 = ~n33719 | ~P2_ADDRESS_REG_29__SCAN_IN;
  assign n33678 = ~n33722 | ~P3_ADDRESS_REG_29__SCAN_IN;
  assign U355 = ~n33679 | ~n33678;
  assign n33681 = ~n33719 | ~P2_ADDRESS_REG_28__SCAN_IN;
  assign n33680 = ~n33700 | ~P3_ADDRESS_REG_28__SCAN_IN;
  assign U356 = ~n33681 | ~n33680;
  assign n33683 = ~n33719 | ~P2_ADDRESS_REG_27__SCAN_IN;
  assign n33682 = ~n33700 | ~P3_ADDRESS_REG_27__SCAN_IN;
  assign U357 = ~n33683 | ~n33682;
  assign n33685 = ~n33719 | ~P2_ADDRESS_REG_26__SCAN_IN;
  assign n33684 = ~n33700 | ~P3_ADDRESS_REG_26__SCAN_IN;
  assign U358 = ~n33685 | ~n33684;
  assign n33687 = ~n33719 | ~P2_ADDRESS_REG_25__SCAN_IN;
  assign n33686 = ~n33700 | ~P3_ADDRESS_REG_25__SCAN_IN;
  assign U359 = ~n33687 | ~n33686;
  assign n33689 = ~n33719 | ~P2_ADDRESS_REG_24__SCAN_IN;
  assign n33688 = ~n33700 | ~P3_ADDRESS_REG_24__SCAN_IN;
  assign U360 = ~n33689 | ~n33688;
  assign n33691 = ~n33719 | ~P2_ADDRESS_REG_23__SCAN_IN;
  assign n33690 = ~n33700 | ~P3_ADDRESS_REG_23__SCAN_IN;
  assign U361 = ~n33691 | ~n33690;
  assign n33693 = ~n33719 | ~P2_ADDRESS_REG_22__SCAN_IN;
  assign n33692 = ~n33700 | ~P3_ADDRESS_REG_22__SCAN_IN;
  assign U362 = ~n33693 | ~n33692;
  assign n33695 = ~n33719 | ~P2_ADDRESS_REG_21__SCAN_IN;
  assign n33694 = ~n33700 | ~P3_ADDRESS_REG_21__SCAN_IN;
  assign U363 = ~n33695 | ~n33694;
  assign n33697 = ~n33719 | ~P2_ADDRESS_REG_20__SCAN_IN;
  assign n33696 = ~n33700 | ~P3_ADDRESS_REG_20__SCAN_IN;
  assign U364 = ~n33697 | ~n33696;
  assign n33699 = ~n33719 | ~P2_ADDRESS_REG_1__SCAN_IN;
  assign n33698 = ~n33700 | ~P3_ADDRESS_REG_1__SCAN_IN;
  assign U365 = ~n33699 | ~n33698;
  assign n33702 = ~n33719 | ~P2_ADDRESS_REG_19__SCAN_IN;
  assign n33701 = ~n33700 | ~P3_ADDRESS_REG_19__SCAN_IN;
  assign U366 = ~n33702 | ~n33701;
  assign n33704 = ~n33719 | ~P2_ADDRESS_REG_18__SCAN_IN;
  assign n33703 = ~n33722 | ~P3_ADDRESS_REG_18__SCAN_IN;
  assign U367 = ~n33704 | ~n33703;
  assign n33706 = ~n33719 | ~P2_ADDRESS_REG_17__SCAN_IN;
  assign n33705 = ~n33722 | ~P3_ADDRESS_REG_17__SCAN_IN;
  assign U368 = ~n33706 | ~n33705;
  assign n33708 = ~n33719 | ~P2_ADDRESS_REG_16__SCAN_IN;
  assign n33707 = ~n33722 | ~P3_ADDRESS_REG_16__SCAN_IN;
  assign U369 = ~n33708 | ~n33707;
  assign n33710 = ~n33719 | ~P2_ADDRESS_REG_15__SCAN_IN;
  assign n33709 = ~n33722 | ~P3_ADDRESS_REG_15__SCAN_IN;
  assign U370 = ~n33710 | ~n33709;
  assign n33712 = ~n33719 | ~P2_ADDRESS_REG_14__SCAN_IN;
  assign n33711 = ~n33722 | ~P3_ADDRESS_REG_14__SCAN_IN;
  assign U371 = ~n33712 | ~n33711;
  assign n33714 = ~n33719 | ~P2_ADDRESS_REG_13__SCAN_IN;
  assign n33713 = ~n33722 | ~P3_ADDRESS_REG_13__SCAN_IN;
  assign U372 = ~n33714 | ~n33713;
  assign n33716 = ~n33719 | ~P2_ADDRESS_REG_12__SCAN_IN;
  assign n33715 = ~n33722 | ~P3_ADDRESS_REG_12__SCAN_IN;
  assign U373 = ~n33716 | ~n33715;
  assign n33718 = ~n33719 | ~P2_ADDRESS_REG_11__SCAN_IN;
  assign n33717 = ~n33722 | ~P3_ADDRESS_REG_11__SCAN_IN;
  assign U374 = ~n33718 | ~n33717;
  assign n33721 = ~n33719 | ~P2_ADDRESS_REG_10__SCAN_IN;
  assign n33720 = ~n33722 | ~P3_ADDRESS_REG_10__SCAN_IN;
  assign U375 = ~n33721 | ~n33720;
  assign n33724 = ~n33719 | ~P2_ADDRESS_REG_0__SCAN_IN;
  assign n33723 = ~n33722 | ~P3_ADDRESS_REG_0__SCAN_IN;
  assign U376 = ~n33724 | ~n33723;
  assign n33727 = ~n38854 | ~n38831;
  assign n38860 = ~P3_STATE_REG_2__SCAN_IN;
  assign n33725 = ~n38854 & ~n38831;
  assign n33726 = ~n38860 | ~n33725;
  assign n39019 = ~n33727 | ~n33726;
  assign n33728 = ~P3_STATE_REG_0__SCAN_IN | ~P3_ADS_N_REG_SCAN_IN;
  assign P3_U2633 = ~n22822 | ~n33728;
  assign n39130 = ~n33729 & ~P3_STATE2_REG_1__SCAN_IN;
  assign n33732 = ~P3_STATE2_REG_0__SCAN_IN | ~n39130;
  assign n33730 = ~n33747 | ~n35945;
  assign n33731 = ~P3_CODEFETCH_REG_SCAN_IN | ~n33730;
  assign P3_U2634 = ~n33732 | ~n33731;
  assign n33733 = ~P3_STATE_REG_0__SCAN_IN & ~P3_STATE_REG_2__SCAN_IN;
  assign n33734 = ~P3_D_C_N_REG_SCAN_IN & ~n33733;
  assign n33736 = ~n39126 & ~n33734;
  assign n33735 = ~P3_CODEFETCH_REG_SCAN_IN & ~n39097;
  assign P3_U2635 = n33736 | n33735;
  assign n33738 = n33737 | BS16;
  assign n39023 = ~n39019 | ~n33738;
  assign n33739 = ~P3_STATEBS16_REG_SCAN_IN | ~n22822;
  assign P3_U2636 = ~n39023 | ~n33739;
  assign n38804 = ~n39114;
  assign n33789 = ~n35811 & ~n35948;
  assign n33741 = ~n33789 & ~n33740;
  assign n33743 = ~n33742 & ~n33741;
  assign n33745 = ~n38804 & ~n33743;
  assign n33744 = ~n38681;
  assign n33746 = ~n33745 & ~n33744;
  assign n38670 = ~n33747 | ~n33746;
  assign n39101 = ~n39105 | ~n38670;
  assign n33748 = ~P3_FLUSH_REG_SCAN_IN | ~n39101;
  assign P3_U2637 = ~n33749 | ~n33748;
  assign n33751 = ~P3_DATAWIDTH_REG_12__SCAN_IN & ~P3_DATAWIDTH_REG_13__SCAN_IN;
  assign n33750 = ~P3_DATAWIDTH_REG_14__SCAN_IN & ~P3_DATAWIDTH_REG_15__SCAN_IN;
  assign n33755 = ~n33751 | ~n33750;
  assign n33753 = ~P3_DATAWIDTH_REG_8__SCAN_IN & ~P3_DATAWIDTH_REG_9__SCAN_IN;
  assign n33752 = ~P3_DATAWIDTH_REG_10__SCAN_IN & ~P3_DATAWIDTH_REG_11__SCAN_IN;
  assign n33754 = ~n33753 | ~n33752;
  assign n33779 = ~n33755 & ~n33754;
  assign n33757 = ~P3_DATAWIDTH_REG_4__SCAN_IN & ~P3_DATAWIDTH_REG_5__SCAN_IN;
  assign n33756 = ~P3_DATAWIDTH_REG_6__SCAN_IN & ~P3_DATAWIDTH_REG_7__SCAN_IN;
  assign n33759 = ~n33757 | ~n33756;
  assign n33758 = P3_DATAWIDTH_REG_0__SCAN_IN & P3_DATAWIDTH_REG_1__SCAN_IN;
  assign n33761 = ~n33759 & ~n33758;
  assign n33760 = ~P3_DATAWIDTH_REG_2__SCAN_IN & ~P3_DATAWIDTH_REG_3__SCAN_IN;
  assign n33777 = ~n33761 | ~n33760;
  assign n33763 = ~P3_DATAWIDTH_REG_28__SCAN_IN & ~P3_DATAWIDTH_REG_29__SCAN_IN;
  assign n33762 = ~P3_DATAWIDTH_REG_30__SCAN_IN & ~P3_DATAWIDTH_REG_31__SCAN_IN;
  assign n33767 = ~n33763 | ~n33762;
  assign n33765 = ~P3_DATAWIDTH_REG_24__SCAN_IN & ~P3_DATAWIDTH_REG_25__SCAN_IN;
  assign n33764 = ~P3_DATAWIDTH_REG_26__SCAN_IN & ~P3_DATAWIDTH_REG_27__SCAN_IN;
  assign n33766 = ~n33765 | ~n33764;
  assign n33775 = ~n33767 & ~n33766;
  assign n33769 = ~P3_DATAWIDTH_REG_20__SCAN_IN & ~P3_DATAWIDTH_REG_21__SCAN_IN;
  assign n33768 = ~P3_DATAWIDTH_REG_22__SCAN_IN & ~P3_DATAWIDTH_REG_23__SCAN_IN;
  assign n33773 = ~n33769 | ~n33768;
  assign n33771 = ~P3_DATAWIDTH_REG_16__SCAN_IN & ~P3_DATAWIDTH_REG_17__SCAN_IN;
  assign n33770 = ~P3_DATAWIDTH_REG_18__SCAN_IN & ~P3_DATAWIDTH_REG_19__SCAN_IN;
  assign n33772 = ~n33771 | ~n33770;
  assign n33774 = ~n33773 & ~n33772;
  assign n33776 = ~n33775 | ~n33774;
  assign n33778 = ~n33777 & ~n33776;
  assign n39092 = ~n33779 | ~n33778;
  assign n33783 = ~P3_BYTEENABLE_REG_1__SCAN_IN | ~n39092;
  assign n39083 = ~P3_REIP_REG_0__SCAN_IN;
  assign n39082 = ~P3_DATAWIDTH_REG_0__SCAN_IN;
  assign n33780 = ~n39083 | ~n39082;
  assign n33784 = ~P3_DATAWIDTH_REG_1__SCAN_IN & ~n33780;
  assign n33781 = ~P3_REIP_REG_1__SCAN_IN & ~n33784;
  assign n33782 = n39092 | n33781;
  assign P3_U2638 = ~n33783 | ~n33782;
  assign n33787 = ~P3_BYTEENABLE_REG_3__SCAN_IN | ~n39092;
  assign n39081 = ~P3_REIP_REG_1__SCAN_IN & ~P3_DATAWIDTH_REG_1__SCAN_IN;
  assign n33785 = ~n33784 & ~n39081;
  assign n33786 = n39092 | n33785;
  assign P3_U2639 = ~n33787 | ~n33786;
  assign n39006 = ~P3_REIP_REG_31__SCAN_IN;
  assign n33847 = ~n36112 | ~n39114;
  assign n34005 = ~P3_REIP_REG_21__SCAN_IN | ~P3_REIP_REG_20__SCAN_IN;
  assign n38950 = ~P3_REIP_REG_19__SCAN_IN;
  assign n38940 = ~P3_REIP_REG_17__SCAN_IN;
  assign n38930 = ~P3_REIP_REG_15__SCAN_IN;
  assign n38920 = ~P3_REIP_REG_13__SCAN_IN;
  assign n38910 = ~P3_REIP_REG_11__SCAN_IN;
  assign n38900 = ~P3_REIP_REG_9__SCAN_IN;
  assign n38880 = ~P3_REIP_REG_5__SCAN_IN;
  assign n39084 = ~P3_REIP_REG_1__SCAN_IN;
  assign n33790 = ~P3_REIP_REG_3__SCAN_IN | ~P3_REIP_REG_2__SCAN_IN;
  assign n34369 = ~n39084 & ~n33790;
  assign n34349 = ~P3_REIP_REG_4__SCAN_IN | ~n34369;
  assign n34325 = ~n38880 & ~n34349;
  assign n34305 = ~P3_REIP_REG_6__SCAN_IN | ~n34325;
  assign n34285 = ~n38890 & ~n34305;
  assign n34243 = ~P3_REIP_REG_8__SCAN_IN | ~n34285;
  assign n34231 = ~n38900 & ~n34243;
  assign n34219 = ~P3_REIP_REG_10__SCAN_IN | ~n34231;
  assign n34191 = ~n38910 & ~n34219;
  assign n34173 = ~P3_REIP_REG_12__SCAN_IN | ~n34191;
  assign n34145 = ~n38920 & ~n34173;
  assign n34127 = ~P3_REIP_REG_14__SCAN_IN | ~n34145;
  assign n34112 = ~n38930 & ~n34127;
  assign n34090 = ~P3_REIP_REG_16__SCAN_IN | ~n34112;
  assign n34077 = ~n38940 & ~n34090;
  assign n34058 = ~P3_REIP_REG_18__SCAN_IN | ~n34077;
  assign n34004 = ~n38950 & ~n34058;
  assign n33791 = ~P3_REIP_REG_22__SCAN_IN | ~n34004;
  assign n33945 = ~n34005 & ~n33791;
  assign n33892 = ~P3_REIP_REG_24__SCAN_IN | ~P3_REIP_REG_23__SCAN_IN;
  assign n33894 = ~P3_REIP_REG_26__SCAN_IN | ~P3_REIP_REG_25__SCAN_IN;
  assign n33792 = ~n33892 & ~n33894;
  assign n33915 = ~n33945 | ~n33792;
  assign n33793 = ~P3_REIP_REG_28__SCAN_IN | ~P3_REIP_REG_27__SCAN_IN;
  assign n33872 = ~n33915 & ~n33793;
  assign n33797 = ~P3_REIP_REG_29__SCAN_IN | ~n33872;
  assign n33840 = n34405 | n33797;
  assign n33865 = ~P3_REIP_REG_30__SCAN_IN & ~n33840;
  assign n33795 = ~n39132 | ~n37197;
  assign n38818 = ~n33794 & ~n38810;
  assign n38808 = ~n38815 | ~n38476;
  assign n33798 = ~n34371 & ~n33797;
  assign n33869 = ~n34468 & ~n33798;
  assign n33799 = ~n33865 & ~n33869;
  assign n33846 = ~n39006 & ~n33799;
  assign n33806 = n34460 | n36107;
  assign n33800 = ~n36109 | ~n33806;
  assign n36106 = ~n33801 | ~n33800;
  assign n33907 = ~n36106;
  assign n36147 = ~P3_PHYADDRPOINTER_REG_27__SCAN_IN;
  assign n36184 = ~n33802;
  assign n33810 = ~n34460 & ~n36184;
  assign n36111 = ~n33803 | ~n33810;
  assign n33804 = n36166 | n36111;
  assign n33805 = ~n36147 | ~n33804;
  assign n36148 = ~n33806 | ~n33805;
  assign n33833 = ~n36148;
  assign n33807 = ~P3_PHYADDRPOINTER_REG_24__SCAN_IN | ~n33810;
  assign n33808 = ~n36183 | ~n33807;
  assign n36180 = ~n36111 | ~n33808;
  assign n33832 = ~n36180;
  assign n36209 = n33810 ^ P3_PHYADDRPOINTER_REG_24__SCAN_IN;
  assign n33814 = P3_PHYADDRPOINTER_REG_1__SCAN_IN & n36260;
  assign n36239 = ~P3_PHYADDRPOINTER_REG_22__SCAN_IN | ~n33814;
  assign n33809 = n36229 & n36239;
  assign n36234 = ~n33810 & ~n33809;
  assign n36272 = P3_PHYADDRPOINTER_REG_22__SCAN_IN ^ n33814;
  assign n33819 = ~n34460 & ~n36347;
  assign n36345 = ~n33819;
  assign n36263 = ~n33811 & ~n36345;
  assign n33812 = P3_PHYADDRPOINTER_REG_20__SCAN_IN & n36263;
  assign n33813 = ~P3_PHYADDRPOINTER_REG_21__SCAN_IN & ~n33812;
  assign n36291 = ~n33814 & ~n33813;
  assign n36311 = n23552 ^ n36263;
  assign n33827 = ~n36311;
  assign n36364 = ~P3_PHYADDRPOINTER_REG_18__SCAN_IN;
  assign n33815 = ~n36364 & ~n36345;
  assign n33816 = ~P3_PHYADDRPOINTER_REG_19__SCAN_IN & ~n33815;
  assign n36342 = ~n36263 & ~n33816;
  assign n33825 = ~P3_PHYADDRPOINTER_REG_1__SCAN_IN | ~n36384;
  assign n33817 = ~n33825;
  assign n33818 = ~P3_PHYADDRPOINTER_REG_17__SCAN_IN & ~n33817;
  assign n36391 = ~n33819 & ~n33818;
  assign n36447 = ~P3_PHYADDRPOINTER_REG_15__SCAN_IN;
  assign n36455 = ~P3_PHYADDRPOINTER_REG_14__SCAN_IN;
  assign n33821 = ~n33820;
  assign n34298 = ~P3_PHYADDRPOINTER_REG_1__SCAN_IN | ~n36536;
  assign n36477 = ~n33821 & ~n34298;
  assign n34179 = ~n33822 | ~n36477;
  assign n36410 = ~n36455 & ~n34179;
  assign n36747 = ~P3_PHYADDRPOINTER_REG_0__SCAN_IN;
  assign n34138 = ~n36410 | ~n36747;
  assign n34107 = ~n36447 & ~n34138;
  assign n36412 = ~P3_PHYADDRPOINTER_REG_16__SCAN_IN;
  assign n33823 = ~P3_PHYADDRPOINTER_REG_15__SCAN_IN | ~n36410;
  assign n33824 = ~n36412 | ~n33823;
  assign n36404 = ~n33825 | ~n33824;
  assign n34086 = ~n34107 | ~n36404;
  assign n34071 = ~n36391 & ~n34086;
  assign n36363 = ~n36364 ^ n36345;
  assign n34051 = ~n34071 | ~n36363;
  assign n33826 = ~n36342 & ~n34051;
  assign n34030 = ~n34320 & ~n33826;
  assign n33828 = ~n33827 & ~n34030;
  assign n33829 = ~n36291 & ~n34024;
  assign n33956 = ~n33831 & ~n34376;
  assign n33834 = ~n33833 & ~n22989;
  assign n33906 = ~n33834 & ~n34376;
  assign n33835 = ~n33863 & ~n33862;
  assign n34463 = ~n38818;
  assign n34421 = ~n34320 & ~n34463;
  assign n33844 = ~n33835 | ~n34421;
  assign n33850 = ~P3_EBX_REG_31__SCAN_IN | ~n35948;
  assign n33836 = ~n33848 | ~n33850;
  assign n34445 = ~n38796 & ~n33836;
  assign n33838 = ~n34445 | ~P3_EBX_REG_31__SCAN_IN;
  assign n33837 = ~n34384 | ~P3_PHYADDRPOINTER_REG_31__SCAN_IN;
  assign n33842 = ~n33838 | ~n33837;
  assign n33839 = ~P3_REIP_REG_30__SCAN_IN | ~n39006;
  assign n33841 = ~n33840 & ~n33839;
  assign n33843 = ~n33842 & ~n33841;
  assign n33845 = ~n33844 | ~n33843;
  assign n33853 = ~n33846 & ~n33845;
  assign n34484 = ~P3_EBX_REG_2__SCAN_IN;
  assign n34401 = ~n34447 | ~n34484;
  assign n34389 = ~P3_EBX_REG_3__SCAN_IN & ~n34401;
  assign n34486 = ~P3_EBX_REG_4__SCAN_IN;
  assign n34352 = ~n34389 | ~n34486;
  assign n34317 = ~P3_EBX_REG_5__SCAN_IN & ~n34352;
  assign n34304 = ~n34317 | ~n35447;
  assign n34276 = ~P3_EBX_REG_7__SCAN_IN & ~n34304;
  assign n34279 = ~P3_EBX_REG_8__SCAN_IN;
  assign n34251 = ~n34276 | ~n34279;
  assign n34227 = ~P3_EBX_REG_9__SCAN_IN & ~n34251;
  assign n34217 = ~n34227 | ~n35353;
  assign n34189 = ~P3_EBX_REG_11__SCAN_IN & ~n34217;
  assign n34167 = ~n34189 | ~n35273;
  assign n34154 = ~P3_EBX_REG_13__SCAN_IN & ~n34167;
  assign n35190 = ~P3_EBX_REG_14__SCAN_IN;
  assign n34128 = ~n34154 | ~n35190;
  assign n35121 = ~P3_EBX_REG_16__SCAN_IN;
  assign n34093 = ~n34116 | ~n35121;
  assign n34074 = ~P3_EBX_REG_17__SCAN_IN & ~n34093;
  assign n34047 = ~n34074 | ~n34492;
  assign n34035 = ~P3_EBX_REG_19__SCAN_IN & ~n34047;
  assign n34493 = ~P3_EBX_REG_20__SCAN_IN;
  assign n34021 = ~n34035 | ~n34493;
  assign n34893 = ~P3_EBX_REG_22__SCAN_IN;
  assign n33980 = ~n34002 | ~n34893;
  assign n33963 = ~P3_EBX_REG_23__SCAN_IN & ~n33980;
  assign n34494 = ~P3_EBX_REG_24__SCAN_IN;
  assign n33948 = ~n33963 | ~n34494;
  assign n33930 = ~P3_EBX_REG_25__SCAN_IN & ~n33948;
  assign n34806 = ~P3_EBX_REG_26__SCAN_IN;
  assign n33912 = ~n33930 | ~n34806;
  assign n33900 = ~P3_EBX_REG_27__SCAN_IN & ~n33912;
  assign n33899 = ~P3_EBX_REG_28__SCAN_IN;
  assign n33898 = ~n33900 | ~n33899;
  assign n33854 = ~P3_EBX_REG_29__SCAN_IN & ~n33898;
  assign n33849 = ~n33848 | ~n33847;
  assign n33851 = ~P3_EBX_REG_30__SCAN_IN & ~n34470;
  assign n33852 = ~n33854 | ~n33851;
  assign P3_U2640 = ~n33853 | ~n33852;
  assign n34507 = ~P3_EBX_REG_30__SCAN_IN;
  assign n33855 = n34507 ^ n33854;
  assign n33857 = ~n33855 | ~n34448;
  assign n33856 = ~P3_EBX_REG_30__SCAN_IN | ~n34445;
  assign n33861 = ~n33857 | ~n33856;
  assign n33859 = ~n33869 | ~P3_REIP_REG_30__SCAN_IN;
  assign n33858 = ~n34384 | ~P3_PHYADDRPOINTER_REG_30__SCAN_IN;
  assign n33860 = ~n33859 | ~n33858;
  assign n33868 = ~n33861 & ~n33860;
  assign n33864 = ~n33863 ^ n33862;
  assign n33866 = ~n34463 & ~n33864;
  assign n33867 = ~n33866 & ~n33865;
  assign P3_U2641 = ~n33868 | ~n33867;
  assign n33871 = ~n33869 | ~P3_REIP_REG_29__SCAN_IN;
  assign n33870 = ~n34384 | ~P3_PHYADDRPOINTER_REG_29__SCAN_IN;
  assign n33875 = ~n33871 | ~n33870;
  assign n33873 = ~n33872 | ~n34430;
  assign n33874 = ~P3_REIP_REG_29__SCAN_IN & ~n33873;
  assign n33885 = ~n33875 & ~n33874;
  assign n33878 = ~P3_EBX_REG_29__SCAN_IN | ~n34445;
  assign n33876 = P3_EBX_REG_29__SCAN_IN ^ n33898;
  assign n33877 = ~n33876 | ~n34448;
  assign n33883 = ~n33878 | ~n33877;
  assign n33881 = ~n33880 ^ n33879;
  assign n33882 = ~n34463 & ~n33881;
  assign n33884 = ~n33883 & ~n33882;
  assign P3_U2642 = ~n33885 | ~n33884;
  assign n33886 = ~n34371 & ~n33915;
  assign n33940 = ~n34468 & ~n33886;
  assign n33917 = ~P3_REIP_REG_27__SCAN_IN & ~n34405;
  assign n33887 = ~n33940 & ~n33917;
  assign n33891 = ~n33887 & ~n33447;
  assign n33889 = ~P3_EBX_REG_28__SCAN_IN | ~n34445;
  assign n33888 = ~n34384 | ~P3_PHYADDRPOINTER_REG_28__SCAN_IN;
  assign n33890 = ~n33889 | ~n33888;
  assign n33897 = ~n33891 & ~n33890;
  assign n33986 = ~n34430 | ~n33945;
  assign n33953 = ~n33892 & ~n33986;
  assign n33893 = ~P3_REIP_REG_27__SCAN_IN | ~n33953;
  assign n33895 = ~n33894 & ~n33893;
  assign n33896 = ~n33895 | ~n33447;
  assign n33904 = ~n33897 | ~n33896;
  assign n33902 = ~n34448 | ~n33898;
  assign n33901 = ~n33900 & ~n33899;
  assign n33903 = ~n33902 & ~n33901;
  assign n33911 = ~n33904 & ~n33903;
  assign n33909 = ~n33905 & ~n34463;
  assign n33908 = ~n33907 | ~n33906;
  assign n33910 = ~n33909 | ~n33908;
  assign P3_U2643 = ~n33911 | ~n33910;
  assign n34827 = ~P3_EBX_REG_27__SCAN_IN;
  assign n33913 = n34827 ^ n33912;
  assign n33925 = ~n34470 & ~n33913;
  assign n33914 = n36148 ^ n22989;
  assign n33921 = ~n34463 & ~n33914;
  assign n33916 = ~n33915;
  assign n33919 = ~n33917 | ~n33916;
  assign n33918 = ~P3_EBX_REG_27__SCAN_IN | ~n34445;
  assign n33920 = ~n33919 | ~n33918;
  assign n33923 = ~n33921 & ~n33920;
  assign n33922 = ~n34384 | ~P3_PHYADDRPOINTER_REG_27__SCAN_IN;
  assign n33924 = ~n33923 | ~n33922;
  assign n33927 = ~n33925 & ~n33924;
  assign n33926 = ~n33940 | ~P3_REIP_REG_27__SCAN_IN;
  assign P3_U2644 = ~n33927 | ~n33926;
  assign n33928 = ~P3_REIP_REG_25__SCAN_IN | ~n33953;
  assign n33939 = ~P3_REIP_REG_26__SCAN_IN & ~n33928;
  assign n33929 = n23066 ^ n22926;
  assign n33935 = ~n34463 & ~n33929;
  assign n33931 = n34806 ^ n33930;
  assign n33933 = ~n33931 | ~n34448;
  assign n33932 = ~P3_EBX_REG_26__SCAN_IN | ~n34445;
  assign n33934 = ~n33933 | ~n33932;
  assign n33937 = ~n33935 & ~n33934;
  assign n33936 = ~n34384 | ~P3_PHYADDRPOINTER_REG_26__SCAN_IN;
  assign n33938 = ~n33937 | ~n33936;
  assign n33942 = ~n33939 & ~n33938;
  assign n33941 = ~P3_REIP_REG_26__SCAN_IN | ~n33940;
  assign P3_U2645 = ~n33942 | ~n33941;
  assign n33965 = ~n34448 | ~n33948;
  assign n33944 = ~n33965 & ~P3_EBX_REG_25__SCAN_IN;
  assign n33943 = ~n36183 & ~n34459;
  assign n33961 = ~n33944 & ~n33943;
  assign n33970 = ~n33945 | ~P3_REIP_REG_23__SCAN_IN;
  assign n33946 = ~n34371 & ~n33970;
  assign n33987 = ~n34468 & ~n33946;
  assign n33972 = ~P3_REIP_REG_24__SCAN_IN & ~n34405;
  assign n33947 = ~n33987 & ~n33972;
  assign n38981 = ~P3_REIP_REG_25__SCAN_IN;
  assign n33952 = ~n33947 & ~n38981;
  assign n34805 = ~P3_EBX_REG_25__SCAN_IN;
  assign n33949 = ~n34470 & ~n33948;
  assign n33950 = ~n34445 & ~n33949;
  assign n33951 = ~n34805 & ~n33950;
  assign n33955 = ~n33952 & ~n33951;
  assign n33954 = ~n33953 | ~n38981;
  assign n33959 = ~n33955 | ~n33954;
  assign n33957 = n36180 ^ n33956;
  assign n33958 = ~n34463 & ~n33957;
  assign n33960 = ~n33959 & ~n33958;
  assign P3_U2646 = ~n33961 | ~n33960;
  assign n33962 = ~n36209 ^ n23038;
  assign n33976 = ~n34463 & ~n33962;
  assign n33964 = ~n33963 & ~n34494;
  assign n33969 = ~n33965 & ~n33964;
  assign n33967 = ~P3_EBX_REG_24__SCAN_IN | ~n34445;
  assign n33966 = ~n34384 | ~P3_PHYADDRPOINTER_REG_24__SCAN_IN;
  assign n33968 = ~n33967 | ~n33966;
  assign n33974 = ~n33969 & ~n33968;
  assign n33971 = ~n33970;
  assign n33973 = ~n33972 | ~n33971;
  assign n33975 = ~n33974 | ~n33973;
  assign n33978 = ~n33976 & ~n33975;
  assign n33977 = ~n33987 | ~P3_REIP_REG_24__SCAN_IN;
  assign P3_U2647 = ~n33978 | ~n33977;
  assign n33979 = ~n36234 ^ n23037;
  assign n33985 = ~n34463 & ~n33979;
  assign n34804 = ~P3_EBX_REG_23__SCAN_IN;
  assign n33981 = ~n34804 ^ n33980;
  assign n33983 = ~n34448 | ~n33981;
  assign n33982 = ~P3_PHYADDRPOINTER_REG_23__SCAN_IN | ~n34384;
  assign n33984 = ~n33983 | ~n33982;
  assign n33993 = ~n33985 & ~n33984;
  assign n33991 = ~n33986 & ~P3_REIP_REG_23__SCAN_IN;
  assign n33989 = ~n34445 | ~P3_EBX_REG_23__SCAN_IN;
  assign n33988 = ~P3_REIP_REG_23__SCAN_IN | ~n33987;
  assign n33990 = ~n33989 | ~n33988;
  assign n33992 = ~n33991 & ~n33990;
  assign P3_U2648 = ~n33993 | ~n33992;
  assign n33995 = ~P3_EBX_REG_22__SCAN_IN | ~n34445;
  assign n33994 = ~n34384 | ~P3_PHYADDRPOINTER_REG_22__SCAN_IN;
  assign n33998 = ~n33995 | ~n33994;
  assign n33997 = ~n34463 & ~n33996;
  assign n34012 = ~n33998 & ~n33997;
  assign n34014 = ~n34004 | ~P3_REIP_REG_20__SCAN_IN;
  assign n33999 = ~n34371 & ~n34014;
  assign n34044 = ~n34468 & ~n33999;
  assign n38960 = ~P3_REIP_REG_21__SCAN_IN;
  assign n34013 = ~n38960 | ~n34430;
  assign n34000 = ~n34013;
  assign n34001 = ~n34044 & ~n34000;
  assign n38965 = ~P3_REIP_REG_22__SCAN_IN;
  assign n34010 = ~n34001 & ~n38965;
  assign n34003 = n34893 ^ n34002;
  assign n34008 = ~n34003 | ~n34448;
  assign n34034 = ~n34430 | ~n34004;
  assign n34006 = ~n34005 & ~n34034;
  assign n34007 = ~n38965 | ~n34006;
  assign n34009 = ~n34008 | ~n34007;
  assign n34011 = ~n34010 & ~n34009;
  assign P3_U2649 = ~n34012 | ~n34011;
  assign n34020 = ~n34014 & ~n34013;
  assign n34037 = ~n34448 | ~n34021;
  assign n34016 = ~n34037 & ~P3_EBX_REG_21__SCAN_IN;
  assign n34015 = ~n36290 & ~n34459;
  assign n34018 = ~n34016 & ~n34015;
  assign n34017 = ~P3_REIP_REG_21__SCAN_IN | ~n34044;
  assign n34019 = ~n34018 | ~n34017;
  assign n34029 = ~n34020 & ~n34019;
  assign n34803 = ~P3_EBX_REG_21__SCAN_IN;
  assign n34022 = ~n34470 & ~n34021;
  assign n34023 = ~n34445 & ~n34022;
  assign n34027 = ~n34803 & ~n34023;
  assign n34025 = ~n36291 ^ n34024;
  assign n34026 = ~n34463 & ~n34025;
  assign n34028 = ~n34027 & ~n34026;
  assign P3_U2650 = ~n34029 | ~n34028;
  assign n34031 = n36311 ^ n34030;
  assign n34043 = ~n34463 & ~n34031;
  assign n34033 = ~n34469 & ~n34493;
  assign n34032 = ~n23552 & ~n34459;
  assign n34041 = ~n34033 & ~n34032;
  assign n34039 = ~P3_REIP_REG_20__SCAN_IN & ~n34034;
  assign n34036 = ~n34035 & ~n34493;
  assign n34038 = ~n34037 & ~n34036;
  assign n34040 = ~n34039 & ~n34038;
  assign n34042 = ~n34041 | ~n34040;
  assign n34046 = ~n34043 & ~n34042;
  assign n34045 = ~n34044 | ~P3_REIP_REG_20__SCAN_IN;
  assign P3_U2651 = ~n34046 | ~n34045;
  assign n34050 = ~P3_EBX_REG_19__SCAN_IN | ~n34445;
  assign n34048 = P3_EBX_REG_19__SCAN_IN ^ n34047;
  assign n34049 = ~n34048 | ~n34448;
  assign n34055 = ~n34050 | ~n34049;
  assign n34052 = ~n34425 | ~n34051;
  assign n34053 = n36342 ^ n34052;
  assign n34054 = ~n34463 & ~n34053;
  assign n34065 = ~n34055 & ~n34054;
  assign n34076 = ~P3_REIP_REG_18__SCAN_IN & ~n34405;
  assign n34089 = n34405 | n34077;
  assign n34102 = ~n34478 | ~n34089;
  assign n34056 = ~n34076 & ~n34102;
  assign n34063 = ~n38950 & ~n34056;
  assign n34057 = ~n34430 | ~n38950;
  assign n34059 = ~n34058 & ~n34057;
  assign n34061 = ~n22843 & ~n34059;
  assign n34060 = ~P3_PHYADDRPOINTER_REG_19__SCAN_IN | ~n34384;
  assign n34062 = ~n34061 | ~n34060;
  assign n34064 = ~n34063 & ~n34062;
  assign P3_U2652 = ~n34065 | ~n34064;
  assign n34067 = ~n34469 & ~n34492;
  assign n34066 = ~n36364 & ~n34459;
  assign n34069 = ~n34067 & ~n34066;
  assign n34068 = ~P3_REIP_REG_18__SCAN_IN | ~n34102;
  assign n34070 = ~n34069 | ~n34068;
  assign n34083 = ~n22843 & ~n34070;
  assign n34072 = ~n34071 & ~n34376;
  assign n34073 = n34072 ^ n36363;
  assign n34081 = ~n34463 & ~n34073;
  assign n34075 = n34074 ^ n34492;
  assign n34079 = ~n34075 | ~n34448;
  assign n34078 = ~n34077 | ~n34076;
  assign n34080 = ~n34079 | ~n34078;
  assign n34082 = ~n34081 & ~n34080;
  assign P3_U2653 = ~n34083 | ~n34082;
  assign n35078 = ~P3_EBX_REG_17__SCAN_IN;
  assign n34084 = ~n34470 & ~n34093;
  assign n34085 = ~n34445 & ~n34084;
  assign n34101 = ~n35078 & ~n34085;
  assign n34087 = ~n34425 | ~n34086;
  assign n34088 = n36391 ^ n34087;
  assign n34097 = ~n34463 & ~n34088;
  assign n34091 = ~n34090 & ~n34089;
  assign n34095 = ~n22843 & ~n34091;
  assign n34092 = ~P3_EBX_REG_17__SCAN_IN & ~n34470;
  assign n34094 = ~n34093 | ~n34092;
  assign n34096 = ~n34095 | ~n34094;
  assign n34099 = ~n34097 & ~n34096;
  assign n34098 = ~n34384 | ~P3_PHYADDRPOINTER_REG_17__SCAN_IN;
  assign n34100 = ~n34099 | ~n34098;
  assign n34104 = ~n34101 & ~n34100;
  assign n34103 = ~P3_REIP_REG_17__SCAN_IN | ~n34102;
  assign P3_U2654 = ~n34104 | ~n34103;
  assign n34126 = ~n34430 | ~n38930;
  assign n34105 = n34127 & n34430;
  assign n34147 = ~n34371 & ~n34105;
  assign n34106 = ~n34126 | ~n34147;
  assign n34125 = ~n34106 | ~P3_REIP_REG_16__SCAN_IN;
  assign n34108 = ~n34107 & ~n34376;
  assign n34109 = n34108 ^ n36404;
  assign n34123 = ~n34463 & ~n34109;
  assign n34110 = ~n34116 | ~n34448;
  assign n34111 = ~n34110 | ~n34469;
  assign n34121 = ~n34111 | ~P3_EBX_REG_16__SCAN_IN;
  assign n34113 = ~n34430 | ~n34112;
  assign n34115 = ~n34113 & ~P3_REIP_REG_16__SCAN_IN;
  assign n34114 = ~n36412 & ~n34459;
  assign n34118 = ~n34115 & ~n34114;
  assign n34130 = ~n34116 & ~n34470;
  assign n34117 = ~n34130 | ~n35121;
  assign n34119 = ~n34118 | ~n34117;
  assign n34120 = ~n22843 & ~n34119;
  assign n34122 = ~n34121 | ~n34120;
  assign n34124 = ~n34123 & ~n34122;
  assign P3_U2655 = ~n34125 | ~n34124;
  assign n34137 = ~n34127 & ~n34126;
  assign n34129 = ~P3_EBX_REG_15__SCAN_IN | ~n34128;
  assign n34135 = ~n34130 | ~n34129;
  assign n34132 = ~P3_EBX_REG_15__SCAN_IN | ~n34445;
  assign n34131 = ~n34384 | ~P3_PHYADDRPOINTER_REG_15__SCAN_IN;
  assign n34133 = ~n34132 | ~n34131;
  assign n34134 = ~n22843 & ~n34133;
  assign n34136 = ~n34135 | ~n34134;
  assign n34144 = ~n34137 & ~n34136;
  assign n34142 = ~n34147 & ~n38930;
  assign n36444 = n36447 ^ n36410;
  assign n34139 = ~n34425 | ~n34138;
  assign n34140 = ~n36444 ^ n34139;
  assign n34141 = ~n34463 & ~n34140;
  assign n34143 = ~n34142 & ~n34141;
  assign P3_U2656 = ~n34144 | ~n34143;
  assign n34146 = ~n34430 | ~n34145;
  assign n38925 = ~P3_REIP_REG_14__SCAN_IN;
  assign n34149 = ~n34146 | ~n38925;
  assign n34148 = ~n34147;
  assign n34153 = ~n34149 | ~n34148;
  assign n34150 = ~n34154 | ~n34448;
  assign n34151 = ~n34150 | ~n34469;
  assign n34152 = ~n34151 | ~P3_EBX_REG_14__SCAN_IN;
  assign n34158 = ~n34153 | ~n34152;
  assign n34156 = ~P3_PHYADDRPOINTER_REG_14__SCAN_IN | ~n34384;
  assign n34169 = ~n34154 & ~n34470;
  assign n34155 = ~n34169 | ~n35190;
  assign n34157 = ~n34156 | ~n34155;
  assign n34164 = ~n34158 & ~n34157;
  assign n36459 = n36455 ^ n34179;
  assign n34159 = ~P3_PHYADDRPOINTER_REG_0__SCAN_IN & ~n34179;
  assign n34160 = ~n34376 & ~n34159;
  assign n34161 = ~n36459 ^ n34160;
  assign n34162 = ~n34463 & ~n34161;
  assign n34163 = ~n22843 & ~n34162;
  assign P3_U2657 = ~n34164 | ~n34163;
  assign n38915 = ~P3_REIP_REG_12__SCAN_IN;
  assign n34193 = ~n34430 | ~n38915;
  assign n34165 = ~n34191 & ~n34405;
  assign n34222 = ~n34371 & ~n34165;
  assign n34166 = ~n34193 | ~n34222;
  assign n34188 = ~n34166 | ~P3_REIP_REG_13__SCAN_IN;
  assign n34168 = ~P3_EBX_REG_13__SCAN_IN | ~n34167;
  assign n34171 = ~n34169 | ~n34168;
  assign n34170 = ~P3_EBX_REG_13__SCAN_IN | ~n34445;
  assign n34186 = ~n34171 | ~n34170;
  assign n34172 = ~n34430 | ~n38920;
  assign n34175 = ~n34173 & ~n34172;
  assign n34174 = ~n36483 & ~n34459;
  assign n34184 = ~n34175 & ~n34174;
  assign n34177 = ~P3_PHYADDRPOINTER_REG_12__SCAN_IN | ~n36477;
  assign n34176 = ~P3_PHYADDRPOINTER_REG_0__SCAN_IN & ~n34177;
  assign n34180 = ~n34376 & ~n34176;
  assign n34178 = ~n36483 | ~n34177;
  assign n36476 = ~n34179 | ~n34178;
  assign n34181 = n34180 ^ n36476;
  assign n34182 = ~n34463 & ~n34181;
  assign n34183 = ~n34182 & ~n22843;
  assign n34185 = ~n34184 | ~n34183;
  assign n34187 = ~n34186 & ~n34185;
  assign P3_U2658 = ~n34188 | ~n34187;
  assign n34200 = ~n36511 & ~n34459;
  assign n34190 = n34189 ^ P3_EBX_REG_12__SCAN_IN;
  assign n34195 = ~n34470 & ~n34190;
  assign n34192 = ~n34191;
  assign n34194 = ~n34193 & ~n34192;
  assign n34198 = ~n34195 & ~n34194;
  assign n34196 = ~n35273 & ~n34469;
  assign n34197 = ~n22843 & ~n34196;
  assign n34199 = ~n34198 | ~n34197;
  assign n34207 = ~n34200 & ~n34199;
  assign n34205 = ~n34222 & ~n38915;
  assign n36507 = n36511 ^ n36477;
  assign n34201 = ~n36477 | ~n36747;
  assign n34202 = ~n34425 | ~n34201;
  assign n34203 = ~n36507 ^ n34202;
  assign n34204 = ~n34463 & ~n34203;
  assign n34206 = ~n34205 & ~n34204;
  assign P3_U2659 = ~n34207 | ~n34206;
  assign n34208 = ~n36538 & ~n34459;
  assign n34210 = ~n34208 & ~n22843;
  assign n34209 = ~P3_EBX_REG_11__SCAN_IN | ~n34445;
  assign n34216 = ~n34210 | ~n34209;
  assign n34235 = ~n36537 & ~n34298;
  assign n34211 = ~P3_PHYADDRPOINTER_REG_11__SCAN_IN & ~n34235;
  assign n36535 = ~n36477 & ~n34211;
  assign n34212 = ~n34235 | ~n36747;
  assign n34213 = ~n34425 | ~n34212;
  assign n34214 = n36535 ^ n34213;
  assign n34215 = ~n34463 & ~n34214;
  assign n34226 = ~n34216 & ~n34215;
  assign n35279 = ~P3_EBX_REG_11__SCAN_IN;
  assign n34218 = n35279 ^ n34217;
  assign n34224 = ~n34470 & ~n34218;
  assign n34220 = ~n34405 & ~n34219;
  assign n34221 = ~P3_REIP_REG_11__SCAN_IN & ~n34220;
  assign n34223 = ~n34222 & ~n34221;
  assign n34225 = ~n34224 & ~n34223;
  assign P3_U2660 = ~n34226 | ~n34225;
  assign n34230 = ~n35353 & ~n34469;
  assign n34228 = P3_EBX_REG_10__SCAN_IN ^ n34227;
  assign n34229 = ~n34470 & ~n34228;
  assign n34248 = ~n34230 & ~n34229;
  assign n34232 = ~n34430 | ~n34231;
  assign n34233 = ~P3_REIP_REG_10__SCAN_IN & ~n34232;
  assign n34242 = ~n22843 & ~n34233;
  assign n36581 = ~P3_PHYADDRPOINTER_REG_10__SCAN_IN;
  assign n34240 = ~n34459 & ~n36581;
  assign n34252 = n36622 | n34298;
  assign n34236 = ~n36590 & ~n34252;
  assign n34234 = ~P3_PHYADDRPOINTER_REG_10__SCAN_IN & ~n34236;
  assign n36565 = ~n34235 & ~n34234;
  assign n34237 = ~n34236 | ~n36747;
  assign n34254 = ~n34425 | ~n34237;
  assign n34238 = n36565 ^ n34254;
  assign n34239 = ~n34463 & ~n34238;
  assign n34241 = ~n34240 & ~n34239;
  assign n34246 = ~n34242 | ~n34241;
  assign n38905 = ~P3_REIP_REG_10__SCAN_IN;
  assign n34266 = ~P3_REIP_REG_9__SCAN_IN & ~n34405;
  assign n34265 = ~n34243;
  assign n34286 = ~n34405 & ~n34265;
  assign n34244 = ~n34266 & ~n34291;
  assign n34245 = ~n38905 & ~n34244;
  assign n34247 = ~n34246 & ~n34245;
  assign P3_U2661 = ~n34248 | ~n34247;
  assign n35346 = ~P3_EBX_REG_9__SCAN_IN;
  assign n34249 = ~n34470 & ~n34251;
  assign n34250 = ~n34445 & ~n34249;
  assign n34270 = ~n35346 & ~n34250;
  assign n34278 = ~n34448 | ~n34251;
  assign n34264 = ~P3_EBX_REG_9__SCAN_IN & ~n34278;
  assign n36596 = n36590 ^ n34252;
  assign n34253 = ~n36596;
  assign n34259 = ~n34254 | ~n34253;
  assign n34422 = ~n34460 & ~P3_PHYADDRPOINTER_REG_0__SCAN_IN;
  assign n34273 = ~n36536 | ~n34422;
  assign n34256 = ~n36622 & ~n34273;
  assign n34255 = ~n34425 | ~n36596;
  assign n34257 = ~n34256 & ~n34255;
  assign n34258 = ~n34463 & ~n34257;
  assign n34262 = ~n34259 | ~n34258;
  assign n34260 = ~n34459 & ~n36590;
  assign n34261 = ~n22843 & ~n34260;
  assign n34263 = ~n34262 | ~n34261;
  assign n34268 = ~n34264 & ~n34263;
  assign n34267 = ~n34266 | ~n34265;
  assign n34269 = ~n34268 | ~n34267;
  assign n34272 = ~n34270 & ~n34269;
  assign n34271 = ~P3_REIP_REG_9__SCAN_IN | ~n34291;
  assign P3_U2662 = ~n34272 | ~n34271;
  assign n36615 = n36622 ^ n34298;
  assign n34274 = ~n34425 | ~n34273;
  assign n34275 = n36615 ^ n34274;
  assign n34290 = ~n34463 & ~n34275;
  assign n34277 = ~n34276 & ~n34279;
  assign n34284 = ~n34278 & ~n34277;
  assign n34280 = ~n34469 & ~n34279;
  assign n34282 = ~n34280 & ~n22843;
  assign n34281 = ~n34384 | ~P3_PHYADDRPOINTER_REG_8__SCAN_IN;
  assign n34283 = ~n34282 | ~n34281;
  assign n34288 = ~n34284 & ~n34283;
  assign n34287 = ~n34286 | ~n34285;
  assign n34289 = ~n34288 | ~n34287;
  assign n34293 = ~n34290 & ~n34289;
  assign n34292 = ~P3_REIP_REG_8__SCAN_IN | ~n34291;
  assign P3_U2663 = ~n34293 | ~n34292;
  assign n35439 = ~P3_EBX_REG_7__SCAN_IN;
  assign n34294 = ~n34470 & ~n34304;
  assign n34295 = ~n34445 & ~n34294;
  assign n34302 = ~n35439 & ~n34295;
  assign n34412 = ~n34460 & ~n36686;
  assign n34342 = ~P3_PHYADDRPOINTER_REG_4__SCAN_IN | ~n34412;
  assign n34321 = ~n34343 & ~n34342;
  assign n34296 = ~P3_PHYADDRPOINTER_REG_6__SCAN_IN | ~n34321;
  assign n34297 = ~n34309 | ~n34296;
  assign n36633 = ~n34298 | ~n34297;
  assign n34374 = ~n34422;
  assign n34299 = ~n36639 & ~n34374;
  assign n34331 = ~n34320 & ~n34299;
  assign n34300 = n36633 ^ n34331;
  assign n34301 = ~n34463 & ~n34300;
  assign n34316 = ~n34302 & ~n34301;
  assign n34326 = ~P3_REIP_REG_6__SCAN_IN & ~n34405;
  assign n34348 = n34405 | n34325;
  assign n34361 = ~n34478 | ~n34348;
  assign n34303 = ~n34326 & ~n34361;
  assign n34314 = ~n34303 & ~n38890;
  assign n34319 = ~n34448 | ~n34304;
  assign n34308 = ~n34319 & ~P3_EBX_REG_7__SCAN_IN;
  assign n34306 = ~n34430 | ~n38890;
  assign n34307 = ~n34306 & ~n34305;
  assign n34312 = ~n34308 & ~n34307;
  assign n34310 = ~n34459 & ~n34309;
  assign n34311 = ~n34310 & ~n22843;
  assign n34313 = ~n34312 | ~n34311;
  assign n34315 = ~n34314 & ~n34313;
  assign P3_U2664 = ~n34316 | ~n34315;
  assign n34318 = ~n34317 & ~n35447;
  assign n34339 = ~n34319 & ~n34318;
  assign n34324 = ~n34320 & ~n34321;
  assign n36654 = ~P3_PHYADDRPOINTER_REG_6__SCAN_IN;
  assign n36649 = ~n36654 ^ n34321;
  assign n34461 = ~n34376 & ~n36747;
  assign n34322 = ~n34461 & ~n34463;
  assign n34323 = ~n36649 | ~n34322;
  assign n34335 = ~n34324 & ~n34323;
  assign n34328 = ~n34326 | ~n34325;
  assign n34327 = ~n34384 | ~P3_PHYADDRPOINTER_REG_6__SCAN_IN;
  assign n34329 = ~n34328 | ~n34327;
  assign n34333 = ~n22843 & ~n34329;
  assign n34330 = ~n36649 & ~n34463;
  assign n34332 = ~n34331 | ~n34330;
  assign n34334 = ~n34333 | ~n34332;
  assign n34337 = ~n34335 & ~n34334;
  assign n34336 = ~P3_EBX_REG_6__SCAN_IN | ~n34445;
  assign n34338 = ~n34337 | ~n34336;
  assign n34341 = ~n34339 & ~n34338;
  assign n34340 = ~P3_REIP_REG_6__SCAN_IN | ~n34361;
  assign P3_U2665 = ~n34341 | ~n34340;
  assign n36670 = n34343 ^ n34342;
  assign n34344 = ~n36665 & ~n34374;
  assign n34372 = ~n34376 & ~n34344;
  assign n34345 = ~n36670 ^ n34372;
  assign n34360 = ~n34463 & ~n34345;
  assign n35455 = ~P3_EBX_REG_5__SCAN_IN;
  assign n34346 = ~n34470 & ~n34352;
  assign n34347 = ~n34445 & ~n34346;
  assign n34356 = ~n35455 & ~n34347;
  assign n34350 = ~n34349 & ~n34348;
  assign n34354 = ~n22843 & ~n34350;
  assign n34351 = ~P3_EBX_REG_5__SCAN_IN & ~n34470;
  assign n34353 = ~n34352 | ~n34351;
  assign n34355 = ~n34354 | ~n34353;
  assign n34358 = ~n34356 & ~n34355;
  assign n34357 = ~n34384 | ~P3_PHYADDRPOINTER_REG_5__SCAN_IN;
  assign n34359 = ~n34358 | ~n34357;
  assign n34363 = ~n34360 & ~n34359;
  assign n34362 = ~P3_REIP_REG_5__SCAN_IN | ~n34361;
  assign P3_U2666 = ~n34363 | ~n34362;
  assign n35815 = ~n39110;
  assign n39136 = ~n35815 & ~n39132;
  assign n37389 = ~P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN;
  assign n34364 = ~n34585 | ~n37389;
  assign n34368 = ~n39136 | ~n34364;
  assign n34365 = ~n34430 | ~n34369;
  assign n34366 = ~P3_REIP_REG_4__SCAN_IN & ~n34365;
  assign n34367 = ~n22843 & ~n34366;
  assign n34388 = ~n34368 | ~n34367;
  assign n38875 = ~P3_REIP_REG_4__SCAN_IN;
  assign n34370 = ~n34369 & ~n34405;
  assign n34404 = ~n34371 & ~n34370;
  assign n34383 = ~n38875 & ~n34404;
  assign n36692 = P3_PHYADDRPOINTER_REG_4__SCAN_IN ^ n34412;
  assign n34373 = ~n36692 & ~n34372;
  assign n34379 = ~n34373 & ~n34463;
  assign n34375 = ~n36686 & ~n34374;
  assign n34377 = ~n34376 & ~n34375;
  assign n34378 = ~n36692 | ~n34377;
  assign n34381 = ~n34379 | ~n34378;
  assign n34403 = ~n34389 & ~n34470;
  assign n34380 = ~n34403 | ~n34486;
  assign n34382 = ~n34381 | ~n34380;
  assign n34386 = ~n34383 & ~n34382;
  assign n34385 = ~P3_PHYADDRPOINTER_REG_4__SCAN_IN | ~n34384;
  assign n34387 = ~n34386 | ~n34385;
  assign n34393 = ~n34388 & ~n34387;
  assign n34390 = ~n34389 | ~n34448;
  assign n34391 = ~n34390 | ~n34469;
  assign n34392 = ~n34391 | ~P3_EBX_REG_4__SCAN_IN;
  assign P3_U2667 = ~n34393 | ~n34392;
  assign n36699 = ~P3_PHYADDRPOINTER_REG_3__SCAN_IN;
  assign n34400 = ~n36699 & ~n34459;
  assign n38742 = ~n23642 & ~n34395;
  assign n38736 = ~n38742 & ~n23643;
  assign n39039 = ~n38736 | ~n22844;
  assign n34398 = ~n39136 | ~n39039;
  assign n34397 = ~n34445 | ~P3_EBX_REG_3__SCAN_IN;
  assign n34399 = ~n34398 | ~n34397;
  assign n34419 = ~n34400 & ~n34399;
  assign n34402 = ~P3_EBX_REG_3__SCAN_IN | ~n34401;
  assign n34410 = ~n34403 | ~n34402;
  assign n38870 = ~P3_REIP_REG_3__SCAN_IN;
  assign n34408 = ~n34404 & ~n38870;
  assign n34429 = ~n34405 & ~n39084;
  assign n34406 = ~P3_REIP_REG_2__SCAN_IN | ~n34429;
  assign n34407 = ~P3_REIP_REG_3__SCAN_IN & ~n34406;
  assign n34409 = ~n34408 & ~n34407;
  assign n34417 = ~n34410 | ~n34409;
  assign n36717 = ~P3_PHYADDRPOINTER_REG_2__SCAN_IN;
  assign n34413 = ~n34460 & ~n36717;
  assign n34411 = ~P3_PHYADDRPOINTER_REG_3__SCAN_IN & ~n34413;
  assign n36703 = ~n34412 & ~n34411;
  assign n34420 = ~n34413 | ~n36747;
  assign n34414 = ~n34425 | ~n34420;
  assign n34415 = n36703 ^ n34414;
  assign n34416 = ~n34463 & ~n34415;
  assign n34418 = ~n34417 & ~n34416;
  assign P3_U2668 = ~n34419 | ~n34418;
  assign n34424 = ~n34421 | ~n34420;
  assign n36720 = n34460 ^ P3_PHYADDRPOINTER_REG_2__SCAN_IN;
  assign n34423 = ~n34422 & ~n36720;
  assign n34428 = ~n34424 & ~n34423;
  assign n34426 = n34463 | n34425;
  assign n34427 = ~n34426 & ~n36720;
  assign n34444 = ~n34428 & ~n34427;
  assign n38865 = ~P3_REIP_REG_2__SCAN_IN;
  assign n34433 = ~n38865 | ~n34429;
  assign n34455 = ~n34430 | ~n39084;
  assign n34431 = ~n34478 | ~n34455;
  assign n34432 = ~n34431 | ~P3_REIP_REG_2__SCAN_IN;
  assign n34442 = ~n34433 | ~n34432;
  assign n34474 = ~n39136;
  assign n39047 = ~n38725 ^ P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n34435 = ~n34474 & ~n39047;
  assign n34434 = ~n36717 & ~n34459;
  assign n34440 = ~n34435 & ~n34434;
  assign n34438 = ~n34484 & ~n34469;
  assign n34436 = P3_EBX_REG_2__SCAN_IN ^ n34447;
  assign n34437 = ~n34470 & ~n34436;
  assign n34439 = ~n34438 & ~n34437;
  assign n34441 = ~n34440 | ~n34439;
  assign n34443 = ~n34442 & ~n34441;
  assign P3_U2669 = ~n34444 | ~n34443;
  assign n34450 = ~P3_EBX_REG_1__SCAN_IN | ~n34445;
  assign n35472 = ~P3_EBX_REG_0__SCAN_IN | ~P3_EBX_REG_1__SCAN_IN;
  assign n34446 = ~n35472;
  assign n35482 = ~n34447 & ~n34446;
  assign n34449 = ~n35482 | ~n34448;
  assign n34458 = ~n34450 | ~n34449;
  assign n34452 = ~n34451;
  assign n39057 = ~n34452 | ~n38723;
  assign n34454 = ~n34474 & ~n39057;
  assign n34453 = ~n34478 & ~n39084;
  assign n34456 = ~n34454 & ~n34453;
  assign n34457 = ~n34456 | ~n34455;
  assign n34467 = ~n34458 & ~n34457;
  assign n34465 = ~n34460 & ~n34459;
  assign n34462 = P3_PHYADDRPOINTER_REG_1__SCAN_IN ^ n34461;
  assign n34464 = ~n34463 & ~n34462;
  assign n34466 = ~n34465 & ~n34464;
  assign P3_U2670 = ~n34467 | ~n34466;
  assign n34473 = n39083 | n34468;
  assign n34471 = ~n34470 | ~n34469;
  assign n34472 = ~P3_EBX_REG_0__SCAN_IN | ~n34471;
  assign n34476 = ~n34473 | ~n34472;
  assign n34475 = ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN & ~n34474;
  assign n34480 = ~n34476 & ~n34475;
  assign n39073 = ~n39056;
  assign n34477 = ~n39073 & ~n36747;
  assign n34479 = ~n34478 | ~n34477;
  assign P3_U2671 = ~n34480 | ~n34479;
  assign n34482 = ~n39105 | ~n34481;
  assign n35192 = ~P3_EBX_REG_14__SCAN_IN | ~P3_EBX_REG_13__SCAN_IN;
  assign n35460 = ~n34484 & ~n35472;
  assign n34485 = ~P3_EBX_REG_3__SCAN_IN | ~n35460;
  assign n35446 = ~n34486 & ~n34485;
  assign n34487 = ~n35447 & ~n35455;
  assign n35441 = ~n35446 | ~n34487;
  assign n34488 = ~n35439 & ~n35441;
  assign n35345 = ~P3_EBX_REG_8__SCAN_IN | ~n34488;
  assign n35119 = ~n35353 & ~n35346;
  assign n35348 = ~n35119;
  assign n34489 = ~n35345 & ~n35348;
  assign n35272 = ~P3_EBX_REG_11__SCAN_IN | ~n34489;
  assign n35200 = ~n35273 & ~n35272;
  assign n34490 = ~P3_EBX_REG_15__SCAN_IN | ~n35200;
  assign n35113 = ~n35192 & ~n34490;
  assign n35046 = ~P3_EBX_REG_16__SCAN_IN | ~n35113;
  assign n35009 = ~n35078 & ~n35046;
  assign n34491 = ~n35394 | ~n35009;
  assign n34802 = ~P3_EBX_REG_19__SCAN_IN | ~n35006;
  assign n34933 = ~n34493 & ~n34802;
  assign n34496 = ~n34494 & ~n34804;
  assign n34495 = ~n34893 & ~n34803;
  assign n34500 = ~n34496 | ~n34495;
  assign n34812 = ~P3_EBX_REG_28__SCAN_IN | ~P3_EBX_REG_27__SCAN_IN;
  assign n34497 = ~P3_EBX_REG_26__SCAN_IN | ~P3_EBX_REG_29__SCAN_IN;
  assign n34498 = ~n34812 & ~n34497;
  assign n34499 = ~P3_EBX_REG_25__SCAN_IN | ~n34498;
  assign n34501 = ~n34500 & ~n34499;
  assign n34508 = ~n34933 | ~n34501;
  assign n34504 = ~n34507 & ~n34508;
  assign n34502 = ~n35477 & ~n34504;
  assign n34506 = ~P3_EBX_REG_31__SCAN_IN | ~n34502;
  assign n34503 = ~P3_EBX_REG_31__SCAN_IN & ~n37514;
  assign n34505 = ~n34504 | ~n34503;
  assign P3_U2672 = ~n34506 | ~n34505;
  assign n34509 = n34508 ^ n34507;
  assign n34801 = ~n34509 | ~n35487;
  assign n34511 = ~n24451 | ~P3_INSTQUEUE_REG_13__7__SCAN_IN;
  assign n34510 = ~n34545 | ~P3_INSTQUEUE_REG_9__7__SCAN_IN;
  assign n34515 = ~n34511 | ~n34510;
  assign n34513 = ~n24470 | ~P3_INSTQUEUE_REG_6__7__SCAN_IN;
  assign n34512 = ~n34564 | ~P3_INSTQUEUE_REG_3__7__SCAN_IN;
  assign n34514 = ~n34513 | ~n34512;
  assign n34524 = ~n34515 & ~n34514;
  assign n34518 = ~n35328 | ~P3_INSTQUEUE_REG_5__7__SCAN_IN;
  assign n34517 = ~n24543 | ~P3_INSTQUEUE_REG_8__7__SCAN_IN;
  assign n34522 = ~n34518 | ~n34517;
  assign n34520 = ~n34993 | ~P3_INSTQUEUE_REG_7__7__SCAN_IN;
  assign n34519 = ~n24516 | ~P3_INSTQUEUE_REG_0__7__SCAN_IN;
  assign n34521 = ~n34520 | ~n34519;
  assign n34523 = ~n34522 & ~n34521;
  assign n34542 = ~n34524 | ~n34523;
  assign n34527 = ~n34872 | ~P3_INSTQUEUE_REG_2__7__SCAN_IN;
  assign n34526 = ~n35405 | ~P3_INSTQUEUE_REG_4__7__SCAN_IN;
  assign n34531 = ~n34527 | ~n34526;
  assign n34529 = ~n35412 | ~P3_INSTQUEUE_REG_10__7__SCAN_IN;
  assign n34528 = ~n24513 | ~P3_INSTQUEUE_REG_14__7__SCAN_IN;
  assign n34530 = ~n34529 | ~n34528;
  assign n34540 = ~n34531 & ~n34530;
  assign n34534 = ~n34717 | ~P3_INSTQUEUE_REG_15__7__SCAN_IN;
  assign n34533 = ~n35319 | ~P3_INSTQUEUE_REG_12__7__SCAN_IN;
  assign n34538 = ~n34534 | ~n34533;
  assign n34536 = ~n35366 | ~P3_INSTQUEUE_REG_11__7__SCAN_IN;
  assign n34535 = ~n35252 | ~P3_INSTQUEUE_REG_1__7__SCAN_IN;
  assign n34537 = ~n34536 | ~n34535;
  assign n34539 = ~n34538 & ~n34537;
  assign n34541 = ~n34540 | ~n34539;
  assign n34799 = ~n34542 & ~n34541;
  assign n34544 = ~n24470 | ~P3_INSTQUEUE_REG_6__5__SCAN_IN;
  assign n34543 = ~n24516 | ~P3_INSTQUEUE_REG_0__5__SCAN_IN;
  assign n34549 = ~n34544 | ~n34543;
  assign n34547 = ~n34545 | ~P3_INSTQUEUE_REG_9__5__SCAN_IN;
  assign n34546 = ~n24513 | ~P3_INSTQUEUE_REG_14__5__SCAN_IN;
  assign n34548 = ~n34547 | ~n34546;
  assign n34557 = ~n34549 & ~n34548;
  assign n34551 = ~n24451 | ~P3_INSTQUEUE_REG_13__5__SCAN_IN;
  assign n34550 = ~n35328 | ~P3_INSTQUEUE_REG_5__5__SCAN_IN;
  assign n34555 = ~n34551 | ~n34550;
  assign n34553 = ~n35319 | ~P3_INSTQUEUE_REG_12__5__SCAN_IN;
  assign n34552 = ~n24543 | ~P3_INSTQUEUE_REG_8__5__SCAN_IN;
  assign n34554 = ~n34553 | ~n34552;
  assign n34556 = ~n34555 & ~n34554;
  assign n34574 = ~n34557 | ~n34556;
  assign n34559 = ~n35366 | ~P3_INSTQUEUE_REG_11__5__SCAN_IN;
  assign n34558 = ~n35252 | ~P3_INSTQUEUE_REG_1__5__SCAN_IN;
  assign n34563 = ~n34559 | ~n34558;
  assign n34561 = ~n35412 | ~P3_INSTQUEUE_REG_10__5__SCAN_IN;
  assign n34560 = ~n34872 | ~P3_INSTQUEUE_REG_2__5__SCAN_IN;
  assign n34562 = ~n34561 | ~n34560;
  assign n34572 = ~n34563 & ~n34562;
  assign n34566 = ~n34717 | ~P3_INSTQUEUE_REG_15__5__SCAN_IN;
  assign n34565 = ~n34564 | ~P3_INSTQUEUE_REG_3__5__SCAN_IN;
  assign n34570 = ~n34566 | ~n34565;
  assign n34568 = ~n35405 | ~P3_INSTQUEUE_REG_4__5__SCAN_IN;
  assign n34567 = ~n34993 | ~P3_INSTQUEUE_REG_7__5__SCAN_IN;
  assign n34569 = ~n34568 | ~n34567;
  assign n34571 = ~n34570 & ~n34569;
  assign n34573 = ~n34572 | ~n34571;
  assign n34819 = ~n34574 & ~n34573;
  assign n34577 = ~n24535 | ~P3_INSTQUEUE_REG_9__3__SCAN_IN;
  assign n34576 = ~n35405 | ~P3_INSTQUEUE_REG_4__3__SCAN_IN;
  assign n34582 = ~n34577 | ~n34576;
  assign n34580 = ~n24513 | ~P3_INSTQUEUE_REG_14__3__SCAN_IN;
  assign n34579 = ~n34993 | ~P3_INSTQUEUE_REG_7__3__SCAN_IN;
  assign n34581 = ~n34580 | ~n34579;
  assign n34591 = ~n34582 & ~n34581;
  assign n34584 = ~n24451 | ~P3_INSTQUEUE_REG_13__3__SCAN_IN;
  assign n34583 = ~n35252 | ~P3_INSTQUEUE_REG_1__3__SCAN_IN;
  assign n34589 = ~n34584 | ~n34583;
  assign n34587 = ~n34717 | ~P3_INSTQUEUE_REG_15__3__SCAN_IN;
  assign n35359 = ~n34585;
  assign n34586 = ~n35359 | ~P3_INSTQUEUE_REG_3__3__SCAN_IN;
  assign n34588 = ~n34587 | ~n34586;
  assign n34590 = ~n34589 & ~n34588;
  assign n34607 = ~n34591 | ~n34590;
  assign n34593 = ~n24543 | ~P3_INSTQUEUE_REG_8__3__SCAN_IN;
  assign n34592 = ~n24516 | ~P3_INSTQUEUE_REG_0__3__SCAN_IN;
  assign n34597 = ~n34593 | ~n34592;
  assign n34595 = ~n35412 | ~P3_INSTQUEUE_REG_10__3__SCAN_IN;
  assign n34594 = ~n34872 | ~P3_INSTQUEUE_REG_2__3__SCAN_IN;
  assign n34596 = ~n34595 | ~n34594;
  assign n34605 = ~n34597 & ~n34596;
  assign n34599 = ~n35366 | ~P3_INSTQUEUE_REG_11__3__SCAN_IN;
  assign n34598 = ~n35319 | ~P3_INSTQUEUE_REG_12__3__SCAN_IN;
  assign n34603 = ~n34599 | ~n34598;
  assign n34601 = ~n35328 | ~P3_INSTQUEUE_REG_5__3__SCAN_IN;
  assign n34600 = ~n24470 | ~P3_INSTQUEUE_REG_6__3__SCAN_IN;
  assign n34602 = ~n34601 | ~n34600;
  assign n34604 = ~n34603 & ~n34602;
  assign n34606 = ~n34605 | ~n34604;
  assign n34834 = ~n34607 & ~n34606;
  assign n34609 = ~n35252 | ~P3_INSTQUEUE_REG_1__1__SCAN_IN;
  assign n34608 = ~n24543 | ~P3_INSTQUEUE_REG_8__1__SCAN_IN;
  assign n34614 = ~n34609 | ~n34608;
  assign n34612 = ~n35405 | ~P3_INSTQUEUE_REG_4__1__SCAN_IN;
  assign n34611 = ~n34993 | ~P3_INSTQUEUE_REG_7__1__SCAN_IN;
  assign n34613 = ~n34612 | ~n34611;
  assign n34622 = ~n34614 & ~n34613;
  assign n34616 = ~n24470 | ~P3_INSTQUEUE_REG_6__1__SCAN_IN;
  assign n34615 = ~n24516 | ~P3_INSTQUEUE_REG_0__1__SCAN_IN;
  assign n34620 = ~n34616 | ~n34615;
  assign n35366 = ~n22844;
  assign n34618 = ~n35366 | ~P3_INSTQUEUE_REG_11__1__SCAN_IN;
  assign n34617 = ~n35359 | ~P3_INSTQUEUE_REG_3__1__SCAN_IN;
  assign n34619 = ~n34618 | ~n34617;
  assign n34621 = ~n34620 & ~n34619;
  assign n34639 = ~n34622 | ~n34621;
  assign n34624 = ~n24513 | ~P3_INSTQUEUE_REG_14__1__SCAN_IN;
  assign n34623 = ~n34872 | ~P3_INSTQUEUE_REG_2__1__SCAN_IN;
  assign n34628 = ~n34624 | ~n34623;
  assign n34626 = ~n35412 | ~P3_INSTQUEUE_REG_10__1__SCAN_IN;
  assign n34625 = ~n35319 | ~P3_INSTQUEUE_REG_12__1__SCAN_IN;
  assign n34627 = ~n34626 | ~n34625;
  assign n34637 = ~n34628 & ~n34627;
  assign n34630 = ~n34717 | ~P3_INSTQUEUE_REG_15__1__SCAN_IN;
  assign n34629 = ~n35328 | ~P3_INSTQUEUE_REG_5__1__SCAN_IN;
  assign n34635 = ~n34630 | ~n34629;
  assign n34633 = ~n24451 | ~P3_INSTQUEUE_REG_13__1__SCAN_IN;
  assign n34632 = ~n24535 | ~P3_INSTQUEUE_REG_9__1__SCAN_IN;
  assign n34634 = ~n34633 | ~n34632;
  assign n34636 = ~n34635 & ~n34634;
  assign n34638 = ~n34637 | ~n34636;
  assign n34848 = ~n34639 & ~n34638;
  assign n34641 = ~n34717 | ~P3_INSTQUEUE_REG_15__0__SCAN_IN;
  assign n34640 = ~n24470 | ~P3_INSTQUEUE_REG_6__0__SCAN_IN;
  assign n34645 = ~n34641 | ~n34640;
  assign n34643 = ~n24451 | ~P3_INSTQUEUE_REG_13__0__SCAN_IN;
  assign n34642 = ~n35252 | ~P3_INSTQUEUE_REG_1__0__SCAN_IN;
  assign n34644 = ~n34643 | ~n34642;
  assign n34670 = ~n34645 & ~n34644;
  assign n34647 = ~n35405 | ~P3_INSTQUEUE_REG_4__0__SCAN_IN;
  assign n34646 = ~n24516 | ~P3_INSTQUEUE_REG_0__0__SCAN_IN;
  assign n34651 = ~n34647 | ~n34646;
  assign n34649 = ~n35319 | ~P3_INSTQUEUE_REG_12__0__SCAN_IN;
  assign n34648 = ~n35359 | ~P3_INSTQUEUE_REG_3__0__SCAN_IN;
  assign n34650 = ~n34649 | ~n34648;
  assign n34668 = n34651 | n34650;
  assign n34653 = ~n24535 | ~P3_INSTQUEUE_REG_9__0__SCAN_IN;
  assign n34652 = ~n35366 | ~P3_INSTQUEUE_REG_11__0__SCAN_IN;
  assign n34657 = ~n34653 | ~n34652;
  assign n34655 = ~n35412 | ~P3_INSTQUEUE_REG_10__0__SCAN_IN;
  assign n34654 = ~n34872 | ~P3_INSTQUEUE_REG_2__0__SCAN_IN;
  assign n34656 = ~n34655 | ~n34654;
  assign n34666 = ~n34657 & ~n34656;
  assign n34659 = ~n24513 | ~P3_INSTQUEUE_REG_14__0__SCAN_IN;
  assign n34658 = ~n34993 | ~P3_INSTQUEUE_REG_7__0__SCAN_IN;
  assign n34664 = ~n34659 | ~n34658;
  assign n34662 = ~n35328 | ~P3_INSTQUEUE_REG_5__0__SCAN_IN;
  assign n34661 = ~n24543 | ~P3_INSTQUEUE_REG_8__0__SCAN_IN;
  assign n34663 = ~n34662 | ~n34661;
  assign n34665 = ~n34664 & ~n34663;
  assign n34667 = ~n34666 | ~n34665;
  assign n34669 = ~n34668 & ~n34667;
  assign n34856 = ~n34670 | ~n34669;
  assign n34672 = ~n35366 | ~P3_INSTQUEUE_REG_10__7__SCAN_IN;
  assign n34671 = ~n35252 | ~P3_INSTQUEUE_REG_0__7__SCAN_IN;
  assign n34676 = ~n34672 | ~n34671;
  assign n34674 = ~n24535 | ~P3_INSTQUEUE_REG_8__7__SCAN_IN;
  assign n34673 = ~n24470 | ~P3_INSTQUEUE_REG_5__7__SCAN_IN;
  assign n34675 = ~n34674 | ~n34673;
  assign n34700 = ~n34676 & ~n34675;
  assign n34678 = ~n35405 | ~P3_INSTQUEUE_REG_3__7__SCAN_IN;
  assign n34677 = ~n24516 | ~P3_INSTQUEUE_REG_15__7__SCAN_IN;
  assign n34682 = ~n34678 | ~n34677;
  assign n34680 = ~n24543 | ~P3_INSTQUEUE_REG_7__7__SCAN_IN;
  assign n34679 = ~n35359 | ~P3_INSTQUEUE_REG_2__7__SCAN_IN;
  assign n34681 = ~n34680 | ~n34679;
  assign n34698 = n34682 | n34681;
  assign n34684 = ~n34717 | ~P3_INSTQUEUE_REG_14__7__SCAN_IN;
  assign n34683 = ~n34993 | ~P3_INSTQUEUE_REG_6__7__SCAN_IN;
  assign n34688 = ~n34684 | ~n34683;
  assign n34686 = ~n35412 | ~P3_INSTQUEUE_REG_9__7__SCAN_IN;
  assign n34685 = ~n34872 | ~P3_INSTQUEUE_REG_1__7__SCAN_IN;
  assign n34687 = ~n34686 | ~n34685;
  assign n34696 = ~n34688 & ~n34687;
  assign n34690 = ~n24513 | ~P3_INSTQUEUE_REG_13__7__SCAN_IN;
  assign n34689 = ~n35328 | ~P3_INSTQUEUE_REG_4__7__SCAN_IN;
  assign n34694 = ~n34690 | ~n34689;
  assign n34692 = ~n24451 | ~P3_INSTQUEUE_REG_12__7__SCAN_IN;
  assign n34691 = ~n35319 | ~P3_INSTQUEUE_REG_11__7__SCAN_IN;
  assign n34693 = ~n34692 | ~n34691;
  assign n34695 = ~n34694 & ~n34693;
  assign n34697 = ~n34696 | ~n34695;
  assign n34699 = ~n34698 & ~n34697;
  assign n34855 = ~n34700 | ~n34699;
  assign n34847 = ~n34856 | ~n34855;
  assign n34841 = ~n34848 & ~n34847;
  assign n34702 = ~n35319 | ~P3_INSTQUEUE_REG_12__2__SCAN_IN;
  assign n34701 = ~n35405 | ~P3_INSTQUEUE_REG_4__2__SCAN_IN;
  assign n34706 = ~n34702 | ~n34701;
  assign n34704 = ~n24535 | ~P3_INSTQUEUE_REG_9__2__SCAN_IN;
  assign n34703 = ~n24543 | ~P3_INSTQUEUE_REG_8__2__SCAN_IN;
  assign n34705 = ~n34704 | ~n34703;
  assign n34731 = ~n34706 & ~n34705;
  assign n34708 = ~n24513 | ~P3_INSTQUEUE_REG_14__2__SCAN_IN;
  assign n34707 = ~n35252 | ~P3_INSTQUEUE_REG_1__2__SCAN_IN;
  assign n34729 = ~n34708 | ~n34707;
  assign n34710 = ~n35412 | ~P3_INSTQUEUE_REG_10__2__SCAN_IN;
  assign n34709 = ~n35366 | ~P3_INSTQUEUE_REG_11__2__SCAN_IN;
  assign n34714 = ~n34710 | ~n34709;
  assign n34712 = ~n34872 | ~P3_INSTQUEUE_REG_2__2__SCAN_IN;
  assign n34711 = ~n35359 | ~P3_INSTQUEUE_REG_3__2__SCAN_IN;
  assign n34713 = ~n34712 | ~n34711;
  assign n34727 = ~n34714 & ~n34713;
  assign n34716 = ~n24451 | ~P3_INSTQUEUE_REG_13__2__SCAN_IN;
  assign n34715 = ~n35328 | ~P3_INSTQUEUE_REG_5__2__SCAN_IN;
  assign n34721 = ~n34716 | ~n34715;
  assign n34719 = ~n34717 | ~P3_INSTQUEUE_REG_15__2__SCAN_IN;
  assign n34718 = ~n24516 | ~P3_INSTQUEUE_REG_0__2__SCAN_IN;
  assign n34720 = ~n34719 | ~n34718;
  assign n34725 = n34721 | n34720;
  assign n34723 = ~n24470 | ~P3_INSTQUEUE_REG_6__2__SCAN_IN;
  assign n34722 = ~n34993 | ~P3_INSTQUEUE_REG_7__2__SCAN_IN;
  assign n34724 = ~n34723 | ~n34722;
  assign n34726 = ~n34725 & ~n34724;
  assign n34728 = ~n34727 | ~n34726;
  assign n34730 = ~n34729 & ~n34728;
  assign n34840 = ~n34731 | ~n34730;
  assign n34833 = ~n34841 | ~n34840;
  assign n34826 = ~n34834 & ~n34833;
  assign n34733 = ~n35366 | ~P3_INSTQUEUE_REG_11__4__SCAN_IN;
  assign n34732 = ~n35319 | ~P3_INSTQUEUE_REG_12__4__SCAN_IN;
  assign n34737 = ~n34733 | ~n34732;
  assign n34735 = ~n24470 | ~P3_INSTQUEUE_REG_6__4__SCAN_IN;
  assign n34734 = ~n34993 | ~P3_INSTQUEUE_REG_7__4__SCAN_IN;
  assign n34736 = ~n34735 | ~n34734;
  assign n34761 = ~n34737 & ~n34736;
  assign n34739 = ~n24513 | ~P3_INSTQUEUE_REG_14__4__SCAN_IN;
  assign n34738 = ~n35252 | ~P3_INSTQUEUE_REG_1__4__SCAN_IN;
  assign n34759 = ~n34739 | ~n34738;
  assign n34741 = ~n24535 | ~P3_INSTQUEUE_REG_9__4__SCAN_IN;
  assign n34740 = ~n35359 | ~P3_INSTQUEUE_REG_3__4__SCAN_IN;
  assign n34745 = ~n34741 | ~n34740;
  assign n34743 = ~n35412 | ~P3_INSTQUEUE_REG_10__4__SCAN_IN;
  assign n34742 = ~n34872 | ~P3_INSTQUEUE_REG_2__4__SCAN_IN;
  assign n34744 = ~n34743 | ~n34742;
  assign n34757 = ~n34745 & ~n34744;
  assign n34747 = ~n24451 | ~P3_INSTQUEUE_REG_13__4__SCAN_IN;
  assign n34746 = ~n35328 | ~P3_INSTQUEUE_REG_5__4__SCAN_IN;
  assign n34751 = ~n34747 | ~n34746;
  assign n34749 = ~n35405 | ~P3_INSTQUEUE_REG_4__4__SCAN_IN;
  assign n34748 = ~n24516 | ~P3_INSTQUEUE_REG_0__4__SCAN_IN;
  assign n34750 = ~n34749 | ~n34748;
  assign n34755 = n34751 | n34750;
  assign n34753 = ~n34717 | ~P3_INSTQUEUE_REG_15__4__SCAN_IN;
  assign n34752 = ~n24543 | ~P3_INSTQUEUE_REG_8__4__SCAN_IN;
  assign n34754 = ~n34753 | ~n34752;
  assign n34756 = ~n34755 & ~n34754;
  assign n34758 = ~n34757 | ~n34756;
  assign n34760 = ~n34759 & ~n34758;
  assign n34825 = ~n34761 | ~n34760;
  assign n34818 = ~n34826 | ~n34825;
  assign n34809 = ~n34819 & ~n34818;
  assign n34763 = ~n24513 | ~P3_INSTQUEUE_REG_14__6__SCAN_IN;
  assign n34762 = ~n35366 | ~P3_INSTQUEUE_REG_11__6__SCAN_IN;
  assign n34767 = ~n34763 | ~n34762;
  assign n34765 = ~n34717 | ~P3_INSTQUEUE_REG_15__6__SCAN_IN;
  assign n34764 = ~n35328 | ~P3_INSTQUEUE_REG_5__6__SCAN_IN;
  assign n34766 = ~n34765 | ~n34764;
  assign n34797 = ~n34767 & ~n34766;
  assign n34769 = ~n24451 | ~P3_INSTQUEUE_REG_13__6__SCAN_IN;
  assign n34768 = ~n24543 | ~P3_INSTQUEUE_REG_8__6__SCAN_IN;
  assign n34795 = ~n34769 | ~n34768;
  assign n34771 = ~n35405 | ~P3_INSTQUEUE_REG_4__6__SCAN_IN;
  assign n34770 = ~n34993 | ~P3_INSTQUEUE_REG_7__6__SCAN_IN;
  assign n34775 = ~n34771 | ~n34770;
  assign n34773 = ~n35412 | ~P3_INSTQUEUE_REG_10__6__SCAN_IN;
  assign n34772 = ~n34872 | ~P3_INSTQUEUE_REG_2__6__SCAN_IN;
  assign n34774 = ~n34773 | ~n34772;
  assign n34793 = ~n34775 & ~n34774;
  assign n34776 = ~P3_INSTQUEUE_REG_9__6__SCAN_IN;
  assign n34781 = ~n34777 & ~n34776;
  assign n34780 = ~n34779 & ~n34778;
  assign n34787 = ~n34781 & ~n34780;
  assign n37505 = ~P3_INSTQUEUE_REG_0__6__SCAN_IN;
  assign n34785 = ~n34782 & ~n37505;
  assign n34784 = ~n34585 & ~n34783;
  assign n34786 = ~n34785 & ~n34784;
  assign n34791 = ~n34787 | ~n34786;
  assign n34789 = ~n35252 | ~P3_INSTQUEUE_REG_1__6__SCAN_IN;
  assign n34788 = ~n35319 | ~P3_INSTQUEUE_REG_12__6__SCAN_IN;
  assign n34790 = ~n34789 | ~n34788;
  assign n34792 = ~n34791 & ~n34790;
  assign n34794 = ~n34793 | ~n34792;
  assign n34796 = ~n34795 & ~n34794;
  assign n34808 = ~n34797 | ~n34796;
  assign n34798 = ~n34809 | ~n34808;
  assign n35511 = n34799 ^ n34798;
  assign n34800 = ~n35477 | ~n35511;
  assign P3_U2673 = ~n34801 | ~n34800;
  assign n34966 = ~n37514 & ~n34802;
  assign n34900 = ~P3_EBX_REG_20__SCAN_IN | ~n34966;
  assign n34895 = ~n34803 & ~n34900;
  assign n34897 = ~P3_EBX_REG_22__SCAN_IN | ~n34895;
  assign n34849 = ~n34804 & ~n34897;
  assign n34851 = ~P3_EBX_REG_24__SCAN_IN | ~n34849;
  assign n34816 = ~n34806 & ~n34843;
  assign n34836 = ~n34816;
  assign n34807 = n34836 | n34812;
  assign n34811 = ~P3_EBX_REG_29__SCAN_IN & ~n34807;
  assign n35520 = ~n34809 ^ n34808;
  assign n34810 = ~n35520 & ~n35391;
  assign n34815 = ~n34811 & ~n34810;
  assign n34828 = ~n35487 | ~n34836;
  assign n35486 = ~n34971 | ~n35394;
  assign n35483 = ~n35486;
  assign n34813 = ~n35483 | ~n34812;
  assign n34822 = ~n34828 | ~n34813;
  assign n34814 = ~P3_EBX_REG_29__SCAN_IN | ~n34822;
  assign P3_U2674 = ~n34815 | ~n34814;
  assign n34817 = ~P3_EBX_REG_27__SCAN_IN | ~n34816;
  assign n34821 = ~P3_EBX_REG_28__SCAN_IN & ~n34817;
  assign n35530 = ~n34819 ^ n34818;
  assign n34820 = ~n35530 & ~n35487;
  assign n34824 = ~n34821 & ~n34820;
  assign n34823 = ~P3_EBX_REG_28__SCAN_IN | ~n34822;
  assign P3_U2675 = ~n34824 | ~n34823;
  assign n35541 = n34826 ^ n34825;
  assign n34832 = ~n35541 | ~n35477;
  assign n34830 = ~n34828 & ~n34827;
  assign n34829 = ~P3_EBX_REG_27__SCAN_IN & ~n34836;
  assign n34831 = ~n34830 & ~n34829;
  assign P3_U2676 = ~n34832 | ~n34831;
  assign n35551 = n34834 ^ n34833;
  assign n34839 = ~n35551 | ~n35477;
  assign n34835 = ~n35391 | ~P3_EBX_REG_26__SCAN_IN;
  assign n34837 = ~n34835 | ~n34843;
  assign n34838 = ~n34837 | ~n34836;
  assign P3_U2677 = ~n34839 | ~n34838;
  assign n35564 = ~n34841 ^ n34840;
  assign n34846 = n35564 | n35391;
  assign n34842 = ~n35391 | ~P3_EBX_REG_25__SCAN_IN;
  assign n34844 = ~n34842 | ~n34851;
  assign n34845 = ~n34844 | ~n34843;
  assign P3_U2678 = ~n34846 | ~n34845;
  assign n35578 = ~n34848 ^ n34847;
  assign n34854 = n35578 | n35391;
  assign n34850 = ~n35391 | ~P3_EBX_REG_24__SCAN_IN;
  assign n34858 = ~n34849;
  assign n34852 = ~n34850 | ~n34858;
  assign n34853 = ~n34852 | ~n34851;
  assign P3_U2679 = ~n34854 | ~n34853;
  assign n35585 = n34856 ^ n34855;
  assign n34861 = ~n35477 | ~n35585;
  assign n34857 = ~n35391 | ~P3_EBX_REG_23__SCAN_IN;
  assign n34859 = ~n34857 | ~n34897;
  assign n34860 = ~n34859 | ~n34858;
  assign P3_U2680 = ~n34861 | ~n34860;
  assign n34863 = ~n24513 | ~P3_INSTQUEUE_REG_13__6__SCAN_IN;
  assign n34862 = ~n24516 | ~P3_INSTQUEUE_REG_15__6__SCAN_IN;
  assign n34867 = ~n34863 | ~n34862;
  assign n34865 = ~n24535 | ~P3_INSTQUEUE_REG_8__6__SCAN_IN;
  assign n34864 = ~n35405 | ~P3_INSTQUEUE_REG_3__6__SCAN_IN;
  assign n34866 = ~n34865 | ~n34864;
  assign n34892 = ~n34867 & ~n34866;
  assign n34869 = ~n35328 | ~P3_INSTQUEUE_REG_4__6__SCAN_IN;
  assign n34868 = ~n24470 | ~P3_INSTQUEUE_REG_5__6__SCAN_IN;
  assign n34890 = ~n34869 | ~n34868;
  assign n34871 = ~n24543 | ~P3_INSTQUEUE_REG_7__6__SCAN_IN;
  assign n34870 = ~n34993 | ~P3_INSTQUEUE_REG_6__6__SCAN_IN;
  assign n34876 = ~n34871 | ~n34870;
  assign n34874 = ~n35412 | ~P3_INSTQUEUE_REG_9__6__SCAN_IN;
  assign n34873 = ~n34872 | ~P3_INSTQUEUE_REG_1__6__SCAN_IN;
  assign n34875 = ~n34874 | ~n34873;
  assign n34888 = ~n34876 & ~n34875;
  assign n34878 = ~n35319 | ~P3_INSTQUEUE_REG_11__6__SCAN_IN;
  assign n34877 = ~n35252 | ~P3_INSTQUEUE_REG_0__6__SCAN_IN;
  assign n34882 = ~n34878 | ~n34877;
  assign n34880 = ~n34717 | ~P3_INSTQUEUE_REG_14__6__SCAN_IN;
  assign n34879 = ~n35359 | ~P3_INSTQUEUE_REG_2__6__SCAN_IN;
  assign n34881 = ~n34880 | ~n34879;
  assign n34886 = n34882 | n34881;
  assign n34884 = ~n24451 | ~P3_INSTQUEUE_REG_12__6__SCAN_IN;
  assign n34883 = ~n35366 | ~P3_INSTQUEUE_REG_10__6__SCAN_IN;
  assign n34885 = ~n34884 | ~n34883;
  assign n34887 = ~n34886 & ~n34885;
  assign n34889 = ~n34888 | ~n34887;
  assign n34891 = ~n34890 & ~n34889;
  assign n35592 = ~n34892 | ~n34891;
  assign n34899 = ~n35477 | ~n35592;
  assign n34894 = ~n35477 & ~n34893;
  assign n34896 = n34895 | n34894;
  assign n34898 = ~n34897 | ~n34896;
  assign P3_U2681 = ~n34899 | ~n34898;
  assign n34932 = ~P3_EBX_REG_21__SCAN_IN & ~n34900;
  assign n34902 = ~n35405 | ~P3_INSTQUEUE_REG_3__5__SCAN_IN;
  assign n34901 = ~n24470 | ~P3_INSTQUEUE_REG_5__5__SCAN_IN;
  assign n34906 = ~n34902 | ~n34901;
  assign n34904 = ~n24535 | ~P3_INSTQUEUE_REG_8__5__SCAN_IN;
  assign n34903 = ~n34993 | ~P3_INSTQUEUE_REG_6__5__SCAN_IN;
  assign n34905 = ~n34904 | ~n34903;
  assign n34914 = ~n34906 & ~n34905;
  assign n34908 = ~n24451 | ~P3_INSTQUEUE_REG_12__5__SCAN_IN;
  assign n34907 = ~n35359 | ~P3_INSTQUEUE_REG_2__5__SCAN_IN;
  assign n34912 = ~n34908 | ~n34907;
  assign n34910 = ~n35366 | ~P3_INSTQUEUE_REG_10__5__SCAN_IN;
  assign n34909 = ~n35252 | ~P3_INSTQUEUE_REG_0__5__SCAN_IN;
  assign n34911 = ~n34910 | ~n34909;
  assign n34913 = ~n34912 & ~n34911;
  assign n34930 = ~n34914 | ~n34913;
  assign n34916 = ~n35412 | ~P3_INSTQUEUE_REG_9__5__SCAN_IN;
  assign n34915 = ~n35319 | ~P3_INSTQUEUE_REG_11__5__SCAN_IN;
  assign n34920 = ~n34916 | ~n34915;
  assign n34918 = ~n24513 | ~P3_INSTQUEUE_REG_13__5__SCAN_IN;
  assign n34917 = ~n34872 | ~P3_INSTQUEUE_REG_1__5__SCAN_IN;
  assign n34919 = ~n34918 | ~n34917;
  assign n34928 = ~n34920 & ~n34919;
  assign n34922 = ~n24543 | ~P3_INSTQUEUE_REG_7__5__SCAN_IN;
  assign n34921 = ~n24516 | ~P3_INSTQUEUE_REG_15__5__SCAN_IN;
  assign n34926 = ~n34922 | ~n34921;
  assign n34924 = ~n34717 | ~P3_INSTQUEUE_REG_14__5__SCAN_IN;
  assign n34923 = ~n35328 | ~P3_INSTQUEUE_REG_4__5__SCAN_IN;
  assign n34925 = ~n34924 | ~n34923;
  assign n34927 = ~n34926 & ~n34925;
  assign n34929 = ~n34928 | ~n34927;
  assign n35607 = ~n34930 & ~n34929;
  assign n34931 = ~n35607 & ~n35391;
  assign n34935 = ~n34932 & ~n34931;
  assign n34968 = ~n35477 & ~n34933;
  assign n34934 = ~P3_EBX_REG_21__SCAN_IN | ~n34968;
  assign P3_U2682 = ~n34935 | ~n34934;
  assign n34937 = ~n24513 | ~P3_INSTQUEUE_REG_13__4__SCAN_IN;
  assign n34936 = ~n35319 | ~P3_INSTQUEUE_REG_11__4__SCAN_IN;
  assign n34941 = ~n34937 | ~n34936;
  assign n34939 = ~n34516 | ~P3_INSTQUEUE_REG_7__4__SCAN_IN;
  assign n34938 = ~n24470 | ~P3_INSTQUEUE_REG_5__4__SCAN_IN;
  assign n34940 = ~n34939 | ~n34938;
  assign n34949 = ~n34941 & ~n34940;
  assign n34943 = ~n35252 | ~P3_INSTQUEUE_REG_0__4__SCAN_IN;
  assign n34942 = ~n35359 | ~P3_INSTQUEUE_REG_2__4__SCAN_IN;
  assign n34947 = ~n34943 | ~n34942;
  assign n34945 = ~n24451 | ~P3_INSTQUEUE_REG_12__4__SCAN_IN;
  assign n34944 = ~n35366 | ~P3_INSTQUEUE_REG_10__4__SCAN_IN;
  assign n34946 = ~n34945 | ~n34944;
  assign n34948 = ~n34947 & ~n34946;
  assign n34965 = ~n34949 | ~n34948;
  assign n34951 = ~n34717 | ~P3_INSTQUEUE_REG_14__4__SCAN_IN;
  assign n34950 = ~n34993 | ~P3_INSTQUEUE_REG_6__4__SCAN_IN;
  assign n34955 = ~n34951 | ~n34950;
  assign n34953 = ~n35412 | ~P3_INSTQUEUE_REG_9__4__SCAN_IN;
  assign n34952 = ~n34872 | ~P3_INSTQUEUE_REG_1__4__SCAN_IN;
  assign n34954 = ~n34953 | ~n34952;
  assign n34963 = ~n34955 & ~n34954;
  assign n34957 = ~n24535 | ~P3_INSTQUEUE_REG_8__4__SCAN_IN;
  assign n34956 = ~n24516 | ~P3_INSTQUEUE_REG_15__4__SCAN_IN;
  assign n34961 = ~n34957 | ~n34956;
  assign n34959 = ~n35328 | ~P3_INSTQUEUE_REG_4__4__SCAN_IN;
  assign n34958 = ~n35405 | ~P3_INSTQUEUE_REG_3__4__SCAN_IN;
  assign n34960 = ~n34959 | ~n34958;
  assign n34962 = ~n34961 & ~n34960;
  assign n34964 = ~n34963 | ~n34962;
  assign n35619 = ~n34965 & ~n34964;
  assign n34970 = n35619 | n35391;
  assign n34967 = n34966 | P3_EBX_REG_20__SCAN_IN;
  assign n34969 = ~n34968 | ~n34967;
  assign P3_U2683 = ~n34970 | ~n34969;
  assign n34972 = ~n34971 | ~n35006;
  assign n35005 = ~P3_EBX_REG_19__SCAN_IN & ~n34972;
  assign n34974 = ~n24513 | ~P3_INSTQUEUE_REG_13__3__SCAN_IN;
  assign n34973 = ~n35328 | ~P3_INSTQUEUE_REG_4__3__SCAN_IN;
  assign n34978 = ~n34974 | ~n34973;
  assign n34976 = ~n24451 | ~P3_INSTQUEUE_REG_12__3__SCAN_IN;
  assign n34975 = ~n35359 | ~P3_INSTQUEUE_REG_2__3__SCAN_IN;
  assign n34977 = ~n34976 | ~n34975;
  assign n34986 = ~n34978 & ~n34977;
  assign n34980 = ~n35405 | ~P3_INSTQUEUE_REG_3__3__SCAN_IN;
  assign n34979 = ~n24516 | ~P3_INSTQUEUE_REG_15__3__SCAN_IN;
  assign n34984 = ~n34980 | ~n34979;
  assign n34982 = ~n24535 | ~P3_INSTQUEUE_REG_8__3__SCAN_IN;
  assign n34981 = ~n24543 | ~P3_INSTQUEUE_REG_7__3__SCAN_IN;
  assign n34983 = ~n34982 | ~n34981;
  assign n34985 = ~n34984 & ~n34983;
  assign n35003 = ~n34986 | ~n34985;
  assign n34988 = ~n35412 | ~P3_INSTQUEUE_REG_9__3__SCAN_IN;
  assign n34987 = ~n35319 | ~P3_INSTQUEUE_REG_11__3__SCAN_IN;
  assign n34992 = ~n34988 | ~n34987;
  assign n34990 = ~n34872 | ~P3_INSTQUEUE_REG_1__3__SCAN_IN;
  assign n34989 = ~n24470 | ~P3_INSTQUEUE_REG_5__3__SCAN_IN;
  assign n34991 = ~n34990 | ~n34989;
  assign n35001 = ~n34992 & ~n34991;
  assign n34995 = ~n35366 | ~P3_INSTQUEUE_REG_10__3__SCAN_IN;
  assign n34994 = ~n34993 | ~P3_INSTQUEUE_REG_6__3__SCAN_IN;
  assign n34999 = ~n34995 | ~n34994;
  assign n34997 = ~n34717 | ~P3_INSTQUEUE_REG_14__3__SCAN_IN;
  assign n34996 = ~n35252 | ~P3_INSTQUEUE_REG_0__3__SCAN_IN;
  assign n34998 = ~n34997 | ~n34996;
  assign n35000 = ~n34999 & ~n34998;
  assign n35002 = ~n35001 | ~n35000;
  assign n35629 = ~n35003 & ~n35002;
  assign n35004 = ~n35629 & ~n35487;
  assign n35008 = ~n35005 & ~n35004;
  assign n35043 = ~n35477 & ~n35006;
  assign n35007 = ~P3_EBX_REG_19__SCAN_IN | ~n35043;
  assign P3_U2684 = ~n35008 | ~n35007;
  assign n35010 = ~n35009 | ~n35483;
  assign n35042 = ~P3_EBX_REG_18__SCAN_IN & ~n35010;
  assign n35012 = ~n24451 | ~P3_INSTQUEUE_REG_12__2__SCAN_IN;
  assign n35011 = ~n35328 | ~P3_INSTQUEUE_REG_4__2__SCAN_IN;
  assign n35016 = ~n35012 | ~n35011;
  assign n35014 = ~n34717 | ~P3_INSTQUEUE_REG_14__2__SCAN_IN;
  assign n35013 = ~n24543 | ~P3_INSTQUEUE_REG_7__2__SCAN_IN;
  assign n35015 = ~n35014 | ~n35013;
  assign n35024 = ~n35016 & ~n35015;
  assign n35018 = ~n24470 | ~P3_INSTQUEUE_REG_5__2__SCAN_IN;
  assign n35017 = ~n35359 | ~P3_INSTQUEUE_REG_2__2__SCAN_IN;
  assign n35022 = ~n35018 | ~n35017;
  assign n35020 = ~n24513 | ~P3_INSTQUEUE_REG_13__2__SCAN_IN;
  assign n35019 = ~n35366 | ~P3_INSTQUEUE_REG_10__2__SCAN_IN;
  assign n35021 = ~n35020 | ~n35019;
  assign n35023 = ~n35022 & ~n35021;
  assign n35040 = ~n35024 | ~n35023;
  assign n35026 = ~n24535 | ~P3_INSTQUEUE_REG_8__2__SCAN_IN;
  assign n35025 = ~n34993 | ~P3_INSTQUEUE_REG_6__2__SCAN_IN;
  assign n35030 = ~n35026 | ~n35025;
  assign n35028 = ~n35412 | ~P3_INSTQUEUE_REG_9__2__SCAN_IN;
  assign n35027 = ~n34872 | ~P3_INSTQUEUE_REG_1__2__SCAN_IN;
  assign n35029 = ~n35028 | ~n35027;
  assign n35038 = ~n35030 & ~n35029;
  assign n35032 = ~n35252 | ~P3_INSTQUEUE_REG_0__2__SCAN_IN;
  assign n35031 = ~n24516 | ~P3_INSTQUEUE_REG_15__2__SCAN_IN;
  assign n35036 = ~n35032 | ~n35031;
  assign n35034 = ~n35319 | ~P3_INSTQUEUE_REG_11__2__SCAN_IN;
  assign n35033 = ~n35405 | ~P3_INSTQUEUE_REG_3__2__SCAN_IN;
  assign n35035 = ~n35034 | ~n35033;
  assign n35037 = ~n35036 & ~n35035;
  assign n35039 = ~n35038 | ~n35037;
  assign n35640 = ~n35040 & ~n35039;
  assign n35041 = ~n35640 & ~n35487;
  assign n35045 = ~n35042 & ~n35041;
  assign n35044 = ~P3_EBX_REG_18__SCAN_IN | ~n35043;
  assign P3_U2685 = ~n35045 | ~n35044;
  assign n35047 = n35046 ^ n35078;
  assign n35082 = ~n35047 | ~n35483;
  assign n35049 = ~n24451 | ~P3_INSTQUEUE_REG_12__1__SCAN_IN;
  assign n35048 = ~n35328 | ~P3_INSTQUEUE_REG_4__1__SCAN_IN;
  assign n35053 = ~n35049 | ~n35048;
  assign n35051 = ~n24513 | ~P3_INSTQUEUE_REG_13__1__SCAN_IN;
  assign n35050 = ~n24543 | ~P3_INSTQUEUE_REG_7__1__SCAN_IN;
  assign n35052 = ~n35051 | ~n35050;
  assign n35061 = ~n35053 & ~n35052;
  assign n35055 = ~n24535 | ~P3_INSTQUEUE_REG_8__1__SCAN_IN;
  assign n35054 = ~n34717 | ~P3_INSTQUEUE_REG_14__1__SCAN_IN;
  assign n35059 = ~n35055 | ~n35054;
  assign n35057 = ~n35366 | ~P3_INSTQUEUE_REG_10__1__SCAN_IN;
  assign n35056 = ~n24516 | ~P3_INSTQUEUE_REG_15__1__SCAN_IN;
  assign n35058 = ~n35057 | ~n35056;
  assign n35060 = ~n35059 & ~n35058;
  assign n35077 = ~n35061 | ~n35060;
  assign n35063 = ~n35252 | ~P3_INSTQUEUE_REG_0__1__SCAN_IN;
  assign n35062 = ~n35319 | ~P3_INSTQUEUE_REG_11__1__SCAN_IN;
  assign n35067 = ~n35063 | ~n35062;
  assign n35065 = ~n35412 | ~P3_INSTQUEUE_REG_9__1__SCAN_IN;
  assign n35064 = ~n34872 | ~P3_INSTQUEUE_REG_1__1__SCAN_IN;
  assign n35066 = ~n35065 | ~n35064;
  assign n35075 = ~n35067 & ~n35066;
  assign n35069 = ~n24470 | ~P3_INSTQUEUE_REG_5__1__SCAN_IN;
  assign n35068 = ~n34993 | ~P3_INSTQUEUE_REG_6__1__SCAN_IN;
  assign n35073 = ~n35069 | ~n35068;
  assign n35071 = ~n35405 | ~P3_INSTQUEUE_REG_3__1__SCAN_IN;
  assign n35070 = ~n35359 | ~P3_INSTQUEUE_REG_2__1__SCAN_IN;
  assign n35072 = ~n35071 | ~n35070;
  assign n35074 = ~n35073 & ~n35072;
  assign n35076 = ~n35075 | ~n35074;
  assign n35651 = ~n35077 & ~n35076;
  assign n35080 = ~n35487 & ~n35651;
  assign n35079 = ~n35078 & ~n35394;
  assign n35081 = ~n35080 & ~n35079;
  assign P3_U2686 = ~n35082 | ~n35081;
  assign n35084 = ~n34993 | ~P3_INSTQUEUE_REG_6__0__SCAN_IN;
  assign n35083 = ~n35359 | ~P3_INSTQUEUE_REG_2__0__SCAN_IN;
  assign n35088 = ~n35084 | ~n35083;
  assign n35086 = ~n35405 | ~P3_INSTQUEUE_REG_3__0__SCAN_IN;
  assign n35085 = ~n24516 | ~P3_INSTQUEUE_REG_15__0__SCAN_IN;
  assign n35087 = ~n35086 | ~n35085;
  assign n35096 = ~n35088 & ~n35087;
  assign n35090 = ~n24451 | ~P3_INSTQUEUE_REG_12__0__SCAN_IN;
  assign n35089 = ~n24513 | ~P3_INSTQUEUE_REG_13__0__SCAN_IN;
  assign n35094 = ~n35090 | ~n35089;
  assign n35092 = ~n34717 | ~P3_INSTQUEUE_REG_14__0__SCAN_IN;
  assign n35091 = ~n24543 | ~P3_INSTQUEUE_REG_7__0__SCAN_IN;
  assign n35093 = ~n35092 | ~n35091;
  assign n35095 = ~n35094 & ~n35093;
  assign n35112 = ~n35096 | ~n35095;
  assign n35098 = ~n35366 | ~P3_INSTQUEUE_REG_10__0__SCAN_IN;
  assign n35097 = ~n35319 | ~P3_INSTQUEUE_REG_11__0__SCAN_IN;
  assign n35102 = ~n35098 | ~n35097;
  assign n35100 = ~n35412 | ~P3_INSTQUEUE_REG_9__0__SCAN_IN;
  assign n35099 = ~n34872 | ~P3_INSTQUEUE_REG_1__0__SCAN_IN;
  assign n35101 = ~n35100 | ~n35099;
  assign n35110 = ~n35102 & ~n35101;
  assign n35104 = ~n24535 | ~P3_INSTQUEUE_REG_8__0__SCAN_IN;
  assign n35103 = ~n35252 | ~P3_INSTQUEUE_REG_0__0__SCAN_IN;
  assign n35108 = ~n35104 | ~n35103;
  assign n35106 = ~n35328 | ~P3_INSTQUEUE_REG_4__0__SCAN_IN;
  assign n35105 = ~n24470 | ~P3_INSTQUEUE_REG_5__0__SCAN_IN;
  assign n35107 = ~n35106 | ~n35105;
  assign n35109 = ~n35108 & ~n35107;
  assign n35111 = ~n35110 | ~n35109;
  assign n35664 = ~n35112 & ~n35111;
  assign n35118 = ~n35664 & ~n35487;
  assign n35116 = ~n35113 & ~P3_EBX_REG_16__SCAN_IN;
  assign n35114 = ~P3_EBX_REG_16__SCAN_IN | ~P3_EBX_REG_15__SCAN_IN;
  assign n35115 = ~n35483 | ~n35114;
  assign n35117 = ~n35116 & ~n35115;
  assign n35124 = ~n35118 & ~n35117;
  assign n35357 = ~n35490 & ~n35345;
  assign n35278 = ~n35119 | ~n35357;
  assign n35120 = ~n35279 & ~n35278;
  assign n35189 = ~P3_EBX_REG_12__SCAN_IN | ~n35120;
  assign n35155 = ~n35192 & ~n35189;
  assign n35122 = ~n35155 & ~n35121;
  assign n35123 = ~n35122 | ~n35487;
  assign P3_U2687 = ~n35124 | ~n35123;
  assign n35126 = ~n34516 | ~P3_INSTQUEUE_REG_6__7__SCAN_IN;
  assign n35125 = ~n24470 | ~P3_INSTQUEUE_REG_4__7__SCAN_IN;
  assign n35130 = ~n35126 | ~n35125;
  assign n35128 = ~n24513 | ~P3_INSTQUEUE_REG_12__7__SCAN_IN;
  assign n35127 = ~n35366 | ~P3_INSTQUEUE_REG_9__7__SCAN_IN;
  assign n35129 = ~n35128 | ~n35127;
  assign n35154 = ~n35130 & ~n35129;
  assign n35132 = ~n24300 | ~P3_INSTQUEUE_REG_7__7__SCAN_IN;
  assign n35131 = ~n35319 | ~P3_INSTQUEUE_REG_10__7__SCAN_IN;
  assign n35152 = ~n35132 | ~n35131;
  assign n35134 = ~n35252 | ~P3_INSTQUEUE_REG_15__7__SCAN_IN;
  assign n35133 = ~n35359 | ~P3_INSTQUEUE_REG_1__7__SCAN_IN;
  assign n35138 = ~n35134 | ~n35133;
  assign n35136 = ~n35412 | ~P3_INSTQUEUE_REG_8__7__SCAN_IN;
  assign n35135 = ~n34872 | ~P3_INSTQUEUE_REG_0__7__SCAN_IN;
  assign n35137 = ~n35136 | ~n35135;
  assign n35150 = ~n35138 & ~n35137;
  assign n35140 = ~n34717 | ~P3_INSTQUEUE_REG_13__7__SCAN_IN;
  assign n35139 = ~n35328 | ~P3_INSTQUEUE_REG_3__7__SCAN_IN;
  assign n35144 = ~n35140 | ~n35139;
  assign n35142 = ~n35405 | ~P3_INSTQUEUE_REG_2__7__SCAN_IN;
  assign n35141 = ~n24516 | ~P3_INSTQUEUE_REG_14__7__SCAN_IN;
  assign n35143 = ~n35142 | ~n35141;
  assign n35148 = n35144 | n35143;
  assign n35146 = ~n24451 | ~P3_INSTQUEUE_REG_11__7__SCAN_IN;
  assign n35145 = ~n34993 | ~P3_INSTQUEUE_REG_5__7__SCAN_IN;
  assign n35147 = ~n35146 | ~n35145;
  assign n35149 = ~n35148 & ~n35147;
  assign n35151 = ~n35150 | ~n35149;
  assign n35153 = ~n35152 & ~n35151;
  assign n35672 = ~n35154 | ~n35153;
  assign n35158 = ~n35477 | ~n35672;
  assign n35156 = P3_EBX_REG_15__SCAN_IN ^ n35155;
  assign n35157 = ~n35156 | ~n35487;
  assign P3_U2688 = ~n35158 | ~n35157;
  assign n35160 = ~n24470 | ~P3_INSTQUEUE_REG_4__6__SCAN_IN;
  assign n35159 = ~n34993 | ~P3_INSTQUEUE_REG_5__6__SCAN_IN;
  assign n35164 = ~n35160 | ~n35159;
  assign n35162 = ~n24516 | ~P3_INSTQUEUE_REG_14__6__SCAN_IN;
  assign n35161 = ~n35359 | ~P3_INSTQUEUE_REG_1__6__SCAN_IN;
  assign n35163 = ~n35162 | ~n35161;
  assign n35188 = ~n35164 & ~n35163;
  assign n35168 = ~n34525 & ~n37505;
  assign n35166 = ~n24535 | ~P3_INSTQUEUE_REG_7__6__SCAN_IN;
  assign n35165 = ~n24513 | ~P3_INSTQUEUE_REG_12__6__SCAN_IN;
  assign n35167 = ~n35166 | ~n35165;
  assign n35170 = ~n35168 & ~n35167;
  assign n35169 = ~n35412 | ~P3_INSTQUEUE_REG_8__6__SCAN_IN;
  assign n35186 = ~n35170 | ~n35169;
  assign n35172 = ~n35366 | ~P3_INSTQUEUE_REG_9__6__SCAN_IN;
  assign n35171 = ~n35405 | ~P3_INSTQUEUE_REG_2__6__SCAN_IN;
  assign n35176 = ~n35172 | ~n35171;
  assign n35174 = ~n35328 | ~P3_INSTQUEUE_REG_3__6__SCAN_IN;
  assign n35173 = ~n35319 | ~P3_INSTQUEUE_REG_10__6__SCAN_IN;
  assign n35175 = ~n35174 | ~n35173;
  assign n35184 = ~n35176 & ~n35175;
  assign n35178 = ~n24451 | ~P3_INSTQUEUE_REG_11__6__SCAN_IN;
  assign n35177 = ~n24543 | ~P3_INSTQUEUE_REG_6__6__SCAN_IN;
  assign n35182 = ~n35178 | ~n35177;
  assign n35180 = ~n34717 | ~P3_INSTQUEUE_REG_13__6__SCAN_IN;
  assign n35179 = ~n35252 | ~P3_INSTQUEUE_REG_15__6__SCAN_IN;
  assign n35181 = ~n35180 | ~n35179;
  assign n35183 = ~n35182 & ~n35181;
  assign n35185 = ~n35184 | ~n35183;
  assign n35187 = ~n35186 & ~n35185;
  assign n35682 = ~n35188 | ~n35187;
  assign n35198 = ~n35477 | ~n35682;
  assign n35201 = ~n35487 | ~n35189;
  assign n35196 = ~n35190 & ~n35201;
  assign n35191 = ~P3_EBX_REG_13__SCAN_IN | ~n35200;
  assign n35193 = ~n35191 | ~n35190;
  assign n35194 = ~n35193 | ~n35192;
  assign n35195 = ~n35486 & ~n35194;
  assign n35197 = ~n35196 & ~n35195;
  assign P3_U2689 = ~n35198 | ~n35197;
  assign n35199 = ~P3_EBX_REG_13__SCAN_IN & ~n35486;
  assign n35236 = ~n35200 | ~n35199;
  assign n35202 = ~P3_EBX_REG_13__SCAN_IN;
  assign n35234 = ~n35202 & ~n35201;
  assign n35204 = ~n35328 | ~P3_INSTQUEUE_REG_3__5__SCAN_IN;
  assign n35203 = ~n24516 | ~P3_INSTQUEUE_REG_14__5__SCAN_IN;
  assign n35208 = ~n35204 | ~n35203;
  assign n35206 = ~n35252 | ~P3_INSTQUEUE_REG_15__5__SCAN_IN;
  assign n35205 = ~n24470 | ~P3_INSTQUEUE_REG_4__5__SCAN_IN;
  assign n35207 = ~n35206 | ~n35205;
  assign n35216 = ~n35208 & ~n35207;
  assign n35210 = ~n24451 | ~P3_INSTQUEUE_REG_11__5__SCAN_IN;
  assign n35209 = ~n35359 | ~P3_INSTQUEUE_REG_1__5__SCAN_IN;
  assign n35214 = ~n35210 | ~n35209;
  assign n35212 = ~n34717 | ~P3_INSTQUEUE_REG_13__5__SCAN_IN;
  assign n35211 = ~n34993 | ~P3_INSTQUEUE_REG_5__5__SCAN_IN;
  assign n35213 = ~n35212 | ~n35211;
  assign n35215 = ~n35214 & ~n35213;
  assign n35232 = ~n35216 | ~n35215;
  assign n35218 = ~n24535 | ~P3_INSTQUEUE_REG_7__5__SCAN_IN;
  assign n35217 = ~n35366 | ~P3_INSTQUEUE_REG_9__5__SCAN_IN;
  assign n35222 = ~n35218 | ~n35217;
  assign n35220 = ~n35412 | ~P3_INSTQUEUE_REG_8__5__SCAN_IN;
  assign n35219 = ~n34872 | ~P3_INSTQUEUE_REG_0__5__SCAN_IN;
  assign n35221 = ~n35220 | ~n35219;
  assign n35230 = ~n35222 & ~n35221;
  assign n35224 = ~n35319 | ~P3_INSTQUEUE_REG_10__5__SCAN_IN;
  assign n35223 = ~n24543 | ~P3_INSTQUEUE_REG_6__5__SCAN_IN;
  assign n35228 = ~n35224 | ~n35223;
  assign n35226 = ~n24513 | ~P3_INSTQUEUE_REG_12__5__SCAN_IN;
  assign n35225 = ~n35405 | ~P3_INSTQUEUE_REG_2__5__SCAN_IN;
  assign n35227 = ~n35226 | ~n35225;
  assign n35229 = ~n35228 & ~n35227;
  assign n35231 = ~n35230 | ~n35229;
  assign n35694 = ~n35232 & ~n35231;
  assign n35233 = ~n35694 & ~n35487;
  assign n35235 = ~n35234 & ~n35233;
  assign P3_U2690 = ~n35236 | ~n35235;
  assign n35237 = ~n35278 | ~P3_EBX_REG_12__SCAN_IN;
  assign n35270 = ~n35391 | ~n35237;
  assign n35239 = ~n35366 | ~P3_INSTQUEUE_REG_9__4__SCAN_IN;
  assign n35238 = ~n24516 | ~P3_INSTQUEUE_REG_14__4__SCAN_IN;
  assign n35243 = ~n35239 | ~n35238;
  assign n35241 = ~n24535 | ~P3_INSTQUEUE_REG_7__4__SCAN_IN;
  assign n35240 = ~n35328 | ~P3_INSTQUEUE_REG_3__4__SCAN_IN;
  assign n35242 = ~n35241 | ~n35240;
  assign n35251 = ~n35243 & ~n35242;
  assign n35245 = ~n35319 | ~P3_INSTQUEUE_REG_10__4__SCAN_IN;
  assign n35244 = ~n35359 | ~P3_INSTQUEUE_REG_1__4__SCAN_IN;
  assign n35249 = ~n35245 | ~n35244;
  assign n35247 = ~n24451 | ~P3_INSTQUEUE_REG_11__4__SCAN_IN;
  assign n35246 = ~n24470 | ~P3_INSTQUEUE_REG_4__4__SCAN_IN;
  assign n35248 = ~n35247 | ~n35246;
  assign n35250 = ~n35249 & ~n35248;
  assign n35268 = ~n35251 | ~n35250;
  assign n35254 = ~n35252 | ~P3_INSTQUEUE_REG_15__4__SCAN_IN;
  assign n35253 = ~n35405 | ~P3_INSTQUEUE_REG_2__4__SCAN_IN;
  assign n35258 = ~n35254 | ~n35253;
  assign n35256 = ~n35412 | ~P3_INSTQUEUE_REG_8__4__SCAN_IN;
  assign n35255 = ~n34872 | ~P3_INSTQUEUE_REG_0__4__SCAN_IN;
  assign n35257 = ~n35256 | ~n35255;
  assign n35266 = ~n35258 & ~n35257;
  assign n35260 = ~n24513 | ~P3_INSTQUEUE_REG_12__4__SCAN_IN;
  assign n35259 = ~n34717 | ~P3_INSTQUEUE_REG_13__4__SCAN_IN;
  assign n35264 = ~n35260 | ~n35259;
  assign n35262 = ~n24543 | ~P3_INSTQUEUE_REG_6__4__SCAN_IN;
  assign n35261 = ~n34993 | ~P3_INSTQUEUE_REG_5__4__SCAN_IN;
  assign n35263 = ~n35262 | ~n35261;
  assign n35265 = ~n35264 & ~n35263;
  assign n35267 = ~n35266 | ~n35265;
  assign n35699 = ~n35268 & ~n35267;
  assign n35269 = ~n35477 | ~n35699;
  assign n35277 = ~n35270 | ~n35269;
  assign n35271 = ~n35273 & ~n35279;
  assign n35275 = ~n35271 & ~n35486;
  assign n35274 = ~n35273 | ~n35272;
  assign n35276 = ~n35275 | ~n35274;
  assign P3_U2691 = ~n35277 | ~n35276;
  assign n35280 = n35279 ^ n35278;
  assign n35312 = ~n35280 | ~n35487;
  assign n35282 = ~n35366 | ~P3_INSTQUEUE_REG_9__3__SCAN_IN;
  assign n35281 = ~n24470 | ~P3_INSTQUEUE_REG_4__3__SCAN_IN;
  assign n35286 = ~n35282 | ~n35281;
  assign n35284 = ~n24451 | ~P3_INSTQUEUE_REG_11__3__SCAN_IN;
  assign n35283 = ~n24535 | ~P3_INSTQUEUE_REG_7__3__SCAN_IN;
  assign n35285 = ~n35284 | ~n35283;
  assign n35294 = ~n35286 & ~n35285;
  assign n35288 = ~n24513 | ~P3_INSTQUEUE_REG_12__3__SCAN_IN;
  assign n35287 = ~n24516 | ~P3_INSTQUEUE_REG_14__3__SCAN_IN;
  assign n35292 = ~n35288 | ~n35287;
  assign n35290 = ~n24543 | ~P3_INSTQUEUE_REG_6__3__SCAN_IN;
  assign n35289 = ~n35359 | ~P3_INSTQUEUE_REG_1__3__SCAN_IN;
  assign n35291 = ~n35290 | ~n35289;
  assign n35293 = ~n35292 & ~n35291;
  assign n35310 = ~n35294 | ~n35293;
  assign n35296 = ~n35319 | ~P3_INSTQUEUE_REG_10__3__SCAN_IN;
  assign n35295 = ~n34993 | ~P3_INSTQUEUE_REG_5__3__SCAN_IN;
  assign n35300 = ~n35296 | ~n35295;
  assign n35298 = ~n35412 | ~P3_INSTQUEUE_REG_8__3__SCAN_IN;
  assign n35297 = ~n34872 | ~P3_INSTQUEUE_REG_0__3__SCAN_IN;
  assign n35299 = ~n35298 | ~n35297;
  assign n35308 = ~n35300 & ~n35299;
  assign n35302 = ~n35252 | ~P3_INSTQUEUE_REG_15__3__SCAN_IN;
  assign n35301 = ~n35405 | ~P3_INSTQUEUE_REG_2__3__SCAN_IN;
  assign n35306 = ~n35302 | ~n35301;
  assign n35304 = ~n34717 | ~P3_INSTQUEUE_REG_13__3__SCAN_IN;
  assign n35303 = ~n35328 | ~P3_INSTQUEUE_REG_3__3__SCAN_IN;
  assign n35305 = ~n35304 | ~n35303;
  assign n35307 = ~n35306 & ~n35305;
  assign n35309 = ~n35308 | ~n35307;
  assign n35708 = ~n35310 & ~n35309;
  assign n35311 = n35391 | n35708;
  assign P3_U2692 = ~n35312 | ~n35311;
  assign n35314 = ~n24292 | ~P3_INSTQUEUE_REG_11__2__SCAN_IN;
  assign n35313 = ~n35252 | ~P3_INSTQUEUE_REG_15__2__SCAN_IN;
  assign n35318 = ~n35314 | ~n35313;
  assign n35316 = ~n24513 | ~P3_INSTQUEUE_REG_12__2__SCAN_IN;
  assign n35315 = ~n24516 | ~P3_INSTQUEUE_REG_14__2__SCAN_IN;
  assign n35317 = ~n35316 | ~n35315;
  assign n35327 = ~n35318 & ~n35317;
  assign n35321 = ~n35319 | ~P3_INSTQUEUE_REG_10__2__SCAN_IN;
  assign n35320 = ~n34993 | ~P3_INSTQUEUE_REG_5__2__SCAN_IN;
  assign n35325 = ~n35321 | ~n35320;
  assign n35323 = ~n35405 | ~P3_INSTQUEUE_REG_2__2__SCAN_IN;
  assign n35322 = ~n35359 | ~P3_INSTQUEUE_REG_1__2__SCAN_IN;
  assign n35324 = ~n35323 | ~n35322;
  assign n35326 = ~n35325 & ~n35324;
  assign n35344 = ~n35327 | ~n35326;
  assign n35330 = ~n35366 | ~P3_INSTQUEUE_REG_9__2__SCAN_IN;
  assign n35329 = ~n35328 | ~P3_INSTQUEUE_REG_3__2__SCAN_IN;
  assign n35334 = ~n35330 | ~n35329;
  assign n35332 = ~n35412 | ~P3_INSTQUEUE_REG_8__2__SCAN_IN;
  assign n35331 = ~n34872 | ~P3_INSTQUEUE_REG_0__2__SCAN_IN;
  assign n35333 = ~n35332 | ~n35331;
  assign n35342 = ~n35334 & ~n35333;
  assign n35336 = ~n24535 | ~P3_INSTQUEUE_REG_7__2__SCAN_IN;
  assign n35335 = ~n24470 | ~P3_INSTQUEUE_REG_4__2__SCAN_IN;
  assign n35340 = ~n35336 | ~n35335;
  assign n35338 = ~n34717 | ~P3_INSTQUEUE_REG_13__2__SCAN_IN;
  assign n35337 = ~n24543 | ~P3_INSTQUEUE_REG_6__2__SCAN_IN;
  assign n35339 = ~n35338 | ~n35337;
  assign n35341 = ~n35340 & ~n35339;
  assign n35343 = ~n35342 | ~n35341;
  assign n35717 = ~n35344 & ~n35343;
  assign n35352 = ~n35717 & ~n35391;
  assign n35347 = ~n35346 & ~n35345;
  assign n35350 = ~P3_EBX_REG_10__SCAN_IN & ~n35347;
  assign n35349 = ~n35348 | ~n35483;
  assign n35351 = ~n35350 & ~n35349;
  assign n35356 = ~n35352 & ~n35351;
  assign n35354 = ~n35357 & ~n35353;
  assign n35355 = ~n35354 | ~n35487;
  assign P3_U2693 = ~n35356 | ~n35355;
  assign n35358 = n35357 ^ P3_EBX_REG_9__SCAN_IN;
  assign n35393 = ~n35358 | ~n35487;
  assign n35361 = ~n24535 | ~P3_INSTQUEUE_REG_7__1__SCAN_IN;
  assign n35360 = ~n35359 | ~P3_INSTQUEUE_REG_1__1__SCAN_IN;
  assign n35365 = ~n35361 | ~n35360;
  assign n35363 = ~n24451 | ~P3_INSTQUEUE_REG_11__1__SCAN_IN;
  assign n35362 = ~n24470 | ~P3_INSTQUEUE_REG_4__1__SCAN_IN;
  assign n35364 = ~n35363 | ~n35362;
  assign n35374 = ~n35365 & ~n35364;
  assign n35368 = ~n35366 | ~P3_INSTQUEUE_REG_9__1__SCAN_IN;
  assign n35367 = ~n35252 | ~P3_INSTQUEUE_REG_15__1__SCAN_IN;
  assign n35372 = ~n35368 | ~n35367;
  assign n35370 = ~n35405 | ~P3_INSTQUEUE_REG_2__1__SCAN_IN;
  assign n35369 = ~n34993 | ~P3_INSTQUEUE_REG_5__1__SCAN_IN;
  assign n35371 = ~n35370 | ~n35369;
  assign n35373 = ~n35372 & ~n35371;
  assign n35390 = ~n35374 | ~n35373;
  assign n35376 = ~n34717 | ~P3_INSTQUEUE_REG_13__1__SCAN_IN;
  assign n35375 = ~n24516 | ~P3_INSTQUEUE_REG_14__1__SCAN_IN;
  assign n35380 = ~n35376 | ~n35375;
  assign n35378 = ~n35412 | ~P3_INSTQUEUE_REG_8__1__SCAN_IN;
  assign n35377 = ~n34872 | ~P3_INSTQUEUE_REG_0__1__SCAN_IN;
  assign n35379 = ~n35378 | ~n35377;
  assign n35388 = ~n35380 & ~n35379;
  assign n35382 = ~n24513 | ~P3_INSTQUEUE_REG_12__1__SCAN_IN;
  assign n35381 = ~n34532 | ~P3_INSTQUEUE_REG_10__1__SCAN_IN;
  assign n35386 = ~n35382 | ~n35381;
  assign n35384 = ~n35328 | ~P3_INSTQUEUE_REG_3__1__SCAN_IN;
  assign n35383 = ~n34516 | ~P3_INSTQUEUE_REG_6__1__SCAN_IN;
  assign n35385 = ~n35384 | ~n35383;
  assign n35387 = ~n35386 & ~n35385;
  assign n35389 = ~n35388 | ~n35387;
  assign n35723 = ~n35390 & ~n35389;
  assign n35392 = n35391 | n35723;
  assign P3_U2694 = ~n35393 | ~n35392;
  assign n35454 = ~n35394 | ~n35446;
  assign n35451 = ~n35455 & ~n35454;
  assign n35437 = ~P3_EBX_REG_6__SCAN_IN | ~n35451;
  assign n35434 = ~n35439 & ~n35437;
  assign n35395 = ~P3_EBX_REG_8__SCAN_IN | ~n35487;
  assign n35432 = ~n35434 & ~n35395;
  assign n35398 = ~n35396 | ~P3_INSTQUEUE_REG_9__0__SCAN_IN;
  assign n35397 = ~n35319 | ~P3_INSTQUEUE_REG_10__0__SCAN_IN;
  assign n35402 = ~n35398 | ~n35397;
  assign n35400 = ~n35328 | ~P3_INSTQUEUE_REG_3__0__SCAN_IN;
  assign n35399 = ~n24289 | ~P3_INSTQUEUE_REG_5__0__SCAN_IN;
  assign n35401 = ~n35400 | ~n35399;
  assign n35411 = ~n35402 & ~n35401;
  assign n35404 = ~n34717 | ~P3_INSTQUEUE_REG_13__0__SCAN_IN;
  assign n35403 = ~n34516 | ~P3_INSTQUEUE_REG_6__0__SCAN_IN;
  assign n35409 = ~n35404 | ~n35403;
  assign n35407 = ~n35252 | ~P3_INSTQUEUE_REG_15__0__SCAN_IN;
  assign n35406 = ~n35405 | ~P3_INSTQUEUE_REG_2__0__SCAN_IN;
  assign n35408 = ~n35407 | ~n35406;
  assign n35410 = ~n35409 & ~n35408;
  assign n35430 = ~n35411 | ~n35410;
  assign n35414 = ~n35412 | ~P3_INSTQUEUE_REG_8__0__SCAN_IN;
  assign n35413 = ~n24513 | ~P3_INSTQUEUE_REG_12__0__SCAN_IN;
  assign n35419 = ~n35414 | ~n35413;
  assign n35417 = ~n34872 | ~P3_INSTQUEUE_REG_0__0__SCAN_IN;
  assign n35416 = ~n35415 | ~P3_INSTQUEUE_REG_14__0__SCAN_IN;
  assign n35418 = ~n35417 | ~n35416;
  assign n35428 = ~n35419 & ~n35418;
  assign n35421 = ~n24292 | ~P3_INSTQUEUE_REG_11__0__SCAN_IN;
  assign n35420 = ~n35359 | ~P3_INSTQUEUE_REG_1__0__SCAN_IN;
  assign n35426 = ~n35421 | ~n35420;
  assign n35424 = ~n35422 | ~P3_INSTQUEUE_REG_7__0__SCAN_IN;
  assign n35423 = ~n24470 | ~P3_INSTQUEUE_REG_4__0__SCAN_IN;
  assign n35425 = ~n35424 | ~n35423;
  assign n35427 = ~n35426 & ~n35425;
  assign n35429 = ~n35428 | ~n35427;
  assign n35733 = ~n35430 & ~n35429;
  assign n35431 = ~n35733 & ~n35487;
  assign n35436 = ~n35432 & ~n35431;
  assign n35433 = ~P3_EBX_REG_8__SCAN_IN & ~n37514;
  assign n35435 = ~n35434 | ~n35433;
  assign P3_U2695 = ~n35436 | ~n35435;
  assign n35438 = ~P3_EBX_REG_7__SCAN_IN | ~n35437;
  assign n35443 = ~n35477 & ~n35438;
  assign n35440 = ~n35483 | ~n35439;
  assign n35442 = ~n35441 & ~n35440;
  assign n35445 = ~n35443 & ~n35442;
  assign n35444 = ~n35477 | ~P3_INSTQUEUE_REG_0__7__SCAN_IN;
  assign P3_U2696 = ~n35445 | ~n35444;
  assign n35462 = ~n35446 | ~n35483;
  assign n35448 = ~P3_EBX_REG_5__SCAN_IN | ~n35447;
  assign n35450 = ~n35462 & ~n35448;
  assign n35449 = ~n37505 & ~n35487;
  assign n35453 = ~n35450 & ~n35449;
  assign n35457 = ~n35477 & ~n35451;
  assign n35452 = ~P3_EBX_REG_6__SCAN_IN | ~n35457;
  assign P3_U2697 = ~n35453 | ~n35452;
  assign n35459 = ~P3_INSTQUEUE_REG_0__5__SCAN_IN | ~n35477;
  assign n35456 = ~n35455 | ~n35454;
  assign n35458 = ~n35457 | ~n35456;
  assign P3_U2698 = ~n35459 | ~n35458;
  assign n35465 = ~P3_INSTQUEUE_REG_0__4__SCAN_IN | ~n35477;
  assign n35461 = ~n35487 | ~P3_EBX_REG_4__SCAN_IN;
  assign n35466 = ~n35460 | ~n35483;
  assign n35475 = ~n35466;
  assign n35468 = ~P3_EBX_REG_3__SCAN_IN | ~n35475;
  assign n35463 = ~n35461 | ~n35468;
  assign n35464 = ~n35463 | ~n35462;
  assign P3_U2699 = ~n35465 | ~n35464;
  assign n35471 = ~P3_INSTQUEUE_REG_0__3__SCAN_IN | ~n35477;
  assign n35467 = ~n35487 | ~P3_EBX_REG_3__SCAN_IN;
  assign n35469 = ~n35467 | ~n35466;
  assign n35470 = ~n35469 | ~n35468;
  assign P3_U2700 = ~n35471 | ~n35470;
  assign n35473 = ~n35490 & ~n35472;
  assign n35474 = ~P3_EBX_REG_2__SCAN_IN & ~n35473;
  assign n35476 = ~n35475 & ~n35474;
  assign n35479 = ~n35476 | ~n35487;
  assign n35478 = ~P3_INSTQUEUE_REG_0__2__SCAN_IN | ~n35477;
  assign P3_U2701 = ~n35479 | ~n35478;
  assign n35481 = P3_EBX_REG_1__SCAN_IN & n35490;
  assign n37456 = ~P3_INSTQUEUE_REG_0__1__SCAN_IN;
  assign n35480 = ~n37456 & ~n35487;
  assign n35485 = ~n35481 & ~n35480;
  assign n35484 = ~n35483 | ~n35482;
  assign P3_U2702 = ~n35485 | ~n35484;
  assign n35489 = ~P3_EBX_REG_0__SCAN_IN & ~n35486;
  assign n37446 = ~P3_INSTQUEUE_REG_0__0__SCAN_IN;
  assign n35488 = ~n37446 & ~n35487;
  assign n35492 = ~n35489 & ~n35488;
  assign n35491 = ~P3_EBX_REG_0__SCAN_IN | ~n35490;
  assign P3_U2703 = ~n35492 | ~n35491;
  assign n36013 = ~P3_EAX_REG_29__SCAN_IN;
  assign n36003 = ~P3_EAX_REG_27__SCAN_IN;
  assign n35994 = ~P3_EAX_REG_25__SCAN_IN;
  assign n36098 = ~P3_EAX_REG_15__SCAN_IN;
  assign n35688 = ~P3_EAX_REG_13__SCAN_IN | ~P3_EAX_REG_12__SCAN_IN;
  assign n35493 = ~P3_EAX_REG_14__SCAN_IN | ~n35504;
  assign n35495 = ~P3_EAX_REG_4__SCAN_IN | ~P3_EAX_REG_7__SCAN_IN;
  assign n35494 = ~P3_EAX_REG_2__SCAN_IN | ~P3_EAX_REG_3__SCAN_IN;
  assign n35497 = ~n35495 & ~n35494;
  assign n35741 = ~P3_EAX_REG_1__SCAN_IN | ~P3_EAX_REG_0__SCAN_IN;
  assign n35742 = ~P3_EAX_REG_6__SCAN_IN | ~P3_EAX_REG_5__SCAN_IN;
  assign n35496 = ~n35741 & ~n35742;
  assign n35744 = ~n35497 | ~n35496;
  assign n35687 = ~n36062 & ~n35744;
  assign n35498 = ~P3_EAX_REG_10__SCAN_IN | ~n35687;
  assign n35596 = ~P3_EAX_REG_16__SCAN_IN | ~n35667;
  assign n35597 = ~P3_EAX_REG_18__SCAN_IN | ~P3_EAX_REG_17__SCAN_IN;
  assign n35975 = ~P3_EAX_REG_21__SCAN_IN;
  assign n35964 = ~P3_EAX_REG_19__SCAN_IN;
  assign n35499 = ~n35975 & ~n35964;
  assign n35595 = ~P3_EAX_REG_20__SCAN_IN | ~n35499;
  assign n35500 = ~n35597 & ~n35595;
  assign n35501 = ~P3_EAX_REG_22__SCAN_IN | ~n35500;
  assign n35502 = ~P3_EAX_REG_23__SCAN_IN | ~n35583;
  assign n35571 = ~n37514 & ~n35502;
  assign n35537 = ~P3_EAX_REG_28__SCAN_IN | ~n35535;
  assign n35503 = ~n35514 | ~P3_EAX_REG_30__SCAN_IN;
  assign n35506 = ~n35503 & ~P3_EAX_REG_31__SCAN_IN;
  assign n40548 = ~BUF2_REG_31__SCAN_IN;
  assign n35505 = ~n40548 & ~n35554;
  assign n35510 = ~n35506 & ~n35505;
  assign n36018 = ~P3_EAX_REG_30__SCAN_IN;
  assign n35507 = ~n36018 | ~n35800;
  assign n35508 = ~n35507 | ~n22933;
  assign n35509 = ~n35508 | ~P3_EAX_REG_31__SCAN_IN;
  assign P3_U2704 = ~n35510 | ~n35509;
  assign n35513 = n35752 & n35511;
  assign n35512 = ~n31973 & ~n35554;
  assign n35516 = ~n35513 & ~n35512;
  assign n35515 = ~n35514 | ~n36018;
  assign n35517 = ~n35516 | ~n35515;
  assign n35660 = ~n37494 & ~n35671;
  assign n35518 = ~BUF2_REG_14__SCAN_IN | ~n35660;
  assign P3_U2705 = ~n35519 | ~n35518;
  assign n35526 = ~P3_EAX_REG_29__SCAN_IN & ~n35537;
  assign n35522 = ~n35784 & ~n35520;
  assign n35521 = ~n40515 & ~n35554;
  assign n35524 = ~n35522 & ~n35521;
  assign n35523 = ~BUF2_REG_13__SCAN_IN | ~n35660;
  assign n35525 = ~n35524 | ~n35523;
  assign n35529 = ~n35526 & ~n35525;
  assign n35527 = ~n35789 & ~n36013;
  assign n35528 = ~n35537 | ~n35527;
  assign P3_U2706 = ~n35529 | ~n35528;
  assign n35532 = n35530 | n35784;
  assign n35531 = ~n35660 | ~BUF2_REG_12__SCAN_IN;
  assign n35534 = ~n35532 | ~n35531;
  assign n35533 = ~n32001 & ~n35554;
  assign n35540 = ~n35534 & ~n35533;
  assign n35536 = ~n35671 | ~P3_EAX_REG_28__SCAN_IN;
  assign n35547 = ~n35535;
  assign n35538 = ~n35536 | ~n35547;
  assign n35539 = ~n35538 | ~n35537;
  assign P3_U2707 = ~n35540 | ~n35539;
  assign n35543 = ~n35541 | ~n35752;
  assign n35542 = ~n35660 | ~BUF2_REG_11__SCAN_IN;
  assign n35545 = ~n35543 | ~n35542;
  assign n35544 = ~n32017 & ~n35554;
  assign n35550 = ~n35545 & ~n35544;
  assign n35546 = ~n35671 | ~P3_EAX_REG_27__SCAN_IN;
  assign n35548 = ~n35546 | ~n35558;
  assign n35549 = ~n35548 | ~n35547;
  assign P3_U2708 = ~n35550 | ~n35549;
  assign n35553 = ~n35551 | ~n35752;
  assign n35552 = ~n35660 | ~BUF2_REG_10__SCAN_IN;
  assign n35556 = ~n35553 | ~n35552;
  assign n35555 = ~n32032 & ~n35554;
  assign n35561 = ~n35556 & ~n35555;
  assign n35557 = ~n35671 | ~P3_EAX_REG_26__SCAN_IN;
  assign n35559 = ~n35557 | ~n22908;
  assign n35560 = ~n35559 | ~n35558;
  assign P3_U2709 = ~n35561 | ~n35560;
  assign n35563 = ~n35660 | ~BUF2_REG_9__SCAN_IN;
  assign n35562 = ~n35661 | ~BUF2_REG_25__SCAN_IN;
  assign n35566 = ~n35563 | ~n35562;
  assign n35565 = ~n35784 & ~n35564;
  assign n35570 = ~n35566 & ~n35565;
  assign n35567 = ~n35671 | ~P3_EAX_REG_25__SCAN_IN;
  assign n35568 = ~n35567 | ~n35574;
  assign n35569 = ~n35568 | ~n22908;
  assign P3_U2710 = ~n35570 | ~n35569;
  assign n35573 = ~P3_EAX_REG_24__SCAN_IN | ~n35671;
  assign n35572 = ~n22830;
  assign n35575 = ~n35573 | ~n35572;
  assign n35582 = ~n35575 | ~n35574;
  assign n35577 = ~n35660 | ~BUF2_REG_8__SCAN_IN;
  assign n35576 = ~n35661 | ~BUF2_REG_24__SCAN_IN;
  assign n35580 = ~n35577 | ~n35576;
  assign n35579 = ~n35784 & ~n35578;
  assign n35581 = ~n35580 & ~n35579;
  assign P3_U2711 = ~n35582 | ~n35581;
  assign n35985 = ~P3_EAX_REG_23__SCAN_IN;
  assign n35584 = n35985 ^ n35583;
  assign n35589 = ~n35789 & ~n35584;
  assign n35587 = ~n35585 | ~n35752;
  assign n35586 = ~n35660 | ~BUF2_REG_7__SCAN_IN;
  assign n35588 = ~n35587 | ~n35586;
  assign n35591 = ~n35589 & ~n35588;
  assign n35590 = ~n35661 | ~BUF2_REG_23__SCAN_IN;
  assign P3_U2712 = ~n35591 | ~n35590;
  assign n35594 = ~BUF2_REG_22__SCAN_IN | ~n35661;
  assign n35593 = ~n35752 | ~n35592;
  assign n35604 = ~n35594 | ~n35593;
  assign n35598 = ~P3_EAX_REG_22__SCAN_IN & ~n35595;
  assign n35643 = ~n37514 & ~n35596;
  assign n35654 = ~n35643;
  assign n35602 = ~n35598 | ~n35632;
  assign n35970 = ~P3_EAX_REG_20__SCAN_IN;
  assign n35634 = ~P3_EAX_REG_19__SCAN_IN | ~n35632;
  assign n35612 = ~n35671 | ~n35623;
  assign n35599 = ~n35800 | ~n35975;
  assign n35600 = ~n35612 | ~n35599;
  assign n35601 = ~P3_EAX_REG_22__SCAN_IN | ~n35600;
  assign n35603 = ~n35602 | ~n35601;
  assign n35606 = ~n35604 & ~n35603;
  assign n35605 = ~BUF2_REG_6__SCAN_IN | ~n35660;
  assign P3_U2713 = ~n35606 | ~n35605;
  assign n35611 = ~n35784 & ~n35607;
  assign n35609 = ~BUF2_REG_21__SCAN_IN | ~n35661;
  assign n35608 = ~BUF2_REG_5__SCAN_IN | ~n35660;
  assign n35610 = ~n35609 | ~n35608;
  assign n35616 = ~n35611 & ~n35610;
  assign n35614 = ~n35612 & ~n35975;
  assign n35613 = ~P3_EAX_REG_21__SCAN_IN & ~n35623;
  assign n35615 = ~n35614 & ~n35613;
  assign P3_U2714 = ~n35616 | ~n35615;
  assign n35618 = ~n35660 | ~BUF2_REG_4__SCAN_IN;
  assign n35617 = ~n35661 | ~BUF2_REG_20__SCAN_IN;
  assign n35621 = ~n35618 | ~n35617;
  assign n35620 = ~n35619 & ~n35784;
  assign n35626 = ~n35621 & ~n35620;
  assign n35622 = ~n35671 | ~P3_EAX_REG_20__SCAN_IN;
  assign n35624 = ~n35622 | ~n35634;
  assign n35625 = ~n35624 | ~n35623;
  assign P3_U2715 = ~n35626 | ~n35625;
  assign n35628 = ~n35660 | ~BUF2_REG_3__SCAN_IN;
  assign n35627 = ~n35661 | ~BUF2_REG_19__SCAN_IN;
  assign n35631 = ~n35628 | ~n35627;
  assign n35630 = ~n35629 & ~n35784;
  assign n35637 = ~n35631 & ~n35630;
  assign n35633 = ~n35671 | ~P3_EAX_REG_19__SCAN_IN;
  assign n35645 = ~n35632;
  assign n35635 = ~n35633 | ~n35645;
  assign n35636 = ~n35635 | ~n35634;
  assign P3_U2716 = ~n35637 | ~n35636;
  assign n35639 = ~n35660 | ~BUF2_REG_2__SCAN_IN;
  assign n35638 = ~n35661 | ~BUF2_REG_18__SCAN_IN;
  assign n35642 = ~n35639 | ~n35638;
  assign n35641 = ~n35640 & ~n35784;
  assign n35648 = ~n35642 & ~n35641;
  assign n35644 = ~n35671 | ~P3_EAX_REG_18__SCAN_IN;
  assign n35656 = ~P3_EAX_REG_17__SCAN_IN | ~n35643;
  assign n35646 = ~n35644 | ~n35656;
  assign n35647 = ~n35646 | ~n35645;
  assign P3_U2717 = ~n35648 | ~n35647;
  assign n35650 = ~n35660 | ~BUF2_REG_1__SCAN_IN;
  assign n35649 = ~n35661 | ~BUF2_REG_17__SCAN_IN;
  assign n35653 = ~n35650 | ~n35649;
  assign n35652 = ~n35651 & ~n35784;
  assign n35659 = ~n35653 & ~n35652;
  assign n35655 = ~n35671 | ~P3_EAX_REG_17__SCAN_IN;
  assign n35657 = ~n35655 | ~n35654;
  assign n35658 = ~n35657 | ~n35656;
  assign P3_U2718 = ~n35659 | ~n35658;
  assign n35663 = ~n35660 | ~BUF2_REG_0__SCAN_IN;
  assign n35662 = ~n35661 | ~BUF2_REG_16__SCAN_IN;
  assign n35666 = ~n35663 | ~n35662;
  assign n35665 = ~n35664 & ~n35784;
  assign n35670 = ~n35666 & ~n35665;
  assign n35947 = ~P3_EAX_REG_16__SCAN_IN;
  assign n35668 = ~n35947 ^ n35667;
  assign n35669 = ~n35668 | ~n35671;
  assign P3_U2719 = ~n35670 | ~n35669;
  assign n35681 = ~n35671 | ~n35677;
  assign n35676 = ~n35681 & ~n36098;
  assign n35674 = ~BUF2_REG_15__SCAN_IN | ~n35807;
  assign n35673 = ~n35752 | ~n35672;
  assign n35675 = ~n35674 | ~n35673;
  assign n35680 = ~n35676 & ~n35675;
  assign n35678 = ~n37514 & ~n35677;
  assign n35679 = ~n35678 | ~n36098;
  assign P3_U2720 = ~n35680 | ~n35679;
  assign n36092 = ~P3_EAX_REG_14__SCAN_IN;
  assign n35686 = ~n35681 & ~n36092;
  assign n35684 = ~BUF2_REG_14__SCAN_IN | ~n35807;
  assign n35683 = ~n35752 | ~n35682;
  assign n35685 = ~n35684 | ~n35683;
  assign n35690 = ~n35686 & ~n35685;
  assign n36072 = ~P3_EAX_REG_10__SCAN_IN;
  assign n35724 = ~P3_EAX_REG_9__SCAN_IN | ~n35726;
  assign n35710 = ~n36072 & ~n35724;
  assign n35700 = ~P3_EAX_REG_11__SCAN_IN | ~n35710;
  assign n35693 = ~n35688 & ~n35700;
  assign n35689 = ~n35693 | ~n36092;
  assign P3_U2721 = ~n35690 | ~n35689;
  assign n36082 = ~P3_EAX_REG_12__SCAN_IN;
  assign n35703 = ~n36082 & ~n35700;
  assign n36087 = ~P3_EAX_REG_13__SCAN_IN;
  assign n35691 = ~n35789 & ~n36087;
  assign n35692 = ~n35703 & ~n35691;
  assign n35696 = ~n35693 & ~n35692;
  assign n35695 = ~n35784 & ~n35694;
  assign n35698 = ~n35696 & ~n35695;
  assign n35697 = ~BUF2_REG_13__SCAN_IN | ~n35807;
  assign P3_U2722 = ~n35698 | ~n35697;
  assign n35705 = ~n35699 & ~n35784;
  assign n35712 = ~n35700;
  assign n35701 = ~n35789 & ~n36082;
  assign n35702 = ~n35712 & ~n35701;
  assign n35704 = ~n35703 & ~n35702;
  assign n35707 = ~n35705 & ~n35704;
  assign n35706 = ~n35807 | ~BUF2_REG_12__SCAN_IN;
  assign P3_U2723 = ~n35707 | ~n35706;
  assign n35714 = ~n35708 & ~n35784;
  assign n36077 = ~P3_EAX_REG_11__SCAN_IN;
  assign n35709 = ~n35789 & ~n36077;
  assign n35711 = ~n35710 & ~n35709;
  assign n35713 = ~n35712 & ~n35711;
  assign n35716 = ~n35714 & ~n35713;
  assign n35715 = ~n35807 | ~BUF2_REG_11__SCAN_IN;
  assign P3_U2724 = ~n35716 | ~n35715;
  assign n35720 = ~n35717 & ~n35784;
  assign n35718 = P3_EAX_REG_10__SCAN_IN ^ n35724;
  assign n35719 = ~n35789 & ~n35718;
  assign n35722 = ~n35720 & ~n35719;
  assign n35721 = ~n35807 | ~BUF2_REG_10__SCAN_IN;
  assign P3_U2725 = ~n35722 | ~n35721;
  assign n35730 = ~n35723 & ~n35784;
  assign n35728 = ~n35724;
  assign n36067 = ~P3_EAX_REG_9__SCAN_IN;
  assign n35725 = ~n35789 & ~n36067;
  assign n35727 = ~n35726 & ~n35725;
  assign n35729 = ~n35728 & ~n35727;
  assign n35732 = ~n35730 & ~n35729;
  assign n35731 = ~n35807 | ~BUF2_REG_9__SCAN_IN;
  assign P3_U2726 = ~n35732 | ~n35731;
  assign n35738 = ~n35733 & ~n35784;
  assign n35734 = n36062 ^ n35744;
  assign n35736 = ~n35734 | ~n35800;
  assign n35735 = ~P3_EAX_REG_8__SCAN_IN | ~n35799;
  assign n35737 = ~n35736 | ~n35735;
  assign n35740 = ~n35738 & ~n35737;
  assign n35739 = ~n35807 | ~BUF2_REG_8__SCAN_IN;
  assign P3_U2727 = ~n35740 | ~n35739;
  assign n35749 = ~n37212 & ~n35784;
  assign n36037 = ~P3_EAX_REG_3__SCAN_IN;
  assign n35791 = ~n35741 & ~n35745;
  assign n35778 = ~P3_EAX_REG_2__SCAN_IN | ~n35791;
  assign n35781 = ~n36037 & ~n35778;
  assign n35762 = ~P3_EAX_REG_4__SCAN_IN | ~n35781;
  assign n35756 = ~n35742 & ~n35762;
  assign n36057 = ~P3_EAX_REG_7__SCAN_IN;
  assign n35743 = ~n35789 & ~n36057;
  assign n35747 = ~n35756 & ~n35743;
  assign n35746 = ~n35745 & ~n35744;
  assign n35748 = ~n35747 & ~n35746;
  assign n35751 = ~n35749 & ~n35748;
  assign n35750 = ~n35807 | ~BUF2_REG_7__SCAN_IN;
  assign P3_U2728 = ~n35751 | ~n35750;
  assign n35758 = n35753 & n35752;
  assign n36047 = ~P3_EAX_REG_5__SCAN_IN;
  assign n35765 = ~n36047 & ~n35762;
  assign n36052 = ~P3_EAX_REG_6__SCAN_IN;
  assign n35754 = ~n35789 & ~n36052;
  assign n35755 = ~n35765 & ~n35754;
  assign n35757 = ~n35756 & ~n35755;
  assign n35760 = ~n35758 & ~n35757;
  assign n35759 = ~n35807 | ~BUF2_REG_6__SCAN_IN;
  assign P3_U2729 = ~n35760 | ~n35759;
  assign n35767 = ~n35761 & ~n35784;
  assign n35772 = ~n35762;
  assign n35763 = ~n35789 & ~n36047;
  assign n35764 = ~n35772 & ~n35763;
  assign n35766 = ~n35765 & ~n35764;
  assign n35769 = ~n35767 & ~n35766;
  assign n35768 = ~n35807 | ~BUF2_REG_5__SCAN_IN;
  assign P3_U2730 = ~n35769 | ~n35768;
  assign n36042 = ~P3_EAX_REG_4__SCAN_IN;
  assign n35770 = ~n35789 & ~n36042;
  assign n35771 = ~n35781 & ~n35770;
  assign n35775 = ~n35772 & ~n35771;
  assign n35774 = ~n35784 & ~n35773;
  assign n35777 = ~n35775 & ~n35774;
  assign n35776 = ~n35807 | ~BUF2_REG_4__SCAN_IN;
  assign P3_U2731 = ~n35777 | ~n35776;
  assign n35793 = ~n35778;
  assign n35779 = ~n35789 & ~n36037;
  assign n35780 = ~n35793 & ~n35779;
  assign n35786 = ~n35781 & ~n35780;
  assign n35783 = ~n35782;
  assign n35785 = ~n35784 & ~n35783;
  assign n35788 = ~n35786 & ~n35785;
  assign n35787 = ~n35807 | ~BUF2_REG_3__SCAN_IN;
  assign P3_U2732 = ~n35788 | ~n35787;
  assign n36032 = ~P3_EAX_REG_2__SCAN_IN;
  assign n35790 = ~n35789 & ~n36032;
  assign n35792 = ~n35791 & ~n35790;
  assign n35796 = ~n35793 & ~n35792;
  assign n35795 = ~n35784 & ~n35794;
  assign n35798 = ~n35796 & ~n35795;
  assign n35797 = ~n35807 | ~BUF2_REG_2__SCAN_IN;
  assign P3_U2733 = ~n35798 | ~n35797;
  assign n35803 = ~P3_EAX_REG_1__SCAN_IN | ~n35799;
  assign n36027 = ~P3_EAX_REG_1__SCAN_IN;
  assign n35801 = ~n36027 ^ P3_EAX_REG_0__SCAN_IN;
  assign n35802 = ~n35801 | ~n35800;
  assign n35806 = ~n35803 | ~n35802;
  assign n35805 = ~n35784 & ~n35804;
  assign n35809 = ~n35806 & ~n35805;
  assign n35808 = ~n35807 | ~BUF2_REG_1__SCAN_IN;
  assign P3_U2734 = ~n35809 | ~n35808;
  assign n35936 = ~n37396 & ~P3_STATE2_REG_0__SCAN_IN;
  assign P3_U2736 = n35940 & P3_DATAO_REG_31__SCAN_IN;
  assign n35814 = ~n35940 | ~P3_DATAO_REG_30__SCAN_IN;
  assign n35813 = ~P3_UWORD_REG_14__SCAN_IN | ~n39106;
  assign n35817 = n35814 & n35813;
  assign n35816 = ~P3_EAX_REG_30__SCAN_IN | ~n35872;
  assign P3_U2737 = ~n35817 | ~n35816;
  assign n35819 = ~n35940 | ~P3_DATAO_REG_29__SCAN_IN;
  assign n35818 = ~P3_UWORD_REG_13__SCAN_IN | ~n39106;
  assign n35821 = n35819 & n35818;
  assign n35820 = ~P3_EAX_REG_29__SCAN_IN | ~n35872;
  assign P3_U2738 = ~n35821 | ~n35820;
  assign n35823 = ~P3_DATAO_REG_28__SCAN_IN | ~n35909;
  assign n35822 = ~P3_UWORD_REG_12__SCAN_IN | ~n39106;
  assign n35825 = n35823 & n35822;
  assign n35824 = ~P3_EAX_REG_28__SCAN_IN | ~n35872;
  assign P3_U2739 = ~n35825 | ~n35824;
  assign n35827 = ~n35940 | ~P3_DATAO_REG_27__SCAN_IN;
  assign n35826 = ~P3_UWORD_REG_11__SCAN_IN | ~n39106;
  assign n35829 = n35827 & n35826;
  assign n35828 = ~P3_EAX_REG_27__SCAN_IN | ~n35872;
  assign P3_U2740 = ~n35829 | ~n35828;
  assign n35831 = ~n35940 | ~P3_DATAO_REG_26__SCAN_IN;
  assign n35830 = ~P3_UWORD_REG_10__SCAN_IN | ~n39106;
  assign n35833 = n35831 & n35830;
  assign n35832 = ~P3_EAX_REG_26__SCAN_IN | ~n35872;
  assign P3_U2741 = ~n35833 | ~n35832;
  assign n35835 = ~n35940 | ~P3_DATAO_REG_25__SCAN_IN;
  assign n35834 = ~P3_UWORD_REG_9__SCAN_IN | ~n39106;
  assign n35837 = n35835 & n35834;
  assign n35836 = ~P3_EAX_REG_25__SCAN_IN | ~n35872;
  assign P3_U2742 = ~n35837 | ~n35836;
  assign n35839 = ~n35940 | ~P3_DATAO_REG_24__SCAN_IN;
  assign n35838 = ~P3_UWORD_REG_8__SCAN_IN | ~n39106;
  assign n35841 = n35839 & n35838;
  assign n35840 = ~P3_EAX_REG_24__SCAN_IN | ~n35872;
  assign P3_U2743 = ~n35841 | ~n35840;
  assign n35843 = ~n35940 | ~P3_DATAO_REG_23__SCAN_IN;
  assign n35842 = ~P3_UWORD_REG_7__SCAN_IN | ~n35936;
  assign n35845 = n35843 & n35842;
  assign n35844 = ~P3_EAX_REG_23__SCAN_IN | ~n35872;
  assign P3_U2744 = ~n35845 | ~n35844;
  assign n35847 = ~n35909 | ~P3_DATAO_REG_22__SCAN_IN;
  assign n35846 = ~P3_UWORD_REG_6__SCAN_IN | ~n39106;
  assign n35849 = n35847 & n35846;
  assign n35848 = ~P3_EAX_REG_22__SCAN_IN | ~n35872;
  assign P3_U2745 = ~n35849 | ~n35848;
  assign n35851 = ~n35909 | ~P3_DATAO_REG_21__SCAN_IN;
  assign n35850 = ~P3_UWORD_REG_5__SCAN_IN | ~n39106;
  assign n35853 = n35851 & n35850;
  assign n35852 = ~P3_EAX_REG_21__SCAN_IN | ~n35872;
  assign P3_U2746 = ~n35853 | ~n35852;
  assign n35855 = ~P3_DATAO_REG_20__SCAN_IN | ~n35909;
  assign n35854 = ~P3_UWORD_REG_4__SCAN_IN | ~n39106;
  assign n35857 = n35855 & n35854;
  assign n35856 = ~P3_EAX_REG_20__SCAN_IN | ~n35872;
  assign P3_U2747 = ~n35857 | ~n35856;
  assign n35859 = ~P3_DATAO_REG_19__SCAN_IN | ~n35909;
  assign n35858 = ~P3_UWORD_REG_3__SCAN_IN | ~n39106;
  assign n35861 = n35859 & n35858;
  assign n35860 = ~P3_EAX_REG_19__SCAN_IN | ~n35872;
  assign P3_U2748 = ~n35861 | ~n35860;
  assign n35863 = ~n35909 | ~P3_DATAO_REG_18__SCAN_IN;
  assign n35862 = ~P3_UWORD_REG_2__SCAN_IN | ~n39106;
  assign n35865 = n35863 & n35862;
  assign n35864 = ~P3_EAX_REG_18__SCAN_IN | ~n35872;
  assign P3_U2749 = ~n35865 | ~n35864;
  assign n35867 = ~n35909 | ~P3_DATAO_REG_17__SCAN_IN;
  assign n35866 = ~P3_UWORD_REG_1__SCAN_IN | ~n39106;
  assign n35869 = n35867 & n35866;
  assign n35868 = ~P3_EAX_REG_17__SCAN_IN | ~n35872;
  assign P3_U2750 = ~n35869 | ~n35868;
  assign n35871 = ~n35909 | ~P3_DATAO_REG_16__SCAN_IN;
  assign n35870 = ~P3_UWORD_REG_0__SCAN_IN | ~n39106;
  assign n35874 = n35871 & n35870;
  assign n35873 = ~P3_EAX_REG_16__SCAN_IN | ~n35872;
  assign P3_U2751 = ~n35874 | ~n35873;
  assign n35876 = ~P3_LWORD_REG_15__SCAN_IN | ~n39106;
  assign n35875 = ~n35937 | ~P3_EAX_REG_15__SCAN_IN;
  assign n35878 = n35876 & n35875;
  assign n35877 = ~n35940 | ~P3_DATAO_REG_15__SCAN_IN;
  assign P3_U2752 = ~n35878 | ~n35877;
  assign n35880 = ~P3_LWORD_REG_14__SCAN_IN | ~n39106;
  assign n35879 = ~n35937 | ~P3_EAX_REG_14__SCAN_IN;
  assign n35882 = n35880 & n35879;
  assign n35881 = ~n35940 | ~P3_DATAO_REG_14__SCAN_IN;
  assign P3_U2753 = ~n35882 | ~n35881;
  assign n35884 = ~P3_LWORD_REG_13__SCAN_IN | ~n39106;
  assign n35883 = ~n35937 | ~P3_EAX_REG_13__SCAN_IN;
  assign n35886 = n35884 & n35883;
  assign n35885 = ~n35940 | ~P3_DATAO_REG_13__SCAN_IN;
  assign P3_U2754 = ~n35886 | ~n35885;
  assign n35888 = ~P3_LWORD_REG_12__SCAN_IN | ~n39106;
  assign n35887 = ~n35937 | ~P3_EAX_REG_12__SCAN_IN;
  assign n35890 = n35888 & n35887;
  assign n35889 = ~n35940 | ~P3_DATAO_REG_12__SCAN_IN;
  assign P3_U2755 = ~n35890 | ~n35889;
  assign n35892 = ~P3_LWORD_REG_11__SCAN_IN | ~n39106;
  assign n35891 = ~n35937 | ~P3_EAX_REG_11__SCAN_IN;
  assign n35894 = n35892 & n35891;
  assign n35893 = ~n35940 | ~P3_DATAO_REG_11__SCAN_IN;
  assign P3_U2756 = ~n35894 | ~n35893;
  assign n35896 = ~P3_LWORD_REG_10__SCAN_IN | ~n35936;
  assign n35895 = ~n35937 | ~P3_EAX_REG_10__SCAN_IN;
  assign n35898 = n35896 & n35895;
  assign n35897 = ~n35940 | ~P3_DATAO_REG_10__SCAN_IN;
  assign P3_U2757 = ~n35898 | ~n35897;
  assign n35900 = ~P3_LWORD_REG_9__SCAN_IN | ~n35936;
  assign n35899 = ~n35937 | ~P3_EAX_REG_9__SCAN_IN;
  assign n35902 = n35900 & n35899;
  assign n35901 = ~n35909 | ~P3_DATAO_REG_9__SCAN_IN;
  assign P3_U2758 = ~n35902 | ~n35901;
  assign n35904 = ~P3_LWORD_REG_8__SCAN_IN | ~n35936;
  assign n35903 = ~n35937 | ~P3_EAX_REG_8__SCAN_IN;
  assign n35906 = n35904 & n35903;
  assign n35905 = ~n35909 | ~P3_DATAO_REG_8__SCAN_IN;
  assign P3_U2759 = ~n35906 | ~n35905;
  assign n35908 = ~P3_LWORD_REG_7__SCAN_IN | ~n35936;
  assign n35907 = ~n35937 | ~P3_EAX_REG_7__SCAN_IN;
  assign n35911 = n35908 & n35907;
  assign n35910 = ~n35909 | ~P3_DATAO_REG_7__SCAN_IN;
  assign P3_U2760 = ~n35911 | ~n35910;
  assign n35913 = ~P3_LWORD_REG_6__SCAN_IN | ~n39106;
  assign n35912 = ~n35937 | ~P3_EAX_REG_6__SCAN_IN;
  assign n35915 = n35913 & n35912;
  assign n35914 = ~n35940 | ~P3_DATAO_REG_6__SCAN_IN;
  assign P3_U2761 = ~n35915 | ~n35914;
  assign n35917 = ~P3_LWORD_REG_5__SCAN_IN | ~n35936;
  assign n35916 = ~n35937 | ~P3_EAX_REG_5__SCAN_IN;
  assign n35919 = n35917 & n35916;
  assign n35918 = ~n35940 | ~P3_DATAO_REG_5__SCAN_IN;
  assign P3_U2762 = ~n35919 | ~n35918;
  assign n35921 = ~P3_LWORD_REG_4__SCAN_IN | ~n35936;
  assign n35920 = ~n35937 | ~P3_EAX_REG_4__SCAN_IN;
  assign n35923 = n35921 & n35920;
  assign n35922 = ~n35940 | ~P3_DATAO_REG_4__SCAN_IN;
  assign P3_U2763 = ~n35923 | ~n35922;
  assign n35925 = ~P3_LWORD_REG_3__SCAN_IN | ~n35936;
  assign n35924 = ~n35937 | ~P3_EAX_REG_3__SCAN_IN;
  assign n35927 = n35925 & n35924;
  assign n35926 = ~n35940 | ~P3_DATAO_REG_3__SCAN_IN;
  assign P3_U2764 = ~n35927 | ~n35926;
  assign n35929 = ~P3_LWORD_REG_2__SCAN_IN | ~n35936;
  assign n35928 = ~n35937 | ~P3_EAX_REG_2__SCAN_IN;
  assign n35931 = n35929 & n35928;
  assign n35930 = ~n35940 | ~P3_DATAO_REG_2__SCAN_IN;
  assign P3_U2765 = ~n35931 | ~n35930;
  assign n35933 = ~P3_LWORD_REG_1__SCAN_IN | ~n35936;
  assign n35932 = ~n35937 | ~P3_EAX_REG_1__SCAN_IN;
  assign n35935 = n35933 & n35932;
  assign n35934 = ~n35940 | ~P3_DATAO_REG_1__SCAN_IN;
  assign P3_U2766 = ~n35935 | ~n35934;
  assign n35939 = ~P3_LWORD_REG_0__SCAN_IN | ~n35936;
  assign n35938 = ~n35937 | ~P3_EAX_REG_0__SCAN_IN;
  assign n35942 = n35939 & n35938;
  assign n35941 = ~n35940 | ~P3_DATAO_REG_0__SCAN_IN;
  assign P3_U2767 = ~n35942 | ~n35941;
  assign n35946 = ~n35944 | ~n38797;
  assign n36103 = ~n35946 | ~n35945;
  assign n35952 = ~P3_UWORD_REG_0__SCAN_IN | ~n36103;
  assign n36097 = ~n37453 | ~n35966;
  assign n35950 = ~n36097 & ~n35947;
  assign n35949 = ~BUF2_REG_0__SCAN_IN;
  assign n36023 = ~n35949 & ~n36099;
  assign n35951 = ~n35950 & ~n36023;
  assign P3_U2768 = ~n35952 | ~n35951;
  assign n35953 = ~BUF2_REG_1__SCAN_IN;
  assign n36028 = ~n35953 & ~n36099;
  assign n35954 = ~P3_EAX_REG_17__SCAN_IN;
  assign n35955 = ~n35954 & ~n36097;
  assign n35957 = ~n36028 & ~n35955;
  assign n35956 = ~P3_UWORD_REG_1__SCAN_IN | ~n36103;
  assign P3_U2769 = ~n35957 | ~n35956;
  assign n35958 = ~BUF2_REG_2__SCAN_IN;
  assign n36033 = ~n35958 & ~n36099;
  assign n35959 = ~P3_EAX_REG_18__SCAN_IN;
  assign n35960 = ~n35959 & ~n36097;
  assign n35962 = ~n36033 & ~n35960;
  assign n35961 = ~P3_UWORD_REG_2__SCAN_IN | ~n36103;
  assign P3_U2770 = ~n35962 | ~n35961;
  assign n35963 = ~BUF2_REG_3__SCAN_IN;
  assign n36038 = ~n35963 & ~n36099;
  assign n35965 = ~n35964 & ~n36097;
  assign n35968 = ~n36038 & ~n35965;
  assign n35967 = ~P3_UWORD_REG_3__SCAN_IN | ~n36103;
  assign P3_U2771 = ~n35968 | ~n35967;
  assign n35969 = ~BUF2_REG_4__SCAN_IN;
  assign n36043 = ~n35969 & ~n36099;
  assign n35971 = ~n35970 & ~n36097;
  assign n35973 = ~n36043 & ~n35971;
  assign n35972 = ~P3_UWORD_REG_4__SCAN_IN | ~n36103;
  assign P3_U2772 = ~n35973 | ~n35972;
  assign n35974 = ~BUF2_REG_5__SCAN_IN;
  assign n36048 = ~n35974 & ~n36099;
  assign n35976 = ~n35975 & ~n36097;
  assign n35978 = ~n36048 & ~n35976;
  assign n35977 = ~P3_UWORD_REG_5__SCAN_IN | ~n36103;
  assign P3_U2773 = ~n35978 | ~n35977;
  assign n35979 = ~BUF2_REG_6__SCAN_IN;
  assign n36053 = ~n35979 & ~n36099;
  assign n35980 = ~P3_EAX_REG_22__SCAN_IN;
  assign n35981 = ~n35980 & ~n36097;
  assign n35983 = ~n36053 & ~n35981;
  assign n35982 = ~P3_UWORD_REG_6__SCAN_IN | ~n36103;
  assign P3_U2774 = ~n35983 | ~n35982;
  assign n35984 = ~BUF2_REG_7__SCAN_IN;
  assign n36058 = ~n35984 & ~n36099;
  assign n35986 = ~n35985 & ~n36097;
  assign n35988 = ~n36058 & ~n35986;
  assign n35987 = ~P3_UWORD_REG_7__SCAN_IN | ~n36103;
  assign P3_U2775 = ~n35988 | ~n35987;
  assign n35989 = ~BUF2_REG_8__SCAN_IN;
  assign n36063 = ~n35989 & ~n36099;
  assign n35990 = ~n23363 & ~n36097;
  assign n35992 = ~n36063 & ~n35990;
  assign n35991 = ~P3_UWORD_REG_8__SCAN_IN | ~n36103;
  assign P3_U2776 = ~n35992 | ~n35991;
  assign n35993 = ~BUF2_REG_9__SCAN_IN;
  assign n36068 = ~n35993 & ~n36099;
  assign n35995 = ~n35994 & ~n36097;
  assign n35997 = ~n36068 & ~n35995;
  assign n35996 = ~P3_UWORD_REG_9__SCAN_IN | ~n36103;
  assign P3_U2777 = ~n35997 | ~n35996;
  assign n35998 = ~BUF2_REG_10__SCAN_IN;
  assign n36073 = ~n35998 & ~n36099;
  assign n35999 = ~n23364 & ~n36097;
  assign n36001 = ~n36073 & ~n35999;
  assign n36000 = ~P3_UWORD_REG_10__SCAN_IN | ~n36103;
  assign P3_U2778 = ~n36001 | ~n36000;
  assign n36002 = ~BUF2_REG_11__SCAN_IN;
  assign n36078 = ~n36002 & ~n36099;
  assign n36004 = ~n36003 & ~n36097;
  assign n36006 = ~n36078 & ~n36004;
  assign n36005 = ~P3_UWORD_REG_11__SCAN_IN | ~n36103;
  assign P3_U2779 = ~n36006 | ~n36005;
  assign n36007 = ~BUF2_REG_12__SCAN_IN;
  assign n36083 = ~n36007 & ~n36099;
  assign n36008 = ~P3_EAX_REG_28__SCAN_IN;
  assign n36009 = ~n36008 & ~n36097;
  assign n36011 = ~n36083 & ~n36009;
  assign n36010 = ~P3_UWORD_REG_12__SCAN_IN | ~n36103;
  assign P3_U2780 = ~n36011 | ~n36010;
  assign n36012 = ~BUF2_REG_13__SCAN_IN;
  assign n36088 = ~n36012 & ~n36099;
  assign n36014 = ~n36013 & ~n36097;
  assign n36016 = ~n36088 & ~n36014;
  assign n36015 = ~P3_UWORD_REG_13__SCAN_IN | ~n36103;
  assign P3_U2781 = ~n36016 | ~n36015;
  assign n36017 = ~BUF2_REG_14__SCAN_IN;
  assign n36093 = ~n36017 & ~n36099;
  assign n36019 = ~n36018 & ~n36097;
  assign n36021 = ~n36093 & ~n36019;
  assign n36020 = ~P3_UWORD_REG_14__SCAN_IN | ~n36103;
  assign P3_U2782 = ~n36021 | ~n36020;
  assign n36022 = ~P3_EAX_REG_0__SCAN_IN;
  assign n36024 = ~n36022 & ~n36097;
  assign n36026 = ~n36024 & ~n36023;
  assign n36025 = ~P3_LWORD_REG_0__SCAN_IN | ~n36103;
  assign P3_U2783 = ~n36026 | ~n36025;
  assign n36029 = ~n36027 & ~n36097;
  assign n36031 = ~n36029 & ~n36028;
  assign n36030 = ~P3_LWORD_REG_1__SCAN_IN | ~n36103;
  assign P3_U2784 = ~n36031 | ~n36030;
  assign n36034 = ~n36032 & ~n36097;
  assign n36036 = ~n36034 & ~n36033;
  assign n36035 = ~P3_LWORD_REG_2__SCAN_IN | ~n36103;
  assign P3_U2785 = ~n36036 | ~n36035;
  assign n36039 = ~n36037 & ~n36097;
  assign n36041 = ~n36039 & ~n36038;
  assign n36040 = ~P3_LWORD_REG_3__SCAN_IN | ~n36103;
  assign P3_U2786 = ~n36041 | ~n36040;
  assign n36044 = ~n36042 & ~n36097;
  assign n36046 = ~n36044 & ~n36043;
  assign n36045 = ~P3_LWORD_REG_4__SCAN_IN | ~n36103;
  assign P3_U2787 = ~n36046 | ~n36045;
  assign n36049 = ~n36047 & ~n36097;
  assign n36051 = ~n36049 & ~n36048;
  assign n36050 = ~P3_LWORD_REG_5__SCAN_IN | ~n36103;
  assign P3_U2788 = ~n36051 | ~n36050;
  assign n36054 = ~n36052 & ~n36097;
  assign n36056 = ~n36054 & ~n36053;
  assign n36055 = ~P3_LWORD_REG_6__SCAN_IN | ~n36103;
  assign P3_U2789 = ~n36056 | ~n36055;
  assign n36059 = ~n36057 & ~n36097;
  assign n36061 = ~n36059 & ~n36058;
  assign n36060 = ~P3_LWORD_REG_7__SCAN_IN | ~n36103;
  assign P3_U2790 = ~n36061 | ~n36060;
  assign n36064 = ~n36062 & ~n36097;
  assign n36066 = ~n36064 & ~n36063;
  assign n36065 = ~P3_LWORD_REG_8__SCAN_IN | ~n36103;
  assign P3_U2791 = ~n36066 | ~n36065;
  assign n36069 = ~n36067 & ~n36097;
  assign n36071 = ~n36069 & ~n36068;
  assign n36070 = ~P3_LWORD_REG_9__SCAN_IN | ~n36103;
  assign P3_U2792 = ~n36071 | ~n36070;
  assign n36074 = ~n36072 & ~n36097;
  assign n36076 = ~n36074 & ~n36073;
  assign n36075 = ~P3_LWORD_REG_10__SCAN_IN | ~n36103;
  assign P3_U2793 = ~n36076 | ~n36075;
  assign n36079 = ~n36077 & ~n36097;
  assign n36081 = ~n36079 & ~n36078;
  assign n36080 = ~P3_LWORD_REG_11__SCAN_IN | ~n36103;
  assign P3_U2794 = ~n36081 | ~n36080;
  assign n36084 = ~n36082 & ~n36097;
  assign n36086 = ~n36084 & ~n36083;
  assign n36085 = ~P3_LWORD_REG_12__SCAN_IN | ~n36103;
  assign P3_U2795 = ~n36086 | ~n36085;
  assign n36089 = ~n36087 & ~n36097;
  assign n36091 = ~n36089 & ~n36088;
  assign n36090 = ~P3_LWORD_REG_13__SCAN_IN | ~n36103;
  assign P3_U2796 = ~n36091 | ~n36090;
  assign n36094 = ~n36092 & ~n36097;
  assign n36096 = ~n36094 & ~n36093;
  assign n36095 = ~P3_LWORD_REG_14__SCAN_IN | ~n36103;
  assign P3_U2797 = ~n36096 | ~n36095;
  assign n36102 = ~n36098 & ~n36097;
  assign n36100 = ~BUF2_REG_15__SCAN_IN;
  assign n36101 = ~n36100 & ~n36099;
  assign n36105 = ~n36102 & ~n36101;
  assign n36104 = ~P3_LWORD_REG_15__SCAN_IN | ~n36103;
  assign P3_U2798 = ~n36105 | ~n36104;
  assign n36121 = ~n36508 & ~n36106;
  assign n36108 = ~n36484 & ~n36107;
  assign n36119 = ~n36109 | ~n36108;
  assign n36110 = ~n36484 & ~P3_PHYADDRPOINTER_REG_27__SCAN_IN;
  assign n36145 = ~n36113 | ~n36110;
  assign n36162 = ~P3_PHYADDRPOINTER_REG_26__SCAN_IN & ~n36262;
  assign n36116 = ~n36745 | ~n36111;
  assign n37401 = ~n39069 & ~n36112;
  assign n38823 = ~n37401;
  assign n36114 = ~n36113 & ~n38823;
  assign n36115 = ~n36114 & ~n36666;
  assign n36168 = ~n36116 | ~n36115;
  assign n36146 = ~n36162 & ~n36168;
  assign n36117 = ~n36145 | ~n36146;
  assign n36118 = ~n36117 | ~P3_PHYADDRPOINTER_REG_28__SCAN_IN;
  assign n36120 = ~n36119 | ~n36118;
  assign n36124 = ~n36121 & ~n36120;
  assign n36123 = ~n36122;
  assign n36127 = ~n36124 | ~n36123;
  assign n36125 = ~n36142 | ~P3_INSTADDRPOINTER_REG_27__SCAN_IN;
  assign n36126 = ~P3_INSTADDRPOINTER_REG_28__SCAN_IN & ~n36125;
  assign n36141 = ~n36127 & ~n36126;
  assign n36131 = ~n36490 & ~n36691;
  assign n36129 = ~n36613 & ~n36766;
  assign n36128 = ~n36731 & ~n36767;
  assign n36161 = ~n36129 & ~n36128;
  assign n36143 = ~P3_INSTADDRPOINTER_REG_27__SCAN_IN | ~n36161;
  assign n36130 = ~n36143 | ~P3_INSTADDRPOINTER_REG_28__SCAN_IN;
  assign n36139 = ~n36131 & ~n36130;
  assign n36133 = ~n36132;
  assign n36137 = ~n36134 & ~n36133;
  assign n36136 = ~n36135 | ~n36629;
  assign n36138 = ~n36137 & ~n36136;
  assign n36140 = ~n36139 & ~n36138;
  assign P3_U2802 = ~n36141 | ~n36140;
  assign n36144 = n36142 | P3_INSTADDRPOINTER_REG_27__SCAN_IN;
  assign n36160 = ~n36144 | ~n36143;
  assign n36757 = ~n22843 | ~P3_REIP_REG_27__SCAN_IN;
  assign n36158 = ~n36145 | ~n36757;
  assign n36150 = ~n36147 & ~n36146;
  assign n36149 = ~n36508 & ~n36148;
  assign n36156 = ~n36150 & ~n36149;
  assign n36153 = ~n36151;
  assign n36154 = ~n36153 | ~n36152;
  assign n36755 = ~n36154 ^ n36497;
  assign n36155 = ~n36629 | ~n36755;
  assign n36157 = ~n36156 | ~n36155;
  assign n36159 = ~n36158 & ~n36157;
  assign P3_U2803 = ~n36160 | ~n36159;
  assign n36177 = ~n36161 & ~n24282;
  assign n36163 = ~n36389 & ~n36162;
  assign n36171 = ~n23066 & ~n36163;
  assign n36802 = ~n22843 | ~P3_REIP_REG_26__SCAN_IN;
  assign n36165 = n38570 | n36164;
  assign n36167 = ~n36166 | ~n36165;
  assign n36169 = ~n36168 | ~n36167;
  assign n36170 = ~n36802 | ~n36169;
  assign n36175 = ~n36171 & ~n36170;
  assign n36173 = ~P3_INSTADDRPOINTER_REG_26__SCAN_IN & ~n36172;
  assign n36174 = ~P3_INSTADDRPOINTER_REG_25__SCAN_IN | ~n36173;
  assign n36176 = ~n36175 | ~n36174;
  assign n36179 = ~n36177 & ~n36176;
  assign n36178 = ~n36800 | ~n36629;
  assign P3_U2804 = ~n36179 | ~n36178;
  assign n36189 = ~n36508 & ~n36180;
  assign n36230 = ~n38115 | ~n36184;
  assign n36181 = ~n36745 | ~n36239;
  assign n36182 = ~n36230 | ~n36181;
  assign n36228 = ~n36666 & ~n36182;
  assign n36240 = ~n36390 | ~n36229;
  assign n36206 = ~n36228 | ~n36240;
  assign n36187 = ~P3_PHYADDRPOINTER_REG_25__SCAN_IN | ~n36206;
  assign n36185 = ~n36183 ^ P3_PHYADDRPOINTER_REG_24__SCAN_IN;
  assign n36204 = ~n36484 & ~n36184;
  assign n36186 = ~n36185 | ~n36204;
  assign n36188 = ~n36187 | ~n36186;
  assign n36190 = ~n36189 & ~n36188;
  assign n36830 = ~P3_REIP_REG_25__SCAN_IN | ~n22843;
  assign n36200 = ~n36190 | ~n36830;
  assign n36820 = ~P3_INSTADDRPOINTER_REG_25__SCAN_IN;
  assign n36192 = ~n36191;
  assign n36194 = ~n36192 | ~n36610;
  assign n36195 = ~n36194 | ~n36193;
  assign n36807 = n36820 ^ n36195;
  assign n36198 = ~n36807 | ~n36629;
  assign n36813 = n36820 ^ n36196;
  assign n36197 = ~n36813 | ~n36490;
  assign n36199 = ~n36198 | ~n36197;
  assign n36203 = ~n36200 & ~n36199;
  assign n36814 = n36820 ^ n36201;
  assign n36202 = ~n36691 | ~n36814;
  assign P3_U2805 = ~n36203 | ~n36202;
  assign n36250 = ~n36832 & ~n36613;
  assign n36248 = ~n36833 & ~n36731;
  assign n36238 = ~n36250 & ~n36248;
  assign n36219 = ~n36238 & ~n36849;
  assign n36208 = ~n36205 | ~n36204;
  assign n36207 = ~P3_PHYADDRPOINTER_REG_24__SCAN_IN | ~n36206;
  assign n36212 = ~n36208 | ~n36207;
  assign n36210 = ~n36389 | ~n36209;
  assign n36853 = ~n22843 | ~P3_REIP_REG_24__SCAN_IN;
  assign n36211 = ~n36210 | ~n36853;
  assign n36217 = ~n36212 & ~n36211;
  assign n36214 = ~n36213 | ~P3_INSTADDRPOINTER_REG_24__SCAN_IN;
  assign n36857 = ~n36215 | ~n36214;
  assign n36216 = ~n36857 | ~n36629;
  assign n36218 = ~n36217 | ~n36216;
  assign n36222 = ~n36219 & ~n36218;
  assign n36221 = ~n36220 | ~n36849;
  assign P3_U2806 = ~n36222 | ~n36221;
  assign n36761 = ~P3_INSTADDRPOINTER_REG_22__SCAN_IN;
  assign n36223 = ~n36278 & ~n36761;
  assign n36226 = ~n36223 & ~n36276;
  assign n36224 = ~n36497 | ~P3_INSTADDRPOINTER_REG_22__SCAN_IN;
  assign n36225 = ~n36333 | ~n36224;
  assign n36227 = ~n36226 & ~n36225;
  assign n36860 = n36869 ^ n36227;
  assign n36246 = ~n36580 & ~n36860;
  assign n38970 = ~P3_REIP_REG_23__SCAN_IN;
  assign n36861 = ~n37197 & ~n38970;
  assign n36233 = ~n36229 & ~n36228;
  assign n36232 = ~n36231 & ~n36230;
  assign n36236 = ~n36233 & ~n36232;
  assign n36235 = ~n36389 | ~n36234;
  assign n36237 = ~n36236 | ~n36235;
  assign n36244 = ~n36861 & ~n36237;
  assign n36242 = ~n36238 & ~n36869;
  assign n36241 = ~n36240 & ~n36239;
  assign n36243 = ~n36242 & ~n36241;
  assign n36245 = ~n36244 | ~n36243;
  assign n36255 = ~n36246 & ~n36245;
  assign n36252 = ~n36248 | ~n36247;
  assign n36251 = ~n36250 | ~n36249;
  assign n36253 = ~n36252 | ~n36251;
  assign n36254 = ~P3_INSTADDRPOINTER_REG_22__SCAN_IN | ~n36253;
  assign P3_U2807 = ~n36255 | ~n36254;
  assign n37009 = ~n36321;
  assign n36257 = ~n36691 | ~n37009;
  assign n36256 = ~n36490 | ~n37008;
  assign n36424 = ~n36257 | ~n36256;
  assign n36259 = ~n36258 | ~n36424;
  assign n36284 = ~P3_INSTADDRPOINTER_REG_22__SCAN_IN & ~n36259;
  assign n36261 = ~P3_PHYADDRPOINTER_REG_22__SCAN_IN & ~n36484;
  assign n36271 = ~n36261 | ~n36260;
  assign n36309 = ~P3_PHYADDRPOINTER_REG_20__SCAN_IN & ~n36262;
  assign n36264 = ~n36263 & ~n36478;
  assign n36266 = ~n36666 & ~n36264;
  assign n36265 = ~n37401 | ~n36267;
  assign n36314 = ~n36266 | ~n36265;
  assign n36289 = ~n36309 & ~n36314;
  assign n36268 = ~n36484 & ~n36267;
  assign n36295 = ~n36268 | ~n36290;
  assign n36269 = ~n36289 | ~n36295;
  assign n36270 = ~P3_PHYADDRPOINTER_REG_22__SCAN_IN | ~n36269;
  assign n36275 = ~n36271 | ~n36270;
  assign n36902 = ~P3_REIP_REG_22__SCAN_IN | ~n22843;
  assign n36273 = ~n36272 | ~n36389;
  assign n36274 = ~n36902 | ~n36273;
  assign n36282 = ~n36275 & ~n36274;
  assign n36277 = ~n36276;
  assign n36279 = ~n36278 | ~n36277;
  assign n36280 = ~n36279 | ~n36333;
  assign n36901 = ~n36280 ^ P3_INSTADDRPOINTER_REG_22__SCAN_IN;
  assign n36281 = ~n36629 | ~n36901;
  assign n36283 = ~n36282 | ~n36281;
  assign n36288 = ~n36284 & ~n36283;
  assign n36286 = ~n36691 | ~n36880;
  assign n36285 = ~n36490 | ~n36881;
  assign n36306 = ~n36286 | ~n36285;
  assign n36287 = ~P3_INSTADDRPOINTER_REG_22__SCAN_IN | ~n36306;
  assign P3_U2808 = ~n36288 | ~n36287;
  assign n36294 = ~n36290 & ~n36289;
  assign n36924 = ~n22843 | ~P3_REIP_REG_21__SCAN_IN;
  assign n36292 = ~n36389 | ~n36291;
  assign n36293 = ~n36924 | ~n36292;
  assign n36296 = ~n36294 & ~n36293;
  assign n36305 = ~n36296 | ~n36295;
  assign n36923 = ~P3_INSTADDRPOINTER_REG_21__SCAN_IN & ~n36951;
  assign n36341 = ~n36863 | ~n36424;
  assign n36319 = ~n36962 & ~n36341;
  assign n36303 = ~n36923 | ~n36319;
  assign n36373 = ~n36297;
  assign n36372 = ~n36610 ^ P3_INSTADDRPOINTER_REG_18__SCAN_IN;
  assign n36375 = ~n36373 | ~n36372;
  assign n36354 = ~n36375 & ~n36610;
  assign n36300 = ~n36298 | ~n36354;
  assign n36330 = ~n36375 | ~P3_INSTADDRPOINTER_REG_18__SCAN_IN;
  assign n36353 = ~n36497 & ~n36330;
  assign n36299 = ~n36909 | ~n36353;
  assign n36301 = ~n36300 | ~n36299;
  assign n36928 = n36301 ^ P3_INSTADDRPOINTER_REG_21__SCAN_IN;
  assign n36302 = ~n36629 | ~n36928;
  assign n36304 = ~n36303 | ~n36302;
  assign n36308 = ~n36305 & ~n36304;
  assign n36307 = ~P3_INSTADDRPOINTER_REG_21__SCAN_IN | ~n36306;
  assign P3_U2809 = ~n36308 | ~n36307;
  assign n36310 = ~n36389 & ~n36309;
  assign n36318 = ~n36311 & ~n36310;
  assign n36313 = ~n38115 | ~n36312;
  assign n36315 = ~n36313 | ~n23552;
  assign n36316 = ~n36315 | ~n36314;
  assign n36948 = ~n22843 | ~P3_REIP_REG_20__SCAN_IN;
  assign n36317 = ~n36316 | ~n36948;
  assign n36340 = ~n36318 & ~n36317;
  assign n36326 = ~n36951 | ~n36319;
  assign n36971 = ~n36320 & ~n36380;
  assign n36936 = ~n36322 | ~n36971;
  assign n36324 = ~n36490 | ~n36936;
  assign n36972 = ~n36380 & ~n36321;
  assign n36935 = ~n36322 | ~n36972;
  assign n36323 = ~n36691 | ~n36935;
  assign n36360 = ~n36324 | ~n36323;
  assign n36325 = ~P3_INSTADDRPOINTER_REG_20__SCAN_IN | ~n36360;
  assign n36338 = ~n36326 | ~n36325;
  assign n36329 = ~P3_INSTADDRPOINTER_REG_19__SCAN_IN & ~n36497;
  assign n36328 = ~n36610 & ~n36327;
  assign n36332 = ~n36329 & ~n36328;
  assign n36331 = ~P3_INSTADDRPOINTER_REG_19__SCAN_IN | ~n36330;
  assign n36335 = ~n36332 | ~n36331;
  assign n36334 = ~n36333;
  assign n36336 = ~n36335 & ~n36334;
  assign n36931 = ~n36336 ^ P3_INSTADDRPOINTER_REG_20__SCAN_IN;
  assign n36337 = ~n36580 & ~n36931;
  assign n36339 = ~n36338 & ~n36337;
  assign P3_U2810 = ~n36340 | ~n36339;
  assign n36359 = ~P3_INSTADDRPOINTER_REG_19__SCAN_IN & ~n36341;
  assign n36958 = ~P3_REIP_REG_19__SCAN_IN | ~n22843;
  assign n36343 = ~n36342 | ~n36389;
  assign n36352 = ~n36958 | ~n36343;
  assign n36344 = n36347 & n37401;
  assign n36387 = ~n36666 & ~n36344;
  assign n36346 = ~n36745 | ~n36345;
  assign n36369 = ~n36387 | ~n36346;
  assign n36350 = ~P3_PHYADDRPOINTER_REG_19__SCAN_IN | ~n36369;
  assign n36348 = ~P3_PHYADDRPOINTER_REG_19__SCAN_IN ^ n36364;
  assign n36365 = ~n36484 & ~n36347;
  assign n36349 = ~n36348 | ~n36365;
  assign n36351 = ~n36350 | ~n36349;
  assign n36357 = ~n36352 & ~n36351;
  assign n36355 = ~n36354 & ~n36353;
  assign n36956 = n36355 ^ n36962;
  assign n36356 = ~n36629 | ~n36956;
  assign n36358 = ~n36357 | ~n36356;
  assign n36362 = ~n36359 & ~n36358;
  assign n36361 = ~P3_INSTADDRPOINTER_REG_19__SCAN_IN | ~n36360;
  assign P3_U2811 = ~n36362 | ~n36361;
  assign n36368 = ~n36508 & ~n36363;
  assign n36967 = ~P3_REIP_REG_18__SCAN_IN | ~n22843;
  assign n36366 = ~n36365 | ~n36364;
  assign n36367 = ~n36967 | ~n36366;
  assign n36371 = ~n36368 & ~n36367;
  assign n36370 = ~P3_PHYADDRPOINTER_REG_18__SCAN_IN | ~n36369;
  assign n36379 = ~n36371 | ~n36370;
  assign n36374 = n36373 | n36372;
  assign n36965 = ~n36375 | ~n36374;
  assign n36377 = ~n36965 | ~n36629;
  assign n36994 = ~P3_INSTADDRPOINTER_REG_18__SCAN_IN & ~n36380;
  assign n36376 = ~n36994 | ~n36424;
  assign n36378 = ~n36377 | ~n36376;
  assign n36383 = ~n36379 & ~n36378;
  assign n36428 = ~n37009 & ~n36731;
  assign n36429 = ~n37008 & ~n36613;
  assign n36403 = ~n36428 & ~n36429;
  assign n36381 = ~n36380 | ~n36424;
  assign n36394 = ~n36403 | ~n36381;
  assign n36382 = ~P3_INSTADDRPOINTER_REG_18__SCAN_IN | ~n36394;
  assign P3_U2812 = ~n36383 | ~n36382;
  assign n37001 = ~n37197 & ~n38940;
  assign n36385 = n38115 & n36384;
  assign n36386 = ~P3_PHYADDRPOINTER_REG_17__SCAN_IN & ~n36385;
  assign n36388 = ~n36387 & ~n36386;
  assign n36393 = ~n37001 & ~n36388;
  assign n36392 = ~n36391 | ~n36702;
  assign n36398 = ~n36393 | ~n36392;
  assign n36396 = ~P3_INSTADDRPOINTER_REG_17__SCAN_IN | ~n36394;
  assign n37024 = ~P3_INSTADDRPOINTER_REG_16__SCAN_IN;
  assign n37003 = ~P3_INSTADDRPOINTER_REG_17__SCAN_IN & ~n37024;
  assign n36395 = ~n37003 | ~n36424;
  assign n36397 = ~n36396 | ~n36395;
  assign n36402 = ~n36398 & ~n36397;
  assign n37002 = ~n36400 ^ P3_INSTADDRPOINTER_REG_17__SCAN_IN;
  assign n36401 = ~n37002 | ~n36629;
  assign P3_U2813 = ~n36402 | ~n36401;
  assign n36423 = ~n36403 & ~n37024;
  assign n36417 = ~n36508 & ~n36404;
  assign n36407 = ~P3_PHYADDRPOINTER_REG_15__SCAN_IN & ~P3_PHYADDRPOINTER_REG_16__SCAN_IN;
  assign n36448 = ~n36484 & ~n36408;
  assign n36406 = ~n36405 | ~n36448;
  assign n36414 = ~n36407 & ~n36406;
  assign n36409 = ~n37401 | ~n36408;
  assign n36457 = ~n36743 | ~n36409;
  assign n36411 = ~n36410 & ~n36478;
  assign n36445 = ~n36457 & ~n36411;
  assign n36413 = ~n36445 & ~n36412;
  assign n36415 = ~n36414 & ~n36413;
  assign n37030 = ~P3_REIP_REG_16__SCAN_IN | ~n22843;
  assign n36416 = ~n36415 | ~n37030;
  assign n36421 = ~n36417 & ~n36416;
  assign n36418 = ~n36497 ^ P3_INSTADDRPOINTER_REG_16__SCAN_IN;
  assign n37023 = ~n36419 ^ n36418;
  assign n36420 = ~n37023 | ~n36629;
  assign n36422 = ~n36421 | ~n36420;
  assign n36426 = ~n36423 & ~n36422;
  assign n36425 = ~n36424 | ~n37024;
  assign P3_U2814 = ~n36426 | ~n36425;
  assign n37047 = ~P3_INSTADDRPOINTER_REG_15__SCAN_IN;
  assign n36427 = ~P3_INSTADDRPOINTER_REG_14__SCAN_IN | ~n36462;
  assign n37034 = ~n37047 | ~n36427;
  assign n36431 = ~n36428 | ~n37034;
  assign n36465 = ~n37183 | ~n36990;
  assign n37032 = ~n37047 | ~n36465;
  assign n36430 = ~n36429 | ~n37032;
  assign n36443 = ~n36431 | ~n36430;
  assign n36433 = ~n36432;
  assign n36434 = ~n36433 & ~P3_INSTADDRPOINTER_REG_13__SCAN_IN;
  assign n36435 = ~n36434 | ~n36574;
  assign n36436 = ~n36554 & ~n36435;
  assign n36471 = ~n36436 | ~n36498;
  assign n36440 = ~n36471 | ~n37080;
  assign n36438 = n36610 & n36437;
  assign n36472 = ~n36515 | ~n36438;
  assign n36439 = ~n36472 | ~P3_INSTADDRPOINTER_REG_14__SCAN_IN;
  assign n36441 = ~n36440 | ~n36439;
  assign n37046 = n36441 ^ P3_INSTADDRPOINTER_REG_15__SCAN_IN;
  assign n36442 = ~n37046 & ~n36580;
  assign n36454 = ~n36443 & ~n36442;
  assign n36452 = ~n36508 & ~n36444;
  assign n36446 = ~n36445 & ~n36447;
  assign n37044 = ~n37197 & ~n38930;
  assign n36450 = ~n36446 & ~n37044;
  assign n36449 = ~n36448 | ~n36447;
  assign n36451 = ~n36450 | ~n36449;
  assign n36453 = ~n36452 & ~n36451;
  assign P3_U2815 = ~n36454 | ~n36453;
  assign n36456 = ~n38115 | ~n23075;
  assign n36458 = ~n36456 | ~n36455;
  assign n36461 = ~n36458 | ~n36457;
  assign n36460 = ~n36459 | ~n36702;
  assign n36470 = ~n36461 | ~n36460;
  assign n37053 = n37080 ^ n36462;
  assign n36467 = ~n36731 & ~n37053;
  assign n36464 = ~n36463 | ~n37080;
  assign n37052 = ~n36465 | ~n36464;
  assign n36466 = ~n36613 & ~n37052;
  assign n36468 = ~n36467 & ~n36466;
  assign n37079 = ~n22843 | ~P3_REIP_REG_14__SCAN_IN;
  assign n36469 = ~n36468 | ~n37079;
  assign n36475 = ~n36470 & ~n36469;
  assign n36473 = ~n36472 | ~n36471;
  assign n37077 = n36473 ^ P3_INSTADDRPOINTER_REG_14__SCAN_IN;
  assign n36474 = ~n36629 | ~n37077;
  assign P3_U2816 = ~n36475 | ~n36474;
  assign n36526 = ~n37091 & ~n36613;
  assign n37142 = ~n37087 | ~n37185;
  assign n37093 = ~n37085 & ~n37142;
  assign n36524 = ~n37093 & ~n36731;
  assign n36523 = ~n36526 & ~n36524;
  assign n36496 = ~n36523 & ~n37066;
  assign n36489 = ~n36508 & ~n36476;
  assign n36481 = ~n36478 & ~n36477;
  assign n36479 = ~n37401 | ~n36540;
  assign n36480 = ~n36743 | ~n36479;
  assign n36509 = ~n36481 & ~n36480;
  assign n36482 = ~n36483 & ~n36509;
  assign n37112 = ~n37197 & ~n38920;
  assign n36487 = ~n36482 & ~n37112;
  assign n36485 = ~n36483 ^ P3_PHYADDRPOINTER_REG_12__SCAN_IN;
  assign n36510 = ~n36484 & ~n36540;
  assign n36486 = ~n36485 | ~n36510;
  assign n36488 = ~n36487 | ~n36486;
  assign n36494 = ~n36489 & ~n36488;
  assign n37106 = ~P3_INSTADDRPOINTER_REG_13__SCAN_IN & ~n37059;
  assign n36492 = ~n37183 | ~n36490;
  assign n36491 = ~n36691 | ~n37185;
  assign n36600 = ~n36492 | ~n36491;
  assign n36493 = ~n37106 | ~n36600;
  assign n36495 = ~n36494 | ~n36493;
  assign n36506 = ~n36496 & ~n36495;
  assign n36503 = ~P3_INSTADDRPOINTER_REG_12__SCAN_IN & ~n36497;
  assign n36571 = ~n36498;
  assign n36499 = ~n36574 | ~n37154;
  assign n36500 = ~n36571 & ~n36499;
  assign n36516 = ~n36500 & ~n36610;
  assign n37123 = ~P3_INSTADDRPOINTER_REG_12__SCAN_IN;
  assign n36501 = ~n36515 & ~n37123;
  assign n36502 = n36516 | n36501;
  assign n36504 = ~n36503 & ~n36502;
  assign n37107 = ~n37066 ^ n36504;
  assign n36505 = ~n37107 | ~n36629;
  assign P3_U2817 = ~n36506 | ~n36505;
  assign n36522 = ~n36508 & ~n36507;
  assign n36514 = ~n36509 & ~n36511;
  assign n37130 = ~n22843 | ~P3_REIP_REG_12__SCAN_IN;
  assign n36512 = ~n36511 | ~n36510;
  assign n36513 = ~n37130 | ~n36512;
  assign n36520 = ~n36514 & ~n36513;
  assign n36518 = ~n36516 & ~n36515;
  assign n36517 = ~n36610 ^ P3_INSTADDRPOINTER_REG_12__SCAN_IN;
  assign n37128 = ~n36518 ^ n36517;
  assign n36519 = ~n36629 | ~n37128;
  assign n36521 = ~n36520 | ~n36519;
  assign n36534 = ~n36522 & ~n36521;
  assign n36532 = ~n36523 & ~n37123;
  assign n36525 = ~n36524;
  assign n36529 = ~n37142 & ~n36525;
  assign n36527 = ~n36526;
  assign n36528 = ~n37146 & ~n36527;
  assign n36530 = ~n36529 & ~n36528;
  assign n36531 = ~n37154 & ~n36530;
  assign n36533 = ~n36532 & ~n36531;
  assign P3_U2818 = ~n36534 | ~n36533;
  assign n36545 = ~n36535 | ~n36702;
  assign n37138 = ~n37197 & ~n38910;
  assign n36614 = ~n38115 | ~n36536;
  assign n36584 = ~n36537 & ~n36614;
  assign n36736 = ~n38823 | ~n36743;
  assign n36591 = ~n36736;
  assign n36539 = ~n36591 & ~n36538;
  assign n36542 = ~n36584 & ~n36539;
  assign n36541 = ~n36540 & ~n38570;
  assign n36543 = ~n36542 & ~n36541;
  assign n36544 = ~n37138 & ~n36543;
  assign n36553 = ~n36545 | ~n36544;
  assign n36546 = ~P3_INSTADDRPOINTER_REG_11__SCAN_IN & ~n37121;
  assign n36551 = ~n36546 | ~n36600;
  assign n36548 = ~n36613 & ~n37183;
  assign n36547 = ~n36731 & ~n37185;
  assign n36589 = ~n36548 & ~n36547;
  assign n36549 = ~n37121 | ~n36600;
  assign n36563 = ~n36589 | ~n36549;
  assign n36550 = ~P3_INSTADDRPOINTER_REG_11__SCAN_IN | ~n36563;
  assign n36552 = ~n36551 | ~n36550;
  assign n36561 = ~n36553 & ~n36552;
  assign n36605 = ~n36554 & ~P3_INSTADDRPOINTER_REG_8__SCAN_IN;
  assign n36558 = ~n36605 | ~n36574;
  assign n36555 = ~n36610 | ~P3_INSTADDRPOINTER_REG_8__SCAN_IN;
  assign n36606 = ~n36556 & ~n36555;
  assign n36557 = ~n36606 | ~n37087;
  assign n36559 = ~n36558 | ~n36557;
  assign n37135 = P3_INSTADDRPOINTER_REG_11__SCAN_IN ^ n36559;
  assign n36560 = ~n36629 | ~n37135;
  assign P3_U2819 = ~n36561 | ~n36560;
  assign n37177 = ~n37197 & ~n38905;
  assign n36562 = ~n36600 | ~P3_INSTADDRPOINTER_REG_9__SCAN_IN;
  assign n37151 = ~P3_INSTADDRPOINTER_REG_10__SCAN_IN;
  assign n36564 = ~n36562 | ~n37151;
  assign n36567 = ~n36564 | ~n36563;
  assign n36566 = ~n36565 | ~n36702;
  assign n36568 = ~n36567 | ~n36566;
  assign n36588 = ~n37177 & ~n36568;
  assign n36569 = ~P3_INSTADDRPOINTER_REG_9__SCAN_IN & ~n36610;
  assign n36570 = ~n36606 & ~n36569;
  assign n36573 = ~n37151 & ~n36570;
  assign n37206 = ~P3_INSTADDRPOINTER_REG_9__SCAN_IN;
  assign n36572 = ~n36571 | ~n37206;
  assign n36579 = ~n36573 | ~n36572;
  assign n37162 = ~P3_INSTADDRPOINTER_REG_9__SCAN_IN | ~n37151;
  assign n36577 = ~n37162 & ~n36606;
  assign n36575 = ~n36574;
  assign n36576 = ~n36575 & ~n36605;
  assign n36578 = ~n36577 & ~n36576;
  assign n37164 = ~n36579 | ~n36578;
  assign n36586 = ~n37164 & ~n36580;
  assign n36593 = ~n36622 & ~n36614;
  assign n36595 = P3_PHYADDRPOINTER_REG_9__SCAN_IN & n36593;
  assign n36582 = ~n36591 & ~n36581;
  assign n36583 = ~n36595 & ~n36582;
  assign n36585 = ~n36584 & ~n36583;
  assign n36587 = ~n36586 & ~n36585;
  assign P3_U2820 = ~n36588 | ~n36587;
  assign n36604 = ~n36589 & ~n37206;
  assign n36592 = ~n36591 & ~n36590;
  assign n36594 = ~n36593 & ~n36592;
  assign n36599 = ~n36595 & ~n36594;
  assign n37203 = ~n22843 | ~P3_REIP_REG_9__SCAN_IN;
  assign n36597 = ~n36596 | ~n36702;
  assign n36598 = ~n37203 | ~n36597;
  assign n36602 = ~n36599 & ~n36598;
  assign n36601 = ~n36600 | ~n37206;
  assign n36603 = ~n36602 | ~n36601;
  assign n36609 = ~n36604 & ~n36603;
  assign n36607 = ~n36606 & ~n36605;
  assign n37200 = n36607 ^ n37206;
  assign n36608 = ~n36629 | ~n37200;
  assign P3_U2821 = ~n36609 | ~n36608;
  assign n36611 = ~n36610 ^ n37210;
  assign n37213 = ~n36612 ^ n36611;
  assign n36628 = ~n37213 & ~n36613;
  assign n36618 = ~n36614 & ~P3_PHYADDRPOINTER_REG_8__SCAN_IN;
  assign n37233 = ~n22843 | ~P3_REIP_REG_8__SCAN_IN;
  assign n36616 = ~n36615 | ~n36702;
  assign n36617 = ~n37233 | ~n36616;
  assign n36626 = ~n36618 & ~n36617;
  assign n37227 = n37210 ^ n36619;
  assign n36624 = ~n37227 & ~n36731;
  assign n36640 = ~P3_PHYADDRPOINTER_REG_7__SCAN_IN & ~n38570;
  assign n36620 = ~n37401 | ~n36639;
  assign n36634 = ~n36743 | ~n36620;
  assign n36621 = ~n36640 & ~n36634;
  assign n36623 = ~n36622 & ~n36621;
  assign n36625 = ~n36624 & ~n36623;
  assign n36627 = ~n36626 | ~n36625;
  assign n36631 = ~n36628 & ~n36627;
  assign n36630 = ~n37213 | ~n36629;
  assign P3_U2822 = ~n36631 | ~n36630;
  assign n37242 = ~n36632 ^ n37235;
  assign n36733 = ~n36727;
  assign n36644 = ~n37242 & ~n36733;
  assign n36638 = ~n36730 & ~n36633;
  assign n37237 = ~n37197 & ~n38890;
  assign n36636 = ~n37237;
  assign n36635 = ~P3_PHYADDRPOINTER_REG_7__SCAN_IN | ~n36634;
  assign n36637 = ~n36636 | ~n36635;
  assign n36642 = ~n36638 & ~n36637;
  assign n36641 = ~n36640 | ~n23795;
  assign n36643 = ~n36642 | ~n36641;
  assign n36648 = ~n36644 & ~n36643;
  assign n36646 = ~n36645 & ~n23059;
  assign n37238 = n36646 ^ P3_INSTADDRPOINTER_REG_7__SCAN_IN;
  assign n36647 = ~n37238 | ~n36691;
  assign P3_U2823 = ~n36648 | ~n36647;
  assign n37272 = ~n22843 | ~P3_REIP_REG_6__SCAN_IN;
  assign n36650 = ~n36649 | ~n36702;
  assign n36661 = ~n37272 | ~n36650;
  assign n37250 = n36652 ^ n36651;
  assign n36659 = ~n36727 | ~n37250;
  assign n36655 = ~n38115 | ~n36653;
  assign n36669 = ~n36736 | ~n36655;
  assign n36657 = ~n36669 & ~n36654;
  assign n36656 = ~P3_PHYADDRPOINTER_REG_6__SCAN_IN & ~n36655;
  assign n36658 = ~n36657 & ~n36656;
  assign n36660 = ~n36659 | ~n36658;
  assign n36664 = ~n36661 & ~n36660;
  assign n37251 = ~n37257 ^ n36662;
  assign n36663 = ~n36691 | ~n37251;
  assign P3_U2824 = ~n36664 | ~n36663;
  assign n36667 = ~n36666 & ~n36665;
  assign n36668 = ~P3_PHYADDRPOINTER_REG_5__SCAN_IN & ~n36667;
  assign n36676 = ~n36669 & ~n36668;
  assign n36671 = n36670 & n36702;
  assign n37287 = ~n37197 & ~n38880;
  assign n36674 = ~n36671 & ~n37287;
  assign n37274 = ~n36672 ^ P3_INSTADDRPOINTER_REG_5__SCAN_IN;
  assign n36673 = ~n36727 | ~n37274;
  assign n36675 = ~n36674 | ~n36673;
  assign n36680 = ~n36676 & ~n36675;
  assign n37275 = n36678 ^ n36677;
  assign n36679 = ~n36691 | ~n37275;
  assign P3_U2825 = ~n36680 | ~n36679;
  assign n37291 = ~n37197 & ~n38875;
  assign n37306 = ~n36683 ^ n36682;
  assign n36684 = ~n36733 & ~n37306;
  assign n36698 = ~n37291 & ~n36684;
  assign n36685 = ~P3_PHYADDRPOINTER_REG_4__SCAN_IN & ~n36686;
  assign n36689 = ~n36685 | ~n38115;
  assign n36687 = ~n37401 | ~n36686;
  assign n36700 = ~n36743 | ~n36687;
  assign n36688 = ~P3_PHYADDRPOINTER_REG_4__SCAN_IN | ~n36700;
  assign n36696 = ~n36689 | ~n36688;
  assign n36694 = ~n36691 | ~n37293;
  assign n36693 = ~n36692 | ~n36702;
  assign n36695 = ~n36694 | ~n36693;
  assign n36697 = ~n36696 & ~n36695;
  assign P3_U2826 = ~n36698 | ~n36697;
  assign n36718 = ~P3_PHYADDRPOINTER_REG_2__SCAN_IN | ~n36743;
  assign n36701 = ~n36718 | ~n36699;
  assign n36714 = ~n36701 | ~n36700;
  assign n37315 = ~n37197 & ~n38870;
  assign n36711 = ~n36703 | ~n36702;
  assign n37321 = ~n36705 ^ n36704;
  assign n36709 = ~n36731 & ~n37321;
  assign n37320 = ~n36707 ^ n36706;
  assign n36708 = ~n36733 & ~n37320;
  assign n36710 = ~n36709 & ~n36708;
  assign n36712 = ~n36711 | ~n36710;
  assign n36713 = ~n37315 & ~n36712;
  assign P3_U2827 = ~n36714 | ~n36713;
  assign n37329 = ~n36716 ^ n36715;
  assign n36725 = ~n36731 & ~n37329;
  assign n36719 = ~n36717 | ~n38570;
  assign n36723 = ~n36719 | ~n36718;
  assign n36721 = ~n36720 & ~n36730;
  assign n37350 = ~n37197 & ~n38865;
  assign n36722 = ~n36721 & ~n37350;
  assign n36724 = ~n36723 | ~n36722;
  assign n36729 = ~n36725 & ~n36724;
  assign n36728 = ~n36727 | ~n37331;
  assign P3_U2828 = ~n36729 | ~n36728;
  assign n36740 = ~n36730 & ~P3_PHYADDRPOINTER_REG_1__SCAN_IN;
  assign n37361 = ~n36732 ^ n36750;
  assign n36735 = ~n36731 & ~n37361;
  assign n37362 = ~n36732 ^ n36749;
  assign n36734 = ~n36733 & ~n37362;
  assign n36738 = ~n36735 & ~n36734;
  assign n36737 = ~P3_PHYADDRPOINTER_REG_1__SCAN_IN | ~n36736;
  assign n36739 = ~n36738 | ~n36737;
  assign n36742 = ~n36740 & ~n36739;
  assign n37371 = ~n37197 & ~n39084;
  assign n36741 = ~n37371;
  assign P3_U2829 = ~n36742 | ~n36741;
  assign n36744 = ~n39069 | ~n36743;
  assign n36746 = ~n36745 & ~n36744;
  assign n36748 = ~n36747 & ~n36746;
  assign n37385 = ~n39083 & ~n37197;
  assign n36754 = ~n36748 & ~n37385;
  assign n37374 = ~n36750 & ~n36749;
  assign n36752 = n37374 ^ n37453;
  assign n36753 = ~n36752 | ~n36751;
  assign P3_U2830 = ~n36754 | ~n36753;
  assign n36756 = ~n37201 | ~n36755;
  assign n36759 = ~n36757 | ~n36756;
  assign n36758 = ~n36764 & ~n37383;
  assign n36790 = ~n36759 & ~n36758;
  assign n36810 = ~n38673 & ~n36842;
  assign n36877 = ~n36760;
  assign n36762 = ~n36877 & ~n36761;
  assign n36850 = ~n36810 & ~n36762;
  assign n36763 = ~P3_INSTADDRPOINTER_REG_25__SCAN_IN | ~n36811;
  assign n36797 = ~n36850 & ~n36763;
  assign n36765 = ~n36797 | ~P3_INSTADDRPOINTER_REG_26__SCAN_IN;
  assign n36788 = ~n36765 | ~n36764;
  assign n36769 = ~n37184 & ~n36766;
  assign n36768 = ~n38674 & ~n36767;
  assign n36779 = ~n36769 & ~n36768;
  assign n36777 = ~P3_INSTADDRPOINTER_REG_25__SCAN_IN & ~n22828;
  assign n36773 = ~n22834 & ~n36770;
  assign n36771 = ~n36864;
  assign n36772 = ~n36916 & ~n36771;
  assign n36840 = ~n22828 & ~n36772;
  assign n36776 = ~n36773 & ~n36840;
  assign n36775 = ~n36774 | ~n38758;
  assign n36817 = ~n36776 | ~n36775;
  assign n36778 = ~n36777 & ~n36817;
  assign n36791 = ~n36779 | ~n36778;
  assign n36783 = ~n36780 & ~n36791;
  assign n36782 = ~n38757 | ~n36781;
  assign n36785 = ~n36783 | ~n36782;
  assign n36784 = ~n22828 & ~P3_INSTADDRPOINTER_REG_26__SCAN_IN;
  assign n36786 = ~n36785 & ~n36784;
  assign n36787 = ~n37349 & ~n36786;
  assign n36789 = ~n36788 | ~n36787;
  assign P3_U2835 = ~n36790 | ~n36789;
  assign n36795 = ~n24282 & ~n36791;
  assign n36818 = ~n36792 & ~n38673;
  assign n36793 = ~P3_INSTADDRPOINTER_REG_25__SCAN_IN & ~n36932;
  assign n36794 = ~n36818 & ~n36793;
  assign n36796 = ~n36795 | ~n36794;
  assign n36799 = ~n36796 | ~n24731;
  assign n36798 = ~P3_INSTADDRPOINTER_REG_26__SCAN_IN & ~n36797;
  assign n36804 = ~n36799 & ~n36798;
  assign n36801 = ~n36800 | ~n37201;
  assign n36803 = ~n36802 | ~n36801;
  assign n36806 = ~n36804 & ~n36803;
  assign n36805 = ~n37352 | ~P3_INSTADDRPOINTER_REG_26__SCAN_IN;
  assign P3_U2836 = ~n36806 | ~n36805;
  assign n36829 = ~n36820 & ~n37383;
  assign n36827 = ~n37201 | ~n36807;
  assign n36809 = n36808 & P3_INSTADDRPOINTER_REG_22__SCAN_IN;
  assign n36865 = ~n36810 & ~n36809;
  assign n36812 = ~P3_INSTADDRPOINTER_REG_25__SCAN_IN & ~n36865;
  assign n36824 = ~n36812 | ~n36811;
  assign n36816 = ~n36813 | ~n37147;
  assign n36815 = ~n36814 | ~n37292;
  assign n36822 = ~n36816 | ~n36815;
  assign n36819 = ~n36818 & ~n36817;
  assign n36821 = ~n36820 & ~n36819;
  assign n36823 = ~n36822 & ~n36821;
  assign n36825 = ~n36824 | ~n36823;
  assign n36826 = ~n24731 | ~n36825;
  assign n36828 = ~n36827 | ~n36826;
  assign n36831 = ~n36829 & ~n36828;
  assign P3_U2837 = ~n36831 | ~n36830;
  assign n36835 = ~n37184 & ~n36832;
  assign n36834 = ~n38674 & ~n36833;
  assign n36838 = ~n36835 & ~n36834;
  assign n36837 = ~n38757 | ~n36836;
  assign n36839 = ~n36838 | ~n36837;
  assign n36841 = ~n36840 & ~n36839;
  assign n36845 = ~n36841 | ~n37383;
  assign n36848 = ~n36845 & ~n37356;
  assign n36843 = ~n38730 | ~n36842;
  assign n36844 = ~P3_INSTADDRPOINTER_REG_23__SCAN_IN | ~n36843;
  assign n36846 = ~n36845 & ~n36844;
  assign n36871 = ~n22843 & ~n36846;
  assign n36847 = ~P3_INSTADDRPOINTER_REG_24__SCAN_IN | ~n36871;
  assign n36856 = ~n36848 & ~n36847;
  assign n36851 = ~n36849 | ~n24731;
  assign n36852 = ~n36851 & ~n36850;
  assign n36854 = ~n36852 | ~P3_INSTADDRPOINTER_REG_23__SCAN_IN;
  assign n36855 = ~n36854 | ~n36853;
  assign n36859 = ~n36856 & ~n36855;
  assign n36858 = ~n36857 | ~n37201;
  assign P3_U2838 = ~n36859 | ~n36858;
  assign n36862 = ~n37165 & ~n36860;
  assign n36873 = ~n36862 & ~n36861;
  assign n36908 = ~n36863;
  assign n36917 = ~n36987 & ~n36908;
  assign n36866 = ~n36864 | ~n36917;
  assign n36867 = ~n36866 | ~n36865;
  assign n36868 = ~n36867 | ~n37383;
  assign n36870 = ~n36869 | ~n36868;
  assign n36872 = ~n36871 | ~n36870;
  assign P3_U2839 = ~n36873 | ~n36872;
  assign n36875 = ~n36874 & ~n36975;
  assign n36876 = ~n36875 | ~n38730;
  assign n36878 = ~n36877 | ~n36876;
  assign n36900 = ~P3_INSTADDRPOINTER_REG_22__SCAN_IN & ~n36878;
  assign n36896 = ~n22834 & ~n36879;
  assign n36883 = ~n37292 | ~n36880;
  assign n36882 = ~n37147 | ~n36881;
  assign n36891 = ~n36883 | ~n36882;
  assign n36886 = ~n22828 & ~n36884;
  assign n36885 = ~n38673 & ~n36919;
  assign n36943 = ~n36886 & ~n36885;
  assign n36888 = ~P3_INSTADDRPOINTER_REG_20__SCAN_IN & ~n22828;
  assign n36887 = ~n38673 & ~n36909;
  assign n36889 = ~n36888 & ~n36887;
  assign n36890 = ~n36943 | ~n36889;
  assign n36911 = ~n36891 & ~n36890;
  assign n36894 = ~n36893 | ~n36892;
  assign n36895 = ~n36911 | ~n36894;
  assign n36897 = ~n36896 & ~n36895;
  assign n36898 = ~n36897 | ~P3_INSTADDRPOINTER_REG_22__SCAN_IN;
  assign n36899 = ~n24731 | ~n36898;
  assign n36905 = ~n36900 & ~n36899;
  assign n36903 = ~n36901 | ~n37201;
  assign n36904 = ~n36903 | ~n36902;
  assign n36907 = ~n36905 & ~n36904;
  assign n36906 = ~n37352 | ~P3_INSTADDRPOINTER_REG_22__SCAN_IN;
  assign P3_U2840 = ~n36907 | ~n36906;
  assign n36934 = ~n36908 & ~n37010;
  assign n36910 = ~n36934 | ~n36909;
  assign n36912 = ~n36910 | ~n38757;
  assign n36913 = ~n36912 | ~n36911;
  assign n36915 = ~n36913 & ~n37349;
  assign n36914 = ~n37197 | ~P3_INSTADDRPOINTER_REG_21__SCAN_IN;
  assign n36927 = ~n36915 & ~n36914;
  assign n37355 = ~n22828 | ~n37382;
  assign n36980 = ~n37338;
  assign n37334 = ~n37355 | ~n36980;
  assign n36918 = ~n36916 & ~n37334;
  assign n36921 = ~n36918 & ~n36917;
  assign n36920 = ~n36919 | ~n38730;
  assign n36922 = ~n36921 | ~n36920;
  assign n36955 = ~n24731 | ~n36922;
  assign n36952 = ~n36962 & ~n36955;
  assign n36925 = ~n36952 | ~n36923;
  assign n36926 = ~n36925 | ~n36924;
  assign n36930 = ~n36927 & ~n36926;
  assign n36929 = ~n37201 | ~n36928;
  assign P3_U2841 = ~n36930 | ~n36929;
  assign n36950 = ~n37165 & ~n36931;
  assign n37358 = ~n36932;
  assign n36933 = ~P3_INSTADDRPOINTER_REG_19__SCAN_IN & ~n38803;
  assign n36945 = ~n37358 | ~n36933;
  assign n36941 = ~n22834 & ~n36934;
  assign n36938 = ~n36935 | ~n37292;
  assign n36937 = ~n37147 | ~n36936;
  assign n36939 = n36938 & n36937;
  assign n36940 = ~n37383 | ~n36939;
  assign n36942 = ~n36941 & ~n36940;
  assign n36944 = ~n36943 | ~n36942;
  assign n36961 = ~n37197 | ~n36944;
  assign n36946 = ~n36945 | ~n36961;
  assign n36947 = ~P3_INSTADDRPOINTER_REG_20__SCAN_IN | ~n36946;
  assign n36949 = ~n36948 | ~n36947;
  assign n36954 = ~n36950 & ~n36949;
  assign n36953 = ~n36952 | ~n36951;
  assign P3_U2842 = ~n36954 | ~n36953;
  assign n36960 = ~P3_INSTADDRPOINTER_REG_19__SCAN_IN & ~n36955;
  assign n36957 = ~n37201 | ~n36956;
  assign n36959 = ~n36958 | ~n36957;
  assign n36964 = ~n36960 & ~n36959;
  assign n36963 = n36962 | n36961;
  assign P3_U2843 = ~n36964 | ~n36963;
  assign n36966 = ~n36965 | ~n37201;
  assign n36986 = ~n36967 | ~n36966;
  assign n37263 = ~n37382 | ~n38757;
  assign n37336 = ~n37263;
  assign n36969 = ~n36968 | ~P3_INSTADDRPOINTER_REG_16__SCAN_IN;
  assign n36970 = ~n37336 & ~n36969;
  assign n36979 = ~n37338 & ~n36970;
  assign n36974 = ~n37184 & ~n36971;
  assign n36973 = ~n38674 & ~n36972;
  assign n36977 = ~n36974 & ~n36973;
  assign n36976 = ~n38730 | ~n36975;
  assign n36978 = ~n36977 | ~n36976;
  assign n36997 = ~n36979 & ~n36978;
  assign n36981 = ~n24269 | ~n36980;
  assign n36982 = ~n36997 | ~n36981;
  assign n36984 = ~n37352 & ~n36982;
  assign n36983 = ~P3_INSTADDRPOINTER_REG_18__SCAN_IN | ~n37197;
  assign n36985 = ~n36984 & ~n36983;
  assign n36996 = ~n36986 & ~n36985;
  assign n36992 = ~n36987;
  assign n36989 = ~n38673 & ~n37218;
  assign n36988 = ~n37188 & ~n37334;
  assign n37211 = ~P3_INSTADDRPOINTER_REG_7__SCAN_IN | ~n37239;
  assign n37105 = ~n37210 & ~n37211;
  assign n37038 = ~n36990 | ~n37105;
  assign n36991 = ~n37047 & ~n37038;
  assign n36993 = ~n36992 & ~n36991;
  assign n37025 = ~n36993 & ~n37349;
  assign n36995 = ~n36994 | ~n37025;
  assign P3_U2844 = ~n36996 | ~n36995;
  assign n36998 = ~n36997 & ~n37349;
  assign n36999 = ~n37352 & ~n36998;
  assign n37000 = ~n24269 & ~n36999;
  assign n37007 = ~n37001 & ~n37000;
  assign n37005 = ~n37002 | ~n37201;
  assign n37004 = ~n37003 | ~n37025;
  assign n37006 = n37005 & n37004;
  assign P3_U2845 = ~n37007 | ~n37006;
  assign n37033 = ~n37008 & ~n37184;
  assign n37020 = ~n37352 & ~n37033;
  assign n37035 = ~n37009 & ~n38674;
  assign n37011 = ~n22834 | ~P3_INSTADDRPOINTER_REG_15__SCAN_IN;
  assign n37014 = ~n37011 | ~n37010;
  assign n37013 = ~n38730 | ~n37012;
  assign n37017 = ~n37014 | ~n37013;
  assign n37015 = ~n37080 & ~n37062;
  assign n37016 = ~n22828 & ~n37015;
  assign n37040 = ~n37017 & ~n37016;
  assign n37018 = ~n37300 & ~n37040;
  assign n37019 = ~n37035 & ~n37018;
  assign n37021 = ~n37020 | ~n37019;
  assign n37022 = ~n37021 | ~P3_INSTADDRPOINTER_REG_16__SCAN_IN;
  assign n37029 = ~n22843 & ~n37022;
  assign n37027 = ~n37023 | ~n37201;
  assign n37026 = ~n37025 | ~n37024;
  assign n37028 = ~n37027 | ~n37026;
  assign n37031 = ~n37029 & ~n37028;
  assign P3_U2846 = ~n37031 | ~n37030;
  assign n37037 = ~n37033 | ~n37032;
  assign n37036 = ~n37035 | ~n37034;
  assign n37042 = ~n37037 | ~n37036;
  assign n37039 = n37047 & n37038;
  assign n37041 = ~n37040 & ~n37039;
  assign n37043 = ~n37042 & ~n37041;
  assign n37045 = ~n37349 & ~n37043;
  assign n37051 = ~n37045 & ~n37044;
  assign n37049 = ~n37165 & ~n37046;
  assign n37048 = ~n37047 & ~n37383;
  assign n37050 = ~n37049 & ~n37048;
  assign P3_U2847 = ~n37051 | ~n37050;
  assign n37055 = ~n37184 & ~n37052;
  assign n37054 = ~n38674 & ~n37053;
  assign n37075 = ~n37055 & ~n37054;
  assign n37057 = ~n37056 | ~n37105;
  assign n37073 = ~n37057 | ~n37080;
  assign n37221 = ~n37382 & ~n37188;
  assign n37182 = ~n37058 | ~n37221;
  assign n37118 = ~n37059 & ~n37182;
  assign n37061 = ~n22834 & ~n37118;
  assign n37060 = ~n38673 & ~P3_INSTADDRPOINTER_REG_12__SCAN_IN;
  assign n37098 = ~n37061 & ~n37060;
  assign n37063 = ~n38758 | ~n37062;
  assign n37070 = ~P3_INSTADDRPOINTER_REG_14__SCAN_IN | ~n37063;
  assign n37191 = ~n37064 & ~n38673;
  assign n37086 = ~n37065 & ~n38673;
  assign n37068 = ~n37191 & ~n37086;
  assign n37067 = ~n37066 | ~n37358;
  assign n37069 = ~n37068 | ~n37067;
  assign n37071 = ~n37070 & ~n37069;
  assign n37072 = ~n37098 | ~n37071;
  assign n37074 = ~n37073 | ~n37072;
  assign n37076 = ~n37075 | ~n37074;
  assign n37084 = ~n37076 | ~n24731;
  assign n37078 = ~n37201 | ~n37077;
  assign n37082 = ~n37079 | ~n37078;
  assign n37081 = ~n37080 & ~n37383;
  assign n37083 = ~n37082 & ~n37081;
  assign P3_U2848 = ~n37084 | ~n37083;
  assign n37115 = ~n37085 | ~n38758;
  assign n37097 = ~n37115 | ~n37383;
  assign n37090 = ~n37086;
  assign n37088 = ~n37087 | ~n37140;
  assign n37089 = ~n38758 | ~n37088;
  assign n37150 = ~n37090 | ~n37089;
  assign n37092 = ~n37091 & ~n37184;
  assign n37096 = ~n37150 & ~n37092;
  assign n37094 = ~n37093 & ~n38674;
  assign n37095 = ~n37094 & ~n37191;
  assign n37120 = ~n37096 | ~n37095;
  assign n37099 = ~n37097 & ~n37120;
  assign n37100 = ~n37099 | ~n37098;
  assign n37101 = ~P3_INSTADDRPOINTER_REG_13__SCAN_IN | ~n37100;
  assign n37111 = ~n22843 & ~n37101;
  assign n37103 = ~n37183 | ~n37147;
  assign n37102 = ~n37292 | ~n37185;
  assign n37104 = ~n37103 | ~n37102;
  assign n37122 = ~n37105 & ~n37104;
  assign n37207 = ~n37122 & ~n37349;
  assign n37109 = ~n37106 | ~n37207;
  assign n37108 = ~n37107 | ~n37201;
  assign n37110 = ~n37109 | ~n37108;
  assign n37114 = ~n37111 & ~n37110;
  assign n37113 = ~n37112;
  assign P3_U2849 = ~n37114 | ~n37113;
  assign n37116 = ~n22834 | ~n37115;
  assign n37117 = ~n37123 & ~n37116;
  assign n37119 = ~n37118 & ~n37117;
  assign n37127 = ~n37120 & ~n37119;
  assign n37156 = ~n37122 & ~n37121;
  assign n37124 = ~n37156 | ~P3_INSTADDRPOINTER_REG_11__SCAN_IN;
  assign n37125 = ~n37124 | ~n37123;
  assign n37126 = ~n37125 | ~n24731;
  assign n37132 = ~n37127 & ~n37126;
  assign n37129 = ~n37201 | ~n37128;
  assign n37131 = ~n37130 | ~n37129;
  assign n37134 = ~n37132 & ~n37131;
  assign n37133 = ~n37352 | ~P3_INSTADDRPOINTER_REG_12__SCAN_IN;
  assign P3_U2850 = ~n37134 | ~n37133;
  assign n37137 = ~P3_INSTADDRPOINTER_REG_11__SCAN_IN | ~n37352;
  assign n37136 = ~n37201 | ~n37135;
  assign n37139 = ~n37137 | ~n37136;
  assign n37161 = ~n37139 & ~n37138;
  assign n37169 = P3_INSTADDRPOINTER_REG_9__SCAN_IN & n37140;
  assign n37141 = ~P3_INSTADDRPOINTER_REG_0__SCAN_IN | ~n37169;
  assign n37144 = ~n37141 | ~n38757;
  assign n37143 = ~n37292 | ~n37142;
  assign n37145 = ~n37144 | ~n37143;
  assign n37149 = ~n37191 & ~n37145;
  assign n37148 = ~n37147 | ~n37146;
  assign n37168 = ~n37149 | ~n37148;
  assign n37153 = ~n37150 & ~n37168;
  assign n37152 = ~n38757 | ~n37151;
  assign n37155 = ~n37153 | ~n37152;
  assign n37158 = ~n37155 & ~n37154;
  assign n37157 = ~P3_INSTADDRPOINTER_REG_11__SCAN_IN & ~n37156;
  assign n37159 = ~n37158 & ~n37157;
  assign n37160 = ~n24731 | ~n37159;
  assign P3_U2851 = ~n37161 | ~n37160;
  assign n37163 = ~n37207;
  assign n37167 = ~n37163 & ~n37162;
  assign n37166 = ~n37165 & ~n37164;
  assign n37179 = ~n37167 & ~n37166;
  assign n37173 = ~n37168 & ~n37352;
  assign n37171 = ~n22828 & ~n37169;
  assign n37170 = ~n38673 & ~P3_INSTADDRPOINTER_REG_9__SCAN_IN;
  assign n37172 = ~n37171 & ~n37170;
  assign n37174 = ~n37173 | ~n37172;
  assign n37175 = ~n37174 | ~P3_INSTADDRPOINTER_REG_10__SCAN_IN;
  assign n37176 = ~n22843 & ~n37175;
  assign n37178 = ~n37177 & ~n37176;
  assign P3_U2852 = ~n37179 | ~n37178;
  assign n37180 = ~n38757 & ~n37210;
  assign n37181 = ~n37338 & ~n37180;
  assign n37196 = ~n37182 | ~n37181;
  assign n37187 = ~n37184 & ~n37183;
  assign n37186 = ~n37185 & ~n38674;
  assign n37193 = ~n37187 & ~n37186;
  assign n37189 = ~n37235 & ~n37188;
  assign n37217 = ~n22828 & ~n37189;
  assign n37192 = ~n37191 & ~n37217;
  assign n37194 = ~n37193 | ~n37192;
  assign n37195 = ~n37352 & ~n37194;
  assign n37198 = ~n37196 | ~n37195;
  assign n37199 = ~n37198 | ~n37197;
  assign n37205 = ~n37199 & ~n37206;
  assign n37202 = ~n37201 | ~n37200;
  assign n37204 = ~n37203 | ~n37202;
  assign n37209 = ~n37205 & ~n37204;
  assign n37208 = ~n37207 | ~n37206;
  assign P3_U2853 = ~n37209 | ~n37208;
  assign n37232 = ~n37210 & ~n37383;
  assign n37216 = ~P3_INSTADDRPOINTER_REG_8__SCAN_IN & ~n37211;
  assign n37214 = ~n37213 ^ n37212;
  assign n37215 = ~n37363 & ~n37214;
  assign n37226 = ~n37216 & ~n37215;
  assign n37220 = ~n37217 & ~n37235;
  assign n37219 = ~n38730 | ~n37218;
  assign n37223 = ~n37220 | ~n37219;
  assign n37222 = ~n22834 & ~n37221;
  assign n37241 = ~n37223 & ~n37222;
  assign n37224 = ~n37300 & ~n37241;
  assign n37225 = ~P3_INSTADDRPOINTER_REG_8__SCAN_IN | ~n37224;
  assign n37229 = ~n37226 | ~n37225;
  assign n37228 = ~n37227 & ~n38674;
  assign n37230 = ~n37229 & ~n37228;
  assign n37231 = ~n37349 & ~n37230;
  assign n37234 = ~n37232 & ~n37231;
  assign P3_U2854 = ~n37234 | ~n37233;
  assign n37236 = ~n37235 & ~n37383;
  assign n37249 = ~n37237 & ~n37236;
  assign n37246 = ~n37238 | ~n37292;
  assign n37240 = ~P3_INSTADDRPOINTER_REG_7__SCAN_IN & ~n37239;
  assign n37244 = ~n37241 & ~n37240;
  assign n37243 = ~n37242 & ~n37363;
  assign n37245 = ~n37244 & ~n37243;
  assign n37247 = ~n37246 | ~n37245;
  assign n37248 = ~n37247 | ~n24731;
  assign P3_U2855 = ~n37249 | ~n37248;
  assign n37271 = ~n37257 & ~n37383;
  assign n37253 = ~n37250 | ~n38678;
  assign n37252 = ~n37251 | ~n37292;
  assign n37268 = ~n37253 | ~n37252;
  assign n37255 = ~n38673 & ~n37294;
  assign n37254 = ~n37295 & ~n37334;
  assign n37316 = ~n37255 & ~n37254;
  assign n37258 = ~n37316 & ~n37256;
  assign n37266 = ~n37258 | ~n37257;
  assign n37262 = ~n37259 & ~n37338;
  assign n37261 = ~n38673 & ~n37260;
  assign n37264 = ~n37262 & ~n37261;
  assign n37280 = ~n37264 | ~n37263;
  assign n37265 = ~P3_INSTADDRPOINTER_REG_6__SCAN_IN | ~n37280;
  assign n37267 = ~n37266 | ~n37265;
  assign n37269 = ~n37268 & ~n37267;
  assign n37270 = ~n37349 & ~n37269;
  assign n37273 = ~n37271 & ~n37270;
  assign P3_U2856 = ~n37273 | ~n37272;
  assign n37277 = ~n37274 | ~n38678;
  assign n37276 = ~n37275 | ~n37292;
  assign n37284 = ~n37277 | ~n37276;
  assign n37279 = ~P3_INSTADDRPOINTER_REG_5__SCAN_IN & ~n37316;
  assign n37282 = ~n37279 | ~n37278;
  assign n37281 = ~P3_INSTADDRPOINTER_REG_5__SCAN_IN | ~n37280;
  assign n37283 = ~n37282 | ~n37281;
  assign n37285 = ~n37284 & ~n37283;
  assign n37286 = ~n37349 & ~n37285;
  assign n37289 = ~n37287 & ~n37286;
  assign n37288 = ~n37352 | ~P3_INSTADDRPOINTER_REG_5__SCAN_IN;
  assign P3_U2857 = ~n37289 | ~n37288;
  assign n37290 = ~n37302 & ~n37383;
  assign n37313 = ~n37291 & ~n37290;
  assign n37310 = ~n37293 | ~n37292;
  assign n37330 = ~n37382 & ~n37295;
  assign n37298 = ~n22834 & ~n37330;
  assign n37345 = ~n38730 | ~n37294;
  assign n37296 = ~n38758 | ~n37295;
  assign n37297 = ~n37345 | ~n37296;
  assign n37299 = ~n37298 & ~n37297;
  assign n37318 = ~P3_INSTADDRPOINTER_REG_3__SCAN_IN | ~n37299;
  assign n37301 = ~n37300 & ~n37302;
  assign n37305 = ~n37318 | ~n37301;
  assign n37303 = ~n37316 & ~n37317;
  assign n37304 = ~n37303 | ~n37302;
  assign n37308 = ~n37305 | ~n37304;
  assign n37307 = ~n37363 & ~n37306;
  assign n37309 = ~n37308 & ~n37307;
  assign n37311 = ~n37310 | ~n37309;
  assign n37312 = ~n37311 | ~n24731;
  assign P3_U2858 = ~n37313 | ~n37312;
  assign n37314 = ~n37317 & ~n37383;
  assign n37328 = ~n37315 & ~n37314;
  assign n37319 = ~n37317 | ~n37316;
  assign n37325 = ~n37319 | ~n37318;
  assign n37323 = ~n37363 & ~n37320;
  assign n37322 = ~n38674 & ~n37321;
  assign n37324 = ~n37323 & ~n37322;
  assign n37326 = ~n37325 | ~n37324;
  assign n37327 = ~n24731 | ~n37326;
  assign P3_U2859 = ~n37328 | ~n37327;
  assign n37347 = ~n37329 & ~n38674;
  assign n37333 = ~n37330 | ~n38730;
  assign n37332 = ~n38678 | ~n37331;
  assign n37343 = ~n37333 | ~n37332;
  assign n37335 = ~P3_INSTADDRPOINTER_REG_2__SCAN_IN & ~n37334;
  assign n37341 = ~n37335 | ~P3_INSTADDRPOINTER_REG_1__SCAN_IN;
  assign n37337 = ~n37336 & ~n37369;
  assign n37339 = ~n37338 & ~n37337;
  assign n37340 = ~P3_INSTADDRPOINTER_REG_2__SCAN_IN | ~n37339;
  assign n37342 = ~n37341 | ~n37340;
  assign n37344 = ~n37343 & ~n37342;
  assign n37346 = ~n37345 | ~n37344;
  assign n37348 = ~n37347 & ~n37346;
  assign n37351 = ~n37349 & ~n37348;
  assign n37354 = ~n37351 & ~n37350;
  assign n37353 = ~P3_INSTADDRPOINTER_REG_2__SCAN_IN | ~n37352;
  assign P3_U2860 = ~n37354 | ~n37353;
  assign n37357 = ~n37356 | ~n37355;
  assign n37360 = ~n37369 | ~n37357;
  assign n37380 = ~n37382 | ~n37358;
  assign n37359 = ~P3_INSTADDRPOINTER_REG_1__SCAN_IN | ~n37380;
  assign n37367 = ~n37360 | ~n37359;
  assign n37365 = ~n38674 & ~n37361;
  assign n37364 = ~n37363 & ~n37362;
  assign n37366 = ~n37365 & ~n37364;
  assign n37368 = ~n37367 | ~n37366;
  assign n37373 = ~n37368 | ~n24731;
  assign n37370 = ~n37369 & ~n37383;
  assign n37372 = ~n37371 & ~n37370;
  assign P3_U2861 = ~n37373 | ~n37372;
  assign n37378 = ~n38674 & ~n37374;
  assign n37376 = ~P3_INSTADDRPOINTER_REG_0__SCAN_IN | ~n38758;
  assign n37375 = ~n38678 | ~n37374;
  assign n37377 = ~n37376 | ~n37375;
  assign n37379 = ~n37378 & ~n37377;
  assign n37381 = ~n37380 | ~n37379;
  assign n37387 = ~n37381 | ~n24731;
  assign n37384 = ~n37383 & ~n37382;
  assign n37386 = ~n37385 & ~n37384;
  assign P3_U2862 = ~n37387 | ~n37386;
  assign n37388 = ~P3_FLUSH_REG_SCAN_IN;
  assign n39026 = n39118 | n37396;
  assign n39028 = ~n37388 & ~n39026;
  assign n37390 = ~n23642 | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n38667 = ~n37390 | ~n37389;
  assign n37394 = ~n35252 & ~n38667;
  assign n37391 = ~n37394 & ~n39026;
  assign n37392 = ~n39028 & ~n37391;
  assign n37435 = ~n37392 | ~n38489;
  assign n37393 = ~n37435 | ~n39104;
  assign n37400 = ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN | ~n37393;
  assign n37395 = ~n37394 & ~P3_FLUSH_REG_SCAN_IN;
  assign n38805 = ~n37396 & ~n37395;
  assign n37397 = ~n38805;
  assign n37525 = ~P3_STATE2_REG_3__SCAN_IN | ~n24681;
  assign n37398 = ~n37397 | ~n37525;
  assign n37399 = ~n37435 | ~n37398;
  assign P3_U2863 = ~n37400 | ~n37399;
  assign n37402 = ~n37401 & ~n39104;
  assign n37425 = ~n37402 | ~n37435;
  assign n37406 = ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & ~n37425;
  assign n38180 = ~n38768 & ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n37414 = ~n37435;
  assign n37813 = ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN | ~n38768;
  assign n37403 = ~n37414 & ~n37813;
  assign n37404 = ~n38180 & ~n37403;
  assign n37405 = ~n38487 & ~n37404;
  assign n37409 = ~n37406 & ~n37405;
  assign n37407 = ~n37441 | ~n37435;
  assign n37408 = ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~n37407;
  assign P3_U2864 = ~n37409 | ~n37408;
  assign n37412 = ~n37441 & ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign n37440 = ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign n37419 = ~n37440;
  assign n37416 = ~n38487 & ~n37419;
  assign n37410 = ~n37416;
  assign n38761 = ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n37411 = ~n37410 & ~n38761;
  assign n37413 = ~n37412 & ~n37411;
  assign n37418 = ~n37414 & ~n37413;
  assign n37415 = ~n37525 | ~n37435;
  assign n37423 = ~n37416 & ~n37415;
  assign n37417 = ~n37428 & ~n37423;
  assign n37422 = ~n37418 & ~n37417;
  assign n37420 = ~n37419 & ~n37425;
  assign n37437 = ~n38768 | ~n37428;
  assign n37421 = ~n37420 | ~n37437;
  assign P3_U2865 = ~n37422 | ~n37421;
  assign n37427 = ~n38781 & ~n37423;
  assign n37424 = P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN ^ n37440;
  assign n37426 = ~n37425 & ~n37424;
  assign n37434 = ~n37427 & ~n37426;
  assign n38114 = ~n37440 & ~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN;
  assign n37431 = ~P3_STATE2_REG_3__SCAN_IN | ~n38248;
  assign n37674 = ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & ~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN;
  assign n37429 = ~n37674 & ~n37441;
  assign n38403 = ~n37428 & ~n38781;
  assign n38328 = ~n38403;
  assign n37430 = ~n37429 | ~n38328;
  assign n37432 = ~n37431 | ~n37430;
  assign n37433 = ~n37435 | ~n37432;
  assign P3_U2866 = ~n37434 | ~n37433;
  assign P3_U2867 = ~n38686 & ~n37435;
  assign n39029 = ~P3_STATE2_REG_0__SCAN_IN & ~n38487;
  assign n38557 = ~n39110 & ~n37501;
  assign n38033 = ~n37437;
  assign n37532 = ~n38033 | ~n38781;
  assign n37732 = ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & ~n37532;
  assign n37439 = ~n38557 | ~n37732;
  assign n38558 = ~BUF2_REG_24__SCAN_IN | ~n38115;
  assign n38458 = ~n37813 & ~n38328;
  assign n37438 = n38558 | n38654;
  assign n37448 = ~n37439 | ~n37438;
  assign n38559 = ~n38781 & ~n37440;
  assign n38652 = ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN | ~n38559;
  assign n38640 = ~n38652;
  assign n37595 = ~n38180;
  assign n38182 = ~n37813 | ~n37595;
  assign n38485 = ~n38403 | ~n38182;
  assign n37442 = ~n37441 & ~n38485;
  assign n37443 = ~n38640 & ~n37442;
  assign n37444 = ~P3_STATE2_REG_3__SCAN_IN & ~n37443;
  assign n37445 = ~n37732 & ~n37444;
  assign n37506 = ~n38489 & ~n37445;
  assign n37447 = ~n37506 & ~n37446;
  assign n37452 = ~n37448 & ~n37447;
  assign n38568 = ~n38559;
  assign n38556 = ~BUF2_REG_16__SCAN_IN | ~n38115;
  assign n37450 = ~n38545 & ~n38556;
  assign n38560 = ~BUF2_REG_0__SCAN_IN | ~n38340;
  assign n37724 = ~n37732;
  assign n37598 = ~n38652 | ~n37724;
  assign n37513 = ~n38814 | ~n37598;
  assign n37449 = ~n38560 & ~n37513;
  assign n37451 = ~n37450 & ~n37449;
  assign P3_U2868 = ~n37452 | ~n37451;
  assign n38579 = ~n37453 & ~n37501;
  assign n37455 = ~n38579 | ~n37732;
  assign n38576 = ~BUF2_REG_25__SCAN_IN | ~n38115;
  assign n37454 = n38576 | n38654;
  assign n37458 = ~n37455 | ~n37454;
  assign n37457 = ~n37506 & ~n37456;
  assign n37462 = ~n37458 & ~n37457;
  assign n38582 = ~BUF2_REG_17__SCAN_IN | ~n38115;
  assign n37460 = ~n38582 & ~n38545;
  assign n38575 = ~BUF2_REG_1__SCAN_IN | ~n38340;
  assign n37459 = ~n37513 & ~n38575;
  assign n37461 = ~n37460 & ~n37459;
  assign P3_U2869 = ~n37462 | ~n37461;
  assign n38591 = ~n37463 & ~n37501;
  assign n37465 = ~n38591 | ~n37732;
  assign n38594 = ~BUF2_REG_26__SCAN_IN | ~n38115;
  assign n37464 = n38594 | n38654;
  assign n37468 = ~n37465 | ~n37464;
  assign n37466 = ~P3_INSTQUEUE_REG_0__2__SCAN_IN;
  assign n37467 = ~n37506 & ~n37466;
  assign n37472 = ~n37468 & ~n37467;
  assign n38588 = ~BUF2_REG_18__SCAN_IN | ~n38115;
  assign n37470 = ~n38588 & ~n38545;
  assign n38587 = ~BUF2_REG_2__SCAN_IN | ~n38340;
  assign n37469 = ~n37513 & ~n38587;
  assign n37471 = ~n37470 & ~n37469;
  assign P3_U2870 = ~n37472 | ~n37471;
  assign n38599 = ~BUF2_REG_3__SCAN_IN | ~n38340;
  assign n37477 = ~n38599 & ~n37513;
  assign n38600 = ~BUF2_REG_27__SCAN_IN | ~n38115;
  assign n37475 = n38654 | n38600;
  assign n38603 = ~n37473 & ~n37501;
  assign n37474 = ~n37732 | ~n38603;
  assign n37476 = ~n37475 | ~n37474;
  assign n37481 = ~n37477 & ~n37476;
  assign n37522 = ~n37506;
  assign n37479 = n37522 & P3_INSTQUEUE_REG_0__3__SCAN_IN;
  assign n38606 = ~BUF2_REG_19__SCAN_IN | ~n38115;
  assign n37478 = ~n38545 & ~n38606;
  assign n37480 = ~n37479 & ~n37478;
  assign P3_U2871 = ~n37481 | ~n37480;
  assign n38611 = ~BUF2_REG_4__SCAN_IN | ~n38340;
  assign n37486 = ~n38611 & ~n37513;
  assign n38612 = ~BUF2_REG_28__SCAN_IN | ~n38115;
  assign n37484 = n38654 | n38612;
  assign n38615 = ~n37482 & ~n37501;
  assign n37483 = ~n37732 | ~n38615;
  assign n37485 = ~n37484 | ~n37483;
  assign n37491 = ~n37486 & ~n37485;
  assign n37487 = ~P3_INSTQUEUE_REG_0__4__SCAN_IN;
  assign n37489 = ~n37506 & ~n37487;
  assign n38618 = ~BUF2_REG_20__SCAN_IN | ~n38115;
  assign n37488 = ~n38545 & ~n38618;
  assign n37490 = ~n37489 & ~n37488;
  assign P3_U2872 = ~n37491 | ~n37490;
  assign n38627 = ~n40515 & ~n38570;
  assign n37493 = ~n38458 | ~n38627;
  assign n37492 = ~P3_INSTQUEUE_REG_0__5__SCAN_IN | ~n37522;
  assign n37496 = ~n37493 | ~n37492;
  assign n37515 = ~n37501;
  assign n38630 = ~n37515 | ~n37494;
  assign n37495 = ~n37724 & ~n38630;
  assign n37500 = ~n37496 & ~n37495;
  assign n38624 = ~BUF2_REG_21__SCAN_IN | ~n38115;
  assign n37498 = ~n38624 & ~n38545;
  assign n38623 = ~BUF2_REG_5__SCAN_IN | ~n38340;
  assign n37497 = ~n37513 & ~n38623;
  assign n37499 = ~n37498 & ~n37497;
  assign P3_U2873 = ~n37500 | ~n37499;
  assign n38641 = ~n37502 & ~n37501;
  assign n37504 = ~n38641 | ~n37732;
  assign n38637 = ~BUF2_REG_30__SCAN_IN | ~n38115;
  assign n37503 = n38637 | n38654;
  assign n37508 = ~n37504 | ~n37503;
  assign n37507 = ~n37506 & ~n37505;
  assign n37512 = ~n37508 & ~n37507;
  assign n38644 = ~BUF2_REG_22__SCAN_IN | ~n38115;
  assign n37510 = ~n38644 & ~n38545;
  assign n38635 = ~BUF2_REG_6__SCAN_IN | ~n38340;
  assign n37509 = ~n37513 & ~n38635;
  assign n37511 = ~n37510 & ~n37509;
  assign P3_U2874 = ~n37512 | ~n37511;
  assign n38653 = ~BUF2_REG_23__SCAN_IN | ~n38115;
  assign n37521 = ~n38545 & ~n38653;
  assign n38650 = ~BUF2_REG_7__SCAN_IN | ~n38340;
  assign n37517 = ~n37513 & ~n38650;
  assign n38651 = ~n37515 | ~n37514;
  assign n37516 = ~n37724 & ~n38651;
  assign n37519 = ~n37517 & ~n37516;
  assign n38658 = ~n40548 & ~n38570;
  assign n37518 = ~n38458 | ~n38658;
  assign n37520 = ~n37519 | ~n37518;
  assign n37524 = ~n37521 & ~n37520;
  assign n37523 = ~P3_INSTQUEUE_REG_0__7__SCAN_IN | ~n37522;
  assign P3_U2875 = ~n37524 | ~n37523;
  assign n37529 = ~n37805 | ~n38557;
  assign n38567 = ~n38340 | ~n37525;
  assign n37527 = ~n37532 & ~n38567;
  assign n37526 = ~n38570 & ~n38568;
  assign n37588 = ~n37527 & ~n37526;
  assign n37528 = ~n37588 | ~P3_INSTQUEUE_REG_1__0__SCAN_IN;
  assign n37531 = ~n37529 | ~n37528;
  assign n37530 = ~n38652 & ~n38556;
  assign n37536 = ~n37531 & ~n37530;
  assign n37534 = ~n38545 & ~n38558;
  assign n37585 = n37532 | n38476;
  assign n37533 = ~n38560 & ~n37585;
  assign n37535 = ~n37534 & ~n37533;
  assign P3_U2876 = ~n37536 | ~n37535;
  assign n37538 = ~n38575 & ~n37585;
  assign n37537 = ~n38652 & ~n38582;
  assign n37544 = ~n37538 & ~n37537;
  assign n37540 = ~n37805 | ~n38579;
  assign n37539 = ~n37588 | ~P3_INSTQUEUE_REG_1__1__SCAN_IN;
  assign n37542 = ~n37540 | ~n37539;
  assign n37541 = ~n38545 & ~n38576;
  assign n37543 = ~n37542 & ~n37541;
  assign P3_U2877 = ~n37544 | ~n37543;
  assign n37546 = ~n38587 & ~n37585;
  assign n37545 = ~n38652 & ~n38588;
  assign n37552 = ~n37546 & ~n37545;
  assign n37548 = ~n37805 | ~n38591;
  assign n37547 = ~n37588 | ~P3_INSTQUEUE_REG_1__2__SCAN_IN;
  assign n37550 = ~n37548 | ~n37547;
  assign n37549 = ~n38545 & ~n38594;
  assign n37551 = ~n37550 & ~n37549;
  assign P3_U2878 = ~n37552 | ~n37551;
  assign n37554 = ~n37805 | ~n38603;
  assign n37553 = ~n37588 | ~P3_INSTQUEUE_REG_1__3__SCAN_IN;
  assign n37556 = ~n37554 | ~n37553;
  assign n37555 = ~n38652 & ~n38606;
  assign n37560 = ~n37556 & ~n37555;
  assign n37558 = ~n38600 & ~n38545;
  assign n37557 = ~n38599 & ~n37585;
  assign n37559 = ~n37558 & ~n37557;
  assign P3_U2879 = ~n37560 | ~n37559;
  assign n37562 = ~n37805 | ~n38615;
  assign n37561 = ~n37588 | ~P3_INSTQUEUE_REG_1__4__SCAN_IN;
  assign n37564 = ~n37562 | ~n37561;
  assign n37563 = ~n38652 & ~n38618;
  assign n37568 = ~n37564 & ~n37563;
  assign n37566 = ~n38612 & ~n38545;
  assign n37565 = ~n38611 & ~n37585;
  assign n37567 = ~n37566 & ~n37565;
  assign P3_U2880 = ~n37568 | ~n37567;
  assign n37574 = ~n38652 & ~n38624;
  assign n37570 = ~n38623 & ~n37585;
  assign n37569 = ~n38630 & ~n37797;
  assign n37572 = ~n37570 & ~n37569;
  assign n37571 = ~n38627 | ~n38537;
  assign n37573 = ~n37572 | ~n37571;
  assign n37576 = ~n37574 & ~n37573;
  assign n37575 = ~n37588 | ~P3_INSTQUEUE_REG_1__5__SCAN_IN;
  assign P3_U2881 = ~n37576 | ~n37575;
  assign n37578 = ~n37805 | ~n38641;
  assign n37577 = ~n37588 | ~P3_INSTQUEUE_REG_1__6__SCAN_IN;
  assign n37580 = ~n37578 | ~n37577;
  assign n37579 = ~n38652 & ~n38644;
  assign n37584 = ~n37580 & ~n37579;
  assign n37582 = ~n38637 & ~n38545;
  assign n37581 = ~n38635 & ~n37585;
  assign n37583 = ~n37582 & ~n37581;
  assign P3_U2882 = ~n37584 | ~n37583;
  assign n37587 = ~n38650 & ~n37585;
  assign n37586 = ~n38652 & ~n38653;
  assign n37594 = ~n37587 & ~n37586;
  assign n37590 = ~n38658 | ~n38537;
  assign n37589 = ~n37588 | ~P3_INSTQUEUE_REG_1__7__SCAN_IN;
  assign n37592 = ~n37590 | ~n37589;
  assign n37591 = ~n38651 & ~n37797;
  assign n37593 = ~n37592 & ~n37591;
  assign P3_U2883 = ~n37594 | ~n37593;
  assign n37740 = ~n37797 | ~n37870;
  assign n37657 = ~n38814 | ~n37740;
  assign n37597 = ~n38560 & ~n37657;
  assign n37596 = ~n37724 & ~n38556;
  assign n37608 = ~n37597 & ~n37596;
  assign n37604 = ~n38557 | ~n37878;
  assign n37599 = ~n38483 | ~n37598;
  assign n37600 = ~n37797 | ~n37599;
  assign n37601 = ~n37600 | ~n38487;
  assign n37602 = ~n37601 | ~n37870;
  assign n37664 = ~n38340 | ~n37602;
  assign n37603 = ~P3_INSTQUEUE_REG_2__0__SCAN_IN | ~n37664;
  assign n37606 = ~n37604 | ~n37603;
  assign n37605 = ~n38558 & ~n38652;
  assign n37607 = ~n37606 & ~n37605;
  assign P3_U2884 = ~n37608 | ~n37607;
  assign n37610 = ~n38575 & ~n37657;
  assign n37609 = ~n38652 & ~n38576;
  assign n37616 = ~n37610 & ~n37609;
  assign n37612 = ~n38579 | ~n37878;
  assign n37611 = ~P3_INSTQUEUE_REG_2__1__SCAN_IN | ~n37664;
  assign n37614 = ~n37612 | ~n37611;
  assign n37613 = ~n37724 & ~n38582;
  assign n37615 = ~n37614 & ~n37613;
  assign P3_U2885 = ~n37616 | ~n37615;
  assign n37618 = ~n38587 & ~n37657;
  assign n37617 = ~n38652 & ~n38594;
  assign n37624 = ~n37618 & ~n37617;
  assign n37620 = ~n38591 | ~n37878;
  assign n37619 = ~P3_INSTQUEUE_REG_2__2__SCAN_IN | ~n37664;
  assign n37622 = ~n37620 | ~n37619;
  assign n37621 = ~n37724 & ~n38588;
  assign n37623 = ~n37622 & ~n37621;
  assign P3_U2886 = ~n37624 | ~n37623;
  assign n37626 = ~n38599 & ~n37657;
  assign n37625 = ~n38652 & ~n38600;
  assign n37632 = ~n37626 & ~n37625;
  assign n37628 = ~n38603 | ~n37878;
  assign n37627 = ~P3_INSTQUEUE_REG_2__3__SCAN_IN | ~n37664;
  assign n37630 = ~n37628 | ~n37627;
  assign n37629 = ~n37724 & ~n38606;
  assign n37631 = ~n37630 & ~n37629;
  assign P3_U2887 = ~n37632 | ~n37631;
  assign n37634 = ~n38611 & ~n37657;
  assign n37633 = ~n38652 & ~n38612;
  assign n37640 = ~n37634 & ~n37633;
  assign n37636 = ~n38615 | ~n37878;
  assign n37635 = ~P3_INSTQUEUE_REG_2__4__SCAN_IN | ~n37664;
  assign n37638 = ~n37636 | ~n37635;
  assign n37637 = ~n37724 & ~n38618;
  assign n37639 = ~n37638 & ~n37637;
  assign P3_U2888 = ~n37640 | ~n37639;
  assign n37642 = ~n38623 & ~n37657;
  assign n37641 = ~n37724 & ~n38624;
  assign n37648 = ~n37642 & ~n37641;
  assign n37644 = ~n38640 | ~n38627;
  assign n37643 = ~P3_INSTQUEUE_REG_2__5__SCAN_IN | ~n37664;
  assign n37646 = ~n37644 | ~n37643;
  assign n37645 = ~n38630 & ~n37870;
  assign n37647 = ~n37646 & ~n37645;
  assign P3_U2889 = ~n37648 | ~n37647;
  assign n37650 = ~n38635 & ~n37657;
  assign n37649 = ~n37724 & ~n38644;
  assign n37656 = ~n37650 & ~n37649;
  assign n37652 = ~n38641 | ~n37878;
  assign n37651 = ~P3_INSTQUEUE_REG_2__6__SCAN_IN | ~n37664;
  assign n37654 = ~n37652 | ~n37651;
  assign n37653 = ~n38652 & ~n38637;
  assign n37655 = ~n37654 & ~n37653;
  assign P3_U2890 = ~n37656 | ~n37655;
  assign n37663 = ~n38650 & ~n37657;
  assign n37659 = ~n38651 & ~n37870;
  assign n37658 = ~n37724 & ~n38653;
  assign n37661 = ~n37659 & ~n37658;
  assign n37660 = ~n38640 | ~n38658;
  assign n37662 = ~n37661 | ~n37660;
  assign n37666 = ~n37663 & ~n37662;
  assign n37665 = ~P3_INSTQUEUE_REG_2__7__SCAN_IN | ~n37664;
  assign P3_U2891 = ~n37666 | ~n37665;
  assign n37673 = ~n38558 & ~n37724;
  assign n37814 = ~n38768 & ~n37667;
  assign n37953 = ~n37941;
  assign n37671 = ~n38557 | ~n37953;
  assign n37729 = ~n37814 | ~n38814;
  assign n37669 = ~n38560 & ~n37729;
  assign n37668 = ~n38556 & ~n37797;
  assign n37670 = ~n37669 & ~n37668;
  assign n37672 = ~n37671 | ~n37670;
  assign n37679 = ~n37673 & ~n37672;
  assign n37675 = ~n38487 | ~n37674;
  assign n37677 = ~n37675 | ~n37941;
  assign n37676 = ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & ~n38483;
  assign n37970 = ~n38489 & ~n37676;
  assign n37733 = ~n37677 | ~n37970;
  assign n37678 = ~P3_INSTQUEUE_REG_3__0__SCAN_IN | ~n37733;
  assign P3_U2892 = ~n37679 | ~n37678;
  assign n37681 = ~n38575 & ~n37729;
  assign n37680 = ~n38582 & ~n37797;
  assign n37687 = ~n37681 & ~n37680;
  assign n37683 = ~n38579 | ~n37953;
  assign n37682 = ~P3_INSTQUEUE_REG_3__1__SCAN_IN | ~n37733;
  assign n37685 = ~n37683 | ~n37682;
  assign n37684 = ~n37724 & ~n38576;
  assign n37686 = ~n37685 & ~n37684;
  assign P3_U2893 = ~n37687 | ~n37686;
  assign n37691 = ~n38587 & ~n37729;
  assign n37689 = ~n38591 | ~n37953;
  assign n37688 = ~P3_INSTQUEUE_REG_3__2__SCAN_IN | ~n37733;
  assign n37690 = ~n37689 | ~n37688;
  assign n37695 = ~n37691 & ~n37690;
  assign n37693 = ~n38588 & ~n37797;
  assign n37692 = ~n37724 & ~n38594;
  assign n37694 = ~n37693 & ~n37692;
  assign P3_U2894 = ~n37695 | ~n37694;
  assign n37697 = ~n38599 & ~n37729;
  assign n37696 = ~n38606 & ~n37797;
  assign n37703 = ~n37697 & ~n37696;
  assign n37699 = ~n38603 | ~n37953;
  assign n37698 = ~P3_INSTQUEUE_REG_3__3__SCAN_IN | ~n37733;
  assign n37701 = ~n37699 | ~n37698;
  assign n37700 = ~n37724 & ~n38600;
  assign n37702 = ~n37701 & ~n37700;
  assign P3_U2895 = ~n37703 | ~n37702;
  assign n37707 = ~n38611 & ~n37729;
  assign n37705 = ~n38615 | ~n37953;
  assign n37704 = ~P3_INSTQUEUE_REG_3__4__SCAN_IN | ~n37733;
  assign n37706 = ~n37705 | ~n37704;
  assign n37711 = ~n37707 & ~n37706;
  assign n37709 = ~n38618 & ~n37797;
  assign n37708 = ~n37724 & ~n38612;
  assign n37710 = ~n37709 & ~n37708;
  assign P3_U2896 = ~n37711 | ~n37710;
  assign n37717 = ~n38623 & ~n37729;
  assign n37713 = ~n38624 & ~n37797;
  assign n37712 = ~n38630 & ~n37941;
  assign n37715 = ~n37713 & ~n37712;
  assign n37714 = ~P3_INSTQUEUE_REG_3__5__SCAN_IN | ~n37733;
  assign n37716 = ~n37715 | ~n37714;
  assign n37719 = ~n37717 & ~n37716;
  assign n37718 = ~n37732 | ~n38627;
  assign P3_U2897 = ~n37719 | ~n37718;
  assign n37723 = ~n38635 & ~n37729;
  assign n37721 = ~n38641 | ~n37953;
  assign n37720 = ~P3_INSTQUEUE_REG_3__6__SCAN_IN | ~n37733;
  assign n37722 = ~n37721 | ~n37720;
  assign n37728 = ~n37723 & ~n37722;
  assign n37726 = ~n38644 & ~n37797;
  assign n37725 = ~n37724 & ~n38637;
  assign n37727 = ~n37726 & ~n37725;
  assign P3_U2898 = ~n37728 | ~n37727;
  assign n37731 = ~n38650 & ~n37729;
  assign n37730 = ~n38653 & ~n37797;
  assign n37739 = ~n37731 & ~n37730;
  assign n37735 = ~n37732 | ~n38658;
  assign n37734 = ~P3_INSTQUEUE_REG_3__7__SCAN_IN | ~n37733;
  assign n37737 = ~n37735 | ~n37734;
  assign n37736 = ~n38651 & ~n37941;
  assign n37738 = ~n37737 & ~n37736;
  assign P3_U2899 = ~n37739 | ~n37738;
  assign n38776 = ~n38768 | ~n24681;
  assign n37968 = ~n38781 | ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign n37889 = ~n37941 | ~n38017;
  assign n37802 = ~n38814 | ~n37889;
  assign n37748 = ~n37802 & ~n38560;
  assign n37741 = ~n38483 | ~n37740;
  assign n37742 = ~n37941 | ~n37741;
  assign n37743 = ~n37742 | ~n38487;
  assign n37744 = ~n37743 | ~n38017;
  assign n37806 = ~n38340 | ~n37744;
  assign n37746 = ~P3_INSTQUEUE_REG_4__0__SCAN_IN | ~n37806;
  assign n37745 = ~n38557 | ~n38025;
  assign n37747 = ~n37746 | ~n37745;
  assign n37752 = ~n37748 & ~n37747;
  assign n37750 = ~n38556 & ~n37870;
  assign n37749 = ~n38558 & ~n37797;
  assign n37751 = ~n37750 & ~n37749;
  assign P3_U2900 = ~n37752 | ~n37751;
  assign n37754 = ~n38575 & ~n37802;
  assign n37753 = ~n38576 & ~n37797;
  assign n37760 = ~n37754 & ~n37753;
  assign n37756 = ~n38579 | ~n38025;
  assign n37755 = ~P3_INSTQUEUE_REG_4__1__SCAN_IN | ~n37806;
  assign n37758 = ~n37756 | ~n37755;
  assign n37757 = ~n38582 & ~n37870;
  assign n37759 = ~n37758 & ~n37757;
  assign P3_U2901 = ~n37760 | ~n37759;
  assign n37764 = ~n38587 & ~n37802;
  assign n37762 = ~n38591 | ~n38025;
  assign n37761 = ~P3_INSTQUEUE_REG_4__2__SCAN_IN | ~n37806;
  assign n37763 = ~n37762 | ~n37761;
  assign n37768 = ~n37764 & ~n37763;
  assign n37766 = ~n38588 & ~n37870;
  assign n37765 = ~n38594 & ~n37797;
  assign n37767 = ~n37766 & ~n37765;
  assign P3_U2902 = ~n37768 | ~n37767;
  assign n37772 = ~n38599 & ~n37802;
  assign n37770 = ~n38603 | ~n38025;
  assign n37769 = ~P3_INSTQUEUE_REG_4__3__SCAN_IN | ~n37806;
  assign n37771 = ~n37770 | ~n37769;
  assign n37776 = ~n37772 & ~n37771;
  assign n37774 = ~n38600 & ~n37797;
  assign n37773 = ~n38606 & ~n37870;
  assign n37775 = ~n37774 & ~n37773;
  assign P3_U2903 = ~n37776 | ~n37775;
  assign n37780 = ~n38611 & ~n37802;
  assign n37778 = ~n38615 | ~n38025;
  assign n37777 = ~P3_INSTQUEUE_REG_4__4__SCAN_IN | ~n37806;
  assign n37779 = ~n37778 | ~n37777;
  assign n37784 = ~n37780 & ~n37779;
  assign n37782 = ~n38612 & ~n37797;
  assign n37781 = ~n38618 & ~n37870;
  assign n37783 = ~n37782 & ~n37781;
  assign P3_U2904 = ~n37784 | ~n37783;
  assign n37786 = ~n38623 & ~n37802;
  assign n37785 = ~n38624 & ~n37870;
  assign n37792 = ~n37786 & ~n37785;
  assign n37788 = ~n38627 | ~n37805;
  assign n37787 = ~P3_INSTQUEUE_REG_4__5__SCAN_IN | ~n37806;
  assign n37790 = ~n37788 | ~n37787;
  assign n37789 = ~n38630 & ~n38017;
  assign n37791 = ~n37790 & ~n37789;
  assign P3_U2905 = ~n37792 | ~n37791;
  assign n37796 = ~n38635 & ~n37802;
  assign n37794 = ~n38641 | ~n38025;
  assign n37793 = ~P3_INSTQUEUE_REG_4__6__SCAN_IN | ~n37806;
  assign n37795 = ~n37794 | ~n37793;
  assign n37801 = ~n37796 & ~n37795;
  assign n37799 = ~n38644 & ~n37870;
  assign n37798 = ~n38637 & ~n37797;
  assign n37800 = ~n37799 & ~n37798;
  assign P3_U2906 = ~n37801 | ~n37800;
  assign n37804 = ~n38650 & ~n37802;
  assign n37803 = ~n38653 & ~n37870;
  assign n37812 = ~n37804 & ~n37803;
  assign n37808 = ~n38658 | ~n37805;
  assign n37807 = ~P3_INSTQUEUE_REG_4__7__SCAN_IN | ~n37806;
  assign n37810 = ~n37808 | ~n37807;
  assign n37809 = ~n38651 & ~n38017;
  assign n37811 = ~n37810 & ~n37809;
  assign P3_U2907 = ~n37812 | ~n37811;
  assign n38099 = ~n37813 & ~n37968;
  assign n37818 = ~n38099 | ~n38557;
  assign n37886 = ~n37968;
  assign n37821 = ~n37886 | ~n38768;
  assign n37816 = ~n38567 & ~n37821;
  assign n37815 = n38115 & n37814;
  assign n37883 = ~n37816 & ~n37815;
  assign n37817 = ~n37883 | ~P3_INSTQUEUE_REG_5__0__SCAN_IN;
  assign n37820 = ~n37818 | ~n37817;
  assign n37819 = ~n38558 & ~n37870;
  assign n37825 = ~n37820 & ~n37819;
  assign n37875 = n37821 | n38476;
  assign n37823 = ~n38560 & ~n37875;
  assign n37822 = ~n38556 & ~n37941;
  assign n37824 = ~n37823 & ~n37822;
  assign P3_U2908 = ~n37825 | ~n37824;
  assign n37827 = ~n38575 & ~n37875;
  assign n37826 = ~n38576 & ~n37870;
  assign n37833 = ~n37827 & ~n37826;
  assign n37829 = ~n38099 | ~n38579;
  assign n37828 = ~n37883 | ~P3_INSTQUEUE_REG_5__1__SCAN_IN;
  assign n37831 = ~n37829 | ~n37828;
  assign n37830 = ~n38582 & ~n37941;
  assign n37832 = ~n37831 & ~n37830;
  assign P3_U2909 = ~n37833 | ~n37832;
  assign n37835 = ~n38587 & ~n37875;
  assign n37834 = ~n38588 & ~n37941;
  assign n37841 = ~n37835 & ~n37834;
  assign n37837 = ~n38099 | ~n38591;
  assign n37836 = ~n37883 | ~P3_INSTQUEUE_REG_5__2__SCAN_IN;
  assign n37839 = ~n37837 | ~n37836;
  assign n37838 = ~n38594 & ~n37870;
  assign n37840 = ~n37839 & ~n37838;
  assign P3_U2910 = ~n37841 | ~n37840;
  assign n37843 = ~n38599 & ~n37875;
  assign n37842 = ~n38600 & ~n37870;
  assign n37849 = ~n37843 & ~n37842;
  assign n37845 = ~n38099 | ~n38603;
  assign n37844 = ~n37883 | ~P3_INSTQUEUE_REG_5__3__SCAN_IN;
  assign n37847 = ~n37845 | ~n37844;
  assign n37846 = ~n38606 & ~n37941;
  assign n37848 = ~n37847 & ~n37846;
  assign P3_U2911 = ~n37849 | ~n37848;
  assign n37851 = ~n38611 & ~n37875;
  assign n37850 = ~n38612 & ~n37870;
  assign n37857 = ~n37851 & ~n37850;
  assign n37853 = ~n38099 | ~n38615;
  assign n37852 = ~n37883 | ~P3_INSTQUEUE_REG_5__4__SCAN_IN;
  assign n37855 = ~n37853 | ~n37852;
  assign n37854 = ~n38618 & ~n37941;
  assign n37856 = ~n37855 & ~n37854;
  assign P3_U2912 = ~n37857 | ~n37856;
  assign n37859 = ~n38623 & ~n37875;
  assign n37858 = ~n38624 & ~n37941;
  assign n37865 = ~n37859 & ~n37858;
  assign n37861 = ~n37878 | ~n38627;
  assign n37860 = ~n37883 | ~P3_INSTQUEUE_REG_5__5__SCAN_IN;
  assign n37863 = ~n37861 | ~n37860;
  assign n37862 = ~n38630 & ~n38087;
  assign n37864 = ~n37863 & ~n37862;
  assign P3_U2913 = ~n37865 | ~n37864;
  assign n37867 = ~n38635 & ~n37875;
  assign n37866 = ~n38644 & ~n37941;
  assign n37874 = ~n37867 & ~n37866;
  assign n37869 = ~n38099 | ~n38641;
  assign n37868 = ~n37883 | ~P3_INSTQUEUE_REG_5__6__SCAN_IN;
  assign n37872 = ~n37869 | ~n37868;
  assign n37871 = ~n38637 & ~n37870;
  assign n37873 = ~n37872 & ~n37871;
  assign P3_U2914 = ~n37874 | ~n37873;
  assign n37882 = ~n38650 & ~n37875;
  assign n37877 = ~n38651 & ~n38087;
  assign n37876 = ~n38653 & ~n37941;
  assign n37880 = ~n37877 & ~n37876;
  assign n37879 = ~n38658 | ~n37878;
  assign n37881 = ~n37880 | ~n37879;
  assign n37885 = ~n37882 & ~n37881;
  assign n37884 = ~P3_INSTQUEUE_REG_5__7__SCAN_IN | ~n37883;
  assign P3_U2915 = ~n37885 | ~n37884;
  assign n37898 = ~n38558 & ~n37941;
  assign n37888 = ~n38556 & ~n38017;
  assign n37890 = ~n37886 | ~n38182;
  assign n38036 = ~n37890;
  assign n37950 = ~n38036 | ~n38814;
  assign n37887 = ~n38560 & ~n37950;
  assign n37896 = ~n37888 & ~n37887;
  assign n37891 = ~n37889 | ~n38483;
  assign n37894 = ~n37891 | ~n37890;
  assign n38160 = ~n24681 | ~n38114;
  assign n38172 = ~n38160;
  assign n37892 = ~n38172 & ~n38487;
  assign n37893 = ~n38489 & ~n37892;
  assign n37958 = ~n37894 | ~n37893;
  assign n37895 = ~P3_INSTQUEUE_REG_6__0__SCAN_IN | ~n37958;
  assign n37897 = ~n37896 | ~n37895;
  assign n37900 = ~n37898 & ~n37897;
  assign n37899 = ~n38172 | ~n38557;
  assign P3_U2916 = ~n37900 | ~n37899;
  assign n37902 = ~n38575 & ~n37950;
  assign n37901 = ~n38576 & ~n37941;
  assign n37908 = ~n37902 & ~n37901;
  assign n37904 = ~n38579 | ~n38172;
  assign n37903 = ~P3_INSTQUEUE_REG_6__1__SCAN_IN | ~n37958;
  assign n37906 = ~n37904 | ~n37903;
  assign n37905 = ~n38582 & ~n38017;
  assign n37907 = ~n37906 & ~n37905;
  assign P3_U2917 = ~n37908 | ~n37907;
  assign n37910 = ~n38587 & ~n37950;
  assign n37909 = ~n38588 & ~n38017;
  assign n37916 = ~n37910 & ~n37909;
  assign n37912 = ~n38591 | ~n38172;
  assign n37911 = ~P3_INSTQUEUE_REG_6__2__SCAN_IN | ~n37958;
  assign n37914 = ~n37912 | ~n37911;
  assign n37913 = ~n38594 & ~n37941;
  assign n37915 = ~n37914 & ~n37913;
  assign P3_U2918 = ~n37916 | ~n37915;
  assign n37918 = ~n38599 & ~n37950;
  assign n37917 = ~n38600 & ~n37941;
  assign n37924 = ~n37918 & ~n37917;
  assign n37920 = ~n38603 | ~n38172;
  assign n37919 = ~P3_INSTQUEUE_REG_6__3__SCAN_IN | ~n37958;
  assign n37922 = ~n37920 | ~n37919;
  assign n37921 = ~n38606 & ~n38017;
  assign n37923 = ~n37922 & ~n37921;
  assign P3_U2919 = ~n37924 | ~n37923;
  assign n37926 = ~n38611 & ~n37950;
  assign n37925 = ~n38618 & ~n38017;
  assign n37932 = ~n37926 & ~n37925;
  assign n37928 = ~n38615 | ~n38172;
  assign n37927 = ~P3_INSTQUEUE_REG_6__4__SCAN_IN | ~n37958;
  assign n37930 = ~n37928 | ~n37927;
  assign n37929 = ~n38612 & ~n37941;
  assign n37931 = ~n37930 & ~n37929;
  assign P3_U2920 = ~n37932 | ~n37931;
  assign n37934 = ~n38623 & ~n37950;
  assign n37933 = ~n38624 & ~n38017;
  assign n37940 = ~n37934 & ~n37933;
  assign n37936 = ~n38627 | ~n37953;
  assign n37935 = ~P3_INSTQUEUE_REG_6__5__SCAN_IN | ~n37958;
  assign n37938 = ~n37936 | ~n37935;
  assign n37937 = ~n38630 & ~n38160;
  assign n37939 = ~n37938 & ~n37937;
  assign P3_U2921 = ~n37940 | ~n37939;
  assign n37943 = ~n38635 & ~n37950;
  assign n37942 = ~n38637 & ~n37941;
  assign n37949 = ~n37943 & ~n37942;
  assign n37945 = ~n38641 | ~n38172;
  assign n37944 = ~P3_INSTQUEUE_REG_6__6__SCAN_IN | ~n37958;
  assign n37947 = ~n37945 | ~n37944;
  assign n37946 = ~n38644 & ~n38017;
  assign n37948 = ~n37947 & ~n37946;
  assign P3_U2922 = ~n37949 | ~n37948;
  assign n37957 = ~n38650 & ~n37950;
  assign n37952 = ~n38651 & ~n38160;
  assign n37951 = ~n38653 & ~n38017;
  assign n37955 = ~n37952 & ~n37951;
  assign n37954 = ~n38658 | ~n37953;
  assign n37956 = ~n37955 | ~n37954;
  assign n37960 = ~n37957 & ~n37956;
  assign n37959 = ~P3_INSTQUEUE_REG_6__7__SCAN_IN | ~n37958;
  assign P3_U2923 = ~n37960 | ~n37959;
  assign n37966 = ~n38558 & ~n38017;
  assign n37964 = ~n38557 | ~n38248;
  assign n38022 = ~n38114 | ~n38814;
  assign n37962 = ~n38560 & ~n38022;
  assign n37961 = ~n38556 & ~n38087;
  assign n37963 = ~n37962 & ~n37961;
  assign n37965 = ~n37964 | ~n37963;
  assign n37972 = ~n37966 & ~n37965;
  assign n37967 = ~n38248 & ~n38487;
  assign n37969 = ~n37968 & ~n37967;
  assign n38030 = ~n37970 | ~n37969;
  assign n37971 = ~P3_INSTQUEUE_REG_7__0__SCAN_IN | ~n38030;
  assign P3_U2924 = ~n37972 | ~n37971;
  assign n37976 = ~n38575 & ~n38022;
  assign n37974 = ~n38579 | ~n38248;
  assign n37973 = ~P3_INSTQUEUE_REG_7__1__SCAN_IN | ~n38030;
  assign n37975 = ~n37974 | ~n37973;
  assign n37980 = ~n37976 & ~n37975;
  assign n37978 = ~n38582 & ~n38087;
  assign n37977 = ~n38576 & ~n38017;
  assign n37979 = ~n37978 & ~n37977;
  assign P3_U2925 = ~n37980 | ~n37979;
  assign n37984 = ~n38587 & ~n38022;
  assign n37982 = ~n38591 | ~n38248;
  assign n37981 = ~P3_INSTQUEUE_REG_7__2__SCAN_IN | ~n38030;
  assign n37983 = ~n37982 | ~n37981;
  assign n37988 = ~n37984 & ~n37983;
  assign n37986 = ~n38588 & ~n38087;
  assign n37985 = ~n38594 & ~n38017;
  assign n37987 = ~n37986 & ~n37985;
  assign P3_U2926 = ~n37988 | ~n37987;
  assign n37992 = ~n38599 & ~n38022;
  assign n37990 = ~n38603 | ~n38248;
  assign n37989 = ~P3_INSTQUEUE_REG_7__3__SCAN_IN | ~n38030;
  assign n37991 = ~n37990 | ~n37989;
  assign n37996 = ~n37992 & ~n37991;
  assign n37994 = ~n38600 & ~n38017;
  assign n37993 = ~n38606 & ~n38087;
  assign n37995 = ~n37994 & ~n37993;
  assign P3_U2927 = ~n37996 | ~n37995;
  assign n37998 = ~n38611 & ~n38022;
  assign n37997 = ~n38612 & ~n38017;
  assign n38004 = ~n37998 & ~n37997;
  assign n38000 = ~n38615 | ~n38248;
  assign n37999 = ~P3_INSTQUEUE_REG_7__4__SCAN_IN | ~n38030;
  assign n38002 = ~n38000 | ~n37999;
  assign n38001 = ~n38618 & ~n38087;
  assign n38003 = ~n38002 & ~n38001;
  assign P3_U2928 = ~n38004 | ~n38003;
  assign n38006 = ~n38623 & ~n38022;
  assign n38005 = ~n38624 & ~n38087;
  assign n38012 = ~n38006 & ~n38005;
  assign n38008 = ~n38627 | ~n38025;
  assign n38007 = ~P3_INSTQUEUE_REG_7__5__SCAN_IN | ~n38030;
  assign n38010 = ~n38008 | ~n38007;
  assign n38009 = ~n38630 & ~n38240;
  assign n38011 = ~n38010 & ~n38009;
  assign P3_U2929 = ~n38012 | ~n38011;
  assign n38014 = ~n38635 & ~n38022;
  assign n38013 = ~n38644 & ~n38087;
  assign n38021 = ~n38014 & ~n38013;
  assign n38016 = ~n38641 | ~n38248;
  assign n38015 = ~P3_INSTQUEUE_REG_7__6__SCAN_IN | ~n38030;
  assign n38019 = ~n38016 | ~n38015;
  assign n38018 = ~n38637 & ~n38017;
  assign n38020 = ~n38019 & ~n38018;
  assign P3_U2930 = ~n38021 | ~n38020;
  assign n38029 = ~n38650 & ~n38022;
  assign n38024 = ~n38651 & ~n38240;
  assign n38023 = ~n38653 & ~n38087;
  assign n38027 = ~n38024 & ~n38023;
  assign n38026 = ~n38658 | ~n38025;
  assign n38028 = ~n38027 | ~n38026;
  assign n38032 = ~n38029 & ~n38028;
  assign n38031 = ~P3_INSTQUEUE_REG_7__7__SCAN_IN | ~n38030;
  assign P3_U2931 = ~n38032 | ~n38031;
  assign n38263 = ~P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | ~n38033;
  assign n38320 = ~n38263 & ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n38181 = ~n38240 | ~n38308;
  assign n38096 = ~n38814 | ~n38181;
  assign n38035 = ~n38560 & ~n38096;
  assign n38034 = ~n38558 & ~n38087;
  assign n38046 = ~n38035 & ~n38034;
  assign n38042 = ~n38557 | ~n38320;
  assign n38037 = ~n38483 | ~n38036;
  assign n38038 = ~n38037 | ~n38240;
  assign n38039 = ~n38038 | ~n38487;
  assign n38040 = ~n38308 | ~n38039;
  assign n38104 = ~n38340 | ~n38040;
  assign n38041 = ~P3_INSTQUEUE_REG_8__0__SCAN_IN | ~n38104;
  assign n38044 = ~n38042 | ~n38041;
  assign n38043 = ~n38556 & ~n38160;
  assign n38045 = ~n38044 & ~n38043;
  assign P3_U2932 = ~n38046 | ~n38045;
  assign n38048 = ~n38575 & ~n38096;
  assign n38047 = ~n38582 & ~n38160;
  assign n38054 = ~n38048 & ~n38047;
  assign n38050 = ~n38579 | ~n38320;
  assign n38049 = ~P3_INSTQUEUE_REG_8__1__SCAN_IN | ~n38104;
  assign n38052 = ~n38050 | ~n38049;
  assign n38051 = ~n38576 & ~n38087;
  assign n38053 = ~n38052 & ~n38051;
  assign P3_U2933 = ~n38054 | ~n38053;
  assign n38056 = ~n38587 & ~n38096;
  assign n38055 = ~n38594 & ~n38087;
  assign n38062 = ~n38056 & ~n38055;
  assign n38058 = ~n38591 | ~n38320;
  assign n38057 = ~P3_INSTQUEUE_REG_8__2__SCAN_IN | ~n38104;
  assign n38060 = ~n38058 | ~n38057;
  assign n38059 = ~n38588 & ~n38160;
  assign n38061 = ~n38060 & ~n38059;
  assign P3_U2934 = ~n38062 | ~n38061;
  assign n38064 = ~n38599 & ~n38096;
  assign n38063 = ~n38606 & ~n38160;
  assign n38070 = ~n38064 & ~n38063;
  assign n38066 = ~n38603 | ~n38320;
  assign n38065 = ~P3_INSTQUEUE_REG_8__3__SCAN_IN | ~n38104;
  assign n38068 = ~n38066 | ~n38065;
  assign n38067 = ~n38600 & ~n38087;
  assign n38069 = ~n38068 & ~n38067;
  assign P3_U2935 = ~n38070 | ~n38069;
  assign n38072 = ~n38611 & ~n38096;
  assign n38071 = ~n38612 & ~n38087;
  assign n38078 = ~n38072 & ~n38071;
  assign n38074 = ~n38615 | ~n38320;
  assign n38073 = ~P3_INSTQUEUE_REG_8__4__SCAN_IN | ~n38104;
  assign n38076 = ~n38074 | ~n38073;
  assign n38075 = ~n38618 & ~n38160;
  assign n38077 = ~n38076 & ~n38075;
  assign P3_U2936 = ~n38078 | ~n38077;
  assign n38080 = ~n38623 & ~n38096;
  assign n38079 = ~n38624 & ~n38160;
  assign n38086 = ~n38080 & ~n38079;
  assign n38082 = ~n38627 | ~n38099;
  assign n38081 = ~P3_INSTQUEUE_REG_8__5__SCAN_IN | ~n38104;
  assign n38084 = ~n38082 | ~n38081;
  assign n38083 = ~n38630 & ~n38308;
  assign n38085 = ~n38084 & ~n38083;
  assign P3_U2937 = ~n38086 | ~n38085;
  assign n38089 = ~n38635 & ~n38096;
  assign n38088 = ~n38637 & ~n38087;
  assign n38095 = ~n38089 & ~n38088;
  assign n38091 = ~n38641 | ~n38320;
  assign n38090 = ~P3_INSTQUEUE_REG_8__6__SCAN_IN | ~n38104;
  assign n38093 = ~n38091 | ~n38090;
  assign n38092 = ~n38644 & ~n38160;
  assign n38094 = ~n38093 & ~n38092;
  assign P3_U2938 = ~n38095 | ~n38094;
  assign n38103 = ~n38650 & ~n38096;
  assign n38098 = ~n38651 & ~n38308;
  assign n38097 = ~n38653 & ~n38160;
  assign n38101 = ~n38098 & ~n38097;
  assign n38100 = ~n38658 | ~n38099;
  assign n38102 = ~n38101 | ~n38100;
  assign n38106 = ~n38103 & ~n38102;
  assign n38105 = ~P3_INSTQUEUE_REG_8__7__SCAN_IN | ~n38104;
  assign P3_U2939 = ~n38106 | ~n38105;
  assign n38113 = ~n38556 & ~n38240;
  assign n38107 = ~n38263;
  assign n38383 = ~P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN | ~n38107;
  assign n38395 = ~n38383;
  assign n38111 = ~n38557 | ~n38395;
  assign n38109 = ~n38558 & ~n38160;
  assign n38169 = ~n38107 | ~n38814;
  assign n38108 = ~n38560 & ~n38169;
  assign n38110 = ~n38109 & ~n38108;
  assign n38112 = ~n38111 | ~n38110;
  assign n38119 = ~n38113 & ~n38112;
  assign n38117 = ~n38567 & ~n38263;
  assign n38116 = n38115 & n38114;
  assign n38173 = ~n38117 & ~n38116;
  assign n38118 = ~n38173 | ~P3_INSTQUEUE_REG_9__0__SCAN_IN;
  assign P3_U2940 = ~n38119 | ~n38118;
  assign n38121 = ~n38575 & ~n38169;
  assign n38120 = ~n38582 & ~n38240;
  assign n38127 = ~n38121 & ~n38120;
  assign n38123 = ~n38395 | ~n38579;
  assign n38122 = ~n38173 | ~P3_INSTQUEUE_REG_9__1__SCAN_IN;
  assign n38125 = ~n38123 | ~n38122;
  assign n38124 = ~n38576 & ~n38160;
  assign n38126 = ~n38125 & ~n38124;
  assign P3_U2941 = ~n38127 | ~n38126;
  assign n38129 = ~n38587 & ~n38169;
  assign n38128 = ~n38588 & ~n38240;
  assign n38135 = ~n38129 & ~n38128;
  assign n38131 = ~n38395 | ~n38591;
  assign n38130 = ~n38173 | ~P3_INSTQUEUE_REG_9__2__SCAN_IN;
  assign n38133 = ~n38131 | ~n38130;
  assign n38132 = ~n38594 & ~n38160;
  assign n38134 = ~n38133 & ~n38132;
  assign P3_U2942 = ~n38135 | ~n38134;
  assign n38137 = ~n38599 & ~n38169;
  assign n38136 = ~n38600 & ~n38160;
  assign n38143 = ~n38137 & ~n38136;
  assign n38139 = ~n38395 | ~n38603;
  assign n38138 = ~n38173 | ~P3_INSTQUEUE_REG_9__3__SCAN_IN;
  assign n38141 = ~n38139 | ~n38138;
  assign n38140 = ~n38606 & ~n38240;
  assign n38142 = ~n38141 & ~n38140;
  assign P3_U2943 = ~n38143 | ~n38142;
  assign n38145 = ~n38611 & ~n38169;
  assign n38144 = ~n38618 & ~n38240;
  assign n38151 = ~n38145 & ~n38144;
  assign n38147 = ~n38395 | ~n38615;
  assign n38146 = ~n38173 | ~P3_INSTQUEUE_REG_9__4__SCAN_IN;
  assign n38149 = ~n38147 | ~n38146;
  assign n38148 = ~n38612 & ~n38160;
  assign n38150 = ~n38149 & ~n38148;
  assign P3_U2944 = ~n38151 | ~n38150;
  assign n38157 = ~n38624 & ~n38240;
  assign n38153 = ~n38623 & ~n38169;
  assign n38152 = ~n38630 & ~n38383;
  assign n38155 = ~n38153 & ~n38152;
  assign n38154 = ~n38172 | ~n38627;
  assign n38156 = ~n38155 | ~n38154;
  assign n38159 = ~n38157 & ~n38156;
  assign n38158 = ~n38173 | ~P3_INSTQUEUE_REG_9__5__SCAN_IN;
  assign P3_U2945 = ~n38159 | ~n38158;
  assign n38162 = ~n38635 & ~n38169;
  assign n38161 = ~n38637 & ~n38160;
  assign n38168 = ~n38162 & ~n38161;
  assign n38164 = ~n38395 | ~n38641;
  assign n38163 = ~n38173 | ~P3_INSTQUEUE_REG_9__6__SCAN_IN;
  assign n38166 = ~n38164 | ~n38163;
  assign n38165 = ~n38644 & ~n38240;
  assign n38167 = ~n38166 & ~n38165;
  assign P3_U2946 = ~n38168 | ~n38167;
  assign n38171 = ~n38650 & ~n38169;
  assign n38170 = ~n38653 & ~n38240;
  assign n38179 = ~n38171 & ~n38170;
  assign n38175 = ~n38172 | ~n38658;
  assign n38174 = ~n38173 | ~P3_INSTQUEUE_REG_9__7__SCAN_IN;
  assign n38177 = ~n38175 | ~n38174;
  assign n38176 = ~n38651 & ~n38383;
  assign n38178 = ~n38177 & ~n38176;
  assign P3_U2947 = ~n38179 | ~n38178;
  assign n38256 = ~n38781 & ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign n38455 = ~n38180 | ~n38256;
  assign n38188 = ~n38557 | ~n38468;
  assign n38183 = ~n38181 | ~n38483;
  assign n38191 = ~n38256 | ~n38182;
  assign n38186 = ~n38183 | ~n38191;
  assign n38184 = ~n38468 & ~n38487;
  assign n38185 = ~n38489 & ~n38184;
  assign n38253 = ~n38186 | ~n38185;
  assign n38187 = ~P3_INSTQUEUE_REG_10__0__SCAN_IN | ~n38253;
  assign n38190 = ~n38188 | ~n38187;
  assign n38189 = ~n38558 & ~n38240;
  assign n38195 = ~n38190 & ~n38189;
  assign n38335 = ~n38191;
  assign n38245 = ~n38335 | ~n38814;
  assign n38193 = ~n38245 & ~n38560;
  assign n38192 = ~n38556 & ~n38308;
  assign n38194 = ~n38193 & ~n38192;
  assign P3_U2948 = ~n38195 | ~n38194;
  assign n38197 = ~n38575 & ~n38245;
  assign n38196 = ~n38582 & ~n38308;
  assign n38203 = ~n38197 & ~n38196;
  assign n38199 = ~n38579 | ~n38468;
  assign n38198 = ~P3_INSTQUEUE_REG_10__1__SCAN_IN | ~n38253;
  assign n38201 = ~n38199 | ~n38198;
  assign n38200 = ~n38576 & ~n38240;
  assign n38202 = ~n38201 & ~n38200;
  assign P3_U2949 = ~n38203 | ~n38202;
  assign n38205 = ~n38587 & ~n38245;
  assign n38204 = ~n38588 & ~n38308;
  assign n38211 = ~n38205 & ~n38204;
  assign n38207 = ~n38591 | ~n38468;
  assign n38206 = ~P3_INSTQUEUE_REG_10__2__SCAN_IN | ~n38253;
  assign n38209 = ~n38207 | ~n38206;
  assign n38208 = ~n38594 & ~n38240;
  assign n38210 = ~n38209 & ~n38208;
  assign P3_U2950 = ~n38211 | ~n38210;
  assign n38213 = ~n38599 & ~n38245;
  assign n38212 = ~n38600 & ~n38240;
  assign n38219 = ~n38213 & ~n38212;
  assign n38215 = ~n38603 | ~n38468;
  assign n38214 = ~P3_INSTQUEUE_REG_10__3__SCAN_IN | ~n38253;
  assign n38217 = ~n38215 | ~n38214;
  assign n38216 = ~n38606 & ~n38308;
  assign n38218 = ~n38217 & ~n38216;
  assign P3_U2951 = ~n38219 | ~n38218;
  assign n38221 = ~n38611 & ~n38245;
  assign n38220 = ~n38612 & ~n38240;
  assign n38227 = ~n38221 & ~n38220;
  assign n38223 = ~n38615 | ~n38468;
  assign n38222 = ~P3_INSTQUEUE_REG_10__4__SCAN_IN | ~n38253;
  assign n38225 = ~n38223 | ~n38222;
  assign n38224 = ~n38618 & ~n38308;
  assign n38226 = ~n38225 & ~n38224;
  assign P3_U2952 = ~n38227 | ~n38226;
  assign n38229 = ~n38623 & ~n38245;
  assign n38228 = ~n38624 & ~n38308;
  assign n38235 = ~n38229 & ~n38228;
  assign n38231 = ~n38627 | ~n38248;
  assign n38230 = ~P3_INSTQUEUE_REG_10__5__SCAN_IN | ~n38253;
  assign n38233 = ~n38231 | ~n38230;
  assign n38232 = ~n38630 & ~n38455;
  assign n38234 = ~n38233 & ~n38232;
  assign P3_U2953 = ~n38235 | ~n38234;
  assign n38237 = ~n38635 & ~n38245;
  assign n38236 = ~n38644 & ~n38308;
  assign n38244 = ~n38237 & ~n38236;
  assign n38239 = ~n38641 | ~n38468;
  assign n38238 = ~P3_INSTQUEUE_REG_10__6__SCAN_IN | ~n38253;
  assign n38242 = ~n38239 | ~n38238;
  assign n38241 = ~n38637 & ~n38240;
  assign n38243 = ~n38242 & ~n38241;
  assign P3_U2954 = ~n38244 | ~n38243;
  assign n38252 = ~n38650 & ~n38245;
  assign n38247 = ~n38651 & ~n38455;
  assign n38246 = ~n38653 & ~n38308;
  assign n38250 = ~n38247 & ~n38246;
  assign n38249 = ~n38658 | ~n38248;
  assign n38251 = ~n38250 | ~n38249;
  assign n38255 = ~n38252 & ~n38251;
  assign n38254 = ~P3_INSTQUEUE_REG_10__7__SCAN_IN | ~n38253;
  assign P3_U2955 = ~n38255 | ~n38254;
  assign n38262 = ~n38556 & ~n38383;
  assign n38406 = ~P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~n38256;
  assign n38317 = n38406 | n38476;
  assign n38258 = ~n38560 & ~n38317;
  assign n38257 = ~n38558 & ~n38308;
  assign n38260 = ~n38258 & ~n38257;
  assign n38548 = ~n24681 & ~n38406;
  assign n38259 = ~n38548 | ~n38557;
  assign n38261 = ~n38260 | ~n38259;
  assign n38267 = ~n38262 & ~n38261;
  assign n38265 = ~n38567 & ~n38406;
  assign n38264 = ~n38263 & ~n38570;
  assign n38325 = ~n38265 & ~n38264;
  assign n38266 = ~P3_INSTQUEUE_REG_11__0__SCAN_IN | ~n38325;
  assign P3_U2956 = ~n38267 | ~n38266;
  assign n38269 = ~n38575 & ~n38317;
  assign n38268 = ~n38576 & ~n38308;
  assign n38275 = ~n38269 & ~n38268;
  assign n38271 = ~n38548 | ~n38579;
  assign n38270 = ~n38325 | ~P3_INSTQUEUE_REG_11__1__SCAN_IN;
  assign n38273 = ~n38271 | ~n38270;
  assign n38272 = ~n38582 & ~n38383;
  assign n38274 = ~n38273 & ~n38272;
  assign P3_U2957 = ~n38275 | ~n38274;
  assign n38277 = ~n38587 & ~n38317;
  assign n38276 = ~n38588 & ~n38383;
  assign n38283 = ~n38277 & ~n38276;
  assign n38279 = ~n38548 | ~n38591;
  assign n38278 = ~n38325 | ~P3_INSTQUEUE_REG_11__2__SCAN_IN;
  assign n38281 = ~n38279 | ~n38278;
  assign n38280 = ~n38594 & ~n38308;
  assign n38282 = ~n38281 & ~n38280;
  assign P3_U2958 = ~n38283 | ~n38282;
  assign n38285 = ~n38599 & ~n38317;
  assign n38284 = ~n38600 & ~n38308;
  assign n38291 = ~n38285 & ~n38284;
  assign n38287 = ~n38548 | ~n38603;
  assign n38286 = ~n38325 | ~P3_INSTQUEUE_REG_11__3__SCAN_IN;
  assign n38289 = ~n38287 | ~n38286;
  assign n38288 = ~n38606 & ~n38383;
  assign n38290 = ~n38289 & ~n38288;
  assign P3_U2959 = ~n38291 | ~n38290;
  assign n38293 = ~n38611 & ~n38317;
  assign n38292 = ~n38618 & ~n38383;
  assign n38299 = ~n38293 & ~n38292;
  assign n38295 = ~n38548 | ~n38615;
  assign n38294 = ~n38325 | ~P3_INSTQUEUE_REG_11__4__SCAN_IN;
  assign n38297 = ~n38295 | ~n38294;
  assign n38296 = ~n38612 & ~n38308;
  assign n38298 = ~n38297 & ~n38296;
  assign P3_U2960 = ~n38299 | ~n38298;
  assign n38305 = ~n38624 & ~n38383;
  assign n38301 = ~n38623 & ~n38317;
  assign n38300 = ~n38630 & ~n38534;
  assign n38303 = ~n38301 & ~n38300;
  assign n38302 = ~n38320 | ~n38627;
  assign n38304 = ~n38303 | ~n38302;
  assign n38307 = ~n38305 & ~n38304;
  assign n38306 = ~n38325 | ~P3_INSTQUEUE_REG_11__5__SCAN_IN;
  assign P3_U2961 = ~n38307 | ~n38306;
  assign n38310 = ~n38635 & ~n38317;
  assign n38309 = ~n38637 & ~n38308;
  assign n38316 = ~n38310 & ~n38309;
  assign n38312 = ~n38548 | ~n38641;
  assign n38311 = ~n38325 | ~P3_INSTQUEUE_REG_11__6__SCAN_IN;
  assign n38314 = ~n38312 | ~n38311;
  assign n38313 = ~n38644 & ~n38383;
  assign n38315 = ~n38314 & ~n38313;
  assign P3_U2962 = ~n38316 | ~n38315;
  assign n38324 = ~n38650 & ~n38317;
  assign n38319 = ~n38651 & ~n38534;
  assign n38318 = ~n38653 & ~n38383;
  assign n38322 = ~n38319 & ~n38318;
  assign n38321 = ~n38658 | ~n38320;
  assign n38323 = ~n38322 | ~n38321;
  assign n38327 = ~n38324 & ~n38323;
  assign n38326 = ~P3_INSTQUEUE_REG_11__7__SCAN_IN | ~n38325;
  assign P3_U2963 = ~n38327 | ~n38326;
  assign n38334 = ~n38558 & ~n38383;
  assign n38657 = ~n38776 & ~n38328;
  assign n38332 = ~n38557 | ~n38657;
  assign n38636 = ~n38657;
  assign n38484 = ~n38534 | ~n38636;
  assign n38392 = ~n38814 | ~n38484;
  assign n38330 = ~n38560 & ~n38392;
  assign n38329 = ~n38556 & ~n38455;
  assign n38331 = ~n38330 & ~n38329;
  assign n38333 = ~n38332 | ~n38331;
  assign n38342 = ~n38334 & ~n38333;
  assign n38336 = ~n38483 | ~n38335;
  assign n38337 = ~n38534 | ~n38336;
  assign n38338 = ~n38337 | ~n38487;
  assign n38339 = ~n38338 | ~n38636;
  assign n38396 = ~n38340 | ~n38339;
  assign n38341 = ~P3_INSTQUEUE_REG_12__0__SCAN_IN | ~n38396;
  assign P3_U2964 = ~n38342 | ~n38341;
  assign n38344 = ~n38575 & ~n38392;
  assign n38343 = ~n38582 & ~n38455;
  assign n38350 = ~n38344 & ~n38343;
  assign n38346 = ~n38579 | ~n38657;
  assign n38345 = ~P3_INSTQUEUE_REG_12__1__SCAN_IN | ~n38396;
  assign n38348 = ~n38346 | ~n38345;
  assign n38347 = ~n38576 & ~n38383;
  assign n38349 = ~n38348 & ~n38347;
  assign P3_U2965 = ~n38350 | ~n38349;
  assign n38354 = ~n38587 & ~n38392;
  assign n38352 = ~n38591 | ~n38657;
  assign n38351 = ~P3_INSTQUEUE_REG_12__2__SCAN_IN | ~n38396;
  assign n38353 = ~n38352 | ~n38351;
  assign n38358 = ~n38354 & ~n38353;
  assign n38356 = ~n38588 & ~n38455;
  assign n38355 = ~n38594 & ~n38383;
  assign n38357 = ~n38356 & ~n38355;
  assign P3_U2966 = ~n38358 | ~n38357;
  assign n38360 = ~n38599 & ~n38392;
  assign n38359 = ~n38600 & ~n38383;
  assign n38366 = ~n38360 & ~n38359;
  assign n38362 = ~n38603 | ~n38657;
  assign n38361 = ~P3_INSTQUEUE_REG_12__3__SCAN_IN | ~n38396;
  assign n38364 = ~n38362 | ~n38361;
  assign n38363 = ~n38606 & ~n38455;
  assign n38365 = ~n38364 & ~n38363;
  assign P3_U2967 = ~n38366 | ~n38365;
  assign n38368 = ~n38611 & ~n38392;
  assign n38367 = ~n38618 & ~n38455;
  assign n38374 = ~n38368 & ~n38367;
  assign n38370 = ~n38615 | ~n38657;
  assign n38369 = ~P3_INSTQUEUE_REG_12__4__SCAN_IN | ~n38396;
  assign n38372 = ~n38370 | ~n38369;
  assign n38371 = ~n38612 & ~n38383;
  assign n38373 = ~n38372 & ~n38371;
  assign P3_U2968 = ~n38374 | ~n38373;
  assign n38380 = ~n38623 & ~n38392;
  assign n38376 = ~n38624 & ~n38455;
  assign n38375 = ~n38630 & ~n38636;
  assign n38378 = ~n38376 & ~n38375;
  assign n38377 = ~n38627 | ~n38395;
  assign n38379 = ~n38378 | ~n38377;
  assign n38382 = ~n38380 & ~n38379;
  assign n38381 = ~P3_INSTQUEUE_REG_12__5__SCAN_IN | ~n38396;
  assign P3_U2969 = ~n38382 | ~n38381;
  assign n38385 = ~n38635 & ~n38392;
  assign n38384 = ~n38637 & ~n38383;
  assign n38391 = ~n38385 & ~n38384;
  assign n38387 = ~n38641 | ~n38657;
  assign n38386 = ~P3_INSTQUEUE_REG_12__6__SCAN_IN | ~n38396;
  assign n38389 = ~n38387 | ~n38386;
  assign n38388 = ~n38644 & ~n38455;
  assign n38390 = ~n38389 & ~n38388;
  assign P3_U2970 = ~n38391 | ~n38390;
  assign n38394 = ~n38650 & ~n38392;
  assign n38393 = ~n38653 & ~n38455;
  assign n38402 = ~n38394 & ~n38393;
  assign n38398 = ~n38658 | ~n38395;
  assign n38397 = ~P3_INSTQUEUE_REG_12__7__SCAN_IN | ~n38396;
  assign n38400 = ~n38398 | ~n38397;
  assign n38399 = ~n38651 & ~n38636;
  assign n38401 = ~n38400 & ~n38399;
  assign P3_U2971 = ~n38402 | ~n38401;
  assign n38569 = ~n38768 | ~n38403;
  assign n38465 = n38569 | n38476;
  assign n38405 = ~n38560 & ~n38465;
  assign n38404 = ~n38558 & ~n38455;
  assign n38414 = ~n38405 & ~n38404;
  assign n38410 = ~n38557 | ~n38458;
  assign n38408 = ~n38567 & ~n38569;
  assign n38407 = ~n38406 & ~n38570;
  assign n38469 = ~n38408 & ~n38407;
  assign n38409 = ~n38469 | ~P3_INSTQUEUE_REG_13__0__SCAN_IN;
  assign n38412 = ~n38410 | ~n38409;
  assign n38411 = ~n38556 & ~n38534;
  assign n38413 = ~n38412 & ~n38411;
  assign P3_U2972 = ~n38414 | ~n38413;
  assign n38416 = ~n38575 & ~n38465;
  assign n38415 = ~n38582 & ~n38534;
  assign n38422 = ~n38416 & ~n38415;
  assign n38418 = ~n38579 | ~n38458;
  assign n38417 = ~n38469 | ~P3_INSTQUEUE_REG_13__1__SCAN_IN;
  assign n38420 = ~n38418 | ~n38417;
  assign n38419 = ~n38576 & ~n38455;
  assign n38421 = ~n38420 & ~n38419;
  assign P3_U2973 = ~n38422 | ~n38421;
  assign n38424 = ~n38587 & ~n38465;
  assign n38423 = ~n38594 & ~n38455;
  assign n38430 = ~n38424 & ~n38423;
  assign n38426 = ~n38591 | ~n38458;
  assign n38425 = ~n38469 | ~P3_INSTQUEUE_REG_13__2__SCAN_IN;
  assign n38428 = ~n38426 | ~n38425;
  assign n38427 = ~n38588 & ~n38534;
  assign n38429 = ~n38428 & ~n38427;
  assign P3_U2974 = ~n38430 | ~n38429;
  assign n38432 = ~n38599 & ~n38465;
  assign n38431 = ~n38606 & ~n38534;
  assign n38438 = ~n38432 & ~n38431;
  assign n38434 = ~n38603 | ~n38458;
  assign n38433 = ~n38469 | ~P3_INSTQUEUE_REG_13__3__SCAN_IN;
  assign n38436 = ~n38434 | ~n38433;
  assign n38435 = ~n38600 & ~n38455;
  assign n38437 = ~n38436 & ~n38435;
  assign P3_U2975 = ~n38438 | ~n38437;
  assign n38440 = ~n38611 & ~n38465;
  assign n38439 = ~n38612 & ~n38455;
  assign n38446 = ~n38440 & ~n38439;
  assign n38442 = ~n38615 | ~n38458;
  assign n38441 = ~n38469 | ~P3_INSTQUEUE_REG_13__4__SCAN_IN;
  assign n38444 = ~n38442 | ~n38441;
  assign n38443 = ~n38618 & ~n38534;
  assign n38445 = ~n38444 & ~n38443;
  assign P3_U2976 = ~n38446 | ~n38445;
  assign n38448 = ~n38623 & ~n38465;
  assign n38447 = ~n38624 & ~n38534;
  assign n38454 = ~n38448 & ~n38447;
  assign n38450 = ~n38468 | ~n38627;
  assign n38449 = ~n38469 | ~P3_INSTQUEUE_REG_13__5__SCAN_IN;
  assign n38452 = ~n38450 | ~n38449;
  assign n38451 = ~n38654 & ~n38630;
  assign n38453 = ~n38452 & ~n38451;
  assign P3_U2977 = ~n38454 | ~n38453;
  assign n38457 = ~n38635 & ~n38465;
  assign n38456 = ~n38637 & ~n38455;
  assign n38464 = ~n38457 & ~n38456;
  assign n38460 = ~n38641 | ~n38458;
  assign n38459 = ~n38469 | ~P3_INSTQUEUE_REG_13__6__SCAN_IN;
  assign n38462 = ~n38460 | ~n38459;
  assign n38461 = ~n38644 & ~n38534;
  assign n38463 = ~n38462 & ~n38461;
  assign P3_U2978 = ~n38464 | ~n38463;
  assign n38467 = ~n38650 & ~n38465;
  assign n38466 = ~n38653 & ~n38534;
  assign n38475 = ~n38467 & ~n38466;
  assign n38471 = ~n38468 | ~n38658;
  assign n38470 = ~n38469 | ~P3_INSTQUEUE_REG_13__7__SCAN_IN;
  assign n38473 = ~n38471 | ~n38470;
  assign n38472 = ~n38654 & ~n38651;
  assign n38474 = ~n38473 & ~n38472;
  assign P3_U2979 = ~n38475 | ~n38474;
  assign n38482 = ~n38558 & ~n38534;
  assign n38544 = n38485 | n38476;
  assign n38478 = ~n38560 & ~n38544;
  assign n38477 = ~n38556 & ~n38636;
  assign n38480 = ~n38478 & ~n38477;
  assign n38479 = ~n38537 | ~n38557;
  assign n38481 = ~n38480 | ~n38479;
  assign n38493 = ~n38482 & ~n38481;
  assign n38486 = ~n38484 | ~n38483;
  assign n38491 = ~n38486 | ~n38485;
  assign n38488 = ~n38537 & ~n38487;
  assign n38490 = ~n38489 & ~n38488;
  assign n38553 = ~n38491 | ~n38490;
  assign n38492 = ~P3_INSTQUEUE_REG_14__0__SCAN_IN | ~n38553;
  assign P3_U2980 = ~n38493 | ~n38492;
  assign n38495 = ~n38575 & ~n38544;
  assign n38494 = ~n38576 & ~n38534;
  assign n38501 = ~n38495 & ~n38494;
  assign n38497 = ~n38537 | ~n38579;
  assign n38496 = ~P3_INSTQUEUE_REG_14__1__SCAN_IN | ~n38553;
  assign n38499 = ~n38497 | ~n38496;
  assign n38498 = ~n38582 & ~n38636;
  assign n38500 = ~n38499 & ~n38498;
  assign P3_U2981 = ~n38501 | ~n38500;
  assign n38503 = ~n38587 & ~n38544;
  assign n38502 = ~n38588 & ~n38636;
  assign n38509 = ~n38503 & ~n38502;
  assign n38505 = ~n38537 | ~n38591;
  assign n38504 = ~P3_INSTQUEUE_REG_14__2__SCAN_IN | ~n38553;
  assign n38507 = ~n38505 | ~n38504;
  assign n38506 = ~n38594 & ~n38534;
  assign n38508 = ~n38507 & ~n38506;
  assign P3_U2982 = ~n38509 | ~n38508;
  assign n38511 = ~n38599 & ~n38544;
  assign n38510 = ~n38600 & ~n38534;
  assign n38517 = ~n38511 & ~n38510;
  assign n38513 = ~n38537 | ~n38603;
  assign n38512 = ~P3_INSTQUEUE_REG_14__3__SCAN_IN | ~n38553;
  assign n38515 = ~n38513 | ~n38512;
  assign n38514 = ~n38606 & ~n38636;
  assign n38516 = ~n38515 & ~n38514;
  assign P3_U2983 = ~n38517 | ~n38516;
  assign n38519 = ~n38611 & ~n38544;
  assign n38518 = ~n38612 & ~n38534;
  assign n38525 = ~n38519 & ~n38518;
  assign n38521 = ~n38537 | ~n38615;
  assign n38520 = ~P3_INSTQUEUE_REG_14__4__SCAN_IN | ~n38553;
  assign n38523 = ~n38521 | ~n38520;
  assign n38522 = ~n38618 & ~n38636;
  assign n38524 = ~n38523 & ~n38522;
  assign P3_U2984 = ~n38525 | ~n38524;
  assign n38527 = ~n38623 & ~n38544;
  assign n38526 = ~n38624 & ~n38636;
  assign n38533 = ~n38527 & ~n38526;
  assign n38529 = ~n38627 | ~n38548;
  assign n38528 = ~P3_INSTQUEUE_REG_14__5__SCAN_IN | ~n38553;
  assign n38531 = ~n38529 | ~n38528;
  assign n38530 = ~n38545 & ~n38630;
  assign n38532 = ~n38531 & ~n38530;
  assign P3_U2985 = ~n38533 | ~n38532;
  assign n38536 = ~n38635 & ~n38544;
  assign n38535 = ~n38637 & ~n38534;
  assign n38543 = ~n38536 & ~n38535;
  assign n38539 = ~n38537 | ~n38641;
  assign n38538 = ~P3_INSTQUEUE_REG_14__6__SCAN_IN | ~n38553;
  assign n38541 = ~n38539 | ~n38538;
  assign n38540 = ~n38644 & ~n38636;
  assign n38542 = ~n38541 & ~n38540;
  assign P3_U2986 = ~n38543 | ~n38542;
  assign n38552 = ~n38650 & ~n38544;
  assign n38547 = ~n38653 & ~n38636;
  assign n38546 = ~n38545 & ~n38651;
  assign n38550 = ~n38547 & ~n38546;
  assign n38549 = ~n38658 | ~n38548;
  assign n38551 = ~n38550 | ~n38549;
  assign n38555 = ~n38552 & ~n38551;
  assign n38554 = ~P3_INSTQUEUE_REG_14__7__SCAN_IN | ~n38553;
  assign P3_U2987 = ~n38555 | ~n38554;
  assign n38566 = ~n38654 & ~n38556;
  assign n38564 = ~n38640 | ~n38557;
  assign n38562 = ~n38558 & ~n38636;
  assign n38649 = ~n38559 | ~n38814;
  assign n38561 = ~n38560 & ~n38649;
  assign n38563 = ~n38562 & ~n38561;
  assign n38565 = ~n38564 | ~n38563;
  assign n38574 = ~n38566 & ~n38565;
  assign n38572 = ~n38568 & ~n38567;
  assign n38571 = ~n38570 & ~n38569;
  assign n38663 = ~n38572 & ~n38571;
  assign n38573 = ~P3_INSTQUEUE_REG_15__0__SCAN_IN | ~n38663;
  assign P3_U2988 = ~n38574 | ~n38573;
  assign n38578 = ~n38575 & ~n38649;
  assign n38577 = ~n38576 & ~n38636;
  assign n38586 = ~n38578 & ~n38577;
  assign n38581 = ~n38579 | ~n38640;
  assign n38580 = ~n38663 | ~P3_INSTQUEUE_REG_15__1__SCAN_IN;
  assign n38584 = ~n38581 | ~n38580;
  assign n38583 = ~n38654 & ~n38582;
  assign n38585 = ~n38584 & ~n38583;
  assign P3_U2989 = ~n38586 | ~n38585;
  assign n38590 = ~n38587 & ~n38649;
  assign n38589 = ~n38654 & ~n38588;
  assign n38598 = ~n38590 & ~n38589;
  assign n38593 = ~n38591 | ~n38640;
  assign n38592 = ~n38663 | ~P3_INSTQUEUE_REG_15__2__SCAN_IN;
  assign n38596 = ~n38593 | ~n38592;
  assign n38595 = ~n38594 & ~n38636;
  assign n38597 = ~n38596 & ~n38595;
  assign P3_U2990 = ~n38598 | ~n38597;
  assign n38602 = ~n38599 & ~n38649;
  assign n38601 = ~n38600 & ~n38636;
  assign n38610 = ~n38602 & ~n38601;
  assign n38605 = ~n38603 | ~n38640;
  assign n38604 = ~n38663 | ~P3_INSTQUEUE_REG_15__3__SCAN_IN;
  assign n38608 = ~n38605 | ~n38604;
  assign n38607 = ~n38654 & ~n38606;
  assign n38609 = ~n38608 & ~n38607;
  assign P3_U2991 = ~n38610 | ~n38609;
  assign n38614 = ~n38611 & ~n38649;
  assign n38613 = ~n38612 & ~n38636;
  assign n38622 = ~n38614 & ~n38613;
  assign n38617 = ~n38615 | ~n38640;
  assign n38616 = ~n38663 | ~P3_INSTQUEUE_REG_15__4__SCAN_IN;
  assign n38620 = ~n38617 | ~n38616;
  assign n38619 = ~n38654 & ~n38618;
  assign n38621 = ~n38620 & ~n38619;
  assign P3_U2992 = ~n38622 | ~n38621;
  assign n38626 = ~n38623 & ~n38649;
  assign n38625 = ~n38654 & ~n38624;
  assign n38634 = ~n38626 & ~n38625;
  assign n38629 = ~n38657 | ~n38627;
  assign n38628 = ~n38663 | ~P3_INSTQUEUE_REG_15__5__SCAN_IN;
  assign n38632 = ~n38629 | ~n38628;
  assign n38631 = ~n38652 & ~n38630;
  assign n38633 = ~n38632 & ~n38631;
  assign P3_U2993 = ~n38634 | ~n38633;
  assign n38639 = ~n38635 & ~n38649;
  assign n38638 = ~n38637 & ~n38636;
  assign n38648 = ~n38639 & ~n38638;
  assign n38643 = ~n38641 | ~n38640;
  assign n38642 = ~n38663 | ~P3_INSTQUEUE_REG_15__6__SCAN_IN;
  assign n38646 = ~n38643 | ~n38642;
  assign n38645 = ~n38654 & ~n38644;
  assign n38647 = ~n38646 & ~n38645;
  assign P3_U2994 = ~n38648 | ~n38647;
  assign n38662 = ~n38650 & ~n38649;
  assign n38656 = ~n38652 & ~n38651;
  assign n38655 = ~n38654 & ~n38653;
  assign n38660 = ~n38656 & ~n38655;
  assign n38659 = ~n38658 | ~n38657;
  assign n38661 = ~n38660 | ~n38659;
  assign n38665 = ~n38662 & ~n38661;
  assign n38664 = ~P3_INSTQUEUE_REG_15__7__SCAN_IN | ~n38663;
  assign P3_U2995 = ~n38665 | ~n38664;
  assign n38666 = ~n38763;
  assign n39033 = ~n38667 | ~n38666;
  assign n38672 = ~n39033 | ~n38668;
  assign n38669 = ~P3_MORE_REG_SCAN_IN & ~P3_FLUSH_REG_SCAN_IN;
  assign n38671 = ~n38670 & ~n38669;
  assign n38685 = ~n38672 & ~n38671;
  assign n38676 = ~n38674 | ~n38673;
  assign n38680 = ~n38676 | ~n38675;
  assign n38679 = ~n38678 | ~n38677;
  assign n38684 = ~n38680 | ~n38679;
  assign n38683 = ~n38682 & ~n38681;
  assign n39100 = ~n38684 & ~n38683;
  assign n38787 = ~n38685 | ~n39100;
  assign n38722 = ~n38686 | ~n38781;
  assign n38690 = ~n38688 & ~n38687;
  assign n38691 = ~n38690 & ~n38689;
  assign n38693 = ~n38692 | ~n38691;
  assign n38698 = n38696 | n38695;
  assign n38697 = ~n38710;
  assign n38762 = n38698 & n38697;
  assign n38700 = ~n38762 & ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n38699 = ~n38763 & ~n23642;
  assign n38702 = ~n38700 & ~n38699;
  assign n38701 = ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN & ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign n38716 = ~n38702 & ~n38701;
  assign n38708 = ~n38704 | ~n38703;
  assign n38707 = ~n38706 | ~n38705;
  assign n38735 = ~n38708 | ~n38707;
  assign n38712 = ~n38732 & ~n38735;
  assign n38711 = ~n38710 | ~n38709;
  assign n38714 = n38712 & n38711;
  assign n38713 = ~n38723 | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign n38715 = ~n38714 & ~n38713;
  assign n38718 = ~n38716 & ~n38715;
  assign n38717 = ~n38730 | ~n39047;
  assign n39045 = ~n38718 | ~n38717;
  assign n38720 = ~n38788 | ~n38719;
  assign n38755 = ~n38721 | ~n38720;
  assign n38754 = ~n38722 | ~n38755;
  assign n38727 = ~n38724 | ~n38723;
  assign n38726 = ~n38725 | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n38729 = ~n38727 | ~n38726;
  assign n38731 = ~n38729 | ~n38728;
  assign n38734 = ~n38731 | ~n38730;
  assign n38733 = ~n38732 | ~n23643;
  assign n38739 = ~n38734 | ~n38733;
  assign n38737 = ~n38735;
  assign n38738 = ~n38737 & ~n38736;
  assign n38751 = ~n38739 & ~n38738;
  assign n38741 = ~n38740;
  assign n38749 = ~n38762 & ~n38741;
  assign n38743 = ~n38744 & ~n38741;
  assign n38747 = ~n38743 & ~n38742;
  assign n38746 = ~n38745 & ~n38744;
  assign n38748 = ~n38747 & ~n38746;
  assign n38750 = ~n38749 & ~n38748;
  assign n39037 = ~n38751 | ~n38750;
  assign n39030 = ~n38788;
  assign n38753 = ~n39037 | ~n39030;
  assign n38752 = ~n38788 | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign n38780 = ~n38753 | ~n38752;
  assign n38785 = ~n38754 | ~n38780;
  assign n38778 = ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN | ~n38755;
  assign n38774 = ~P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & ~n38755;
  assign n38765 = ~n38757 & ~n38756;
  assign n38760 = P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | n38765;
  assign n38759 = ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~n38758;
  assign n39072 = ~n38760 | ~n38759;
  assign n38771 = n39072 | n38761;
  assign n38764 = n38763 & n38762;
  assign n38767 = ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN & ~n38764;
  assign n38766 = ~n38765 & ~n39057;
  assign n39055 = ~n38767 & ~n38766;
  assign n38769 = ~n39072 | ~n38768;
  assign n38770 = ~n39055 | ~n38769;
  assign n38772 = ~n38771 | ~n38770;
  assign n38773 = ~n38788 & ~n38772;
  assign n38777 = ~n38776 | ~n38775;
  assign n38779 = ~n38778 | ~n38777;
  assign n38783 = ~P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN & ~n38779;
  assign n38782 = n38781 | n38780;
  assign n38784 = ~n38783 | ~n38782;
  assign n38786 = ~n38785 | ~n38784;
  assign n38789 = ~P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN | ~n38788;
  assign n38795 = ~n38790 | ~n38789;
  assign n38794 = ~n39105 | ~n38795;
  assign n38813 = n38804 & n39106;
  assign n38791 = ~n38811 & ~n39068;
  assign n38792 = ~n38813 & ~n38791;
  assign n38793 = ~n38792 | ~n39118;
  assign n38807 = ~n38794 | ~n38793;
  assign n38802 = ~n38795;
  assign n38798 = ~n38796;
  assign n38800 = ~n38798 & ~n38797;
  assign n38801 = ~n38800 & ~n38799;
  assign n39024 = ~n38802 | ~n38801;
  assign n38812 = ~n38804 | ~n38803;
  assign n38817 = ~n39024 | ~n38812;
  assign n38809 = ~n38807 & ~n38806;
  assign P3_U2996 = ~n38809 | ~n38808;
  assign n38822 = ~n38811 | ~n38810;
  assign n38826 = ~n38812 & ~n38822;
  assign n38821 = ~n38813 & ~n38826;
  assign n38816 = ~n38815 | ~n38814;
  assign n38819 = ~n38817 & ~n38816;
  assign n38820 = ~n38819 & ~n38818;
  assign P3_U2997 = ~n38821 | ~n38820;
  assign n38824 = ~n38823 | ~n38822;
  assign n38825 = ~n39026 | ~n38824;
  assign P3_U2998 = ~n38826 & ~n38825;
  assign P3_U2999 = P3_DATAWIDTH_REG_31__SCAN_IN & n22822;
  assign P3_U3000 = P3_DATAWIDTH_REG_30__SCAN_IN & n22822;
  assign P3_U3001 = P3_DATAWIDTH_REG_29__SCAN_IN & n22823;
  assign P3_U3002 = P3_DATAWIDTH_REG_28__SCAN_IN & n22823;
  assign P3_U3003 = P3_DATAWIDTH_REG_27__SCAN_IN & n22822;
  assign P3_U3004 = P3_DATAWIDTH_REG_26__SCAN_IN & n22822;
  assign P3_U3005 = P3_DATAWIDTH_REG_25__SCAN_IN & n22823;
  assign P3_U3006 = P3_DATAWIDTH_REG_24__SCAN_IN & n22822;
  assign P3_U3007 = P3_DATAWIDTH_REG_23__SCAN_IN & n22823;
  assign P3_U3008 = P3_DATAWIDTH_REG_22__SCAN_IN & n22822;
  assign P3_U3009 = P3_DATAWIDTH_REG_21__SCAN_IN & n22823;
  assign P3_U3010 = P3_DATAWIDTH_REG_20__SCAN_IN & n22822;
  assign P3_U3011 = P3_DATAWIDTH_REG_19__SCAN_IN & n22823;
  assign P3_U3012 = P3_DATAWIDTH_REG_18__SCAN_IN & n22822;
  assign P3_U3013 = P3_DATAWIDTH_REG_17__SCAN_IN & n22823;
  assign P3_U3014 = P3_DATAWIDTH_REG_16__SCAN_IN & n22822;
  assign P3_U3015 = P3_DATAWIDTH_REG_15__SCAN_IN & n22823;
  assign P3_U3016 = P3_DATAWIDTH_REG_14__SCAN_IN & n22822;
  assign P3_U3017 = P3_DATAWIDTH_REG_13__SCAN_IN & n22823;
  assign P3_U3018 = P3_DATAWIDTH_REG_12__SCAN_IN & n22822;
  assign P3_U3019 = P3_DATAWIDTH_REG_11__SCAN_IN & n22823;
  assign P3_U3020 = P3_DATAWIDTH_REG_10__SCAN_IN & n22822;
  assign P3_U3021 = P3_DATAWIDTH_REG_9__SCAN_IN & n22823;
  assign P3_U3022 = P3_DATAWIDTH_REG_8__SCAN_IN & n22823;
  assign P3_U3023 = P3_DATAWIDTH_REG_7__SCAN_IN & n22822;
  assign P3_U3024 = P3_DATAWIDTH_REG_6__SCAN_IN & n22823;
  assign P3_U3025 = P3_DATAWIDTH_REG_5__SCAN_IN & n22822;
  assign P3_U3026 = P3_DATAWIDTH_REG_4__SCAN_IN & n22823;
  assign P3_U3027 = P3_DATAWIDTH_REG_3__SCAN_IN & n22822;
  assign P3_U3028 = P3_DATAWIDTH_REG_2__SCAN_IN & n22823;
  assign n38850 = ~P3_STATE_REG_2__SCAN_IN | ~HOLD;
  assign n38836 = ~P3_REQUESTPENDING_REG_SCAN_IN | ~n38850;
  assign n38828 = ~n38831 & ~n41918;
  assign n38829 = ~n38836 & ~n38828;
  assign n38834 = n39126 | n38829;
  assign n44540 = ~NA;
  assign n38830 = ~P3_STATE_REG_1__SCAN_IN & ~n44540;
  assign n38848 = ~n38860 & ~n38830;
  assign n38832 = ~n38848;
  assign n38849 = ~n39114 & ~n38831;
  assign n38847 = n38854 | n38849;
  assign n38833 = ~n38832 | ~n38847;
  assign P3_U3029 = ~n38834 | ~n38833;
  assign n38835 = ~n39114 | ~P3_STATE_REG_2__SCAN_IN;
  assign n38846 = ~n38835 | ~n39126;
  assign n38837 = ~n38854 & ~n38836;
  assign n38842 = ~P3_STATE_REG_0__SCAN_IN & ~n38860;
  assign n38838 = ~n38837 & ~n38842;
  assign n38844 = ~P3_STATE_REG_1__SCAN_IN & ~n38838;
  assign n38856 = P3_REQUESTPENDING_REG_SCAN_IN | HOLD;
  assign n38839 = ~n38856 | ~n38850;
  assign n38840 = ~n38839 | ~n39114;
  assign n38841 = ~n38840 | ~P3_STATE_REG_1__SCAN_IN;
  assign n38843 = ~n38842 & ~n38841;
  assign n38845 = ~n38844 & ~n38843;
  assign P3_U3030 = ~n38846 | ~n38845;
  assign n38859 = ~n38848 | ~n38847;
  assign n38853 = ~P3_STATE_REG_1__SCAN_IN & ~P3_REQUESTPENDING_REG_SCAN_IN;
  assign n38851 = ~n38849 | ~n44540;
  assign n38852 = ~n38851 | ~n38850;
  assign n38855 = ~n38853 & ~n38852;
  assign n38857 = ~n38855 & ~n38854;
  assign n38858 = ~n38857 | ~n38856;
  assign P3_U3031 = ~n38859 | ~n38858;
  assign n38975 = ~n39126 | ~n38860;
  assign n38862 = ~n38865 & ~n38975;
  assign n38861 = ~n39005 & ~n39084;
  assign n38864 = ~n38862 & ~n38861;
  assign n38863 = ~P3_ADDRESS_REG_0__SCAN_IN | ~n39097;
  assign P3_U3032 = ~n38864 | ~n38863;
  assign n38867 = ~n38870 & ~n38975;
  assign n38866 = ~n39005 & ~n38865;
  assign n38869 = ~n38867 & ~n38866;
  assign n39125 = ~n39126;
  assign n38868 = ~P3_ADDRESS_REG_1__SCAN_IN | ~n39125;
  assign P3_U3033 = ~n38869 | ~n38868;
  assign n38872 = ~n38875 & ~n38975;
  assign n38871 = ~n39005 & ~n38870;
  assign n38874 = ~n38872 & ~n38871;
  assign n38873 = ~P3_ADDRESS_REG_2__SCAN_IN | ~n39125;
  assign P3_U3034 = ~n38874 | ~n38873;
  assign n38877 = ~n38880 & ~n38975;
  assign n38876 = ~n39005 & ~n38875;
  assign n38879 = ~n38877 & ~n38876;
  assign n38878 = ~P3_ADDRESS_REG_3__SCAN_IN | ~n39125;
  assign P3_U3035 = ~n38879 | ~n38878;
  assign n38885 = ~P3_REIP_REG_6__SCAN_IN;
  assign n38882 = ~n38885 & ~n38975;
  assign n38881 = ~n39005 & ~n38880;
  assign n38884 = ~n38882 & ~n38881;
  assign n38883 = ~P3_ADDRESS_REG_4__SCAN_IN | ~n39125;
  assign P3_U3036 = ~n38884 | ~n38883;
  assign n38887 = ~n38890 & ~n38975;
  assign n38886 = ~n39005 & ~n38885;
  assign n38889 = ~n38887 & ~n38886;
  assign n38888 = ~P3_ADDRESS_REG_5__SCAN_IN | ~n39125;
  assign P3_U3037 = ~n38889 | ~n38888;
  assign n38895 = ~P3_REIP_REG_8__SCAN_IN;
  assign n38892 = ~n38895 & ~n38975;
  assign n38891 = ~n39005 & ~n38890;
  assign n38894 = ~n38892 & ~n38891;
  assign n38893 = ~P3_ADDRESS_REG_6__SCAN_IN | ~n39125;
  assign P3_U3038 = ~n38894 | ~n38893;
  assign n38897 = ~n38900 & ~n38975;
  assign n38896 = ~n39005 & ~n38895;
  assign n38899 = ~n38897 & ~n38896;
  assign n38898 = ~P3_ADDRESS_REG_7__SCAN_IN | ~n39125;
  assign P3_U3039 = ~n38899 | ~n38898;
  assign n38902 = ~n38905 & ~n38975;
  assign n38901 = ~n39005 & ~n38900;
  assign n38904 = ~n38902 & ~n38901;
  assign n38903 = ~P3_ADDRESS_REG_8__SCAN_IN | ~n39125;
  assign P3_U3040 = ~n38904 | ~n38903;
  assign n38907 = ~n38910 & ~n38975;
  assign n38906 = ~n39005 & ~n38905;
  assign n38909 = ~n38907 & ~n38906;
  assign n38908 = ~P3_ADDRESS_REG_9__SCAN_IN | ~n39125;
  assign P3_U3041 = ~n38909 | ~n38908;
  assign n38912 = ~n38915 & ~n38975;
  assign n38911 = ~n39005 & ~n38910;
  assign n38914 = ~n38912 & ~n38911;
  assign n38913 = ~P3_ADDRESS_REG_10__SCAN_IN | ~n39125;
  assign P3_U3042 = ~n38914 | ~n38913;
  assign n38917 = ~n38920 & ~n38975;
  assign n38916 = ~n39005 & ~n38915;
  assign n38919 = ~n38917 & ~n38916;
  assign n38918 = ~P3_ADDRESS_REG_11__SCAN_IN | ~n39125;
  assign P3_U3043 = ~n38919 | ~n38918;
  assign n38922 = ~n38925 & ~n38975;
  assign n38921 = ~n39005 & ~n38920;
  assign n38924 = ~n38922 & ~n38921;
  assign n38923 = ~P3_ADDRESS_REG_12__SCAN_IN | ~n39125;
  assign P3_U3044 = ~n38924 | ~n38923;
  assign n38927 = ~n38930 & ~n38975;
  assign n38926 = ~n39005 & ~n38925;
  assign n38929 = ~n38927 & ~n38926;
  assign n38928 = ~P3_ADDRESS_REG_13__SCAN_IN | ~n39125;
  assign P3_U3045 = ~n38929 | ~n38928;
  assign n38935 = ~P3_REIP_REG_16__SCAN_IN;
  assign n38932 = ~n38935 & ~n38975;
  assign n38931 = ~n39005 & ~n38930;
  assign n38934 = ~n38932 & ~n38931;
  assign n38933 = ~P3_ADDRESS_REG_14__SCAN_IN | ~n39125;
  assign P3_U3046 = ~n38934 | ~n38933;
  assign n38937 = ~n38940 & ~n38975;
  assign n38936 = ~n39005 & ~n38935;
  assign n38939 = ~n38937 & ~n38936;
  assign n38938 = ~P3_ADDRESS_REG_15__SCAN_IN | ~n39125;
  assign P3_U3047 = ~n38939 | ~n38938;
  assign n38945 = ~P3_REIP_REG_18__SCAN_IN;
  assign n38942 = ~n38945 & ~n38975;
  assign n38941 = ~n39005 & ~n38940;
  assign n38944 = ~n38942 & ~n38941;
  assign n38943 = ~P3_ADDRESS_REG_16__SCAN_IN | ~n39125;
  assign P3_U3048 = ~n38944 | ~n38943;
  assign n38947 = ~n38950 & ~n38975;
  assign n38946 = ~n39005 & ~n38945;
  assign n38949 = ~n38947 & ~n38946;
  assign n38948 = ~P3_ADDRESS_REG_17__SCAN_IN | ~n39125;
  assign P3_U3049 = ~n38949 | ~n38948;
  assign n38955 = ~P3_REIP_REG_20__SCAN_IN;
  assign n38952 = ~n38955 & ~n38975;
  assign n38951 = ~n39005 & ~n38950;
  assign n38954 = ~n38952 & ~n38951;
  assign n38953 = ~P3_ADDRESS_REG_18__SCAN_IN | ~n39125;
  assign P3_U3050 = ~n38954 | ~n38953;
  assign n38957 = ~n38960 & ~n38975;
  assign n38956 = ~n39005 & ~n38955;
  assign n38959 = ~n38957 & ~n38956;
  assign n38958 = ~P3_ADDRESS_REG_19__SCAN_IN | ~n39125;
  assign P3_U3051 = ~n38959 | ~n38958;
  assign n38962 = ~n38965 & ~n38975;
  assign n38961 = ~n39005 & ~n38960;
  assign n38964 = ~n38962 & ~n38961;
  assign n38963 = ~P3_ADDRESS_REG_20__SCAN_IN | ~n39125;
  assign P3_U3052 = ~n38964 | ~n38963;
  assign n38967 = ~n38970 & ~n38975;
  assign n38966 = ~n39005 & ~n38965;
  assign n38969 = ~n38967 & ~n38966;
  assign n38968 = ~P3_ADDRESS_REG_21__SCAN_IN | ~n39097;
  assign P3_U3053 = ~n38969 | ~n38968;
  assign n38976 = ~P3_REIP_REG_24__SCAN_IN;
  assign n38972 = ~n38976 & ~n38975;
  assign n38971 = ~n39005 & ~n38970;
  assign n38974 = ~n38972 & ~n38971;
  assign n38973 = ~P3_ADDRESS_REG_22__SCAN_IN | ~n39097;
  assign P3_U3054 = ~n38974 | ~n38973;
  assign n38978 = ~n38981 & ~n38975;
  assign n38977 = ~n39005 & ~n38976;
  assign n38980 = ~n38978 & ~n38977;
  assign n38979 = ~P3_ADDRESS_REG_23__SCAN_IN | ~n39097;
  assign P3_U3055 = ~n38980 | ~n38979;
  assign n38986 = ~P3_REIP_REG_26__SCAN_IN;
  assign n38983 = ~n38986 & ~n38975;
  assign n38982 = ~n39005 & ~n38981;
  assign n38985 = ~n38983 & ~n38982;
  assign n38984 = ~P3_ADDRESS_REG_24__SCAN_IN | ~n39097;
  assign P3_U3056 = ~n38985 | ~n38984;
  assign n38991 = ~P3_REIP_REG_27__SCAN_IN;
  assign n38988 = ~n38991 & ~n38975;
  assign n38987 = ~n39005 & ~n38986;
  assign n38990 = ~n38988 & ~n38987;
  assign n38989 = ~P3_ADDRESS_REG_25__SCAN_IN | ~n39097;
  assign P3_U3057 = ~n38990 | ~n38989;
  assign n38993 = ~n33447 & ~n38975;
  assign n38992 = ~n39005 & ~n38991;
  assign n38995 = ~n38993 & ~n38992;
  assign n38994 = ~P3_ADDRESS_REG_26__SCAN_IN | ~n39097;
  assign P3_U3058 = ~n38995 | ~n38994;
  assign n38997 = ~n33351 & ~n38975;
  assign n38996 = ~n39005 & ~n33447;
  assign n38999 = ~n38997 & ~n38996;
  assign n38998 = ~P3_ADDRESS_REG_27__SCAN_IN | ~n39097;
  assign P3_U3059 = ~n38999 | ~n38998;
  assign n39004 = ~P3_REIP_REG_30__SCAN_IN;
  assign n39001 = ~n39004 & ~n38975;
  assign n39000 = ~n39005 & ~n33351;
  assign n39003 = ~n39001 & ~n39000;
  assign n39002 = ~P3_ADDRESS_REG_28__SCAN_IN | ~n39097;
  assign P3_U3060 = ~n39003 | ~n39002;
  assign n39008 = ~n39005 & ~n39004;
  assign n39007 = ~n39006 & ~n38975;
  assign n39010 = ~n39008 & ~n39007;
  assign n39009 = ~P3_ADDRESS_REG_29__SCAN_IN | ~n39097;
  assign P3_U3061 = ~n39010 | ~n39009;
  assign n39012 = ~n39125 | ~P3_BE_N_REG_3__SCAN_IN;
  assign n39011 = ~n39126 | ~P3_BYTEENABLE_REG_3__SCAN_IN;
  assign P3_U3274 = ~n39012 | ~n39011;
  assign n39014 = ~n39125 | ~P3_BE_N_REG_2__SCAN_IN;
  assign n39013 = ~n39126 | ~P3_BYTEENABLE_REG_2__SCAN_IN;
  assign P3_U3275 = ~n39014 | ~n39013;
  assign n39016 = ~n39097 | ~P3_BE_N_REG_1__SCAN_IN;
  assign n39015 = ~n39126 | ~P3_BYTEENABLE_REG_1__SCAN_IN;
  assign P3_U3276 = ~n39016 | ~n39015;
  assign n39018 = ~n39125 | ~P3_BE_N_REG_0__SCAN_IN;
  assign n39017 = ~n39126 | ~P3_BYTEENABLE_REG_0__SCAN_IN;
  assign P3_U3277 = ~n39018 | ~n39017;
  assign n39021 = ~n39023;
  assign n39020 = ~P3_DATAWIDTH_REG_0__SCAN_IN & ~n39019;
  assign P3_U3280 = ~n39021 & ~n39020;
  assign n39022 = ~P3_DATAWIDTH_REG_1__SCAN_IN | ~n22823;
  assign P3_U3281 = ~n39023 | ~n39022;
  assign n39025 = ~n39024 | ~P3_STATE2_REG_0__SCAN_IN;
  assign n39027 = ~n39025 | ~P3_STATE2_REG_3__SCAN_IN;
  assign P3_U3282 = ~n39027 | ~n39026;
  assign n39032 = ~n39029 & ~n39028;
  assign n39031 = ~n39105 | ~n39030;
  assign n39034 = ~n39078 & ~n39033;
  assign n39036 = ~n39034 | ~n39073;
  assign n39035 = ~n39078 | ~P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN;
  assign P3_U3284 = ~n39036 | ~n39035;
  assign n39041 = ~n39073 | ~n39037;
  assign n39040 = ~n39039 | ~n39038;
  assign n39042 = ~n39041 | ~n39040;
  assign n39044 = ~n39077 | ~n39042;
  assign n39043 = ~n39078 | ~P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign P3_U3285 = ~n39044 | ~n39043;
  assign n39051 = ~n39073 | ~n39045;
  assign n39061 = n39046 ^ P3_INSTADDRPOINTER_REG_1__SCAN_IN;
  assign n39060 = ~P3_INSTADDRPOINTER_REG_0__SCAN_IN | ~P3_STATE2_REG_1__SCAN_IN;
  assign n39049 = ~n39061 & ~n39060;
  assign n39048 = ~n39047 & ~n39068;
  assign n39050 = ~n39049 & ~n39048;
  assign n39052 = ~n39051 | ~n39050;
  assign n39054 = ~n39077 | ~n39052;
  assign n39053 = ~n39078 | ~P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign P3_U3288 = ~n39054 | ~n39053;
  assign n39059 = ~n39056 & ~n39055;
  assign n39058 = ~n39057 & ~n39068;
  assign n39064 = ~n39059 & ~n39058;
  assign n39062 = ~n39060;
  assign n39063 = ~n39062 | ~n39061;
  assign n39065 = ~n39064 | ~n39063;
  assign n39067 = ~n39077 | ~n39065;
  assign n39066 = ~n39078 | ~P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign P3_U3289 = ~n39067 | ~n39066;
  assign n39071 = ~n39068 & ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN;
  assign n39070 = ~n39069 & ~P3_INSTADDRPOINTER_REG_0__SCAN_IN;
  assign n39075 = ~n39071 & ~n39070;
  assign n39074 = ~n39073 | ~n39072;
  assign n39076 = ~n39075 | ~n39074;
  assign n39080 = ~n39077 | ~n39076;
  assign n39079 = ~P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~n39078;
  assign P3_U3290 = ~n39080 | ~n39079;
  assign n39091 = ~n39092 | ~P3_BYTEENABLE_REG_2__SCAN_IN;
  assign n39088 = ~n39081 | ~n39082;
  assign n39093 = ~n39084 | ~n39083;
  assign n39086 = ~n39082 & ~n39093;
  assign n39085 = ~n39084 & ~n39083;
  assign n39087 = ~n39086 & ~n39085;
  assign n39089 = ~n39088 | ~n39087;
  assign n39094 = ~n39092;
  assign n39090 = ~n39089 | ~n39094;
  assign P3_U3292 = ~n39091 | ~n39090;
  assign n39096 = ~n39092 | ~P3_BYTEENABLE_REG_0__SCAN_IN;
  assign n39095 = ~n39094 | ~n39093;
  assign P3_U3293 = ~n39096 | ~n39095;
  assign n39099 = ~P3_W_R_N_REG_SCAN_IN | ~n39097;
  assign n39098 = n39125 | P3_READREQUEST_REG_SCAN_IN;
  assign P3_U3294 = ~n39099 | ~n39098;
  assign n39103 = ~P3_MORE_REG_SCAN_IN | ~n39101;
  assign n39102 = n39101 | n39100;
  assign P3_U3295 = ~n39103 | ~n39102;
  assign n39109 = ~n39105 & ~n39104;
  assign n39107 = ~n39106 | ~n39114;
  assign n39108 = ~n39107 | ~n39132;
  assign n39122 = ~n39109 & ~n39108;
  assign n39124 = ~P3_REQUESTPENDING_REG_SCAN_IN | ~n39122;
  assign n39111 = ~n39110 & ~P3_STATEBS16_REG_SCAN_IN;
  assign n39113 = ~n39112 & ~n39111;
  assign n39116 = ~n39129 & ~n39113;
  assign n39115 = ~P3_STATE2_REG_2__SCAN_IN | ~n39114;
  assign n39117 = ~n39116 & ~n39115;
  assign n39119 = ~n39118 & ~n39117;
  assign n39121 = ~n39120 & ~n39119;
  assign n39123 = n39122 | n39121;
  assign P3_U3296 = ~n39124 | ~n39123;
  assign n39128 = ~n39125 | ~P3_M_IO_N_REG_SCAN_IN;
  assign n39127 = ~n39126 | ~P3_MEMORYFETCH_REG_SCAN_IN;
  assign P3_U3297 = ~n39128 | ~n39127;
  assign n39134 = ~n39132 & ~n39129;
  assign n39131 = ~n39130;
  assign n39135 = ~n39132 | ~n39131;
  assign n39133 = ~n39135 & ~P3_READREQUEST_REG_SCAN_IN;
  assign P3_U3298 = ~n39134 & ~n39133;
  assign n39137 = ~n39135 & ~P3_MEMORYFETCH_REG_SCAN_IN;
  assign P3_U3299 = ~n39137 & ~n39136;
  assign n39139 = ~n39138;
  assign n39142 = ~n39140;
  assign n39143 = ~n39142 | ~n39141;
  assign n39144 = ~n39143 | ~P2_MEMORYFETCH_REG_SCAN_IN;
  assign n39146 = n40117 & n39144;
  assign n39145 = ~n39150;
  assign P2_U2814 = ~n39146 | ~n39145;
  assign n39147 = ~P2_STATE_REG_2__SCAN_IN & ~n41920;
  assign n39148 = ~P2_STATE_REG_1__SCAN_IN | ~n39147;
  assign n41897 = ~n41920 | ~n39153;
  assign n42070 = ~n39148 | ~n41897;
  assign n39149 = ~P2_STATE_REG_0__SCAN_IN | ~P2_ADS_N_REG_SCAN_IN;
  assign P2_U2815 = ~n22819 | ~n39149;
  assign n39152 = ~P2_STATE2_REG_0__SCAN_IN | ~n39150;
  assign n39151 = ~P2_CODEFETCH_REG_SCAN_IN | ~n42200;
  assign P2_U2816 = ~n39152 | ~n39151;
  assign n42224 = ~n42065;
  assign n42223 = ~n42224;
  assign n39155 = ~P2_CODEFETCH_REG_SCAN_IN & ~n42223;
  assign n41911 = ~n39153 | ~n41926;
  assign n39154 = ~P2_STATE_REG_0__SCAN_IN & ~n41911;
  assign n39157 = ~n39155 & ~n39154;
  assign n39156 = ~P2_D_C_N_REG_SCAN_IN | ~n42223;
  assign P2_U2817 = ~n39157 | ~n39156;
  assign n42245 = ~BS16;
  assign n39158 = ~n41911 | ~n42245;
  assign n42074 = ~n42070 | ~n39158;
  assign n39159 = ~P2_STATEBS16_REG_SCAN_IN | ~n22820;
  assign P2_U2818 = ~n42074 | ~n39159;
  assign n42193 = n39161 & n39160;
  assign n42191 = ~n42193;
  assign n39162 = ~P2_FLUSH_REG_SCAN_IN | ~n42191;
  assign P2_U2819 = ~n39163 | ~n39162;
  assign n39165 = ~P2_DATAWIDTH_REG_4__SCAN_IN & ~P2_DATAWIDTH_REG_5__SCAN_IN;
  assign n39164 = ~P2_DATAWIDTH_REG_6__SCAN_IN & ~P2_DATAWIDTH_REG_7__SCAN_IN;
  assign n39169 = ~n39165 | ~n39164;
  assign n39167 = ~P2_DATAWIDTH_REG_3__SCAN_IN & ~P2_DATAWIDTH_REG_2__SCAN_IN;
  assign n39166 = ~P2_DATAWIDTH_REG_0__SCAN_IN | ~P2_DATAWIDTH_REG_1__SCAN_IN;
  assign n39168 = ~n39167 | ~n39166;
  assign n39193 = ~n39169 & ~n39168;
  assign n39171 = ~P2_DATAWIDTH_REG_12__SCAN_IN & ~P2_DATAWIDTH_REG_13__SCAN_IN;
  assign n39170 = ~P2_DATAWIDTH_REG_14__SCAN_IN & ~P2_DATAWIDTH_REG_15__SCAN_IN;
  assign n39175 = ~n39171 | ~n39170;
  assign n39173 = ~P2_DATAWIDTH_REG_8__SCAN_IN & ~P2_DATAWIDTH_REG_9__SCAN_IN;
  assign n39172 = ~P2_DATAWIDTH_REG_10__SCAN_IN & ~P2_DATAWIDTH_REG_11__SCAN_IN;
  assign n39174 = ~n39173 | ~n39172;
  assign n39191 = n39175 | n39174;
  assign n39177 = ~P2_DATAWIDTH_REG_20__SCAN_IN & ~P2_DATAWIDTH_REG_21__SCAN_IN;
  assign n39176 = ~P2_DATAWIDTH_REG_22__SCAN_IN & ~P2_DATAWIDTH_REG_23__SCAN_IN;
  assign n39181 = ~n39177 | ~n39176;
  assign n39179 = ~P2_DATAWIDTH_REG_16__SCAN_IN & ~P2_DATAWIDTH_REG_17__SCAN_IN;
  assign n39178 = ~P2_DATAWIDTH_REG_18__SCAN_IN & ~P2_DATAWIDTH_REG_19__SCAN_IN;
  assign n39180 = ~n39179 | ~n39178;
  assign n39189 = ~n39181 & ~n39180;
  assign n39183 = ~P2_DATAWIDTH_REG_28__SCAN_IN & ~P2_DATAWIDTH_REG_29__SCAN_IN;
  assign n39182 = ~P2_DATAWIDTH_REG_30__SCAN_IN & ~P2_DATAWIDTH_REG_31__SCAN_IN;
  assign n39187 = ~n39183 | ~n39182;
  assign n39185 = ~P2_DATAWIDTH_REG_24__SCAN_IN & ~P2_DATAWIDTH_REG_25__SCAN_IN;
  assign n39184 = ~P2_DATAWIDTH_REG_26__SCAN_IN & ~P2_DATAWIDTH_REG_27__SCAN_IN;
  assign n39186 = ~n39185 | ~n39184;
  assign n39188 = ~n39187 & ~n39186;
  assign n39190 = ~n39189 | ~n39188;
  assign n39192 = ~n39191 & ~n39190;
  assign n39210 = ~n39193 | ~n39192;
  assign n39207 = ~n39210;
  assign n39195 = ~n39207 & ~P2_BYTEENABLE_REG_0__SCAN_IN;
  assign n39200 = ~n27692 | ~n39207;
  assign n39194 = ~P2_REIP_REG_0__SCAN_IN & ~n39200;
  assign P2_U2820 = ~n39195 & ~n39194;
  assign n39198 = ~n39207 & ~P2_BYTEENABLE_REG_1__SCAN_IN;
  assign n39196 = P2_DATAWIDTH_REG_1__SCAN_IN | P2_DATAWIDTH_REG_0__SCAN_IN;
  assign n39206 = ~P2_REIP_REG_0__SCAN_IN & ~n39196;
  assign n39197 = ~n39200 & ~n39206;
  assign P2_U2821 = ~n39198 & ~n39197;
  assign n39199 = ~P2_REIP_REG_1__SCAN_IN | ~P2_REIP_REG_0__SCAN_IN;
  assign n39203 = ~n39199 & ~n39210;
  assign n39208 = n39200 | P2_DATAWIDTH_REG_1__SCAN_IN;
  assign n39201 = P2_REIP_REG_0__SCAN_IN & P2_DATAWIDTH_REG_0__SCAN_IN;
  assign n39202 = ~n39208 & ~n39201;
  assign n39205 = ~n39203 & ~n39202;
  assign n39204 = ~P2_BYTEENABLE_REG_2__SCAN_IN | ~n39210;
  assign P2_U2822 = ~n39205 | ~n39204;
  assign n39209 = ~n39207 | ~n39206;
  assign n39212 = n39209 & n39208;
  assign n39211 = ~n39210 | ~P2_BYTEENABLE_REG_3__SCAN_IN;
  assign P2_U2823 = ~n39212 | ~n39211;
  assign n39213 = ~P2_EBX_REG_22__SCAN_IN;
  assign n39223 = ~n39214 | ~n39639;
  assign n39221 = ~n32310 & ~n39516;
  assign n39216 = ~n42097 & ~n39215;
  assign n39218 = ~P2_PHYADDRPOINTER_REG_22__SCAN_IN | ~n39672;
  assign n39220 = ~n39219 | ~n39218;
  assign n39222 = ~n39221 & ~n39220;
  assign n39227 = ~n39224 & ~n39628;
  assign n39226 = ~n39225 & ~n39683;
  assign n39228 = ~n39227 & ~n39226;
  assign n39229 = ~P2_EBX_REG_21__SCAN_IN;
  assign n39241 = ~n39229 & ~n39495;
  assign n39239 = ~n39230 | ~n39639;
  assign n39237 = ~n28457 & ~n39516;
  assign n39232 = ~n42095 | ~n39261;
  assign n39233 = ~n39232 ^ n39231;
  assign n39235 = ~n39233 | ~n39647;
  assign n39234 = ~P2_PHYADDRPOINTER_REG_21__SCAN_IN | ~n39672;
  assign n39236 = ~n39235 | ~n39234;
  assign n39238 = ~n39237 & ~n39236;
  assign n39240 = ~n39239 | ~n39238;
  assign n39247 = ~n39241 & ~n39240;
  assign n39245 = ~n39242 & ~n39628;
  assign n39244 = ~n39243 & ~n39683;
  assign n39246 = ~n39245 & ~n39244;
  assign P2_U2834 = ~n39247 | ~n39246;
  assign n39266 = n39248 & n39686;
  assign n39673 = ~n42095 & ~n41893;
  assign n39252 = ~n39258 & ~n39335;
  assign n39250 = ~n39672 | ~P2_PHYADDRPOINTER_REG_20__SCAN_IN;
  assign n39249 = ~n39678 | ~P2_EBX_REG_20__SCAN_IN;
  assign n39251 = ~n39250 | ~n39249;
  assign n39254 = ~n39252 & ~n39251;
  assign n39253 = ~n39677 | ~P2_REIP_REG_20__SCAN_IN;
  assign n39257 = ~n39254 | ~n39253;
  assign n39256 = ~n39255 & ~n39683;
  assign n39264 = ~n39257 & ~n39256;
  assign n39260 = ~n39259 & ~n39258;
  assign n39262 = ~n39653 & ~n39260;
  assign n39263 = ~n39262 | ~n39261;
  assign n39265 = ~n39264 | ~n39263;
  assign n39269 = ~n39266 & ~n39265;
  assign n39268 = ~n39267 | ~n39639;
  assign P2_U2835 = ~n39269 | ~n39268;
  assign n39279 = ~n39270 & ~n39628;
  assign n39273 = ~n42095 | ~n39271;
  assign n39274 = ~n39273 ^ n39272;
  assign n39277 = ~n39274 | ~n39647;
  assign n39276 = ~n39275 | ~n39639;
  assign n39278 = ~n39277 | ~n39276;
  assign n39289 = ~n39279 & ~n39278;
  assign n39287 = ~n39280 & ~n39683;
  assign n39282 = ~n39672 | ~P2_PHYADDRPOINTER_REG_19__SCAN_IN;
  assign n39281 = ~n39678 | ~P2_EBX_REG_19__SCAN_IN;
  assign n39283 = ~n39282 | ~n39281;
  assign n39285 = ~n40325 & ~n39283;
  assign n39284 = ~n39677 | ~P2_REIP_REG_19__SCAN_IN;
  assign n39286 = ~n39285 | ~n39284;
  assign n39288 = ~n39287 & ~n39286;
  assign P2_U2836 = ~n39289 | ~n39288;
  assign n39307 = ~n39290 & ~n39628;
  assign n39292 = ~n39291 ^ n39297;
  assign n39303 = ~n39653 & ~n39292;
  assign n39294 = ~n39677 | ~P2_REIP_REG_18__SCAN_IN;
  assign n39293 = ~n39672 | ~P2_PHYADDRPOINTER_REG_18__SCAN_IN;
  assign n39295 = ~n39294 | ~n39293;
  assign n39301 = ~n40325 & ~n39295;
  assign n39299 = ~n39296 & ~n39683;
  assign n39298 = ~n39297 & ~n39335;
  assign n39300 = ~n39299 & ~n39298;
  assign n39302 = ~n39301 | ~n39300;
  assign n39305 = ~n39303 & ~n39302;
  assign n39304 = ~n39678 | ~P2_EBX_REG_18__SCAN_IN;
  assign n39306 = ~n39305 | ~n39304;
  assign n39310 = ~n39307 & ~n39306;
  assign n39309 = ~n39308 | ~n39639;
  assign P2_U2837 = ~n39310 | ~n39309;
  assign n39312 = ~n39677 | ~P2_REIP_REG_17__SCAN_IN;
  assign n39311 = ~n39672 | ~P2_PHYADDRPOINTER_REG_17__SCAN_IN;
  assign n39323 = ~n39312 | ~n39311;
  assign n39316 = ~n39313 & ~n39683;
  assign n39314 = ~P2_EBX_REG_17__SCAN_IN;
  assign n39315 = ~n39495 & ~n39314;
  assign n39321 = ~n39316 & ~n39315;
  assign n39318 = ~n39324 ^ n39317;
  assign n39319 = ~n39653 & ~n39318;
  assign n39320 = ~n39319 & ~n40325;
  assign n39322 = ~n39321 | ~n39320;
  assign n39332 = ~n39323 & ~n39322;
  assign n39327 = ~n39673 | ~n39324;
  assign n39326 = ~n39325 | ~n39639;
  assign n39330 = ~n39327 | ~n39326;
  assign n39329 = ~n39328 & ~n39628;
  assign n39331 = ~n39330 & ~n39329;
  assign P2_U2838 = ~n39332 | ~n39331;
  assign n39334 = ~n39333 ^ n39336;
  assign n39350 = ~n39653 & ~n39334;
  assign n39346 = ~n39336 & ~n39335;
  assign n39338 = ~n39677 | ~P2_REIP_REG_16__SCAN_IN;
  assign n39337 = ~n39672 | ~P2_PHYADDRPOINTER_REG_16__SCAN_IN;
  assign n39339 = ~n39338 | ~n39337;
  assign n39344 = ~n40325 & ~n39339;
  assign n39342 = ~n39340 & ~n39683;
  assign n39697 = ~P2_EBX_REG_16__SCAN_IN;
  assign n39341 = ~n39495 & ~n39697;
  assign n39343 = ~n39342 & ~n39341;
  assign n39345 = ~n39344 | ~n39343;
  assign n39348 = ~n39346 & ~n39345;
  assign n39347 = ~n39704 | ~n39639;
  assign n39349 = ~n39348 | ~n39347;
  assign n39353 = ~n39350 & ~n39349;
  assign n39829 = ~n39351;
  assign n39352 = ~n39829 | ~n39686;
  assign P2_U2839 = ~n39353 | ~n39352;
  assign n39355 = ~n39677 | ~P2_REIP_REG_15__SCAN_IN;
  assign n39354 = ~n39672 | ~P2_PHYADDRPOINTER_REG_15__SCAN_IN;
  assign n39366 = ~n39355 | ~n39354;
  assign n39357 = ~n39356;
  assign n39359 = ~n39357 & ~n39683;
  assign n39707 = ~P2_EBX_REG_15__SCAN_IN;
  assign n39358 = ~n39495 & ~n39707;
  assign n39364 = ~n39359 & ~n39358;
  assign n39361 = ~n39367 ^ n39360;
  assign n39362 = ~n39653 & ~n39361;
  assign n39363 = ~n39362 & ~n40325;
  assign n39365 = ~n39364 | ~n39363;
  assign n39373 = ~n39366 & ~n39365;
  assign n39369 = ~n39673 | ~n39367;
  assign n39368 = ~n39713 | ~n39639;
  assign n39371 = ~n39369 | ~n39368;
  assign n39370 = ~n39846 & ~n39628;
  assign n39372 = ~n39371 & ~n39370;
  assign P2_U2840 = ~n39373 | ~n39372;
  assign n39375 = ~n39677 | ~P2_REIP_REG_14__SCAN_IN;
  assign n39374 = ~n39656 | ~P2_PHYADDRPOINTER_REG_14__SCAN_IN;
  assign n39386 = ~n39375 | ~n39374;
  assign n39378 = ~n39376 & ~n39683;
  assign n39716 = ~P2_EBX_REG_14__SCAN_IN;
  assign n39377 = ~n39495 & ~n39716;
  assign n39384 = ~n39378 & ~n39377;
  assign n39387 = ~n39379;
  assign n39381 = n39380 ^ n39387;
  assign n39382 = ~n39653 & ~n39381;
  assign n39383 = ~n39382 & ~n40325;
  assign n39385 = ~n39384 | ~n39383;
  assign n39393 = ~n39386 & ~n39385;
  assign n39389 = ~n39673 | ~n39387;
  assign n39388 = ~n39721 | ~n39639;
  assign n39391 = ~n39389 | ~n39388;
  assign n39390 = ~n39855 & ~n39628;
  assign n39392 = ~n39391 & ~n39390;
  assign P2_U2841 = ~n39393 | ~n39392;
  assign n39395 = ~n39396 ^ n39394;
  assign n39411 = ~n39653 & ~n39395;
  assign n39401 = ~n39396 | ~n39673;
  assign n39398 = ~n39677 | ~P2_REIP_REG_13__SCAN_IN;
  assign n39397 = ~n39656 | ~P2_PHYADDRPOINTER_REG_13__SCAN_IN;
  assign n39399 = ~n39398 | ~n39397;
  assign n39400 = ~n40325 & ~n39399;
  assign n39404 = ~n39401 | ~n39400;
  assign n39403 = ~n39402 & ~n39683;
  assign n39409 = ~n39404 & ~n39403;
  assign n39724 = ~P2_EBX_REG_13__SCAN_IN;
  assign n39407 = ~n39495 & ~n39724;
  assign n39860 = ~n39405;
  assign n39406 = ~n39860 & ~n39628;
  assign n39408 = ~n39407 & ~n39406;
  assign n39410 = ~n39409 | ~n39408;
  assign n39413 = ~n39411 & ~n39410;
  assign n39412 = ~n39732 | ~n39639;
  assign P2_U2842 = ~n39413 | ~n39412;
  assign n39415 = ~n39677 | ~P2_REIP_REG_12__SCAN_IN;
  assign n39414 = ~n39656 | ~P2_PHYADDRPOINTER_REG_12__SCAN_IN;
  assign n39425 = ~n39415 | ~n39414;
  assign n39418 = n39416 | n39683;
  assign n39417 = ~n39678 | ~P2_EBX_REG_12__SCAN_IN;
  assign n39423 = n39418 & n39417;
  assign n39426 = ~n39419;
  assign n39420 = n39443 ^ n39426;
  assign n39421 = ~n39653 & ~n39420;
  assign n39422 = ~n39421 & ~n40325;
  assign n39424 = ~n39423 | ~n39422;
  assign n39433 = ~n39425 & ~n39424;
  assign n39428 = ~n39673 | ~n39426;
  assign n39427 = ~n39741 | ~n39639;
  assign n39431 = ~n39428 | ~n39427;
  assign n39865 = ~n39429;
  assign n39430 = ~n39865 & ~n39628;
  assign n39432 = ~n39431 & ~n39430;
  assign P2_U2843 = ~n39433 | ~n39432;
  assign n39435 = ~n39677 | ~P2_REIP_REG_11__SCAN_IN;
  assign n39434 = ~n39656 | ~P2_PHYADDRPOINTER_REG_11__SCAN_IN;
  assign n39436 = ~n39435 | ~n39434;
  assign n39438 = ~n40325 & ~n39436;
  assign n39437 = ~P2_EBX_REG_11__SCAN_IN | ~n39678;
  assign n39442 = ~n39438 | ~n39437;
  assign n39440 = ~n39439;
  assign n39441 = ~n39440 & ~n39683;
  assign n39448 = ~n39442 & ~n39441;
  assign n39446 = ~n39443 & ~n39653;
  assign n39445 = ~n39453 | ~n39444;
  assign n39447 = ~n39446 | ~n39445;
  assign n39452 = ~n39448 | ~n39447;
  assign n39450 = ~n39870 | ~n39686;
  assign n39449 = ~n39751 | ~n39639;
  assign n39451 = ~n39450 | ~n39449;
  assign n39455 = ~n39452 & ~n39451;
  assign n39454 = ~n39453 | ~n39673;
  assign P2_U2844 = ~n39455 | ~n39454;
  assign n39457 = ~n39677 | ~P2_REIP_REG_10__SCAN_IN;
  assign n39456 = ~n39656 | ~P2_PHYADDRPOINTER_REG_10__SCAN_IN;
  assign n39468 = ~n39457 | ~n39456;
  assign n39460 = ~n39458 & ~n39683;
  assign n39754 = ~P2_EBX_REG_10__SCAN_IN;
  assign n39459 = ~n39495 & ~n39754;
  assign n39466 = ~n39460 & ~n39459;
  assign n39469 = ~n39461;
  assign n39463 = n39462 ^ n39469;
  assign n39464 = ~n39653 & ~n39463;
  assign n39465 = ~n39464 & ~n40325;
  assign n39467 = ~n39466 | ~n39465;
  assign n39475 = ~n39468 & ~n39467;
  assign n39471 = ~n39673 | ~n39469;
  assign n39470 = ~n39759 | ~n39639;
  assign n39473 = ~n39471 | ~n39470;
  assign n39472 = ~n39876 & ~n39628;
  assign n39474 = ~n39473 & ~n39472;
  assign P2_U2845 = ~n39475 | ~n39474;
  assign n39477 = ~n39677 | ~P2_REIP_REG_9__SCAN_IN;
  assign n39476 = ~n39656 | ~P2_PHYADDRPOINTER_REG_9__SCAN_IN;
  assign n39478 = ~n39477 | ~n39476;
  assign n39483 = ~n40325 & ~n39478;
  assign n39481 = ~n39881 | ~n39686;
  assign n39480 = ~n39479 | ~n39520;
  assign n39482 = n39481 & n39480;
  assign n39491 = ~n39483 | ~n39482;
  assign n39486 = ~n42095 | ~n39484;
  assign n39487 = ~n39486 ^ n39485;
  assign n39489 = ~n39487 | ~n39647;
  assign n39488 = ~P2_EBX_REG_9__SCAN_IN | ~n39678;
  assign n39490 = ~n39489 | ~n39488;
  assign n39494 = ~n39491 & ~n39490;
  assign n39768 = ~n39492;
  assign n39493 = ~n39768 | ~n39639;
  assign P2_U2846 = ~n39494 | ~n39493;
  assign n39771 = ~P2_EBX_REG_8__SCAN_IN;
  assign n39509 = ~n39771 & ~n39495;
  assign n39777 = ~n39496;
  assign n39507 = ~n39777 | ~n39639;
  assign n39887 = ~n39497;
  assign n39500 = ~n39887 & ~n39628;
  assign n39499 = ~n39498 & ~n39683;
  assign n39505 = ~n39500 & ~n39499;
  assign n39502 = ~n39677 | ~P2_REIP_REG_8__SCAN_IN;
  assign n39501 = ~n39656 | ~P2_PHYADDRPOINTER_REG_8__SCAN_IN;
  assign n39503 = ~n39502 | ~n39501;
  assign n39504 = ~n40325 & ~n39503;
  assign n39506 = n39505 & n39504;
  assign n39508 = ~n39507 | ~n39506;
  assign n39515 = ~n39509 & ~n39508;
  assign n39512 = ~n42097 & ~n39510;
  assign n39513 = ~n39512 ^ n39511;
  assign n39514 = ~n39647 | ~n39513;
  assign P2_U2847 = ~n39515 | ~n39514;
  assign n39517 = ~n28361 & ~n39516;
  assign n39519 = ~n39517 & ~n40325;
  assign n39518 = ~n39656 | ~P2_PHYADDRPOINTER_REG_7__SCAN_IN;
  assign n39529 = ~n39519 | ~n39518;
  assign n39523 = ~n39521 | ~n39520;
  assign n39522 = ~n39678 | ~P2_EBX_REG_7__SCAN_IN;
  assign n39525 = ~n39523 | ~n39522;
  assign n39524 = ~n39893 & ~n39628;
  assign n39527 = ~n39525 & ~n39524;
  assign n39526 = ~n39787 | ~n39639;
  assign n39528 = ~n39527 | ~n39526;
  assign n39535 = ~n39529 & ~n39528;
  assign n39532 = ~n42095 | ~n39530;
  assign n39533 = ~n39532 ^ n39531;
  assign n39534 = ~n39533 | ~n39647;
  assign P2_U2848 = ~n39535 | ~n39534;
  assign n39542 = ~n39899 & ~n39628;
  assign n39537 = ~n39677 | ~P2_REIP_REG_6__SCAN_IN;
  assign n39536 = ~n39656 | ~P2_PHYADDRPOINTER_REG_6__SCAN_IN;
  assign n39538 = ~n39537 | ~n39536;
  assign n39540 = ~n40325 & ~n39538;
  assign n39539 = ~P2_EBX_REG_6__SCAN_IN | ~n39678;
  assign n39541 = ~n39540 | ~n39539;
  assign n39548 = ~n39542 & ~n39541;
  assign n39546 = ~n39543 & ~n39681;
  assign n39545 = ~n39544 & ~n39683;
  assign n39547 = ~n39546 & ~n39545;
  assign n39554 = n39548 & n39547;
  assign n39551 = ~n42097 & ~n39549;
  assign n39552 = ~n39551 ^ n39550;
  assign n39553 = ~n39647 | ~n39552;
  assign P2_U2849 = ~n39554 | ~n39553;
  assign n39556 = ~n39677 | ~P2_REIP_REG_5__SCAN_IN;
  assign n39555 = ~n39656 | ~P2_PHYADDRPOINTER_REG_5__SCAN_IN;
  assign n39557 = ~n39556 | ~n39555;
  assign n39563 = ~n40325 & ~n39557;
  assign n39917 = ~n39558;
  assign n39561 = ~n39917 & ~n39628;
  assign n39560 = ~n39559 & ~n39683;
  assign n39562 = ~n39561 & ~n39560;
  assign n39571 = ~n39563 | ~n39562;
  assign n39566 = ~n42095 | ~n39564;
  assign n39567 = ~n39566 ^ n39565;
  assign n39569 = ~n39567 | ~n39647;
  assign n39568 = ~P2_EBX_REG_5__SCAN_IN | ~n39678;
  assign n39570 = ~n39569 | ~n39568;
  assign n39573 = ~n39571 & ~n39570;
  assign n39572 = ~n39802 | ~n39639;
  assign P2_U2850 = ~n39573 | ~n39572;
  assign n39575 = ~n39677 | ~P2_REIP_REG_4__SCAN_IN;
  assign n39574 = ~n39678 | ~P2_EBX_REG_4__SCAN_IN;
  assign n39576 = ~n39575 | ~n39574;
  assign n39578 = ~n40325 & ~n39576;
  assign n39577 = ~n39656 | ~P2_PHYADDRPOINTER_REG_4__SCAN_IN;
  assign n39597 = ~n39578 | ~n39577;
  assign n39581 = ~n39579 | ~n39580;
  assign n40278 = ~n39582 | ~n39581;
  assign n39585 = ~n40278 & ~n39681;
  assign n39584 = ~n39583 & ~n39683;
  assign n39592 = n39585 | n39584;
  assign n39590 = ~n39586;
  assign n39589 = ~n39588 | ~n39587;
  assign n40357 = ~n39590 | ~n39589;
  assign n39591 = ~n40357 & ~n39628;
  assign n39595 = ~n39592 & ~n39591;
  assign n39780 = ~n22922 & ~n40497;
  assign n39916 = ~n39926;
  assign n39676 = n27370 & n39593;
  assign n39594 = ~n39916 | ~n39676;
  assign n39596 = ~n39595 | ~n39594;
  assign n39602 = ~n39597 & ~n39596;
  assign n39599 = ~n42097 & ~n39598;
  assign n39600 = ~n39599 ^ n40293;
  assign n39601 = ~n39647 | ~n39600;
  assign P2_U2851 = ~n39602 | ~n39601;
  assign n39604 = ~n39677 | ~P2_REIP_REG_3__SCAN_IN;
  assign n39603 = ~n39678 | ~P2_EBX_REG_3__SCAN_IN;
  assign n39611 = ~n39604 | ~n39603;
  assign n39607 = ~n42147 & ~n39628;
  assign n39606 = ~n39683 & ~n39605;
  assign n39609 = ~n39607 & ~n39606;
  assign n39608 = ~P2_PHYADDRPOINTER_REG_3__SCAN_IN | ~n39656;
  assign n39610 = ~n39609 | ~n39608;
  assign n39617 = ~n39611 & ~n39610;
  assign n39614 = ~n42095 | ~n39612;
  assign n39615 = ~n39614 ^ n39613;
  assign n39616 = ~n39615 | ~n39647;
  assign n39619 = ~n39617 | ~n39616;
  assign n39623 = ~n39619 & ~n39618;
  assign n42141 = ~n41490;
  assign n39622 = ~n42141 | ~n39676;
  assign P2_U2852 = ~n39623 | ~n39622;
  assign n39625 = ~n39677 | ~P2_REIP_REG_2__SCAN_IN;
  assign n39624 = ~n39678 | ~P2_EBX_REG_2__SCAN_IN;
  assign n39635 = ~n39625 | ~n39624;
  assign n39908 = ~n39627 ^ n39626;
  assign n42158 = ~n39908;
  assign n39631 = ~n42158 & ~n39628;
  assign n39630 = ~n39683 & ~n39629;
  assign n39633 = ~n39631 & ~n39630;
  assign n39632 = ~P2_PHYADDRPOINTER_REG_2__SCAN_IN | ~n39656;
  assign n39634 = ~n39633 | ~n39632;
  assign n39643 = ~n39635 & ~n39634;
  assign n42156 = ~n39637 ^ n39636;
  assign n39638 = ~n39676;
  assign n39641 = n42156 | n39638;
  assign n39640 = ~n27757 | ~n39639;
  assign n39642 = n39641 & n39640;
  assign n39649 = n39643 & n39642;
  assign n39645 = ~n42097 & ~n39644;
  assign n39646 = ~n39645 ^ n40303;
  assign n39648 = ~n39647 | ~n39646;
  assign P2_U2853 = ~n39649 | ~n39648;
  assign n39651 = ~n42170 | ~n39676;
  assign n39650 = ~n39673 | ~n40329;
  assign n39655 = ~n39651 | ~n39650;
  assign n42094 = ~n39675 ^ n39652;
  assign n39654 = ~n39653 & ~n42094;
  assign n39671 = ~n39655 & ~n39654;
  assign n39658 = ~n39677 | ~P2_REIP_REG_1__SCAN_IN;
  assign n39657 = ~n39656 | ~P2_PHYADDRPOINTER_REG_1__SCAN_IN;
  assign n39664 = ~n39658 | ~n39657;
  assign n39662 = ~P2_EBX_REG_1__SCAN_IN | ~n39678;
  assign n39959 = ~n39660 ^ n39659;
  assign n39661 = ~n39686 | ~n39959;
  assign n39663 = ~n39662 | ~n39661;
  assign n39669 = ~n39664 & ~n39663;
  assign n39666 = ~n39683 & ~n39665;
  assign n39668 = ~n39667 & ~n39666;
  assign n39670 = n39669 & n39668;
  assign P2_U2854 = ~n39671 | ~n39670;
  assign n39674 = n39673 | n39672;
  assign n39696 = ~n39674 | ~P2_PHYADDRPOINTER_REG_0__SCAN_IN;
  assign n42093 = ~n42095 | ~n39675;
  assign n39694 = ~n41893 & ~n42093;
  assign n39692 = ~n42177 | ~n39676;
  assign n39680 = ~n39677 | ~P2_REIP_REG_0__SCAN_IN;
  assign n39679 = ~n39678 | ~P2_EBX_REG_0__SCAN_IN;
  assign n39690 = ~n39680 | ~n39679;
  assign n39685 = ~n40343 & ~n39681;
  assign n39684 = ~n39683 & ~n39682;
  assign n39688 = ~n39685 & ~n39684;
  assign n39687 = ~n39686 | ~n39963;
  assign n39689 = ~n39688 | ~n39687;
  assign n39691 = ~n39690 & ~n39689;
  assign n39693 = ~n39692 | ~n39691;
  assign n39695 = ~n39694 & ~n39693;
  assign P2_U2855 = ~n39696 | ~n39695;
  assign n39703 = ~n31948 & ~n39697;
  assign n39700 = n39699 | n39698;
  assign n39832 = ~n39701 | ~n39700;
  assign n39702 = ~n39832 & ~n39814;
  assign n39706 = ~n39703 & ~n39702;
  assign n39705 = ~n39704 | ~n31948;
  assign P2_U2871 = ~n39706 | ~n39705;
  assign n39712 = ~n31948 & ~n39707;
  assign n39710 = ~n39709 ^ n39708;
  assign n39711 = ~n39710 & ~n39814;
  assign n39715 = ~n39712 & ~n39711;
  assign n39714 = ~n39713 | ~n31948;
  assign P2_U2872 = ~n39715 | ~n39714;
  assign n39720 = ~n31948 & ~n39716;
  assign n39718 = ~n39729 ^ n39717;
  assign n39719 = ~n39718 & ~n39814;
  assign n39723 = ~n39720 & ~n39719;
  assign n39722 = ~n39721 | ~n31948;
  assign P2_U2873 = ~n39723 | ~n39722;
  assign n39731 = ~n31948 & ~n39724;
  assign n39727 = ~n39726 | ~n39725;
  assign n39728 = ~n39727 | ~n39782;
  assign n39730 = ~n39729 & ~n39728;
  assign n39734 = ~n39731 & ~n39730;
  assign n39733 = ~n39732 | ~n31948;
  assign P2_U2874 = ~n39734 | ~n39733;
  assign n39735 = ~P2_EBX_REG_12__SCAN_IN;
  assign n39740 = ~n31948 & ~n39735;
  assign n39764 = ~n22907 | ~n39762;
  assign n39755 = ~n39736;
  assign n39745 = ~n39764 & ~n39755;
  assign n39747 = ~n39745 | ~n39744;
  assign n39738 = n39737 ^ n39747;
  assign n39739 = ~n39738 & ~n39814;
  assign n39743 = ~n39740 & ~n39739;
  assign n39742 = ~n39741 | ~n31948;
  assign P2_U2875 = ~n39743 | ~n39742;
  assign n39750 = n39817 & P2_EBX_REG_11__SCAN_IN;
  assign n39746 = ~n39745 & ~n39744;
  assign n39748 = ~n39746 & ~n39814;
  assign n39749 = n39748 & n39747;
  assign n39753 = ~n39750 & ~n39749;
  assign n39752 = ~n39751 | ~n31948;
  assign P2_U2876 = ~n39753 | ~n39752;
  assign n39758 = ~n31948 & ~n39754;
  assign n39756 = ~n39764 ^ n39755;
  assign n39757 = ~n39756 & ~n39814;
  assign n39761 = ~n39758 & ~n39757;
  assign n39760 = ~n39759 | ~n31948;
  assign P2_U2877 = ~n39761 | ~n39760;
  assign n39767 = n39817 & P2_EBX_REG_9__SCAN_IN;
  assign n39763 = ~n22907 & ~n39762;
  assign n39765 = ~n39763 & ~n39814;
  assign n39766 = n39765 & n39764;
  assign n39770 = ~n39767 & ~n39766;
  assign n39769 = ~n39768 | ~n31948;
  assign P2_U2878 = ~n39770 | ~n39769;
  assign n39776 = ~n31948 & ~n39771;
  assign n39774 = ~n39772 ^ n39773;
  assign n39775 = ~n39774 & ~n39814;
  assign n39779 = ~n39776 & ~n39775;
  assign n39778 = ~n39777 | ~n31948;
  assign P2_U2879 = ~n39779 | ~n39778;
  assign n39786 = n39817 & P2_EBX_REG_7__SCAN_IN;
  assign n39798 = ~n23056 | ~P2_INSTQUEUE_REG_0__5__SCAN_IN;
  assign n39781 = ~n39798 & ~n40530;
  assign n39784 = ~n39781 & ~P2_INSTQUEUE_REG_0__7__SCAN_IN;
  assign n39783 = ~n39772 | ~n39782;
  assign n39785 = ~n39784 & ~n39783;
  assign n39789 = ~n39786 & ~n39785;
  assign n39788 = ~n39787 | ~n31948;
  assign P2_U2880 = ~n39789 | ~n39788;
  assign n39793 = ~n31948 & ~n39790;
  assign n39791 = P2_INSTQUEUE_REG_0__6__SCAN_IN ^ n39798;
  assign n39792 = ~n39791 & ~n39814;
  assign n39796 = ~n39793 & ~n39792;
  assign n39795 = ~n39794 | ~n31948;
  assign P2_U2881 = ~n39796 | ~n39795;
  assign n39801 = n39817 & P2_EBX_REG_5__SCAN_IN;
  assign n39797 = ~n23056 & ~P2_INSTQUEUE_REG_0__5__SCAN_IN;
  assign n39799 = ~n39797 & ~n39814;
  assign n39800 = n39799 & n39798;
  assign n39804 = ~n39801 & ~n39800;
  assign n39803 = ~n39802 | ~n31948;
  assign P2_U2882 = ~n39804 | ~n39803;
  assign n39806 = ~n39916 | ~n39805;
  assign n39807 = ~n39806 | ~n40278;
  assign n39809 = ~n39807 | ~n31948;
  assign n39808 = ~P2_EBX_REG_4__SCAN_IN | ~n39817;
  assign P2_U2883 = ~n39809 | ~n39808;
  assign n39811 = ~n41490 & ~n39814;
  assign n39813 = ~n39811 & ~n39810;
  assign n39812 = ~P2_EBX_REG_3__SCAN_IN | ~n39817;
  assign P2_U2884 = ~n39813 | ~n39812;
  assign n39816 = n42156 | n39814;
  assign n39815 = ~n27757 | ~n31948;
  assign n39819 = n39816 & n39815;
  assign n39818 = ~P2_EBX_REG_2__SCAN_IN | ~n39817;
  assign P2_U2885 = ~n39819 | ~n39818;
  assign n39821 = ~n39820;
  assign n39825 = ~n39821 & ~n39945;
  assign n39823 = ~n39839 | ~BUF1_REG_31__SCAN_IN;
  assign n39822 = ~P2_EAX_REG_31__SCAN_IN | ~n39970;
  assign n39824 = ~n39823 | ~n39822;
  assign n39827 = ~n39825 & ~n39824;
  assign n39826 = ~BUF2_REG_31__SCAN_IN | ~n39828;
  assign P2_U2888 = ~n39827 | ~n39826;
  assign n39831 = ~BUF2_REG_16__SCAN_IN | ~n39828;
  assign n39830 = ~n39829 | ~n31972;
  assign n39834 = ~n39831 | ~n39830;
  assign n39952 = ~n39964;
  assign n39833 = ~n39832 & ~n39952;
  assign n39845 = ~n39834 & ~n39833;
  assign n39838 = ~n39835;
  assign n39837 = ~n40435 | ~BUF1_REG_0__SCAN_IN;
  assign n39836 = ~BUF2_REG_0__SCAN_IN | ~n40437;
  assign n39843 = ~n39838 & ~n40429;
  assign n39841 = ~n39839 | ~BUF1_REG_16__SCAN_IN;
  assign n39840 = ~P2_EAX_REG_16__SCAN_IN | ~n39970;
  assign n39842 = ~n39841 | ~n39840;
  assign n39844 = ~n39843 & ~n39842;
  assign P2_U2903 = ~n39845 | ~n39844;
  assign n39848 = ~n39846 & ~n39898;
  assign n39847 = ~n28956 & ~n39888;
  assign n39854 = ~n39848 & ~n39847;
  assign n39962 = ~n39850 | ~n39849;
  assign n39852 = ~n40437 | ~BUF2_REG_15__SCAN_IN;
  assign n39851 = ~n40435 | ~BUF1_REG_15__SCAN_IN;
  assign n40271 = ~n39852 | ~n39851;
  assign n39853 = ~n39954 | ~n40271;
  assign P2_U2904 = ~n39854 | ~n39853;
  assign n39857 = ~n39855 & ~n39898;
  assign n39856 = ~n28912 & ~n39888;
  assign n39859 = ~n39857 & ~n39856;
  assign n39858 = ~n39954 | ~n40195;
  assign P2_U2905 = ~n39859 | ~n39858;
  assign n39862 = ~n39860 & ~n39898;
  assign n39861 = ~n28872 & ~n39888;
  assign n39864 = ~n39862 & ~n39861;
  assign n39863 = ~n39954 | ~n40189;
  assign P2_U2906 = ~n39864 | ~n39863;
  assign n39867 = ~n39865 & ~n39898;
  assign n39866 = ~n28828 & ~n39888;
  assign n39869 = ~n39867 & ~n39866;
  assign n39868 = ~n39954 | ~n40183;
  assign P2_U2907 = ~n39869 | ~n39868;
  assign n39871 = ~n39870;
  assign n39873 = ~n39871 & ~n39898;
  assign n39872 = ~n28791 & ~n39888;
  assign n39875 = ~n39873 & ~n39872;
  assign n39874 = ~n39954 | ~n40177;
  assign P2_U2908 = ~n39875 | ~n39874;
  assign n39878 = ~n39876 & ~n39898;
  assign n39877 = ~n28748 & ~n39888;
  assign n39880 = ~n39878 & ~n39877;
  assign n39879 = ~n39954 | ~n40171;
  assign P2_U2909 = ~n39880 | ~n39879;
  assign n39882 = ~n39881;
  assign n39884 = ~n39882 & ~n39898;
  assign n39883 = ~n28707 & ~n39888;
  assign n39886 = ~n39884 & ~n39883;
  assign n39885 = ~n39954 | ~n40165;
  assign P2_U2910 = ~n39886 | ~n39885;
  assign n39890 = ~n39887 & ~n39898;
  assign n39889 = ~n28661 & ~n39888;
  assign n39892 = ~n39890 & ~n39889;
  assign n39891 = ~n39954 | ~n40159;
  assign P2_U2911 = ~n39892 | ~n39891;
  assign n39895 = ~n39893 & ~n39898;
  assign n40154 = ~n40565;
  assign n39894 = ~n39962 & ~n40154;
  assign n39897 = ~n39895 & ~n39894;
  assign n39896 = ~P2_EAX_REG_7__SCAN_IN | ~n39970;
  assign P2_U2912 = ~n39897 | ~n39896;
  assign n39901 = ~n39899 & ~n39898;
  assign n40149 = ~n40543;
  assign n39900 = ~n39962 & ~n40149;
  assign n39903 = ~n39901 & ~n39900;
  assign n39902 = ~P2_EAX_REG_6__SCAN_IN | ~n39970;
  assign P2_U2913 = ~n39903 | ~n39902;
  assign n39907 = ~n39917 & ~n39945;
  assign n39905 = ~P2_EAX_REG_5__SCAN_IN | ~n39970;
  assign n39904 = ~n39954 | ~n40528;
  assign n39906 = ~n39905 | ~n39904;
  assign n39921 = ~n39907 & ~n39906;
  assign n39914 = ~n41490 | ~n42147;
  assign n39935 = n42147 ^ n41490;
  assign n39912 = ~n42156 | ~n42158;
  assign n39940 = ~n42156 ^ n39908;
  assign n42166 = ~n39959;
  assign n39910 = ~n42112 | ~n42166;
  assign n39950 = ~n42112 ^ n39959;
  assign n39951 = ~n42177 | ~n39963;
  assign n39909 = ~n39950 | ~n39951;
  assign n39941 = ~n39910 | ~n39909;
  assign n39911 = ~n39940 | ~n39941;
  assign n39936 = ~n39912 | ~n39911;
  assign n39913 = ~n39935 | ~n39936;
  assign n39915 = ~n39914 | ~n39913;
  assign n39927 = ~n39915 | ~n40357;
  assign n39918 = ~n39916 | ~n39927;
  assign n39919 = ~n39918 | ~n39917;
  assign n39920 = ~n39919 | ~n39964;
  assign P2_U2914 = ~n39921 | ~n39920;
  assign n39923 = ~P2_EAX_REG_4__SCAN_IN | ~n39970;
  assign n39922 = ~n39954 | ~n40510;
  assign n39925 = ~n39923 | ~n39922;
  assign n39924 = ~n40357 & ~n39945;
  assign n39930 = ~n39925 & ~n39924;
  assign n39928 = ~n39927 ^ n39926;
  assign n39929 = ~n39928 | ~n39964;
  assign P2_U2915 = ~n39930 | ~n39929;
  assign n39932 = ~P2_EAX_REG_3__SCAN_IN | ~n39970;
  assign n39931 = ~n39954 | ~n40495;
  assign n39934 = ~n39932 | ~n39931;
  assign n39933 = ~n42147 & ~n39945;
  assign n39939 = ~n39934 & ~n39933;
  assign n39937 = ~n39936 ^ n39935;
  assign n39938 = ~n39937 | ~n39964;
  assign P2_U2916 = ~n39939 | ~n39938;
  assign n39942 = ~n39941 ^ n39940;
  assign n39949 = ~n39942 | ~n39964;
  assign n39944 = ~P2_EAX_REG_2__SCAN_IN | ~n39970;
  assign n39943 = ~n39954 | ~n40480;
  assign n39947 = ~n39944 | ~n39943;
  assign n39946 = ~n42158 & ~n39945;
  assign n39948 = ~n39947 & ~n39946;
  assign P2_U2917 = ~n39949 | ~n39948;
  assign n39953 = n39951 ^ n39950;
  assign n39958 = ~n39953 & ~n39952;
  assign n39956 = ~P2_EAX_REG_1__SCAN_IN | ~n39970;
  assign n39955 = ~n39954 | ~n40465;
  assign n39957 = ~n39956 | ~n39955;
  assign n39961 = ~n39958 & ~n39957;
  assign n39960 = ~n31972 | ~n39959;
  assign P2_U2918 = ~n39961 | ~n39960;
  assign n39969 = ~n39962 & ~n40429;
  assign n39967 = ~n31972 | ~n39963;
  assign n39965 = ~n41491 ^ n39963;
  assign n39966 = ~n39965 | ~n39964;
  assign n39968 = ~n39967 | ~n39966;
  assign n39972 = ~n39969 & ~n39968;
  assign n39971 = ~P2_EAX_REG_0__SCAN_IN | ~n39970;
  assign P2_U2919 = ~n39972 | ~n39971;
  assign n39974 = ~n39973 & ~n42075;
  assign n42213 = ~n41909;
  assign P2_U2920 = ~n40076 & ~n39977;
  assign n39979 = ~P2_DATAO_REG_30__SCAN_IN | ~n40114;
  assign n39978 = ~P2_UWORD_REG_14__SCAN_IN | ~n42199;
  assign n39981 = n39979 & n39978;
  assign n39980 = ~n40037 | ~P2_EAX_REG_30__SCAN_IN;
  assign P2_U2921 = ~n39981 | ~n39980;
  assign n39983 = ~n40114 | ~P2_DATAO_REG_29__SCAN_IN;
  assign n39982 = ~P2_UWORD_REG_13__SCAN_IN | ~n40022;
  assign n39985 = n39983 & n39982;
  assign n39984 = ~n40037 | ~P2_EAX_REG_29__SCAN_IN;
  assign P2_U2922 = ~n39985 | ~n39984;
  assign n39987 = ~P2_DATAO_REG_28__SCAN_IN | ~n40114;
  assign n39986 = ~P2_UWORD_REG_12__SCAN_IN | ~n40022;
  assign n39989 = n39987 & n39986;
  assign n39988 = ~n40037 | ~P2_EAX_REG_28__SCAN_IN;
  assign P2_U2923 = ~n39989 | ~n39988;
  assign n39991 = ~n40108 | ~P2_DATAO_REG_27__SCAN_IN;
  assign n39990 = ~P2_UWORD_REG_11__SCAN_IN | ~n40022;
  assign n39993 = n39991 & n39990;
  assign n39992 = ~n40037 | ~P2_EAX_REG_27__SCAN_IN;
  assign P2_U2924 = ~n39993 | ~n39992;
  assign n39995 = ~n40114 | ~P2_DATAO_REG_26__SCAN_IN;
  assign n39994 = ~P2_UWORD_REG_10__SCAN_IN | ~n40022;
  assign n39997 = n39995 & n39994;
  assign n39996 = ~n40037 | ~P2_EAX_REG_26__SCAN_IN;
  assign P2_U2925 = ~n39997 | ~n39996;
  assign n39999 = ~P2_DATAO_REG_25__SCAN_IN | ~n40114;
  assign n39998 = ~P2_UWORD_REG_9__SCAN_IN | ~n40022;
  assign n40001 = n39999 & n39998;
  assign n40000 = ~n40037 | ~P2_EAX_REG_25__SCAN_IN;
  assign P2_U2926 = ~n40001 | ~n40000;
  assign n40003 = ~n40114 | ~P2_DATAO_REG_24__SCAN_IN;
  assign n40002 = ~P2_UWORD_REG_8__SCAN_IN | ~n40022;
  assign n40005 = n40003 & n40002;
  assign n40004 = ~n40037 | ~P2_EAX_REG_24__SCAN_IN;
  assign P2_U2927 = ~n40005 | ~n40004;
  assign n40007 = ~P2_DATAO_REG_23__SCAN_IN | ~n40114;
  assign n40006 = ~P2_UWORD_REG_7__SCAN_IN | ~n40022;
  assign n40009 = n40007 & n40006;
  assign n40008 = ~n40037 | ~P2_EAX_REG_23__SCAN_IN;
  assign P2_U2928 = ~n40009 | ~n40008;
  assign n40011 = ~n40114 | ~P2_DATAO_REG_22__SCAN_IN;
  assign n40010 = ~P2_UWORD_REG_6__SCAN_IN | ~n40022;
  assign n40013 = n40011 & n40010;
  assign n40012 = ~n40037 | ~P2_EAX_REG_22__SCAN_IN;
  assign P2_U2929 = ~n40013 | ~n40012;
  assign n40015 = ~P2_DATAO_REG_21__SCAN_IN | ~n40114;
  assign n40014 = ~P2_UWORD_REG_5__SCAN_IN | ~n40022;
  assign n40017 = n40015 & n40014;
  assign n40016 = ~n40037 | ~P2_EAX_REG_21__SCAN_IN;
  assign P2_U2930 = ~n40017 | ~n40016;
  assign n40019 = ~P2_DATAO_REG_20__SCAN_IN | ~n40114;
  assign n40018 = ~P2_UWORD_REG_4__SCAN_IN | ~n40022;
  assign n40021 = n40019 & n40018;
  assign n40020 = ~n40037 | ~P2_EAX_REG_20__SCAN_IN;
  assign P2_U2931 = ~n40021 | ~n40020;
  assign n40024 = ~P2_DATAO_REG_19__SCAN_IN | ~n40114;
  assign n40023 = ~P2_UWORD_REG_3__SCAN_IN | ~n40022;
  assign n40026 = n40024 & n40023;
  assign n40025 = ~n40037 | ~P2_EAX_REG_19__SCAN_IN;
  assign P2_U2932 = ~n40026 | ~n40025;
  assign n40028 = ~n40108 | ~P2_DATAO_REG_18__SCAN_IN;
  assign n40027 = ~P2_UWORD_REG_2__SCAN_IN | ~n42199;
  assign n40030 = n40028 & n40027;
  assign n40029 = ~n40037 | ~P2_EAX_REG_18__SCAN_IN;
  assign P2_U2933 = ~n40030 | ~n40029;
  assign n40032 = ~P2_DATAO_REG_17__SCAN_IN | ~n40114;
  assign n40031 = ~P2_UWORD_REG_1__SCAN_IN | ~n42199;
  assign n40034 = n40032 & n40031;
  assign n40033 = ~n40037 | ~P2_EAX_REG_17__SCAN_IN;
  assign P2_U2934 = ~n40034 | ~n40033;
  assign n40036 = ~P2_DATAO_REG_16__SCAN_IN | ~n40114;
  assign n40035 = ~P2_UWORD_REG_0__SCAN_IN | ~n42199;
  assign n40039 = n40036 & n40035;
  assign n40038 = ~n40037 | ~P2_EAX_REG_16__SCAN_IN;
  assign P2_U2935 = ~n40039 | ~n40038;
  assign n40042 = ~n40076 & ~n40040;
  assign n40041 = ~n28956 & ~n40077;
  assign n40044 = ~n40042 & ~n40041;
  assign n40043 = ~n42199 | ~P2_LWORD_REG_15__SCAN_IN;
  assign P2_U2936 = ~n40044 | ~n40043;
  assign n40047 = ~n40076 & ~n40045;
  assign n40046 = ~n28912 & ~n40077;
  assign n40049 = ~n40047 & ~n40046;
  assign n40048 = ~n42199 | ~P2_LWORD_REG_14__SCAN_IN;
  assign P2_U2937 = ~n40049 | ~n40048;
  assign n40052 = ~n40076 & ~n40050;
  assign n40051 = ~n28872 & ~n40077;
  assign n40054 = ~n40052 & ~n40051;
  assign n40053 = ~n42199 | ~P2_LWORD_REG_13__SCAN_IN;
  assign P2_U2938 = ~n40054 | ~n40053;
  assign n40057 = ~n40076 & ~n40055;
  assign n40056 = ~n28828 & ~n40077;
  assign n40059 = ~n40057 & ~n40056;
  assign n40058 = ~n42199 | ~P2_LWORD_REG_12__SCAN_IN;
  assign P2_U2939 = ~n40059 | ~n40058;
  assign n40062 = ~n40076 & ~n40060;
  assign n40061 = ~n28791 & ~n40077;
  assign n40064 = ~n40062 & ~n40061;
  assign n40063 = ~n42199 | ~P2_LWORD_REG_11__SCAN_IN;
  assign P2_U2940 = ~n40064 | ~n40063;
  assign n40067 = ~n40076 & ~n40065;
  assign n40066 = ~n28748 & ~n40077;
  assign n40069 = ~n40067 & ~n40066;
  assign n40068 = ~n42199 | ~P2_LWORD_REG_10__SCAN_IN;
  assign P2_U2941 = ~n40069 | ~n40068;
  assign n40072 = ~n40076 & ~n40070;
  assign n40071 = ~n28707 & ~n40077;
  assign n40074 = ~n40072 & ~n40071;
  assign n40073 = ~n42199 | ~P2_LWORD_REG_9__SCAN_IN;
  assign P2_U2942 = ~n40074 | ~n40073;
  assign n40079 = ~n40076 & ~n40075;
  assign n40078 = ~n28661 & ~n40077;
  assign n40081 = ~n40079 & ~n40078;
  assign n40080 = ~n42199 | ~P2_LWORD_REG_8__SCAN_IN;
  assign P2_U2943 = ~n40081 | ~n40080;
  assign n40083 = ~P2_LWORD_REG_7__SCAN_IN | ~n42199;
  assign n40082 = ~n40111 | ~P2_EAX_REG_7__SCAN_IN;
  assign n40085 = n40083 & n40082;
  assign n40084 = ~n40114 | ~P2_DATAO_REG_7__SCAN_IN;
  assign P2_U2944 = ~n40085 | ~n40084;
  assign n40087 = ~P2_LWORD_REG_6__SCAN_IN | ~n42199;
  assign n40086 = ~n40111 | ~P2_EAX_REG_6__SCAN_IN;
  assign n40089 = n40087 & n40086;
  assign n40088 = ~n40108 | ~P2_DATAO_REG_6__SCAN_IN;
  assign P2_U2945 = ~n40089 | ~n40088;
  assign n40091 = ~P2_LWORD_REG_5__SCAN_IN | ~n42199;
  assign n40090 = ~n40111 | ~P2_EAX_REG_5__SCAN_IN;
  assign n40093 = n40091 & n40090;
  assign n40092 = ~n40108 | ~P2_DATAO_REG_5__SCAN_IN;
  assign P2_U2946 = ~n40093 | ~n40092;
  assign n40095 = ~P2_LWORD_REG_4__SCAN_IN | ~n42199;
  assign n40094 = ~n40111 | ~P2_EAX_REG_4__SCAN_IN;
  assign n40097 = n40095 & n40094;
  assign n40096 = ~n40108 | ~P2_DATAO_REG_4__SCAN_IN;
  assign P2_U2947 = ~n40097 | ~n40096;
  assign n40099 = ~P2_LWORD_REG_3__SCAN_IN | ~n42199;
  assign n40098 = ~n40111 | ~P2_EAX_REG_3__SCAN_IN;
  assign n40101 = n40099 & n40098;
  assign n40100 = ~n40108 | ~P2_DATAO_REG_3__SCAN_IN;
  assign P2_U2948 = ~n40101 | ~n40100;
  assign n40103 = ~P2_LWORD_REG_2__SCAN_IN | ~n42199;
  assign n40102 = ~n40111 | ~P2_EAX_REG_2__SCAN_IN;
  assign n40105 = n40103 & n40102;
  assign n40104 = ~n40108 | ~P2_DATAO_REG_2__SCAN_IN;
  assign P2_U2949 = ~n40105 | ~n40104;
  assign n40107 = ~P2_LWORD_REG_1__SCAN_IN | ~n42199;
  assign n40106 = ~n40111 | ~P2_EAX_REG_1__SCAN_IN;
  assign n40110 = n40107 & n40106;
  assign n40109 = ~n40108 | ~P2_DATAO_REG_1__SCAN_IN;
  assign P2_U2950 = ~n40110 | ~n40109;
  assign n40113 = ~P2_LWORD_REG_0__SCAN_IN | ~n42199;
  assign n40112 = ~n40111 | ~P2_EAX_REG_0__SCAN_IN;
  assign n40116 = n40113 & n40112;
  assign n40115 = ~n40114 | ~P2_DATAO_REG_0__SCAN_IN;
  assign P2_U2951 = ~n40116 | ~n40115;
  assign n40120 = ~n40117 & ~n41895;
  assign n40201 = ~n40273 & ~n40429;
  assign n40119 = ~n40226 & ~n40118;
  assign n40122 = ~n40201 & ~n40119;
  assign n40270 = ~n40120 & ~n40200;
  assign n40121 = ~P2_UWORD_REG_0__SCAN_IN | ~n40270;
  assign P2_U2952 = ~n40122 | ~n40121;
  assign n40125 = ~n40226 & ~n40123;
  assign n40124 = ~n40465;
  assign n40206 = ~n40273 & ~n40124;
  assign n40127 = ~n40125 & ~n40206;
  assign n40126 = ~n40270 | ~P2_UWORD_REG_1__SCAN_IN;
  assign P2_U2953 = ~n40127 | ~n40126;
  assign n40130 = ~n40226 & ~n40128;
  assign n40129 = ~n40480;
  assign n40211 = ~n40273 & ~n40129;
  assign n40132 = ~n40130 & ~n40211;
  assign n40131 = ~n40270 | ~P2_UWORD_REG_2__SCAN_IN;
  assign P2_U2954 = ~n40132 | ~n40131;
  assign n40135 = ~n40226 & ~n40133;
  assign n40134 = ~n40495;
  assign n40216 = ~n40273 & ~n40134;
  assign n40137 = ~n40135 & ~n40216;
  assign n40136 = ~n40270 | ~P2_UWORD_REG_3__SCAN_IN;
  assign P2_U2955 = ~n40137 | ~n40136;
  assign n40140 = ~n40226 & ~n40138;
  assign n40139 = ~n40510;
  assign n40221 = ~n40273 & ~n40139;
  assign n40142 = ~n40140 & ~n40221;
  assign n40141 = ~n40270 | ~P2_UWORD_REG_4__SCAN_IN;
  assign P2_U2956 = ~n40142 | ~n40141;
  assign n40226 = ~n40200;
  assign n40145 = ~n40226 & ~n40143;
  assign n40144 = ~n40528;
  assign n40227 = ~n40273 & ~n40144;
  assign n40147 = ~n40145 & ~n40227;
  assign n40146 = ~n40270 | ~P2_UWORD_REG_5__SCAN_IN;
  assign P2_U2957 = ~n40147 | ~n40146;
  assign n40150 = ~n40226 & ~n40148;
  assign n40232 = ~n40273 & ~n40149;
  assign n40152 = ~n40150 & ~n40232;
  assign n40151 = ~n40270 | ~P2_UWORD_REG_6__SCAN_IN;
  assign P2_U2958 = ~n40152 | ~n40151;
  assign n40155 = ~n40226 & ~n40153;
  assign n40237 = ~n40273 & ~n40154;
  assign n40157 = ~n40155 & ~n40237;
  assign n40156 = ~n40270 | ~P2_UWORD_REG_7__SCAN_IN;
  assign P2_U2959 = ~n40157 | ~n40156;
  assign n40161 = ~n40226 & ~n40158;
  assign n40160 = ~n40159;
  assign n40241 = ~n40273 & ~n40160;
  assign n40163 = ~n40161 & ~n40241;
  assign n40162 = ~n40270 | ~P2_UWORD_REG_8__SCAN_IN;
  assign P2_U2960 = ~n40163 | ~n40162;
  assign n40167 = ~n40226 & ~n40164;
  assign n40166 = ~n40165;
  assign n40245 = ~n40273 & ~n40166;
  assign n40169 = ~n40167 & ~n40245;
  assign n40168 = ~n40270 | ~P2_UWORD_REG_9__SCAN_IN;
  assign P2_U2961 = ~n40169 | ~n40168;
  assign n40173 = ~n40226 & ~n40170;
  assign n40172 = ~n40171;
  assign n40250 = ~n40273 & ~n40172;
  assign n40175 = ~n40173 & ~n40250;
  assign n40174 = ~n40270 | ~P2_UWORD_REG_10__SCAN_IN;
  assign P2_U2962 = ~n40175 | ~n40174;
  assign n40176 = ~P2_EAX_REG_27__SCAN_IN;
  assign n40179 = ~n40249 & ~n40176;
  assign n40178 = ~n40177;
  assign n40254 = ~n40273 & ~n40178;
  assign n40181 = ~n40179 & ~n40254;
  assign n40180 = ~n40270 | ~P2_UWORD_REG_11__SCAN_IN;
  assign P2_U2963 = ~n40181 | ~n40180;
  assign n40185 = ~n40226 & ~n40182;
  assign n40184 = ~n40183;
  assign n40258 = ~n40273 & ~n40184;
  assign n40187 = ~n40185 & ~n40258;
  assign n40186 = ~n40270 | ~P2_UWORD_REG_12__SCAN_IN;
  assign P2_U2964 = ~n40187 | ~n40186;
  assign n40188 = ~P2_EAX_REG_29__SCAN_IN;
  assign n40191 = ~n40226 & ~n40188;
  assign n40190 = ~n40189;
  assign n40262 = ~n40273 & ~n40190;
  assign n40193 = ~n40191 & ~n40262;
  assign n40192 = ~n40270 | ~P2_UWORD_REG_13__SCAN_IN;
  assign P2_U2965 = ~n40193 | ~n40192;
  assign n40197 = ~n40249 & ~n40194;
  assign n40196 = ~n40195;
  assign n40266 = ~n40273 & ~n40196;
  assign n40199 = ~n40197 & ~n40266;
  assign n40198 = ~n40270 | ~P2_UWORD_REG_14__SCAN_IN;
  assign P2_U2966 = ~n40199 | ~n40198;
  assign n40202 = n40200 & P2_EAX_REG_0__SCAN_IN;
  assign n40204 = ~n40202 & ~n40201;
  assign n40203 = ~P2_LWORD_REG_0__SCAN_IN | ~n40270;
  assign P2_U2967 = ~n40204 | ~n40203;
  assign n40207 = ~n40226 & ~n40205;
  assign n40209 = ~n40207 & ~n40206;
  assign n40208 = ~n40270 | ~P2_LWORD_REG_1__SCAN_IN;
  assign P2_U2968 = ~n40209 | ~n40208;
  assign n40212 = ~n40226 & ~n40210;
  assign n40214 = ~n40212 & ~n40211;
  assign n40213 = ~n40270 | ~P2_LWORD_REG_2__SCAN_IN;
  assign P2_U2969 = ~n40214 | ~n40213;
  assign n40217 = ~n40226 & ~n40215;
  assign n40219 = ~n40217 & ~n40216;
  assign n40218 = ~n40270 | ~P2_LWORD_REG_3__SCAN_IN;
  assign P2_U2970 = ~n40219 | ~n40218;
  assign n40222 = ~n40226 & ~n40220;
  assign n40224 = ~n40222 & ~n40221;
  assign n40223 = ~n40270 | ~P2_LWORD_REG_4__SCAN_IN;
  assign P2_U2971 = ~n40224 | ~n40223;
  assign n40228 = ~n40226 & ~n40225;
  assign n40230 = ~n40228 & ~n40227;
  assign n40229 = ~n40270 | ~P2_LWORD_REG_5__SCAN_IN;
  assign P2_U2972 = ~n40230 | ~n40229;
  assign n40233 = ~n40249 & ~n40231;
  assign n40235 = ~n40233 & ~n40232;
  assign n40234 = ~n40270 | ~P2_LWORD_REG_6__SCAN_IN;
  assign P2_U2973 = ~n40235 | ~n40234;
  assign n40238 = ~n40226 & ~n40236;
  assign n40240 = ~n40238 & ~n40237;
  assign n40239 = ~n40270 | ~P2_LWORD_REG_7__SCAN_IN;
  assign P2_U2974 = ~n40240 | ~n40239;
  assign n40242 = ~n40249 & ~n28661;
  assign n40244 = ~n40242 & ~n40241;
  assign n40243 = ~n40270 | ~P2_LWORD_REG_8__SCAN_IN;
  assign P2_U2975 = ~n40244 | ~n40243;
  assign n40246 = ~n40249 & ~n28707;
  assign n40248 = ~n40246 & ~n40245;
  assign n40247 = ~n40270 | ~P2_LWORD_REG_9__SCAN_IN;
  assign P2_U2976 = ~n40248 | ~n40247;
  assign n40251 = ~n40249 & ~n28748;
  assign n40253 = ~n40251 & ~n40250;
  assign n40252 = ~n40270 | ~P2_LWORD_REG_10__SCAN_IN;
  assign P2_U2977 = ~n40253 | ~n40252;
  assign n40255 = ~n40226 & ~n28791;
  assign n40257 = ~n40255 & ~n40254;
  assign n40256 = ~n40270 | ~P2_LWORD_REG_11__SCAN_IN;
  assign P2_U2978 = ~n40257 | ~n40256;
  assign n40259 = ~n40226 & ~n28828;
  assign n40261 = ~n40259 & ~n40258;
  assign n40260 = ~n40270 | ~P2_LWORD_REG_12__SCAN_IN;
  assign P2_U2979 = ~n40261 | ~n40260;
  assign n40263 = ~n40226 & ~n28872;
  assign n40265 = ~n40263 & ~n40262;
  assign n40264 = ~n40270 | ~P2_LWORD_REG_13__SCAN_IN;
  assign P2_U2980 = ~n40265 | ~n40264;
  assign n40267 = ~n40226 & ~n28912;
  assign n40269 = ~n40267 & ~n40266;
  assign n40268 = ~n40270 | ~P2_LWORD_REG_14__SCAN_IN;
  assign P2_U2981 = ~n40269 | ~n40268;
  assign n40277 = ~P2_LWORD_REG_15__SCAN_IN | ~n40270;
  assign n40275 = ~n40226 & ~n28956;
  assign n40272 = ~n40271;
  assign n40274 = ~n40273 & ~n40272;
  assign n40276 = ~n40275 & ~n40274;
  assign P2_U2982 = ~n40277 | ~n40276;
  assign n40358 = ~n40278;
  assign n40283 = ~n40358 | ~n40324;
  assign n40280 = n40279;
  assign n40355 = ~n40281 ^ P2_INSTADDRPOINTER_REG_4__SCAN_IN;
  assign n40282 = ~n40355 | ~n40348;
  assign n40292 = ~n40283 | ~n40282;
  assign n40288 = ~n40285 & ~n40284;
  assign n40287 = ~n40286;
  assign n40290 = ~n40288 & ~n40287;
  assign n40369 = ~n40290 ^ n40289;
  assign n40291 = ~n40369 & ~n40342;
  assign n40300 = ~n40292 & ~n40291;
  assign n40298 = ~n40304 & ~n40293;
  assign n40366 = ~n40294 & ~n28339;
  assign n40296 = ~n40366;
  assign n40295 = ~n40337 | ~P2_PHYADDRPOINTER_REG_4__SCAN_IN;
  assign n40297 = ~n40296 | ~n40295;
  assign n40299 = ~n40298 & ~n40297;
  assign P2_U3010 = ~n40300 | ~n40299;
  assign n40381 = ~n40302 ^ n40301;
  assign n40314 = ~n40342 & ~n40381;
  assign n40310 = ~n40304 & ~n40303;
  assign n40307 = ~n40306 | ~n40305;
  assign n40374 = ~n40308 | ~n40307;
  assign n40309 = ~n40323 & ~n40374;
  assign n40312 = ~n40310 & ~n40309;
  assign n40311 = ~P2_PHYADDRPOINTER_REG_2__SCAN_IN | ~n40337;
  assign n40313 = ~n40312 | ~n40311;
  assign n40318 = ~n40314 & ~n40313;
  assign n40379 = ~n40325 | ~P2_REIP_REG_2__SCAN_IN;
  assign n40315 = ~n40379;
  assign n40317 = ~n40316 & ~n40315;
  assign P2_U3012 = ~n40318 | ~n40317;
  assign n40321 = ~n40320 | ~n40319;
  assign n40398 = ~n40321 ^ n42096;
  assign n40334 = ~n40342 & ~n40398;
  assign n40400 = ~n40322 ^ n42096;
  assign n40328 = ~n40323 & ~n40400;
  assign n40326 = ~n33176 | ~n40324;
  assign n40409 = ~n40325 | ~P2_REIP_REG_1__SCAN_IN;
  assign n40327 = ~n40326 | ~n40409;
  assign n40332 = ~n40328 & ~n40327;
  assign n40331 = ~n40330 | ~n40329;
  assign n40333 = ~n40332 | ~n40331;
  assign n40336 = ~n40334 & ~n40333;
  assign n40335 = ~n40337 | ~P2_PHYADDRPOINTER_REG_1__SCAN_IN;
  assign P2_U3013 = ~n40336 | ~n40335;
  assign n40339 = ~n40337;
  assign n40340 = ~n40339 | ~n40338;
  assign n40354 = ~n40340 | ~P2_PHYADDRPOINTER_REG_0__SCAN_IN;
  assign n40352 = ~n40342 & ~n40341;
  assign n40345 = ~n40344 & ~n40343;
  assign n40350 = ~n40346 & ~n40345;
  assign n40349 = ~n40348 | ~n40347;
  assign n40351 = ~n40350 | ~n40349;
  assign n40353 = ~n40352 & ~n40351;
  assign P2_U3014 = ~n40354 | ~n40353;
  assign n40364 = ~n40356 | ~n40355;
  assign n40362 = ~n40357 & ~n40399;
  assign n40359 = ~n40358 | ~n40408;
  assign n40361 = ~n40360 | ~n40359;
  assign n40363 = ~n40362 & ~n40361;
  assign n40365 = ~n40364 | ~n40363;
  assign n40373 = ~n40366 & ~n40365;
  assign n40371 = ~n40368 & ~n40367;
  assign n40370 = ~n40369 & ~n40397;
  assign n40372 = ~n40371 & ~n40370;
  assign P2_U3042 = ~n40373 | ~n40372;
  assign n40376 = ~n40399 & ~n42158;
  assign n40375 = ~n23239 & ~n40374;
  assign n40396 = ~n40376 & ~n40375;
  assign n40394 = n40378 & n40377;
  assign n40380 = ~n27757 | ~n40408;
  assign n40383 = ~n40380 | ~n40379;
  assign n40382 = ~n40397 & ~n40381;
  assign n40386 = ~n40383 & ~n40382;
  assign n40385 = ~P2_INSTADDRPOINTER_REG_2__SCAN_IN | ~n40384;
  assign n40387 = ~n40386 | ~n40385;
  assign n40392 = ~n40388 & ~n40387;
  assign n40391 = n40390 | n40389;
  assign n40393 = ~n40392 | ~n40391;
  assign n40395 = ~n40394 & ~n40393;
  assign P2_U3044 = ~n40396 | ~n40395;
  assign n40407 = ~n40398 & ~n40397;
  assign n40402 = ~n40399 & ~n42166;
  assign n40401 = ~n23239 & ~n40400;
  assign n40405 = ~n40402 & ~n40401;
  assign n40404 = ~P2_INSTADDRPOINTER_REG_1__SCAN_IN | ~n40403;
  assign n40406 = ~n40405 | ~n40404;
  assign n40416 = ~n40407 & ~n40406;
  assign n40410 = ~n33176 | ~n40408;
  assign n40414 = ~n40410 | ~n40409;
  assign n40411 = ~P2_INSTADDRPOINTER_REG_0__SCAN_IN ^ P2_INSTADDRPOINTER_REG_1__SCAN_IN;
  assign n40413 = ~n40412 & ~n40411;
  assign n40415 = ~n40414 & ~n40413;
  assign P2_U3045 = ~n40416 | ~n40415;
  assign n40448 = ~n41788 & ~n41491;
  assign n41155 = ~n42156 | ~n42112;
  assign n40417 = ~n41155;
  assign n40580 = ~n41490 | ~n40417;
  assign n40418 = ~n40448 & ~n40560;
  assign n40419 = ~n41789 & ~n40418;
  assign n40431 = ~n41002 & ~n40419;
  assign n40420 = ~n40431;
  assign n40427 = ~n40432 & ~n40420;
  assign n40424 = ~n40421 | ~n42196;
  assign n40422 = ~n40553;
  assign n40423 = ~n40422 & ~n41785;
  assign n40425 = ~n40424 | ~n40423;
  assign n40426 = ~n41686 | ~n40425;
  assign n40443 = n40546 | n40428;
  assign n41773 = ~n40429 & ~n41786;
  assign n40430 = ~n27883 | ~n40553;
  assign n40434 = ~n40430 | ~P2_STATE2_REG_2__SCAN_IN;
  assign n40433 = ~n40432 | ~n40431;
  assign n40441 = ~n41773 | ~n40566;
  assign n40439 = ~n40556 | ~BUF2_REG_16__SCAN_IN;
  assign n40438 = ~n40557 | ~BUF1_REG_16__SCAN_IN;
  assign n40440 = ~n40560 | ~n41675;
  assign n40442 = n40441 & n40440;
  assign n41775 = ~n40444 | ~n40518;
  assign n40450 = ~n41775 & ~n40553;
  assign n40447 = BUF2_REG_24__SCAN_IN & n40556;
  assign n40446 = ~n40531 & ~n40445;
  assign n41774 = ~n40447 & ~n40446;
  assign n40449 = ~n41774 & ~n41868;
  assign n40451 = ~n40450 & ~n40449;
  assign P2_U3048 = ~n23949 | ~n40451;
  assign n40464 = n40546 | n40452;
  assign n40455 = BUF2_REG_25__SCAN_IN & n40556;
  assign n40454 = ~n40453 & ~n40531;
  assign n41802 = ~n40455 & ~n40454;
  assign n40458 = ~n41802 & ~n41868;
  assign n41597 = n40456 & n40518;
  assign n40457 = ~n41796 & ~n40553;
  assign n40462 = ~n40458 & ~n40457;
  assign n40460 = ~n40556 | ~BUF2_REG_17__SCAN_IN;
  assign n40459 = ~n40557 | ~BUF1_REG_17__SCAN_IN;
  assign n40461 = ~n40560 | ~n41693;
  assign n40463 = n40462 & n40461;
  assign n41799 = ~n41690;
  assign n40466 = ~n41799 | ~n40566;
  assign P2_U3049 = ~n23965 | ~n40466;
  assign n40479 = n40546 | n40467;
  assign n40470 = ~n32032 & ~n40547;
  assign n40469 = ~n40468 & ~n40531;
  assign n41807 = ~n40470 & ~n40469;
  assign n40473 = ~n41807 & ~n41868;
  assign n40551 = ~n40518;
  assign n40472 = ~n41808 & ~n40553;
  assign n40477 = ~n40473 & ~n40472;
  assign n40475 = ~n40556 | ~BUF2_REG_18__SCAN_IN;
  assign n40474 = ~n40557 | ~BUF1_REG_18__SCAN_IN;
  assign n40476 = ~n40560 | ~n41703;
  assign n40478 = n40477 & n40476;
  assign n41811 = ~n41700;
  assign n40481 = ~n41811 | ~n40566;
  assign P2_U3050 = ~n22972 | ~n40481;
  assign n40494 = n40546 | n40482;
  assign n40485 = ~n32017 & ~n40547;
  assign n40484 = ~n40483 & ~n40531;
  assign n41826 = ~n40485 & ~n40484;
  assign n40488 = ~n41826 & ~n41868;
  assign n41820 = ~n40486 | ~n40518;
  assign n40487 = ~n41820 & ~n40553;
  assign n40492 = ~n40488 & ~n40487;
  assign n40490 = ~n40556 | ~BUF2_REG_19__SCAN_IN;
  assign n40489 = ~n40557 | ~BUF1_REG_19__SCAN_IN;
  assign n40491 = ~n40560 | ~n41710;
  assign n40493 = n40492 & n40491;
  assign n41823 = ~n41715;
  assign n40496 = ~n41823 | ~n40566;
  assign P2_U3051 = ~n22973 | ~n40496;
  assign n40509 = ~n40546 & ~n40497;
  assign n40500 = ~n32001 & ~n40547;
  assign n40499 = ~n40498 & ~n40531;
  assign n41831 = ~n40500 & ~n40499;
  assign n40503 = ~n41831 & ~n41868;
  assign n40502 = ~n41832 & ~n40553;
  assign n40507 = ~n40503 & ~n40502;
  assign n40505 = ~n40556 | ~BUF2_REG_20__SCAN_IN;
  assign n40504 = ~n40557 | ~BUF1_REG_20__SCAN_IN;
  assign n40506 = ~n40560 | ~n41720;
  assign n40508 = ~n40507 | ~n40506;
  assign n40512 = ~n40509 & ~n40508;
  assign n41725 = ~n40510 | ~n41686;
  assign n41835 = ~n41725;
  assign n40511 = ~n41835 | ~n40566;
  assign P2_U3052 = ~n40512 | ~n40511;
  assign n40527 = n40546 | n40513;
  assign n40517 = ~n40514 & ~n40531;
  assign n40516 = ~n40515 & ~n40547;
  assign n41843 = ~n40517 & ~n40516;
  assign n40521 = ~n41843 & ~n41868;
  assign n41844 = ~n40519 | ~n40518;
  assign n40520 = ~n41844 & ~n40553;
  assign n40525 = ~n40521 & ~n40520;
  assign n40523 = ~n40556 | ~BUF2_REG_21__SCAN_IN;
  assign n40522 = ~n40557 | ~BUF1_REG_21__SCAN_IN;
  assign n40524 = ~n40560 | ~n41733;
  assign n40526 = n40525 & n40524;
  assign n41730 = ~n40528 | ~n41686;
  assign n41847 = ~n41730;
  assign n40529 = ~n41847 | ~n40566;
  assign P2_U3053 = ~n22974 | ~n40529;
  assign n40542 = n40546 | n40530;
  assign n40534 = ~n40532 & ~n40531;
  assign n40533 = ~n31973 & ~n40547;
  assign n41862 = ~n40534 & ~n40533;
  assign n40536 = ~n41862 & ~n41868;
  assign n40535 = ~n41856 & ~n40553;
  assign n40540 = ~n40536 & ~n40535;
  assign n40538 = ~n40556 | ~BUF2_REG_22__SCAN_IN;
  assign n40537 = ~n40557 | ~BUF1_REG_22__SCAN_IN;
  assign n40539 = ~n40560 | ~n41740;
  assign n40541 = n40540 & n40539;
  assign n41859 = ~n41745;
  assign n40544 = ~n41859 | ~n40566;
  assign P2_U3054 = ~n22975 | ~n40544;
  assign n40564 = n40546 | n40545;
  assign n40550 = ~n40548 & ~n40547;
  assign n40549 = BUF1_REG_31__SCAN_IN & n40557;
  assign n41879 = ~n40550 & ~n40549;
  assign n40555 = ~n41879 & ~n41868;
  assign n40554 = ~n41870 & ~n40553;
  assign n40562 = ~n40555 & ~n40554;
  assign n40559 = ~n40556 | ~BUF2_REG_23__SCAN_IN;
  assign n40558 = ~n40557 | ~BUF1_REG_23__SCAN_IN;
  assign n40561 = ~n40560 | ~n41756;
  assign n40563 = n40562 & n40561;
  assign n41753 = ~n40565 | ~n41686;
  assign n41875 = ~n41753;
  assign n40567 = ~n41875 | ~n40566;
  assign P2_U3055 = ~n22976 | ~n40567;
  assign n40576 = ~n41774 & ~n40637;
  assign n40636 = ~n40582 | ~P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n40570 = ~n40568 | ~P2_STATE2_REG_2__SCAN_IN;
  assign n40569 = ~n41785 | ~n40582;
  assign n40640 = ~n40570 | ~n40569;
  assign n40574 = ~n41773 | ~n40640;
  assign n40572 = ~n41765 & ~n40729;
  assign n40571 = ~n41775 & ~n40636;
  assign n40573 = ~n40572 & ~n40571;
  assign n40575 = ~n40574 | ~n40573;
  assign n40587 = ~n40576 & ~n40575;
  assign n40578 = ~n40577 | ~n42196;
  assign n40579 = ~n40578 | ~n40636;
  assign n40584 = ~n41785 & ~n40579;
  assign n40581 = ~n41789 & ~n40580;
  assign n40583 = ~n40582 & ~n40581;
  assign n40585 = ~n40584 & ~n40583;
  assign n40586 = ~P2_INSTQUEUE_REG_1__0__SCAN_IN | ~n40645;
  assign P2_U3056 = ~n40587 | ~n40586;
  assign n40593 = ~n41796 & ~n40636;
  assign n40589 = ~n40729 & ~n41795;
  assign n40588 = ~n40637 & ~n41802;
  assign n40591 = ~n40589 & ~n40588;
  assign n40590 = ~n41799 | ~n40640;
  assign n40592 = ~n40591 | ~n40590;
  assign n40595 = ~n40593 & ~n40592;
  assign n40594 = ~P2_INSTQUEUE_REG_1__1__SCAN_IN | ~n40645;
  assign P2_U3057 = ~n40595 | ~n40594;
  assign n40601 = ~n41808 & ~n40636;
  assign n40597 = ~n40729 & ~n41814;
  assign n40596 = ~n40637 & ~n41807;
  assign n40599 = ~n40597 & ~n40596;
  assign n40598 = ~n41811 | ~n40640;
  assign n40600 = ~n40599 | ~n40598;
  assign n40603 = ~n40601 & ~n40600;
  assign n40602 = ~P2_INSTQUEUE_REG_1__2__SCAN_IN | ~n40645;
  assign P2_U3058 = ~n40603 | ~n40602;
  assign n40609 = ~n41820 & ~n40636;
  assign n40605 = ~n40729 & ~n41819;
  assign n40604 = ~n40637 & ~n41826;
  assign n40607 = ~n40605 & ~n40604;
  assign n40606 = ~n41823 | ~n40640;
  assign n40608 = ~n40607 | ~n40606;
  assign n40611 = ~n40609 & ~n40608;
  assign n40610 = ~P2_INSTQUEUE_REG_1__3__SCAN_IN | ~n40645;
  assign P2_U3059 = ~n40611 | ~n40610;
  assign n40617 = ~n41832 & ~n40636;
  assign n40613 = ~n40729 & ~n41838;
  assign n40612 = ~n40637 & ~n41831;
  assign n40615 = ~n40613 & ~n40612;
  assign n40614 = ~n41835 | ~n40640;
  assign n40616 = ~n40615 | ~n40614;
  assign n40619 = ~n40617 & ~n40616;
  assign n40618 = ~P2_INSTQUEUE_REG_1__4__SCAN_IN | ~n40645;
  assign P2_U3060 = ~n40619 | ~n40618;
  assign n40625 = ~n41844 & ~n40636;
  assign n40621 = ~n40729 & ~n41850;
  assign n40620 = ~n40637 & ~n41843;
  assign n40623 = ~n40621 & ~n40620;
  assign n40622 = ~n41847 | ~n40640;
  assign n40624 = ~n40623 | ~n40622;
  assign n40627 = ~n40625 & ~n40624;
  assign n40626 = ~P2_INSTQUEUE_REG_1__5__SCAN_IN | ~n40645;
  assign P2_U3061 = ~n40627 | ~n40626;
  assign n40633 = ~n41856 & ~n40636;
  assign n40629 = ~n40729 & ~n41855;
  assign n40628 = ~n40637 & ~n41862;
  assign n40631 = ~n40629 & ~n40628;
  assign n40630 = ~n41859 | ~n40640;
  assign n40632 = ~n40631 | ~n40630;
  assign n40635 = ~n40633 & ~n40632;
  assign n40634 = ~P2_INSTQUEUE_REG_1__6__SCAN_IN | ~n40645;
  assign P2_U3062 = ~n40635 | ~n40634;
  assign n40644 = ~n41870 & ~n40636;
  assign n40639 = ~n40729 & ~n41867;
  assign n40638 = ~n40637 & ~n41879;
  assign n40642 = ~n40639 & ~n40638;
  assign n40641 = ~n41875 | ~n40640;
  assign n40643 = ~n40642 | ~n40641;
  assign n40647 = ~n40644 & ~n40643;
  assign n40646 = ~P2_INSTQUEUE_REG_1__7__SCAN_IN | ~n40645;
  assign P2_U3063 = ~n40647 | ~n40646;
  assign n40671 = ~n41774 & ~n40729;
  assign n40723 = ~n40746 | ~n41575;
  assign n40656 = ~n41775 & ~n40723;
  assign n40650 = ~n40992;
  assign n40649 = ~n41785 | ~n40648;
  assign n40662 = ~n40650 & ~n40649;
  assign n40652 = ~n40657;
  assign n40651 = ~n40723;
  assign n40653 = ~n40652 & ~n40651;
  assign n40654 = ~n40653 & ~n41664;
  assign n40655 = ~n40722 & ~n41672;
  assign n40669 = ~n40656 & ~n40655;
  assign n40658 = ~n40657 | ~P2_STATE2_REG_2__SCAN_IN;
  assign n40659 = ~n40658 | ~n42196;
  assign n40667 = ~n40659 | ~n40723;
  assign n40660 = ~n40729;
  assign n40661 = ~n40740 & ~n40660;
  assign n40664 = ~n41789 & ~n40661;
  assign n40663 = n40662 | n41002;
  assign n40665 = ~n40664 & ~n40663;
  assign n40666 = ~n41786 & ~n40665;
  assign n40726 = ~n40667 | ~n40666;
  assign n40668 = ~P2_INSTQUEUE_REG_2__0__SCAN_IN | ~n40726;
  assign n40670 = ~n40669 | ~n40668;
  assign n40673 = ~n40671 & ~n40670;
  assign n40672 = ~n40740 | ~n41675;
  assign P2_U3064 = ~n40673 | ~n40672;
  assign n40675 = ~n41690 & ~n40722;
  assign n40674 = ~n41796 & ~n40723;
  assign n40681 = ~n40675 & ~n40674;
  assign n40677 = ~P2_INSTQUEUE_REG_2__1__SCAN_IN | ~n40726;
  assign n40676 = ~n40740 | ~n41693;
  assign n40679 = ~n40677 | ~n40676;
  assign n40678 = ~n41802 & ~n40729;
  assign n40680 = ~n40679 & ~n40678;
  assign P2_U3065 = ~n40681 | ~n40680;
  assign n40683 = ~n41700 & ~n40722;
  assign n40682 = ~n41808 & ~n40723;
  assign n40689 = ~n40683 & ~n40682;
  assign n40685 = ~P2_INSTQUEUE_REG_2__2__SCAN_IN | ~n40726;
  assign n40684 = ~n40740 | ~n41703;
  assign n40687 = ~n40685 | ~n40684;
  assign n40686 = ~n41807 & ~n40729;
  assign n40688 = ~n40687 & ~n40686;
  assign P2_U3066 = ~n40689 | ~n40688;
  assign n40691 = ~n41715 & ~n40722;
  assign n40690 = ~n41820 & ~n40723;
  assign n40697 = ~n40691 & ~n40690;
  assign n40693 = ~P2_INSTQUEUE_REG_2__3__SCAN_IN | ~n40726;
  assign n40692 = ~n40740 | ~n41710;
  assign n40695 = ~n40693 | ~n40692;
  assign n40694 = ~n41826 & ~n40729;
  assign n40696 = ~n40695 & ~n40694;
  assign P2_U3067 = ~n40697 | ~n40696;
  assign n40699 = ~n41725 & ~n40722;
  assign n40698 = ~n41832 & ~n40723;
  assign n40705 = ~n40699 & ~n40698;
  assign n40701 = ~P2_INSTQUEUE_REG_2__4__SCAN_IN | ~n40726;
  assign n40700 = ~n40740 | ~n41720;
  assign n40703 = ~n40701 | ~n40700;
  assign n40702 = ~n41831 & ~n40729;
  assign n40704 = ~n40703 & ~n40702;
  assign P2_U3068 = ~n40705 | ~n40704;
  assign n40707 = ~n41730 & ~n40722;
  assign n40706 = ~n41844 & ~n40723;
  assign n40713 = ~n40707 & ~n40706;
  assign n40709 = ~P2_INSTQUEUE_REG_2__5__SCAN_IN | ~n40726;
  assign n40708 = ~n40740 | ~n41733;
  assign n40711 = ~n40709 | ~n40708;
  assign n40710 = ~n41843 & ~n40729;
  assign n40712 = ~n40711 & ~n40710;
  assign P2_U3069 = ~n40713 | ~n40712;
  assign n40715 = ~n41745 & ~n40722;
  assign n40714 = ~n41856 & ~n40723;
  assign n40721 = ~n40715 & ~n40714;
  assign n40717 = ~P2_INSTQUEUE_REG_2__6__SCAN_IN | ~n40726;
  assign n40716 = ~n40740 | ~n41740;
  assign n40719 = ~n40717 | ~n40716;
  assign n40718 = ~n41862 & ~n40729;
  assign n40720 = ~n40719 & ~n40718;
  assign P2_U3070 = ~n40721 | ~n40720;
  assign n40725 = ~n41753 & ~n40722;
  assign n40724 = ~n41870 & ~n40723;
  assign n40733 = ~n40725 & ~n40724;
  assign n40728 = ~P2_INSTQUEUE_REG_2__7__SCAN_IN | ~n40726;
  assign n40727 = ~n40740 | ~n41756;
  assign n40731 = ~n40728 | ~n40727;
  assign n40730 = ~n41879 & ~n40729;
  assign n40732 = ~n40731 & ~n40730;
  assign P2_U3071 = ~n40733 | ~n40732;
  assign n40735 = ~n23291 & ~n40741;
  assign n40739 = ~n40735 & ~n41664;
  assign n40737 = ~n40746;
  assign n40736 = ~P2_STATEBS16_REG_SCAN_IN | ~n40755;
  assign n40747 = ~n41785 | ~n40736;
  assign n40738 = ~n40737 & ~n40747;
  assign n40754 = ~n40808 & ~n41672;
  assign n40743 = ~n40807 & ~n41774;
  assign n40742 = ~n41775 & ~n40806;
  assign n40752 = ~n40743 & ~n40742;
  assign n40744 = ~n23291 | ~n42196;
  assign n40745 = ~n40744 | ~n40806;
  assign n40749 = ~n41785 & ~n40745;
  assign n40748 = ~n40747 & ~n40746;
  assign n40750 = ~n40749 & ~n40748;
  assign n40815 = ~n40750 | ~n41686;
  assign n40751 = ~P2_INSTQUEUE_REG_3__0__SCAN_IN | ~n40815;
  assign n40753 = ~n40752 | ~n40751;
  assign n40757 = ~n40754 & ~n40753;
  assign n40756 = ~n40820 | ~n41675;
  assign P2_U3072 = ~n40757 | ~n40756;
  assign n40761 = ~n41796 & ~n40806;
  assign n40759 = ~P2_INSTQUEUE_REG_3__1__SCAN_IN | ~n40815;
  assign n40758 = ~n40820 | ~n41693;
  assign n40760 = ~n40759 | ~n40758;
  assign n40765 = ~n40761 & ~n40760;
  assign n40763 = ~n40807 & ~n41802;
  assign n40762 = ~n41690 & ~n40808;
  assign n40764 = ~n40763 & ~n40762;
  assign P2_U3073 = ~n40765 | ~n40764;
  assign n40767 = ~n40807 & ~n41807;
  assign n40766 = ~n41808 & ~n40806;
  assign n40773 = ~n40767 & ~n40766;
  assign n40769 = ~P2_INSTQUEUE_REG_3__2__SCAN_IN | ~n40815;
  assign n40768 = ~n40820 | ~n41703;
  assign n40771 = ~n40769 | ~n40768;
  assign n40770 = ~n40808 & ~n41700;
  assign n40772 = ~n40771 & ~n40770;
  assign P2_U3074 = ~n40773 | ~n40772;
  assign n40777 = ~n41820 & ~n40806;
  assign n40775 = ~P2_INSTQUEUE_REG_3__3__SCAN_IN | ~n40815;
  assign n40774 = ~n40820 | ~n41710;
  assign n40776 = ~n40775 | ~n40774;
  assign n40781 = ~n40777 & ~n40776;
  assign n40779 = ~n40807 & ~n41826;
  assign n40778 = ~n41715 & ~n40808;
  assign n40780 = ~n40779 & ~n40778;
  assign P2_U3075 = ~n40781 | ~n40780;
  assign n40783 = ~n40807 & ~n41831;
  assign n40782 = ~n41832 & ~n40806;
  assign n40789 = ~n40783 & ~n40782;
  assign n40785 = ~P2_INSTQUEUE_REG_3__4__SCAN_IN | ~n40815;
  assign n40784 = ~n40820 | ~n41720;
  assign n40787 = ~n40785 | ~n40784;
  assign n40786 = ~n40808 & ~n41725;
  assign n40788 = ~n40787 & ~n40786;
  assign P2_U3076 = ~n40789 | ~n40788;
  assign n40793 = ~n41844 & ~n40806;
  assign n40791 = ~P2_INSTQUEUE_REG_3__5__SCAN_IN | ~n40815;
  assign n40790 = ~n40820 | ~n41733;
  assign n40792 = ~n40791 | ~n40790;
  assign n40797 = ~n40793 & ~n40792;
  assign n40795 = ~n40807 & ~n41843;
  assign n40794 = ~n41730 & ~n40808;
  assign n40796 = ~n40795 & ~n40794;
  assign P2_U3077 = ~n40797 | ~n40796;
  assign n40803 = ~n41856 & ~n40806;
  assign n40799 = ~n40807 & ~n41862;
  assign n40798 = ~n41745 & ~n40808;
  assign n40801 = ~n40799 & ~n40798;
  assign n40800 = ~n40820 | ~n41740;
  assign n40802 = ~n40801 | ~n40800;
  assign n40805 = ~n40803 & ~n40802;
  assign n40804 = ~P2_INSTQUEUE_REG_3__6__SCAN_IN | ~n40815;
  assign P2_U3078 = ~n40805 | ~n40804;
  assign n40814 = ~n41870 & ~n40806;
  assign n40810 = ~n40807 & ~n41879;
  assign n40809 = ~n41753 & ~n40808;
  assign n40812 = ~n40810 & ~n40809;
  assign n40811 = ~n40820 | ~n41756;
  assign n40813 = ~n40812 | ~n40811;
  assign n40817 = ~n40814 & ~n40813;
  assign n40816 = ~P2_INSTQUEUE_REG_3__7__SCAN_IN | ~n40815;
  assign P2_U3079 = ~n40817 | ~n40816;
  assign n40834 = ~n41774 & ~n40894;
  assign n40838 = n40922 & n41575;
  assign n40895 = ~n40838;
  assign n40830 = ~n41775 & ~n40895;
  assign n40835 = ~n27905;
  assign n40818 = ~n40835 & ~n40838;
  assign n40828 = ~n40818 & ~n41664;
  assign n40819 = ~n41489;
  assign n40913 = ~n41490 | ~n40819;
  assign n40977 = n40913 | n42177;
  assign n40899 = ~n40977;
  assign n40821 = ~n40899 & ~n40820;
  assign n40822 = ~n41789 & ~n40821;
  assign n40841 = ~n41002 & ~n40822;
  assign n40826 = ~n40841;
  assign n40825 = ~n41493;
  assign n40824 = ~n40823;
  assign n41494 = ~n40824 & ~n40992;
  assign n40840 = ~n40825 | ~n41494;
  assign n40827 = ~n40826 & ~n40840;
  assign n40896 = ~n40828 & ~n40827;
  assign n40829 = ~n40896 & ~n41672;
  assign n40832 = ~n40830 & ~n40829;
  assign n40831 = ~n40899 | ~n41675;
  assign n40833 = ~n40832 | ~n40831;
  assign n40845 = ~n40834 & ~n40833;
  assign n40836 = ~n40835 | ~n42196;
  assign n40837 = ~n40836 | ~n41002;
  assign n40839 = ~n40838 & ~n40837;
  assign n40843 = ~n41786 & ~n40839;
  assign n40842 = ~n40841 | ~n40840;
  assign n40844 = ~P2_INSTQUEUE_REG_4__0__SCAN_IN | ~n40904;
  assign P2_U3080 = ~n40845 | ~n40844;
  assign n40851 = ~n41802 & ~n40894;
  assign n40847 = ~n41796 & ~n40895;
  assign n40846 = ~n40896 & ~n41690;
  assign n40849 = ~n40847 & ~n40846;
  assign n40848 = ~n40899 | ~n41693;
  assign n40850 = ~n40849 | ~n40848;
  assign n40853 = ~n40851 & ~n40850;
  assign n40852 = ~P2_INSTQUEUE_REG_4__1__SCAN_IN | ~n40904;
  assign P2_U3081 = ~n40853 | ~n40852;
  assign n40855 = ~n40894 & ~n41807;
  assign n40854 = ~n41808 & ~n40895;
  assign n40861 = ~n40855 & ~n40854;
  assign n40857 = ~P2_INSTQUEUE_REG_4__2__SCAN_IN | ~n40904;
  assign n40856 = ~n40899 | ~n41703;
  assign n40859 = ~n40857 | ~n40856;
  assign n40858 = ~n40896 & ~n41700;
  assign n40860 = ~n40859 & ~n40858;
  assign P2_U3082 = ~n40861 | ~n40860;
  assign n40863 = ~n40894 & ~n41826;
  assign n40862 = ~n41820 & ~n40895;
  assign n40869 = ~n40863 & ~n40862;
  assign n40865 = ~P2_INSTQUEUE_REG_4__3__SCAN_IN | ~n40904;
  assign n40864 = ~n40899 | ~n41710;
  assign n40867 = ~n40865 | ~n40864;
  assign n40866 = ~n40896 & ~n41715;
  assign n40868 = ~n40867 & ~n40866;
  assign P2_U3083 = ~n40869 | ~n40868;
  assign n40875 = ~n41831 & ~n40894;
  assign n40871 = ~n41832 & ~n40895;
  assign n40870 = ~n40896 & ~n41725;
  assign n40873 = ~n40871 & ~n40870;
  assign n40872 = ~n40899 | ~n41720;
  assign n40874 = ~n40873 | ~n40872;
  assign n40877 = ~n40875 & ~n40874;
  assign n40876 = ~P2_INSTQUEUE_REG_4__4__SCAN_IN | ~n40904;
  assign P2_U3084 = ~n40877 | ~n40876;
  assign n40883 = ~n41843 & ~n40894;
  assign n40879 = ~n41844 & ~n40895;
  assign n40878 = ~n40896 & ~n41730;
  assign n40881 = ~n40879 & ~n40878;
  assign n40880 = ~n40899 | ~n41733;
  assign n40882 = ~n40881 | ~n40880;
  assign n40885 = ~n40883 & ~n40882;
  assign n40884 = ~P2_INSTQUEUE_REG_4__5__SCAN_IN | ~n40904;
  assign P2_U3085 = ~n40885 | ~n40884;
  assign n40887 = ~n40894 & ~n41862;
  assign n40886 = ~n41856 & ~n40895;
  assign n40893 = ~n40887 & ~n40886;
  assign n40889 = ~P2_INSTQUEUE_REG_4__6__SCAN_IN | ~n40904;
  assign n40888 = ~n40899 | ~n41740;
  assign n40891 = ~n40889 | ~n40888;
  assign n40890 = ~n40896 & ~n41745;
  assign n40892 = ~n40891 & ~n40890;
  assign P2_U3086 = ~n40893 | ~n40892;
  assign n40903 = ~n41879 & ~n40894;
  assign n40898 = ~n41870 & ~n40895;
  assign n40897 = ~n40896 & ~n41753;
  assign n40901 = ~n40898 & ~n40897;
  assign n40900 = ~n40899 | ~n41756;
  assign n40902 = ~n40901 | ~n40900;
  assign n40906 = ~n40903 & ~n40902;
  assign n40905 = ~P2_INSTQUEUE_REG_4__7__SCAN_IN | ~n40904;
  assign P2_U3087 = ~n40906 | ~n40905;
  assign n40917 = ~n41774 & ~n40977;
  assign n40978 = ~n40920;
  assign n40912 = ~n41775 & ~n40978;
  assign n40907 = ~n27869 & ~n40920;
  assign n40910 = ~n40907 & ~n41664;
  assign n40908 = ~n41789 & ~n40913;
  assign n40923 = ~n41002 & ~n40908;
  assign n40909 = n40923 & n40922;
  assign n40911 = ~n40985 & ~n41672;
  assign n40915 = ~n40912 & ~n40911;
  assign n40914 = ~n40982 | ~n41675;
  assign n40916 = ~n40915 | ~n40914;
  assign n40928 = ~n40917 & ~n40916;
  assign n40918 = ~n27869 | ~n42196;
  assign n40919 = ~n40918 | ~n41002;
  assign n40921 = ~n40920 & ~n40919;
  assign n40926 = ~n41786 & ~n40921;
  assign n40924 = ~n40922;
  assign n40925 = ~n40924 | ~n40923;
  assign n40927 = ~P2_INSTQUEUE_REG_5__0__SCAN_IN | ~n40981;
  assign P2_U3088 = ~n40928 | ~n40927;
  assign n40930 = ~n40977 & ~n41802;
  assign n40929 = ~n41796 & ~n40978;
  assign n40936 = ~n40930 & ~n40929;
  assign n40932 = ~P2_INSTQUEUE_REG_5__1__SCAN_IN | ~n40981;
  assign n40931 = ~n40982 | ~n41693;
  assign n40934 = ~n40932 | ~n40931;
  assign n40933 = ~n40985 & ~n41690;
  assign n40935 = ~n40934 & ~n40933;
  assign P2_U3089 = ~n40936 | ~n40935;
  assign n40942 = ~n41808 & ~n40978;
  assign n40938 = ~n40977 & ~n41807;
  assign n40937 = ~n41700 & ~n40985;
  assign n40940 = ~n40938 & ~n40937;
  assign n40939 = ~n40982 | ~n41703;
  assign n40941 = ~n40940 | ~n40939;
  assign n40944 = ~n40942 & ~n40941;
  assign n40943 = ~P2_INSTQUEUE_REG_5__2__SCAN_IN | ~n40981;
  assign P2_U3090 = ~n40944 | ~n40943;
  assign n40946 = ~n40977 & ~n41826;
  assign n40945 = ~n41820 & ~n40978;
  assign n40952 = ~n40946 & ~n40945;
  assign n40948 = ~P2_INSTQUEUE_REG_5__3__SCAN_IN | ~n40981;
  assign n40947 = ~n40982 | ~n41710;
  assign n40950 = ~n40948 | ~n40947;
  assign n40949 = ~n40985 & ~n41715;
  assign n40951 = ~n40950 & ~n40949;
  assign P2_U3091 = ~n40952 | ~n40951;
  assign n40954 = ~n40977 & ~n41831;
  assign n40953 = ~n41832 & ~n40978;
  assign n40960 = ~n40954 & ~n40953;
  assign n40956 = ~P2_INSTQUEUE_REG_5__4__SCAN_IN | ~n40981;
  assign n40955 = ~n40982 | ~n41720;
  assign n40958 = ~n40956 | ~n40955;
  assign n40957 = ~n40985 & ~n41725;
  assign n40959 = ~n40958 & ~n40957;
  assign P2_U3092 = ~n40960 | ~n40959;
  assign n40962 = ~n40977 & ~n41843;
  assign n40961 = ~n41844 & ~n40978;
  assign n40968 = ~n40962 & ~n40961;
  assign n40964 = ~P2_INSTQUEUE_REG_5__5__SCAN_IN | ~n40981;
  assign n40963 = ~n40982 | ~n41733;
  assign n40966 = ~n40964 | ~n40963;
  assign n40965 = ~n40985 & ~n41730;
  assign n40967 = ~n40966 & ~n40965;
  assign P2_U3093 = ~n40968 | ~n40967;
  assign n40970 = ~n40977 & ~n41862;
  assign n40969 = ~n41856 & ~n40978;
  assign n40976 = ~n40970 & ~n40969;
  assign n40972 = ~P2_INSTQUEUE_REG_5__6__SCAN_IN | ~n40981;
  assign n40971 = ~n40982 | ~n41740;
  assign n40974 = ~n40972 | ~n40971;
  assign n40973 = ~n40985 & ~n41745;
  assign n40975 = ~n40974 & ~n40973;
  assign P2_U3094 = ~n40976 | ~n40975;
  assign n40980 = ~n40977 & ~n41879;
  assign n40979 = ~n41870 & ~n40978;
  assign n40989 = ~n40980 & ~n40979;
  assign n40984 = ~P2_INSTQUEUE_REG_5__7__SCAN_IN | ~n40981;
  assign n40983 = ~n40982 | ~n41756;
  assign n40987 = ~n40984 | ~n40983;
  assign n40986 = ~n40985 & ~n41753;
  assign n40988 = ~n40987 & ~n40986;
  assign P2_U3095 = ~n40989 | ~n40988;
  assign n41012 = ~n41774 & ~n41071;
  assign n41005 = ~n41089 & ~P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n41064 = ~n41005;
  assign n40996 = ~n41775 & ~n41064;
  assign n41001 = ~n27904;
  assign n40990 = ~n41001 & ~n41005;
  assign n40994 = ~n40990 & ~n41664;
  assign n40999 = ~n40992 | ~n40991;
  assign n40993 = ~n40999 & ~n41002;
  assign n40995 = ~n41063 & ~n41672;
  assign n41010 = ~n40996 & ~n40995;
  assign n40997 = ~n42140;
  assign n40998 = ~n41071 | ~n41144;
  assign n41000 = ~n40998 | ~P2_STATEBS16_REG_SCAN_IN;
  assign n41008 = ~n41000 | ~n40999;
  assign n41003 = ~n41001 | ~n42196;
  assign n41004 = ~n41003 | ~n41002;
  assign n41006 = ~n41005 & ~n41004;
  assign n41007 = ~n41006 & ~n41786;
  assign n41067 = ~n41008 | ~n41007;
  assign n41009 = ~P2_INSTQUEUE_REG_6__0__SCAN_IN | ~n41067;
  assign n41011 = ~n41010 | ~n41009;
  assign n41014 = ~n41012 & ~n41011;
  assign n41013 = ~n41068 | ~n41675;
  assign P2_U3096 = ~n41014 | ~n41013;
  assign n41016 = ~n41690 & ~n41063;
  assign n41015 = ~n41796 & ~n41064;
  assign n41022 = ~n41016 & ~n41015;
  assign n41018 = ~P2_INSTQUEUE_REG_6__1__SCAN_IN | ~n41067;
  assign n41017 = ~n41068 | ~n41693;
  assign n41020 = ~n41018 | ~n41017;
  assign n41019 = ~n41802 & ~n41071;
  assign n41021 = ~n41020 & ~n41019;
  assign P2_U3097 = ~n41022 | ~n41021;
  assign n41024 = ~n41700 & ~n41063;
  assign n41023 = ~n41808 & ~n41064;
  assign n41030 = ~n41024 & ~n41023;
  assign n41026 = ~P2_INSTQUEUE_REG_6__2__SCAN_IN | ~n41067;
  assign n41025 = ~n41068 | ~n41703;
  assign n41028 = ~n41026 | ~n41025;
  assign n41027 = ~n41807 & ~n41071;
  assign n41029 = ~n41028 & ~n41027;
  assign P2_U3098 = ~n41030 | ~n41029;
  assign n41032 = ~n41715 & ~n41063;
  assign n41031 = ~n41820 & ~n41064;
  assign n41038 = ~n41032 & ~n41031;
  assign n41034 = ~P2_INSTQUEUE_REG_6__3__SCAN_IN | ~n41067;
  assign n41033 = ~n41068 | ~n41710;
  assign n41036 = ~n41034 | ~n41033;
  assign n41035 = ~n41826 & ~n41071;
  assign n41037 = ~n41036 & ~n41035;
  assign P2_U3099 = ~n41038 | ~n41037;
  assign n41040 = ~n41725 & ~n41063;
  assign n41039 = ~n41832 & ~n41064;
  assign n41046 = ~n41040 & ~n41039;
  assign n41042 = ~P2_INSTQUEUE_REG_6__4__SCAN_IN | ~n41067;
  assign n41041 = ~n41068 | ~n41720;
  assign n41044 = ~n41042 | ~n41041;
  assign n41043 = ~n41831 & ~n41071;
  assign n41045 = ~n41044 & ~n41043;
  assign P2_U3100 = ~n41046 | ~n41045;
  assign n41048 = ~n41730 & ~n41063;
  assign n41047 = ~n41844 & ~n41064;
  assign n41054 = ~n41048 & ~n41047;
  assign n41050 = ~P2_INSTQUEUE_REG_6__5__SCAN_IN | ~n41067;
  assign n41049 = ~n41068 | ~n41733;
  assign n41052 = ~n41050 | ~n41049;
  assign n41051 = ~n41843 & ~n41071;
  assign n41053 = ~n41052 & ~n41051;
  assign P2_U3101 = ~n41054 | ~n41053;
  assign n41056 = ~n41745 & ~n41063;
  assign n41055 = ~n41856 & ~n41064;
  assign n41062 = ~n41056 & ~n41055;
  assign n41058 = ~P2_INSTQUEUE_REG_6__6__SCAN_IN | ~n41067;
  assign n41057 = ~n41068 | ~n41740;
  assign n41060 = ~n41058 | ~n41057;
  assign n41059 = ~n41862 & ~n41071;
  assign n41061 = ~n41060 & ~n41059;
  assign P2_U3102 = ~n41062 | ~n41061;
  assign n41066 = ~n41753 & ~n41063;
  assign n41065 = ~n41870 & ~n41064;
  assign n41075 = ~n41066 & ~n41065;
  assign n41070 = ~P2_INSTQUEUE_REG_6__7__SCAN_IN | ~n41067;
  assign n41069 = ~n41068 | ~n41756;
  assign n41073 = ~n41070 | ~n41069;
  assign n41072 = ~n41879 & ~n41071;
  assign n41074 = ~n41073 & ~n41072;
  assign P2_U3103 = ~n41075 | ~n41074;
  assign n41085 = ~n27897;
  assign n41076 = ~n41085 & ~n41158;
  assign n41078 = ~n41076 & ~n41664;
  assign n41077 = ~n41089 & ~n41002;
  assign n41084 = ~n41143 & ~n41672;
  assign n41080 = ~n41228 & ~n41765;
  assign n41079 = ~n41144 & ~n41774;
  assign n41082 = ~n41080 & ~n41079;
  assign n41579 = ~n41775;
  assign n41081 = ~n41579 | ~n41158;
  assign n41083 = ~n41082 | ~n41081;
  assign n41094 = ~n41084 & ~n41083;
  assign n41086 = ~n41085 | ~n42196;
  assign n41087 = ~n41086 | ~n41002;
  assign n41088 = ~n41158 & ~n41087;
  assign n41092 = ~n41088 & ~n41786;
  assign n41090 = ~P2_STATEBS16_REG_SCAN_IN | ~n42139;
  assign n41091 = ~n41090 | ~n41089;
  assign n41093 = ~P2_INSTQUEUE_REG_7__0__SCAN_IN | ~n41151;
  assign P2_U3104 = ~n41094 | ~n41093;
  assign n41100 = ~n41143 & ~n41690;
  assign n41096 = ~n41228 & ~n41795;
  assign n41095 = ~n41144 & ~n41802;
  assign n41098 = ~n41096 & ~n41095;
  assign n41097 = ~n41597 | ~n41158;
  assign n41099 = ~n41098 | ~n41097;
  assign n41102 = ~n41100 & ~n41099;
  assign n41101 = ~P2_INSTQUEUE_REG_7__1__SCAN_IN | ~n41151;
  assign P2_U3105 = ~n41102 | ~n41101;
  assign n41108 = ~n41143 & ~n41700;
  assign n41104 = ~n41228 & ~n41814;
  assign n41103 = ~n41144 & ~n41807;
  assign n41106 = ~n41104 & ~n41103;
  assign n41105 = ~n41606 | ~n41158;
  assign n41107 = ~n41106 | ~n41105;
  assign n41110 = ~n41108 & ~n41107;
  assign n41109 = ~P2_INSTQUEUE_REG_7__2__SCAN_IN | ~n41151;
  assign P2_U3106 = ~n41110 | ~n41109;
  assign n41116 = ~n41143 & ~n41715;
  assign n41112 = ~n41228 & ~n41819;
  assign n41111 = ~n41144 & ~n41826;
  assign n41114 = ~n41112 & ~n41111;
  assign n41615 = ~n41820;
  assign n41113 = ~n41615 | ~n41158;
  assign n41115 = ~n41114 | ~n41113;
  assign n41118 = ~n41116 & ~n41115;
  assign n41117 = ~P2_INSTQUEUE_REG_7__3__SCAN_IN | ~n41151;
  assign P2_U3107 = ~n41118 | ~n41117;
  assign n41124 = ~n41143 & ~n41725;
  assign n41120 = ~n41228 & ~n41838;
  assign n41119 = ~n41144 & ~n41831;
  assign n41122 = ~n41120 & ~n41119;
  assign n41121 = ~n41624 | ~n41158;
  assign n41123 = ~n41122 | ~n41121;
  assign n41126 = ~n41124 & ~n41123;
  assign n41125 = ~P2_INSTQUEUE_REG_7__4__SCAN_IN | ~n41151;
  assign P2_U3108 = ~n41126 | ~n41125;
  assign n41132 = ~n41143 & ~n41730;
  assign n41128 = ~n41228 & ~n41850;
  assign n41127 = ~n41144 & ~n41843;
  assign n41130 = ~n41128 & ~n41127;
  assign n41633 = ~n41844;
  assign n41129 = ~n41633 | ~n41158;
  assign n41131 = ~n41130 | ~n41129;
  assign n41134 = ~n41132 & ~n41131;
  assign n41133 = ~P2_INSTQUEUE_REG_7__5__SCAN_IN | ~n41151;
  assign P2_U3109 = ~n41134 | ~n41133;
  assign n41140 = ~n41143 & ~n41745;
  assign n41136 = ~n41228 & ~n41855;
  assign n41135 = ~n41144 & ~n41862;
  assign n41138 = ~n41136 & ~n41135;
  assign n41137 = ~n41642 | ~n41158;
  assign n41139 = ~n41138 | ~n41137;
  assign n41142 = ~n41140 & ~n41139;
  assign n41141 = ~P2_INSTQUEUE_REG_7__6__SCAN_IN | ~n41151;
  assign P2_U3110 = ~n41142 | ~n41141;
  assign n41150 = ~n41143 & ~n41753;
  assign n41146 = ~n41228 & ~n41867;
  assign n41145 = ~n41144 & ~n41879;
  assign n41148 = ~n41146 & ~n41145;
  assign n41652 = ~n41870;
  assign n41147 = ~n41652 | ~n41158;
  assign n41149 = ~n41148 | ~n41147;
  assign n41153 = ~n41150 & ~n41149;
  assign n41152 = ~P2_INSTQUEUE_REG_7__7__SCAN_IN | ~n41151;
  assign P2_U3111 = ~n41153 | ~n41152;
  assign n41167 = ~n41774 & ~n41228;
  assign n41154 = ~P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN & ~P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN;
  assign n41172 = n41255 & n41575;
  assign n41163 = ~n41775 & ~n41227;
  assign n41232 = ~n41242 & ~n42177;
  assign n41156 = ~n41310 | ~n41228;
  assign n41157 = ~n41156 | ~P2_STATEBS16_REG_SCAN_IN;
  assign n41170 = ~n41157 | ~n41785;
  assign n41168 = ~n41158 & ~n41172;
  assign n41161 = ~n41170 & ~n41168;
  assign n41159 = ~n27881 & ~n41172;
  assign n41160 = ~n41159 & ~n41664;
  assign n41229 = ~n41161 & ~n41160;
  assign n41162 = ~n41229 & ~n41672;
  assign n41165 = ~n41163 & ~n41162;
  assign n41164 = ~n41232 | ~n41675;
  assign n41166 = ~n41165 | ~n41164;
  assign n41178 = ~n41167 & ~n41166;
  assign n41169 = ~n41168;
  assign n41171 = ~n41170 & ~n41169;
  assign n41176 = ~n41171 & ~n41786;
  assign n41173 = ~n23107 & ~P2_STATE2_REG_3__SCAN_IN;
  assign n41174 = ~n41173 & ~n41172;
  assign n41175 = ~n41174 | ~n41002;
  assign n41177 = ~P2_INSTQUEUE_REG_8__0__SCAN_IN | ~n41237;
  assign P2_U3112 = ~n41178 | ~n41177;
  assign n41182 = ~n41796 & ~n41227;
  assign n41180 = ~P2_INSTQUEUE_REG_8__1__SCAN_IN | ~n41237;
  assign n41179 = ~n41232 | ~n41693;
  assign n41181 = ~n41180 | ~n41179;
  assign n41186 = ~n41182 & ~n41181;
  assign n41184 = ~n41228 & ~n41802;
  assign n41183 = ~n41690 & ~n41229;
  assign n41185 = ~n41184 & ~n41183;
  assign P2_U3113 = ~n41186 | ~n41185;
  assign n41190 = ~n41808 & ~n41227;
  assign n41188 = ~P2_INSTQUEUE_REG_8__2__SCAN_IN | ~n41237;
  assign n41187 = ~n41232 | ~n41703;
  assign n41189 = ~n41188 | ~n41187;
  assign n41194 = ~n41190 & ~n41189;
  assign n41192 = ~n41228 & ~n41807;
  assign n41191 = ~n41700 & ~n41229;
  assign n41193 = ~n41192 & ~n41191;
  assign P2_U3114 = ~n41194 | ~n41193;
  assign n41198 = ~n41820 & ~n41227;
  assign n41196 = ~P2_INSTQUEUE_REG_8__3__SCAN_IN | ~n41237;
  assign n41195 = ~n41232 | ~n41710;
  assign n41197 = ~n41196 | ~n41195;
  assign n41202 = ~n41198 & ~n41197;
  assign n41200 = ~n41228 & ~n41826;
  assign n41199 = ~n41715 & ~n41229;
  assign n41201 = ~n41200 & ~n41199;
  assign P2_U3115 = ~n41202 | ~n41201;
  assign n41208 = ~n41832 & ~n41227;
  assign n41204 = ~n41228 & ~n41831;
  assign n41203 = ~n41725 & ~n41229;
  assign n41206 = ~n41204 & ~n41203;
  assign n41205 = ~n41232 | ~n41720;
  assign n41207 = ~n41206 | ~n41205;
  assign n41210 = ~n41208 & ~n41207;
  assign n41209 = ~P2_INSTQUEUE_REG_8__4__SCAN_IN | ~n41237;
  assign P2_U3116 = ~n41210 | ~n41209;
  assign n41216 = ~n41844 & ~n41227;
  assign n41212 = ~n41228 & ~n41843;
  assign n41211 = ~n41730 & ~n41229;
  assign n41214 = ~n41212 & ~n41211;
  assign n41213 = ~n41232 | ~n41733;
  assign n41215 = ~n41214 | ~n41213;
  assign n41218 = ~n41216 & ~n41215;
  assign n41217 = ~P2_INSTQUEUE_REG_8__5__SCAN_IN | ~n41237;
  assign P2_U3117 = ~n41218 | ~n41217;
  assign n41224 = ~n41856 & ~n41227;
  assign n41220 = ~n41228 & ~n41862;
  assign n41219 = ~n41745 & ~n41229;
  assign n41222 = ~n41220 & ~n41219;
  assign n41221 = ~n41232 | ~n41740;
  assign n41223 = ~n41222 | ~n41221;
  assign n41226 = ~n41224 & ~n41223;
  assign n41225 = ~P2_INSTQUEUE_REG_8__6__SCAN_IN | ~n41237;
  assign P2_U3118 = ~n41226 | ~n41225;
  assign n41236 = ~n41870 & ~n41227;
  assign n41231 = ~n41228 & ~n41879;
  assign n41230 = ~n41753 & ~n41229;
  assign n41234 = ~n41231 & ~n41230;
  assign n41233 = ~n41232 | ~n41756;
  assign n41235 = ~n41234 | ~n41233;
  assign n41239 = ~n41236 & ~n41235;
  assign n41238 = ~P2_INSTQUEUE_REG_8__7__SCAN_IN | ~n41237;
  assign P2_U3119 = ~n41239 | ~n41238;
  assign n41240 = ~n41242;
  assign n41395 = ~n41240 | ~n42177;
  assign n41251 = ~n41765 & ~n41395;
  assign n41249 = ~n41579 | ~n41326;
  assign n41241 = ~n27956 & ~n41326;
  assign n41245 = ~n41241 & ~n41664;
  assign n41243 = ~n41789 & ~n41242;
  assign n41257 = ~n41002 & ~n41243;
  assign n41244 = n41257 & n41255;
  assign n41247 = ~n41311 & ~n41672;
  assign n41246 = ~n41774 & ~n41310;
  assign n41248 = ~n41247 & ~n41246;
  assign n41250 = ~n41249 | ~n41248;
  assign n41261 = ~n41251 & ~n41250;
  assign n41252 = ~n27956 | ~n42196;
  assign n41253 = ~n41252 | ~n41002;
  assign n41254 = ~n41326 & ~n41253;
  assign n41259 = ~n41786 & ~n41254;
  assign n41256 = ~n41255;
  assign n41258 = ~n41257 | ~n41256;
  assign n41260 = ~P2_INSTQUEUE_REG_9__0__SCAN_IN | ~n41318;
  assign P2_U3120 = ~n41261 | ~n41260;
  assign n41265 = ~n41795 & ~n41395;
  assign n41263 = ~n41597 | ~n41326;
  assign n41262 = ~P2_INSTQUEUE_REG_9__1__SCAN_IN | ~n41318;
  assign n41264 = ~n41263 | ~n41262;
  assign n41269 = ~n41265 & ~n41264;
  assign n41267 = ~n41310 & ~n41802;
  assign n41266 = ~n41690 & ~n41311;
  assign n41268 = ~n41267 & ~n41266;
  assign P2_U3121 = ~n41269 | ~n41268;
  assign n41273 = ~n41814 & ~n41395;
  assign n41271 = ~n41606 | ~n41326;
  assign n41270 = ~P2_INSTQUEUE_REG_9__2__SCAN_IN | ~n41318;
  assign n41272 = ~n41271 | ~n41270;
  assign n41277 = ~n41273 & ~n41272;
  assign n41275 = ~n41310 & ~n41807;
  assign n41274 = ~n41700 & ~n41311;
  assign n41276 = ~n41275 & ~n41274;
  assign P2_U3122 = ~n41277 | ~n41276;
  assign n41283 = ~n41819 & ~n41395;
  assign n41281 = ~n41615 | ~n41326;
  assign n41279 = ~n41311 & ~n41715;
  assign n41278 = ~n41826 & ~n41310;
  assign n41280 = ~n41279 & ~n41278;
  assign n41282 = ~n41281 | ~n41280;
  assign n41285 = ~n41283 & ~n41282;
  assign n41284 = ~P2_INSTQUEUE_REG_9__3__SCAN_IN | ~n41318;
  assign P2_U3123 = ~n41285 | ~n41284;
  assign n41291 = ~n41838 & ~n41395;
  assign n41289 = ~n41624 | ~n41326;
  assign n41287 = ~n41311 & ~n41725;
  assign n41286 = ~n41831 & ~n41310;
  assign n41288 = ~n41287 & ~n41286;
  assign n41290 = ~n41289 | ~n41288;
  assign n41293 = ~n41291 & ~n41290;
  assign n41292 = ~P2_INSTQUEUE_REG_9__4__SCAN_IN | ~n41318;
  assign P2_U3124 = ~n41293 | ~n41292;
  assign n41299 = ~n41850 & ~n41395;
  assign n41297 = ~n41633 | ~n41326;
  assign n41295 = ~n41311 & ~n41730;
  assign n41294 = ~n41843 & ~n41310;
  assign n41296 = ~n41295 & ~n41294;
  assign n41298 = ~n41297 | ~n41296;
  assign n41301 = ~n41299 & ~n41298;
  assign n41300 = ~P2_INSTQUEUE_REG_9__5__SCAN_IN | ~n41318;
  assign P2_U3125 = ~n41301 | ~n41300;
  assign n41305 = ~n41855 & ~n41395;
  assign n41303 = ~n41642 | ~n41326;
  assign n41302 = ~P2_INSTQUEUE_REG_9__6__SCAN_IN | ~n41318;
  assign n41304 = ~n41303 | ~n41302;
  assign n41309 = ~n41305 & ~n41304;
  assign n41307 = ~n41310 & ~n41862;
  assign n41306 = ~n41745 & ~n41311;
  assign n41308 = ~n41307 & ~n41306;
  assign P2_U3126 = ~n41309 | ~n41308;
  assign n41317 = ~n41395 & ~n41867;
  assign n41315 = ~n41652 | ~n41326;
  assign n41313 = ~n41310 & ~n41879;
  assign n41312 = ~n41753 & ~n41311;
  assign n41314 = ~n41313 & ~n41312;
  assign n41316 = ~n41315 | ~n41314;
  assign n41320 = ~n41317 & ~n41316;
  assign n41319 = ~P2_INSTQUEUE_REG_9__7__SCAN_IN | ~n41318;
  assign P2_U3127 = ~n41320 | ~n41319;
  assign n41321 = ~n42153;
  assign n41400 = ~n41411 & ~n42177;
  assign n41322 = ~n41395 | ~n41479;
  assign n41323 = ~n41322 | ~P2_STATEBS16_REG_SCAN_IN;
  assign n41334 = ~n41323 | ~n41785;
  assign n41325 = n41324 & P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN;
  assign n41423 = ~n41325 | ~P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN;
  assign n41338 = ~n41423 & ~P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n41332 = ~n41338 & ~n41326;
  assign n41327 = ~n41336 & ~n41338;
  assign n41328 = ~n41327 & ~n41664;
  assign n41403 = ~n41329 & ~n41328;
  assign n41346 = ~n41403 & ~n41672;
  assign n41331 = ~n41774 & ~n41395;
  assign n41396 = ~n41338;
  assign n41330 = ~n41775 & ~n41396;
  assign n41344 = ~n41331 & ~n41330;
  assign n41333 = ~n41332;
  assign n41335 = ~n41334 & ~n41333;
  assign n41342 = ~n41335 & ~n41786;
  assign n41337 = ~n41336;
  assign n41339 = ~n41337 & ~P2_STATE2_REG_3__SCAN_IN;
  assign n41340 = ~n41339 & ~n41338;
  assign n41341 = ~n41340 | ~n41002;
  assign n41343 = ~P2_INSTQUEUE_REG_10__0__SCAN_IN | ~n41399;
  assign n41345 = ~n41344 | ~n41343;
  assign n41348 = ~n41346 & ~n41345;
  assign n41347 = ~n41400 | ~n41675;
  assign P2_U3128 = ~n41348 | ~n41347;
  assign n41352 = ~n41796 & ~n41396;
  assign n41350 = ~P2_INSTQUEUE_REG_10__1__SCAN_IN | ~n41399;
  assign n41349 = ~n41400 | ~n41693;
  assign n41351 = ~n41350 | ~n41349;
  assign n41356 = ~n41352 & ~n41351;
  assign n41354 = ~n41395 & ~n41802;
  assign n41353 = ~n41690 & ~n41403;
  assign n41355 = ~n41354 & ~n41353;
  assign P2_U3129 = ~n41356 | ~n41355;
  assign n41358 = ~n41395 & ~n41807;
  assign n41357 = ~n41808 & ~n41396;
  assign n41364 = ~n41358 & ~n41357;
  assign n41360 = ~P2_INSTQUEUE_REG_10__2__SCAN_IN | ~n41399;
  assign n41359 = ~n41400 | ~n41703;
  assign n41362 = ~n41360 | ~n41359;
  assign n41361 = ~n41403 & ~n41700;
  assign n41363 = ~n41362 & ~n41361;
  assign P2_U3130 = ~n41364 | ~n41363;
  assign n41366 = ~n41395 & ~n41826;
  assign n41365 = ~n41820 & ~n41396;
  assign n41372 = ~n41366 & ~n41365;
  assign n41368 = ~P2_INSTQUEUE_REG_10__3__SCAN_IN | ~n41399;
  assign n41367 = ~n41400 | ~n41710;
  assign n41370 = ~n41368 | ~n41367;
  assign n41369 = ~n41403 & ~n41715;
  assign n41371 = ~n41370 & ~n41369;
  assign P2_U3131 = ~n41372 | ~n41371;
  assign n41376 = ~n41832 & ~n41396;
  assign n41374 = ~n41395 & ~n41831;
  assign n41373 = ~n41725 & ~n41403;
  assign n41375 = ~n41374 & ~n41373;
  assign n41377 = ~P2_INSTQUEUE_REG_10__4__SCAN_IN | ~n41399;
  assign P2_U3132 = ~n41378 | ~n41377;
  assign n41380 = ~n41395 & ~n41843;
  assign n41379 = ~n41844 & ~n41396;
  assign n41386 = ~n41380 & ~n41379;
  assign n41382 = ~P2_INSTQUEUE_REG_10__5__SCAN_IN | ~n41399;
  assign n41381 = ~n41400 | ~n41733;
  assign n41384 = ~n41382 | ~n41381;
  assign n41383 = ~n41403 & ~n41730;
  assign n41385 = ~n41384 & ~n41383;
  assign P2_U3133 = ~n41386 | ~n41385;
  assign n41392 = ~n41856 & ~n41396;
  assign n41388 = ~n41395 & ~n41862;
  assign n41387 = ~n41745 & ~n41403;
  assign n41390 = ~n41388 & ~n41387;
  assign n41389 = ~n41400 | ~n41740;
  assign n41391 = ~n41390 | ~n41389;
  assign n41394 = ~n41392 & ~n41391;
  assign n41393 = ~P2_INSTQUEUE_REG_10__6__SCAN_IN | ~n41399;
  assign P2_U3134 = ~n41394 | ~n41393;
  assign n41398 = ~n41395 & ~n41879;
  assign n41397 = ~n41870 & ~n41396;
  assign n41407 = ~n41398 & ~n41397;
  assign n41402 = ~P2_INSTQUEUE_REG_10__7__SCAN_IN | ~n41399;
  assign n41401 = ~n41400 | ~n41756;
  assign n41405 = ~n41402 | ~n41401;
  assign n41404 = ~n41403 & ~n41753;
  assign n41406 = ~n41405 & ~n41404;
  assign P2_U3135 = ~n41407 | ~n41406;
  assign n41478 = ~n41423 & ~n41575;
  assign n41408 = ~n41418 & ~n41478;
  assign n41410 = ~n41408 & ~n41664;
  assign n41409 = ~n41002 & ~n41423;
  assign n41417 = ~n41672 & ~n41477;
  assign n41415 = ~n41579 | ~n41478;
  assign n41413 = ~n41569 & ~n41765;
  assign n41412 = ~n41479 & ~n41774;
  assign n41414 = ~n41413 & ~n41412;
  assign n41416 = ~n41415 | ~n41414;
  assign n41428 = ~n41417 & ~n41416;
  assign n41419 = ~n41418 | ~n42196;
  assign n41420 = ~n41419 | ~n41002;
  assign n41421 = ~n41478 & ~n41420;
  assign n41426 = ~n41786 & ~n41421;
  assign n41424 = ~P2_STATEBS16_REG_SCAN_IN | ~n41422;
  assign n41425 = ~n41424 | ~n41423;
  assign n41427 = ~P2_INSTQUEUE_REG_11__0__SCAN_IN | ~n41486;
  assign P2_U3136 = ~n41428 | ~n41427;
  assign n41434 = ~n41690 & ~n41477;
  assign n41432 = ~n41597 | ~n41478;
  assign n41430 = ~n41569 & ~n41795;
  assign n41429 = ~n41479 & ~n41802;
  assign n41431 = ~n41430 & ~n41429;
  assign n41433 = ~n41432 | ~n41431;
  assign n41436 = ~n41434 & ~n41433;
  assign n41435 = ~P2_INSTQUEUE_REG_11__1__SCAN_IN | ~n41486;
  assign P2_U3137 = ~n41436 | ~n41435;
  assign n41442 = ~n41700 & ~n41477;
  assign n41440 = ~n41606 | ~n41478;
  assign n41438 = ~n41569 & ~n41814;
  assign n41437 = ~n41479 & ~n41807;
  assign n41439 = ~n41438 & ~n41437;
  assign n41441 = ~n41440 | ~n41439;
  assign n41444 = ~n41442 & ~n41441;
  assign n41443 = ~P2_INSTQUEUE_REG_11__2__SCAN_IN | ~n41486;
  assign P2_U3138 = ~n41444 | ~n41443;
  assign n41450 = ~n41715 & ~n41477;
  assign n41448 = ~n41615 | ~n41478;
  assign n41446 = ~n41569 & ~n41819;
  assign n41445 = ~n41479 & ~n41826;
  assign n41447 = ~n41446 & ~n41445;
  assign n41449 = ~n41448 | ~n41447;
  assign n41452 = ~n41450 & ~n41449;
  assign n41451 = ~P2_INSTQUEUE_REG_11__3__SCAN_IN | ~n41486;
  assign P2_U3139 = ~n41452 | ~n41451;
  assign n41458 = ~n41725 & ~n41477;
  assign n41456 = ~n41624 | ~n41478;
  assign n41454 = ~n41569 & ~n41838;
  assign n41453 = ~n41479 & ~n41831;
  assign n41455 = ~n41454 & ~n41453;
  assign n41457 = ~n41456 | ~n41455;
  assign n41460 = ~n41458 & ~n41457;
  assign n41459 = ~P2_INSTQUEUE_REG_11__4__SCAN_IN | ~n41486;
  assign P2_U3140 = ~n41460 | ~n41459;
  assign n41466 = ~n41730 & ~n41477;
  assign n41464 = ~n41633 | ~n41478;
  assign n41462 = ~n41569 & ~n41850;
  assign n41461 = ~n41479 & ~n41843;
  assign n41463 = ~n41462 & ~n41461;
  assign n41465 = ~n41464 | ~n41463;
  assign n41468 = ~n41466 & ~n41465;
  assign n41467 = ~P2_INSTQUEUE_REG_11__5__SCAN_IN | ~n41486;
  assign P2_U3141 = ~n41468 | ~n41467;
  assign n41474 = ~n41745 & ~n41477;
  assign n41472 = ~n41642 | ~n41478;
  assign n41470 = ~n41569 & ~n41855;
  assign n41469 = ~n41479 & ~n41862;
  assign n41471 = ~n41470 & ~n41469;
  assign n41473 = ~n41472 | ~n41471;
  assign n41476 = ~n41474 & ~n41473;
  assign n41475 = ~P2_INSTQUEUE_REG_11__6__SCAN_IN | ~n41486;
  assign P2_U3142 = ~n41476 | ~n41475;
  assign n41485 = ~n41753 & ~n41477;
  assign n41483 = ~n41652 | ~n41478;
  assign n41481 = ~n41569 & ~n41867;
  assign n41480 = ~n41479 & ~n41879;
  assign n41482 = ~n41481 & ~n41480;
  assign n41484 = ~n41483 | ~n41482;
  assign n41488 = ~n41485 & ~n41484;
  assign n41487 = ~P2_INSTQUEUE_REG_11__7__SCAN_IN | ~n41486;
  assign P2_U3143 = ~n41488 | ~n41487;
  assign n41502 = ~n41774 & ~n41569;
  assign n41564 = ~P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & ~n41591;
  assign n41500 = ~n41579 | ~n41564;
  assign n41498 = ~n41765 & ~n41653;
  assign n41492 = ~n41503 & ~n41564;
  assign n41496 = ~n41492 & ~n41664;
  assign n41508 = ~n41494 | ~n41493;
  assign n41495 = ~n41508 & ~n41002;
  assign n41497 = ~n41562 & ~n41672;
  assign n41499 = ~n41498 & ~n41497;
  assign n41501 = ~n41500 | ~n41499;
  assign n41513 = ~n41502 & ~n41501;
  assign n41504 = ~n41503 | ~n42196;
  assign n41505 = ~n41504 | ~n41002;
  assign n41506 = ~n41564 & ~n41505;
  assign n41511 = ~n41786 & ~n41506;
  assign n41507 = ~n41569 | ~n41653;
  assign n41509 = ~P2_STATEBS16_REG_SCAN_IN | ~n41507;
  assign n41510 = ~n41509 | ~n41508;
  assign n41512 = ~P2_INSTQUEUE_REG_12__0__SCAN_IN | ~n41563;
  assign P2_U3144 = ~n41513 | ~n41512;
  assign n41517 = ~n41690 & ~n41562;
  assign n41515 = ~P2_INSTQUEUE_REG_12__1__SCAN_IN | ~n41563;
  assign n41514 = ~n41564 | ~n41597;
  assign n41516 = ~n41515 | ~n41514;
  assign n41521 = ~n41517 & ~n41516;
  assign n41519 = ~n41653 & ~n41795;
  assign n41518 = ~n41569 & ~n41802;
  assign n41520 = ~n41519 & ~n41518;
  assign P2_U3145 = ~n41521 | ~n41520;
  assign n41525 = ~n41700 & ~n41562;
  assign n41523 = ~P2_INSTQUEUE_REG_12__2__SCAN_IN | ~n41563;
  assign n41522 = ~n41564 | ~n41606;
  assign n41524 = ~n41523 | ~n41522;
  assign n41529 = ~n41525 & ~n41524;
  assign n41527 = ~n41653 & ~n41814;
  assign n41526 = ~n41569 & ~n41807;
  assign n41528 = ~n41527 & ~n41526;
  assign P2_U3146 = ~n41529 | ~n41528;
  assign n41533 = ~n41715 & ~n41562;
  assign n41531 = ~P2_INSTQUEUE_REG_12__3__SCAN_IN | ~n41563;
  assign n41530 = ~n41615 | ~n41564;
  assign n41532 = ~n41531 | ~n41530;
  assign n41537 = ~n41533 & ~n41532;
  assign n41535 = ~n41653 & ~n41819;
  assign n41534 = ~n41569 & ~n41826;
  assign n41536 = ~n41535 & ~n41534;
  assign P2_U3147 = ~n41537 | ~n41536;
  assign n41541 = ~n41725 & ~n41562;
  assign n41539 = ~P2_INSTQUEUE_REG_12__4__SCAN_IN | ~n41563;
  assign n41538 = ~n41564 | ~n41624;
  assign n41540 = ~n41539 | ~n41538;
  assign n41545 = ~n41541 & ~n41540;
  assign n41543 = ~n41653 & ~n41838;
  assign n41542 = ~n41569 & ~n41831;
  assign n41544 = ~n41543 & ~n41542;
  assign P2_U3148 = ~n41545 | ~n41544;
  assign n41549 = ~n41730 & ~n41562;
  assign n41547 = ~P2_INSTQUEUE_REG_12__5__SCAN_IN | ~n41563;
  assign n41546 = ~n41633 | ~n41564;
  assign n41548 = ~n41547 | ~n41546;
  assign n41553 = ~n41549 & ~n41548;
  assign n41551 = ~n41653 & ~n41850;
  assign n41550 = ~n41569 & ~n41843;
  assign n41552 = ~n41551 & ~n41550;
  assign P2_U3149 = ~n41553 | ~n41552;
  assign n41557 = ~n41745 & ~n41562;
  assign n41555 = ~P2_INSTQUEUE_REG_12__6__SCAN_IN | ~n41563;
  assign n41554 = ~n41564 | ~n41642;
  assign n41556 = ~n41555 | ~n41554;
  assign n41561 = ~n41557 & ~n41556;
  assign n41559 = ~n41653 & ~n41855;
  assign n41558 = ~n41569 & ~n41862;
  assign n41560 = ~n41559 & ~n41558;
  assign P2_U3150 = ~n41561 | ~n41560;
  assign n41568 = ~n41753 & ~n41562;
  assign n41566 = ~P2_INSTQUEUE_REG_12__7__SCAN_IN | ~n41563;
  assign n41565 = ~n41564 | ~n41652;
  assign n41567 = ~n41566 | ~n41565;
  assign n41573 = ~n41568 & ~n41567;
  assign n41571 = ~n41653 & ~n41867;
  assign n41570 = ~n41569 & ~n41879;
  assign n41572 = ~n41571 & ~n41570;
  assign P2_U3151 = ~n41573 | ~n41572;
  assign n41586 = ~n41574;
  assign n41576 = ~n41586 & ~n41680;
  assign n41578 = ~n41576 & ~n41664;
  assign n41577 = ~n41002 & ~n41591;
  assign n41585 = ~n41672 & ~n41651;
  assign n41583 = ~n41579 | ~n41680;
  assign n41581 = ~n41751 & ~n41765;
  assign n41580 = ~n41653 & ~n41774;
  assign n41582 = ~n41581 & ~n41580;
  assign n41584 = ~n41583 | ~n41582;
  assign n41596 = ~n41585 & ~n41584;
  assign n41587 = ~n41586 | ~n42196;
  assign n41588 = ~n41587 | ~n41002;
  assign n41589 = ~n41680 & ~n41588;
  assign n41594 = ~n41786 & ~n41589;
  assign n41592 = ~P2_STATEBS16_REG_SCAN_IN | ~n41590;
  assign n41593 = ~n41592 | ~n41591;
  assign n41595 = ~P2_INSTQUEUE_REG_13__0__SCAN_IN | ~n41660;
  assign P2_U3152 = ~n41596 | ~n41595;
  assign n41603 = ~n41690 & ~n41651;
  assign n41601 = ~n41680 | ~n41597;
  assign n41599 = ~n41751 & ~n41795;
  assign n41598 = ~n41653 & ~n41802;
  assign n41600 = ~n41599 & ~n41598;
  assign n41602 = ~n41601 | ~n41600;
  assign n41605 = ~n41603 & ~n41602;
  assign n41604 = ~P2_INSTQUEUE_REG_13__1__SCAN_IN | ~n41660;
  assign P2_U3153 = ~n41605 | ~n41604;
  assign n41612 = ~n41700 & ~n41651;
  assign n41610 = ~n41680 | ~n41606;
  assign n41608 = ~n41751 & ~n41814;
  assign n41607 = ~n41653 & ~n41807;
  assign n41609 = ~n41608 & ~n41607;
  assign n41611 = ~n41610 | ~n41609;
  assign n41614 = ~n41612 & ~n41611;
  assign n41613 = ~P2_INSTQUEUE_REG_13__2__SCAN_IN | ~n41660;
  assign P2_U3154 = ~n41614 | ~n41613;
  assign n41621 = ~n41715 & ~n41651;
  assign n41619 = ~n41615 | ~n41680;
  assign n41617 = ~n41751 & ~n41819;
  assign n41616 = ~n41653 & ~n41826;
  assign n41618 = ~n41617 & ~n41616;
  assign n41620 = ~n41619 | ~n41618;
  assign n41623 = ~n41621 & ~n41620;
  assign n41622 = ~P2_INSTQUEUE_REG_13__3__SCAN_IN | ~n41660;
  assign P2_U3155 = ~n41623 | ~n41622;
  assign n41630 = ~n41725 & ~n41651;
  assign n41628 = ~n41680 | ~n41624;
  assign n41626 = ~n41751 & ~n41838;
  assign n41625 = ~n41653 & ~n41831;
  assign n41627 = ~n41626 & ~n41625;
  assign n41629 = ~n41628 | ~n41627;
  assign n41632 = ~n41630 & ~n41629;
  assign n41631 = ~P2_INSTQUEUE_REG_13__4__SCAN_IN | ~n41660;
  assign P2_U3156 = ~n41632 | ~n41631;
  assign n41639 = ~n41730 & ~n41651;
  assign n41637 = ~n41633 | ~n41680;
  assign n41635 = ~n41751 & ~n41850;
  assign n41634 = ~n41653 & ~n41843;
  assign n41636 = ~n41635 & ~n41634;
  assign n41638 = ~n41637 | ~n41636;
  assign n41641 = ~n41639 & ~n41638;
  assign n41640 = ~P2_INSTQUEUE_REG_13__5__SCAN_IN | ~n41660;
  assign P2_U3157 = ~n41641 | ~n41640;
  assign n41648 = ~n41745 & ~n41651;
  assign n41646 = ~n41680 | ~n41642;
  assign n41644 = ~n41751 & ~n41855;
  assign n41643 = ~n41653 & ~n41862;
  assign n41645 = ~n41644 & ~n41643;
  assign n41647 = ~n41646 | ~n41645;
  assign n41650 = ~n41648 & ~n41647;
  assign n41649 = ~P2_INSTQUEUE_REG_13__6__SCAN_IN | ~n41660;
  assign P2_U3158 = ~n41650 | ~n41649;
  assign n41659 = ~n41753 & ~n41651;
  assign n41657 = ~n41680 | ~n41652;
  assign n41655 = ~n41751 & ~n41867;
  assign n41654 = ~n41653 & ~n41879;
  assign n41656 = ~n41655 & ~n41654;
  assign n41658 = ~n41657 | ~n41656;
  assign n41662 = ~n41659 & ~n41658;
  assign n41661 = ~P2_INSTQUEUE_REG_13__7__SCAN_IN | ~n41660;
  assign P2_U3159 = ~n41662 | ~n41661;
  assign n41663 = ~P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & ~n41768;
  assign n41750 = ~n41663 | ~P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN;
  assign n41679 = ~n41775 & ~n41750;
  assign n41674 = ~n41751 & ~n41774;
  assign n41668 = ~n41750;
  assign n41665 = ~n27889 & ~n41668;
  assign n41671 = ~n41665 & ~n41664;
  assign n41757 = ~n41788 & ~n42177;
  assign n41666 = ~n41878 | ~n41751;
  assign n41667 = ~n41666 | ~P2_STATEBS16_REG_SCAN_IN;
  assign n41681 = ~n41667 | ~n41785;
  assign n41669 = ~n41668 & ~n41680;
  assign n41670 = ~n41681 & ~n41669;
  assign n41752 = ~n41671 & ~n41670;
  assign n41673 = ~n41672 & ~n41752;
  assign n41677 = ~n41674 & ~n41673;
  assign n41676 = ~n41757 | ~n41675;
  assign n41678 = ~n41677 | ~n41676;
  assign n41689 = ~n41679 & ~n41678;
  assign n41684 = n41681 | n41680;
  assign n41682 = ~n27889 | ~n42196;
  assign n41683 = ~n41682 | ~n41002;
  assign n41685 = ~n41684 | ~n41683;
  assign n41687 = ~n41685 | ~n41750;
  assign n41688 = ~P2_INSTQUEUE_REG_14__0__SCAN_IN | ~n41762;
  assign P2_U3160 = ~n41689 | ~n41688;
  assign n41697 = ~n41796 & ~n41750;
  assign n41692 = ~n41751 & ~n41802;
  assign n41691 = ~n41690 & ~n41752;
  assign n41695 = ~n41692 & ~n41691;
  assign n41694 = ~n41757 | ~n41693;
  assign n41696 = ~n41695 | ~n41694;
  assign n41699 = ~n41697 & ~n41696;
  assign n41698 = ~P2_INSTQUEUE_REG_14__1__SCAN_IN | ~n41762;
  assign P2_U3161 = ~n41699 | ~n41698;
  assign n41707 = ~n41808 & ~n41750;
  assign n41702 = ~n41751 & ~n41807;
  assign n41701 = ~n41700 & ~n41752;
  assign n41705 = ~n41702 & ~n41701;
  assign n41704 = ~n41757 | ~n41703;
  assign n41706 = ~n41705 | ~n41704;
  assign n41709 = ~n41707 & ~n41706;
  assign n41708 = ~P2_INSTQUEUE_REG_14__2__SCAN_IN | ~n41762;
  assign P2_U3162 = ~n41709 | ~n41708;
  assign n41714 = ~n41820 & ~n41750;
  assign n41712 = ~P2_INSTQUEUE_REG_14__3__SCAN_IN | ~n41762;
  assign n41711 = ~n41757 | ~n41710;
  assign n41713 = ~n41712 | ~n41711;
  assign n41719 = ~n41714 & ~n41713;
  assign n41717 = ~n41751 & ~n41826;
  assign n41716 = ~n41715 & ~n41752;
  assign n41718 = ~n41717 & ~n41716;
  assign P2_U3163 = ~n41719 | ~n41718;
  assign n41724 = ~n41832 & ~n41750;
  assign n41722 = ~P2_INSTQUEUE_REG_14__4__SCAN_IN | ~n41762;
  assign n41721 = ~n41757 | ~n41720;
  assign n41723 = ~n41722 | ~n41721;
  assign n41729 = ~n41724 & ~n41723;
  assign n41727 = ~n41751 & ~n41831;
  assign n41726 = ~n41725 & ~n41752;
  assign n41728 = ~n41727 & ~n41726;
  assign P2_U3164 = ~n41729 | ~n41728;
  assign n41737 = ~n41844 & ~n41750;
  assign n41732 = ~n41751 & ~n41843;
  assign n41731 = ~n41730 & ~n41752;
  assign n41735 = ~n41732 & ~n41731;
  assign n41734 = ~n41757 | ~n41733;
  assign n41736 = ~n41735 | ~n41734;
  assign n41739 = ~n41737 & ~n41736;
  assign n41738 = ~P2_INSTQUEUE_REG_14__5__SCAN_IN | ~n41762;
  assign P2_U3165 = ~n41739 | ~n41738;
  assign n41744 = ~n41856 & ~n41750;
  assign n41742 = ~P2_INSTQUEUE_REG_14__6__SCAN_IN | ~n41762;
  assign n41741 = ~n41757 | ~n41740;
  assign n41743 = ~n41742 | ~n41741;
  assign n41749 = ~n41744 & ~n41743;
  assign n41747 = ~n41751 & ~n41862;
  assign n41746 = ~n41745 & ~n41752;
  assign n41748 = ~n41747 & ~n41746;
  assign P2_U3166 = ~n41749 | ~n41748;
  assign n41761 = ~n41870 & ~n41750;
  assign n41755 = ~n41751 & ~n41879;
  assign n41754 = ~n41753 & ~n41752;
  assign n41759 = ~n41755 & ~n41754;
  assign n41758 = ~n41757 | ~n41756;
  assign n41760 = ~n41759 | ~n41758;
  assign n41764 = ~n41761 & ~n41760;
  assign n41763 = ~P2_INSTQUEUE_REG_14__7__SCAN_IN | ~n41762;
  assign P2_U3167 = ~n41764 | ~n41763;
  assign n41781 = ~n41868 & ~n41765;
  assign n41767 = ~n41766 | ~n41869;
  assign n41772 = ~n41767 | ~P2_STATE2_REG_2__SCAN_IN;
  assign n41791 = ~n41769 & ~n41768;
  assign n41770 = ~n41791;
  assign n41771 = n41002 | n41770;
  assign n41874 = ~n41772 | ~n41771;
  assign n41779 = ~n41773 | ~n41874;
  assign n41777 = ~n41878 & ~n41774;
  assign n41776 = ~n41775 & ~n41869;
  assign n41778 = ~n41777 & ~n41776;
  assign n41780 = ~n41779 | ~n41778;
  assign n41794 = ~n41781 & ~n41780;
  assign n41783 = ~n41782 | ~n42196;
  assign n41784 = ~n41783 | ~n41869;
  assign n41787 = ~n41785 & ~n41784;
  assign n41792 = ~n41787 & ~n41786;
  assign n41790 = ~n41789 & ~n41788;
  assign n41793 = ~P2_INSTQUEUE_REG_15__0__SCAN_IN | ~n41873;
  assign P2_U3168 = ~n41794 | ~n41793;
  assign n41798 = ~n41868 & ~n41795;
  assign n41797 = ~n41796 & ~n41869;
  assign n41806 = ~n41798 & ~n41797;
  assign n41801 = ~P2_INSTQUEUE_REG_15__1__SCAN_IN | ~n41873;
  assign n41800 = ~n41799 | ~n41874;
  assign n41804 = ~n41801 | ~n41800;
  assign n41803 = ~n41802 & ~n41878;
  assign n41805 = ~n41804 & ~n41803;
  assign P2_U3169 = ~n41806 | ~n41805;
  assign n41810 = ~n41878 & ~n41807;
  assign n41809 = ~n41808 & ~n41869;
  assign n41818 = ~n41810 & ~n41809;
  assign n41813 = ~P2_INSTQUEUE_REG_15__2__SCAN_IN | ~n41873;
  assign n41812 = ~n41811 | ~n41874;
  assign n41816 = ~n41813 | ~n41812;
  assign n41815 = ~n41814 & ~n41868;
  assign n41817 = ~n41816 & ~n41815;
  assign P2_U3170 = ~n41818 | ~n41817;
  assign n41822 = ~n41868 & ~n41819;
  assign n41821 = ~n41820 & ~n41869;
  assign n41830 = ~n41822 & ~n41821;
  assign n41825 = ~P2_INSTQUEUE_REG_15__3__SCAN_IN | ~n41873;
  assign n41824 = ~n41823 | ~n41874;
  assign n41828 = ~n41825 | ~n41824;
  assign n41827 = ~n41826 & ~n41878;
  assign n41829 = ~n41828 & ~n41827;
  assign P2_U3171 = ~n41830 | ~n41829;
  assign n41834 = ~n41878 & ~n41831;
  assign n41833 = ~n41832 & ~n41869;
  assign n41842 = ~n41834 & ~n41833;
  assign n41837 = ~P2_INSTQUEUE_REG_15__4__SCAN_IN | ~n41873;
  assign n41836 = ~n41835 | ~n41874;
  assign n41840 = ~n41837 | ~n41836;
  assign n41839 = ~n41838 & ~n41868;
  assign n41841 = ~n41840 & ~n41839;
  assign P2_U3172 = ~n41842 | ~n41841;
  assign n41846 = ~n41878 & ~n41843;
  assign n41845 = ~n41844 & ~n41869;
  assign n41854 = ~n41846 & ~n41845;
  assign n41849 = ~P2_INSTQUEUE_REG_15__5__SCAN_IN | ~n41873;
  assign n41848 = ~n41847 | ~n41874;
  assign n41852 = ~n41849 | ~n41848;
  assign n41851 = ~n41850 & ~n41868;
  assign n41853 = ~n41852 & ~n41851;
  assign P2_U3173 = ~n41854 | ~n41853;
  assign n41858 = ~n41868 & ~n41855;
  assign n41857 = ~n41856 & ~n41869;
  assign n41866 = ~n41858 & ~n41857;
  assign n41861 = ~P2_INSTQUEUE_REG_15__6__SCAN_IN | ~n41873;
  assign n41860 = ~n41859 | ~n41874;
  assign n41864 = ~n41861 | ~n41860;
  assign n41863 = ~n41862 & ~n41878;
  assign n41865 = ~n41864 & ~n41863;
  assign P2_U3174 = ~n41866 | ~n41865;
  assign n41872 = ~n41868 & ~n41867;
  assign n41871 = ~n41870 & ~n41869;
  assign n41883 = ~n41872 & ~n41871;
  assign n41877 = ~P2_INSTQUEUE_REG_15__7__SCAN_IN | ~n41873;
  assign n41876 = ~n41875 | ~n41874;
  assign n41881 = ~n41877 | ~n41876;
  assign n41880 = ~n41879 & ~n41878;
  assign n41882 = ~n41881 & ~n41880;
  assign P2_U3175 = ~n41883 | ~n41882;
  assign n41886 = ~n41885 & ~n41884;
  assign n41892 = n41886 | n42123;
  assign n41888 = n42137 | n41887;
  assign n41889 = ~n41888 | ~n42075;
  assign n41891 = ~n41890 | ~n41889;
  assign P2_U3177 = ~n22977 | ~n41893;
  assign P2_U3179 = P2_DATAWIDTH_REG_31__SCAN_IN & n22820;
  assign P2_U3180 = P2_DATAWIDTH_REG_30__SCAN_IN & n22819;
  assign P2_U3181 = P2_DATAWIDTH_REG_29__SCAN_IN & n22820;
  assign P2_U3182 = P2_DATAWIDTH_REG_28__SCAN_IN & n22819;
  assign P2_U3183 = P2_DATAWIDTH_REG_27__SCAN_IN & n22820;
  assign P2_U3184 = P2_DATAWIDTH_REG_26__SCAN_IN & n22819;
  assign P2_U3185 = P2_DATAWIDTH_REG_25__SCAN_IN & n22820;
  assign P2_U3186 = P2_DATAWIDTH_REG_24__SCAN_IN & n22819;
  assign P2_U3187 = P2_DATAWIDTH_REG_23__SCAN_IN & n22820;
  assign P2_U3188 = P2_DATAWIDTH_REG_22__SCAN_IN & n22819;
  assign P2_U3189 = P2_DATAWIDTH_REG_21__SCAN_IN & n22820;
  assign P2_U3190 = P2_DATAWIDTH_REG_20__SCAN_IN & n22819;
  assign P2_U3191 = P2_DATAWIDTH_REG_19__SCAN_IN & n22820;
  assign P2_U3192 = P2_DATAWIDTH_REG_18__SCAN_IN & n22819;
  assign P2_U3193 = P2_DATAWIDTH_REG_17__SCAN_IN & n22820;
  assign P2_U3194 = P2_DATAWIDTH_REG_16__SCAN_IN & n22819;
  assign P2_U3195 = P2_DATAWIDTH_REG_15__SCAN_IN & n22820;
  assign P2_U3196 = P2_DATAWIDTH_REG_14__SCAN_IN & n22819;
  assign P2_U3197 = P2_DATAWIDTH_REG_13__SCAN_IN & n22819;
  assign P2_U3198 = P2_DATAWIDTH_REG_12__SCAN_IN & n22820;
  assign P2_U3199 = P2_DATAWIDTH_REG_11__SCAN_IN & n22819;
  assign P2_U3200 = P2_DATAWIDTH_REG_10__SCAN_IN & n22820;
  assign P2_U3201 = P2_DATAWIDTH_REG_9__SCAN_IN & n22820;
  assign P2_U3202 = P2_DATAWIDTH_REG_8__SCAN_IN & n22819;
  assign P2_U3203 = P2_DATAWIDTH_REG_7__SCAN_IN & n22820;
  assign P2_U3204 = P2_DATAWIDTH_REG_6__SCAN_IN & n22819;
  assign P2_U3205 = P2_DATAWIDTH_REG_5__SCAN_IN & n22820;
  assign P2_U3206 = P2_DATAWIDTH_REG_4__SCAN_IN & n22819;
  assign P2_U3207 = P2_DATAWIDTH_REG_3__SCAN_IN & n22820;
  assign P2_U3208 = P2_DATAWIDTH_REG_2__SCAN_IN & n22819;
  assign n41917 = ~n41895 | ~P2_STATE_REG_1__SCAN_IN;
  assign n41903 = P2_STATE_REG_0__SCAN_IN & P2_REQUESTPENDING_REG_SCAN_IN;
  assign n41896 = ~n41917 | ~n41903;
  assign n41902 = ~n41896 | ~n41926;
  assign n41921 = ~n44540 & ~n41897;
  assign n41898 = ~P2_REQUESTPENDING_REG_SCAN_IN | ~n41918;
  assign n41899 = ~n41911 | ~n41898;
  assign n41900 = ~n42224 & ~n41899;
  assign n41901 = ~n41921 & ~n41900;
  assign P2_U3209 = ~n41902 | ~n41901;
  assign n41904 = ~HOLD | ~P2_STATE_REG_2__SCAN_IN;
  assign n41905 = ~n41904 | ~n41903;
  assign n41908 = ~n41905 | ~n41917;
  assign n41914 = ~P2_REQUESTPENDING_REG_SCAN_IN & ~HOLD;
  assign n41906 = ~P2_STATE_REG_1__SCAN_IN | ~n41926;
  assign n41907 = ~n41914 & ~n41906;
  assign n41910 = ~n41908 & ~n41907;
  assign P2_U3210 = ~n41910 | ~n41909;
  assign n41913 = ~NA & ~n41917;
  assign n41912 = ~P2_REQUESTPENDING_REG_SCAN_IN & ~n41911;
  assign n41915 = ~n41913 & ~n41912;
  assign n41916 = ~n41915 & ~n41914;
  assign n41925 = ~P2_STATE_REG_0__SCAN_IN | ~n41916;
  assign n41919 = ~n41918 | ~n41917;
  assign n41922 = ~n41920 & ~n41919;
  assign n41923 = ~n41922 & ~n41921;
  assign n41924 = ~P2_STATE_REG_2__SCAN_IN | ~n41923;
  assign P2_U3211 = ~n41925 | ~n41924;
  assign n41928 = ~n27692 & ~n42024;
  assign n42023 = ~n42224 | ~n41926;
  assign n41927 = ~n27699 & ~n42023;
  assign n41930 = ~n41928 & ~n41927;
  assign n41929 = ~P2_ADDRESS_REG_0__SCAN_IN | ~n42065;
  assign P2_U3212 = ~n41930 | ~n41929;
  assign n41932 = ~n27699 & ~n42024;
  assign n41935 = ~P2_REIP_REG_3__SCAN_IN;
  assign n41931 = ~n41935 & ~n42023;
  assign n41934 = ~n41932 & ~n41931;
  assign n41933 = ~P2_ADDRESS_REG_1__SCAN_IN | ~n42065;
  assign P2_U3213 = ~n41934 | ~n41933;
  assign n41937 = ~n28339 & ~n42023;
  assign n41936 = ~n41935 & ~n42024;
  assign n41939 = ~n41937 & ~n41936;
  assign n41938 = ~P2_ADDRESS_REG_2__SCAN_IN | ~n42065;
  assign P2_U3214 = ~n41939 | ~n41938;
  assign n41943 = ~P2_ADDRESS_REG_3__SCAN_IN | ~n42223;
  assign n41941 = ~n28339 & ~n42024;
  assign n41940 = ~n32586 & ~n42023;
  assign n41942 = ~n41941 & ~n41940;
  assign P2_U3215 = ~n41943 | ~n41942;
  assign n41945 = ~n28354 & ~n42023;
  assign n41944 = ~n32586 & ~n42024;
  assign n41947 = ~n41945 & ~n41944;
  assign n41946 = ~P2_ADDRESS_REG_4__SCAN_IN | ~n42065;
  assign P2_U3216 = ~n41947 | ~n41946;
  assign n41949 = ~n28361 & ~n42023;
  assign n41948 = ~n28354 & ~n42024;
  assign n41951 = ~n41949 & ~n41948;
  assign n41950 = ~P2_ADDRESS_REG_5__SCAN_IN | ~n42065;
  assign P2_U3217 = ~n41951 | ~n41950;
  assign n41955 = ~P2_ADDRESS_REG_6__SCAN_IN | ~n42065;
  assign n41953 = ~n28361 & ~n42024;
  assign n41952 = ~n28369 & ~n42023;
  assign n41954 = ~n41953 & ~n41952;
  assign P2_U3218 = ~n41955 | ~n41954;
  assign n41959 = ~P2_ADDRESS_REG_7__SCAN_IN | ~n42065;
  assign n41957 = ~n28369 & ~n42024;
  assign n41956 = ~n32974 & ~n42023;
  assign n41958 = ~n41957 & ~n41956;
  assign P2_U3219 = ~n41959 | ~n41958;
  assign n41961 = ~n28382 & ~n42023;
  assign n41960 = ~n32974 & ~n42024;
  assign n41963 = ~n41961 & ~n41960;
  assign n41962 = ~P2_ADDRESS_REG_8__SCAN_IN | ~n42223;
  assign P2_U3220 = ~n41963 | ~n41962;
  assign n41967 = ~P2_ADDRESS_REG_9__SCAN_IN | ~n42223;
  assign n41965 = ~n28382 & ~n42024;
  assign n41964 = ~n28389 & ~n42023;
  assign n41966 = ~n41965 & ~n41964;
  assign P2_U3221 = ~n41967 | ~n41966;
  assign n41971 = ~P2_ADDRESS_REG_10__SCAN_IN | ~n42065;
  assign n41969 = ~n28389 & ~n42024;
  assign n41968 = ~n28396 & ~n42023;
  assign n41970 = ~n41969 & ~n41968;
  assign P2_U3222 = ~n41971 | ~n41970;
  assign n41973 = ~n28396 & ~n42024;
  assign n41972 = ~n28403 & ~n42023;
  assign n41975 = ~n41973 & ~n41972;
  assign n41974 = ~P2_ADDRESS_REG_11__SCAN_IN | ~n42223;
  assign P2_U3223 = ~n41975 | ~n41974;
  assign n41979 = ~P2_ADDRESS_REG_12__SCAN_IN | ~n42065;
  assign n41977 = ~n28403 & ~n42024;
  assign n41976 = ~n32422 & ~n42023;
  assign n41978 = ~n41977 & ~n41976;
  assign P2_U3224 = ~n41979 | ~n41978;
  assign n41981 = ~n41984 & ~n42023;
  assign n41980 = ~n32422 & ~n42024;
  assign n41983 = ~n41981 & ~n41980;
  assign n41982 = ~P2_ADDRESS_REG_13__SCAN_IN | ~n42223;
  assign P2_U3225 = ~n41983 | ~n41982;
  assign n41986 = ~n41984 & ~n42024;
  assign n41985 = ~n28422 & ~n42023;
  assign n41988 = ~n41986 & ~n41985;
  assign n41987 = ~P2_ADDRESS_REG_14__SCAN_IN | ~n42065;
  assign P2_U3226 = ~n41988 | ~n41987;
  assign n41990 = ~n28430 & ~n42023;
  assign n41989 = ~n28422 & ~n42024;
  assign n41992 = ~n41990 & ~n41989;
  assign n41991 = ~P2_ADDRESS_REG_15__SCAN_IN | ~n42065;
  assign P2_U3227 = ~n41992 | ~n41991;
  assign n41994 = ~n41997 & ~n42023;
  assign n41993 = ~n28430 & ~n42024;
  assign n41996 = ~n41994 & ~n41993;
  assign n41995 = ~P2_ADDRESS_REG_16__SCAN_IN | ~n42065;
  assign P2_U3228 = ~n41996 | ~n41995;
  assign n41999 = ~n28443 & ~n42023;
  assign n41998 = ~n41997 & ~n42024;
  assign n42001 = ~n41999 & ~n41998;
  assign n42000 = ~P2_ADDRESS_REG_17__SCAN_IN | ~n42065;
  assign P2_U3229 = ~n42001 | ~n42000;
  assign n42005 = ~P2_ADDRESS_REG_18__SCAN_IN | ~n42065;
  assign n42003 = ~n28443 & ~n42024;
  assign n42002 = ~n28450 & ~n42023;
  assign n42004 = ~n42003 & ~n42002;
  assign P2_U3230 = ~n42005 | ~n42004;
  assign n42007 = ~n28457 & ~n42023;
  assign n42006 = ~n28450 & ~n42024;
  assign n42009 = ~n42007 & ~n42006;
  assign n42008 = ~P2_ADDRESS_REG_19__SCAN_IN | ~n42065;
  assign P2_U3231 = ~n42009 | ~n42008;
  assign n42011 = ~n32310 & ~n42023;
  assign n42010 = ~n28457 & ~n42024;
  assign n42013 = ~n42011 & ~n42010;
  assign n42012 = ~P2_ADDRESS_REG_20__SCAN_IN | ~n42065;
  assign P2_U3232 = ~n42013 | ~n42012;
  assign n42015 = ~n42018 & ~n42023;
  assign n42014 = ~n32310 & ~n42024;
  assign n42017 = ~n42015 & ~n42014;
  assign n42016 = ~P2_ADDRESS_REG_21__SCAN_IN | ~n42223;
  assign P2_U3233 = ~n42017 | ~n42016;
  assign n42020 = ~n42025 & ~n42023;
  assign n42019 = ~n42018 & ~n42024;
  assign n42022 = ~n42020 & ~n42019;
  assign n42021 = ~P2_ADDRESS_REG_22__SCAN_IN | ~n42223;
  assign P2_U3234 = ~n42022 | ~n42021;
  assign n42027 = ~n42030 & ~n42023;
  assign n42026 = ~n42025 & ~n42024;
  assign n42029 = ~n42027 & ~n42026;
  assign n42028 = ~P2_ADDRESS_REG_23__SCAN_IN | ~n42223;
  assign P2_U3235 = ~n42029 | ~n42028;
  assign n42032 = ~n42035 & ~n42023;
  assign n42031 = ~n42030 & ~n42024;
  assign n42034 = ~n42032 & ~n42031;
  assign n42033 = ~P2_ADDRESS_REG_24__SCAN_IN | ~n42223;
  assign P2_U3236 = ~n42034 | ~n42033;
  assign n42037 = ~n42040 & ~n42023;
  assign n42036 = ~n42035 & ~n42024;
  assign n42039 = ~n42037 & ~n42036;
  assign n42038 = ~P2_ADDRESS_REG_25__SCAN_IN | ~n42223;
  assign P2_U3237 = ~n42039 | ~n42038;
  assign n42042 = ~n42045 & ~n42023;
  assign n42041 = ~n42040 & ~n42024;
  assign n42044 = ~n42042 & ~n42041;
  assign n42043 = ~P2_ADDRESS_REG_26__SCAN_IN | ~n42223;
  assign P2_U3238 = ~n42044 | ~n42043;
  assign n42047 = ~n42050 & ~n42023;
  assign n42046 = ~n42045 & ~n42024;
  assign n42049 = ~n42047 & ~n42046;
  assign n42048 = ~P2_ADDRESS_REG_27__SCAN_IN | ~n42223;
  assign P2_U3239 = ~n42049 | ~n42048;
  assign n42052 = ~n42056 & ~n42023;
  assign n42051 = ~n42050 & ~n42024;
  assign n42054 = ~n42052 & ~n42051;
  assign n42053 = ~P2_ADDRESS_REG_28__SCAN_IN | ~n42223;
  assign P2_U3240 = ~n42054 | ~n42053;
  assign n42058 = ~n42055 & ~n42023;
  assign n42057 = ~n42056 & ~n42024;
  assign n42060 = ~n42058 & ~n42057;
  assign n42059 = ~P2_ADDRESS_REG_29__SCAN_IN | ~n42223;
  assign P2_U3241 = ~n42060 | ~n42059;
  assign n42062 = ~n42223 | ~P2_BE_N_REG_3__SCAN_IN;
  assign n42061 = ~n42224 | ~P2_BYTEENABLE_REG_3__SCAN_IN;
  assign P2_U3585 = ~n42062 | ~n42061;
  assign n42064 = ~n42065 | ~P2_BE_N_REG_2__SCAN_IN;
  assign n42063 = ~n42224 | ~P2_BYTEENABLE_REG_2__SCAN_IN;
  assign P2_U3586 = ~n42064 | ~n42063;
  assign n42067 = ~n42065 | ~P2_BE_N_REG_1__SCAN_IN;
  assign n42066 = ~n42224 | ~P2_BYTEENABLE_REG_1__SCAN_IN;
  assign P2_U3587 = ~n42067 | ~n42066;
  assign n42069 = ~n42223 | ~P2_BE_N_REG_0__SCAN_IN;
  assign n42068 = ~n42224 | ~P2_BYTEENABLE_REG_0__SCAN_IN;
  assign P2_U3588 = ~n42069 | ~n42068;
  assign n42072 = ~n42074;
  assign n42071 = ~P2_DATAWIDTH_REG_0__SCAN_IN & ~n42070;
  assign P2_U3591 = ~n42072 & ~n42071;
  assign n42073 = ~P2_DATAWIDTH_REG_1__SCAN_IN | ~n22819;
  assign P2_U3592 = ~n42074 | ~n42073;
  assign n42078 = ~n42076 & ~n42075;
  assign n42077 = ~P2_STATE2_REG_0__SCAN_IN & ~n42196;
  assign n42081 = ~n42078 & ~n42077;
  assign n42080 = ~n42079 | ~P2_FLUSH_REG_SCAN_IN;
  assign n42132 = ~n42081 | ~n42080;
  assign n42083 = ~n42133 & ~n42137;
  assign n42085 = ~n42083 | ~n42082;
  assign n42084 = ~n42133 | ~P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN;
  assign P2_U3595 = ~n42085 | ~n42084;
  assign n42128 = ~n42111;
  assign n42088 = ~n42141 | ~n42128;
  assign n42087 = n42086 | n42137;
  assign n42089 = ~n42088 | ~n42087;
  assign n42091 = ~n42132 | ~n42089;
  assign n42090 = ~P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN | ~n42133;
  assign P2_U3596 = ~n42091 | ~n42090;
  assign n42092 = ~P2_INSTADDRPOINTER_REG_0__SCAN_IN | ~n42097;
  assign n42124 = ~n42093 | ~n42092;
  assign n42109 = ~P2_STATE2_REG_1__SCAN_IN | ~n42124;
  assign n42099 = ~n42095 | ~n42094;
  assign n42098 = ~n42097 | ~n42096;
  assign n42108 = ~n42099 | ~n42098;
  assign n42101 = ~n42109 & ~n42108;
  assign n42100 = ~n42156 & ~n42111;
  assign n42104 = ~n42101 & ~n42100;
  assign n42115 = ~n42137;
  assign n42103 = ~n42102 | ~n42115;
  assign n42105 = ~n42104 | ~n42103;
  assign n42107 = ~n42132 | ~n42105;
  assign n42106 = ~n42133 | ~P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign P2_U3599 = ~n42107 | ~n42106;
  assign n42110 = ~n42108;
  assign n42114 = ~n42110 & ~n42109;
  assign n42113 = ~n42112 & ~n42111;
  assign n42118 = ~n42114 & ~n42113;
  assign n42117 = ~n42116 | ~n42115;
  assign n42119 = ~n42118 | ~n42117;
  assign n42122 = ~n42132 | ~n42119;
  assign n42121 = ~n42133 | ~n42120;
  assign P2_U3600 = ~n42122 | ~n42121;
  assign n42127 = ~n42124 & ~n42123;
  assign n42126 = ~n42125 & ~n42137;
  assign n42130 = ~n42127 & ~n42126;
  assign n42129 = ~n42177 | ~n42128;
  assign n42131 = ~n42130 | ~n42129;
  assign n42136 = ~n42132 | ~n42131;
  assign n42135 = ~n42134 | ~n42133;
  assign P2_U3601 = ~n42136 | ~n42135;
  assign n42152 = ~P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | ~n42186;
  assign n42138 = n41002 | P2_STATEBS16_REG_SCAN_IN;
  assign n42169 = ~n42138 | ~n42137;
  assign n42146 = ~n42141 | ~n42169;
  assign n42143 = ~n42139;
  assign n42142 = ~n42141 | ~n42140;
  assign n42144 = ~n42143 | ~n42142;
  assign n42145 = ~n42144 | ~n42154;
  assign n42149 = ~n42146 | ~n42145;
  assign n42148 = ~n42147 & ~n42196;
  assign n42150 = ~n42149 & ~n42148;
  assign n42151 = n42186 | n42150;
  assign P2_U3602 = ~n42152 | ~n42151;
  assign n42185 = ~n42186;
  assign n42162 = ~n42154 | ~n42153;
  assign n42155 = ~n42154;
  assign n42168 = ~n42170 & ~n42155;
  assign n42157 = ~n42168 & ~n42169;
  assign n42160 = ~n42157 & ~n42156;
  assign n42159 = ~n42158 & ~n42196;
  assign n42161 = ~n42160 & ~n42159;
  assign n42163 = ~n42162 | ~n42161;
  assign n42165 = ~n42185 | ~n42163;
  assign n42164 = ~n42186 | ~P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign P2_U3603 = ~n42165 | ~n42164;
  assign n42167 = ~n42166 & ~n42196;
  assign n42172 = ~n42168 & ~n42167;
  assign n42171 = ~n42170 | ~n42169;
  assign n42173 = ~n42172 | ~n42171;
  assign n42175 = ~n42185 | ~n42173;
  assign n42174 = ~n42186 | ~P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN;
  assign P2_U3604 = ~n42175 | ~n42174;
  assign n42178 = n42177 & n42176;
  assign n42183 = ~n42179 & ~n42178;
  assign n42182 = ~n42181 | ~n42180;
  assign n42184 = ~n42183 | ~n42182;
  assign n42188 = ~n42185 | ~n42184;
  assign n42187 = ~n42186 | ~P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign P2_U3605 = ~n42188 | ~n42187;
  assign n42190 = ~P2_W_R_N_REG_SCAN_IN | ~n42223;
  assign n42189 = n42223 | P2_READREQUEST_REG_SCAN_IN;
  assign P2_U3608 = ~n42190 | ~n42189;
  assign n42195 = ~P2_MORE_REG_SCAN_IN | ~n42191;
  assign n42194 = ~n42193 | ~n42192;
  assign P2_U3609 = ~n42195 | ~n42194;
  assign n42198 = ~n42197 | ~n42196;
  assign n42203 = ~n42198 | ~n41002;
  assign n42201 = ~n42199 | ~n42204;
  assign n42202 = ~n42201 | ~n42200;
  assign n42220 = ~n42203 & ~n42202;
  assign n42222 = ~P2_REQUESTPENDING_REG_SCAN_IN | ~n42220;
  assign n42205 = ~n42204 | ~P2_STATE2_REG_2__SCAN_IN;
  assign n42212 = ~n42206 | ~n42205;
  assign n42207 = ~P2_STATEBS16_REG_SCAN_IN | ~n42213;
  assign n42210 = ~n42208 | ~n42207;
  assign n42211 = n42210 | n42209;
  assign n42218 = ~n42212 | ~n42211;
  assign n42215 = n42214 | n42213;
  assign n42217 = ~n42216 & ~n42215;
  assign n42219 = ~n42218 & ~n42217;
  assign n42221 = n42220 | n42219;
  assign P2_U3610 = ~n42222 | ~n42221;
  assign n42226 = ~n42223 | ~P2_M_IO_N_REG_SCAN_IN;
  assign n42225 = ~n42224 | ~P2_MEMORYFETCH_REG_SCAN_IN;
  assign P2_U3611 = ~n42226 | ~n42225;
  assign n42231 = ~n42759 & ~n42234;
  assign n42229 = ~n42228 | ~n44514;
  assign n42230 = ~P1_MEMORYFETCH_REG_SCAN_IN | ~n42229;
  assign P1_U2801 = ~n42231 | ~n42230;
  assign n42233 = ~P1_ADS_N_REG_SCAN_IN & ~n42243;
  assign P1_U2802 = ~n44859 & ~n42233;
  assign n42238 = ~P1_STATE2_REG_0__SCAN_IN | ~n42234;
  assign n42236 = ~n42235 | ~n44514;
  assign n42237 = ~P1_CODEFETCH_REG_SCAN_IN | ~n42236;
  assign P1_U2803 = ~n42238 | ~n42237;
  assign n42239 = ~P1_STATE_REG_2__SCAN_IN & ~P1_STATE_REG_0__SCAN_IN;
  assign n42240 = ~P1_D_C_N_REG_SCAN_IN & ~n42239;
  assign n42242 = ~n44859 & ~n42240;
  assign n44828 = ~n44859;
  assign n42241 = ~P1_CODEFETCH_REG_SCAN_IN & ~n44828;
  assign P1_U2804 = n42242 | n42241;
  assign n44706 = ~n44521;
  assign n44523 = ~n44546 | ~n42244;
  assign n42246 = ~n42245 | ~n44523;
  assign n44711 = ~n44706 | ~n42246;
  assign n44709 = ~n44706;
  assign n42247 = ~P1_STATEBS16_REG_SCAN_IN | ~n44709;
  assign P1_U2805 = ~n44711 | ~n42247;
  assign n44831 = ~n42248 | ~n44514;
  assign n42249 = ~P1_FLUSH_REG_SCAN_IN | ~n44831;
  assign P1_U2806 = ~n42932 | ~n42249;
  assign n42251 = ~P1_DATAWIDTH_REG_12__SCAN_IN & ~P1_DATAWIDTH_REG_13__SCAN_IN;
  assign n42250 = ~P1_DATAWIDTH_REG_14__SCAN_IN & ~P1_DATAWIDTH_REG_15__SCAN_IN;
  assign n42255 = ~n42251 | ~n42250;
  assign n42253 = ~P1_DATAWIDTH_REG_8__SCAN_IN & ~P1_DATAWIDTH_REG_9__SCAN_IN;
  assign n42252 = ~P1_DATAWIDTH_REG_10__SCAN_IN & ~P1_DATAWIDTH_REG_11__SCAN_IN;
  assign n42254 = ~n42253 | ~n42252;
  assign n42279 = ~n42255 & ~n42254;
  assign n42257 = ~P1_DATAWIDTH_REG_4__SCAN_IN & ~P1_DATAWIDTH_REG_5__SCAN_IN;
  assign n42256 = ~P1_DATAWIDTH_REG_6__SCAN_IN & ~P1_DATAWIDTH_REG_7__SCAN_IN;
  assign n42259 = ~n42257 | ~n42256;
  assign n42258 = P1_DATAWIDTH_REG_0__SCAN_IN & P1_DATAWIDTH_REG_1__SCAN_IN;
  assign n42261 = ~n42259 & ~n42258;
  assign n42260 = ~P1_DATAWIDTH_REG_2__SCAN_IN & ~P1_DATAWIDTH_REG_3__SCAN_IN;
  assign n42277 = ~n42261 | ~n42260;
  assign n42263 = ~P1_DATAWIDTH_REG_28__SCAN_IN & ~P1_DATAWIDTH_REG_29__SCAN_IN;
  assign n42262 = ~P1_DATAWIDTH_REG_30__SCAN_IN & ~P1_DATAWIDTH_REG_31__SCAN_IN;
  assign n42267 = ~n42263 | ~n42262;
  assign n42265 = ~P1_DATAWIDTH_REG_24__SCAN_IN & ~P1_DATAWIDTH_REG_25__SCAN_IN;
  assign n42264 = ~P1_DATAWIDTH_REG_26__SCAN_IN & ~P1_DATAWIDTH_REG_27__SCAN_IN;
  assign n42266 = ~n42265 | ~n42264;
  assign n42275 = ~n42267 & ~n42266;
  assign n42269 = ~P1_DATAWIDTH_REG_20__SCAN_IN & ~P1_DATAWIDTH_REG_21__SCAN_IN;
  assign n42268 = ~P1_DATAWIDTH_REG_22__SCAN_IN & ~P1_DATAWIDTH_REG_23__SCAN_IN;
  assign n42273 = ~n42269 | ~n42268;
  assign n42271 = ~P1_DATAWIDTH_REG_16__SCAN_IN & ~P1_DATAWIDTH_REG_17__SCAN_IN;
  assign n42270 = ~P1_DATAWIDTH_REG_18__SCAN_IN & ~P1_DATAWIDTH_REG_19__SCAN_IN;
  assign n42272 = ~n42271 | ~n42270;
  assign n42274 = ~n42273 & ~n42272;
  assign n42276 = ~n42275 | ~n42274;
  assign n42278 = ~n42277 & ~n42276;
  assign n44823 = ~n42279 | ~n42278;
  assign n42283 = ~P1_BYTEENABLE_REG_1__SCAN_IN | ~n44823;
  assign n44814 = ~P1_REIP_REG_0__SCAN_IN;
  assign n44813 = ~P1_DATAWIDTH_REG_0__SCAN_IN;
  assign n42280 = ~n44814 | ~n44813;
  assign n42284 = ~P1_DATAWIDTH_REG_1__SCAN_IN & ~n42280;
  assign n42281 = ~P1_REIP_REG_1__SCAN_IN & ~n42284;
  assign n42282 = n44823 | n42281;
  assign P1_U2807 = ~n42283 | ~n42282;
  assign n42287 = ~P1_BYTEENABLE_REG_3__SCAN_IN | ~n44823;
  assign n44812 = ~P1_REIP_REG_1__SCAN_IN & ~P1_DATAWIDTH_REG_1__SCAN_IN;
  assign n42285 = ~n42284 & ~n44812;
  assign n42286 = n44823 | n42285;
  assign P1_U2808 = ~n42287 | ~n42286;
  assign n42289 = ~n42481 | ~P1_EBX_REG_9__SCAN_IN;
  assign n42288 = ~n42470 | ~P1_PHYADDRPOINTER_REG_9__SCAN_IN;
  assign n42292 = ~n42289 | ~n42288;
  assign n42291 = ~n42290 & ~n22835;
  assign n42294 = ~n42292 & ~n42291;
  assign n42311 = ~n42411 | ~n42296;
  assign n42315 = ~n42469 | ~n42311;
  assign n42293 = ~P1_REIP_REG_9__SCAN_IN | ~n42315;
  assign n42295 = ~n42294 | ~n42293;
  assign n42303 = ~n42389 & ~n42295;
  assign n42301 = ~n42572 & ~n42373;
  assign n42297 = ~P1_REIP_REG_9__SCAN_IN & ~n42296;
  assign n42299 = ~n42297 | ~n42411;
  assign n42298 = ~n42512 | ~n42488;
  assign n42300 = ~n42299 | ~n42298;
  assign n42302 = ~n42301 & ~n42300;
  assign P1_U2831 = ~n42303 | ~n42302;
  assign n42305 = ~n42518 | ~n42488;
  assign n42304 = ~n42481 | ~P1_EBX_REG_8__SCAN_IN;
  assign n42310 = ~n42305 | ~n42304;
  assign n42308 = ~n42413 | ~n42306;
  assign n42307 = ~n42470 | ~P1_PHYADDRPOINTER_REG_8__SCAN_IN;
  assign n42309 = ~n42308 | ~n42307;
  assign n42321 = ~n42310 & ~n42309;
  assign n42312 = ~n42311;
  assign n42314 = ~n42313 | ~n42312;
  assign n42319 = ~n42367 | ~n42314;
  assign n42317 = ~n42579 | ~n42343;
  assign n42316 = ~P1_REIP_REG_8__SCAN_IN | ~n42315;
  assign n42318 = ~n42317 | ~n42316;
  assign n42320 = ~n42319 & ~n42318;
  assign P1_U2832 = ~n42321 | ~n42320;
  assign n42322 = ~n42411 | ~n44576;
  assign n42325 = ~n42334 & ~n42322;
  assign n42523 = ~n42323;
  assign n42324 = ~n42523 & ~n42440;
  assign n42341 = ~n42325 & ~n42324;
  assign n42339 = ~n42582 & ~n42373;
  assign n42330 = ~n42327 & ~n22835;
  assign n42329 = ~n42328 & ~n42494;
  assign n42332 = ~n42330 & ~n42329;
  assign n42331 = ~P1_EBX_REG_7__SCAN_IN | ~n42481;
  assign n42333 = ~n42332 | ~n42331;
  assign n42337 = ~n42389 & ~n42333;
  assign n42335 = ~n42411 | ~n42334;
  assign n42358 = ~n42469 | ~n42335;
  assign n42336 = ~P1_REIP_REG_7__SCAN_IN | ~n42358;
  assign n42338 = ~n42337 | ~n42336;
  assign n42340 = ~n42339 & ~n42338;
  assign P1_U2833 = ~n42341 | ~n42340;
  assign n42528 = ~n42342;
  assign n42348 = ~n42528 & ~n42440;
  assign n42344 = ~n42587;
  assign n42346 = ~n42344 | ~n42343;
  assign n42345 = ~P1_EBX_REG_6__SCAN_IN | ~n42481;
  assign n42347 = ~n42346 | ~n42345;
  assign n42349 = ~n42348 & ~n42347;
  assign n42354 = ~n42367 | ~n42349;
  assign n42352 = ~n42413 | ~n42350;
  assign n42351 = ~n42470 | ~P1_PHYADDRPOINTER_REG_6__SCAN_IN;
  assign n42353 = ~n42352 | ~n42351;
  assign n42360 = ~n42354 & ~n42353;
  assign n44571 = ~P1_REIP_REG_6__SCAN_IN;
  assign n42356 = ~n42411 | ~n42355;
  assign n42357 = ~n44571 | ~n42356;
  assign n42359 = ~n42358 | ~n42357;
  assign P1_U2834 = ~n42360 | ~n42359;
  assign n42362 = ~n42533 | ~n42488;
  assign n42361 = ~n42481 | ~P1_EBX_REG_5__SCAN_IN;
  assign n42378 = ~n42362 | ~n42361;
  assign n42365 = ~n42413 | ~n42363;
  assign n42364 = ~n42470 | ~P1_PHYADDRPOINTER_REG_5__SCAN_IN;
  assign n42370 = ~n42365 | ~n42364;
  assign n42366 = ~P1_REIP_REG_5__SCAN_IN & ~n42379;
  assign n42368 = ~n42411 | ~n42366;
  assign n42369 = ~n42368 | ~n42367;
  assign n42376 = ~n42370 & ~n42369;
  assign n42595 = ~n42371;
  assign n42374 = ~n42372 | ~n42391;
  assign n42460 = ~n42374 | ~n42373;
  assign n42375 = ~n42595 | ~n42460;
  assign n42377 = ~n42376 | ~n42375;
  assign n42381 = ~n42378 & ~n42377;
  assign n42405 = ~n42411 | ~n42379;
  assign n42401 = ~n42469 | ~n42405;
  assign n42380 = ~P1_REIP_REG_5__SCAN_IN | ~n42401;
  assign P1_U2835 = ~n42381 | ~n42380;
  assign n42383 = ~n42481 | ~P1_EBX_REG_4__SCAN_IN;
  assign n42382 = ~n42413 | ~n42894;
  assign n42398 = ~n42383 | ~n42382;
  assign n42957 = n42384 ^ n42385;
  assign n42387 = ~n42957 | ~n42488;
  assign n42386 = ~n42470 | ~P1_PHYADDRPOINTER_REG_4__SCAN_IN;
  assign n42388 = ~n42387 | ~n42386;
  assign n42396 = ~n42389 & ~n42388;
  assign n42394 = ~n42390;
  assign n42392 = ~n42391;
  assign n42484 = ~n42393 & ~n42392;
  assign n42395 = ~n42394 | ~n42484;
  assign n42397 = ~n42396 | ~n42395;
  assign n42410 = ~n42398 & ~n42397;
  assign n42903 = n42399 ^ n42400;
  assign n42403 = ~n42903 | ~n42460;
  assign n42402 = ~P1_REIP_REG_4__SCAN_IN | ~n42401;
  assign n42408 = ~n42403 | ~n42402;
  assign n42406 = ~n42404;
  assign n42407 = ~n42406 & ~n42405;
  assign n42409 = ~n42408 & ~n42407;
  assign P1_U2836 = ~n42410 | ~n42409;
  assign n44556 = ~P1_REIP_REG_3__SCAN_IN;
  assign n42416 = ~n42411 | ~P1_REIP_REG_1__SCAN_IN;
  assign n42450 = ~P1_REIP_REG_2__SCAN_IN & ~n42416;
  assign n42465 = ~n42411 | ~n44815;
  assign n42455 = ~n42469 | ~n42465;
  assign n42412 = ~n42450 & ~n42455;
  assign n42430 = ~n44556 & ~n42412;
  assign n42415 = ~n42481 | ~P1_EBX_REG_3__SCAN_IN;
  assign n42414 = ~n42413 | ~n42906;
  assign n42419 = ~n42415 | ~n42414;
  assign n44551 = ~P1_REIP_REG_2__SCAN_IN;
  assign n42417 = n42416 | n44551;
  assign n42418 = ~P1_REIP_REG_3__SCAN_IN & ~n42417;
  assign n42428 = ~n42419 & ~n42418;
  assign n42422 = n42421 | n42420;
  assign n42983 = ~n42384 | ~n42422;
  assign n42426 = ~n42983 & ~n42440;
  assign n42424 = ~n23619 | ~n42484;
  assign n42423 = ~n42470 | ~P1_PHYADDRPOINTER_REG_3__SCAN_IN;
  assign n42425 = ~n42424 | ~n42423;
  assign n42427 = ~n42426 & ~n42425;
  assign n42429 = ~n42428 | ~n42427;
  assign n42435 = ~n42430 & ~n42429;
  assign n42433 = n42432 | n42431;
  assign n42605 = ~n42399 | ~n42433;
  assign n42916 = ~n42605;
  assign n42434 = ~n42916 | ~n42460;
  assign P1_U2837 = ~n42435 | ~n42434;
  assign n42437 = ~n44784 | ~n42484;
  assign n42436 = ~n42481 | ~P1_EBX_REG_2__SCAN_IN;
  assign n42454 = ~n42437 | ~n42436;
  assign n43000 = ~n42439 ^ n42438;
  assign n42442 = ~n43000 & ~n42440;
  assign n42441 = ~n42919 & ~n22835;
  assign n42448 = ~n42442 & ~n42441;
  assign n42445 = n42444 | n42443;
  assign n42547 = n42446 & n42445;
  assign n42447 = ~n42547 | ~n42460;
  assign n42449 = ~n42448 | ~n42447;
  assign n42452 = ~n42450 & ~n42449;
  assign n42451 = ~P1_PHYADDRPOINTER_REG_2__SCAN_IN | ~n42470;
  assign n42453 = ~n42452 | ~n42451;
  assign n42457 = ~n42454 & ~n42453;
  assign n42456 = ~P1_REIP_REG_2__SCAN_IN | ~n42455;
  assign P1_U2838 = ~n42457 | ~n42456;
  assign n42478 = ~P1_PHYADDRPOINTER_REG_1__SCAN_IN & ~n42493;
  assign n42933 = ~n42459 ^ n42458;
  assign n42483 = ~n42460;
  assign n42468 = ~n42933 & ~n42483;
  assign n42463 = ~n42462 | ~n42461;
  assign n43021 = ~n42464 | ~n42463;
  assign n42466 = ~n43021 | ~n42488;
  assign n42467 = ~n42466 | ~n42465;
  assign n42476 = ~n42468 & ~n42467;
  assign n42474 = ~n42469 & ~n44815;
  assign n42472 = ~n31534 | ~n42484;
  assign n42471 = ~n42470 | ~P1_PHYADDRPOINTER_REG_1__SCAN_IN;
  assign n42473 = ~n42472 | ~n42471;
  assign n42475 = ~n42474 & ~n42473;
  assign n42477 = ~n42476 | ~n42475;
  assign n42480 = ~n42478 & ~n42477;
  assign n42479 = ~n42481 | ~P1_EBX_REG_1__SCAN_IN;
  assign P1_U2839 = ~n42480 | ~n42479;
  assign n42499 = P1_EBX_REG_0__SCAN_IN & n42481;
  assign n42952 = ~n23975 ^ n42482;
  assign n42492 = ~n42952 & ~n42483;
  assign n42490 = ~n23393 | ~n42484;
  assign n42487 = ~n42485 & ~P1_INSTADDRPOINTER_REG_0__SCAN_IN;
  assign n43036 = ~n42487 & ~n42486;
  assign n42489 = ~n43036 | ~n42488;
  assign n42491 = ~n42490 | ~n42489;
  assign n42497 = ~n42492 & ~n42491;
  assign n42495 = ~n42494 | ~n42493;
  assign n42496 = ~P1_PHYADDRPOINTER_REG_0__SCAN_IN | ~n42495;
  assign n42498 = ~n42497 | ~n42496;
  assign n42502 = ~n42499 & ~n42498;
  assign n42501 = ~P1_REIP_REG_0__SCAN_IN | ~n42500;
  assign P1_U2840 = ~n42502 | ~n42501;
  assign n42505 = ~n42503 | ~n42559;
  assign n42504 = ~P1_EBX_REG_31__SCAN_IN | ~n42556;
  assign P1_U2841 = ~n42505 | ~n42504;
  assign n42567 = ~n42506;
  assign n42509 = ~n42567 & ~n42562;
  assign n42508 = ~n42553 & ~n42507;
  assign n42511 = ~n42509 & ~n42508;
  assign n42510 = ~P1_EBX_REG_10__SCAN_IN | ~n42556;
  assign P1_U2862 = ~n42511 | ~n42510;
  assign n42515 = ~n42572 & ~n42562;
  assign n42513 = ~n42512;
  assign n42514 = ~n42553 & ~n42513;
  assign n42517 = ~n42515 & ~n42514;
  assign n42516 = ~P1_EBX_REG_9__SCAN_IN | ~n42556;
  assign P1_U2863 = ~n42517 | ~n42516;
  assign n42520 = ~n42556 | ~P1_EBX_REG_8__SCAN_IN;
  assign n42519 = ~n42559 | ~n42518;
  assign n42522 = n42520 & n42519;
  assign n42521 = ~n42579 | ~n42540;
  assign P1_U2864 = ~n42522 | ~n42521;
  assign n42525 = ~n42553 & ~n42523;
  assign n42524 = ~n42582 & ~n42562;
  assign n42527 = ~n42525 & ~n42524;
  assign n42526 = ~P1_EBX_REG_7__SCAN_IN | ~n42556;
  assign P1_U2865 = ~n42527 | ~n42526;
  assign n42530 = ~n42553 & ~n42528;
  assign n42529 = ~n42587 & ~n42562;
  assign n42532 = ~n42530 & ~n42529;
  assign n42531 = ~P1_EBX_REG_6__SCAN_IN | ~n42556;
  assign P1_U2866 = ~n42532 | ~n42531;
  assign n42535 = ~n42556 | ~P1_EBX_REG_5__SCAN_IN;
  assign n42534 = ~n42559 | ~n42533;
  assign n42537 = n42535 & n42534;
  assign n42536 = ~n42595 | ~n42540;
  assign P1_U2867 = ~n42537 | ~n42536;
  assign n42539 = ~n42556 | ~P1_EBX_REG_4__SCAN_IN;
  assign n42538 = ~n42559 | ~n42957;
  assign n42542 = n42539 & n42538;
  assign n42541 = ~n42903 | ~n42540;
  assign P1_U2868 = ~n42542 | ~n42541;
  assign n42544 = ~n42553 & ~n42983;
  assign n42543 = ~n42605 & ~n42562;
  assign n42546 = ~n42544 & ~n42543;
  assign n42545 = ~P1_EBX_REG_3__SCAN_IN | ~n42556;
  assign P1_U2869 = ~n42546 | ~n42545;
  assign n42549 = ~n42553 & ~n43000;
  assign n42922 = ~n42547;
  assign n42548 = ~n42922 & ~n42562;
  assign n42551 = ~n42549 & ~n42548;
  assign n42550 = ~P1_EBX_REG_2__SCAN_IN | ~n42556;
  assign P1_U2870 = ~n42551 | ~n42550;
  assign n42552 = ~n43021;
  assign n42555 = ~n42553 & ~n42552;
  assign n42554 = ~n42562 & ~n42933;
  assign n42558 = ~n42555 & ~n42554;
  assign n42557 = ~P1_EBX_REG_1__SCAN_IN | ~n42556;
  assign P1_U2871 = ~n42558 | ~n42557;
  assign n42566 = ~n42559 | ~n43036;
  assign n42560 = ~P1_EBX_REG_0__SCAN_IN;
  assign n42564 = ~n42561 & ~n42560;
  assign n42563 = ~n42562 & ~n42952;
  assign n42565 = ~n42564 & ~n42563;
  assign P1_U2872 = ~n42566 | ~n42565;
  assign n42569 = ~n42567 & ~n42622;
  assign n42568 = ~n42599 & ~n25989;
  assign n42571 = ~n42569 & ~n42568;
  assign n42570 = ~n42592 | ~n42800;
  assign P1_U2894 = ~n42571 | ~n42570;
  assign n42574 = ~n42572 & ~n42622;
  assign n42573 = ~n42599 & ~n25979;
  assign n42576 = ~n42574 & ~n42573;
  assign n42575 = ~n42592 | ~n42795;
  assign P1_U2895 = ~n42576 | ~n42575;
  assign n42578 = ~n42625 | ~P1_EAX_REG_8__SCAN_IN;
  assign n42577 = ~n42592 | ~n42790;
  assign n42581 = n42578 & n42577;
  assign n42580 = ~n42579 | ~n30615;
  assign P1_U2896 = ~n42581 | ~n42580;
  assign n42584 = ~n42599 & ~n25927;
  assign n42583 = ~n42582 & ~n42622;
  assign n42586 = ~n42584 & ~n42583;
  assign n42585 = ~n42592 | ~n42785;
  assign P1_U2897 = ~n42586 | ~n42585;
  assign n42589 = ~n42599 & ~n25917;
  assign n42588 = ~n42587 & ~n42622;
  assign n42591 = ~n42589 & ~n42588;
  assign n42590 = ~n42592 | ~n42781;
  assign P1_U2898 = ~n42591 | ~n42590;
  assign n42594 = ~n42625 | ~P1_EAX_REG_5__SCAN_IN;
  assign n42593 = ~n42592 | ~n42777;
  assign n42597 = n42594 & n42593;
  assign n42596 = ~n42595 | ~n30615;
  assign P1_U2899 = ~n42597 | ~n42596;
  assign n42601 = ~n42621 & ~n43152;
  assign n42600 = ~n42599 & ~n25896;
  assign n42603 = ~n42601 & ~n42600;
  assign n42602 = ~n42903 | ~n30615;
  assign P1_U2900 = ~n42603 | ~n42602;
  assign n42607 = ~n42621 & ~n43137;
  assign n42606 = ~n42605 & ~n42622;
  assign n42609 = ~n42607 & ~n42606;
  assign n42608 = ~n42625 | ~P1_EAX_REG_3__SCAN_IN;
  assign P1_U2901 = ~n42609 | ~n42608;
  assign n42612 = ~n42621 & ~n43122;
  assign n42611 = ~n42922 & ~n42622;
  assign n42614 = ~n42612 & ~n42611;
  assign n42613 = ~n42625 | ~P1_EAX_REG_2__SCAN_IN;
  assign P1_U2902 = ~n42614 | ~n42613;
  assign n42617 = ~n42621 & ~n43113;
  assign n42616 = ~n42622 & ~n42933;
  assign n42619 = ~n42617 & ~n42616;
  assign n42618 = ~n42625 | ~P1_EAX_REG_1__SCAN_IN;
  assign P1_U2903 = ~n42619 | ~n42618;
  assign n42624 = ~n42621 & ~n43070;
  assign n42623 = ~n42622 & ~n42952;
  assign n42627 = ~n42624 & ~n42623;
  assign n42626 = ~n42625 | ~P1_EAX_REG_0__SCAN_IN;
  assign P1_U2904 = ~n42627 | ~n42626;
  assign n42629 = ~n42755 | ~P1_DATAO_REG_30__SCAN_IN;
  assign n42628 = ~P1_UWORD_REG_14__SCAN_IN | ~n42746;
  assign n42633 = n42629 & n42628;
  assign n42630 = ~n42752;
  assign n42632 = ~n42631 | ~P1_EAX_REG_30__SCAN_IN;
  assign P1_U2906 = ~n42633 | ~n42632;
  assign n42635 = ~P1_DATAO_REG_29__SCAN_IN | ~n42749;
  assign n42634 = ~P1_UWORD_REG_13__SCAN_IN | ~n44835;
  assign n42637 = n42635 & n42634;
  assign n42636 = ~n42631 | ~P1_EAX_REG_29__SCAN_IN;
  assign P1_U2907 = ~n42637 | ~n42636;
  assign n42639 = ~n42755 | ~P1_DATAO_REG_28__SCAN_IN;
  assign n42638 = ~P1_UWORD_REG_12__SCAN_IN | ~n42746;
  assign n42641 = n42639 & n42638;
  assign n42640 = ~n42631 | ~P1_EAX_REG_28__SCAN_IN;
  assign P1_U2908 = ~n42641 | ~n42640;
  assign n42643 = ~P1_DATAO_REG_27__SCAN_IN | ~n42749;
  assign n42642 = ~P1_UWORD_REG_11__SCAN_IN | ~n42746;
  assign n42645 = n42643 & n42642;
  assign n42644 = ~n42631 | ~P1_EAX_REG_27__SCAN_IN;
  assign P1_U2909 = ~n42645 | ~n42644;
  assign n42647 = ~n42755 | ~P1_DATAO_REG_26__SCAN_IN;
  assign n42646 = ~P1_UWORD_REG_10__SCAN_IN | ~n42746;
  assign n42649 = n42647 & n42646;
  assign n42648 = ~n42631 | ~P1_EAX_REG_26__SCAN_IN;
  assign P1_U2910 = ~n42649 | ~n42648;
  assign n42651 = ~n42755 | ~P1_DATAO_REG_25__SCAN_IN;
  assign n42650 = ~P1_UWORD_REG_9__SCAN_IN | ~n42746;
  assign n42653 = n42651 & n42650;
  assign n42652 = ~n42631 | ~P1_EAX_REG_25__SCAN_IN;
  assign P1_U2911 = ~n42653 | ~n42652;
  assign n42655 = ~n42755 | ~P1_DATAO_REG_24__SCAN_IN;
  assign n42654 = ~P1_UWORD_REG_8__SCAN_IN | ~n42746;
  assign n42657 = n42655 & n42654;
  assign n42656 = ~n42631 | ~P1_EAX_REG_24__SCAN_IN;
  assign P1_U2912 = ~n42657 | ~n42656;
  assign n42659 = ~n42755 | ~P1_DATAO_REG_23__SCAN_IN;
  assign n42658 = ~P1_UWORD_REG_7__SCAN_IN | ~n44835;
  assign n42661 = n42659 & n42658;
  assign n42660 = ~n42631 | ~P1_EAX_REG_23__SCAN_IN;
  assign P1_U2913 = ~n42661 | ~n42660;
  assign n42663 = ~n42755 | ~P1_DATAO_REG_22__SCAN_IN;
  assign n42662 = ~P1_UWORD_REG_6__SCAN_IN | ~n44835;
  assign n42665 = n42663 & n42662;
  assign n42664 = ~n42631 | ~P1_EAX_REG_22__SCAN_IN;
  assign P1_U2914 = ~n42665 | ~n42664;
  assign n42667 = ~n42749 | ~P1_DATAO_REG_21__SCAN_IN;
  assign n42666 = ~P1_UWORD_REG_5__SCAN_IN | ~n42746;
  assign n42669 = n42667 & n42666;
  assign n42668 = ~n42631 | ~P1_EAX_REG_21__SCAN_IN;
  assign P1_U2915 = ~n42669 | ~n42668;
  assign n42671 = ~n42749 | ~P1_DATAO_REG_20__SCAN_IN;
  assign n42670 = ~P1_UWORD_REG_4__SCAN_IN | ~n42746;
  assign n42673 = n42671 & n42670;
  assign n42672 = ~n42631 | ~P1_EAX_REG_20__SCAN_IN;
  assign P1_U2916 = ~n42673 | ~n42672;
  assign n42675 = ~n42755 | ~P1_DATAO_REG_19__SCAN_IN;
  assign n42674 = ~P1_UWORD_REG_3__SCAN_IN | ~n42746;
  assign n42677 = n42675 & n42674;
  assign n42676 = ~n42631 | ~P1_EAX_REG_19__SCAN_IN;
  assign P1_U2917 = ~n42677 | ~n42676;
  assign n42679 = ~n42755 | ~P1_DATAO_REG_18__SCAN_IN;
  assign n42678 = ~P1_UWORD_REG_2__SCAN_IN | ~n44835;
  assign n42681 = n42679 & n42678;
  assign n42680 = ~n42631 | ~P1_EAX_REG_18__SCAN_IN;
  assign P1_U2918 = ~n42681 | ~n42680;
  assign n42683 = ~n42749 | ~P1_DATAO_REG_17__SCAN_IN;
  assign n42682 = ~P1_UWORD_REG_1__SCAN_IN | ~n42746;
  assign n42685 = n42683 & n42682;
  assign n42684 = ~n42631 | ~P1_EAX_REG_17__SCAN_IN;
  assign P1_U2919 = ~n42685 | ~n42684;
  assign n42687 = ~n42755 | ~P1_DATAO_REG_16__SCAN_IN;
  assign n42686 = ~P1_UWORD_REG_0__SCAN_IN | ~n42746;
  assign n42689 = n42687 & n42686;
  assign n42688 = ~n42631 | ~P1_EAX_REG_16__SCAN_IN;
  assign P1_U2920 = ~n42689 | ~n42688;
  assign n42691 = ~P1_LWORD_REG_15__SCAN_IN | ~n42746;
  assign n42690 = ~n42752 | ~P1_EAX_REG_15__SCAN_IN;
  assign n42693 = n42691 & n42690;
  assign n42692 = ~n42755 | ~P1_DATAO_REG_15__SCAN_IN;
  assign P1_U2921 = ~n42693 | ~n42692;
  assign n42695 = ~P1_LWORD_REG_14__SCAN_IN | ~n44835;
  assign n42694 = ~n42752 | ~P1_EAX_REG_14__SCAN_IN;
  assign n42697 = n42695 & n42694;
  assign n42696 = ~n42755 | ~P1_DATAO_REG_14__SCAN_IN;
  assign P1_U2922 = ~n42697 | ~n42696;
  assign n42699 = ~P1_LWORD_REG_13__SCAN_IN | ~n44835;
  assign n42698 = ~n42752 | ~P1_EAX_REG_13__SCAN_IN;
  assign n42701 = n42699 & n42698;
  assign n42700 = ~n42755 | ~P1_DATAO_REG_13__SCAN_IN;
  assign P1_U2923 = ~n42701 | ~n42700;
  assign n42703 = ~P1_LWORD_REG_12__SCAN_IN | ~n42746;
  assign n42702 = ~n42752 | ~P1_EAX_REG_12__SCAN_IN;
  assign n42705 = n42703 & n42702;
  assign n42704 = ~n42755 | ~P1_DATAO_REG_12__SCAN_IN;
  assign P1_U2924 = ~n42705 | ~n42704;
  assign n42707 = ~P1_LWORD_REG_11__SCAN_IN | ~n42746;
  assign n42706 = ~n42752 | ~P1_EAX_REG_11__SCAN_IN;
  assign n42709 = n42707 & n42706;
  assign n42708 = ~n42755 | ~P1_DATAO_REG_11__SCAN_IN;
  assign P1_U2925 = ~n42709 | ~n42708;
  assign n42711 = ~P1_LWORD_REG_10__SCAN_IN | ~n42746;
  assign n42710 = ~n42752 | ~P1_EAX_REG_10__SCAN_IN;
  assign n42713 = n42711 & n42710;
  assign n42712 = ~n42749 | ~P1_DATAO_REG_10__SCAN_IN;
  assign P1_U2926 = ~n42713 | ~n42712;
  assign n42715 = ~P1_LWORD_REG_9__SCAN_IN | ~n44835;
  assign n42714 = ~n42752 | ~P1_EAX_REG_9__SCAN_IN;
  assign n42717 = n42715 & n42714;
  assign n42716 = ~n42749 | ~P1_DATAO_REG_9__SCAN_IN;
  assign P1_U2927 = ~n42717 | ~n42716;
  assign n42719 = ~P1_LWORD_REG_8__SCAN_IN | ~n42746;
  assign n42718 = ~n42752 | ~P1_EAX_REG_8__SCAN_IN;
  assign n42721 = n42719 & n42718;
  assign n42720 = ~n42749 | ~P1_DATAO_REG_8__SCAN_IN;
  assign P1_U2928 = ~n42721 | ~n42720;
  assign n42723 = ~P1_LWORD_REG_7__SCAN_IN | ~n42746;
  assign n42722 = ~n42752 | ~P1_EAX_REG_7__SCAN_IN;
  assign n42725 = n42723 & n42722;
  assign n42724 = ~n42749 | ~P1_DATAO_REG_7__SCAN_IN;
  assign P1_U2929 = ~n42725 | ~n42724;
  assign n42727 = ~P1_LWORD_REG_6__SCAN_IN | ~n42746;
  assign n42726 = ~n42752 | ~P1_EAX_REG_6__SCAN_IN;
  assign n42729 = n42727 & n42726;
  assign n42728 = ~n42749 | ~P1_DATAO_REG_6__SCAN_IN;
  assign P1_U2930 = ~n42729 | ~n42728;
  assign n42731 = ~P1_LWORD_REG_5__SCAN_IN | ~n44835;
  assign n42730 = ~n42752 | ~P1_EAX_REG_5__SCAN_IN;
  assign n42733 = n42731 & n42730;
  assign n42732 = ~n42749 | ~P1_DATAO_REG_5__SCAN_IN;
  assign P1_U2931 = ~n42733 | ~n42732;
  assign n42735 = ~P1_LWORD_REG_4__SCAN_IN | ~n44835;
  assign n42734 = ~n42752 | ~P1_EAX_REG_4__SCAN_IN;
  assign n42737 = n42735 & n42734;
  assign n42736 = ~n42749 | ~P1_DATAO_REG_4__SCAN_IN;
  assign P1_U2932 = ~n42737 | ~n42736;
  assign n42739 = ~P1_LWORD_REG_3__SCAN_IN | ~n42746;
  assign n42738 = ~n42752 | ~P1_EAX_REG_3__SCAN_IN;
  assign n42741 = n42739 & n42738;
  assign n42740 = ~n42749 | ~P1_DATAO_REG_3__SCAN_IN;
  assign P1_U2933 = ~n42741 | ~n42740;
  assign n42743 = ~P1_LWORD_REG_2__SCAN_IN | ~n42746;
  assign n42742 = ~n42752 | ~P1_EAX_REG_2__SCAN_IN;
  assign n42745 = n42743 & n42742;
  assign n42744 = ~n42749 | ~P1_DATAO_REG_2__SCAN_IN;
  assign P1_U2934 = ~n42745 | ~n42744;
  assign n42748 = ~P1_LWORD_REG_1__SCAN_IN | ~n42746;
  assign n42747 = ~n42752 | ~P1_EAX_REG_1__SCAN_IN;
  assign n42751 = n42748 & n42747;
  assign n42750 = ~n42749 | ~P1_DATAO_REG_1__SCAN_IN;
  assign P1_U2935 = ~n42751 | ~n42750;
  assign n42754 = ~P1_LWORD_REG_0__SCAN_IN | ~n44835;
  assign n42753 = ~n42752 | ~P1_EAX_REG_0__SCAN_IN;
  assign n42757 = n42754 & n42753;
  assign n42756 = ~n42755 | ~P1_DATAO_REG_0__SCAN_IN;
  assign P1_U2936 = ~n42757 | ~n42756;
  assign n42888 = ~n42761 | ~n42760;
  assign n42824 = ~n42888 & ~n43070;
  assign n42762 = ~n42855 & ~n26225;
  assign n42764 = ~n42824 & ~n42762;
  assign n42763 = ~P1_UWORD_REG_0__SCAN_IN | ~n42891;
  assign P1_U2937 = ~n42764 | ~n42763;
  assign n42828 = ~n42888 & ~n43113;
  assign n42765 = ~n42855 & ~n26266;
  assign n42767 = ~n42828 & ~n42765;
  assign n42766 = ~P1_UWORD_REG_1__SCAN_IN | ~n42891;
  assign P1_U2938 = ~n42767 | ~n42766;
  assign n42832 = ~n42888 & ~n43122;
  assign n42768 = ~n42855 & ~n26309;
  assign n42770 = ~n42832 & ~n42768;
  assign n42769 = ~P1_UWORD_REG_2__SCAN_IN | ~n42891;
  assign P1_U2939 = ~n42770 | ~n42769;
  assign n42836 = ~n42888 & ~n43137;
  assign n42771 = ~n42855 & ~n26471;
  assign n42773 = ~n42836 & ~n42771;
  assign n42772 = ~P1_UWORD_REG_3__SCAN_IN | ~n42891;
  assign P1_U2940 = ~n42773 | ~n42772;
  assign n42840 = ~n42888 & ~n43152;
  assign n42774 = ~n42855 & ~n26558;
  assign n42776 = ~n42840 & ~n42774;
  assign n42775 = ~P1_UWORD_REG_4__SCAN_IN | ~n42891;
  assign P1_U2941 = ~n42776 | ~n42775;
  assign n43173 = ~n42777;
  assign n42844 = ~n42888 & ~n43173;
  assign n42778 = ~n42855 & ~n26431;
  assign n42780 = ~n42844 & ~n42778;
  assign n42779 = ~P1_UWORD_REG_5__SCAN_IN | ~n42891;
  assign P1_U2942 = ~n42780 | ~n42779;
  assign n43187 = ~n42781;
  assign n42848 = ~n42888 & ~n43187;
  assign n42782 = ~n42855 & ~n26601;
  assign n42784 = ~n42848 & ~n42782;
  assign n42783 = ~P1_UWORD_REG_6__SCAN_IN | ~n42891;
  assign P1_U2943 = ~n42784 | ~n42783;
  assign n43197 = ~n42785;
  assign n42852 = ~n42888 & ~n43197;
  assign n42786 = ~P1_EAX_REG_23__SCAN_IN;
  assign n42787 = ~n42855 & ~n42786;
  assign n42789 = ~n42852 & ~n42787;
  assign n42788 = ~P1_UWORD_REG_7__SCAN_IN | ~n42891;
  assign P1_U2944 = ~n42789 | ~n42788;
  assign n42791 = ~n42790;
  assign n42857 = ~n42888 & ~n42791;
  assign n42792 = ~n42855 & ~n26516;
  assign n42794 = ~n42857 & ~n42792;
  assign n42793 = ~P1_UWORD_REG_8__SCAN_IN | ~n42891;
  assign P1_U2945 = ~n42794 | ~n42793;
  assign n42796 = ~n42795;
  assign n42861 = ~n42888 & ~n42796;
  assign n42797 = ~n42855 & ~n26650;
  assign n42799 = ~n42861 & ~n42797;
  assign n42798 = ~P1_UWORD_REG_9__SCAN_IN | ~n42891;
  assign P1_U2946 = ~n42799 | ~n42798;
  assign n42801 = ~n42800;
  assign n42865 = ~n42888 & ~n42801;
  assign n42802 = ~n42855 & ~n26696;
  assign n42804 = ~n42865 & ~n42802;
  assign n42803 = ~P1_UWORD_REG_10__SCAN_IN | ~n42891;
  assign P1_U2947 = ~n42804 | ~n42803;
  assign n42806 = ~n42805;
  assign n42869 = ~n42888 & ~n42806;
  assign n42807 = ~n42855 & ~n26739;
  assign n42809 = ~n42869 & ~n42807;
  assign n42808 = ~P1_UWORD_REG_11__SCAN_IN | ~n42891;
  assign P1_U2948 = ~n42809 | ~n42808;
  assign n42874 = ~n42888 & ~n42810;
  assign n42811 = ~n42855 & ~n26788;
  assign n42813 = ~n42874 & ~n42811;
  assign n42812 = ~P1_UWORD_REG_12__SCAN_IN | ~n42891;
  assign P1_U2949 = ~n42813 | ~n42812;
  assign n42879 = ~n42888 & ~n42814;
  assign n42815 = ~n42855 & ~n26836;
  assign n42817 = ~n42879 & ~n42815;
  assign n42816 = ~P1_UWORD_REG_13__SCAN_IN | ~n42891;
  assign P1_U2950 = ~n42817 | ~n42816;
  assign n42819 = ~n42818;
  assign n42884 = ~n42888 & ~n42819;
  assign n42820 = ~n42855 & ~n26892;
  assign n42822 = ~n42884 & ~n42820;
  assign n42821 = ~P1_UWORD_REG_14__SCAN_IN | ~n42891;
  assign P1_U2951 = ~n42822 | ~n42821;
  assign n42823 = ~n42855 & ~n25870;
  assign n42826 = ~n42824 & ~n42823;
  assign n42825 = ~P1_LWORD_REG_0__SCAN_IN | ~n42891;
  assign P1_U2952 = ~n42826 | ~n42825;
  assign n42827 = ~n42855 & ~n25861;
  assign n42830 = ~n42828 & ~n42827;
  assign n42829 = ~P1_LWORD_REG_1__SCAN_IN | ~n42891;
  assign P1_U2953 = ~n42830 | ~n42829;
  assign n42831 = ~n42855 & ~n25851;
  assign n42834 = ~n42832 & ~n42831;
  assign n42833 = ~P1_LWORD_REG_2__SCAN_IN | ~n42891;
  assign P1_U2954 = ~n42834 | ~n42833;
  assign n42835 = ~n42855 & ~n25886;
  assign n42838 = ~n42836 & ~n42835;
  assign n42837 = ~P1_LWORD_REG_3__SCAN_IN | ~n42891;
  assign P1_U2955 = ~n42838 | ~n42837;
  assign n42839 = ~n42855 & ~n25896;
  assign n42842 = ~n42840 & ~n42839;
  assign n42841 = ~P1_LWORD_REG_4__SCAN_IN | ~n42891;
  assign P1_U2956 = ~n42842 | ~n42841;
  assign n42843 = ~n42855 & ~n25909;
  assign n42846 = ~n42844 & ~n42843;
  assign n42845 = ~P1_LWORD_REG_5__SCAN_IN | ~n42891;
  assign P1_U2957 = ~n42846 | ~n42845;
  assign n42847 = ~n42855 & ~n25917;
  assign n42850 = ~n42848 & ~n42847;
  assign n42849 = ~P1_LWORD_REG_6__SCAN_IN | ~n42891;
  assign P1_U2958 = ~n42850 | ~n42849;
  assign n42851 = ~n42855 & ~n25927;
  assign n42854 = ~n42852 & ~n42851;
  assign n42853 = ~P1_LWORD_REG_7__SCAN_IN | ~n42891;
  assign P1_U2959 = ~n42854 | ~n42853;
  assign n42856 = ~n42855 & ~n25937;
  assign n42859 = ~n42857 & ~n42856;
  assign n42858 = ~P1_LWORD_REG_8__SCAN_IN | ~n42891;
  assign P1_U2960 = ~n42859 | ~n42858;
  assign n42860 = ~n42855 & ~n25979;
  assign n42863 = ~n42861 & ~n42860;
  assign n42862 = ~P1_LWORD_REG_9__SCAN_IN | ~n42891;
  assign P1_U2961 = ~n42863 | ~n42862;
  assign n42864 = ~n42855 & ~n25989;
  assign n42867 = ~n42865 & ~n42864;
  assign n42866 = ~P1_LWORD_REG_10__SCAN_IN | ~n42891;
  assign P1_U2962 = ~n42867 | ~n42866;
  assign n42868 = ~n42855 & ~n26067;
  assign n42871 = ~n42869 & ~n42868;
  assign n42870 = ~P1_LWORD_REG_11__SCAN_IN | ~n42891;
  assign P1_U2963 = ~n42871 | ~n42870;
  assign n42873 = ~n42855 & ~n42872;
  assign n42876 = ~n42874 & ~n42873;
  assign n42875 = ~P1_LWORD_REG_12__SCAN_IN | ~n42891;
  assign P1_U2964 = ~n42876 | ~n42875;
  assign n42878 = ~n42855 & ~n42877;
  assign n42881 = ~n42879 & ~n42878;
  assign n42880 = ~P1_LWORD_REG_13__SCAN_IN | ~n42891;
  assign P1_U2965 = ~n42881 | ~n42880;
  assign n42883 = ~n42855 & ~n42882;
  assign n42886 = ~n42884 & ~n42883;
  assign n42885 = ~P1_LWORD_REG_14__SCAN_IN | ~n42891;
  assign P1_U2966 = ~n42886 | ~n42885;
  assign n42890 = ~n42888 & ~n42887;
  assign n42889 = ~n42855 & ~n30606;
  assign n42893 = ~n42890 & ~n42889;
  assign n42892 = ~P1_LWORD_REG_15__SCAN_IN | ~n42891;
  assign P1_U2967 = ~n42893 | ~n42892;
  assign n42897 = ~n42895 | ~n42894;
  assign n42896 = ~n42937 | ~P1_PHYADDRPOINTER_REG_4__SCAN_IN;
  assign n42902 = ~n42897 | ~n42896;
  assign n42958 = ~n42929 | ~P1_REIP_REG_4__SCAN_IN;
  assign n42978 = n23083 ^ n42898;
  assign n42900 = ~n42978 | ~n42949;
  assign n42901 = ~n42958 | ~n42900;
  assign n42905 = ~n42902 & ~n42901;
  assign n42904 = ~n42903 | ~n42915;
  assign P1_U2995 = ~n42905 | ~n42904;
  assign n42909 = ~n42907 | ~n42906;
  assign n42908 = ~n42937 | ~P1_PHYADDRPOINTER_REG_3__SCAN_IN;
  assign n42914 = ~n42909 | ~n42908;
  assign n42985 = ~n42947 & ~n44556;
  assign n42912 = ~n42985;
  assign n42982 = n31012 ^ n42910;
  assign n42911 = ~n42982 | ~n42949;
  assign n42913 = ~n42912 | ~n42911;
  assign n42918 = ~n42914 & ~n42913;
  assign n42917 = ~n42916 | ~n42915;
  assign P1_U2996 = ~n42918 | ~n42917;
  assign n42928 = ~n42919 & ~n42936;
  assign n43008 = ~n42920 ^ n42921;
  assign n42924 = ~n43008 & ~n42932;
  assign n42923 = ~n42922 & ~n43061;
  assign n42926 = ~n42924 & ~n42923;
  assign n42925 = ~P1_PHYADDRPOINTER_REG_2__SCAN_IN | ~n42937;
  assign n42927 = ~n42926 | ~n42925;
  assign n42930 = ~n42928 & ~n42927;
  assign n43002 = ~n42929 | ~P1_REIP_REG_2__SCAN_IN;
  assign P1_U2997 = ~n42930 | ~n43002;
  assign n43017 = ~n42931 ^ n25405;
  assign n42935 = ~n42932 & ~n43017;
  assign n42934 = ~n42933 & ~n43061;
  assign n42943 = ~n42935 & ~n42934;
  assign n42941 = ~P1_PHYADDRPOINTER_REG_1__SCAN_IN & ~n42936;
  assign n43019 = ~n42947 & ~n44815;
  assign n42939 = ~n43019;
  assign n42938 = ~n42937 | ~P1_PHYADDRPOINTER_REG_1__SCAN_IN;
  assign n42940 = ~n42939 | ~n42938;
  assign n42942 = ~n42941 & ~n42940;
  assign P1_U2998 = ~n42943 | ~n42942;
  assign n42946 = ~n42945 | ~n42944;
  assign n42956 = ~n42946 | ~P1_PHYADDRPOINTER_REG_0__SCAN_IN;
  assign n43035 = ~n42947 & ~n44814;
  assign n42951 = ~n43035;
  assign n43041 = P1_INSTADDRPOINTER_REG_0__SCAN_IN ^ n42948;
  assign n42950 = ~n42949 | ~n43041;
  assign n42954 = ~n42951 | ~n42950;
  assign n42953 = ~n42952 & ~n43061;
  assign n42955 = ~n42954 & ~n42953;
  assign P1_U2999 = ~n42956 | ~n42955;
  assign n42959 = ~n25838 | ~n42957;
  assign n42977 = ~n42959 | ~n42958;
  assign n42998 = ~P1_INSTADDRPOINTER_REG_2__SCAN_IN & ~n42960;
  assign n42962 = ~n25405 | ~n42961;
  assign n42994 = ~n42963 | ~n42962;
  assign n42964 = ~n42998 & ~n42994;
  assign n43003 = ~n43014 | ~n42965;
  assign n42990 = ~n42964 | ~n43003;
  assign n42975 = ~P1_INSTADDRPOINTER_REG_4__SCAN_IN | ~n42990;
  assign n42970 = ~n42966 & ~n42965;
  assign n42969 = ~n42968 & ~n42967;
  assign n42981 = ~n42970 & ~n42969;
  assign n42971 = ~P1_INSTADDRPOINTER_REG_4__SCAN_IN & ~P1_INSTADDRPOINTER_REG_3__SCAN_IN;
  assign n42973 = ~n42981 & ~n42971;
  assign n42974 = ~n42973 | ~n42972;
  assign n42976 = ~n42975 | ~n42974;
  assign n42980 = ~n42977 & ~n42976;
  assign n42979 = ~n42978 | ~n43042;
  assign P1_U3027 = ~n42980 | ~n42979;
  assign n42989 = ~P1_INSTADDRPOINTER_REG_3__SCAN_IN & ~n42981;
  assign n42987 = ~n42982 | ~n43042;
  assign n42984 = ~n43001 & ~n42983;
  assign n42986 = ~n42985 & ~n42984;
  assign n42988 = ~n42987 | ~n42986;
  assign n42992 = ~n42989 & ~n42988;
  assign n42991 = ~P1_INSTADDRPOINTER_REG_3__SCAN_IN | ~n42990;
  assign P1_U3028 = ~n42992 | ~n42991;
  assign n42996 = ~n43014 | ~n42993;
  assign n42995 = ~n42994;
  assign n42997 = ~n42996 | ~n42995;
  assign n43012 = ~n42997 | ~P1_INSTADDRPOINTER_REG_2__SCAN_IN;
  assign n42999 = ~n25405 & ~n43026;
  assign n43007 = ~n42999 | ~n42998;
  assign n43005 = ~n43001 & ~n43000;
  assign n43004 = ~n43003 | ~n43002;
  assign n43006 = ~n43005 & ~n43004;
  assign n43010 = ~n43007 | ~n43006;
  assign n43009 = ~n43018 & ~n43008;
  assign n43011 = ~n43010 & ~n43009;
  assign P1_U3029 = ~n43012 | ~n43011;
  assign n43015 = ~n43014 & ~n43013;
  assign n43040 = ~P1_INSTADDRPOINTER_REG_0__SCAN_IN & ~n43015;
  assign n43016 = ~n43032 & ~n43040;
  assign n43025 = ~n43016 & ~n25405;
  assign n43020 = ~n43018 & ~n43017;
  assign n43023 = ~n43020 & ~n43019;
  assign n43022 = ~n25838 | ~n43021;
  assign n43024 = ~n43023 | ~n43022;
  assign n43030 = ~n43025 & ~n43024;
  assign n43028 = ~n43027 & ~n43026;
  assign n43029 = ~n43028 | ~n25405;
  assign P1_U3030 = ~n43030 | ~n43029;
  assign n43033 = ~n43032 & ~n43031;
  assign n43034 = ~n44753 & ~n43033;
  assign n43038 = ~n43035 & ~n43034;
  assign n43037 = ~n43036 | ~n25838;
  assign n43039 = ~n43038 | ~n43037;
  assign n43044 = ~n43040 & ~n43039;
  assign n43043 = ~n43042 | ~n43041;
  assign P1_U3031 = ~n43044 | ~n43043;
  assign n43045 = ~n24764;
  assign n43048 = ~n43046 | ~n43045;
  assign n44509 = ~n43048 | ~n43047;
  assign n43050 = ~P1_FLUSH_REG_SCAN_IN & ~n44509;
  assign n43052 = ~n44508 | ~n44853;
  assign n44808 = ~n43054 | ~n43471;
  assign P1_U3032 = ~n43055 & ~n44808;
  assign n43058 = ~n43191 & ~n43057;
  assign n43294 = ~P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & ~P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign n43059 = ~n43294;
  assign n43221 = ~P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN & ~n43059;
  assign n43087 = ~n43221 | ~n44308;
  assign n43192 = ~n43087;
  assign n43069 = ~n44394 | ~n43192;
  assign n43064 = ~n43199 | ~DATAI_24_;
  assign n43200 = ~n43062 & ~n43061;
  assign n43063 = ~n43200 | ~BUF1_REG_24__SCAN_IN;
  assign n44411 = ~n43065 & ~n44781;
  assign n44317 = ~n44411 | ~n43066;
  assign n43068 = ~n44406 | ~n43067;
  assign n43096 = ~n43069 | ~n43068;
  assign n44402 = ~n43471 & ~n43070;
  assign n43470 = ~n43081 & ~n43082;
  assign n43977 = ~n43470;
  assign n43071 = ~n43977 & ~n44153;
  assign n43080 = ~n43071 | ~n44152;
  assign n43075 = ~n43067;
  assign n43073 = ~n44781 | ~n44792;
  assign n43285 = ~n43225 & ~n44801;
  assign n43074 = ~n43285;
  assign n43076 = ~n43075 | ~n43074;
  assign n43077 = ~n43076 | ~P1_STATEBS16_REG_SCAN_IN;
  assign n43085 = ~n43077 | ~n44800;
  assign n43078 = ~n43085;
  assign n43084 = ~n43380 & ~n31534;
  assign n43079 = ~n43078 | ~n43084;
  assign n43094 = ~n44402 | ~n43198;
  assign n43083 = ~n43081;
  assign n43636 = ~n43083 & ~n43082;
  assign n43091 = ~n43085 & ~n43084;
  assign n44136 = ~n44153;
  assign n43086 = ~n44136 | ~n44152;
  assign n43089 = ~n43086 | ~P1_STATE2_REG_2__SCAN_IN;
  assign n43088 = ~n43087 | ~P1_STATE2_REG_3__SCAN_IN;
  assign n43090 = ~n43089 | ~n43088;
  assign n43092 = ~n43091 & ~n43090;
  assign n43093 = ~P1_INSTQUEUE_REG_0__0__SCAN_IN | ~n43207;
  assign n43095 = ~n43094 | ~n43093;
  assign n43100 = ~n43096 & ~n43095;
  assign n43098 = ~n43199 | ~DATAI_16_;
  assign n43097 = ~n43200 | ~BUF1_REG_16__SCAN_IN;
  assign n43099 = ~n44405 | ~n43285;
  assign P1_U3033 = ~n43100 | ~n43099;
  assign n43106 = ~n43102 | ~n43192;
  assign n43104 = ~n43200 | ~BUF1_REG_25__SCAN_IN;
  assign n43103 = ~n43199 | ~DATAI_25_;
  assign n44428 = ~n43104 | ~n43103;
  assign n43105 = ~n44428 | ~n43067;
  assign n43112 = ~n43106 | ~n43105;
  assign n43110 = ~P1_INSTQUEUE_REG_0__1__SCAN_IN | ~n43207;
  assign n43108 = ~n43199 | ~DATAI_17_;
  assign n43107 = ~n43200 | ~BUF1_REG_17__SCAN_IN;
  assign n44427 = ~n43108 | ~n43107;
  assign n43109 = ~n44427 | ~n43285;
  assign n43111 = ~n43110 | ~n43109;
  assign n43115 = ~n43112 & ~n43111;
  assign n44424 = ~n43471 & ~n43113;
  assign n43114 = ~n44424 | ~n43198;
  assign P1_U3034 = ~n43115 | ~n43114;
  assign n43121 = ~n43117 | ~n43192;
  assign n43119 = ~n43200 | ~BUF1_REG_26__SCAN_IN;
  assign n43118 = ~n43199 | ~DATAI_26_;
  assign n44439 = ~n43119 | ~n43118;
  assign n43120 = ~n44439 | ~n43067;
  assign n43128 = ~n43121 | ~n43120;
  assign n44435 = ~n43471 & ~n43122;
  assign n43126 = ~n44435 | ~n43198;
  assign n43124 = ~n43199 | ~DATAI_18_;
  assign n43123 = ~n43200 | ~BUF1_REG_18__SCAN_IN;
  assign n44438 = ~n43124 | ~n43123;
  assign n43125 = ~n44438 | ~n43285;
  assign n43127 = ~n43126 | ~n43125;
  assign n43130 = ~n43128 & ~n43127;
  assign n43129 = ~P1_INSTQUEUE_REG_0__2__SCAN_IN | ~n43207;
  assign P1_U3035 = ~n43130 | ~n43129;
  assign n43136 = ~n43132 | ~n43192;
  assign n43134 = ~n43199 | ~DATAI_27_;
  assign n43133 = ~n43200 | ~BUF1_REG_27__SCAN_IN;
  assign n44450 = ~n43134 | ~n43133;
  assign n43135 = ~n44450 | ~n43067;
  assign n43143 = ~n43136 | ~n43135;
  assign n44446 = ~n43471 & ~n43137;
  assign n43141 = ~n44446 | ~n43198;
  assign n43139 = ~n43200 | ~BUF1_REG_19__SCAN_IN;
  assign n43138 = ~n43199 | ~DATAI_19_;
  assign n44449 = ~n43139 | ~n43138;
  assign n43140 = ~n44449 | ~n43285;
  assign n43142 = ~n43141 | ~n43140;
  assign n43145 = ~n43143 & ~n43142;
  assign n43144 = ~P1_INSTQUEUE_REG_0__3__SCAN_IN | ~n43207;
  assign P1_U3036 = ~n43145 | ~n43144;
  assign n43151 = ~n43147 | ~n43192;
  assign n43149 = ~n43199 | ~DATAI_28_;
  assign n43148 = ~n43200 | ~BUF1_REG_28__SCAN_IN;
  assign n44461 = ~n43149 | ~n43148;
  assign n43150 = ~n44461 | ~n43067;
  assign n43158 = ~n43151 | ~n43150;
  assign n44457 = ~n43471 & ~n43152;
  assign n43156 = ~n44457 | ~n43198;
  assign n43154 = ~n43200 | ~BUF1_REG_20__SCAN_IN;
  assign n43153 = ~n43199 | ~DATAI_20_;
  assign n44460 = ~n43154 | ~n43153;
  assign n43155 = ~n44460 | ~n43285;
  assign n43157 = ~n43156 | ~n43155;
  assign n43160 = ~n43158 & ~n43157;
  assign n43159 = ~P1_INSTQUEUE_REG_0__4__SCAN_IN | ~n43207;
  assign P1_U3037 = ~n43160 | ~n43159;
  assign n43162 = ~n43191 & ~n43161;
  assign n43166 = ~n44468 | ~n43192;
  assign n43164 = ~n43199 | ~DATAI_29_;
  assign n43163 = ~n43200 | ~BUF1_REG_29__SCAN_IN;
  assign n44473 = ~n43164 | ~n43163;
  assign n43165 = ~n44473 | ~n43067;
  assign n43172 = ~n43166 | ~n43165;
  assign n43170 = ~P1_INSTQUEUE_REG_0__5__SCAN_IN | ~n43207;
  assign n43168 = ~n43200 | ~BUF1_REG_21__SCAN_IN;
  assign n43167 = ~n43199 | ~DATAI_21_;
  assign n44472 = ~n43168 | ~n43167;
  assign n43169 = ~n44472 | ~n43285;
  assign n43171 = ~n43170 | ~n43169;
  assign n43175 = ~n43172 & ~n43171;
  assign n44469 = ~n43471 & ~n43173;
  assign n43174 = ~n44469 | ~n43198;
  assign P1_U3038 = ~n43175 | ~n43174;
  assign n43180 = ~n22825 | ~n43192;
  assign n43178 = ~n43199 | ~DATAI_30_;
  assign n43177 = ~n43200 | ~BUF1_REG_30__SCAN_IN;
  assign n44484 = ~n43178 | ~n43177;
  assign n43179 = ~n44484 | ~n43067;
  assign n43186 = ~n43180 | ~n43179;
  assign n43184 = ~P1_INSTQUEUE_REG_0__6__SCAN_IN | ~n43207;
  assign n43182 = ~n43200 | ~BUF1_REG_22__SCAN_IN;
  assign n43181 = ~n43199 | ~DATAI_22_;
  assign n44483 = ~n43182 | ~n43181;
  assign n43183 = ~n44483 | ~n43285;
  assign n43185 = ~n43184 | ~n43183;
  assign n43189 = ~n43186 & ~n43185;
  assign n44480 = ~n43471 & ~n43187;
  assign n43188 = ~n44480 | ~n43198;
  assign P1_U3039 = ~n43189 | ~n43188;
  assign n44492 = ~n43191 & ~n43190;
  assign n43196 = ~n44492 | ~n43192;
  assign n43194 = ~n43200 | ~BUF1_REG_31__SCAN_IN;
  assign n43193 = ~n43199 | ~DATAI_31_;
  assign n44500 = ~n43194 | ~n43193;
  assign n43195 = ~n44500 | ~n43067;
  assign n43206 = ~n43196 | ~n43195;
  assign n44494 = ~n43471 & ~n43197;
  assign n43204 = ~n44494 | ~n43198;
  assign n43202 = ~n43199 | ~DATAI_23_;
  assign n43201 = ~n43200 | ~BUF1_REG_23__SCAN_IN;
  assign n44498 = ~n43202 | ~n43201;
  assign n43203 = ~n44498 | ~n43285;
  assign n43205 = ~n43204 | ~n43203;
  assign n43209 = ~n43206 & ~n43205;
  assign n43208 = ~P1_INSTQUEUE_REG_0__7__SCAN_IN | ~n43207;
  assign P1_U3040 = ~n43209 | ~n43208;
  assign n43215 = ~n44394 | ~n43281;
  assign n43211 = ~n43380 & ~n43880;
  assign n43216 = n43211 | n43281;
  assign n43213 = ~n43216 | ~n44800;
  assign n43212 = ~n43221 | ~P1_STATE2_REG_2__SCAN_IN;
  assign n43282 = ~n43213 | ~n43212;
  assign n43214 = ~n44402 | ~n43282;
  assign n43230 = ~n43215 | ~n43214;
  assign n43218 = ~n43225 & ~n44765;
  assign n43217 = n43216 | n44418;
  assign n43220 = ~n43218 & ~n43217;
  assign n43219 = ~n44766 & ~P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n43224 = ~n43220 & ~n44415;
  assign n43222 = ~n43221;
  assign n43223 = ~n44418 | ~n43222;
  assign n43228 = ~P1_INSTQUEUE_REG_1__0__SCAN_IN | ~n43290;
  assign n43226 = ~n43225 & ~n44230;
  assign n43372 = n43226;
  assign n43227 = ~n44405 | ~n43372;
  assign n43229 = ~n43228 | ~n43227;
  assign n43232 = ~n43230 & ~n43229;
  assign n43231 = ~n44406 | ~n43285;
  assign P1_U3041 = ~n43232 | ~n43231;
  assign n43234 = ~n43102 | ~n43281;
  assign n43233 = ~n44424 | ~n43282;
  assign n43238 = ~n43234 | ~n43233;
  assign n43236 = ~n44427 | ~n43372;
  assign n43235 = ~n44428 | ~n43285;
  assign n43237 = ~n43236 | ~n43235;
  assign n43240 = ~n43238 & ~n43237;
  assign n43239 = ~P1_INSTQUEUE_REG_1__1__SCAN_IN | ~n43290;
  assign P1_U3042 = ~n43240 | ~n43239;
  assign n43242 = ~n43117 | ~n43281;
  assign n43241 = ~n44435 | ~n43282;
  assign n43246 = ~n43242 | ~n43241;
  assign n43244 = ~n44438 | ~n43372;
  assign n43243 = ~n44439 | ~n43285;
  assign n43245 = ~n43244 | ~n43243;
  assign n43248 = ~n43246 & ~n43245;
  assign n43247 = ~P1_INSTQUEUE_REG_1__2__SCAN_IN | ~n43290;
  assign P1_U3043 = ~n43248 | ~n43247;
  assign n43250 = ~n43132 | ~n43281;
  assign n43249 = ~n44446 | ~n43282;
  assign n43254 = ~n43250 | ~n43249;
  assign n43252 = ~n44449 | ~n43372;
  assign n43251 = ~n44450 | ~n43285;
  assign n43253 = ~n43252 | ~n43251;
  assign n43256 = ~n43254 & ~n43253;
  assign n43255 = ~P1_INSTQUEUE_REG_1__3__SCAN_IN | ~n43290;
  assign P1_U3044 = ~n43256 | ~n43255;
  assign n43258 = ~n43147 | ~n43281;
  assign n43257 = ~n44457 | ~n43282;
  assign n43262 = ~n43258 | ~n43257;
  assign n43260 = ~n44460 | ~n43372;
  assign n43259 = ~n44461 | ~n43285;
  assign n43261 = ~n43260 | ~n43259;
  assign n43264 = ~n43262 & ~n43261;
  assign n43263 = ~P1_INSTQUEUE_REG_1__4__SCAN_IN | ~n43290;
  assign P1_U3045 = ~n43264 | ~n43263;
  assign n43266 = ~n44468 | ~n43281;
  assign n43265 = ~n44469 | ~n43282;
  assign n43270 = ~n43266 | ~n43265;
  assign n43268 = ~n44472 | ~n43372;
  assign n43267 = ~n44473 | ~n43285;
  assign n43269 = ~n43268 | ~n43267;
  assign n43272 = ~n43270 & ~n43269;
  assign n43271 = ~P1_INSTQUEUE_REG_1__5__SCAN_IN | ~n43290;
  assign P1_U3046 = ~n43272 | ~n43271;
  assign n43274 = ~n22825 | ~n43281;
  assign n43273 = ~n44480 | ~n43282;
  assign n43278 = ~n43274 | ~n43273;
  assign n43276 = ~n44483 | ~n43372;
  assign n43275 = ~n44484 | ~n43285;
  assign n43277 = ~n43276 | ~n43275;
  assign n43280 = ~n43278 & ~n43277;
  assign n43279 = ~P1_INSTQUEUE_REG_1__6__SCAN_IN | ~n43290;
  assign P1_U3047 = ~n43280 | ~n43279;
  assign n43284 = ~n44492 | ~n43281;
  assign n43283 = ~n44494 | ~n43282;
  assign n43289 = ~n43284 | ~n43283;
  assign n43287 = ~n44498 | ~n43372;
  assign n43286 = ~n44500 | ~n43285;
  assign n43288 = ~n43287 | ~n43286;
  assign n43292 = ~n43289 & ~n43288;
  assign n43291 = ~P1_INSTQUEUE_REG_1__7__SCAN_IN | ~n43290;
  assign P1_U3048 = ~n43292 | ~n43291;
  assign n43293 = ~n44781 | ~n43066;
  assign n43296 = ~n44405 | ~n43450;
  assign n43375 = ~P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN | ~n43294;
  assign n43363 = ~P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN & ~n43375;
  assign n43295 = ~n44394 | ~n43363;
  assign n43305 = ~n43296 | ~n43295;
  assign n43308 = n44152 | P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN;
  assign n43635 = ~n43308;
  assign n43301 = ~n43470 | ~n43635;
  assign n43297 = n43372 | n43450;
  assign n43298 = ~n43297 | ~P1_STATEBS16_REG_SCAN_IN;
  assign n43307 = ~n43298 | ~n44800;
  assign n43299 = ~n43307;
  assign n43306 = ~n43380 & ~n44311;
  assign n43300 = ~n43299 | ~n43306;
  assign n43367 = ~n43301 | ~n43300;
  assign n43303 = ~n44402 | ~n43367;
  assign n43302 = ~n44406 | ~n43372;
  assign n43304 = ~n43303 | ~n43302;
  assign n43314 = ~n43305 & ~n43304;
  assign n43311 = ~n43307 & ~n43306;
  assign n43650 = ~n43308 | ~P1_STATE2_REG_2__SCAN_IN;
  assign n43309 = n44766 | n43363;
  assign n43310 = ~n43650 | ~n43309;
  assign n43313 = ~P1_INSTQUEUE_REG_2__0__SCAN_IN | ~n43366;
  assign P1_U3049 = ~n43314 | ~n43313;
  assign n43316 = ~n43102 | ~n43363;
  assign n43315 = ~n44427 | ~n43450;
  assign n43320 = ~n43316 | ~n43315;
  assign n43318 = ~P1_INSTQUEUE_REG_2__1__SCAN_IN | ~n43366;
  assign n43317 = ~n44424 | ~n43367;
  assign n43319 = ~n43318 | ~n43317;
  assign n43322 = ~n43320 & ~n43319;
  assign n43321 = ~n44428 | ~n43372;
  assign P1_U3050 = ~n43322 | ~n43321;
  assign n43324 = ~n43117 | ~n43363;
  assign n43323 = ~n44438 | ~n43450;
  assign n43328 = ~n43324 | ~n43323;
  assign n43326 = ~P1_INSTQUEUE_REG_2__2__SCAN_IN | ~n43366;
  assign n43325 = ~n44435 | ~n43367;
  assign n43327 = ~n43326 | ~n43325;
  assign n43330 = ~n43328 & ~n43327;
  assign n43329 = ~n44439 | ~n43372;
  assign P1_U3051 = ~n43330 | ~n43329;
  assign n43332 = ~n43132 | ~n43363;
  assign n43331 = ~n44449 | ~n43450;
  assign n43336 = ~n43332 | ~n43331;
  assign n43334 = ~P1_INSTQUEUE_REG_2__3__SCAN_IN | ~n43366;
  assign n43333 = ~n44446 | ~n43367;
  assign n43335 = ~n43334 | ~n43333;
  assign n43338 = ~n43336 & ~n43335;
  assign n43337 = ~n44450 | ~n43372;
  assign P1_U3052 = ~n43338 | ~n43337;
  assign n43340 = ~n43147 | ~n43363;
  assign n43339 = ~n44460 | ~n43450;
  assign n43344 = ~n43340 | ~n43339;
  assign n43342 = ~P1_INSTQUEUE_REG_2__4__SCAN_IN | ~n43366;
  assign n43341 = ~n44457 | ~n43367;
  assign n43343 = ~n43342 | ~n43341;
  assign n43346 = ~n43344 & ~n43343;
  assign n43345 = ~n44461 | ~n43372;
  assign P1_U3053 = ~n43346 | ~n43345;
  assign n43348 = ~n44468 | ~n43363;
  assign n43347 = ~n44472 | ~n43450;
  assign n43352 = ~n43348 | ~n43347;
  assign n43350 = ~P1_INSTQUEUE_REG_2__5__SCAN_IN | ~n43366;
  assign n43349 = ~n44469 | ~n43367;
  assign n43351 = ~n43350 | ~n43349;
  assign n43354 = ~n43352 & ~n43351;
  assign n43353 = ~n44473 | ~n43372;
  assign P1_U3054 = ~n43354 | ~n43353;
  assign n43356 = ~n22825 | ~n43363;
  assign n43355 = ~n44483 | ~n43450;
  assign n43360 = ~n43356 | ~n43355;
  assign n43358 = ~P1_INSTQUEUE_REG_2__6__SCAN_IN | ~n43366;
  assign n43357 = ~n44480 | ~n43367;
  assign n43359 = ~n43358 | ~n43357;
  assign n43362 = ~n43360 & ~n43359;
  assign n43361 = ~n44484 | ~n43372;
  assign P1_U3055 = ~n43362 | ~n43361;
  assign n43365 = ~n44492 | ~n43363;
  assign n43364 = ~n44498 | ~n43450;
  assign n43371 = ~n43365 | ~n43364;
  assign n43369 = ~P1_INSTQUEUE_REG_2__7__SCAN_IN | ~n43366;
  assign n43368 = ~n44494 | ~n43367;
  assign n43370 = ~n43369 | ~n43368;
  assign n43374 = ~n43371 & ~n43370;
  assign n43373 = ~n44500 | ~n43372;
  assign P1_U3056 = ~n43374 | ~n43373;
  assign n43387 = ~n43375;
  assign n43377 = ~n44394 | ~n43449;
  assign n43376 = ~n44406 | ~n43450;
  assign n43396 = ~n43377 | ~n43376;
  assign n43378 = ~n44399 & ~n43387;
  assign n43386 = ~n43378 & ~n44415;
  assign n43382 = n43380 | n43716;
  assign n43381 = ~n43449;
  assign n43383 = ~n44781 | ~n44775;
  assign n43384 = ~n43072 & ~n43383;
  assign n43390 = ~n43384 & ~n44418;
  assign n43385 = ~n43388 | ~n43390;
  assign n43394 = ~P1_INSTQUEUE_REG_3__0__SCAN_IN | ~n43458;
  assign n43392 = ~P1_STATE2_REG_2__SCAN_IN | ~n43387;
  assign n43389 = ~n43388;
  assign n43391 = ~n43390 | ~n43389;
  assign n43453 = ~n43392 | ~n43391;
  assign n43393 = ~n44402 | ~n43453;
  assign n43395 = ~n43394 | ~n43393;
  assign n43400 = ~n43396 & ~n43395;
  assign n43399 = ~n44405 | ~n43398;
  assign P1_U3057 = ~n43400 | ~n43399;
  assign n43402 = ~n43102 | ~n43449;
  assign n43401 = ~n44428 | ~n43450;
  assign n43406 = ~n43402 | ~n43401;
  assign n43404 = ~n44424 | ~n43453;
  assign n43403 = ~n44427 | ~n43398;
  assign n43405 = ~n43404 | ~n43403;
  assign n43408 = ~n43406 & ~n43405;
  assign n43407 = ~P1_INSTQUEUE_REG_3__1__SCAN_IN | ~n43458;
  assign P1_U3058 = ~n43408 | ~n43407;
  assign n43410 = ~n43117 | ~n43449;
  assign n43409 = ~n44439 | ~n43450;
  assign n43414 = ~n43410 | ~n43409;
  assign n43412 = ~n44435 | ~n43453;
  assign n43411 = ~n44438 | ~n43398;
  assign n43413 = ~n43412 | ~n43411;
  assign n43416 = ~n43414 & ~n43413;
  assign n43415 = ~P1_INSTQUEUE_REG_3__2__SCAN_IN | ~n43458;
  assign P1_U3059 = ~n43416 | ~n43415;
  assign n43418 = ~n43132 | ~n43449;
  assign n43417 = ~n44450 | ~n43450;
  assign n43422 = ~n43418 | ~n43417;
  assign n43420 = ~n44446 | ~n43453;
  assign n43419 = ~n44449 | ~n43398;
  assign n43421 = ~n43420 | ~n43419;
  assign n43424 = ~n43422 & ~n43421;
  assign n43423 = ~P1_INSTQUEUE_REG_3__3__SCAN_IN | ~n43458;
  assign P1_U3060 = ~n43424 | ~n43423;
  assign n43426 = ~n43147 | ~n43449;
  assign n43425 = ~n44461 | ~n43450;
  assign n43430 = ~n43426 | ~n43425;
  assign n43428 = ~P1_INSTQUEUE_REG_3__4__SCAN_IN | ~n43458;
  assign n43427 = ~n44460 | ~n43398;
  assign n43429 = ~n43428 | ~n43427;
  assign n43432 = ~n43430 & ~n43429;
  assign n43431 = ~n44457 | ~n43453;
  assign P1_U3061 = ~n43432 | ~n43431;
  assign n43434 = ~n44468 | ~n43449;
  assign n43433 = ~n44473 | ~n43450;
  assign n43438 = ~n43434 | ~n43433;
  assign n43436 = ~n44469 | ~n43453;
  assign n43435 = ~n44472 | ~n43398;
  assign n43437 = ~n43436 | ~n43435;
  assign n43440 = ~n43438 & ~n43437;
  assign n43439 = ~P1_INSTQUEUE_REG_3__5__SCAN_IN | ~n43458;
  assign P1_U3062 = ~n43440 | ~n43439;
  assign n43442 = ~n22825 | ~n43449;
  assign n43441 = ~n44483 | ~n43398;
  assign n43446 = ~n43442 | ~n43441;
  assign n43444 = ~P1_INSTQUEUE_REG_3__6__SCAN_IN | ~n43458;
  assign n43443 = ~n44484 | ~n43450;
  assign n43445 = ~n43444 | ~n43443;
  assign n43448 = ~n43446 & ~n43445;
  assign n43447 = ~n44480 | ~n43453;
  assign P1_U3063 = ~n43448 | ~n43447;
  assign n43452 = ~n44492 | ~n43449;
  assign n43451 = ~n44500 | ~n43450;
  assign n43457 = ~n43452 | ~n43451;
  assign n43455 = ~n44494 | ~n43453;
  assign n43454 = ~n44498 | ~n43398;
  assign n43456 = ~n43455 | ~n43454;
  assign n43460 = ~n43457 & ~n43456;
  assign n43459 = ~P1_INSTQUEUE_REG_3__7__SCAN_IN | ~n43458;
  assign P1_U3064 = ~n43460 | ~n43459;
  assign n43461 = ~P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN & ~P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN;
  assign n43547 = ~n43461 | ~P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign n43478 = n43547 | P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign n43535 = ~n43478;
  assign n43467 = ~n44394 | ~n43535;
  assign n44137 = ~n43636;
  assign n43462 = ~n44137 & ~n44153;
  assign n43465 = ~n43462 | ~n44152;
  assign n43475 = ~n43717 | ~n44311;
  assign n43463 = ~n43475;
  assign n43464 = ~n43463 | ~n44800;
  assign n43536 = ~n43465 | ~n43464;
  assign n43466 = ~n44402 | ~n43536;
  assign n43484 = ~n43467 | ~n43466;
  assign n43468 = ~n43065;
  assign n43469 = ~n43468 & ~n43066;
  assign n44778 = ~n44781;
  assign n43568 = ~n43469 | ~n44778;
  assign n43624 = ~n43568 & ~n44801;
  assign n43482 = ~n44405 | ~n43624;
  assign n43473 = ~n43624;
  assign n43472 = ~n43398;
  assign n43474 = ~n43473 | ~n43472;
  assign n43476 = ~n43474 | ~P1_STATEBS16_REG_SCAN_IN;
  assign n43477 = ~n43476 | ~n43475;
  assign n43479 = ~n43477 | ~n44766;
  assign n43480 = ~n43479 | ~n43478;
  assign n43481 = ~P1_INSTQUEUE_REG_4__0__SCAN_IN | ~n43544;
  assign n43483 = ~n43482 | ~n43481;
  assign n43486 = ~n43484 & ~n43483;
  assign n43485 = ~n44406 | ~n43398;
  assign P1_U3065 = ~n43486 | ~n43485;
  assign n43488 = ~n43102 | ~n43535;
  assign n43487 = ~n44424 | ~n43536;
  assign n43492 = ~n43488 | ~n43487;
  assign n43490 = ~n44427 | ~n43624;
  assign n43489 = ~n44428 | ~n43398;
  assign n43491 = ~n43490 | ~n43489;
  assign n43494 = ~n43492 & ~n43491;
  assign n43493 = ~P1_INSTQUEUE_REG_4__1__SCAN_IN | ~n43544;
  assign P1_U3066 = ~n43494 | ~n43493;
  assign n43496 = ~n43117 | ~n43535;
  assign n43495 = ~n44435 | ~n43536;
  assign n43500 = ~n43496 | ~n43495;
  assign n43498 = ~n44438 | ~n43624;
  assign n43497 = ~n44439 | ~n43398;
  assign n43499 = ~n43498 | ~n43497;
  assign n43502 = ~n43500 & ~n43499;
  assign n43501 = ~P1_INSTQUEUE_REG_4__2__SCAN_IN | ~n43544;
  assign P1_U3067 = ~n43502 | ~n43501;
  assign n43504 = ~n43132 | ~n43535;
  assign n43503 = ~n44446 | ~n43536;
  assign n43508 = ~n43504 | ~n43503;
  assign n43506 = ~n44449 | ~n43624;
  assign n43505 = ~n44450 | ~n43398;
  assign n43507 = ~n43506 | ~n43505;
  assign n43510 = ~n43508 & ~n43507;
  assign n43509 = ~P1_INSTQUEUE_REG_4__3__SCAN_IN | ~n43544;
  assign P1_U3068 = ~n43510 | ~n43509;
  assign n43512 = ~n43147 | ~n43535;
  assign n43511 = ~n44457 | ~n43536;
  assign n43516 = ~n43512 | ~n43511;
  assign n43514 = ~n44460 | ~n43624;
  assign n43513 = ~n44461 | ~n43398;
  assign n43515 = ~n43514 | ~n43513;
  assign n43518 = ~n43516 & ~n43515;
  assign n43517 = ~P1_INSTQUEUE_REG_4__4__SCAN_IN | ~n43544;
  assign P1_U3069 = ~n43518 | ~n43517;
  assign n43520 = ~n44468 | ~n43535;
  assign n43519 = ~n44469 | ~n43536;
  assign n43524 = ~n43520 | ~n43519;
  assign n43522 = ~n44472 | ~n43624;
  assign n43521 = ~n44473 | ~n43398;
  assign n43523 = ~n43522 | ~n43521;
  assign n43526 = ~n43524 & ~n43523;
  assign n43525 = ~P1_INSTQUEUE_REG_4__5__SCAN_IN | ~n43544;
  assign P1_U3070 = ~n43526 | ~n43525;
  assign n43528 = ~n22825 | ~n43535;
  assign n43527 = ~n44480 | ~n43536;
  assign n43532 = ~n43528 | ~n43527;
  assign n43530 = ~n44483 | ~n43624;
  assign n43529 = ~n44484 | ~n43398;
  assign n43531 = ~n43530 | ~n43529;
  assign n43534 = ~n43532 & ~n43531;
  assign n43533 = ~P1_INSTQUEUE_REG_4__6__SCAN_IN | ~n43544;
  assign P1_U3071 = ~n43534 | ~n43533;
  assign n43538 = ~n44492 | ~n43535;
  assign n43537 = ~n44494 | ~n43536;
  assign n43543 = ~n43538 | ~n43537;
  assign n43541 = ~n44498 | ~n43624;
  assign n43540 = ~n44500 | ~n43398;
  assign n43542 = ~n43541 | ~n43540;
  assign n43546 = ~n43543 & ~n43542;
  assign n43545 = ~P1_INSTQUEUE_REG_4__7__SCAN_IN | ~n43544;
  assign P1_U3072 = ~n43546 | ~n43545;
  assign n43620 = ~n43547 & ~n44308;
  assign n43553 = ~n44394 | ~n43620;
  assign n43554 = ~n43547;
  assign n43551 = ~n43554 | ~P1_STATE2_REG_2__SCAN_IN;
  assign n43559 = ~n43548 & ~n43880;
  assign n43549 = n43559 | n43620;
  assign n43550 = ~n43549 | ~n44800;
  assign n43621 = ~n43551 | ~n43550;
  assign n43552 = ~n44402 | ~n43621;
  assign n43567 = ~n43553 | ~n43552;
  assign n43555 = ~n43554 & ~n44399;
  assign n43563 = ~n43555 & ~n44415;
  assign n43556 = ~n43568;
  assign n43561 = ~n43556 | ~P1_STATEBS16_REG_SCAN_IN;
  assign n43557 = ~n43620;
  assign n43558 = ~n43557 | ~n44800;
  assign n43560 = ~n43559 & ~n43558;
  assign n43562 = ~n43561 | ~n43560;
  assign n43565 = ~P1_INSTQUEUE_REG_5__0__SCAN_IN | ~n43629;
  assign n43564 = ~n44406 | ~n43624;
  assign n43566 = ~n43565 | ~n43564;
  assign n43571 = ~n43567 & ~n43566;
  assign n43570 = ~n44405 | ~n43569;
  assign P1_U3073 = ~n43571 | ~n43570;
  assign n43573 = ~n43102 | ~n43620;
  assign n43572 = ~n44424 | ~n43621;
  assign n43577 = ~n43573 | ~n43572;
  assign n43575 = ~n44427 | ~n43569;
  assign n43574 = ~n44428 | ~n43624;
  assign n43576 = ~n43575 | ~n43574;
  assign n43579 = ~n43577 & ~n43576;
  assign n43578 = ~P1_INSTQUEUE_REG_5__1__SCAN_IN | ~n43629;
  assign P1_U3074 = ~n43579 | ~n43578;
  assign n43581 = ~n43117 | ~n43620;
  assign n43580 = ~n44435 | ~n43621;
  assign n43585 = ~n43581 | ~n43580;
  assign n43583 = ~n44438 | ~n43569;
  assign n43582 = ~n44439 | ~n43624;
  assign n43584 = ~n43583 | ~n43582;
  assign n43587 = ~n43585 & ~n43584;
  assign n43586 = ~P1_INSTQUEUE_REG_5__2__SCAN_IN | ~n43629;
  assign P1_U3075 = ~n43587 | ~n43586;
  assign n43589 = ~n43132 | ~n43620;
  assign n43588 = ~n44446 | ~n43621;
  assign n43593 = ~n43589 | ~n43588;
  assign n43591 = ~n44449 | ~n43569;
  assign n43590 = ~n44450 | ~n43624;
  assign n43592 = ~n43591 | ~n43590;
  assign n43595 = ~n43593 & ~n43592;
  assign n43594 = ~P1_INSTQUEUE_REG_5__3__SCAN_IN | ~n43629;
  assign P1_U3076 = ~n43595 | ~n43594;
  assign n43597 = ~n43147 | ~n43620;
  assign n43596 = ~n44457 | ~n43621;
  assign n43601 = ~n43597 | ~n43596;
  assign n43599 = ~n44460 | ~n43569;
  assign n43598 = ~n44461 | ~n43624;
  assign n43600 = ~n43599 | ~n43598;
  assign n43603 = ~n43601 & ~n43600;
  assign n43602 = ~P1_INSTQUEUE_REG_5__4__SCAN_IN | ~n43629;
  assign P1_U3077 = ~n43603 | ~n43602;
  assign n43605 = ~n44468 | ~n43620;
  assign n43604 = ~n44469 | ~n43621;
  assign n43609 = ~n43605 | ~n43604;
  assign n43607 = ~n44472 | ~n43569;
  assign n43606 = ~n44473 | ~n43624;
  assign n43608 = ~n43607 | ~n43606;
  assign n43611 = ~n43609 & ~n43608;
  assign n43610 = ~P1_INSTQUEUE_REG_5__5__SCAN_IN | ~n43629;
  assign P1_U3078 = ~n43611 | ~n43610;
  assign n43613 = ~n22825 | ~n43620;
  assign n43612 = ~n44480 | ~n43621;
  assign n43617 = ~n43613 | ~n43612;
  assign n43615 = ~n44483 | ~n43569;
  assign n43614 = ~n44484 | ~n43624;
  assign n43616 = ~n43615 | ~n43614;
  assign n43619 = ~n43617 & ~n43616;
  assign n43618 = ~P1_INSTQUEUE_REG_5__6__SCAN_IN | ~n43629;
  assign P1_U3079 = ~n43619 | ~n43618;
  assign n43623 = ~n44492 | ~n43620;
  assign n43622 = ~n44494 | ~n43621;
  assign n43628 = ~n43623 | ~n43622;
  assign n43626 = ~n44498 | ~n43569;
  assign n43625 = ~n44500 | ~n43624;
  assign n43627 = ~n43626 | ~n43625;
  assign n43631 = ~n43628 & ~n43627;
  assign n43630 = ~P1_INSTQUEUE_REG_5__7__SCAN_IN | ~n43629;
  assign P1_U3080 = ~n43631 | ~n43630;
  assign n43648 = ~n43729 | ~n44308;
  assign n43705 = ~n43648;
  assign n43634 = ~n44394 | ~n43705;
  assign n43632 = ~n43065 | ~n43066;
  assign n43791 = ~n44760 & ~n44801;
  assign n43633 = ~n44405 | ~n43791;
  assign n43645 = ~n43634 | ~n43633;
  assign n43641 = ~n43636 | ~n43635;
  assign n43637 = ~n43569 & ~n43791;
  assign n43638 = ~n43637 & ~n44765;
  assign n43647 = ~n43638 & ~n44418;
  assign n43646 = ~n43717 | ~n31534;
  assign n43639 = ~n43646;
  assign n43640 = ~n43647 | ~n43639;
  assign n43643 = ~n44402 | ~n43713;
  assign n43642 = ~n44406 | ~n43569;
  assign n43644 = ~n43643 | ~n43642;
  assign n43656 = ~n43645 & ~n43644;
  assign n43654 = ~n43647 | ~n43646;
  assign n43652 = ~n44327;
  assign n43649 = ~n43648 | ~P1_STATE2_REG_3__SCAN_IN;
  assign n43651 = ~n43650 | ~n43649;
  assign n43653 = ~n43652 & ~n43651;
  assign n43655 = ~P1_INSTQUEUE_REG_6__0__SCAN_IN | ~n43708;
  assign P1_U3081 = ~n43656 | ~n43655;
  assign n43658 = ~n43102 | ~n43705;
  assign n43657 = ~n44427 | ~n43791;
  assign n43662 = ~n43658 | ~n43657;
  assign n43660 = ~P1_INSTQUEUE_REG_6__1__SCAN_IN | ~n43708;
  assign n43659 = ~n44428 | ~n43569;
  assign n43661 = ~n43660 | ~n43659;
  assign n43664 = ~n43662 & ~n43661;
  assign n43663 = ~n44424 | ~n43713;
  assign P1_U3082 = ~n43664 | ~n43663;
  assign n43666 = ~n43117 | ~n43705;
  assign n43665 = ~n44438 | ~n43791;
  assign n43670 = ~n43666 | ~n43665;
  assign n43668 = ~n44435 | ~n43713;
  assign n43667 = ~n44439 | ~n43569;
  assign n43669 = ~n43668 | ~n43667;
  assign n43672 = ~n43670 & ~n43669;
  assign n43671 = ~P1_INSTQUEUE_REG_6__2__SCAN_IN | ~n43708;
  assign P1_U3083 = ~n43672 | ~n43671;
  assign n43674 = ~n43132 | ~n43705;
  assign n43673 = ~n44449 | ~n43791;
  assign n43678 = ~n43674 | ~n43673;
  assign n43676 = ~n44446 | ~n43713;
  assign n43675 = ~n44450 | ~n43569;
  assign n43677 = ~n43676 | ~n43675;
  assign n43680 = ~n43678 & ~n43677;
  assign n43679 = ~P1_INSTQUEUE_REG_6__3__SCAN_IN | ~n43708;
  assign P1_U3084 = ~n43680 | ~n43679;
  assign n43682 = ~n43147 | ~n43705;
  assign n43681 = ~n44460 | ~n43791;
  assign n43686 = ~n43682 | ~n43681;
  assign n43684 = ~n44457 | ~n43713;
  assign n43683 = ~n44461 | ~n43569;
  assign n43685 = ~n43684 | ~n43683;
  assign n43688 = ~n43686 & ~n43685;
  assign n43687 = ~P1_INSTQUEUE_REG_6__4__SCAN_IN | ~n43708;
  assign P1_U3085 = ~n43688 | ~n43687;
  assign n43690 = ~n44468 | ~n43705;
  assign n43689 = ~n44472 | ~n43791;
  assign n43694 = ~n43690 | ~n43689;
  assign n43692 = ~P1_INSTQUEUE_REG_6__5__SCAN_IN | ~n43708;
  assign n43691 = ~n44473 | ~n43569;
  assign n43693 = ~n43692 | ~n43691;
  assign n43696 = ~n43694 & ~n43693;
  assign n43695 = ~n44469 | ~n43713;
  assign P1_U3086 = ~n43696 | ~n43695;
  assign n43698 = ~n22825 | ~n43705;
  assign n43697 = ~n44483 | ~n43791;
  assign n43702 = ~n43698 | ~n43697;
  assign n43700 = ~P1_INSTQUEUE_REG_6__6__SCAN_IN | ~n43708;
  assign n43699 = ~n44484 | ~n43569;
  assign n43701 = ~n43700 | ~n43699;
  assign n43704 = ~n43702 & ~n43701;
  assign n43703 = ~n44480 | ~n43713;
  assign P1_U3087 = ~n43704 | ~n43703;
  assign n43707 = ~n44492 | ~n43705;
  assign n43706 = ~n44498 | ~n43791;
  assign n43712 = ~n43707 | ~n43706;
  assign n43710 = ~P1_INSTQUEUE_REG_6__7__SCAN_IN | ~n43708;
  assign n43709 = ~n44500 | ~n43569;
  assign n43711 = ~n43710 | ~n43709;
  assign n43715 = ~n43712 & ~n43711;
  assign n43714 = ~n44494 | ~n43713;
  assign P1_U3088 = ~n43715 | ~n43714;
  assign n43787 = ~n43718;
  assign n43723 = ~n44394 | ~n43787;
  assign n44395 = ~n43716;
  assign n43719 = ~n43717 | ~n44395;
  assign n43730 = ~n43719 | ~n43718;
  assign n43721 = ~n43730 | ~n44800;
  assign n43720 = ~n43729 | ~P1_STATE2_REG_2__SCAN_IN;
  assign n43788 = ~n43721 | ~n43720;
  assign n43722 = ~n44402 | ~n43788;
  assign n43728 = ~n43723 | ~n43722;
  assign n43724 = ~n44760 & ~n44230;
  assign n43726 = ~n44405 | ~n43871;
  assign n43725 = ~n44406 | ~n43791;
  assign n43727 = ~n43726 | ~n43725;
  assign n43738 = ~n43728 & ~n43727;
  assign n43736 = ~n44415;
  assign n43734 = ~n43729 & ~n44399;
  assign n43732 = ~n44765 & ~n44760;
  assign n43731 = n44418 | n43730;
  assign n43733 = ~n43732 & ~n43731;
  assign n43735 = ~n43734 & ~n43733;
  assign n43737 = ~P1_INSTQUEUE_REG_7__0__SCAN_IN | ~n43796;
  assign P1_U3089 = ~n43738 | ~n43737;
  assign n43740 = ~n43102 | ~n43787;
  assign n43739 = ~n44424 | ~n43788;
  assign n43744 = ~n43740 | ~n43739;
  assign n43742 = ~n44427 | ~n43871;
  assign n43741 = ~n44428 | ~n43791;
  assign n43743 = ~n43742 | ~n43741;
  assign n43746 = ~n43744 & ~n43743;
  assign n43745 = ~P1_INSTQUEUE_REG_7__1__SCAN_IN | ~n43796;
  assign P1_U3090 = ~n43746 | ~n43745;
  assign n43748 = ~n43117 | ~n43787;
  assign n43747 = ~n44435 | ~n43788;
  assign n43752 = ~n43748 | ~n43747;
  assign n43750 = ~n44438 | ~n43871;
  assign n43749 = ~n44439 | ~n43791;
  assign n43751 = ~n43750 | ~n43749;
  assign n43754 = ~n43752 & ~n43751;
  assign n43753 = ~P1_INSTQUEUE_REG_7__2__SCAN_IN | ~n43796;
  assign P1_U3091 = ~n43754 | ~n43753;
  assign n43756 = ~n43132 | ~n43787;
  assign n43755 = ~n44446 | ~n43788;
  assign n43760 = ~n43756 | ~n43755;
  assign n43758 = ~n44449 | ~n43871;
  assign n43757 = ~n44450 | ~n43791;
  assign n43759 = ~n43758 | ~n43757;
  assign n43762 = ~n43760 & ~n43759;
  assign n43761 = ~P1_INSTQUEUE_REG_7__3__SCAN_IN | ~n43796;
  assign P1_U3092 = ~n43762 | ~n43761;
  assign n43764 = ~n43147 | ~n43787;
  assign n43763 = ~n44457 | ~n43788;
  assign n43768 = ~n43764 | ~n43763;
  assign n43766 = ~n44460 | ~n43871;
  assign n43765 = ~n44461 | ~n43791;
  assign n43767 = ~n43766 | ~n43765;
  assign n43770 = ~n43768 & ~n43767;
  assign n43769 = ~P1_INSTQUEUE_REG_7__4__SCAN_IN | ~n43796;
  assign P1_U3093 = ~n43770 | ~n43769;
  assign n43772 = ~n44468 | ~n43787;
  assign n43771 = ~n44469 | ~n43788;
  assign n43776 = ~n43772 | ~n43771;
  assign n43774 = ~n44472 | ~n43871;
  assign n43773 = ~n44473 | ~n43791;
  assign n43775 = ~n43774 | ~n43773;
  assign n43778 = ~n43776 & ~n43775;
  assign n43777 = ~P1_INSTQUEUE_REG_7__5__SCAN_IN | ~n43796;
  assign P1_U3094 = ~n43778 | ~n43777;
  assign n43780 = ~n22825 | ~n43787;
  assign n43779 = ~n44480 | ~n43788;
  assign n43784 = ~n43780 | ~n43779;
  assign n43782 = ~n44483 | ~n43871;
  assign n43781 = ~n44484 | ~n43791;
  assign n43783 = ~n43782 | ~n43781;
  assign n43786 = ~n43784 & ~n43783;
  assign n43785 = ~P1_INSTQUEUE_REG_7__6__SCAN_IN | ~n43796;
  assign P1_U3095 = ~n43786 | ~n43785;
  assign n43790 = ~n44492 | ~n43787;
  assign n43789 = ~n44494 | ~n43788;
  assign n43795 = ~n43790 | ~n43789;
  assign n43793 = ~n44498 | ~n43871;
  assign n43792 = ~n44500 | ~n43791;
  assign n43794 = ~n43793 | ~n43792;
  assign n43798 = ~n43795 & ~n43794;
  assign n43797 = ~P1_INSTQUEUE_REG_7__7__SCAN_IN | ~n43796;
  assign P1_U3096 = ~n43798 | ~n43797;
  assign n44133 = ~n43799 | ~P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN;
  assign n43879 = ~n44133 & ~P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign n43898 = ~n43879;
  assign n43806 = ~n44394 | ~n43867;
  assign n43800 = ~n43977 & ~n44136;
  assign n43804 = ~n43800 | ~n44152;
  assign n43802 = ~n44051 | ~n44311;
  assign n43801 = ~n43867;
  assign n43809 = ~n43802 | ~n43801;
  assign n43803 = ~n43809 | ~n44800;
  assign n43868 = ~n43804 | ~n43803;
  assign n43805 = ~n44402 | ~n43868;
  assign n43816 = ~n43806 | ~n43805;
  assign n44070 = ~n43072 | ~n44781;
  assign n43955 = ~n43892 & ~n44801;
  assign n43807 = ~n43955 & ~n43871;
  assign n43808 = ~n44765 & ~n43807;
  assign n43811 = ~n43809 & ~n43808;
  assign n43810 = ~n43867 & ~n44766;
  assign n43812 = ~n43811 & ~n43810;
  assign n43814 = ~P1_INSTQUEUE_REG_8__0__SCAN_IN | ~n43876;
  assign n43813 = ~n44406 | ~n43871;
  assign n43815 = ~n43814 | ~n43813;
  assign n43818 = ~n43816 & ~n43815;
  assign n43817 = ~n44405 | ~n43955;
  assign P1_U3097 = ~n43818 | ~n43817;
  assign n43820 = ~n43102 | ~n43867;
  assign n43819 = ~n44424 | ~n43868;
  assign n43824 = ~n43820 | ~n43819;
  assign n43822 = ~n44427 | ~n43955;
  assign n43821 = ~n44428 | ~n43871;
  assign n43823 = ~n43822 | ~n43821;
  assign n43826 = ~n43824 & ~n43823;
  assign n43825 = ~P1_INSTQUEUE_REG_8__1__SCAN_IN | ~n43876;
  assign P1_U3098 = ~n43826 | ~n43825;
  assign n43828 = ~n43117 | ~n43867;
  assign n43827 = ~n44435 | ~n43868;
  assign n43832 = ~n43828 | ~n43827;
  assign n43830 = ~n44438 | ~n43955;
  assign n43829 = ~n44439 | ~n43871;
  assign n43831 = ~n43830 | ~n43829;
  assign n43834 = ~n43832 & ~n43831;
  assign n43833 = ~P1_INSTQUEUE_REG_8__2__SCAN_IN | ~n43876;
  assign P1_U3099 = ~n43834 | ~n43833;
  assign n43836 = ~n43132 | ~n43867;
  assign n43835 = ~n44446 | ~n43868;
  assign n43840 = ~n43836 | ~n43835;
  assign n43838 = ~n44449 | ~n43955;
  assign n43837 = ~n44450 | ~n43871;
  assign n43839 = ~n43838 | ~n43837;
  assign n43842 = ~n43840 & ~n43839;
  assign n43841 = ~P1_INSTQUEUE_REG_8__3__SCAN_IN | ~n43876;
  assign P1_U3100 = ~n43842 | ~n43841;
  assign n43844 = ~n43147 | ~n43867;
  assign n43843 = ~n44457 | ~n43868;
  assign n43848 = ~n43844 | ~n43843;
  assign n43846 = ~n44460 | ~n43955;
  assign n43845 = ~n44461 | ~n43871;
  assign n43847 = ~n43846 | ~n43845;
  assign n43850 = ~n43848 & ~n43847;
  assign n43849 = ~P1_INSTQUEUE_REG_8__4__SCAN_IN | ~n43876;
  assign P1_U3101 = ~n43850 | ~n43849;
  assign n43852 = ~n44468 | ~n43867;
  assign n43851 = ~n44469 | ~n43868;
  assign n43856 = ~n43852 | ~n43851;
  assign n43854 = ~n44472 | ~n43955;
  assign n43853 = ~n44473 | ~n43871;
  assign n43855 = ~n43854 | ~n43853;
  assign n43858 = ~n43856 & ~n43855;
  assign n43857 = ~P1_INSTQUEUE_REG_8__5__SCAN_IN | ~n43876;
  assign P1_U3102 = ~n43858 | ~n43857;
  assign n43860 = ~n22825 | ~n43867;
  assign n43859 = ~n44480 | ~n43868;
  assign n43864 = ~n43860 | ~n43859;
  assign n43862 = ~n44483 | ~n43955;
  assign n43861 = ~n44484 | ~n43871;
  assign n43863 = ~n43862 | ~n43861;
  assign n43866 = ~n43864 & ~n43863;
  assign n43865 = ~P1_INSTQUEUE_REG_8__6__SCAN_IN | ~n43876;
  assign P1_U3103 = ~n43866 | ~n43865;
  assign n43870 = ~n44492 | ~n43867;
  assign n43869 = ~n44494 | ~n43868;
  assign n43875 = ~n43870 | ~n43869;
  assign n43873 = ~n44498 | ~n43955;
  assign n43872 = ~n44500 | ~n43871;
  assign n43874 = ~n43873 | ~n43872;
  assign n43878 = ~n43875 & ~n43874;
  assign n43877 = ~P1_INSTQUEUE_REG_8__7__SCAN_IN | ~n43876;
  assign P1_U3104 = ~n43878 | ~n43877;
  assign n43886 = ~n44394 | ~n43951;
  assign n43884 = ~P1_STATE2_REG_2__SCAN_IN | ~n43879;
  assign n44223 = ~n43880;
  assign n43894 = ~n44051 | ~n44223;
  assign n43881 = ~n43951;
  assign n43882 = ~n43894 | ~n43881;
  assign n43883 = ~n43882 | ~n44399;
  assign n43952 = ~n43884 | ~n43883;
  assign n43885 = ~n44402 | ~n43952;
  assign n43891 = ~n43886 | ~n43885;
  assign n43887 = ~n43892 & ~n44230;
  assign n44039 = n43887;
  assign n43889 = ~n44405 | ~n44039;
  assign n43888 = ~n44406 | ~n43955;
  assign n43890 = ~n43889 | ~n43888;
  assign n43902 = ~n43891 & ~n43890;
  assign n43896 = ~n43892 & ~n44765;
  assign n43893 = ~n43951 & ~n44418;
  assign n43895 = ~n43894 | ~n43893;
  assign n43897 = ~n43896 & ~n43895;
  assign n43900 = ~n43897 & ~n44415;
  assign n43899 = ~n43898 | ~n44418;
  assign n43901 = ~P1_INSTQUEUE_REG_9__0__SCAN_IN | ~n43960;
  assign P1_U3105 = ~n43902 | ~n43901;
  assign n43904 = ~n43102 | ~n43951;
  assign n43903 = ~n44424 | ~n43952;
  assign n43908 = ~n43904 | ~n43903;
  assign n43906 = ~n44427 | ~n44039;
  assign n43905 = ~n44428 | ~n43955;
  assign n43907 = ~n43906 | ~n43905;
  assign n43910 = ~n43908 & ~n43907;
  assign n43909 = ~P1_INSTQUEUE_REG_9__1__SCAN_IN | ~n43960;
  assign P1_U3106 = ~n43910 | ~n43909;
  assign n43912 = ~n43117 | ~n43951;
  assign n43911 = ~n44435 | ~n43952;
  assign n43916 = ~n43912 | ~n43911;
  assign n43914 = ~n44438 | ~n44039;
  assign n43913 = ~n44439 | ~n43955;
  assign n43915 = ~n43914 | ~n43913;
  assign n43918 = ~n43916 & ~n43915;
  assign n43917 = ~P1_INSTQUEUE_REG_9__2__SCAN_IN | ~n43960;
  assign P1_U3107 = ~n43918 | ~n43917;
  assign n43920 = ~n43132 | ~n43951;
  assign n43919 = ~n44446 | ~n43952;
  assign n43924 = ~n43920 | ~n43919;
  assign n43922 = ~n44449 | ~n44039;
  assign n43921 = ~n44450 | ~n43955;
  assign n43923 = ~n43922 | ~n43921;
  assign n43926 = ~n43924 & ~n43923;
  assign n43925 = ~P1_INSTQUEUE_REG_9__3__SCAN_IN | ~n43960;
  assign P1_U3108 = ~n43926 | ~n43925;
  assign n43928 = ~n43147 | ~n43951;
  assign n43927 = ~n44457 | ~n43952;
  assign n43932 = ~n43928 | ~n43927;
  assign n43930 = ~n44460 | ~n44039;
  assign n43929 = ~n44461 | ~n43955;
  assign n43931 = ~n43930 | ~n43929;
  assign n43934 = ~n43932 & ~n43931;
  assign n43933 = ~P1_INSTQUEUE_REG_9__4__SCAN_IN | ~n43960;
  assign P1_U3109 = ~n43934 | ~n43933;
  assign n43936 = ~n44468 | ~n43951;
  assign n43935 = ~n44469 | ~n43952;
  assign n43940 = ~n43936 | ~n43935;
  assign n43938 = ~n44472 | ~n44039;
  assign n43937 = ~n44473 | ~n43955;
  assign n43939 = ~n43938 | ~n43937;
  assign n43942 = ~n43940 & ~n43939;
  assign n43941 = ~P1_INSTQUEUE_REG_9__5__SCAN_IN | ~n43960;
  assign P1_U3110 = ~n43942 | ~n43941;
  assign n43944 = ~n22825 | ~n43951;
  assign n43943 = ~n44480 | ~n43952;
  assign n43948 = ~n43944 | ~n43943;
  assign n43946 = ~n44483 | ~n44039;
  assign n43945 = ~n44484 | ~n43955;
  assign n43947 = ~n43946 | ~n43945;
  assign n43950 = ~n43948 & ~n43947;
  assign n43949 = ~P1_INSTQUEUE_REG_9__6__SCAN_IN | ~n43960;
  assign P1_U3111 = ~n43950 | ~n43949;
  assign n43954 = ~n44492 | ~n43951;
  assign n43953 = ~n44494 | ~n43952;
  assign n43959 = ~n43954 | ~n43953;
  assign n43957 = ~n44498 | ~n44039;
  assign n43956 = ~n44500 | ~n43955;
  assign n43958 = ~n43957 | ~n43956;
  assign n43962 = ~n43959 & ~n43958;
  assign n43961 = ~P1_INSTQUEUE_REG_9__7__SCAN_IN | ~n43960;
  assign P1_U3112 = ~n43962 | ~n43961;
  assign n43965 = ~n44406 | ~n44039;
  assign n43963 = ~P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | ~P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN;
  assign n44058 = ~n43963 & ~P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN;
  assign n43971 = ~n44058 | ~n44308;
  assign n44038 = ~n43971;
  assign n43964 = ~n44394 | ~n44038;
  assign n43987 = ~n43965 | ~n43964;
  assign n43966 = ~n43066 | ~n44230;
  assign n43968 = ~n43967 | ~P1_STATEBS16_REG_SCAN_IN;
  assign n43979 = ~n43968 | ~n44800;
  assign n43980 = ~n43969 & ~n44311;
  assign n43974 = ~n43979 & ~n43980;
  assign n43970 = n44152 | n44306;
  assign n44323 = ~n43970 | ~P1_STATE2_REG_2__SCAN_IN;
  assign n43972 = ~n43971 | ~P1_STATE2_REG_3__SCAN_IN;
  assign n43973 = ~n44323 | ~n43972;
  assign n43975 = ~n43974 & ~n43973;
  assign n43985 = ~P1_INSTQUEUE_REG_10__0__SCAN_IN | ~n44047;
  assign n43978 = ~n43977 & ~n44306;
  assign n44309 = ~n44152;
  assign n43983 = ~n43978 | ~n44309;
  assign n43981 = ~n43979;
  assign n43982 = ~n43981 | ~n43980;
  assign n43984 = ~n44402 | ~n44042;
  assign n43986 = ~n43985 | ~n43984;
  assign n43989 = ~n43987 & ~n43986;
  assign n43988 = ~n44405 | ~n22905;
  assign P1_U3113 = ~n43989 | ~n43988;
  assign n43991 = ~n43102 | ~n44038;
  assign n43990 = ~n44427 | ~n22905;
  assign n43995 = ~n43991 | ~n43990;
  assign n43993 = ~P1_INSTQUEUE_REG_10__1__SCAN_IN | ~n44047;
  assign n43992 = ~n44428 | ~n44039;
  assign n43994 = ~n43993 | ~n43992;
  assign n43997 = ~n43995 & ~n43994;
  assign n43996 = ~n44424 | ~n44042;
  assign P1_U3114 = ~n43997 | ~n43996;
  assign n43999 = ~n43117 | ~n44038;
  assign n43998 = ~n44439 | ~n44039;
  assign n44003 = ~n43999 | ~n43998;
  assign n44001 = ~P1_INSTQUEUE_REG_10__2__SCAN_IN | ~n44047;
  assign n44000 = ~n44438 | ~n22905;
  assign n44002 = ~n44001 | ~n44000;
  assign n44005 = ~n44003 & ~n44002;
  assign n44004 = ~n44435 | ~n44042;
  assign P1_U3115 = ~n44005 | ~n44004;
  assign n44007 = ~n43132 | ~n44038;
  assign n44006 = ~n44449 | ~n22905;
  assign n44011 = ~n44007 | ~n44006;
  assign n44009 = ~P1_INSTQUEUE_REG_10__3__SCAN_IN | ~n44047;
  assign n44008 = ~n44450 | ~n44039;
  assign n44010 = ~n44009 | ~n44008;
  assign n44013 = ~n44011 & ~n44010;
  assign n44012 = ~n44446 | ~n44042;
  assign P1_U3116 = ~n44013 | ~n44012;
  assign n44015 = ~n43147 | ~n44038;
  assign n44014 = ~n44461 | ~n44039;
  assign n44019 = ~n44015 | ~n44014;
  assign n44017 = ~n44457 | ~n44042;
  assign n44016 = ~n44460 | ~n22905;
  assign n44018 = ~n44017 | ~n44016;
  assign n44021 = ~n44019 & ~n44018;
  assign n44020 = ~P1_INSTQUEUE_REG_10__4__SCAN_IN | ~n44047;
  assign P1_U3117 = ~n44021 | ~n44020;
  assign n44023 = ~n44468 | ~n44038;
  assign n44022 = ~n44472 | ~n22905;
  assign n44027 = ~n44023 | ~n44022;
  assign n44025 = ~n44469 | ~n44042;
  assign n44024 = ~n44473 | ~n44039;
  assign n44026 = ~n44025 | ~n44024;
  assign n44029 = ~n44027 & ~n44026;
  assign n44028 = ~P1_INSTQUEUE_REG_10__5__SCAN_IN | ~n44047;
  assign P1_U3118 = ~n44029 | ~n44028;
  assign n44031 = ~n22825 | ~n44038;
  assign n44030 = ~n44483 | ~n22905;
  assign n44035 = ~n44031 | ~n44030;
  assign n44033 = ~n44480 | ~n44042;
  assign n44032 = ~n44484 | ~n44039;
  assign n44034 = ~n44033 | ~n44032;
  assign n44037 = ~n44035 & ~n44034;
  assign n44036 = ~P1_INSTQUEUE_REG_10__6__SCAN_IN | ~n44047;
  assign P1_U3119 = ~n44037 | ~n44036;
  assign n44041 = ~n44492 | ~n44038;
  assign n44040 = ~n44500 | ~n44039;
  assign n44046 = ~n44041 | ~n44040;
  assign n44044 = ~n44494 | ~n44042;
  assign n44043 = ~n44498 | ~n22905;
  assign n44045 = ~n44044 | ~n44043;
  assign n44049 = ~n44046 & ~n44045;
  assign n44048 = ~P1_INSTQUEUE_REG_10__7__SCAN_IN | ~n44047;
  assign P1_U3120 = ~n44049 | ~n44048;
  assign n44050 = ~n44058;
  assign n44121 = ~n44050 & ~n44308;
  assign n44057 = ~n44394 | ~n44121;
  assign n44055 = ~n44058 | ~P1_STATE2_REG_2__SCAN_IN;
  assign n44053 = ~n44051 | ~n44395;
  assign n44052 = ~n44121;
  assign n44060 = ~n44053 | ~n44052;
  assign n44054 = ~n44060 | ~n44399;
  assign n44122 = ~n44055 | ~n44054;
  assign n44056 = ~n44402 | ~n44122;
  assign n44068 = ~n44057 | ~n44056;
  assign n44059 = ~n44058 & ~n44399;
  assign n44064 = ~n44059 & ~n44415;
  assign n44762 = ~n44070;
  assign n44062 = ~n44762 | ~n44775;
  assign n44061 = ~n44060 & ~n44418;
  assign n44063 = ~n44062 | ~n44061;
  assign n44066 = ~P1_INSTQUEUE_REG_11__0__SCAN_IN | ~n44129;
  assign n44065 = ~n44406 | ~n22905;
  assign n44067 = ~n44066 | ~n44065;
  assign n44072 = ~n44068 & ~n44067;
  assign n44069 = ~n43066 | ~n44801;
  assign n44071 = ~n44405 | ~n44215;
  assign P1_U3121 = ~n44072 | ~n44071;
  assign n44074 = ~n43102 | ~n44121;
  assign n44073 = ~n44424 | ~n44122;
  assign n44078 = ~n44074 | ~n44073;
  assign n44076 = ~n44427 | ~n44215;
  assign n44075 = ~n44428 | ~n22905;
  assign n44077 = ~n44076 | ~n44075;
  assign n44080 = ~n44078 & ~n44077;
  assign n44079 = ~P1_INSTQUEUE_REG_11__1__SCAN_IN | ~n44129;
  assign P1_U3122 = ~n44080 | ~n44079;
  assign n44082 = ~n43117 | ~n44121;
  assign n44081 = ~n44435 | ~n44122;
  assign n44086 = ~n44082 | ~n44081;
  assign n44084 = ~n44438 | ~n44215;
  assign n44083 = ~n44439 | ~n22905;
  assign n44085 = ~n44084 | ~n44083;
  assign n44088 = ~n44086 & ~n44085;
  assign n44087 = ~P1_INSTQUEUE_REG_11__2__SCAN_IN | ~n44129;
  assign P1_U3123 = ~n44088 | ~n44087;
  assign n44090 = ~n43132 | ~n44121;
  assign n44089 = ~n44446 | ~n44122;
  assign n44094 = ~n44090 | ~n44089;
  assign n44092 = ~n44449 | ~n44215;
  assign n44091 = ~n44450 | ~n22905;
  assign n44093 = ~n44092 | ~n44091;
  assign n44096 = ~n44094 & ~n44093;
  assign n44095 = ~P1_INSTQUEUE_REG_11__3__SCAN_IN | ~n44129;
  assign P1_U3124 = ~n44096 | ~n44095;
  assign n44098 = ~n43147 | ~n44121;
  assign n44097 = ~n44457 | ~n44122;
  assign n44102 = ~n44098 | ~n44097;
  assign n44100 = ~n44460 | ~n44215;
  assign n44099 = ~n44461 | ~n22905;
  assign n44101 = ~n44100 | ~n44099;
  assign n44104 = ~n44102 & ~n44101;
  assign n44103 = ~P1_INSTQUEUE_REG_11__4__SCAN_IN | ~n44129;
  assign P1_U3125 = ~n44104 | ~n44103;
  assign n44106 = ~n44468 | ~n44121;
  assign n44105 = ~n44469 | ~n44122;
  assign n44110 = ~n44106 | ~n44105;
  assign n44108 = ~n44472 | ~n44215;
  assign n44107 = ~n44473 | ~n22905;
  assign n44109 = ~n44108 | ~n44107;
  assign n44112 = ~n44110 & ~n44109;
  assign n44111 = ~P1_INSTQUEUE_REG_11__5__SCAN_IN | ~n44129;
  assign P1_U3126 = ~n44112 | ~n44111;
  assign n44114 = ~n22825 | ~n44121;
  assign n44113 = ~n44480 | ~n44122;
  assign n44118 = ~n44114 | ~n44113;
  assign n44116 = ~n44483 | ~n44215;
  assign n44115 = ~n44484 | ~n22905;
  assign n44117 = ~n44116 | ~n44115;
  assign n44120 = ~n44118 & ~n44117;
  assign n44119 = ~P1_INSTQUEUE_REG_11__6__SCAN_IN | ~n44129;
  assign P1_U3127 = ~n44120 | ~n44119;
  assign n44124 = ~n44492 | ~n44121;
  assign n44123 = ~n44494 | ~n44122;
  assign n44128 = ~n44124 | ~n44123;
  assign n44126 = ~n44498 | ~n44215;
  assign n44125 = ~n44500 | ~n22905;
  assign n44127 = ~n44126 | ~n44125;
  assign n44131 = ~n44128 & ~n44127;
  assign n44130 = ~P1_INSTQUEUE_REG_11__7__SCAN_IN | ~n44129;
  assign P1_U3128 = ~n44131 | ~n44130;
  assign n44240 = ~n44133 & ~n44132;
  assign n44155 = ~n44240 | ~n44308;
  assign n44211 = ~n44155;
  assign n44135 = ~n44394 | ~n44211;
  assign n44761 = ~n44411 | ~n44792;
  assign n44134 = ~n44405 | ~n44298;
  assign n44149 = ~n44135 | ~n44134;
  assign n44310 = ~n44137 & ~n44136;
  assign n44145 = ~n44310 | ~n44152;
  assign n44139 = ~n44298;
  assign n44140 = ~n44139 | ~n44138;
  assign n44141 = ~n44140 | ~P1_STATEBS16_REG_SCAN_IN;
  assign n44151 = ~n44141 | ~n44399;
  assign n44143 = ~n44151;
  assign n44312 = n31479 | n44142;
  assign n44150 = ~n44312 & ~n31534;
  assign n44144 = ~n44143 | ~n44150;
  assign n44147 = ~n44402 | ~n44220;
  assign n44146 = ~n44406 | ~n44215;
  assign n44148 = ~n44147 | ~n44146;
  assign n44162 = ~n44149 & ~n44148;
  assign n44159 = ~n44151 & ~n44150;
  assign n44154 = ~n44153 | ~n44152;
  assign n44157 = ~n44154 | ~P1_STATE2_REG_2__SCAN_IN;
  assign n44156 = ~n44155 | ~P1_STATE2_REG_3__SCAN_IN;
  assign n44158 = ~n44157 | ~n44156;
  assign n44160 = ~n44159 & ~n44158;
  assign n44161 = ~P1_INSTQUEUE_REG_12__0__SCAN_IN | ~n44214;
  assign P1_U3129 = ~n44162 | ~n44161;
  assign n44164 = ~n43102 | ~n44211;
  assign n44163 = ~n44427 | ~n44298;
  assign n44168 = ~n44164 | ~n44163;
  assign n44166 = ~P1_INSTQUEUE_REG_12__1__SCAN_IN | ~n44214;
  assign n44165 = ~n44428 | ~n44215;
  assign n44167 = ~n44166 | ~n44165;
  assign n44170 = ~n44168 & ~n44167;
  assign n44169 = ~n44424 | ~n44220;
  assign P1_U3130 = ~n44170 | ~n44169;
  assign n44172 = ~n43117 | ~n44211;
  assign n44171 = ~n44438 | ~n44298;
  assign n44176 = ~n44172 | ~n44171;
  assign n44174 = ~n44435 | ~n44220;
  assign n44173 = ~n44439 | ~n44215;
  assign n44175 = ~n44174 | ~n44173;
  assign n44178 = ~n44176 & ~n44175;
  assign n44177 = ~P1_INSTQUEUE_REG_12__2__SCAN_IN | ~n44214;
  assign P1_U3131 = ~n44178 | ~n44177;
  assign n44180 = ~n43132 | ~n44211;
  assign n44179 = ~n44449 | ~n44298;
  assign n44184 = ~n44180 | ~n44179;
  assign n44182 = ~n44446 | ~n44220;
  assign n44181 = ~n44450 | ~n44215;
  assign n44183 = ~n44182 | ~n44181;
  assign n44186 = ~n44184 & ~n44183;
  assign n44185 = ~P1_INSTQUEUE_REG_12__3__SCAN_IN | ~n44214;
  assign P1_U3132 = ~n44186 | ~n44185;
  assign n44188 = ~n43147 | ~n44211;
  assign n44187 = ~n44460 | ~n44298;
  assign n44192 = ~n44188 | ~n44187;
  assign n44190 = ~n44457 | ~n44220;
  assign n44189 = ~n44461 | ~n44215;
  assign n44191 = ~n44190 | ~n44189;
  assign n44194 = ~n44192 & ~n44191;
  assign n44193 = ~P1_INSTQUEUE_REG_12__4__SCAN_IN | ~n44214;
  assign P1_U3133 = ~n44194 | ~n44193;
  assign n44196 = ~n44468 | ~n44211;
  assign n44195 = ~n44472 | ~n44298;
  assign n44200 = ~n44196 | ~n44195;
  assign n44198 = ~n44469 | ~n44220;
  assign n44197 = ~n44473 | ~n44215;
  assign n44199 = ~n44198 | ~n44197;
  assign n44202 = ~n44200 & ~n44199;
  assign n44201 = ~P1_INSTQUEUE_REG_12__5__SCAN_IN | ~n44214;
  assign P1_U3134 = ~n44202 | ~n44201;
  assign n44204 = ~n22825 | ~n44211;
  assign n44203 = ~n44483 | ~n44298;
  assign n44208 = ~n44204 | ~n44203;
  assign n44206 = ~n44480 | ~n44220;
  assign n44205 = ~n44484 | ~n44215;
  assign n44207 = ~n44206 | ~n44205;
  assign n44210 = ~n44208 & ~n44207;
  assign n44209 = ~P1_INSTQUEUE_REG_12__6__SCAN_IN | ~n44214;
  assign P1_U3135 = ~n44210 | ~n44209;
  assign n44213 = ~n44492 | ~n44211;
  assign n44212 = ~n44498 | ~n44298;
  assign n44219 = ~n44213 | ~n44212;
  assign n44217 = ~P1_INSTQUEUE_REG_12__7__SCAN_IN | ~n44214;
  assign n44216 = ~n44500 | ~n44215;
  assign n44218 = ~n44217 | ~n44216;
  assign n44222 = ~n44219 & ~n44218;
  assign n44221 = ~n44494 | ~n44220;
  assign P1_U3136 = ~n44222 | ~n44221;
  assign n44229 = ~n44394 | ~n44294;
  assign n44396 = ~n44312;
  assign n44225 = ~n44396 | ~n44223;
  assign n44224 = ~n44294;
  assign n44236 = ~n44225 | ~n44224;
  assign n44227 = ~n44236 | ~n44399;
  assign n44226 = ~n44240 | ~P1_STATE2_REG_2__SCAN_IN;
  assign n44295 = ~n44227 | ~n44226;
  assign n44228 = ~n44402 | ~n44295;
  assign n44235 = ~n44229 | ~n44228;
  assign n44231 = ~n44761 & ~n44230;
  assign n44386 = n44231;
  assign n44233 = ~n44405 | ~n44386;
  assign n44232 = ~n44406 | ~n44298;
  assign n44234 = ~n44233 | ~n44232;
  assign n44245 = ~n44235 & ~n44234;
  assign n44238 = ~n44761 & ~n44765;
  assign n44237 = n44236 | n44418;
  assign n44239 = ~n44238 & ~n44237;
  assign n44243 = ~n44239 & ~n44415;
  assign n44241 = ~n44240;
  assign n44242 = ~n44241 | ~n44418;
  assign n44244 = ~P1_INSTQUEUE_REG_13__0__SCAN_IN | ~n44303;
  assign P1_U3137 = ~n44245 | ~n44244;
  assign n44247 = ~n43102 | ~n44294;
  assign n44246 = ~n44424 | ~n44295;
  assign n44251 = ~n44247 | ~n44246;
  assign n44249 = ~n44427 | ~n44386;
  assign n44248 = ~n44428 | ~n44298;
  assign n44250 = ~n44249 | ~n44248;
  assign n44253 = ~n44251 & ~n44250;
  assign n44252 = ~P1_INSTQUEUE_REG_13__1__SCAN_IN | ~n44303;
  assign P1_U3138 = ~n44253 | ~n44252;
  assign n44255 = ~n43117 | ~n44294;
  assign n44254 = ~n44435 | ~n44295;
  assign n44259 = ~n44255 | ~n44254;
  assign n44257 = ~n44438 | ~n44386;
  assign n44256 = ~n44439 | ~n44298;
  assign n44258 = ~n44257 | ~n44256;
  assign n44261 = ~n44259 & ~n44258;
  assign n44260 = ~P1_INSTQUEUE_REG_13__2__SCAN_IN | ~n44303;
  assign P1_U3139 = ~n44261 | ~n44260;
  assign n44263 = ~n43132 | ~n44294;
  assign n44262 = ~n44446 | ~n44295;
  assign n44267 = ~n44263 | ~n44262;
  assign n44265 = ~n44449 | ~n44386;
  assign n44264 = ~n44450 | ~n44298;
  assign n44266 = ~n44265 | ~n44264;
  assign n44269 = ~n44267 & ~n44266;
  assign n44268 = ~P1_INSTQUEUE_REG_13__3__SCAN_IN | ~n44303;
  assign P1_U3140 = ~n44269 | ~n44268;
  assign n44271 = ~n43147 | ~n44294;
  assign n44270 = ~n44457 | ~n44295;
  assign n44275 = ~n44271 | ~n44270;
  assign n44273 = ~n44460 | ~n44386;
  assign n44272 = ~n44461 | ~n44298;
  assign n44274 = ~n44273 | ~n44272;
  assign n44277 = ~n44275 & ~n44274;
  assign n44276 = ~P1_INSTQUEUE_REG_13__4__SCAN_IN | ~n44303;
  assign P1_U3141 = ~n44277 | ~n44276;
  assign n44279 = ~n44468 | ~n44294;
  assign n44278 = ~n44469 | ~n44295;
  assign n44283 = ~n44279 | ~n44278;
  assign n44281 = ~n44472 | ~n44386;
  assign n44280 = ~n44473 | ~n44298;
  assign n44282 = ~n44281 | ~n44280;
  assign n44285 = ~n44283 & ~n44282;
  assign n44284 = ~P1_INSTQUEUE_REG_13__5__SCAN_IN | ~n44303;
  assign P1_U3142 = ~n44285 | ~n44284;
  assign n44287 = ~n22825 | ~n44294;
  assign n44286 = ~n44480 | ~n44295;
  assign n44291 = ~n44287 | ~n44286;
  assign n44289 = ~n44483 | ~n44386;
  assign n44288 = ~n44484 | ~n44298;
  assign n44290 = ~n44289 | ~n44288;
  assign n44293 = ~n44291 & ~n44290;
  assign n44292 = ~P1_INSTQUEUE_REG_13__6__SCAN_IN | ~n44303;
  assign P1_U3143 = ~n44293 | ~n44292;
  assign n44297 = ~n44492 | ~n44294;
  assign n44296 = ~n44494 | ~n44295;
  assign n44302 = ~n44297 | ~n44296;
  assign n44300 = ~n44498 | ~n44386;
  assign n44299 = ~n44500 | ~n44298;
  assign n44301 = ~n44300 | ~n44299;
  assign n44305 = ~n44302 & ~n44301;
  assign n44304 = ~P1_INSTQUEUE_REG_13__7__SCAN_IN | ~n44303;
  assign P1_U3144 = ~n44305 | ~n44304;
  assign n44417 = ~n44307 & ~n44306;
  assign n44316 = ~n44394 | ~n44382;
  assign n44314 = ~n44310 | ~n44309;
  assign n44319 = ~n44312 & ~n44311;
  assign n44313 = ~n44319 | ~n44399;
  assign n44383 = ~n44314 | ~n44313;
  assign n44315 = ~n44402 | ~n44383;
  assign n44331 = ~n44316 | ~n44315;
  assign n44329 = ~n44405 | ~n44499;
  assign n44318 = ~n44386 & ~n44499;
  assign n44320 = ~n44318 & ~n44765;
  assign n44321 = ~n44320 & ~n44319;
  assign n44322 = ~P1_STATE2_REG_3__SCAN_IN & ~n44321;
  assign n44325 = ~n44382 & ~n44322;
  assign n44324 = ~n44323;
  assign n44328 = ~P1_INSTQUEUE_REG_14__0__SCAN_IN | ~n44391;
  assign n44330 = ~n44329 | ~n44328;
  assign n44333 = ~n44331 & ~n44330;
  assign n44332 = ~n44406 | ~n44386;
  assign P1_U3145 = ~n44333 | ~n44332;
  assign n44335 = ~n43102 | ~n44382;
  assign n44334 = ~n44424 | ~n44383;
  assign n44339 = ~n44335 | ~n44334;
  assign n44337 = ~n44427 | ~n44499;
  assign n44336 = ~n44428 | ~n44386;
  assign n44338 = ~n44337 | ~n44336;
  assign n44341 = ~n44339 & ~n44338;
  assign n44340 = ~P1_INSTQUEUE_REG_14__1__SCAN_IN | ~n44391;
  assign P1_U3146 = ~n44341 | ~n44340;
  assign n44343 = ~n43117 | ~n44382;
  assign n44342 = ~n44435 | ~n44383;
  assign n44347 = ~n44343 | ~n44342;
  assign n44345 = ~n44438 | ~n44499;
  assign n44344 = ~n44439 | ~n44386;
  assign n44346 = ~n44345 | ~n44344;
  assign n44349 = ~n44347 & ~n44346;
  assign n44348 = ~P1_INSTQUEUE_REG_14__2__SCAN_IN | ~n44391;
  assign P1_U3147 = ~n44349 | ~n44348;
  assign n44351 = ~n43132 | ~n44382;
  assign n44350 = ~n44446 | ~n44383;
  assign n44355 = ~n44351 | ~n44350;
  assign n44353 = ~n44449 | ~n44499;
  assign n44352 = ~n44450 | ~n44386;
  assign n44354 = ~n44353 | ~n44352;
  assign n44357 = ~n44355 & ~n44354;
  assign n44356 = ~P1_INSTQUEUE_REG_14__3__SCAN_IN | ~n44391;
  assign P1_U3148 = ~n44357 | ~n44356;
  assign n44359 = ~n43147 | ~n44382;
  assign n44358 = ~n44457 | ~n44383;
  assign n44363 = ~n44359 | ~n44358;
  assign n44361 = ~n44460 | ~n44499;
  assign n44360 = ~n44461 | ~n44386;
  assign n44362 = ~n44361 | ~n44360;
  assign n44365 = ~n44363 & ~n44362;
  assign n44364 = ~P1_INSTQUEUE_REG_14__4__SCAN_IN | ~n44391;
  assign P1_U3149 = ~n44365 | ~n44364;
  assign n44367 = ~n44468 | ~n44382;
  assign n44366 = ~n44469 | ~n44383;
  assign n44371 = ~n44367 | ~n44366;
  assign n44369 = ~n44472 | ~n44499;
  assign n44368 = ~n44473 | ~n44386;
  assign n44370 = ~n44369 | ~n44368;
  assign n44373 = ~n44371 & ~n44370;
  assign n44372 = ~P1_INSTQUEUE_REG_14__5__SCAN_IN | ~n44391;
  assign P1_U3150 = ~n44373 | ~n44372;
  assign n44375 = ~n22825 | ~n44382;
  assign n44374 = ~n44480 | ~n44383;
  assign n44379 = ~n44375 | ~n44374;
  assign n44377 = ~n44483 | ~n44499;
  assign n44376 = ~n44484 | ~n44386;
  assign n44378 = ~n44377 | ~n44376;
  assign n44381 = ~n44379 & ~n44378;
  assign n44380 = ~P1_INSTQUEUE_REG_14__6__SCAN_IN | ~n44391;
  assign P1_U3151 = ~n44381 | ~n44380;
  assign n44385 = ~n44492 | ~n44382;
  assign n44384 = ~n44494 | ~n44383;
  assign n44390 = ~n44385 | ~n44384;
  assign n44388 = ~n44498 | ~n44499;
  assign n44387 = ~n44500 | ~n44386;
  assign n44389 = ~n44388 | ~n44387;
  assign n44393 = ~n44390 & ~n44389;
  assign n44392 = ~P1_INSTQUEUE_REG_14__7__SCAN_IN | ~n44391;
  assign P1_U3152 = ~n44393 | ~n44392;
  assign n44404 = ~n44394 | ~n44491;
  assign n44398 = ~n44396 | ~n44395;
  assign n44397 = ~n44491;
  assign n44412 = ~n44398 | ~n44397;
  assign n44401 = ~n44412 | ~n44399;
  assign n44400 = ~n44417 | ~P1_STATE2_REG_2__SCAN_IN;
  assign n44493 = ~n44401 | ~n44400;
  assign n44403 = ~n44402 | ~n44493;
  assign n44410 = ~n44404 | ~n44403;
  assign n44408 = ~n44405 | ~n43067;
  assign n44407 = ~n44406 | ~n44499;
  assign n44409 = ~n44408 | ~n44407;
  assign n44423 = ~n44410 & ~n44409;
  assign n44414 = n44411 & n44775;
  assign n44413 = n44412 | n44418;
  assign n44416 = ~n44414 & ~n44413;
  assign n44421 = ~n44416 & ~n44415;
  assign n44419 = ~n44417;
  assign n44420 = ~n44419 | ~n44418;
  assign n44422 = ~P1_INSTQUEUE_REG_15__0__SCAN_IN | ~n44505;
  assign P1_U3153 = ~n44423 | ~n44422;
  assign n44426 = ~n43102 | ~n44491;
  assign n44425 = ~n44424 | ~n44493;
  assign n44432 = ~n44426 | ~n44425;
  assign n44430 = ~n44427 | ~n43067;
  assign n44429 = ~n44428 | ~n44499;
  assign n44431 = ~n44430 | ~n44429;
  assign n44434 = ~n44432 & ~n44431;
  assign n44433 = ~P1_INSTQUEUE_REG_15__1__SCAN_IN | ~n44505;
  assign P1_U3154 = ~n44434 | ~n44433;
  assign n44437 = ~n43117 | ~n44491;
  assign n44436 = ~n44435 | ~n44493;
  assign n44443 = ~n44437 | ~n44436;
  assign n44441 = ~n44438 | ~n43067;
  assign n44440 = ~n44439 | ~n44499;
  assign n44442 = ~n44441 | ~n44440;
  assign n44445 = ~n44443 & ~n44442;
  assign n44444 = ~P1_INSTQUEUE_REG_15__2__SCAN_IN | ~n44505;
  assign P1_U3155 = ~n44445 | ~n44444;
  assign n44448 = ~n43132 | ~n44491;
  assign n44447 = ~n44446 | ~n44493;
  assign n44454 = ~n44448 | ~n44447;
  assign n44452 = ~n44449 | ~n43067;
  assign n44451 = ~n44450 | ~n44499;
  assign n44453 = ~n44452 | ~n44451;
  assign n44456 = ~n44454 & ~n44453;
  assign n44455 = ~P1_INSTQUEUE_REG_15__3__SCAN_IN | ~n44505;
  assign P1_U3156 = ~n44456 | ~n44455;
  assign n44459 = ~n43147 | ~n44491;
  assign n44458 = ~n44457 | ~n44493;
  assign n44465 = ~n44459 | ~n44458;
  assign n44463 = ~n44460 | ~n43067;
  assign n44462 = ~n44461 | ~n44499;
  assign n44464 = ~n44463 | ~n44462;
  assign n44467 = ~n44465 & ~n44464;
  assign n44466 = ~P1_INSTQUEUE_REG_15__4__SCAN_IN | ~n44505;
  assign P1_U3157 = ~n44467 | ~n44466;
  assign n44471 = ~n44468 | ~n44491;
  assign n44470 = ~n44469 | ~n44493;
  assign n44477 = ~n44471 | ~n44470;
  assign n44475 = ~n44472 | ~n43067;
  assign n44474 = ~n44473 | ~n44499;
  assign n44476 = ~n44475 | ~n44474;
  assign n44479 = ~n44477 & ~n44476;
  assign n44478 = ~P1_INSTQUEUE_REG_15__5__SCAN_IN | ~n44505;
  assign P1_U3158 = ~n44479 | ~n44478;
  assign n44482 = ~n22825 | ~n44491;
  assign n44481 = ~n44480 | ~n44493;
  assign n44488 = ~n44482 | ~n44481;
  assign n44486 = ~n44483 | ~n43067;
  assign n44485 = ~n44484 | ~n44499;
  assign n44487 = ~n44486 | ~n44485;
  assign n44490 = ~n44488 & ~n44487;
  assign n44489 = ~P1_INSTQUEUE_REG_15__6__SCAN_IN | ~n44505;
  assign P1_U3159 = ~n44490 | ~n44489;
  assign n44496 = ~n44492 | ~n44491;
  assign n44495 = ~n44494 | ~n44493;
  assign n44504 = ~n44496 | ~n44495;
  assign n44502 = ~n44498 | ~n43067;
  assign n44501 = ~n44500 | ~n44499;
  assign n44503 = ~n44502 | ~n44501;
  assign n44507 = ~n44504 & ~n44503;
  assign n44506 = ~P1_INSTQUEUE_REG_15__7__SCAN_IN | ~n44505;
  assign P1_U3160 = ~n44507 | ~n44506;
  assign n44806 = ~n44509 & ~n44508;
  assign n44511 = ~n44853 & ~n44750;
  assign n44513 = ~n44512 & ~n44511;
  assign n44516 = ~n44515 | ~n44514;
  assign n44518 = ~n44517 | ~P1_STATE2_REG_1__SCAN_IN;
  assign n44520 = ~n44518 | ~P1_STATE2_REG_2__SCAN_IN;
  assign P1_U3163 = ~n44520 | ~n44519;
  assign P1_U3164 = P1_DATAWIDTH_REG_31__SCAN_IN & n44709;
  assign P1_U3165 = P1_DATAWIDTH_REG_30__SCAN_IN & n44521;
  assign P1_U3166 = P1_DATAWIDTH_REG_29__SCAN_IN & n44709;
  assign P1_U3167 = P1_DATAWIDTH_REG_28__SCAN_IN & n44521;
  assign P1_U3168 = P1_DATAWIDTH_REG_27__SCAN_IN & n44521;
  assign P1_U3169 = P1_DATAWIDTH_REG_26__SCAN_IN & n44521;
  assign P1_U3170 = P1_DATAWIDTH_REG_25__SCAN_IN & n44521;
  assign P1_U3171 = P1_DATAWIDTH_REG_24__SCAN_IN & n44521;
  assign P1_U3172 = P1_DATAWIDTH_REG_23__SCAN_IN & n44521;
  assign P1_U3173 = P1_DATAWIDTH_REG_22__SCAN_IN & n44521;
  assign P1_U3174 = P1_DATAWIDTH_REG_21__SCAN_IN & n44521;
  assign P1_U3175 = P1_DATAWIDTH_REG_20__SCAN_IN & n44521;
  assign P1_U3176 = P1_DATAWIDTH_REG_19__SCAN_IN & n44521;
  assign P1_U3177 = P1_DATAWIDTH_REG_18__SCAN_IN & n44521;
  assign P1_U3178 = P1_DATAWIDTH_REG_17__SCAN_IN & n44521;
  assign P1_U3179 = P1_DATAWIDTH_REG_16__SCAN_IN & n44521;
  assign P1_U3180 = P1_DATAWIDTH_REG_15__SCAN_IN & n44521;
  assign P1_U3181 = P1_DATAWIDTH_REG_14__SCAN_IN & n44709;
  assign P1_U3182 = P1_DATAWIDTH_REG_13__SCAN_IN & n44709;
  assign P1_U3183 = P1_DATAWIDTH_REG_12__SCAN_IN & n44709;
  assign P1_U3184 = P1_DATAWIDTH_REG_11__SCAN_IN & n44709;
  assign P1_U3185 = P1_DATAWIDTH_REG_10__SCAN_IN & n44709;
  assign P1_U3186 = P1_DATAWIDTH_REG_9__SCAN_IN & n44521;
  assign P1_U3187 = P1_DATAWIDTH_REG_8__SCAN_IN & n44709;
  assign P1_U3188 = P1_DATAWIDTH_REG_7__SCAN_IN & n44709;
  assign P1_U3189 = P1_DATAWIDTH_REG_6__SCAN_IN & n44709;
  assign P1_U3190 = P1_DATAWIDTH_REG_5__SCAN_IN & n44709;
  assign P1_U3191 = P1_DATAWIDTH_REG_4__SCAN_IN & n44709;
  assign P1_U3192 = P1_DATAWIDTH_REG_3__SCAN_IN & n44709;
  assign P1_U3193 = P1_DATAWIDTH_REG_2__SCAN_IN & n44709;
  assign n44533 = ~P1_REQUESTPENDING_REG_SCAN_IN;
  assign n44525 = ~NA | ~n44522;
  assign n44524 = ~n44523 | ~HOLD;
  assign n44526 = ~n44525 | ~n44524;
  assign n44527 = ~n44533 & ~n44526;
  assign n44529 = ~n44859 & ~n44527;
  assign n44541 = n44530 & P1_STATE_REG_0__SCAN_IN;
  assign n44528 = ~P1_STATE_REG_2__SCAN_IN & ~n44541;
  assign P1_U3194 = n44529 | n44528;
  assign n44531 = ~NA & ~n44530;
  assign n44538 = ~n44531 | ~P1_REQUESTPENDING_REG_SCAN_IN;
  assign n44532 = ~n44850 | ~n44540;
  assign n44534 = ~P1_STATE_REG_1__SCAN_IN | ~n44532;
  assign n44535 = ~n44534 | ~n44533;
  assign n44536 = ~n44535 | ~n44546;
  assign n44537 = ~n44536 | ~HOLD;
  assign n44539 = ~n44538 | ~n44537;
  assign n44545 = ~n44539 | ~P1_STATE_REG_0__SCAN_IN;
  assign n44542 = ~P1_STATE_REG_1__SCAN_IN & ~n44540;
  assign n44543 = ~n44542 & ~n44541;
  assign n44544 = ~P1_STATE_REG_2__SCAN_IN | ~n44543;
  assign P1_U3196 = ~n44545 | ~n44544;
  assign n44548 = ~n44597 & ~n44551;
  assign n44547 = ~n44815 & ~n44691;
  assign n44550 = ~n44548 & ~n44547;
  assign n44549 = ~P1_ADDRESS_REG_0__SCAN_IN | ~n44828;
  assign P1_U3197 = ~n44550 | ~n44549;
  assign n44553 = ~n44551 & ~n44691;
  assign n44552 = ~n44597 & ~n44556;
  assign n44555 = ~n44553 & ~n44552;
  assign n44554 = ~P1_ADDRESS_REG_1__SCAN_IN | ~n44828;
  assign P1_U3198 = ~n44555 | ~n44554;
  assign n44561 = ~P1_REIP_REG_4__SCAN_IN;
  assign n44558 = ~n44597 & ~n44561;
  assign n44557 = ~n44556 & ~n44691;
  assign n44560 = ~n44558 & ~n44557;
  assign n44559 = ~P1_ADDRESS_REG_2__SCAN_IN | ~n44828;
  assign P1_U3199 = ~n44560 | ~n44559;
  assign n44563 = ~n44561 & ~n44691;
  assign n44562 = ~n44597 & ~n44566;
  assign n44565 = ~n44563 & ~n44562;
  assign n44564 = ~P1_ADDRESS_REG_3__SCAN_IN | ~n44828;
  assign P1_U3200 = ~n44565 | ~n44564;
  assign n44568 = ~n44566 & ~n44691;
  assign n44567 = ~n44597 & ~n44571;
  assign n44570 = ~n44568 & ~n44567;
  assign n44569 = ~P1_ADDRESS_REG_4__SCAN_IN | ~n44828;
  assign P1_U3201 = ~n44570 | ~n44569;
  assign n44573 = ~n44571 & ~n44691;
  assign n44572 = ~n44597 & ~n44576;
  assign n44575 = ~n44573 & ~n44572;
  assign n44574 = ~P1_ADDRESS_REG_5__SCAN_IN | ~n44828;
  assign P1_U3202 = ~n44575 | ~n44574;
  assign n44580 = ~P1_ADDRESS_REG_6__SCAN_IN | ~n44828;
  assign n44581 = ~P1_REIP_REG_8__SCAN_IN;
  assign n44578 = ~n44597 & ~n44581;
  assign n44577 = ~n44576 & ~n44691;
  assign n44579 = ~n44578 & ~n44577;
  assign P1_U3203 = ~n44580 | ~n44579;
  assign n44583 = ~n44581 & ~n44691;
  assign n44582 = ~n44597 & ~n44586;
  assign n44585 = ~n44583 & ~n44582;
  assign n44584 = ~P1_ADDRESS_REG_7__SCAN_IN | ~n44828;
  assign P1_U3204 = ~n44585 | ~n44584;
  assign n44588 = ~n44586 & ~n44691;
  assign n44587 = ~n44597 & ~n44591;
  assign n44590 = ~n44588 & ~n44587;
  assign n44589 = ~P1_ADDRESS_REG_8__SCAN_IN | ~n44828;
  assign P1_U3205 = ~n44590 | ~n44589;
  assign n44593 = ~n44597 & ~n44596;
  assign n44592 = ~n44591 & ~n44691;
  assign n44595 = ~n44593 & ~n44592;
  assign n44594 = ~P1_ADDRESS_REG_9__SCAN_IN | ~n44828;
  assign P1_U3206 = ~n44595 | ~n44594;
  assign n44599 = ~n44596 & ~n44691;
  assign n44598 = ~n44597 & ~n44602;
  assign n44601 = ~n44599 & ~n44598;
  assign n44600 = ~P1_ADDRESS_REG_10__SCAN_IN | ~n44828;
  assign P1_U3207 = ~n44601 | ~n44600;
  assign n44604 = ~n44597 & ~n30890;
  assign n44603 = ~n44602 & ~n44691;
  assign n44606 = ~n44604 & ~n44603;
  assign n44605 = ~P1_ADDRESS_REG_11__SCAN_IN | ~n44828;
  assign P1_U3208 = ~n44606 | ~n44605;
  assign n44608 = ~n30890 & ~n44691;
  assign n44607 = ~n44597 & ~n44611;
  assign n44610 = ~n44608 & ~n44607;
  assign n44609 = ~P1_ADDRESS_REG_12__SCAN_IN | ~n44828;
  assign P1_U3209 = ~n44610 | ~n44609;
  assign n44613 = ~n44611 & ~n44691;
  assign n44612 = ~n44597 & ~n44616;
  assign n44615 = ~n44613 & ~n44612;
  assign n44614 = ~P1_ADDRESS_REG_13__SCAN_IN | ~n44828;
  assign P1_U3210 = ~n44615 | ~n44614;
  assign n44618 = ~n44616 & ~n44691;
  assign n44617 = ~n44597 & ~n44621;
  assign n44620 = ~n44618 & ~n44617;
  assign n44619 = ~P1_ADDRESS_REG_14__SCAN_IN | ~n44828;
  assign P1_U3211 = ~n44620 | ~n44619;
  assign n44623 = ~n44621 & ~n44691;
  assign n44626 = ~P1_REIP_REG_17__SCAN_IN;
  assign n44622 = ~n44597 & ~n44626;
  assign n44625 = ~n44623 & ~n44622;
  assign n44624 = ~P1_ADDRESS_REG_15__SCAN_IN | ~n44828;
  assign P1_U3212 = ~n44625 | ~n44624;
  assign n44630 = ~P1_ADDRESS_REG_16__SCAN_IN | ~n44828;
  assign n44631 = ~P1_REIP_REG_18__SCAN_IN;
  assign n44628 = ~n44597 & ~n44631;
  assign n44627 = ~n44626 & ~n44691;
  assign n44629 = ~n44628 & ~n44627;
  assign P1_U3213 = ~n44630 | ~n44629;
  assign n44633 = ~n44631 & ~n44691;
  assign n44632 = ~n44597 & ~n44636;
  assign n44635 = ~n44633 & ~n44632;
  assign n44634 = ~P1_ADDRESS_REG_17__SCAN_IN | ~n44828;
  assign P1_U3214 = ~n44635 | ~n44634;
  assign n44638 = ~n44636 & ~n44691;
  assign n44637 = ~n44597 & ~n44641;
  assign n44640 = ~n44638 & ~n44637;
  assign n44639 = ~P1_ADDRESS_REG_18__SCAN_IN | ~n44828;
  assign P1_U3215 = ~n44640 | ~n44639;
  assign n44643 = ~n44641 & ~n44691;
  assign n44642 = ~n44597 & ~n44646;
  assign n44645 = ~n44643 & ~n44642;
  assign n44644 = ~P1_ADDRESS_REG_19__SCAN_IN | ~n44828;
  assign P1_U3216 = ~n44645 | ~n44644;
  assign n44648 = ~n44646 & ~n44691;
  assign n44647 = ~n44597 & ~n44651;
  assign n44650 = ~n44648 & ~n44647;
  assign n44649 = ~P1_ADDRESS_REG_20__SCAN_IN | ~n44828;
  assign P1_U3217 = ~n44650 | ~n44649;
  assign n44653 = ~n44651 & ~n44691;
  assign n44656 = ~P1_REIP_REG_23__SCAN_IN;
  assign n44652 = ~n44597 & ~n44656;
  assign n44655 = ~n44653 & ~n44652;
  assign n44654 = ~P1_ADDRESS_REG_21__SCAN_IN | ~n44828;
  assign P1_U3218 = ~n44655 | ~n44654;
  assign n44658 = ~n44656 & ~n44691;
  assign n44657 = ~n44597 & ~n44661;
  assign n44660 = ~n44658 & ~n44657;
  assign n44659 = ~P1_ADDRESS_REG_22__SCAN_IN | ~n44828;
  assign P1_U3219 = ~n44660 | ~n44659;
  assign n44663 = ~n44661 & ~n44691;
  assign n44662 = ~n44597 & ~n44666;
  assign n44665 = ~n44663 & ~n44662;
  assign n44664 = ~P1_ADDRESS_REG_23__SCAN_IN | ~n44828;
  assign P1_U3220 = ~n44665 | ~n44664;
  assign n44668 = ~n44597 & ~n44671;
  assign n44667 = ~n44666 & ~n44691;
  assign n44670 = ~n44668 & ~n44667;
  assign n44669 = ~P1_ADDRESS_REG_24__SCAN_IN | ~n44828;
  assign P1_U3221 = ~n44670 | ~n44669;
  assign n44673 = ~n44671 & ~n44691;
  assign n44672 = ~n44597 & ~n44676;
  assign n44675 = ~n44673 & ~n44672;
  assign n44674 = ~P1_ADDRESS_REG_25__SCAN_IN | ~n44828;
  assign P1_U3222 = ~n44675 | ~n44674;
  assign n44678 = ~n44597 & ~n44681;
  assign n44677 = ~n44676 & ~n44691;
  assign n44680 = ~n44678 & ~n44677;
  assign n44679 = ~P1_ADDRESS_REG_26__SCAN_IN | ~n44828;
  assign P1_U3223 = ~n44680 | ~n44679;
  assign n44683 = ~n44681 & ~n44691;
  assign n44682 = ~n44597 & ~n44686;
  assign n44685 = ~n44683 & ~n44682;
  assign n44684 = ~P1_ADDRESS_REG_27__SCAN_IN | ~n44828;
  assign P1_U3224 = ~n44685 | ~n44684;
  assign n44690 = ~P1_ADDRESS_REG_28__SCAN_IN | ~n44828;
  assign n44688 = ~n44597 & ~n44692;
  assign n44687 = ~n44686 & ~n44691;
  assign n44689 = ~n44688 & ~n44687;
  assign P1_U3225 = ~n44690 | ~n44689;
  assign n44695 = ~n44692 & ~n44691;
  assign n44693 = ~P1_REIP_REG_31__SCAN_IN;
  assign n44694 = ~n44597 & ~n44693;
  assign n44697 = ~n44695 & ~n44694;
  assign n44696 = ~P1_ADDRESS_REG_29__SCAN_IN | ~n44828;
  assign P1_U3226 = ~n44697 | ~n44696;
  assign n44699 = ~n44828 | ~P1_BE_N_REG_3__SCAN_IN;
  assign n44698 = ~n44859 | ~P1_BYTEENABLE_REG_3__SCAN_IN;
  assign P1_U3458 = ~n44699 | ~n44698;
  assign n44701 = ~n44828 | ~P1_BE_N_REG_2__SCAN_IN;
  assign n44700 = ~n44859 | ~P1_BYTEENABLE_REG_2__SCAN_IN;
  assign P1_U3459 = ~n44701 | ~n44700;
  assign n44703 = ~n44828 | ~P1_BE_N_REG_1__SCAN_IN;
  assign n44702 = ~n44859 | ~P1_BYTEENABLE_REG_1__SCAN_IN;
  assign P1_U3460 = ~n44703 | ~n44702;
  assign n44705 = ~n44828 | ~P1_BE_N_REG_0__SCAN_IN;
  assign n44704 = ~n44859 | ~P1_BYTEENABLE_REG_0__SCAN_IN;
  assign P1_U3461 = ~n44705 | ~n44704;
  assign n44708 = ~n44711;
  assign n44707 = ~P1_DATAWIDTH_REG_0__SCAN_IN & ~n44706;
  assign P1_U3464 = ~n44708 & ~n44707;
  assign n44710 = ~P1_DATAWIDTH_REG_1__SCAN_IN | ~n44709;
  assign P1_U3465 = ~n44711 | ~n44710;
  assign n44715 = n44750 | n44712;
  assign n44714 = ~n44713 | ~n44744;
  assign n44716 = ~n44715 | ~n44714;
  assign n44718 = ~n44716 | ~n44757;
  assign n44717 = ~n44741 | ~P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN;
  assign P1_U3469 = ~n44718 | ~n44717;
  assign n44731 = ~n44750;
  assign n44720 = ~n44719;
  assign n44725 = ~n44731 | ~n44720;
  assign n44723 = n44721 & n44744;
  assign n44733 = P1_INSTADDRPOINTER_REG_31__SCAN_IN ^ n25405;
  assign n44734 = ~P1_STATE2_REG_1__SCAN_IN | ~P1_INSTADDRPOINTER_REG_0__SCAN_IN;
  assign n44722 = ~n44733 & ~n44734;
  assign n44724 = ~n44723 & ~n44722;
  assign n44726 = ~n44725 | ~n44724;
  assign n44728 = ~n44757 | ~n44726;
  assign n44727 = ~n44741 | ~P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN;
  assign P1_U3472 = ~n44728 | ~n44727;
  assign n44730 = ~n44729;
  assign n44739 = ~n44731 | ~n44730;
  assign n44737 = n44732 & n44744;
  assign n44735 = ~n44733;
  assign n44736 = ~n44735 & ~n44734;
  assign n44738 = ~n44737 & ~n44736;
  assign n44740 = ~n44739 | ~n44738;
  assign n44743 = ~n44757 | ~n44740;
  assign n44742 = ~n44741 | ~P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN;
  assign P1_U3473 = ~n44743 | ~n44742;
  assign n44746 = ~n44745 | ~n44744;
  assign n44747 = ~n44757 | ~n44746;
  assign n44759 = ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN | ~n44747;
  assign n44752 = ~n44749 & ~n44748;
  assign n44751 = ~P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN & ~n44750;
  assign n44755 = ~n44752 & ~n44751;
  assign n44754 = ~P1_STATE2_REG_1__SCAN_IN | ~n44753;
  assign n44756 = ~n44755 | ~n44754;
  assign n44758 = ~n44757 | ~n44756;
  assign P1_U3474 = ~n44759 | ~n44758;
  assign n44774 = ~P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN | ~n44809;
  assign n44763 = ~n44761 | ~n44760;
  assign n44764 = ~n44763 & ~n44762;
  assign n44771 = ~n44791 & ~n44764;
  assign n44790 = n44800 & n44765;
  assign n44769 = ~n43072 | ~n44790;
  assign n44802 = ~n44766 | ~P1_STATE2_REG_1__SCAN_IN;
  assign n44768 = ~n23619 | ~n44802;
  assign n44770 = ~n44769 | ~n44768;
  assign n44772 = ~n44771 & ~n44770;
  assign n44773 = n44809 | n44772;
  assign P1_U3475 = ~n44774 | ~n44773;
  assign n44776 = ~n44775;
  assign n44777 = ~n44776 | ~n44800;
  assign n44783 = ~n44778 | ~n44777;
  assign n44779 = ~n44791;
  assign n44780 = ~n43066 | ~n44779;
  assign n44782 = ~n44781 | ~n44780;
  assign n44786 = ~n44783 | ~n44782;
  assign n44785 = ~n44784 | ~n44802;
  assign n44787 = ~n44786 | ~n44785;
  assign n44789 = ~n44808 | ~n44787;
  assign n44788 = ~P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN | ~n44809;
  assign P1_U3476 = ~n44789 | ~n44788;
  assign n44794 = n44792 | n44790;
  assign n44793 = ~n44792 | ~n44791;
  assign n44796 = ~n44794 | ~n44793;
  assign n44795 = ~n31534 | ~n44802;
  assign n44797 = ~n44796 | ~n44795;
  assign n44799 = ~n44808 | ~n44797;
  assign n44798 = ~n44809 | ~P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN;
  assign P1_U3477 = ~n44799 | ~n44798;
  assign n44804 = ~n44801 | ~n44800;
  assign n44803 = ~n23393 | ~n44802;
  assign n44805 = ~n44804 | ~n44803;
  assign n44807 = n44806 | n44805;
  assign n44811 = ~n44808 | ~n44807;
  assign n44810 = ~n44809 | ~P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN;
  assign P1_U3478 = ~n44811 | ~n44810;
  assign n44822 = ~n44823 | ~P1_BYTEENABLE_REG_2__SCAN_IN;
  assign n44819 = ~n44812 | ~n44813;
  assign n44824 = ~n44815 | ~n44814;
  assign n44817 = ~n44813 & ~n44824;
  assign n44816 = ~n44815 & ~n44814;
  assign n44818 = ~n44817 & ~n44816;
  assign n44820 = ~n44819 | ~n44818;
  assign n44825 = ~n44823;
  assign n44821 = ~n44820 | ~n44825;
  assign P1_U3481 = ~n44822 | ~n44821;
  assign n44827 = ~n44823 | ~P1_BYTEENABLE_REG_0__SCAN_IN;
  assign n44826 = ~n44825 | ~n44824;
  assign P1_U3482 = ~n44827 | ~n44826;
  assign n44830 = ~P1_W_R_N_REG_SCAN_IN | ~n44828;
  assign n44829 = n44828 | P1_READREQUEST_REG_SCAN_IN;
  assign P1_U3483 = ~n44830 | ~n44829;
  assign n44834 = ~P1_MORE_REG_SCAN_IN | ~n44831;
  assign n44833 = n44832 | n44831;
  assign P1_U3484 = ~n44834 | ~n44833;
  assign n44836 = ~n44835;
  assign n44840 = ~n44836 & ~n44850;
  assign n44839 = n44838 | n44837;
  assign n44856 = ~n44840 & ~n44839;
  assign n44858 = ~P1_REQUESTPENDING_REG_SCAN_IN | ~n44856;
  assign n44844 = ~n44842 | ~n44841;
  assign n44847 = ~n44844 | ~n44843;
  assign n44846 = ~n44845 | ~P1_STATEBS16_REG_SCAN_IN;
  assign n44848 = ~n44847 | ~n44846;
  assign n44849 = ~n44848 | ~P1_STATE2_REG_2__SCAN_IN;
  assign n44852 = ~n44850 & ~n44849;
  assign n44854 = n44852 | n44851;
  assign n44855 = n44854 & n44853;
  assign n44857 = n44856 | n44855;
  assign P1_U3485 = ~n44858 | ~n44857;
  assign n44861 = ~n44828 | ~P1_M_IO_N_REG_SCAN_IN;
  assign n44860 = ~n44859 | ~P1_MEMORYFETCH_REG_SCAN_IN;
  assign P1_U3486 = ~n44861 | ~n44860;
  assign n34993 = ~n34610;
  assign n36497 = ~n36610;
  assign n23304 = n25411 & n25233;
  assign n37463 = ~n24326 & ~n24325;
  assign n30741 = n30054 ^ n30053;
  assign n44863 = n43191 | n25042;
  assign n44864 = n25011 | n25014;
  assign n44865 = ~n42622;
  assign n30615 = ~n42625 & ~n30602;
endmodule


