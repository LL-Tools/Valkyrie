

module b14_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, U3352, U3351, U3350, U3349, 
        U3348, U3347, U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, 
        U3338, U3337, U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, 
        U3328, U3327, U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, 
        U3320, U3319, U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, 
        U3310, U3309, U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, 
        U3300, U3299, U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, 
        U3467, U3469, U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, 
        U3487, U3489, U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, 
        U3506, U3507, U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, 
        U3516, U3517, U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, 
        U3526, U3527, U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, 
        U3536, U3537, U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, 
        U3546, U3547, U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, 
        U3284, U3283, U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, 
        U3274, U3273, U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, 
        U3264, U3263, U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, 
        U3255, U3254, U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, 
        U3245, U3244, U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, 
        U3554, U3555, U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, 
        U3564, U3565, U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, 
        U3574, U3575, U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, 
        U3237, U3236, U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, 
        U3227, U3226, U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, 
        U3217, U3216, U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, 
        U4043, keyinput63, keyinput62, keyinput61, keyinput60, keyinput59, 
        keyinput58, keyinput57, keyinput56, keyinput55, keyinput54, keyinput53, 
        keyinput52, keyinput51, keyinput50, keyinput49, keyinput48, keyinput47, 
        keyinput46, keyinput45, keyinput44, keyinput43, keyinput42, keyinput41, 
        keyinput40, keyinput39, keyinput38, keyinput37, keyinput36, keyinput35, 
        keyinput34, keyinput33, keyinput32, keyinput31, keyinput30, keyinput29, 
        keyinput28, keyinput27, keyinput26, keyinput25, keyinput24, keyinput23, 
        keyinput22, keyinput21, keyinput20, keyinput19, keyinput18, keyinput17, 
        keyinput16, keyinput15, keyinput14, keyinput13, keyinput12, keyinput11, 
        keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, keyinput5, 
        keyinput4, keyinput3, keyinput2, keyinput1, keyinput0 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput63, keyinput62, keyinput61, keyinput60,
         keyinput59, keyinput58, keyinput57, keyinput56, keyinput55,
         keyinput54, keyinput53, keyinput52, keyinput51, keyinput50,
         keyinput49, keyinput48, keyinput47, keyinput46, keyinput45,
         keyinput44, keyinput43, keyinput42, keyinput41, keyinput40,
         keyinput39, keyinput38, keyinput37, keyinput36, keyinput35,
         keyinput34, keyinput33, keyinput32, keyinput31, keyinput30,
         keyinput29, keyinput28, keyinput27, keyinput26, keyinput25,
         keyinput24, keyinput23, keyinput22, keyinput21, keyinput20,
         keyinput19, keyinput18, keyinput17, keyinput16, keyinput15,
         keyinput14, keyinput13, keyinput12, keyinput11, keyinput10, keyinput9,
         keyinput8, keyinput7, keyinput6, keyinput5, keyinput4, keyinput3,
         keyinput2, keyinput1, keyinput0;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903,
         n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913,
         n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923,
         n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933,
         n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943,
         n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953,
         n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963,
         n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973,
         n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983,
         n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993,
         n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003,
         n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013,
         n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023,
         n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033,
         n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043,
         n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053,
         n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063,
         n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073,
         n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083,
         n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093,
         n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103,
         n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113,
         n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123,
         n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133,
         n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143,
         n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153,
         n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163,
         n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173,
         n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183,
         n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193,
         n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203,
         n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213,
         n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223,
         n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233,
         n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243,
         n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253,
         n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263,
         n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273,
         n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283,
         n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293,
         n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303,
         n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313,
         n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323,
         n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333,
         n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
         n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353,
         n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363,
         n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373,
         n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383,
         n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393,
         n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403,
         n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413,
         n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423,
         n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433,
         n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443,
         n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453,
         n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463,
         n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473,
         n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483,
         n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493,
         n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503,
         n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513,
         n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523,
         n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533,
         n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543,
         n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553,
         n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563,
         n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
         n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
         n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593,
         n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
         n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
         n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
         n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
         n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
         n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
         n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
         n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
         n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
         n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
         n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
         n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713,
         n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723,
         n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733,
         n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743,
         n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753,
         n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763,
         n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773,
         n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783,
         n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793,
         n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803,
         n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813,
         n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823,
         n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833,
         n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843,
         n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853,
         n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863,
         n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873,
         n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883,
         n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893,
         n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903,
         n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913,
         n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923,
         n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933,
         n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943,
         n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953,
         n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963,
         n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973,
         n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983,
         n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993,
         n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003,
         n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013,
         n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023,
         n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033,
         n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043,
         n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053,
         n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063,
         n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073,
         n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083,
         n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093,
         n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103,
         n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113,
         n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123,
         n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133,
         n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143,
         n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153,
         n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163,
         n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173,
         n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183,
         n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193,
         n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203,
         n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213,
         n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223,
         n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233,
         n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243,
         n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253,
         n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263,
         n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273,
         n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283,
         n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293,
         n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303,
         n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
         n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
         n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333,
         n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
         n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353,
         n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
         n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373,
         n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383,
         n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
         n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403,
         n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413,
         n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423,
         n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433,
         n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443,
         n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453,
         n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
         n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473,
         n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
         n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
         n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
         n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588;

  CLKBUF_X2 U2245 ( .A(n2022), .Z(n3610) );
  INV_X1 U2246 ( .A(n3487), .ZN(n2789) );
  NAND4_X1 U2247 ( .A1(n2281), .A2(n2280), .A3(n2279), .A4(n2278), .ZN(n2879)
         );
  NAND4_X2 U2248 ( .A1(n2025), .A2(n2277), .A3(n2067), .A4(n2066), .ZN(n3763)
         );
  AND2_X1 U2249 ( .A1(n2630), .A2(n2627), .ZN(n2282) );
  NOR4_X1 U2250 ( .A1(n3619), .A2(n3618), .A3(n3617), .A4(n3616), .ZN(n3624)
         );
  NOR4_X1 U2251 ( .A1(n3850), .A2(n3632), .A3(n3631), .A4(n3630), .ZN(n3633)
         );
  INV_X1 U2252 ( .A(n2007), .ZN(n2862) );
  INV_X1 U2253 ( .A(n3425), .ZN(n2860) );
  OR2_X1 U2254 ( .A1(n3835), .A2(n2520), .ZN(n3439) );
  NAND2_X1 U2255 ( .A1(n2191), .A2(n2193), .ZN(n3861) );
  NAND2_X1 U2256 ( .A1(n2576), .A2(n3643), .ZN(n2728) );
  XNOR2_X1 U2257 ( .A(n2258), .B(n2257), .ZN(n2260) );
  CLKBUF_X2 U2259 ( .A(n2283), .Z(n2008) );
  AND4_X1 U2260 ( .A1(n2287), .A2(n2288), .A3(n2285), .A4(n2286), .ZN(n3487)
         );
  NAND2_X1 U2261 ( .A1(n4047), .A2(n2222), .ZN(n4030) );
  OAI21_X1 U2262 ( .B1(n3874), .B2(n2525), .A(n2509), .ZN(n3883) );
  INV_X2 U2263 ( .A(IR_REG_31__SCAN_IN), .ZN(n2457) );
  NAND2_X1 U2264 ( .A1(n2727), .A2(n2726), .ZN(n2003) );
  OAI21_X2 U2265 ( .B1(n3439), .B2(n2525), .A(n2524), .ZN(n3423) );
  AND2_X2 U2266 ( .A1(n2272), .A2(n2236), .ZN(n2247) );
  NOR2_X2 U2267 ( .A1(n2315), .A2(n2235), .ZN(n2272) );
  OAI22_X2 U2268 ( .A1(n3811), .A2(n3810), .B1(n3809), .B2(
        REG2_REG_13__SCAN_IN), .ZN(n3812) );
  XNOR2_X2 U2269 ( .A(n2289), .B(IR_REG_2__SCAN_IN), .ZN(n4338) );
  INV_X1 U2270 ( .A(n3760), .ZN(n3486) );
  INV_X1 U2271 ( .A(n2008), .ZN(n2004) );
  AND2_X1 U2272 ( .A1(n2829), .A2(n4559), .ZN(n2005) );
  AND2_X1 U2273 ( .A1(n2829), .A2(n4559), .ZN(n3353) );
  AND2_X1 U2274 ( .A1(n2120), .A2(n2119), .ZN(n4441) );
  NAND4_X1 U2275 ( .A1(n2306), .A2(n2305), .A3(n2304), .A4(n2303), .ZN(n3760)
         );
  CLKBUF_X2 U2276 ( .A(n2282), .Z(n2006) );
  XNOR2_X1 U2277 ( .A(n2253), .B(n3449), .ZN(n2259) );
  NOR3_X1 U2278 ( .A1(IR_REG_16__SCAN_IN), .A2(IR_REG_14__SCAN_IN), .A3(
        IR_REG_15__SCAN_IN), .ZN(n2246) );
  NOR2_X1 U2279 ( .A1(n4085), .A2(n2089), .ZN(n2088) );
  OAI21_X1 U2280 ( .B1(n2620), .B2(n4586), .A(n2077), .ZN(n2618) );
  MUX2_X1 U2281 ( .A(REG0_REG_28__SCAN_IN), .B(n2620), .S(n4577), .Z(n2621) );
  AND2_X1 U2282 ( .A1(n2149), .A2(n2145), .ZN(n3574) );
  OAI21_X1 U2283 ( .B1(n3510), .B2(n3503), .A(n3504), .ZN(n3553) );
  NAND2_X1 U2284 ( .A1(n3543), .A2(n3546), .ZN(n3510) );
  AOI211_X1 U2285 ( .C1(n4091), .C2(n4561), .A(n4090), .B(n4089), .ZN(n4298)
         );
  NAND2_X1 U2286 ( .A1(n2139), .A2(n2136), .ZN(n3341) );
  NAND2_X1 U2287 ( .A1(n3112), .A2(n3111), .ZN(n3178) );
  NAND2_X1 U2288 ( .A1(n3028), .A2(n3027), .ZN(n2168) );
  OR2_X1 U2289 ( .A1(n2839), .A2(n2135), .ZN(n2134) );
  OR2_X1 U2290 ( .A1(n2495), .A2(n4096), .ZN(n2504) );
  INV_X1 U2291 ( .A(n2829), .ZN(n3427) );
  NAND2_X2 U2292 ( .A1(n2782), .A2(n2728), .ZN(n3425) );
  NAND4_X1 U2293 ( .A1(n2295), .A2(n2294), .A3(n2293), .A4(n2292), .ZN(n3761)
         );
  NAND3_X2 U2294 ( .A1(n2594), .A2(n2641), .A3(n2593), .ZN(n2727) );
  INV_X1 U2295 ( .A(n2597), .ZN(n3643) );
  INV_X1 U2296 ( .A(n2259), .ZN(n2630) );
  OR2_X1 U2297 ( .A1(n2580), .A2(n2457), .ZN(n2581) );
  AND2_X1 U2298 ( .A1(n2461), .A2(n2526), .ZN(n4334) );
  AND2_X1 U2299 ( .A1(n2531), .A2(n2579), .ZN(n2580) );
  XNOR2_X1 U2300 ( .A(n2530), .B(n2240), .ZN(n2597) );
  NAND3_X2 U2301 ( .A1(n2087), .A2(n2086), .A3(n2245), .ZN(n2462) );
  NAND2_X1 U2302 ( .A1(n3448), .A2(IR_REG_31__SCAN_IN), .ZN(n2253) );
  AND2_X1 U2303 ( .A1(n2255), .A2(n2200), .ZN(n2258) );
  AND3_X1 U2304 ( .A1(n2243), .A2(n2015), .A3(n2228), .ZN(n2244) );
  NOR2_X1 U2305 ( .A1(n2241), .A2(n2582), .ZN(n2579) );
  NAND3_X2 U2306 ( .A1(n2100), .A2(n2099), .A3(n2098), .ZN(n4339) );
  NAND2_X1 U2307 ( .A1(n2457), .A2(IR_REG_1__SCAN_IN), .ZN(n2098) );
  AND2_X1 U2308 ( .A1(n2246), .A2(n2242), .ZN(n2174) );
  NOR2_X1 U2309 ( .A1(IR_REG_18__SCAN_IN), .A2(n2029), .ZN(n2015) );
  NOR2_X1 U2310 ( .A1(IR_REG_12__SCAN_IN), .A2(IR_REG_10__SCAN_IN), .ZN(n2234)
         );
  NOR2_X1 U2311 ( .A1(IR_REG_9__SCAN_IN), .A2(IR_REG_8__SCAN_IN), .ZN(n2232)
         );
  NOR2_X1 U2312 ( .A1(IR_REG_5__SCAN_IN), .A2(IR_REG_7__SCAN_IN), .ZN(n2233)
         );
  INV_X1 U2313 ( .A(IR_REG_24__SCAN_IN), .ZN(n2585) );
  INV_X1 U2314 ( .A(IR_REG_23__SCAN_IN), .ZN(n2596) );
  NOR2_X1 U2315 ( .A1(IR_REG_11__SCAN_IN), .A2(IR_REG_6__SCAN_IN), .ZN(n2231)
         );
  INV_X1 U2316 ( .A(IR_REG_3__SCAN_IN), .ZN(n2297) );
  INV_X1 U2317 ( .A(IR_REG_2__SCAN_IN), .ZN(n4169) );
  NAND2_X1 U2318 ( .A1(n4427), .A2(REG2_REG_12__SCAN_IN), .ZN(n4426) );
  NAND2_X1 U2319 ( .A1(n2260), .A2(n2630), .ZN(n2283) );
  INV_X1 U2320 ( .A(n2260), .ZN(n2627) );
  AOI21_X2 U2321 ( .B1(n3958), .B2(n2479), .A(n2478), .ZN(n3941) );
  OAI21_X2 U2322 ( .B1(n3051), .B2(n2212), .A(n2210), .ZN(n3128) );
  NAND2_X2 U2323 ( .A1(n2354), .A2(n2353), .ZN(n3051) );
  AND2_X4 U2325 ( .A1(n2728), .A2(n2727), .ZN(n2829) );
  NAND2_X1 U2326 ( .A1(n2918), .A2(n2300), .ZN(n2203) );
  NAND2_X1 U2327 ( .A1(n3487), .A2(n3459), .ZN(n3644) );
  OR2_X1 U2328 ( .A1(n2042), .A2(n2017), .ZN(n2167) );
  AOI21_X1 U2329 ( .B1(REG1_REG_11__SCAN_IN), .B2(n3235), .A(n4411), .ZN(n3236) );
  AND2_X1 U2330 ( .A1(n3575), .A2(n3855), .ZN(n3732) );
  OR2_X1 U2331 ( .A1(n3895), .A2(n3695), .ZN(n2071) );
  INV_X1 U2332 ( .A(n2218), .ZN(n2211) );
  AND2_X1 U2333 ( .A1(n2579), .A2(n4201), .ZN(n2243) );
  INV_X1 U2334 ( .A(n4016), .ZN(n3565) );
  OR2_X1 U2335 ( .A1(n2255), .A2(IR_REG_27__SCAN_IN), .ZN(n2087) );
  NAND2_X1 U2336 ( .A1(n2255), .A2(IR_REG_28__SCAN_IN), .ZN(n2086) );
  NOR2_X1 U2337 ( .A1(n2536), .A2(n4334), .ZN(n2781) );
  INV_X1 U2338 ( .A(n2006), .ZN(n2525) );
  OR2_X1 U2339 ( .A1(n4421), .A2(n4422), .ZN(n2104) );
  INV_X1 U2340 ( .A(n2194), .ZN(n2193) );
  OAI21_X1 U2341 ( .B1(n2196), .B2(n2195), .A(n2503), .ZN(n2194) );
  AND2_X1 U2342 ( .A1(n2615), .A2(n3836), .ZN(n3841) );
  AND2_X1 U2343 ( .A1(n2535), .A2(n2536), .ZN(n4554) );
  AND2_X1 U2344 ( .A1(n2449), .A2(n2448), .ZN(n4483) );
  OAI21_X1 U2345 ( .B1(n4339), .B2(n2663), .A(n2101), .ZN(n3764) );
  NAND2_X1 U2346 ( .A1(n4339), .A2(n2663), .ZN(n2101) );
  OR2_X1 U2347 ( .A1(n3472), .A2(n3473), .ZN(n2159) );
  NOR2_X1 U2348 ( .A1(n3693), .A2(n3694), .ZN(n2070) );
  AND2_X1 U2349 ( .A1(n2076), .A2(n3637), .ZN(n2075) );
  AND2_X1 U2350 ( .A1(n2367), .A2(n2034), .ZN(n2218) );
  NOR2_X1 U2351 ( .A1(n3628), .A2(n2214), .ZN(n2213) );
  INV_X1 U2352 ( .A(n2216), .ZN(n2214) );
  AOI21_X1 U2353 ( .B1(n2024), .B2(n2218), .A(n2217), .ZN(n2216) );
  NOR2_X1 U2354 ( .A1(n3181), .A2(n3142), .ZN(n2217) );
  OAI21_X1 U2355 ( .B1(n3052), .B2(n3663), .A(n3661), .ZN(n3139) );
  INV_X1 U2356 ( .A(n3667), .ZN(n2057) );
  INV_X1 U2357 ( .A(n3653), .ZN(n2063) );
  AOI21_X1 U2358 ( .B1(n2062), .B2(n2549), .A(n2060), .ZN(n2059) );
  INV_X1 U2359 ( .A(n3665), .ZN(n2060) );
  AND2_X1 U2360 ( .A1(n2546), .A2(n2761), .ZN(n2290) );
  NAND2_X1 U2361 ( .A1(n3629), .A2(n2084), .ZN(n2878) );
  INV_X1 U2362 ( .A(IR_REG_26__SCAN_IN), .ZN(n4201) );
  NOR2_X1 U2363 ( .A1(n3130), .A2(n3326), .ZN(n2093) );
  AND2_X1 U2364 ( .A1(n2019), .A2(n3053), .ZN(n2092) );
  NAND2_X1 U2365 ( .A1(n2188), .A2(n2187), .ZN(n2186) );
  NAND2_X1 U2366 ( .A1(n2320), .A2(n2189), .ZN(n2185) );
  NOR2_X1 U2367 ( .A1(n2190), .A2(n2329), .ZN(n2189) );
  INV_X1 U2368 ( .A(n2319), .ZN(n2190) );
  NAND2_X1 U2369 ( .A1(n2247), .A2(n2174), .ZN(n2447) );
  INV_X1 U2370 ( .A(IR_REG_6__SCAN_IN), .ZN(n2336) );
  NAND2_X1 U2371 ( .A1(n2141), .A2(n2143), .ZN(n2138) );
  NOR2_X1 U2372 ( .A1(n2142), .A2(n3278), .ZN(n2140) );
  INV_X1 U2373 ( .A(n3188), .ZN(n2143) );
  NAND2_X1 U2374 ( .A1(n2167), .A2(n2041), .ZN(n2163) );
  NAND2_X1 U2375 ( .A1(n2158), .A2(n2038), .ZN(n2155) );
  XNOR2_X1 U2376 ( .A(n2832), .B(n3425), .ZN(n2836) );
  NOR2_X1 U2377 ( .A1(n3096), .A2(n2170), .ZN(n2169) );
  INV_X1 U2378 ( .A(n2172), .ZN(n2170) );
  NAND2_X1 U2379 ( .A1(n3093), .A2(n2173), .ZN(n2171) );
  OR2_X1 U2380 ( .A1(n3091), .A2(n3092), .ZN(n2173) );
  AOI22_X1 U2381 ( .A1(n3763), .A2(n2005), .B1(n2007), .B2(n2790), .ZN(n2816)
         );
  XNOR2_X1 U2382 ( .A(n2788), .B(n3425), .ZN(n2818) );
  XNOR2_X1 U2383 ( .A(n2823), .B(n2860), .ZN(n2824) );
  NAND2_X1 U2384 ( .A1(n2822), .A2(n2821), .ZN(n2823) );
  NOR2_X1 U2385 ( .A1(n2167), .A2(n2165), .ZN(n2164) );
  AND2_X1 U2386 ( .A1(n4356), .A2(n2166), .ZN(n2165) );
  NAND2_X1 U2387 ( .A1(n2157), .A2(n2018), .ZN(n2152) );
  INV_X1 U2388 ( .A(n3517), .ZN(n2147) );
  NAND2_X1 U2389 ( .A1(n2151), .A2(n3516), .ZN(n2150) );
  INV_X1 U2390 ( .A(n2153), .ZN(n2151) );
  NAND2_X1 U2391 ( .A1(n2807), .A2(REG1_REG_8__SCAN_IN), .ZN(n2109) );
  AOI21_X1 U2392 ( .B1(REG1_REG_9__SCAN_IN), .B2(n4335), .A(n3232), .ZN(n3233)
         );
  NAND2_X1 U2393 ( .A1(n2104), .A2(n2028), .ZN(n2103) );
  NAND2_X1 U2394 ( .A1(n2103), .A2(n2102), .ZN(n3797) );
  INV_X1 U2395 ( .A(n3239), .ZN(n2102) );
  AND2_X1 U2396 ( .A1(n3797), .A2(n3796), .ZN(n3799) );
  OR2_X1 U2397 ( .A1(n4431), .A2(n4432), .ZN(n2117) );
  INV_X1 U2398 ( .A(n4442), .ZN(n2119) );
  NOR2_X1 U2399 ( .A1(n4446), .A2(n3802), .ZN(n3803) );
  AND2_X1 U2400 ( .A1(n3814), .A2(REG1_REG_15__SCAN_IN), .ZN(n3802) );
  NAND2_X1 U2401 ( .A1(n3841), .A2(n4083), .ZN(n4078) );
  OAI21_X1 U2402 ( .B1(n3849), .B2(n3850), .A(n2575), .ZN(n3829) );
  INV_X1 U2403 ( .A(n3423), .ZN(n3853) );
  NAND2_X1 U2404 ( .A1(n2033), .A2(n2010), .ZN(n2196) );
  NOR2_X2 U2405 ( .A1(n2480), .A2(n4196), .ZN(n2485) );
  AND2_X1 U2406 ( .A1(n3974), .A2(n3963), .ZN(n2478) );
  AOI21_X1 U2407 ( .B1(n2181), .B2(n2179), .A(n2030), .ZN(n2178) );
  INV_X1 U2408 ( .A(n2438), .ZN(n2179) );
  INV_X1 U2409 ( .A(n2181), .ZN(n2180) );
  INV_X1 U2410 ( .A(n3966), .ZN(n3995) );
  AND2_X1 U2411 ( .A1(n4014), .A2(n2043), .ZN(n2181) );
  NAND2_X1 U2412 ( .A1(n4030), .A2(n2438), .ZN(n2182) );
  OAI21_X1 U2413 ( .B1(n2561), .B2(n2074), .A(n2072), .ZN(n4058) );
  INV_X1 U2414 ( .A(n2073), .ZN(n2072) );
  OAI21_X1 U2415 ( .B1(n2075), .B2(n2074), .A(n4059), .ZN(n2073) );
  INV_X1 U2416 ( .A(n3635), .ZN(n2074) );
  NAND2_X1 U2417 ( .A1(n2561), .A2(n2075), .ZN(n3309) );
  NOR2_X1 U2418 ( .A1(n3302), .A2(n4278), .ZN(n4050) );
  NAND2_X1 U2419 ( .A1(n2400), .A2(n2208), .ZN(n2206) );
  AND2_X1 U2420 ( .A1(n2399), .A2(n2209), .ZN(n2208) );
  NAND2_X1 U2421 ( .A1(n2401), .A2(n3267), .ZN(n2209) );
  OR2_X1 U2422 ( .A1(n2957), .A2(n3658), .ZN(n2552) );
  INV_X1 U2423 ( .A(n4064), .ZN(n3994) );
  AND2_X1 U2424 ( .A1(n2577), .A2(n3738), .ZN(n3998) );
  INV_X1 U2425 ( .A(n4018), .ZN(n4061) );
  NAND2_X1 U2426 ( .A1(n2727), .A2(n4518), .ZN(n2753) );
  OR2_X1 U2427 ( .A1(n4341), .A2(n2742), .ZN(n4018) );
  INV_X1 U2428 ( .A(n3998), .ZN(n4057) );
  INV_X1 U2429 ( .A(n2790), .ZN(n2882) );
  INV_X1 U2430 ( .A(n2543), .ZN(n3629) );
  NAND2_X1 U2431 ( .A1(n4078), .A2(n2090), .ZN(n4084) );
  OR2_X1 U2432 ( .A1(n4083), .A2(n3841), .ZN(n2090) );
  NAND2_X1 U2433 ( .A1(n4050), .A2(n4348), .ZN(n4051) );
  NAND2_X1 U2434 ( .A1(n4038), .A2(n4021), .ZN(n2085) );
  NOR3_X1 U2435 ( .A1(n4051), .A2(n2085), .A3(n3607), .ZN(n4000) );
  AND2_X1 U2436 ( .A1(n3163), .A2(n3162), .ZN(n3160) );
  OR2_X1 U2437 ( .A1(n3006), .A2(n2617), .ZN(n4559) );
  INV_X1 U2438 ( .A(n2753), .ZN(n2873) );
  NOR2_X1 U2439 ( .A1(n2201), .A2(n2256), .ZN(n2200) );
  AND2_X1 U2440 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_28__SCAN_IN), .ZN(n2256)
         );
  INV_X1 U2441 ( .A(IR_REG_28__SCAN_IN), .ZN(n2538) );
  INV_X1 U2442 ( .A(IR_REG_25__SCAN_IN), .ZN(n2238) );
  NAND2_X1 U2443 ( .A1(n2532), .A2(IR_REG_31__SCAN_IN), .ZN(n2533) );
  OR2_X1 U2444 ( .A1(n2458), .A2(n2457), .ZN(n2459) );
  NAND2_X1 U2445 ( .A1(n2459), .A2(n2460), .ZN(n2526) );
  NOR2_X1 U2446 ( .A1(n2365), .A2(IR_REG_9__SCAN_IN), .ZN(n2384) );
  AND2_X1 U2447 ( .A1(n2504), .A2(n2496), .ZN(n3889) );
  INV_X1 U2448 ( .A(n3000), .ZN(n2993) );
  INV_X1 U2449 ( .A(n3283), .ZN(n3587) );
  INV_X1 U2450 ( .A(n4034), .ZN(n3586) );
  OR2_X1 U2451 ( .A1(n3934), .A2(n2525), .ZN(n2488) );
  NAND4_X1 U2452 ( .A1(n2456), .A2(n2455), .A3(n2454), .A4(n2453), .ZN(n4016)
         );
  NAND4_X1 U2453 ( .A1(n2410), .A2(n2409), .A3(n2408), .A4(n2407), .ZN(n4062)
         );
  NAND2_X1 U2454 ( .A1(n2022), .A2(REG1_REG_0__SCAN_IN), .ZN(n2281) );
  NAND2_X1 U2455 ( .A1(n2665), .A2(n2664), .ZN(n3790) );
  XNOR2_X1 U2456 ( .A(n3799), .B(n3798), .ZN(n4431) );
  NAND2_X1 U2457 ( .A1(n4467), .A2(n4468), .ZN(n4466) );
  NAND2_X1 U2458 ( .A1(n4466), .A2(n2107), .ZN(n4478) );
  OR2_X1 U2459 ( .A1(n3817), .A2(REG1_REG_17__SCAN_IN), .ZN(n2107) );
  INV_X1 U2460 ( .A(n4480), .ZN(n2129) );
  AOI21_X1 U2461 ( .B1(n4481), .B2(n4482), .A(n4479), .ZN(n2128) );
  OAI211_X1 U2462 ( .C1(n4488), .C2(n4489), .A(n4487), .B(n2054), .ZN(n2127)
         );
  INV_X1 U2463 ( .A(n4470), .ZN(n4476) );
  INV_X1 U2464 ( .A(n4272), .ZN(n4348) );
  NAND2_X1 U2465 ( .A1(n2081), .A2(n2078), .ZN(n2620) );
  INV_X1 U2466 ( .A(n3445), .ZN(n2081) );
  INV_X1 U2467 ( .A(n2079), .ZN(n2078) );
  OAI21_X1 U2468 ( .B1(n3447), .B2(n4569), .A(n2080), .ZN(n2079) );
  OR2_X1 U2469 ( .A1(n3841), .A2(n2616), .ZN(n3443) );
  NOR2_X1 U2470 ( .A1(n4441), .A2(n2118), .ZN(n3815) );
  AND2_X1 U2471 ( .A1(n3814), .A2(REG2_REG_15__SCAN_IN), .ZN(n2118) );
  AND2_X1 U2472 ( .A1(n2502), .A2(n2013), .ZN(n2192) );
  NAND2_X1 U2473 ( .A1(n3650), .A2(n3653), .ZN(n2933) );
  INV_X1 U2474 ( .A(n2254), .ZN(n2201) );
  NAND2_X1 U2475 ( .A1(n2240), .A2(n2239), .ZN(n2582) );
  INV_X1 U2476 ( .A(IR_REG_4__SCAN_IN), .ZN(n2229) );
  NOR2_X1 U2477 ( .A1(n2219), .A2(n2729), .ZN(n2783) );
  NAND2_X1 U2478 ( .A1(n2154), .A2(n2018), .ZN(n2153) );
  INV_X1 U2479 ( .A(n2159), .ZN(n2154) );
  NAND2_X1 U2480 ( .A1(n3091), .A2(n3092), .ZN(n2172) );
  INV_X1 U2481 ( .A(REG3_REG_9__SCAN_IN), .ZN(n2355) );
  NAND2_X1 U2482 ( .A1(n3377), .A2(n3376), .ZN(n3378) );
  INV_X1 U2483 ( .A(n3374), .ZN(n3377) );
  INV_X1 U2484 ( .A(n3375), .ZN(n3376) );
  NAND2_X1 U2485 ( .A1(n2463), .A2(REG3_REG_20__SCAN_IN), .ZN(n2471) );
  OR2_X1 U2486 ( .A1(n2471), .A2(n3511), .ZN(n2480) );
  OR2_X1 U2487 ( .A1(n2428), .A2(n4181), .ZN(n2439) );
  NOR2_X1 U2488 ( .A1(n2321), .A2(n2912), .ZN(n2330) );
  NOR2_X1 U2489 ( .A1(n2404), .A2(n2403), .ZN(n2415) );
  NAND2_X1 U2490 ( .A1(n2122), .A2(n2121), .ZN(n2682) );
  AOI21_X1 U2491 ( .B1(n2124), .B2(n2125), .A(n2709), .ZN(n2121) );
  INV_X1 U2492 ( .A(REG3_REG_13__SCAN_IN), .ZN(n3231) );
  NAND2_X1 U2493 ( .A1(n4415), .A2(n3225), .ZN(n3227) );
  XNOR2_X1 U2494 ( .A(n3815), .B(n2427), .ZN(n4453) );
  NOR2_X1 U2495 ( .A1(n4078), .A2(n4080), .ZN(n4077) );
  AND2_X1 U2496 ( .A1(n3699), .A2(n3828), .ZN(n3837) );
  AND2_X1 U2497 ( .A1(n2516), .A2(n2515), .ZN(n3575) );
  AND2_X1 U2498 ( .A1(n2462), .A2(DATAI_27_), .ZN(n3855) );
  OAI21_X1 U2499 ( .B1(n2071), .B2(n2574), .A(n2068), .ZN(n3849) );
  NOR2_X1 U2500 ( .A1(n2069), .A2(n2027), .ZN(n2068) );
  NOR2_X1 U2501 ( .A1(n2574), .A2(n2070), .ZN(n2069) );
  NAND2_X1 U2502 ( .A1(n2071), .A2(n3603), .ZN(n3881) );
  NAND2_X1 U2503 ( .A1(n2485), .A2(REG3_REG_23__SCAN_IN), .ZN(n2491) );
  OR2_X1 U2504 ( .A1(n2009), .A2(n4250), .ZN(n3959) );
  OR2_X1 U2505 ( .A1(n4033), .A2(n3916), .ZN(n3918) );
  AND4_X1 U2506 ( .A1(n2477), .A2(n2476), .A3(n2475), .A4(n2474), .ZN(n3974)
         );
  AOI21_X2 U2507 ( .B1(n2175), .B2(n2177), .A(n2176), .ZN(n3978) );
  NOR2_X1 U2508 ( .A1(n2180), .A2(n2011), .ZN(n2177) );
  OAI21_X1 U2509 ( .B1(n2178), .B2(n2011), .A(n2032), .ZN(n2176) );
  INV_X1 U2510 ( .A(n4063), .ZN(n4345) );
  NAND2_X1 U2511 ( .A1(n4058), .A2(n3683), .ZN(n4033) );
  NOR2_X1 U2512 ( .A1(n2207), .A2(n2205), .ZN(n2204) );
  INV_X1 U2513 ( .A(n3754), .ZN(n3323) );
  AOI21_X1 U2514 ( .B1(n2213), .B2(n2211), .A(n2031), .ZN(n2210) );
  INV_X1 U2515 ( .A(n2213), .ZN(n2212) );
  INV_X1 U2516 ( .A(REG3_REG_12__SCAN_IN), .ZN(n2386) );
  NAND2_X1 U2517 ( .A1(n2554), .A2(n3671), .ZN(n3152) );
  NAND2_X1 U2518 ( .A1(n2215), .A2(n2216), .ZN(n3153) );
  NAND2_X1 U2519 ( .A1(n3051), .A2(n2218), .ZN(n2215) );
  AND2_X1 U2520 ( .A1(n2368), .A2(REG3_REG_10__SCAN_IN), .ZN(n2376) );
  INV_X1 U2521 ( .A(n3154), .ZN(n3181) );
  NAND2_X1 U2522 ( .A1(n2082), .A2(n3668), .ZN(n3052) );
  NAND2_X1 U2523 ( .A1(n3076), .A2(n3660), .ZN(n2082) );
  INV_X1 U2524 ( .A(REG3_REG_8__SCAN_IN), .ZN(n2342) );
  INV_X1 U2525 ( .A(n3757), .ZN(n3097) );
  OAI21_X1 U2526 ( .B1(n2934), .B2(n2058), .A(n2056), .ZN(n2550) );
  AOI21_X1 U2527 ( .B1(n2059), .B2(n2061), .A(n2057), .ZN(n2056) );
  INV_X1 U2528 ( .A(n2059), .ZN(n2058) );
  NAND2_X1 U2529 ( .A1(n2055), .A2(n2059), .ZN(n2973) );
  NAND2_X1 U2530 ( .A1(n2934), .A2(n2062), .ZN(n2055) );
  NAND2_X1 U2531 ( .A1(n2064), .A2(n3653), .ZN(n2992) );
  NAND2_X1 U2532 ( .A1(n2065), .A2(n3650), .ZN(n2064) );
  INV_X1 U2533 ( .A(n2934), .ZN(n2065) );
  INV_X1 U2534 ( .A(n2938), .ZN(n2931) );
  NAND2_X1 U2535 ( .A1(n2932), .A2(n2931), .ZN(n2998) );
  AND2_X1 U2536 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n2310) );
  INV_X1 U2537 ( .A(n2933), .ZN(n3597) );
  AND3_X1 U2538 ( .A1(n2882), .A2(n3015), .A3(n2091), .ZN(n2932) );
  NOR2_X1 U2539 ( .A1(n3459), .A2(n2926), .ZN(n2091) );
  NAND2_X1 U2540 ( .A1(n2543), .A2(n3640), .ZN(n2877) );
  NAND2_X1 U2541 ( .A1(n4277), .A2(n3441), .ZN(n2080) );
  AND2_X1 U2542 ( .A1(n3870), .A2(n4087), .ZN(n2615) );
  NOR2_X1 U2543 ( .A1(n3887), .A2(n2614), .ZN(n3870) );
  NOR3_X1 U2544 ( .A1(n3959), .A2(n3605), .A3(n3953), .ZN(n3931) );
  AND2_X1 U2545 ( .A1(n2462), .A2(DATAI_21_), .ZN(n4250) );
  NAND2_X1 U2546 ( .A1(n3160), .A2(n2020), .ZN(n3302) );
  NAND2_X1 U2547 ( .A1(n3160), .A2(n2093), .ZN(n3247) );
  NAND2_X1 U2548 ( .A1(n3160), .A2(n3257), .ZN(n3214) );
  INV_X1 U2549 ( .A(n3183), .ZN(n3162) );
  AND2_X1 U2550 ( .A1(n2981), .A2(n2045), .ZN(n3163) );
  NAND2_X1 U2551 ( .A1(n2981), .A2(n2019), .ZN(n3073) );
  AND2_X1 U2552 ( .A1(n2981), .A2(n3064), .ZN(n3074) );
  INV_X1 U2553 ( .A(n4561), .ZN(n4569) );
  NOR2_X1 U2554 ( .A1(n3627), .A2(n2184), .ZN(n2183) );
  INV_X1 U2555 ( .A(n2186), .ZN(n2184) );
  NAND2_X1 U2556 ( .A1(n2185), .A2(n2186), .ZN(n2964) );
  OR2_X1 U2557 ( .A1(n2998), .A2(n2993), .ZN(n2999) );
  NOR2_X1 U2558 ( .A1(n2999), .A2(n2979), .ZN(n2981) );
  NAND2_X1 U2559 ( .A1(n3212), .A2(n4545), .ZN(n4561) );
  NAND2_X1 U2560 ( .A1(n2882), .A2(n3015), .ZN(n2876) );
  INV_X1 U2561 ( .A(n4554), .ZN(n4545) );
  NAND2_X1 U2562 ( .A1(n2593), .A2(n2590), .ZN(n2646) );
  NAND2_X1 U2563 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_27__SCAN_IN), .ZN(n2254) );
  AND2_X1 U2564 ( .A1(n2246), .A2(n2242), .ZN(n2228) );
  XNOR2_X1 U2565 ( .A(n2528), .B(n2527), .ZN(n2576) );
  INV_X1 U2566 ( .A(IR_REG_20__SCAN_IN), .ZN(n2527) );
  NAND2_X1 U2567 ( .A1(n2526), .A2(IR_REG_31__SCAN_IN), .ZN(n2528) );
  XNOR2_X1 U2568 ( .A(n2396), .B(IR_REG_11__SCAN_IN), .ZN(n3235) );
  INV_X1 U2569 ( .A(IR_REG_7__SCAN_IN), .ZN(n2338) );
  INV_X1 U2570 ( .A(IR_REG_5__SCAN_IN), .ZN(n4162) );
  NAND2_X1 U2571 ( .A1(n2168), .A2(n3029), .ZN(n3067) );
  INV_X1 U2572 ( .A(n3033), .ZN(n3064) );
  INV_X1 U2573 ( .A(n2137), .ZN(n2136) );
  NAND2_X1 U2574 ( .A1(n3178), .A2(n2140), .ZN(n2139) );
  OAI21_X1 U2575 ( .B1(n3278), .B2(n2138), .A(n3277), .ZN(n2137) );
  INV_X1 U2576 ( .A(n3755), .ZN(n3115) );
  NAND2_X1 U2577 ( .A1(n3065), .A2(n3039), .ZN(n3093) );
  NAND2_X1 U2578 ( .A1(n2144), .A2(n2152), .ZN(n3519) );
  OR2_X1 U2579 ( .A1(n3471), .A2(n2153), .ZN(n2144) );
  NAND2_X1 U2580 ( .A1(n2857), .A2(n2856), .ZN(n2895) );
  OAI21_X1 U2581 ( .B1(n3352), .B2(n2164), .A(n2163), .ZN(n3528) );
  NAND2_X1 U2582 ( .A1(n2155), .A2(n3404), .ZN(n3534) );
  NAND2_X1 U2583 ( .A1(n2840), .A2(n2839), .ZN(n2857) );
  NAND2_X1 U2584 ( .A1(n2171), .A2(n2172), .ZN(n3095) );
  NAND2_X1 U2585 ( .A1(n3178), .A2(n3177), .ZN(n3189) );
  NAND2_X1 U2586 ( .A1(n2162), .A2(n2160), .ZN(n3564) );
  AOI21_X1 U2587 ( .B1(n2014), .B2(n2164), .A(n2161), .ZN(n2160) );
  NOR2_X1 U2588 ( .A1(n3365), .A2(n3364), .ZN(n2161) );
  AND2_X1 U2589 ( .A1(n2754), .A2(n3950), .ZN(n4349) );
  INV_X1 U2590 ( .A(n2146), .ZN(n2145) );
  OAI21_X1 U2591 ( .B1(n2152), .B2(n2148), .A(n2147), .ZN(n2146) );
  NAND2_X1 U2592 ( .A1(n2791), .A2(n4341), .ZN(n4344) );
  NAND2_X1 U2593 ( .A1(n2791), .A2(n3772), .ZN(n4343) );
  AND2_X1 U2594 ( .A1(n2847), .A2(n2846), .ZN(n4362) );
  INV_X1 U2595 ( .A(n3581), .ZN(n4357) );
  MUX2_X1 U2596 ( .A(n3814), .B(DATAI_15_), .S(n2462), .Z(n4278) );
  INV_X1 U2597 ( .A(n4349), .ZN(n3589) );
  AND2_X1 U2598 ( .A1(n2007), .A2(n2747), .ZN(n3744) );
  INV_X1 U2599 ( .A(n3575), .ZN(n3867) );
  NAND2_X1 U2600 ( .A1(n2501), .A2(n2500), .ZN(n3898) );
  OAI211_X1 U2601 ( .C1(n2008), .C2(n3906), .A(n2494), .B(n2493), .ZN(n3928)
         );
  OR2_X1 U2602 ( .A1(n3905), .A2(n2525), .ZN(n2494) );
  OAI211_X1 U2603 ( .C1(n3951), .C2(n2525), .A(n2484), .B(n2483), .ZN(n3967)
         );
  NAND4_X1 U2604 ( .A1(n2469), .A2(n2468), .A3(n2467), .A4(n2466), .ZN(n3966)
         );
  NAND2_X1 U2605 ( .A1(n2022), .A2(REG1_REG_1__SCAN_IN), .ZN(n2067) );
  OR2_X1 U2606 ( .A1(n2283), .A2(n2276), .ZN(n2066) );
  NAND2_X1 U2607 ( .A1(n3764), .A2(n3765), .ZN(n3787) );
  OR2_X1 U2608 ( .A1(n4372), .A2(n2125), .ZN(n2123) );
  NAND2_X1 U2609 ( .A1(n2023), .A2(n2807), .ZN(n4393) );
  INV_X1 U2610 ( .A(n2109), .ZN(n2108) );
  AND2_X1 U2611 ( .A1(n2109), .A2(n2023), .ZN(n2810) );
  XNOR2_X1 U2612 ( .A(n3233), .B(n4533), .ZN(n4403) );
  NOR2_X1 U2613 ( .A1(n4403), .A2(n4404), .ZN(n4402) );
  NAND2_X1 U2614 ( .A1(n4416), .A2(n4417), .ZN(n4415) );
  OAI21_X1 U2615 ( .B1(n4403), .B2(n2111), .A(n2110), .ZN(n4411) );
  NAND2_X1 U2616 ( .A1(n2112), .A2(REG1_REG_10__SCAN_IN), .ZN(n2111) );
  NAND2_X1 U2617 ( .A1(n3234), .A2(n2112), .ZN(n2110) );
  INV_X1 U2618 ( .A(n4412), .ZN(n2112) );
  XNOR2_X1 U2619 ( .A(n3227), .B(n4529), .ZN(n4427) );
  INV_X1 U2620 ( .A(n2104), .ZN(n4420) );
  INV_X1 U2621 ( .A(n2103), .ZN(n3240) );
  OAI21_X1 U2622 ( .B1(n4431), .B2(n2116), .A(n2114), .ZN(n4446) );
  OR2_X1 U2623 ( .A1(n4447), .A2(n4432), .ZN(n2116) );
  INV_X1 U2624 ( .A(n4447), .ZN(n2115) );
  INV_X1 U2625 ( .A(n3800), .ZN(n2113) );
  INV_X1 U2626 ( .A(n2120), .ZN(n4443) );
  AND2_X1 U2627 ( .A1(n2667), .A2(n3832), .ZN(n4470) );
  AND2_X1 U2628 ( .A1(n2667), .A2(n3745), .ZN(n4472) );
  AND2_X1 U2629 ( .A1(n2106), .A2(n2105), .ZN(n3806) );
  NAND2_X1 U2630 ( .A1(n4483), .A2(REG1_REG_18__SCAN_IN), .ZN(n2105) );
  OR2_X1 U2631 ( .A1(n2505), .A2(n2519), .ZN(n3874) );
  NAND2_X1 U2632 ( .A1(n2197), .A2(n2196), .ZN(n3879) );
  NAND2_X1 U2633 ( .A1(n3914), .A2(n2013), .ZN(n2197) );
  AND2_X1 U2634 ( .A1(n2198), .A2(n2199), .ZN(n3904) );
  NAND2_X1 U2635 ( .A1(n3914), .A2(n2490), .ZN(n2198) );
  OAI21_X1 U2636 ( .B1(n4030), .B2(n2180), .A(n2178), .ZN(n3986) );
  NAND2_X1 U2637 ( .A1(n2182), .A2(n2181), .ZN(n4010) );
  AND2_X1 U2638 ( .A1(n2182), .A2(n2043), .ZN(n4011) );
  NAND2_X1 U2639 ( .A1(n3309), .A2(n3635), .ZN(n4060) );
  NAND2_X1 U2640 ( .A1(n2561), .A2(n3637), .ZN(n3307) );
  NAND2_X1 U2641 ( .A1(n2320), .A2(n2319), .ZN(n2972) );
  OR2_X1 U2642 ( .A1(n2753), .A2(n2752), .ZN(n3950) );
  INV_X1 U2643 ( .A(n4501), .ZN(n4006) );
  NAND2_X1 U2644 ( .A1(n3629), .A2(n2083), .ZN(n2886) );
  INV_X1 U2645 ( .A(n2885), .ZN(n2083) );
  INV_X1 U2646 ( .A(n3950), .ZN(n4497) );
  INV_X1 U2647 ( .A(n2733), .ZN(n3015) );
  INV_X1 U2648 ( .A(n2950), .ZN(n4502) );
  OAI21_X1 U2649 ( .B1(n4084), .B2(n4559), .A(n2088), .ZN(n4296) );
  NAND2_X1 U2650 ( .A1(n4086), .A2(n2053), .ZN(n2089) );
  NOR2_X1 U2651 ( .A1(n4051), .A2(n2085), .ZN(n4003) );
  AND2_X2 U2652 ( .A1(n2874), .A2(n2619), .ZN(n4577) );
  NAND2_X1 U2653 ( .A1(n2873), .A2(n2646), .ZN(n4517) );
  AND2_X1 U2654 ( .A1(n2251), .A2(n2015), .ZN(n2252) );
  AND2_X1 U2655 ( .A1(n2250), .A2(n2249), .ZN(n2251) );
  INV_X1 U2656 ( .A(IR_REG_30__SCAN_IN), .ZN(n3449) );
  INV_X1 U2657 ( .A(n2592), .ZN(n2641) );
  INV_X1 U2658 ( .A(n2536), .ZN(n3747) );
  OR2_X1 U2659 ( .A1(n2459), .A2(n2460), .ZN(n2461) );
  INV_X1 U2660 ( .A(n3817), .ZN(n4522) );
  NOR2_X1 U2661 ( .A1(n2366), .A2(n2384), .ZN(n4335) );
  AND2_X1 U2662 ( .A1(n2307), .A2(n2299), .ZN(n4337) );
  OAI21_X1 U2663 ( .B1(IR_REG_0__SCAN_IN), .B2(IR_REG_1__SCAN_IN), .A(
        IR_REG_31__SCAN_IN), .ZN(n2289) );
  NAND3_X1 U2664 ( .A1(n2131), .A2(IR_REG_0__SCAN_IN), .A3(IR_REG_31__SCAN_IN), 
        .ZN(n2100) );
  NAND2_X1 U2665 ( .A1(n2132), .A2(IR_REG_1__SCAN_IN), .ZN(n2099) );
  NAND2_X1 U2666 ( .A1(n2130), .A2(n2126), .ZN(U3258) );
  NAND2_X1 U2667 ( .A1(n2106), .A2(n4485), .ZN(n2130) );
  AOI21_X1 U2668 ( .B1(n2129), .B2(n2128), .A(n2127), .ZN(n2126) );
  OR2_X1 U2669 ( .A1(n4588), .A2(REG1_REG_28__SCAN_IN), .ZN(n2077) );
  INV_X1 U2670 ( .A(n3758), .ZN(n2188) );
  OR3_X1 U2671 ( .A1(n4051), .A2(n2047), .A3(n2085), .ZN(n2009) );
  OR2_X1 U2672 ( .A1(n3928), .A2(n3910), .ZN(n2010) );
  AND2_X1 U2673 ( .A1(n4016), .A2(n3607), .ZN(n2011) );
  NAND2_X1 U2674 ( .A1(n3753), .A2(n3326), .ZN(n2012) );
  AND2_X1 U2675 ( .A1(n2010), .A2(n2490), .ZN(n2013) );
  AND2_X1 U2676 ( .A1(n2163), .A2(n2039), .ZN(n2014) );
  NAND2_X1 U2677 ( .A1(n2158), .A2(n2044), .ZN(n2016) );
  NOR2_X1 U2678 ( .A1(n3358), .A2(n3357), .ZN(n2017) );
  AND2_X1 U2679 ( .A1(n3944), .A2(n3605), .ZN(n2489) );
  NAND2_X1 U2680 ( .A1(n3535), .A2(n2156), .ZN(n2018) );
  AND2_X1 U2681 ( .A1(n3064), .A2(n3077), .ZN(n2019) );
  AND2_X1 U2682 ( .A1(n2093), .A2(n4285), .ZN(n2020) );
  AND2_X1 U2683 ( .A1(n2123), .A2(n2124), .ZN(n2021) );
  AND2_X1 U2684 ( .A1(n2627), .A2(n2259), .ZN(n2022) );
  OR2_X1 U2685 ( .A1(n2806), .A2(n4534), .ZN(n2023) );
  AND2_X1 U2686 ( .A1(n2259), .A2(n2260), .ZN(n2284) );
  XNOR2_X1 U2687 ( .A(n2533), .B(n2239), .ZN(n2536) );
  AND2_X1 U2688 ( .A1(n3756), .A2(n3100), .ZN(n2024) );
  OR2_X1 U2689 ( .A1(n4478), .A2(n4477), .ZN(n2106) );
  NAND2_X1 U2690 ( .A1(n2284), .A2(REG0_REG_1__SCAN_IN), .ZN(n2025) );
  AND2_X1 U2691 ( .A1(n3928), .A2(n3910), .ZN(n2026) );
  AND2_X1 U2692 ( .A1(n3883), .A2(n3872), .ZN(n2027) );
  INV_X1 U2693 ( .A(IR_REG_29__SCAN_IN), .ZN(n2257) );
  OR2_X1 U2694 ( .A1(n3236), .A2(n4529), .ZN(n2028) );
  OR2_X1 U2695 ( .A1(IR_REG_20__SCAN_IN), .A2(IR_REG_19__SCAN_IN), .ZN(n2029)
         );
  AND2_X1 U2696 ( .A1(n2551), .A2(n3655), .ZN(n3627) );
  AND2_X1 U2697 ( .A1(n3122), .A2(n3124), .ZN(n3628) );
  NOR2_X1 U2698 ( .A1(n4035), .A2(n4015), .ZN(n2030) );
  AND2_X1 U2699 ( .A1(n3115), .A2(n3162), .ZN(n2031) );
  NAND2_X1 U2700 ( .A1(n3565), .A2(n4002), .ZN(n2032) );
  NAND2_X1 U2701 ( .A1(n3644), .A2(n3647), .ZN(n2546) );
  OR2_X1 U2702 ( .A1(n2489), .A2(n2026), .ZN(n2033) );
  OR2_X1 U2703 ( .A1(n3154), .A2(n3118), .ZN(n2034) );
  AND2_X1 U2704 ( .A1(n2856), .A2(n3483), .ZN(n2035) );
  AND2_X1 U2705 ( .A1(n2071), .A2(n2070), .ZN(n2036) );
  AND2_X1 U2706 ( .A1(n3034), .A2(n3029), .ZN(n2037) );
  INV_X1 U2707 ( .A(n2502), .ZN(n2195) );
  INV_X1 U2708 ( .A(IR_REG_17__SCAN_IN), .ZN(n2242) );
  OAI21_X1 U2709 ( .B1(n3178), .B2(n2143), .A(n2141), .ZN(n3279) );
  OR2_X1 U2710 ( .A1(n3400), .A2(n3399), .ZN(n2038) );
  INV_X1 U2711 ( .A(n2979), .ZN(n2187) );
  INV_X1 U2712 ( .A(n3621), .ZN(n2205) );
  INV_X1 U2713 ( .A(IR_REG_22__SCAN_IN), .ZN(n2239) );
  INV_X1 U2714 ( .A(n3351), .ZN(n2166) );
  NOR2_X1 U2715 ( .A1(n3553), .A2(n3554), .ZN(n3471) );
  INV_X1 U2716 ( .A(IR_REG_21__SCAN_IN), .ZN(n2240) );
  NAND2_X1 U2717 ( .A1(n2400), .A2(n2399), .ZN(n3202) );
  INV_X1 U2718 ( .A(n3516), .ZN(n2148) );
  INV_X1 U2719 ( .A(n3640), .ZN(n2084) );
  OR2_X1 U2720 ( .A1(n3526), .A2(n3525), .ZN(n2039) );
  NOR2_X1 U2721 ( .A1(n2447), .A2(IR_REG_18__SCAN_IN), .ZN(n2458) );
  NAND2_X1 U2722 ( .A1(n2247), .A2(n2246), .ZN(n2435) );
  INV_X1 U2723 ( .A(n2142), .ZN(n2141) );
  OAI21_X1 U2724 ( .B1(n3177), .B2(n2143), .A(n3190), .ZN(n2142) );
  AND2_X1 U2725 ( .A1(n2215), .A2(n2213), .ZN(n2040) );
  OR2_X1 U2726 ( .A1(n2017), .A2(n2166), .ZN(n2041) );
  AND2_X1 U2727 ( .A1(n4356), .A2(n4354), .ZN(n2042) );
  NAND2_X1 U2728 ( .A1(n4063), .A2(n4042), .ZN(n2043) );
  OR2_X1 U2729 ( .A1(n3471), .A2(n2159), .ZN(n2158) );
  OAI21_X1 U2730 ( .B1(n3535), .B2(n2156), .A(n2038), .ZN(n2157) );
  INV_X1 U2731 ( .A(n3404), .ZN(n2156) );
  AND2_X1 U2732 ( .A1(n2038), .A2(n2156), .ZN(n2044) );
  AND2_X1 U2733 ( .A1(n2092), .A2(n3142), .ZN(n2045) );
  AND2_X1 U2734 ( .A1(n2117), .A2(n2113), .ZN(n2046) );
  INV_X1 U2735 ( .A(n2489), .ZN(n2199) );
  INV_X1 U2736 ( .A(n4507), .ZN(n4027) );
  INV_X1 U2737 ( .A(n4588), .ZN(n4586) );
  INV_X1 U2738 ( .A(n3306), .ZN(n2076) );
  XNOR2_X1 U2739 ( .A(n2588), .B(IR_REG_25__SCAN_IN), .ZN(n2592) );
  NAND2_X1 U2740 ( .A1(n2171), .A2(n2169), .ZN(n3112) );
  OR2_X1 U2741 ( .A1(n3607), .A2(n3609), .ZN(n2047) );
  OR2_X1 U2742 ( .A1(n4051), .A2(n4042), .ZN(n2048) );
  OAI21_X1 U2743 ( .B1(n3051), .B2(n2024), .A(n2367), .ZN(n3136) );
  NOR3_X1 U2744 ( .A1(n3959), .A2(n2095), .A3(n3882), .ZN(n2097) );
  NAND2_X1 U2745 ( .A1(n2203), .A2(n2301), .ZN(n2936) );
  NOR2_X1 U2746 ( .A1(n4402), .A2(n3234), .ZN(n2049) );
  INV_X1 U2747 ( .A(n2062), .ZN(n2061) );
  NOR2_X1 U2748 ( .A1(n2991), .A2(n2063), .ZN(n2062) );
  INV_X1 U2749 ( .A(n2096), .ZN(n4246) );
  NOR2_X1 U2750 ( .A1(n3959), .A2(n3953), .ZN(n2096) );
  INV_X1 U2751 ( .A(n2094), .ZN(n3907) );
  NOR2_X1 U2752 ( .A1(n3959), .A2(n2095), .ZN(n2094) );
  INV_X1 U2753 ( .A(n2012), .ZN(n2207) );
  AND2_X1 U2754 ( .A1(n2108), .A2(n2023), .ZN(n2050) );
  AND2_X1 U2755 ( .A1(n2206), .A2(n2012), .ZN(n2051) );
  AND2_X1 U2756 ( .A1(n2981), .A2(n2092), .ZN(n2052) );
  NAND2_X1 U2757 ( .A1(n2202), .A2(IR_REG_31__SCAN_IN), .ZN(n2255) );
  NAND2_X1 U2758 ( .A1(n2255), .A2(n2254), .ZN(n2537) );
  NAND2_X1 U2759 ( .A1(n2543), .A2(n2885), .ZN(n2760) );
  OR2_X1 U2760 ( .A1(n4284), .A2(n4083), .ZN(n2053) );
  XNOR2_X1 U2761 ( .A(n2818), .B(n2816), .ZN(n2815) );
  NAND2_X1 U2762 ( .A1(n4484), .A2(n4483), .ZN(n2054) );
  INV_X1 U2763 ( .A(n3763), .ZN(n2755) );
  XNOR2_X1 U2764 ( .A(n2255), .B(n2625), .ZN(n3832) );
  NAND3_X1 U2765 ( .A1(n2882), .A2(n3015), .A3(n2764), .ZN(n2925) );
  NAND3_X1 U2766 ( .A1(n3933), .A2(n3947), .A3(n4236), .ZN(n2095) );
  INV_X1 U2767 ( .A(n2097), .ZN(n3887) );
  NAND2_X1 U2768 ( .A1(n3800), .A2(n2115), .ZN(n2114) );
  INV_X1 U2769 ( .A(n2117), .ZN(n4430) );
  NAND3_X1 U2770 ( .A1(n4169), .A2(n2132), .A3(n2131), .ZN(n2296) );
  OAI22_X1 U2771 ( .A1(n2805), .A2(n2804), .B1(n4336), .B2(REG1_REG_7__SCAN_IN), .ZN(n2806) );
  XNOR2_X1 U2772 ( .A(n3803), .B(n2427), .ZN(n4456) );
  AOI21_X1 U2773 ( .B1(n2696), .B2(REG1_REG_5__SCAN_IN), .A(n2710), .ZN(n2698)
         );
  OR2_X2 U2774 ( .A1(n4433), .A2(n3813), .ZN(n2120) );
  NAND2_X1 U2775 ( .A1(n4372), .A2(n2124), .ZN(n2122) );
  INV_X1 U2776 ( .A(n2682), .ZN(n2708) );
  NAND2_X1 U2777 ( .A1(n2681), .A2(n4377), .ZN(n2124) );
  INV_X1 U2778 ( .A(REG2_REG_4__SCAN_IN), .ZN(n2125) );
  INV_X1 U2779 ( .A(IR_REG_0__SCAN_IN), .ZN(n2132) );
  INV_X1 U2780 ( .A(IR_REG_1__SCAN_IN), .ZN(n2131) );
  INV_X1 U2781 ( .A(n2296), .ZN(n2230) );
  NAND2_X1 U2782 ( .A1(n3482), .A2(n3483), .ZN(n2840) );
  NAND3_X1 U2783 ( .A1(n2134), .A2(n2894), .A3(n2133), .ZN(n2900) );
  NAND2_X1 U2784 ( .A1(n3482), .A2(n2035), .ZN(n2133) );
  INV_X1 U2785 ( .A(n2856), .ZN(n2135) );
  OR2_X1 U2786 ( .A1(n3471), .A2(n2150), .ZN(n2149) );
  NAND2_X1 U2787 ( .A1(n3352), .A2(n2014), .ZN(n2162) );
  NAND2_X1 U2788 ( .A1(n3352), .A2(n3351), .ZN(n4353) );
  NOR2_X1 U2789 ( .A1(n3352), .A2(n3351), .ZN(n4352) );
  NAND2_X1 U2790 ( .A1(n2168), .A2(n2037), .ZN(n3065) );
  INV_X1 U2791 ( .A(n2447), .ZN(n2529) );
  INV_X1 U2792 ( .A(n4030), .ZN(n2175) );
  NAND2_X1 U2793 ( .A1(n2185), .A2(n2183), .ZN(n2963) );
  NAND2_X1 U2794 ( .A1(n3914), .A2(n2192), .ZN(n2191) );
  NAND2_X1 U2795 ( .A1(n2247), .A2(n2244), .ZN(n2202) );
  NAND3_X1 U2796 ( .A1(n2203), .A2(n2301), .A3(n2933), .ZN(n2935) );
  NAND2_X1 U2797 ( .A1(n2206), .A2(n2204), .ZN(n3246) );
  XNOR2_X1 U2798 ( .A(n2586), .B(n2585), .ZN(n2591) );
  NAND2_X1 U2799 ( .A1(n2584), .A2(IR_REG_31__SCAN_IN), .ZN(n2586) );
  AOI21_X2 U2800 ( .B1(n3301), .B2(n2414), .A(n2413), .ZN(n4049) );
  AOI21_X2 U2801 ( .B1(n2517), .B2(n2226), .A(n2225), .ZN(n3838) );
  AOI22_X2 U2802 ( .A1(n3978), .A2(n2470), .B1(n3609), .B2(n3966), .ZN(n3958)
         );
  AND2_X1 U2803 ( .A1(n2879), .A2(n2007), .ZN(n2219) );
  AND2_X1 U2804 ( .A1(n2297), .A2(n2229), .ZN(n2220) );
  OR2_X1 U2805 ( .A1(n3323), .A2(n3257), .ZN(n2221) );
  OR2_X1 U2806 ( .A1(n3586), .A2(n4348), .ZN(n2222) );
  OR2_X1 U2807 ( .A1(n3443), .A2(n4332), .ZN(n2223) );
  OR2_X1 U2808 ( .A1(n3443), .A2(n4289), .ZN(n2224) );
  AND2_X1 U2809 ( .A1(n3867), .A2(n3855), .ZN(n2225) );
  OR2_X1 U2810 ( .A1(n3867), .A2(n3855), .ZN(n2226) );
  OR2_X1 U2811 ( .A1(n3926), .A2(n3947), .ZN(n2227) );
  OAI21_X2 U2812 ( .B1(n2583), .B2(n2582), .A(IR_REG_31__SCAN_IN), .ZN(n2595)
         );
  NAND2_X1 U2813 ( .A1(n2529), .A2(n2015), .ZN(n2583) );
  NAND2_X1 U2814 ( .A1(n2787), .A2(n2786), .ZN(n2788) );
  OR2_X1 U2815 ( .A1(n3754), .A2(n3130), .ZN(n2399) );
  INV_X1 U2816 ( .A(n2546), .ZN(n3596) );
  AND2_X1 U2817 ( .A1(n2829), .A2(n2733), .ZN(n2729) );
  INV_X1 U2818 ( .A(IR_REG_13__SCAN_IN), .ZN(n2236) );
  INV_X1 U2819 ( .A(n3068), .ZN(n3034) );
  INV_X1 U2820 ( .A(n2854), .ZN(n2855) );
  INV_X1 U2821 ( .A(n4437), .ZN(n3798) );
  AND2_X1 U2822 ( .A1(n3898), .A2(n3888), .ZN(n3694) );
  OR2_X1 U2823 ( .A1(n2491), .A2(n3537), .ZN(n2495) );
  NAND2_X1 U2824 ( .A1(n2310), .A2(REG3_REG_5__SCAN_IN), .ZN(n2321) );
  NAND2_X1 U2825 ( .A1(n2330), .A2(REG3_REG_7__SCAN_IN), .ZN(n2343) );
  AND2_X1 U2826 ( .A1(n3276), .A2(n3314), .ZN(n3277) );
  OR2_X1 U2827 ( .A1(n2387), .A2(n2386), .ZN(n2389) );
  INV_X1 U2828 ( .A(n4062), .ZN(n4342) );
  NOR2_X1 U2829 ( .A1(n2356), .A2(n2355), .ZN(n2368) );
  NAND2_X1 U2830 ( .A1(n2376), .A2(REG3_REG_11__SCAN_IN), .ZN(n2387) );
  NOR2_X1 U2831 ( .A1(n2439), .A2(n4202), .ZN(n2450) );
  INV_X1 U2832 ( .A(n3898), .ZN(n3865) );
  OR2_X1 U2833 ( .A1(n2389), .A2(n3231), .ZN(n2404) );
  INV_X1 U2834 ( .A(REG3_REG_6__SCAN_IN), .ZN(n2912) );
  INV_X1 U2835 ( .A(REG3_REG_18__SCAN_IN), .ZN(n4202) );
  NOR2_X1 U2836 ( .A1(n2504), .A2(n4094), .ZN(n2519) );
  AND2_X1 U2837 ( .A1(n4342), .A2(n3305), .ZN(n2413) );
  OR2_X1 U2838 ( .A1(n2343), .A2(n2342), .ZN(n2356) );
  INV_X1 U2839 ( .A(n2646), .ZN(n2740) );
  OR2_X1 U2840 ( .A1(n3697), .A2(n3732), .ZN(n3850) );
  OR2_X1 U2841 ( .A1(n3006), .A2(n2576), .ZN(n4284) );
  XNOR2_X1 U2842 ( .A(n2581), .B(IR_REG_26__SCAN_IN), .ZN(n2593) );
  OR3_X1 U2843 ( .A1(n2362), .A2(IR_REG_7__SCAN_IN), .A3(IR_REG_8__SCAN_IN), 
        .ZN(n2365) );
  INV_X1 U2844 ( .A(n3933), .ZN(n3605) );
  AND2_X1 U2845 ( .A1(n2450), .A2(REG3_REG_19__SCAN_IN), .ZN(n2463) );
  NAND2_X1 U2846 ( .A1(n2415), .A2(REG3_REG_16__SCAN_IN), .ZN(n2428) );
  INV_X1 U2847 ( .A(n4038), .ZN(n4042) );
  INV_X1 U2848 ( .A(n3267), .ZN(n3326) );
  INV_X1 U2849 ( .A(n4362), .ZN(n3578) );
  NAND4_X1 U2850 ( .A1(n2265), .A2(n2264), .A3(n2263), .A4(n2262), .ZN(n3283)
         );
  AND2_X1 U2851 ( .A1(n2654), .A2(n2655), .ZN(n2667) );
  AND2_X1 U2852 ( .A1(n2667), .A2(n4341), .ZN(n4484) );
  INV_X1 U2853 ( .A(n4284), .ZN(n4277) );
  NAND2_X1 U2854 ( .A1(n3941), .A2(n3942), .ZN(n3940) );
  AND2_X1 U2855 ( .A1(n4341), .A2(n2651), .ZN(n4064) );
  INV_X1 U2856 ( .A(n4070), .ZN(n3979) );
  AND2_X1 U2857 ( .A1(n3649), .A2(n3646), .ZN(n3595) );
  AOI21_X1 U2858 ( .B1(n2740), .B2(n3454), .A(n2613), .ZN(n2741) );
  INV_X1 U2859 ( .A(n3607), .ZN(n4002) );
  INV_X1 U2860 ( .A(n4559), .ZN(n4574) );
  AND3_X1 U2861 ( .A1(n2611), .A2(n2610), .A3(n2609), .ZN(n2619) );
  XNOR2_X1 U2862 ( .A(n2316), .B(n4162), .ZN(n2714) );
  AND2_X1 U2863 ( .A1(n2656), .A2(n2655), .ZN(n4462) );
  OR2_X1 U2864 ( .A1(n2751), .A2(n2743), .ZN(n3581) );
  NOR2_X1 U2865 ( .A1(n2727), .A2(n3452), .ZN(U4043) );
  OAI211_X1 U2866 ( .C1(n2008), .C2(n3935), .A(n2488), .B(n2487), .ZN(n3944)
         );
  NAND4_X1 U2867 ( .A1(n2271), .A2(n2270), .A3(n2269), .A4(n2268), .ZN(n3753)
         );
  INV_X1 U2868 ( .A(n4337), .ZN(n2676) );
  INV_X1 U2869 ( .A(n4484), .ZN(n4475) );
  AND2_X1 U2870 ( .A1(n3127), .A2(n3126), .ZN(n3256) );
  OR2_X1 U2871 ( .A1(n4507), .A2(n2966), .ZN(n4070) );
  AND2_X1 U2872 ( .A1(n2875), .A2(n3950), .ZN(n4507) );
  NAND2_X1 U2873 ( .A1(n4588), .A2(n4574), .ZN(n4289) );
  AND2_X2 U2874 ( .A1(n2619), .A2(n2741), .ZN(n4588) );
  NAND2_X1 U2875 ( .A1(n4577), .A2(n4574), .ZN(n4332) );
  INV_X1 U2876 ( .A(n4577), .ZN(n4575) );
  INV_X1 U2877 ( .A(n4517), .ZN(n4516) );
  AND2_X1 U2878 ( .A1(n2843), .A2(STATE_REG_SCAN_IN), .ZN(n4518) );
  INV_X1 U2879 ( .A(n3226), .ZN(n4529) );
  AND2_X1 U2880 ( .A1(n2349), .A2(n2340), .ZN(n4336) );
  NAND2_X1 U2881 ( .A1(n2230), .A2(n2220), .ZN(n2315) );
  NAND4_X1 U2882 ( .A1(n2234), .A2(n2233), .A3(n2232), .A4(n2231), .ZN(n2235)
         );
  OR2_X1 U2883 ( .A1(n2247), .A2(n2457), .ZN(n2237) );
  XNOR2_X1 U2884 ( .A(n2237), .B(IR_REG_14__SCAN_IN), .ZN(n4437) );
  NAND3_X1 U2885 ( .A1(n2596), .A2(n2585), .A3(n2238), .ZN(n2241) );
  NAND2_X1 U2886 ( .A1(n2538), .A2(IR_REG_27__SCAN_IN), .ZN(n2245) );
  MUX2_X1 U2887 ( .A(n4437), .B(DATAI_14_), .S(n2462), .Z(n3284) );
  AND2_X1 U2888 ( .A1(n2538), .A2(n2257), .ZN(n2250) );
  NOR2_X1 U2889 ( .A1(IR_REG_27__SCAN_IN), .A2(IR_REG_26__SCAN_IN), .ZN(n2248)
         );
  AND2_X1 U2890 ( .A1(n2248), .A2(n2579), .ZN(n2249) );
  NAND2_X1 U2891 ( .A1(n2529), .A2(n2252), .ZN(n3448) );
  NAND2_X1 U2892 ( .A1(n3611), .A2(REG0_REG_14__SCAN_IN), .ZN(n2265) );
  NAND2_X1 U2893 ( .A1(n3610), .A2(REG1_REG_14__SCAN_IN), .ZN(n2264) );
  XNOR2_X1 U2894 ( .A(n2404), .B(REG3_REG_14__SCAN_IN), .ZN(n3290) );
  NAND2_X1 U2895 ( .A1(n2006), .A2(n3290), .ZN(n2263) );
  INV_X1 U2896 ( .A(REG2_REG_14__SCAN_IN), .ZN(n2261) );
  OR2_X1 U2897 ( .A1(n2008), .A2(n2261), .ZN(n2262) );
  NAND2_X1 U2898 ( .A1(n3611), .A2(REG0_REG_13__SCAN_IN), .ZN(n2271) );
  NAND2_X1 U2899 ( .A1(n3610), .A2(REG1_REG_13__SCAN_IN), .ZN(n2270) );
  NAND2_X1 U2900 ( .A1(n2389), .A2(n3231), .ZN(n2266) );
  AND2_X1 U2901 ( .A1(n2404), .A2(n2266), .ZN(n3327) );
  NAND2_X1 U2902 ( .A1(n2006), .A2(n3327), .ZN(n2269) );
  INV_X1 U2903 ( .A(REG2_REG_13__SCAN_IN), .ZN(n2267) );
  OR2_X1 U2904 ( .A1(n2008), .A2(n2267), .ZN(n2268) );
  INV_X1 U2905 ( .A(n3753), .ZN(n2401) );
  NOR2_X1 U2906 ( .A1(n2272), .A2(n2457), .ZN(n2273) );
  MUX2_X1 U2907 ( .A(n2457), .B(n2273), .S(IR_REG_13__SCAN_IN), .Z(n2274) );
  OR2_X1 U2908 ( .A1(n2274), .A2(n2247), .ZN(n3244) );
  INV_X1 U2909 ( .A(DATAI_13_), .ZN(n2275) );
  MUX2_X1 U2910 ( .A(n3244), .B(n2275), .S(n2462), .Z(n3267) );
  INV_X1 U2911 ( .A(REG2_REG_1__SCAN_IN), .ZN(n2276) );
  NAND2_X1 U2912 ( .A1(n2282), .A2(REG3_REG_1__SCAN_IN), .ZN(n2277) );
  MUX2_X1 U2913 ( .A(n4339), .B(DATAI_1_), .S(n2462), .Z(n2790) );
  NAND2_X1 U2914 ( .A1(n3763), .A2(n2882), .ZN(n3641) );
  NAND2_X1 U2915 ( .A1(n2755), .A2(n2790), .ZN(n2545) );
  NAND2_X1 U2916 ( .A1(n3641), .A2(n2545), .ZN(n2543) );
  INV_X1 U2917 ( .A(REG2_REG_0__SCAN_IN), .ZN(n3011) );
  OR2_X1 U2918 ( .A1(n2283), .A2(n3011), .ZN(n2280) );
  NAND2_X1 U2919 ( .A1(n2282), .A2(REG3_REG_0__SCAN_IN), .ZN(n2279) );
  NAND2_X1 U2920 ( .A1(n2284), .A2(REG0_REG_0__SCAN_IN), .ZN(n2278) );
  MUX2_X1 U2921 ( .A(IR_REG_0__SCAN_IN), .B(DATAI_0_), .S(n2462), .Z(n2733) );
  AND2_X1 U2922 ( .A1(n2879), .A2(n2733), .ZN(n2885) );
  NAND2_X1 U2923 ( .A1(n2282), .A2(REG3_REG_2__SCAN_IN), .ZN(n2288) );
  INV_X1 U2924 ( .A(REG2_REG_2__SCAN_IN), .ZN(n2668) );
  OR2_X1 U2925 ( .A1(n2283), .A2(n2668), .ZN(n2287) );
  NAND2_X1 U2926 ( .A1(n2022), .A2(REG1_REG_2__SCAN_IN), .ZN(n2286) );
  NAND2_X1 U2927 ( .A1(n2284), .A2(REG0_REG_2__SCAN_IN), .ZN(n2285) );
  MUX2_X1 U2928 ( .A(n4338), .B(DATAI_2_), .S(n2462), .Z(n3459) );
  INV_X1 U2929 ( .A(n3459), .ZN(n2764) );
  NAND2_X1 U2930 ( .A1(n2789), .A2(n2764), .ZN(n3647) );
  NAND2_X1 U2931 ( .A1(n3763), .A2(n2790), .ZN(n2761) );
  NAND2_X1 U2932 ( .A1(n2760), .A2(n2290), .ZN(n2759) );
  NAND2_X1 U2933 ( .A1(n3487), .A2(n2764), .ZN(n2291) );
  NAND2_X1 U2934 ( .A1(n2759), .A2(n2291), .ZN(n2918) );
  INV_X1 U2935 ( .A(REG2_REG_3__SCAN_IN), .ZN(n2927) );
  OR2_X1 U2936 ( .A1(n2008), .A2(n2927), .ZN(n2295) );
  NAND2_X1 U2937 ( .A1(n2022), .A2(REG1_REG_3__SCAN_IN), .ZN(n2294) );
  NAND2_X1 U2938 ( .A1(n2284), .A2(REG0_REG_3__SCAN_IN), .ZN(n2293) );
  INV_X1 U2939 ( .A(REG3_REG_3__SCAN_IN), .ZN(n3490) );
  NAND2_X1 U2940 ( .A1(n2006), .A2(n3490), .ZN(n2292) );
  NAND2_X1 U2941 ( .A1(n2296), .A2(IR_REG_31__SCAN_IN), .ZN(n2298) );
  NAND2_X1 U2942 ( .A1(n2298), .A2(n2297), .ZN(n2307) );
  OR2_X1 U2943 ( .A1(n2298), .A2(n2297), .ZN(n2299) );
  MUX2_X1 U2944 ( .A(n4337), .B(DATAI_3_), .S(n2462), .Z(n2926) );
  NAND2_X1 U2945 ( .A1(n3761), .A2(n2926), .ZN(n2300) );
  INV_X1 U2946 ( .A(n3761), .ZN(n2548) );
  INV_X1 U2947 ( .A(n2926), .ZN(n3485) );
  NAND2_X1 U2948 ( .A1(n2548), .A2(n3485), .ZN(n2301) );
  NAND2_X1 U2949 ( .A1(n2284), .A2(REG0_REG_4__SCAN_IN), .ZN(n2306) );
  NAND2_X1 U2950 ( .A1(n3610), .A2(REG1_REG_4__SCAN_IN), .ZN(n2305) );
  NOR2_X1 U2951 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n2302) );
  NOR2_X1 U2952 ( .A1(n2310), .A2(n2302), .ZN(n2945) );
  NAND2_X1 U2953 ( .A1(n2006), .A2(n2945), .ZN(n2304) );
  OR2_X1 U2954 ( .A1(n2283), .A2(n2125), .ZN(n2303) );
  NAND2_X1 U2955 ( .A1(n2307), .A2(IR_REG_31__SCAN_IN), .ZN(n2308) );
  XNOR2_X1 U2956 ( .A(n2308), .B(IR_REG_4__SCAN_IN), .ZN(n4377) );
  MUX2_X1 U2957 ( .A(n4377), .B(DATAI_4_), .S(n2462), .Z(n2938) );
  NAND2_X1 U2958 ( .A1(n3486), .A2(n2938), .ZN(n3650) );
  NAND2_X1 U2959 ( .A1(n3760), .A2(n2931), .ZN(n3653) );
  NAND2_X1 U2960 ( .A1(n3760), .A2(n2938), .ZN(n2309) );
  NAND2_X1 U2961 ( .A1(n2935), .A2(n2309), .ZN(n2997) );
  NAND2_X1 U2962 ( .A1(n2284), .A2(REG0_REG_5__SCAN_IN), .ZN(n2314) );
  NAND2_X1 U2963 ( .A1(n3610), .A2(REG1_REG_5__SCAN_IN), .ZN(n2313) );
  OAI21_X1 U2964 ( .B1(n2310), .B2(REG3_REG_5__SCAN_IN), .A(n2321), .ZN(n3002)
         );
  INV_X1 U2965 ( .A(n3002), .ZN(n2867) );
  NAND2_X1 U2966 ( .A1(n2006), .A2(n2867), .ZN(n2312) );
  INV_X1 U2967 ( .A(REG2_REG_5__SCAN_IN), .ZN(n2683) );
  OR2_X1 U2968 ( .A1(n2008), .A2(n2683), .ZN(n2311) );
  NAND4_X1 U2969 ( .A1(n2314), .A2(n2313), .A3(n2312), .A4(n2311), .ZN(n3759)
         );
  INV_X1 U2970 ( .A(n3759), .ZN(n2913) );
  NAND2_X1 U2971 ( .A1(n2315), .A2(IR_REG_31__SCAN_IN), .ZN(n2316) );
  INV_X1 U2972 ( .A(DATAI_5_), .ZN(n2317) );
  MUX2_X1 U2973 ( .A(n2714), .B(n2317), .S(n2462), .Z(n3000) );
  NAND2_X1 U2974 ( .A1(n2913), .A2(n3000), .ZN(n2318) );
  NAND2_X1 U2975 ( .A1(n2997), .A2(n2318), .ZN(n2320) );
  NAND2_X1 U2976 ( .A1(n3759), .A2(n2993), .ZN(n2319) );
  NAND2_X1 U2977 ( .A1(n2284), .A2(REG0_REG_6__SCAN_IN), .ZN(n2327) );
  NAND2_X1 U2978 ( .A1(n3610), .A2(REG1_REG_6__SCAN_IN), .ZN(n2326) );
  AND2_X1 U2979 ( .A1(n2321), .A2(n2912), .ZN(n2322) );
  NOR2_X1 U2980 ( .A1(n2330), .A2(n2322), .ZN(n3018) );
  NAND2_X1 U2981 ( .A1(n2006), .A2(n3018), .ZN(n2325) );
  INV_X1 U2982 ( .A(REG2_REG_6__SCAN_IN), .ZN(n2323) );
  OR2_X1 U2983 ( .A1(n2008), .A2(n2323), .ZN(n2324) );
  NAND4_X1 U2984 ( .A1(n2327), .A2(n2326), .A3(n2325), .A4(n2324), .ZN(n3758)
         );
  NOR2_X1 U2985 ( .A1(n2315), .A2(IR_REG_5__SCAN_IN), .ZN(n2337) );
  OR2_X1 U2986 ( .A1(n2337), .A2(n2457), .ZN(n2328) );
  XNOR2_X1 U2987 ( .A(n2328), .B(IR_REG_6__SCAN_IN), .ZN(n2697) );
  MUX2_X1 U2988 ( .A(n2697), .B(DATAI_6_), .S(n2462), .Z(n2979) );
  AND2_X1 U2989 ( .A1(n3758), .A2(n2979), .ZN(n2329) );
  NAND2_X1 U2990 ( .A1(n2284), .A2(REG0_REG_7__SCAN_IN), .ZN(n2335) );
  NAND2_X1 U2991 ( .A1(n3610), .A2(REG1_REG_7__SCAN_IN), .ZN(n2334) );
  OR2_X1 U2992 ( .A1(n2330), .A2(REG3_REG_7__SCAN_IN), .ZN(n2331) );
  AND2_X1 U2993 ( .A1(n2343), .A2(n2331), .ZN(n3071) );
  NAND2_X1 U2994 ( .A1(n2006), .A2(n3071), .ZN(n2333) );
  INV_X1 U2995 ( .A(REG2_REG_7__SCAN_IN), .ZN(n2686) );
  OR2_X1 U2996 ( .A1(n2008), .A2(n2686), .ZN(n2332) );
  NAND4_X1 U2997 ( .A1(n2335), .A2(n2334), .A3(n2333), .A4(n2332), .ZN(n3046)
         );
  INV_X1 U2998 ( .A(n3046), .ZN(n3078) );
  NAND2_X1 U2999 ( .A1(n2337), .A2(n2336), .ZN(n2362) );
  NAND2_X1 U3000 ( .A1(n2362), .A2(IR_REG_31__SCAN_IN), .ZN(n2339) );
  NAND2_X1 U3001 ( .A1(n2339), .A2(n2338), .ZN(n2349) );
  OR2_X1 U3002 ( .A1(n2339), .A2(n2338), .ZN(n2340) );
  MUX2_X1 U3003 ( .A(n4336), .B(DATAI_7_), .S(n2462), .Z(n3033) );
  NAND2_X1 U3004 ( .A1(n3078), .A2(n3033), .ZN(n2551) );
  NAND2_X1 U3005 ( .A1(n3046), .A2(n3064), .ZN(n3655) );
  NAND2_X1 U3006 ( .A1(n3046), .A2(n3033), .ZN(n2341) );
  NAND2_X1 U3007 ( .A1(n2963), .A2(n2341), .ZN(n3075) );
  NAND2_X1 U3008 ( .A1(n3611), .A2(REG0_REG_8__SCAN_IN), .ZN(n2348) );
  NAND2_X1 U3009 ( .A1(n3610), .A2(REG1_REG_8__SCAN_IN), .ZN(n2347) );
  NAND2_X1 U3010 ( .A1(n2343), .A2(n2342), .ZN(n2344) );
  AND2_X1 U3011 ( .A1(n2356), .A2(n2344), .ZN(n4498) );
  NAND2_X1 U3012 ( .A1(n2006), .A2(n4498), .ZN(n2346) );
  INV_X1 U3013 ( .A(REG2_REG_8__SCAN_IN), .ZN(n4211) );
  OR2_X1 U3014 ( .A1(n2008), .A2(n4211), .ZN(n2345) );
  NAND4_X1 U3015 ( .A1(n2348), .A2(n2347), .A3(n2346), .A4(n2345), .ZN(n3757)
         );
  NAND2_X1 U3016 ( .A1(n2349), .A2(IR_REG_31__SCAN_IN), .ZN(n2351) );
  INV_X1 U3017 ( .A(IR_REG_8__SCAN_IN), .ZN(n2350) );
  XNOR2_X1 U3018 ( .A(n2351), .B(n2350), .ZN(n4534) );
  INV_X1 U3019 ( .A(DATAI_8_), .ZN(n4214) );
  MUX2_X1 U3020 ( .A(n4534), .B(n4214), .S(n2462), .Z(n3077) );
  NAND2_X1 U3021 ( .A1(n3097), .A2(n3077), .ZN(n2352) );
  NAND2_X1 U3022 ( .A1(n3075), .A2(n2352), .ZN(n2354) );
  INV_X1 U3023 ( .A(n3077), .ZN(n2553) );
  NAND2_X1 U3024 ( .A1(n3757), .A2(n2553), .ZN(n2353) );
  NAND2_X1 U3025 ( .A1(n3611), .A2(REG0_REG_9__SCAN_IN), .ZN(n2361) );
  NAND2_X1 U3026 ( .A1(n3610), .A2(REG1_REG_9__SCAN_IN), .ZN(n2360) );
  AND2_X1 U3027 ( .A1(n2356), .A2(n2355), .ZN(n2357) );
  NOR2_X1 U3028 ( .A1(n2368), .A2(n2357), .ZN(n3101) );
  NAND2_X1 U3029 ( .A1(n2006), .A2(n3101), .ZN(n2359) );
  INV_X1 U3030 ( .A(REG2_REG_9__SCAN_IN), .ZN(n3058) );
  OR2_X1 U3031 ( .A1(n2008), .A2(n3058), .ZN(n2358) );
  NAND4_X1 U3032 ( .A1(n2361), .A2(n2360), .A3(n2359), .A4(n2358), .ZN(n3756)
         );
  NAND2_X1 U3033 ( .A1(n2365), .A2(IR_REG_31__SCAN_IN), .ZN(n2363) );
  MUX2_X1 U3034 ( .A(IR_REG_31__SCAN_IN), .B(n2363), .S(IR_REG_9__SCAN_IN), 
        .Z(n2364) );
  INV_X1 U3035 ( .A(n2364), .ZN(n2366) );
  MUX2_X1 U3036 ( .A(n4335), .B(DATAI_9_), .S(n2462), .Z(n3100) );
  INV_X1 U3037 ( .A(n3756), .ZN(n3116) );
  INV_X1 U3038 ( .A(n3100), .ZN(n3053) );
  NAND2_X1 U3039 ( .A1(n3116), .A2(n3053), .ZN(n2367) );
  NOR2_X1 U3040 ( .A1(n2368), .A2(REG3_REG_10__SCAN_IN), .ZN(n2369) );
  OR2_X1 U3041 ( .A1(n2376), .A2(n2369), .ZN(n3121) );
  INV_X1 U3042 ( .A(n3121), .ZN(n4490) );
  NAND2_X1 U3043 ( .A1(n2006), .A2(n4490), .ZN(n2374) );
  NAND2_X1 U3044 ( .A1(n3610), .A2(REG1_REG_10__SCAN_IN), .ZN(n2373) );
  NAND2_X1 U3045 ( .A1(n3611), .A2(REG0_REG_10__SCAN_IN), .ZN(n2372) );
  INV_X1 U3046 ( .A(REG2_REG_10__SCAN_IN), .ZN(n2370) );
  OR2_X1 U3047 ( .A1(n2008), .A2(n2370), .ZN(n2371) );
  NAND4_X1 U3048 ( .A1(n2374), .A2(n2373), .A3(n2372), .A4(n2371), .ZN(n3154)
         );
  OR2_X1 U3049 ( .A1(n2384), .A2(n2457), .ZN(n2375) );
  XNOR2_X1 U3050 ( .A(n2375), .B(IR_REG_10__SCAN_IN), .ZN(n3222) );
  MUX2_X1 U3051 ( .A(n3222), .B(DATAI_10_), .S(n2462), .Z(n3118) );
  INV_X1 U3052 ( .A(n3118), .ZN(n3142) );
  NAND2_X1 U3053 ( .A1(n3611), .A2(REG0_REG_11__SCAN_IN), .ZN(n2382) );
  NAND2_X1 U3054 ( .A1(n3610), .A2(REG1_REG_11__SCAN_IN), .ZN(n2381) );
  OR2_X1 U3055 ( .A1(n2376), .A2(REG3_REG_11__SCAN_IN), .ZN(n2377) );
  AND2_X1 U3056 ( .A1(n2387), .A2(n2377), .ZN(n3184) );
  NAND2_X1 U3057 ( .A1(n2006), .A2(n3184), .ZN(n2380) );
  INV_X1 U3058 ( .A(REG2_REG_11__SCAN_IN), .ZN(n2378) );
  OR2_X1 U3059 ( .A1(n2008), .A2(n2378), .ZN(n2379) );
  NAND4_X1 U3060 ( .A1(n2382), .A2(n2381), .A3(n2380), .A4(n2379), .ZN(n3755)
         );
  INV_X1 U3061 ( .A(IR_REG_10__SCAN_IN), .ZN(n2383) );
  NAND2_X1 U3062 ( .A1(n2384), .A2(n2383), .ZN(n2385) );
  NAND2_X1 U3063 ( .A1(n2385), .A2(IR_REG_31__SCAN_IN), .ZN(n2396) );
  MUX2_X1 U3064 ( .A(n3235), .B(DATAI_11_), .S(n2462), .Z(n3183) );
  NAND2_X1 U3065 ( .A1(n3115), .A2(n3183), .ZN(n3122) );
  NAND2_X1 U3066 ( .A1(n3755), .A2(n3162), .ZN(n3124) );
  NAND2_X1 U3067 ( .A1(n3611), .A2(REG0_REG_12__SCAN_IN), .ZN(n2394) );
  NAND2_X1 U3068 ( .A1(n3610), .A2(REG1_REG_12__SCAN_IN), .ZN(n2393) );
  NAND2_X1 U3069 ( .A1(n2387), .A2(n2386), .ZN(n2388) );
  AND2_X1 U3070 ( .A1(n2389), .A2(n2388), .ZN(n3199) );
  NAND2_X1 U3071 ( .A1(n2006), .A2(n3199), .ZN(n2392) );
  INV_X1 U3072 ( .A(REG2_REG_12__SCAN_IN), .ZN(n2390) );
  OR2_X1 U3073 ( .A1(n2008), .A2(n2390), .ZN(n2391) );
  NAND4_X1 U3074 ( .A1(n2394), .A2(n2393), .A3(n2392), .A4(n2391), .ZN(n3754)
         );
  INV_X1 U3075 ( .A(IR_REG_11__SCAN_IN), .ZN(n2395) );
  NAND2_X1 U3076 ( .A1(n2396), .A2(n2395), .ZN(n2397) );
  NAND2_X1 U3077 ( .A1(n2397), .A2(IR_REG_31__SCAN_IN), .ZN(n2398) );
  XNOR2_X1 U3078 ( .A(n2398), .B(IR_REG_12__SCAN_IN), .ZN(n3226) );
  INV_X1 U3079 ( .A(DATAI_12_), .ZN(n4528) );
  MUX2_X1 U3080 ( .A(n4529), .B(n4528), .S(n2462), .Z(n3257) );
  NAND2_X1 U3081 ( .A1(n3128), .A2(n2221), .ZN(n2400) );
  INV_X1 U3082 ( .A(n3257), .ZN(n3130) );
  NAND2_X1 U3083 ( .A1(n3587), .A2(n3284), .ZN(n3637) );
  INV_X1 U3084 ( .A(n3284), .ZN(n4285) );
  NAND2_X1 U3085 ( .A1(n3283), .A2(n4285), .ZN(n3634) );
  NAND2_X1 U3086 ( .A1(n3637), .A2(n3634), .ZN(n3621) );
  OAI21_X1 U3087 ( .B1(n3284), .B2(n3283), .A(n3246), .ZN(n3301) );
  NAND2_X1 U3088 ( .A1(n3611), .A2(REG0_REG_15__SCAN_IN), .ZN(n2410) );
  NAND2_X1 U3089 ( .A1(n2022), .A2(REG1_REG_15__SCAN_IN), .ZN(n2409) );
  INV_X1 U3090 ( .A(n2404), .ZN(n2402) );
  AOI21_X1 U3091 ( .B1(n2402), .B2(REG3_REG_14__SCAN_IN), .A(
        REG3_REG_15__SCAN_IN), .ZN(n2405) );
  NAND2_X1 U3092 ( .A1(REG3_REG_14__SCAN_IN), .A2(REG3_REG_15__SCAN_IN), .ZN(
        n2403) );
  OR2_X1 U3093 ( .A1(n2405), .A2(n2415), .ZN(n3592) );
  INV_X1 U3094 ( .A(n3592), .ZN(n3303) );
  NAND2_X1 U3095 ( .A1(n2006), .A2(n3303), .ZN(n2408) );
  INV_X1 U3096 ( .A(REG2_REG_15__SCAN_IN), .ZN(n2406) );
  OR2_X1 U3097 ( .A1(n2008), .A2(n2406), .ZN(n2407) );
  INV_X1 U3098 ( .A(IR_REG_14__SCAN_IN), .ZN(n2411) );
  NAND2_X1 U3099 ( .A1(n2247), .A2(n2411), .ZN(n2412) );
  NAND2_X1 U3100 ( .A1(n2412), .A2(IR_REG_31__SCAN_IN), .ZN(n2423) );
  XNOR2_X1 U3101 ( .A(n2423), .B(IR_REG_15__SCAN_IN), .ZN(n3814) );
  NAND2_X1 U3102 ( .A1(n4062), .A2(n4278), .ZN(n2414) );
  INV_X1 U3103 ( .A(n4278), .ZN(n3305) );
  OR2_X1 U3104 ( .A1(n2415), .A2(REG3_REG_16__SCAN_IN), .ZN(n2416) );
  NAND2_X1 U3105 ( .A1(n2428), .A2(n2416), .ZN(n4361) );
  INV_X1 U3106 ( .A(n4361), .ZN(n4054) );
  NAND2_X1 U3107 ( .A1(n2006), .A2(n4054), .ZN(n2421) );
  NAND2_X1 U3108 ( .A1(n2022), .A2(REG1_REG_16__SCAN_IN), .ZN(n2420) );
  NAND2_X1 U3109 ( .A1(n3611), .A2(REG0_REG_16__SCAN_IN), .ZN(n2419) );
  INV_X1 U3110 ( .A(REG2_REG_16__SCAN_IN), .ZN(n2417) );
  OR2_X1 U3111 ( .A1(n2008), .A2(n2417), .ZN(n2418) );
  NAND4_X1 U3112 ( .A1(n2421), .A2(n2420), .A3(n2419), .A4(n2418), .ZN(n4034)
         );
  INV_X1 U3113 ( .A(IR_REG_15__SCAN_IN), .ZN(n2422) );
  NAND2_X1 U3114 ( .A1(n2423), .A2(n2422), .ZN(n2424) );
  NAND2_X1 U3115 ( .A1(n2424), .A2(IR_REG_31__SCAN_IN), .ZN(n2426) );
  INV_X1 U3116 ( .A(IR_REG_16__SCAN_IN), .ZN(n2425) );
  XNOR2_X1 U3117 ( .A(n2426), .B(n2425), .ZN(n4524) );
  INV_X1 U3118 ( .A(n4524), .ZN(n2427) );
  MUX2_X1 U3119 ( .A(n2427), .B(DATAI_16_), .S(n2462), .Z(n4272) );
  NAND2_X1 U3120 ( .A1(n3586), .A2(n4272), .ZN(n3722) );
  NAND2_X1 U3121 ( .A1(n4034), .A2(n4348), .ZN(n3683) );
  NAND2_X1 U3122 ( .A1(n3722), .A2(n3683), .ZN(n4048) );
  NAND2_X1 U3123 ( .A1(n4049), .A2(n4048), .ZN(n4047) );
  NAND2_X1 U3124 ( .A1(n2428), .A2(n4181), .ZN(n2429) );
  AND2_X1 U3125 ( .A1(n2439), .A2(n2429), .ZN(n4041) );
  NAND2_X1 U3126 ( .A1(n2006), .A2(n4041), .ZN(n2434) );
  NAND2_X1 U3127 ( .A1(n3610), .A2(REG1_REG_17__SCAN_IN), .ZN(n2433) );
  NAND2_X1 U3128 ( .A1(n3611), .A2(REG0_REG_17__SCAN_IN), .ZN(n2432) );
  INV_X1 U3129 ( .A(REG2_REG_17__SCAN_IN), .ZN(n2430) );
  OR2_X1 U3130 ( .A1(n2008), .A2(n2430), .ZN(n2431) );
  NAND4_X1 U3131 ( .A1(n2434), .A2(n2433), .A3(n2432), .A4(n2431), .ZN(n4063)
         );
  NAND2_X1 U3132 ( .A1(n2435), .A2(IR_REG_31__SCAN_IN), .ZN(n2436) );
  XNOR2_X1 U3133 ( .A(n2436), .B(IR_REG_17__SCAN_IN), .ZN(n3817) );
  INV_X1 U3134 ( .A(DATAI_17_), .ZN(n2437) );
  MUX2_X1 U3135 ( .A(n4522), .B(n2437), .S(n2462), .Z(n4038) );
  NAND2_X1 U3136 ( .A1(n4345), .A2(n4038), .ZN(n2438) );
  NAND2_X1 U3137 ( .A1(n3611), .A2(REG0_REG_18__SCAN_IN), .ZN(n2445) );
  NAND2_X1 U3138 ( .A1(n3610), .A2(REG1_REG_18__SCAN_IN), .ZN(n2444) );
  AND2_X1 U3139 ( .A1(n2439), .A2(n4202), .ZN(n2440) );
  NOR2_X1 U3140 ( .A1(n2450), .A2(n2440), .ZN(n4023) );
  NAND2_X1 U3141 ( .A1(n2006), .A2(n4023), .ZN(n2443) );
  INV_X1 U3142 ( .A(REG2_REG_18__SCAN_IN), .ZN(n2441) );
  OR2_X1 U3143 ( .A1(n2008), .A2(n2441), .ZN(n2442) );
  NAND4_X1 U3144 ( .A1(n2445), .A2(n2444), .A3(n2443), .A4(n2442), .ZN(n4035)
         );
  INV_X1 U3145 ( .A(n4035), .ZN(n3529) );
  NAND2_X1 U3146 ( .A1(n2447), .A2(IR_REG_31__SCAN_IN), .ZN(n2446) );
  MUX2_X1 U3147 ( .A(IR_REG_31__SCAN_IN), .B(n2446), .S(IR_REG_18__SCAN_IN), 
        .Z(n2449) );
  INV_X1 U31480 ( .A(n2458), .ZN(n2448) );
  MUX2_X1 U31490 ( .A(n4483), .B(DATAI_18_), .S(n2462), .Z(n4015) );
  NAND2_X1 U3150 ( .A1(n3529), .A2(n4015), .ZN(n3989) );
  INV_X1 U3151 ( .A(n4015), .ZN(n4021) );
  NAND2_X1 U3152 ( .A1(n4035), .A2(n4021), .ZN(n3990) );
  NAND2_X1 U3153 ( .A1(n3989), .A2(n3990), .ZN(n4014) );
  NAND2_X1 U3154 ( .A1(n3611), .A2(REG0_REG_19__SCAN_IN), .ZN(n2456) );
  NAND2_X1 U3155 ( .A1(n3610), .A2(REG1_REG_19__SCAN_IN), .ZN(n2455) );
  NOR2_X1 U3156 ( .A1(n2450), .A2(REG3_REG_19__SCAN_IN), .ZN(n2451) );
  OR2_X1 U3157 ( .A1(n2463), .A2(n2451), .ZN(n3502) );
  INV_X1 U3158 ( .A(n3502), .ZN(n4004) );
  NAND2_X1 U3159 ( .A1(n2006), .A2(n4004), .ZN(n2454) );
  INV_X1 U3160 ( .A(REG2_REG_19__SCAN_IN), .ZN(n2452) );
  OR2_X1 U3161 ( .A1(n2008), .A2(n2452), .ZN(n2453) );
  INV_X1 U3162 ( .A(IR_REG_19__SCAN_IN), .ZN(n2460) );
  MUX2_X1 U3163 ( .A(n4334), .B(DATAI_19_), .S(n2462), .Z(n3607) );
  NAND2_X1 U3164 ( .A1(n3611), .A2(REG0_REG_20__SCAN_IN), .ZN(n2469) );
  NAND2_X1 U3165 ( .A1(n3610), .A2(REG1_REG_20__SCAN_IN), .ZN(n2468) );
  OR2_X1 U3166 ( .A1(n2463), .A2(REG3_REG_20__SCAN_IN), .ZN(n2464) );
  AND2_X1 U3167 ( .A1(n2471), .A2(n2464), .ZN(n3980) );
  NAND2_X1 U3168 ( .A1(n2006), .A2(n3980), .ZN(n2467) );
  INV_X1 U3169 ( .A(REG2_REG_20__SCAN_IN), .ZN(n2465) );
  OR2_X1 U3170 ( .A1(n2008), .A2(n2465), .ZN(n2466) );
  NAND2_X1 U3171 ( .A1(n2462), .A2(DATAI_20_), .ZN(n4256) );
  NAND2_X1 U3172 ( .A1(n3995), .A2(n4256), .ZN(n2470) );
  INV_X1 U3173 ( .A(n4256), .ZN(n3609) );
  INV_X1 U3174 ( .A(REG3_REG_21__SCAN_IN), .ZN(n3511) );
  NAND2_X1 U3175 ( .A1(n2471), .A2(n3511), .ZN(n2472) );
  AND2_X1 U3176 ( .A1(n2480), .A2(n2472), .ZN(n3961) );
  NAND2_X1 U3177 ( .A1(n3961), .A2(n2006), .ZN(n2477) );
  NAND2_X1 U3178 ( .A1(n3611), .A2(REG0_REG_21__SCAN_IN), .ZN(n2476) );
  NAND2_X1 U3179 ( .A1(n3610), .A2(REG1_REG_21__SCAN_IN), .ZN(n2475) );
  INV_X1 U3180 ( .A(REG2_REG_21__SCAN_IN), .ZN(n2473) );
  OR2_X1 U3181 ( .A1(n2008), .A2(n2473), .ZN(n2474) );
  INV_X1 U3182 ( .A(n3974), .ZN(n3752) );
  NAND2_X1 U3183 ( .A1(n3752), .A2(n4250), .ZN(n2479) );
  INV_X1 U3184 ( .A(n4250), .ZN(n3963) );
  INV_X1 U3185 ( .A(REG3_REG_22__SCAN_IN), .ZN(n4196) );
  AND2_X1 U3186 ( .A1(n2480), .A2(n4196), .ZN(n2481) );
  OR2_X1 U3187 ( .A1(n2481), .A2(n2485), .ZN(n3951) );
  AOI22_X1 U3188 ( .A1(n3610), .A2(REG1_REG_22__SCAN_IN), .B1(n3611), .B2(
        REG0_REG_22__SCAN_IN), .ZN(n2484) );
  INV_X1 U3189 ( .A(REG2_REG_22__SCAN_IN), .ZN(n2482) );
  OR2_X1 U3190 ( .A1(n2008), .A2(n2482), .ZN(n2483) );
  NAND2_X1 U3191 ( .A1(n2462), .A2(DATAI_22_), .ZN(n3947) );
  OR2_X1 U3192 ( .A1(n3967), .A2(n3947), .ZN(n3923) );
  NAND2_X1 U3193 ( .A1(n3967), .A2(n3947), .ZN(n2568) );
  NAND2_X1 U3194 ( .A1(n3923), .A2(n2568), .ZN(n3942) );
  INV_X1 U3195 ( .A(n3967), .ZN(n3926) );
  NAND2_X1 U3196 ( .A1(n3940), .A2(n2227), .ZN(n3914) );
  INV_X1 U3197 ( .A(REG2_REG_23__SCAN_IN), .ZN(n3935) );
  OR2_X1 U3198 ( .A1(n2485), .A2(REG3_REG_23__SCAN_IN), .ZN(n2486) );
  NAND2_X1 U3199 ( .A1(n2491), .A2(n2486), .ZN(n3934) );
  AOI22_X1 U3200 ( .A1(n3610), .A2(REG1_REG_23__SCAN_IN), .B1(n3611), .B2(
        REG0_REG_23__SCAN_IN), .ZN(n2487) );
  INV_X1 U3201 ( .A(n3944), .ZN(n3900) );
  NAND2_X1 U3202 ( .A1(n2462), .A2(DATAI_23_), .ZN(n3933) );
  NAND2_X1 U3203 ( .A1(n3900), .A2(n3933), .ZN(n2490) );
  INV_X1 U3204 ( .A(REG2_REG_24__SCAN_IN), .ZN(n3906) );
  INV_X1 U3205 ( .A(REG3_REG_24__SCAN_IN), .ZN(n3537) );
  NAND2_X1 U3206 ( .A1(n2491), .A2(n3537), .ZN(n2492) );
  NAND2_X1 U3207 ( .A1(n2495), .A2(n2492), .ZN(n3905) );
  AOI22_X1 U3208 ( .A1(n3610), .A2(REG1_REG_24__SCAN_IN), .B1(n3611), .B2(
        REG0_REG_24__SCAN_IN), .ZN(n2493) );
  NAND2_X1 U3209 ( .A1(n2462), .A2(DATAI_24_), .ZN(n4236) );
  INV_X1 U32100 ( .A(n4236), .ZN(n3910) );
  INV_X1 U32110 ( .A(REG3_REG_25__SCAN_IN), .ZN(n4096) );
  NAND2_X1 U32120 ( .A1(n2495), .A2(n4096), .ZN(n2496) );
  NAND2_X1 U32130 ( .A1(n3889), .A2(n2006), .ZN(n2501) );
  NAND2_X1 U32140 ( .A1(n3611), .A2(REG0_REG_25__SCAN_IN), .ZN(n2498) );
  NAND2_X1 U32150 ( .A1(n3610), .A2(REG1_REG_25__SCAN_IN), .ZN(n2497) );
  OAI211_X1 U32160 ( .C1(n4149), .C2(n2008), .A(n2498), .B(n2497), .ZN(n2499)
         );
  INV_X1 U32170 ( .A(n2499), .ZN(n2500) );
  NAND2_X1 U32180 ( .A1(n2462), .A2(DATAI_25_), .ZN(n3888) );
  NAND2_X1 U32190 ( .A1(n3865), .A2(n3888), .ZN(n2502) );
  INV_X1 U32200 ( .A(n3888), .ZN(n3882) );
  NAND2_X1 U32210 ( .A1(n3898), .A2(n3882), .ZN(n2503) );
  INV_X1 U32220 ( .A(REG3_REG_26__SCAN_IN), .ZN(n4094) );
  AND2_X1 U32230 ( .A1(n2504), .A2(n4094), .ZN(n2505) );
  INV_X1 U32240 ( .A(REG2_REG_26__SCAN_IN), .ZN(n3873) );
  NAND2_X1 U32250 ( .A1(n3611), .A2(REG0_REG_26__SCAN_IN), .ZN(n2507) );
  NAND2_X1 U32260 ( .A1(n3610), .A2(REG1_REG_26__SCAN_IN), .ZN(n2506) );
  OAI211_X1 U32270 ( .C1(n3873), .C2(n2008), .A(n2507), .B(n2506), .ZN(n2508)
         );
  INV_X1 U32280 ( .A(n2508), .ZN(n2509) );
  INV_X1 U32290 ( .A(n3883), .ZN(n3852) );
  NAND2_X1 U32300 ( .A1(n2462), .A2(DATAI_26_), .ZN(n3872) );
  NOR2_X1 U32310 ( .A1(n3852), .A2(n3872), .ZN(n2510) );
  INV_X1 U32320 ( .A(n3872), .ZN(n2614) );
  OAI22_X2 U32330 ( .A1(n3861), .A2(n2510), .B1(n2614), .B2(n3883), .ZN(n3848)
         );
  INV_X1 U32340 ( .A(n3848), .ZN(n2517) );
  INV_X1 U32350 ( .A(REG3_REG_27__SCAN_IN), .ZN(n3466) );
  XNOR2_X1 U32360 ( .A(n2519), .B(n3466), .ZN(n3854) );
  NAND2_X1 U32370 ( .A1(n3854), .A2(n2282), .ZN(n2516) );
  INV_X1 U32380 ( .A(REG2_REG_27__SCAN_IN), .ZN(n2513) );
  NAND2_X1 U32390 ( .A1(n3611), .A2(REG0_REG_27__SCAN_IN), .ZN(n2512) );
  NAND2_X1 U32400 ( .A1(n3610), .A2(REG1_REG_27__SCAN_IN), .ZN(n2511) );
  OAI211_X1 U32410 ( .C1(n2513), .C2(n2008), .A(n2512), .B(n2511), .ZN(n2514)
         );
  INV_X1 U32420 ( .A(n2514), .ZN(n2515) );
  AND2_X1 U32430 ( .A1(REG3_REG_27__SCAN_IN), .A2(REG3_REG_28__SCAN_IN), .ZN(
        n2518) );
  AND2_X1 U32440 ( .A1(n2519), .A2(n2518), .ZN(n3835) );
  AOI21_X1 U32450 ( .B1(n2519), .B2(REG3_REG_27__SCAN_IN), .A(
        REG3_REG_28__SCAN_IN), .ZN(n2520) );
  INV_X1 U32460 ( .A(REG2_REG_28__SCAN_IN), .ZN(n3438) );
  NAND2_X1 U32470 ( .A1(n3611), .A2(REG0_REG_28__SCAN_IN), .ZN(n2522) );
  NAND2_X1 U32480 ( .A1(n3610), .A2(REG1_REG_28__SCAN_IN), .ZN(n2521) );
  OAI211_X1 U32490 ( .C1(n3438), .C2(n2008), .A(n2522), .B(n2521), .ZN(n2523)
         );
  INV_X1 U32500 ( .A(n2523), .ZN(n2524) );
  NAND2_X1 U32510 ( .A1(n2462), .A2(DATAI_28_), .ZN(n3836) );
  OR2_X1 U32520 ( .A1(n3423), .A2(n3836), .ZN(n3699) );
  NAND2_X1 U32530 ( .A1(n3423), .A2(n3836), .ZN(n3828) );
  XNOR2_X1 U32540 ( .A(n3838), .B(n3837), .ZN(n3447) );
  NAND2_X1 U32550 ( .A1(n2583), .A2(IR_REG_31__SCAN_IN), .ZN(n2530) );
  INV_X1 U32560 ( .A(n2583), .ZN(n2531) );
  NAND2_X1 U32570 ( .A1(n2531), .A2(n2240), .ZN(n2532) );
  XNOR2_X1 U32580 ( .A(n2728), .B(n3747), .ZN(n2534) );
  INV_X1 U32590 ( .A(n4334), .ZN(n3822) );
  NAND2_X1 U32600 ( .A1(n2534), .A2(n3822), .ZN(n3212) );
  AND2_X1 U32610 ( .A1(n2576), .A2(n4334), .ZN(n2535) );
  INV_X1 U32620 ( .A(n3836), .ZN(n3441) );
  NAND2_X1 U32630 ( .A1(n2536), .A2(n2597), .ZN(n3006) );
  INV_X1 U32640 ( .A(n2537), .ZN(n2539) );
  MUX2_X1 U32650 ( .A(n2537), .B(n2539), .S(n2538), .Z(n4341) );
  NAND2_X1 U32660 ( .A1(n3747), .A2(n3643), .ZN(n2742) );
  INV_X1 U32670 ( .A(n2742), .ZN(n2651) );
  INV_X1 U32680 ( .A(REG2_REG_29__SCAN_IN), .ZN(n3842) );
  NAND2_X1 U32690 ( .A1(n3610), .A2(REG1_REG_29__SCAN_IN), .ZN(n2541) );
  NAND2_X1 U32700 ( .A1(n3611), .A2(REG0_REG_29__SCAN_IN), .ZN(n2540) );
  OAI211_X1 U32710 ( .C1(n3842), .C2(n2008), .A(n2541), .B(n2540), .ZN(n2542)
         );
  AOI21_X1 U32720 ( .B1(n3835), .B2(n2006), .A(n2542), .ZN(n3702) );
  INV_X1 U32730 ( .A(n2879), .ZN(n2544) );
  NAND2_X1 U32740 ( .A1(n2544), .A2(n2733), .ZN(n3640) );
  NAND2_X1 U32750 ( .A1(n2878), .A2(n2545), .ZN(n2547) );
  NAND2_X1 U32760 ( .A1(n2547), .A2(n3596), .ZN(n2766) );
  NAND2_X1 U32770 ( .A1(n2766), .A2(n3644), .ZN(n2920) );
  NAND2_X1 U32780 ( .A1(n2548), .A2(n2926), .ZN(n3649) );
  NAND2_X1 U32790 ( .A1(n3761), .A2(n3485), .ZN(n3646) );
  NAND2_X1 U32800 ( .A1(n2920), .A2(n3595), .ZN(n2919) );
  NAND2_X1 U32810 ( .A1(n2919), .A2(n3649), .ZN(n2934) );
  INV_X1 U32820 ( .A(n3650), .ZN(n2549) );
  AND2_X1 U32830 ( .A1(n3759), .A2(n3000), .ZN(n2991) );
  NAND2_X1 U32840 ( .A1(n2913), .A2(n2993), .ZN(n3665) );
  NAND2_X1 U32850 ( .A1(n3758), .A2(n2187), .ZN(n3667) );
  NAND2_X1 U32860 ( .A1(n2188), .A2(n2979), .ZN(n3656) );
  NAND2_X1 U32870 ( .A1(n2550), .A2(n3656), .ZN(n2957) );
  INV_X1 U32880 ( .A(n2551), .ZN(n3658) );
  NAND2_X1 U32890 ( .A1(n2552), .A2(n3655), .ZN(n3076) );
  NAND2_X1 U32900 ( .A1(n3097), .A2(n2553), .ZN(n3660) );
  NAND2_X1 U32910 ( .A1(n3757), .A2(n3077), .ZN(n3668) );
  AND2_X1 U32920 ( .A1(n3756), .A2(n3053), .ZN(n3663) );
  NAND2_X1 U32930 ( .A1(n3116), .A2(n3100), .ZN(n3661) );
  NAND2_X1 U32940 ( .A1(n3154), .A2(n3142), .ZN(n3676) );
  NAND2_X1 U32950 ( .A1(n3139), .A2(n3676), .ZN(n2554) );
  NAND2_X1 U32960 ( .A1(n3181), .A2(n3118), .ZN(n3671) );
  NAND2_X1 U32970 ( .A1(n3754), .A2(n3257), .ZN(n3203) );
  NAND2_X1 U32980 ( .A1(n3753), .A2(n3267), .ZN(n2555) );
  NAND2_X1 U32990 ( .A1(n3203), .A2(n2555), .ZN(n3677) );
  INV_X1 U33000 ( .A(n3124), .ZN(n3679) );
  NOR2_X1 U33010 ( .A1(n3677), .A2(n3679), .ZN(n2556) );
  NAND2_X1 U33020 ( .A1(n3152), .A2(n2556), .ZN(n2560) );
  NAND2_X1 U33030 ( .A1(n3323), .A2(n3130), .ZN(n3205) );
  NAND2_X1 U33040 ( .A1(n3122), .A2(n3205), .ZN(n2559) );
  INV_X1 U33050 ( .A(n3677), .ZN(n2558) );
  NOR2_X1 U33060 ( .A1(n3753), .A2(n3267), .ZN(n2557) );
  AOI21_X1 U33070 ( .B1(n2559), .B2(n2558), .A(n2557), .ZN(n3639) );
  NAND2_X1 U33080 ( .A1(n2560), .A2(n3639), .ZN(n3719) );
  NAND2_X1 U33090 ( .A1(n3719), .A2(n2205), .ZN(n2561) );
  NAND2_X1 U33100 ( .A1(n4342), .A2(n4278), .ZN(n3636) );
  NAND2_X1 U33110 ( .A1(n4062), .A2(n3305), .ZN(n3635) );
  NAND2_X1 U33120 ( .A1(n3636), .A2(n3635), .ZN(n3306) );
  INV_X1 U33130 ( .A(n4048), .ZN(n4059) );
  NAND2_X1 U33140 ( .A1(n4345), .A2(n4042), .ZN(n3987) );
  NAND2_X1 U33150 ( .A1(n3989), .A2(n3987), .ZN(n2564) );
  NAND2_X1 U33160 ( .A1(n4016), .A2(n4002), .ZN(n2562) );
  AND2_X1 U33170 ( .A1(n3990), .A2(n2562), .ZN(n2566) );
  NOR2_X1 U33180 ( .A1(n4016), .A2(n4002), .ZN(n2563) );
  AOI21_X1 U33190 ( .B1(n2564), .B2(n2566), .A(n2563), .ZN(n3917) );
  NAND2_X1 U33200 ( .A1(n3995), .A2(n3609), .ZN(n3920) );
  NAND2_X1 U33210 ( .A1(n3917), .A2(n3920), .ZN(n2565) );
  NAND2_X1 U33220 ( .A1(n3966), .A2(n4256), .ZN(n3919) );
  NAND2_X1 U33230 ( .A1(n2565), .A2(n3919), .ZN(n3685) );
  NAND2_X1 U33240 ( .A1(n3974), .A2(n4250), .ZN(n3606) );
  AND2_X1 U33250 ( .A1(n3923), .A2(n3606), .ZN(n3691) );
  NAND2_X1 U33260 ( .A1(n3685), .A2(n3691), .ZN(n3725) );
  INV_X1 U33270 ( .A(n3725), .ZN(n2573) );
  INV_X1 U33280 ( .A(n2566), .ZN(n2567) );
  AND2_X1 U33290 ( .A1(n4063), .A2(n4038), .ZN(n3988) );
  NOR2_X1 U33300 ( .A1(n2567), .A2(n3988), .ZN(n3915) );
  AND2_X1 U33310 ( .A1(n3915), .A2(n3919), .ZN(n3687) );
  OR2_X1 U33320 ( .A1(n3725), .A2(n3687), .ZN(n2572) );
  NOR2_X1 U33330 ( .A1(n3974), .A2(n4250), .ZN(n3692) );
  AND2_X1 U33340 ( .A1(n3923), .A2(n3692), .ZN(n2570) );
  NAND2_X1 U33350 ( .A1(n3944), .A2(n3933), .ZN(n2569) );
  NAND2_X1 U33360 ( .A1(n2569), .A2(n2568), .ZN(n3689) );
  NOR2_X1 U33370 ( .A1(n2570), .A2(n3689), .ZN(n2571) );
  NAND2_X1 U33380 ( .A1(n2572), .A2(n2571), .ZN(n3723) );
  AOI21_X1 U33390 ( .B1(n4033), .B2(n2573), .A(n3723), .ZN(n3895) );
  NOR2_X1 U33400 ( .A1(n3928), .A2(n4236), .ZN(n3604) );
  NOR2_X1 U33410 ( .A1(n3944), .A2(n3933), .ZN(n3894) );
  NOR2_X1 U33420 ( .A1(n3604), .A2(n3894), .ZN(n3729) );
  INV_X1 U33430 ( .A(n3729), .ZN(n3695) );
  NAND2_X1 U33440 ( .A1(n3928), .A2(n4236), .ZN(n3603) );
  NOR2_X1 U33450 ( .A1(n3883), .A2(n3872), .ZN(n3602) );
  NOR2_X1 U33460 ( .A1(n3898), .A2(n3888), .ZN(n3862) );
  NOR2_X1 U33470 ( .A1(n3602), .A2(n3862), .ZN(n3727) );
  INV_X1 U33480 ( .A(n3727), .ZN(n2574) );
  NOR2_X1 U33490 ( .A1(n3575), .A2(n3855), .ZN(n3697) );
  INV_X1 U33500 ( .A(n3732), .ZN(n2575) );
  XOR2_X1 U33510 ( .A(n3837), .B(n3829), .Z(n2578) );
  NAND2_X1 U33520 ( .A1(n3747), .A2(n4334), .ZN(n2577) );
  INV_X1 U3353 ( .A(n2576), .ZN(n2617) );
  NAND2_X1 U33540 ( .A1(n2617), .A2(n3643), .ZN(n3738) );
  OAI222_X1 U3355 ( .A1(n3994), .A2(n3702), .B1(n4018), .B2(n3575), .C1(n2578), 
        .C2(n3998), .ZN(n3445) );
  NAND2_X1 U3356 ( .A1(n2595), .A2(n2596), .ZN(n2584) );
  OAI21_X1 U3357 ( .B1(IR_REG_23__SCAN_IN), .B2(IR_REG_24__SCAN_IN), .A(
        IR_REG_31__SCAN_IN), .ZN(n2587) );
  NAND2_X1 U3358 ( .A1(n2595), .A2(n2587), .ZN(n2588) );
  NAND2_X1 U3359 ( .A1(n2591), .A2(n2592), .ZN(n2589) );
  MUX2_X1 U3360 ( .A(n2591), .B(n2589), .S(B_REG_SCAN_IN), .Z(n2590) );
  INV_X1 U3361 ( .A(n2593), .ZN(n2612) );
  NAND2_X1 U3362 ( .A1(n2612), .A2(n2592), .ZN(n2647) );
  OAI21_X1 U3363 ( .B1(n2646), .B2(D_REG_1__SCAN_IN), .A(n2647), .ZN(n2611) );
  INV_X1 U3364 ( .A(n2591), .ZN(n2594) );
  XNOR2_X1 U3365 ( .A(n2595), .B(n2596), .ZN(n2843) );
  NAND2_X1 U3366 ( .A1(n4554), .A2(n2597), .ZN(n2752) );
  AND2_X1 U3367 ( .A1(n2576), .A2(n3822), .ZN(n2598) );
  OR2_X1 U3368 ( .A1(n2598), .A2(n2742), .ZN(n2871) );
  NAND2_X1 U3369 ( .A1(n2752), .A2(n2871), .ZN(n2599) );
  NOR2_X1 U3370 ( .A1(n2753), .A2(n2599), .ZN(n2610) );
  NOR2_X1 U3371 ( .A1(D_REG_26__SCAN_IN), .A2(D_REG_27__SCAN_IN), .ZN(n2602)
         );
  NOR4_X1 U3372 ( .A1(D_REG_19__SCAN_IN), .A2(D_REG_28__SCAN_IN), .A3(
        D_REG_6__SCAN_IN), .A4(D_REG_3__SCAN_IN), .ZN(n4221) );
  NOR4_X1 U3373 ( .A1(D_REG_2__SCAN_IN), .A2(D_REG_4__SCAN_IN), .A3(
        D_REG_7__SCAN_IN), .A4(D_REG_8__SCAN_IN), .ZN(n2601) );
  NOR4_X1 U3374 ( .A1(D_REG_10__SCAN_IN), .A2(D_REG_29__SCAN_IN), .A3(
        D_REG_30__SCAN_IN), .A4(D_REG_5__SCAN_IN), .ZN(n2600) );
  AND4_X1 U3375 ( .A1(n2602), .A2(n4221), .A3(n2601), .A4(n2600), .ZN(n2608)
         );
  NOR4_X1 U3376 ( .A1(D_REG_14__SCAN_IN), .A2(D_REG_15__SCAN_IN), .A3(
        D_REG_16__SCAN_IN), .A4(D_REG_17__SCAN_IN), .ZN(n2606) );
  NOR4_X1 U3377 ( .A1(D_REG_12__SCAN_IN), .A2(D_REG_9__SCAN_IN), .A3(
        D_REG_11__SCAN_IN), .A4(D_REG_13__SCAN_IN), .ZN(n2605) );
  NOR4_X1 U3378 ( .A1(D_REG_23__SCAN_IN), .A2(D_REG_24__SCAN_IN), .A3(
        D_REG_25__SCAN_IN), .A4(D_REG_31__SCAN_IN), .ZN(n2604) );
  NOR4_X1 U3379 ( .A1(D_REG_18__SCAN_IN), .A2(D_REG_20__SCAN_IN), .A3(
        D_REG_21__SCAN_IN), .A4(D_REG_22__SCAN_IN), .ZN(n2603) );
  AND4_X1 U3380 ( .A1(n2606), .A2(n2605), .A3(n2604), .A4(n2603), .ZN(n2607)
         );
  NAND2_X1 U3381 ( .A1(n2608), .A2(n2607), .ZN(n2736) );
  NAND2_X1 U3382 ( .A1(n2740), .A2(n2736), .ZN(n2609) );
  INV_X1 U3383 ( .A(D_REG_0__SCAN_IN), .ZN(n3454) );
  AND2_X1 U3384 ( .A1(n2612), .A2(n2591), .ZN(n2613) );
  INV_X1 U3385 ( .A(n3947), .ZN(n3953) );
  INV_X1 U3386 ( .A(n3855), .ZN(n4087) );
  NOR2_X1 U3387 ( .A1(n2615), .A2(n3836), .ZN(n2616) );
  NAND2_X1 U3388 ( .A1(n2618), .A2(n2224), .ZN(U3546) );
  INV_X1 U3389 ( .A(n2741), .ZN(n2874) );
  INV_X1 U3390 ( .A(n2621), .ZN(n2622) );
  NAND2_X1 U3391 ( .A1(n2622), .A2(n2223), .ZN(U3514) );
  INV_X1 U3392 ( .A(n4518), .ZN(n3452) );
  INV_X2 U3393 ( .A(U4043), .ZN(n3762) );
  INV_X2 U3394 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  MUX2_X1 U3395 ( .A(n2714), .B(n2317), .S(U3149), .Z(n2623) );
  INV_X1 U3396 ( .A(n2623), .ZN(U3347) );
  INV_X1 U3397 ( .A(n3244), .ZN(n3809) );
  NAND2_X1 U3398 ( .A1(n3809), .A2(STATE_REG_SCAN_IN), .ZN(n2624) );
  OAI21_X1 U3399 ( .B1(STATE_REG_SCAN_IN), .B2(n2275), .A(n2624), .ZN(U3339)
         );
  INV_X1 U3400 ( .A(DATAI_27_), .ZN(n4184) );
  INV_X1 U3401 ( .A(IR_REG_27__SCAN_IN), .ZN(n2625) );
  INV_X1 U3402 ( .A(n3832), .ZN(n2649) );
  NAND2_X1 U3403 ( .A1(n2649), .A2(STATE_REG_SCAN_IN), .ZN(n2626) );
  OAI21_X1 U3404 ( .B1(STATE_REG_SCAN_IN), .B2(n4184), .A(n2626), .ZN(U3325)
         );
  INV_X1 U3405 ( .A(DATAI_29_), .ZN(n2629) );
  NAND2_X1 U3406 ( .A1(n2627), .A2(STATE_REG_SCAN_IN), .ZN(n2628) );
  OAI21_X1 U3407 ( .B1(STATE_REG_SCAN_IN), .B2(n2629), .A(n2628), .ZN(U3323)
         );
  INV_X1 U3408 ( .A(DATAI_30_), .ZN(n2632) );
  NAND2_X1 U3409 ( .A1(n2630), .A2(STATE_REG_SCAN_IN), .ZN(n2631) );
  OAI21_X1 U3410 ( .B1(STATE_REG_SCAN_IN), .B2(n2632), .A(n2631), .ZN(U3322)
         );
  INV_X1 U3411 ( .A(DATAI_21_), .ZN(n2634) );
  NAND2_X1 U3412 ( .A1(n3643), .A2(STATE_REG_SCAN_IN), .ZN(n2633) );
  OAI21_X1 U3413 ( .B1(STATE_REG_SCAN_IN), .B2(n2634), .A(n2633), .ZN(U3331)
         );
  INV_X1 U3414 ( .A(DATAI_26_), .ZN(n2636) );
  NAND2_X1 U3415 ( .A1(n2593), .A2(STATE_REG_SCAN_IN), .ZN(n2635) );
  OAI21_X1 U3416 ( .B1(STATE_REG_SCAN_IN), .B2(n2636), .A(n2635), .ZN(U3326)
         );
  INV_X1 U3417 ( .A(DATAI_20_), .ZN(n2638) );
  NAND2_X1 U3418 ( .A1(n2617), .A2(STATE_REG_SCAN_IN), .ZN(n2637) );
  OAI21_X1 U3419 ( .B1(STATE_REG_SCAN_IN), .B2(n2638), .A(n2637), .ZN(U3332)
         );
  INV_X1 U3420 ( .A(DATAI_22_), .ZN(n2640) );
  NAND2_X1 U3421 ( .A1(n3747), .A2(STATE_REG_SCAN_IN), .ZN(n2639) );
  OAI21_X1 U3422 ( .B1(STATE_REG_SCAN_IN), .B2(n2640), .A(n2639), .ZN(U3330)
         );
  INV_X1 U3423 ( .A(DATAI_25_), .ZN(n2643) );
  NAND2_X1 U3424 ( .A1(n2641), .A2(STATE_REG_SCAN_IN), .ZN(n2642) );
  OAI21_X1 U3425 ( .B1(STATE_REG_SCAN_IN), .B2(n2643), .A(n2642), .ZN(U3327)
         );
  INV_X1 U3426 ( .A(DATAI_24_), .ZN(n2644) );
  MUX2_X1 U3427 ( .A(n2591), .B(n2644), .S(U3149), .Z(n2645) );
  INV_X1 U3428 ( .A(n2645), .ZN(U3328) );
  INV_X1 U3429 ( .A(D_REG_1__SCAN_IN), .ZN(n2648) );
  INV_X1 U3430 ( .A(n2647), .ZN(n2738) );
  AOI22_X1 U3431 ( .A1(n4517), .A2(n2648), .B1(n2738), .B2(n4518), .ZN(U3459)
         );
  AOI21_X1 U3432 ( .B1(n2649), .B2(n3011), .A(n4341), .ZN(n3777) );
  OAI21_X1 U3433 ( .B1(REG1_REG_0__SCAN_IN), .B2(n2649), .A(n3777), .ZN(n2650)
         );
  MUX2_X1 U3434 ( .A(n2650), .B(n3777), .S(IR_REG_0__SCAN_IN), .Z(n2661) );
  NAND2_X1 U3435 ( .A1(n2651), .A2(n2843), .ZN(n2652) );
  AND2_X1 U3436 ( .A1(n2462), .A2(n2652), .ZN(n2654) );
  INV_X1 U3437 ( .A(n2843), .ZN(n2653) );
  NAND2_X1 U3438 ( .A1(n2653), .A2(STATE_REG_SCAN_IN), .ZN(n3749) );
  NAND2_X1 U3439 ( .A1(n2753), .A2(n3749), .ZN(n2655) );
  INV_X1 U3440 ( .A(n2667), .ZN(n2660) );
  INV_X1 U3441 ( .A(n2654), .ZN(n2656) );
  AOI22_X1 U3442 ( .A1(n4462), .A2(ADDR_REG_0__SCAN_IN), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n2659) );
  INV_X1 U3443 ( .A(REG1_REG_0__SCAN_IN), .ZN(n2657) );
  NAND3_X1 U3444 ( .A1(n4470), .A2(IR_REG_0__SCAN_IN), .A3(n2657), .ZN(n2658)
         );
  OAI211_X1 U3445 ( .C1(n2661), .C2(n2660), .A(n2659), .B(n2658), .ZN(U3240)
         );
  AOI222_X1 U3446 ( .A1(n2004), .A2(REG2_REG_30__SCAN_IN), .B1(n2022), .B2(
        REG1_REG_30__SCAN_IN), .C1(n3611), .C2(REG0_REG_30__SCAN_IN), .ZN(
        n3833) );
  NAND2_X1 U3447 ( .A1(n3762), .A2(DATAO_REG_30__SCAN_IN), .ZN(n2662) );
  OAI21_X1 U3448 ( .B1(n3833), .B2(n3762), .A(n2662), .ZN(U3580) );
  INV_X1 U3449 ( .A(REG1_REG_2__SCAN_IN), .ZN(n3785) );
  MUX2_X1 U3450 ( .A(REG1_REG_2__SCAN_IN), .B(n3785), .S(n4338), .Z(n2665) );
  INV_X1 U3451 ( .A(REG1_REG_1__SCAN_IN), .ZN(n2663) );
  AND2_X1 U3452 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n3765)
         );
  NAND2_X1 U3453 ( .A1(n4339), .A2(REG1_REG_1__SCAN_IN), .ZN(n3786) );
  NAND2_X1 U3454 ( .A1(n3787), .A2(n3786), .ZN(n2664) );
  NAND2_X1 U3455 ( .A1(n4338), .A2(REG1_REG_2__SCAN_IN), .ZN(n2666) );
  NAND2_X1 U3456 ( .A1(n3790), .A2(n2666), .ZN(n2691) );
  XNOR2_X1 U3457 ( .A(n2691), .B(n2676), .ZN(n2690) );
  XOR2_X1 U34580 ( .A(n2690), .B(REG1_REG_3__SCAN_IN), .Z(n2673) );
  NOR2_X1 U34590 ( .A1(n4341), .A2(n3832), .ZN(n3745) );
  MUX2_X1 U3460 ( .A(REG2_REG_2__SCAN_IN), .B(n2668), .S(n4338), .Z(n2670) );
  MUX2_X1 U3461 ( .A(REG2_REG_1__SCAN_IN), .B(n2276), .S(n4339), .Z(n3766) );
  AND2_X1 U3462 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n3774)
         );
  NAND2_X1 U3463 ( .A1(n3766), .A2(n3774), .ZN(n3779) );
  NAND2_X1 U3464 ( .A1(n4339), .A2(REG2_REG_1__SCAN_IN), .ZN(n3778) );
  NAND2_X1 U3465 ( .A1(n3779), .A2(n3778), .ZN(n2669) );
  NAND2_X1 U3466 ( .A1(n2670), .A2(n2669), .ZN(n3781) );
  NAND2_X1 U34670 ( .A1(n4338), .A2(REG2_REG_2__SCAN_IN), .ZN(n2671) );
  NAND2_X1 U3468 ( .A1(n3781), .A2(n2671), .ZN(n2678) );
  XNOR2_X1 U34690 ( .A(n2678), .B(n2676), .ZN(n2677) );
  XNOR2_X1 U3470 ( .A(n2677), .B(n2927), .ZN(n2672) );
  AOI22_X1 U34710 ( .A1(n4470), .A2(n2673), .B1(n4472), .B2(n2672), .ZN(n2675)
         );
  AOI22_X1 U3472 ( .A1(n4462), .A2(ADDR_REG_3__SCAN_IN), .B1(
        REG3_REG_3__SCAN_IN), .B2(U3149), .ZN(n2674) );
  OAI211_X1 U34730 ( .C1(n2676), .C2(n4475), .A(n2675), .B(n2674), .ZN(U3243)
         );
  INV_X1 U3474 ( .A(n3762), .ZN(n3775) );
  NOR2_X1 U34750 ( .A1(n4462), .A2(n3775), .ZN(U3148) );
  INV_X1 U3476 ( .A(n4462), .ZN(n4488) );
  INV_X1 U34770 ( .A(ADDR_REG_7__SCAN_IN), .ZN(n4101) );
  NAND2_X1 U3478 ( .A1(REG3_REG_7__SCAN_IN), .A2(U3149), .ZN(n3062) );
  NAND2_X1 U34790 ( .A1(n2677), .A2(REG2_REG_3__SCAN_IN), .ZN(n2680) );
  NAND2_X1 U3480 ( .A1(n2678), .A2(n4337), .ZN(n2679) );
  NAND2_X1 U34810 ( .A1(n2680), .A2(n2679), .ZN(n2681) );
  XNOR2_X1 U3482 ( .A(n2681), .B(n4377), .ZN(n4372) );
  MUX2_X1 U34830 ( .A(REG2_REG_5__SCAN_IN), .B(n2683), .S(n2714), .Z(n2709) );
  OAI21_X1 U3484 ( .B1(n2683), .B2(n2714), .A(n2682), .ZN(n2684) );
  NAND2_X1 U34850 ( .A1(n2697), .A2(n2684), .ZN(n2685) );
  XOR2_X1 U3486 ( .A(n2684), .B(n2697), .Z(n4387) );
  NAND2_X1 U34870 ( .A1(REG2_REG_6__SCAN_IN), .A2(n4387), .ZN(n4386) );
  NAND2_X1 U3488 ( .A1(n2685), .A2(n4386), .ZN(n2688) );
  MUX2_X1 U34890 ( .A(REG2_REG_7__SCAN_IN), .B(n2686), .S(n4336), .Z(n2687) );
  NAND2_X1 U3490 ( .A1(n2688), .A2(n2687), .ZN(n2796) );
  OAI211_X1 U34910 ( .C1(n2688), .C2(n2687), .A(n2796), .B(n4472), .ZN(n2689)
         );
  OAI211_X1 U3492 ( .C1(n4488), .C2(n4101), .A(n3062), .B(n2689), .ZN(n2702)
         );
  NAND2_X1 U34930 ( .A1(n4336), .A2(REG1_REG_7__SCAN_IN), .ZN(n2803) );
  OAI21_X1 U3494 ( .B1(n4336), .B2(REG1_REG_7__SCAN_IN), .A(n2803), .ZN(n2699)
         );
  INV_X1 U34950 ( .A(n2714), .ZN(n2696) );
  NAND2_X1 U3496 ( .A1(n2690), .A2(REG1_REG_3__SCAN_IN), .ZN(n2693) );
  NAND2_X1 U34970 ( .A1(n2691), .A2(n4337), .ZN(n2692) );
  NAND2_X1 U3498 ( .A1(n2693), .A2(n2692), .ZN(n2695) );
  INV_X1 U34990 ( .A(n4377), .ZN(n2694) );
  XNOR2_X1 U3500 ( .A(n2695), .B(n2694), .ZN(n4375) );
  AOI22_X1 U35010 ( .A1(n4375), .A2(REG1_REG_4__SCAN_IN), .B1(n4377), .B2(
        n2695), .ZN(n2712) );
  INV_X1 U3502 ( .A(REG1_REG_5__SCAN_IN), .ZN(n4582) );
  MUX2_X1 U35030 ( .A(REG1_REG_5__SCAN_IN), .B(n4582), .S(n2714), .Z(n2711) );
  NOR2_X1 U3504 ( .A1(n2712), .A2(n2711), .ZN(n2710) );
  INV_X1 U35050 ( .A(n2697), .ZN(n4536) );
  XNOR2_X1 U35060 ( .A(n2698), .B(n2697), .ZN(n4385) );
  NAND2_X1 U35070 ( .A1(REG1_REG_6__SCAN_IN), .A2(n4385), .ZN(n4384) );
  OAI21_X1 U35080 ( .B1(n2698), .B2(n4536), .A(n4384), .ZN(n2805) );
  XOR2_X1 U35090 ( .A(n2699), .B(n2805), .Z(n2700) );
  INV_X1 U35100 ( .A(n4336), .ZN(n2797) );
  OAI22_X1 U35110 ( .A1(n2700), .A2(n4476), .B1(n4475), .B2(n2797), .ZN(n2701)
         );
  OR2_X1 U35120 ( .A1(n2702), .A2(n2701), .ZN(U3247) );
  INV_X1 U35130 ( .A(DATAO_REG_10__SCAN_IN), .ZN(n4106) );
  NAND2_X1 U35140 ( .A1(n3154), .A2(U4043), .ZN(n2703) );
  OAI21_X1 U35150 ( .B1(n3775), .B2(n4106), .A(n2703), .ZN(U3560) );
  INV_X1 U35160 ( .A(DATAO_REG_14__SCAN_IN), .ZN(n2705) );
  NAND2_X1 U35170 ( .A1(n3283), .A2(U4043), .ZN(n2704) );
  OAI21_X1 U35180 ( .B1(n3775), .B2(n2705), .A(n2704), .ZN(U3564) );
  INV_X1 U35190 ( .A(DATAO_REG_15__SCAN_IN), .ZN(n2707) );
  NAND2_X1 U35200 ( .A1(n4062), .A2(n3775), .ZN(n2706) );
  OAI21_X1 U35210 ( .B1(n3775), .B2(n2707), .A(n2706), .ZN(U3565) );
  INV_X1 U35220 ( .A(n4472), .ZN(n4479) );
  AOI211_X1 U35230 ( .C1(n2021), .C2(n2709), .A(n2708), .B(n4479), .ZN(n2717)
         );
  AOI211_X1 U35240 ( .C1(n2712), .C2(n2711), .A(n2710), .B(n4476), .ZN(n2716)
         );
  AND2_X1 U35250 ( .A1(U3149), .A2(REG3_REG_5__SCAN_IN), .ZN(n2866) );
  AOI21_X1 U35260 ( .B1(n4462), .B2(ADDR_REG_5__SCAN_IN), .A(n2866), .ZN(n2713) );
  OAI21_X1 U35270 ( .B1(n4475), .B2(n2714), .A(n2713), .ZN(n2715) );
  OR3_X1 U35280 ( .A1(n2717), .A2(n2716), .A3(n2715), .ZN(U3245) );
  INV_X1 U35290 ( .A(DATAO_REG_7__SCAN_IN), .ZN(n2719) );
  NAND2_X1 U35300 ( .A1(n3046), .A2(U4043), .ZN(n2718) );
  OAI21_X1 U35310 ( .B1(U4043), .B2(n2719), .A(n2718), .ZN(U3557) );
  INV_X1 U35320 ( .A(DATAO_REG_0__SCAN_IN), .ZN(n2721) );
  NAND2_X1 U35330 ( .A1(n2879), .A2(U4043), .ZN(n2720) );
  OAI21_X1 U35340 ( .B1(U4043), .B2(n2721), .A(n2720), .ZN(U3550) );
  INV_X1 U35350 ( .A(DATAO_REG_20__SCAN_IN), .ZN(n4099) );
  NAND2_X1 U35360 ( .A1(n3966), .A2(U4043), .ZN(n2722) );
  OAI21_X1 U35370 ( .B1(n3775), .B2(n4099), .A(n2722), .ZN(U3570) );
  NAND2_X1 U35380 ( .A1(n2879), .A2(n3015), .ZN(n3642) );
  AND2_X1 U35390 ( .A1(n3640), .A2(n3642), .ZN(n3625) );
  INV_X1 U35400 ( .A(n3212), .ZN(n3137) );
  NOR2_X1 U35410 ( .A1(n3137), .A2(n4057), .ZN(n2723) );
  OAI22_X1 U35420 ( .A1(n3625), .A2(n2723), .B1(n2755), .B2(n3994), .ZN(n3009)
         );
  OAI22_X1 U35430 ( .A1(n3625), .A2(n4545), .B1(n3015), .B2(n3006), .ZN(n2724)
         );
  NOR2_X1 U35440 ( .A1(n3009), .A2(n2724), .ZN(n4539) );
  NAND2_X1 U35450 ( .A1(n4586), .A2(REG1_REG_0__SCAN_IN), .ZN(n2725) );
  OAI21_X1 U35460 ( .B1(n4539), .B2(n4586), .A(n2725), .ZN(U3518) );
  INV_X1 U35470 ( .A(n2728), .ZN(n2726) );
  INV_X1 U35480 ( .A(n2727), .ZN(n2730) );
  NAND2_X1 U35490 ( .A1(n2730), .A2(REG1_REG_0__SCAN_IN), .ZN(n2731) );
  NAND2_X1 U35500 ( .A1(n2783), .A2(n2731), .ZN(n2780) );
  NOR2_X1 U35510 ( .A1(n2727), .A2(n2132), .ZN(n2732) );
  AOI21_X1 U35520 ( .B1(n2733), .B2(n2007), .A(n2732), .ZN(n2735) );
  NAND2_X1 U35530 ( .A1(n2879), .A2(n3353), .ZN(n2734) );
  NAND2_X1 U35540 ( .A1(n2735), .A2(n2734), .ZN(n2779) );
  XOR2_X1 U35550 ( .A(n2780), .B(n2779), .Z(n3771) );
  INV_X1 U35560 ( .A(n3771), .ZN(n2758) );
  INV_X1 U35570 ( .A(n2736), .ZN(n2737) );
  NAND2_X1 U35580 ( .A1(n2737), .A2(D_REG_1__SCAN_IN), .ZN(n2739) );
  AOI21_X1 U35590 ( .B1(n2740), .B2(n2739), .A(n2738), .ZN(n2872) );
  NAND2_X1 U35600 ( .A1(n2872), .A2(n2741), .ZN(n2751) );
  OAI211_X1 U35610 ( .C1(n3006), .C2(n3822), .A(n4284), .B(n2742), .ZN(n2744)
         );
  OR2_X1 U35620 ( .A1(n2753), .A2(n2744), .ZN(n2743) );
  NAND2_X1 U35630 ( .A1(n2744), .A2(n4284), .ZN(n2745) );
  NAND2_X1 U35640 ( .A1(n2751), .A2(n2745), .ZN(n2746) );
  NAND2_X1 U35650 ( .A1(n2746), .A2(n2871), .ZN(n2845) );
  INV_X1 U35660 ( .A(n2845), .ZN(n2748) );
  AND2_X1 U35670 ( .A1(n4518), .A2(n2781), .ZN(n2747) );
  NAND2_X1 U35680 ( .A1(n2751), .A2(n3744), .ZN(n2846) );
  NAND3_X1 U35690 ( .A1(n2748), .A2(n2873), .A3(n2846), .ZN(n3460) );
  INV_X1 U35700 ( .A(n3744), .ZN(n2749) );
  NOR2_X1 U35710 ( .A1(n2751), .A2(n2749), .ZN(n2791) );
  NAND2_X1 U35720 ( .A1(n2873), .A2(n4277), .ZN(n2750) );
  OR2_X1 U35730 ( .A1(n2751), .A2(n2750), .ZN(n2754) );
  OAI22_X1 U35740 ( .A1(n4344), .A2(n2755), .B1(n4349), .B2(n3015), .ZN(n2756)
         );
  AOI21_X1 U35750 ( .B1(REG3_REG_0__SCAN_IN), .B2(n3460), .A(n2756), .ZN(n2757) );
  OAI21_X1 U35760 ( .B1(n2758), .B2(n3581), .A(n2757), .ZN(U3229) );
  NAND2_X1 U35770 ( .A1(n2760), .A2(n2761), .ZN(n2762) );
  NAND2_X1 U35780 ( .A1(n2762), .A2(n3596), .ZN(n2763) );
  NAND2_X1 U35790 ( .A1(n2759), .A2(n2763), .ZN(n2771) );
  INV_X1 U35800 ( .A(n2771), .ZN(n2951) );
  OAI22_X1 U35810 ( .A1(n2951), .A2(n4545), .B1(n2764), .B2(n4284), .ZN(n2774)
         );
  NAND3_X1 U3582 ( .A1(n2546), .A2(n2545), .A3(n2878), .ZN(n2765) );
  NAND2_X1 U3583 ( .A1(n2766), .A2(n2765), .ZN(n2770) );
  NAND2_X1 U3584 ( .A1(n3763), .A2(n4061), .ZN(n2768) );
  NAND2_X1 U3585 ( .A1(n3761), .A2(n4064), .ZN(n2767) );
  NAND2_X1 U3586 ( .A1(n2768), .A2(n2767), .ZN(n2769) );
  AOI21_X1 U3587 ( .B1(n2770), .B2(n4057), .A(n2769), .ZN(n2773) );
  NAND2_X1 U3588 ( .A1(n2771), .A2(n3137), .ZN(n2772) );
  NAND2_X1 U3589 ( .A1(n2773), .A2(n2772), .ZN(n2952) );
  NOR2_X1 U3590 ( .A1(n2774), .A2(n2952), .ZN(n2778) );
  INV_X1 U3591 ( .A(n4332), .ZN(n2982) );
  NAND2_X1 U3592 ( .A1(n2876), .A2(n3459), .ZN(n2775) );
  AND2_X1 U3593 ( .A1(n2925), .A2(n2775), .ZN(n2955) );
  AOI22_X1 U3594 ( .A1(n2982), .A2(n2955), .B1(REG0_REG_2__SCAN_IN), .B2(n4575), .ZN(n2776) );
  OAI21_X1 U3595 ( .B1(n2778), .B2(n4575), .A(n2776), .ZN(U3471) );
  INV_X1 U3596 ( .A(n4289), .ZN(n2987) );
  AOI22_X1 U3597 ( .A1(n2987), .A2(n2955), .B1(n4586), .B2(REG1_REG_2__SCAN_IN), .ZN(n2777) );
  OAI21_X1 U3598 ( .B1(n2778), .B2(n4586), .A(n2777), .ZN(U3520) );
  NAND2_X1 U3599 ( .A1(n2780), .A2(n2779), .ZN(n2785) );
  INV_X1 U3600 ( .A(n2781), .ZN(n2782) );
  NAND2_X1 U3601 ( .A1(n2783), .A2(n2860), .ZN(n2784) );
  NAND2_X1 U3602 ( .A1(n2785), .A2(n2784), .ZN(n2814) );
  NAND2_X1 U3603 ( .A1(n2007), .A2(n3763), .ZN(n2787) );
  NAND2_X1 U3604 ( .A1(n2790), .A2(n2829), .ZN(n2786) );
  XNOR2_X1 U3605 ( .A(n2814), .B(n2815), .ZN(n2794) );
  INV_X1 U3606 ( .A(n4344), .ZN(n3475) );
  AOI22_X1 U3607 ( .A1(n3475), .A2(n2789), .B1(n3589), .B2(n2790), .ZN(n2793)
         );
  INV_X1 U3608 ( .A(n4341), .ZN(n3772) );
  INV_X1 U3609 ( .A(n4343), .ZN(n3476) );
  AOI22_X1 U3610 ( .A1(REG3_REG_1__SCAN_IN), .A2(n3460), .B1(n3476), .B2(n2879), .ZN(n2792) );
  OAI211_X1 U3611 ( .C1(n2794), .C2(n3581), .A(n2793), .B(n2792), .ZN(U3219)
         );
  NAND2_X1 U3612 ( .A1(n3762), .A2(DATAO_REG_29__SCAN_IN), .ZN(n2795) );
  OAI21_X1 U3613 ( .B1(n3702), .B2(n3762), .A(n2795), .ZN(U3579) );
  INV_X1 U3614 ( .A(n4335), .ZN(n3221) );
  OAI21_X1 U3615 ( .B1(n2686), .B2(n2797), .A(n2796), .ZN(n2799) );
  INV_X1 U3616 ( .A(n4534), .ZN(n2798) );
  NAND2_X1 U3617 ( .A1(n2799), .A2(n2798), .ZN(n2800) );
  XNOR2_X1 U3618 ( .A(n2799), .B(n4534), .ZN(n4399) );
  NAND2_X1 U3619 ( .A1(REG2_REG_8__SCAN_IN), .A2(n4399), .ZN(n4398) );
  NAND2_X1 U3620 ( .A1(n2800), .A2(n4398), .ZN(n2802) );
  MUX2_X1 U3621 ( .A(REG2_REG_9__SCAN_IN), .B(n3058), .S(n4335), .Z(n2801) );
  NAND2_X1 U3622 ( .A1(n2802), .A2(n2801), .ZN(n3220) );
  OAI211_X1 U3623 ( .C1(n2802), .C2(n2801), .A(n3220), .B(n4472), .ZN(n2813)
         );
  AND2_X1 U3624 ( .A1(U3149), .A2(REG3_REG_9__SCAN_IN), .ZN(n3099) );
  INV_X1 U3625 ( .A(REG1_REG_8__SCAN_IN), .ZN(n4394) );
  INV_X1 U3626 ( .A(n2803), .ZN(n2804) );
  NAND2_X1 U3627 ( .A1(n2806), .A2(n4534), .ZN(n2807) );
  INV_X1 U3628 ( .A(REG1_REG_9__SCAN_IN), .ZN(n2808) );
  MUX2_X1 U3629 ( .A(n2808), .B(REG1_REG_9__SCAN_IN), .S(n4335), .Z(n2809) );
  NOR2_X1 U3630 ( .A1(n2810), .A2(n2809), .ZN(n3232) );
  AOI211_X1 U3631 ( .C1(n2810), .C2(n2809), .A(n3232), .B(n4476), .ZN(n2811)
         );
  AOI211_X1 U3632 ( .C1(n4462), .C2(ADDR_REG_9__SCAN_IN), .A(n3099), .B(n2811), 
        .ZN(n2812) );
  OAI211_X1 U3633 ( .C1(n4475), .C2(n3221), .A(n2813), .B(n2812), .ZN(U3249)
         );
  NAND2_X1 U3634 ( .A1(n2815), .A2(n2814), .ZN(n2820) );
  INV_X1 U3635 ( .A(n2816), .ZN(n2817) );
  NAND2_X1 U3636 ( .A1(n2818), .A2(n2817), .ZN(n2819) );
  NAND2_X1 U3637 ( .A1(n2820), .A2(n2819), .ZN(n3455) );
  INV_X1 U3638 ( .A(n3455), .ZN(n2827) );
  AOI22_X1 U3639 ( .A1(n2789), .A2(n3353), .B1(n3459), .B2(n2007), .ZN(n2825)
         );
  NAND2_X1 U3640 ( .A1(n2007), .A2(n2789), .ZN(n2822) );
  NAND2_X1 U3641 ( .A1(n3459), .A2(n2829), .ZN(n2821) );
  NAND2_X1 U3642 ( .A1(n2824), .A2(n2825), .ZN(n2828) );
  OAI21_X1 U3643 ( .B1(n2825), .B2(n2824), .A(n2828), .ZN(n3458) );
  INV_X1 U3644 ( .A(n3458), .ZN(n2826) );
  NAND2_X1 U3645 ( .A1(n2827), .A2(n2826), .ZN(n3456) );
  NAND2_X1 U3646 ( .A1(n3456), .A2(n2828), .ZN(n3482) );
  NAND2_X1 U3647 ( .A1(n3761), .A2(n2007), .ZN(n2831) );
  NAND2_X1 U3648 ( .A1(n2926), .A2(n2829), .ZN(n2830) );
  NAND2_X1 U3649 ( .A1(n2831), .A2(n2830), .ZN(n2832) );
  AOI22_X1 U3650 ( .A1(n3761), .A2(n3353), .B1(n2926), .B2(n2007), .ZN(n2837)
         );
  XNOR2_X1 U3651 ( .A(n2836), .B(n2837), .ZN(n3483) );
  NAND2_X1 U3652 ( .A1(n3760), .A2(n2007), .ZN(n2834) );
  NAND2_X1 U3653 ( .A1(n2938), .A2(n2829), .ZN(n2833) );
  NAND2_X1 U3654 ( .A1(n2834), .A2(n2833), .ZN(n2835) );
  XNOR2_X1 U3655 ( .A(n2835), .B(n3425), .ZN(n2853) );
  AOI22_X1 U3656 ( .A1(n3760), .A2(n3353), .B1(n2938), .B2(n2007), .ZN(n2854)
         );
  XNOR2_X1 U3657 ( .A(n2853), .B(n2854), .ZN(n2841) );
  INV_X1 U3658 ( .A(n2836), .ZN(n2838) );
  NAND2_X1 U3659 ( .A1(n2838), .A2(n2837), .ZN(n2842) );
  AND2_X1 U3660 ( .A1(n2841), .A2(n2842), .ZN(n2839) );
  NAND2_X1 U3661 ( .A1(n2857), .A2(n4357), .ZN(n2852) );
  AOI21_X1 U3662 ( .B1(n2840), .B2(n2842), .A(n2841), .ZN(n2851) );
  NAND2_X1 U3663 ( .A1(n2727), .A2(n2843), .ZN(n2844) );
  OAI21_X1 U3664 ( .B1(n2845), .B2(n2844), .A(STATE_REG_SCAN_IN), .ZN(n2847)
         );
  AOI22_X1 U3665 ( .A1(n3475), .A2(n3759), .B1(n3476), .B2(n3761), .ZN(n2848)
         );
  NAND2_X1 U3666 ( .A1(U3149), .A2(REG3_REG_4__SCAN_IN), .ZN(n4370) );
  OAI211_X1 U3667 ( .C1(n4349), .C2(n2931), .A(n2848), .B(n4370), .ZN(n2849)
         );
  AOI21_X1 U3668 ( .B1(n2945), .B2(n3578), .A(n2849), .ZN(n2850) );
  OAI21_X1 U3669 ( .B1(n2852), .B2(n2851), .A(n2850), .ZN(U3227) );
  NAND2_X1 U3670 ( .A1(n2853), .A2(n2855), .ZN(n2856) );
  NAND2_X1 U3671 ( .A1(n3759), .A2(n2007), .ZN(n2859) );
  OR2_X1 U3672 ( .A1(n3000), .A2(n3427), .ZN(n2858) );
  NAND2_X1 U3673 ( .A1(n2859), .A2(n2858), .ZN(n2861) );
  XNOR2_X1 U3674 ( .A(n2861), .B(n2860), .ZN(n2896) );
  NAND2_X1 U3675 ( .A1(n3759), .A2(n3353), .ZN(n2864) );
  OR2_X1 U3676 ( .A1(n3000), .A2(n2862), .ZN(n2863) );
  NAND2_X1 U3677 ( .A1(n2864), .A2(n2863), .ZN(n2897) );
  XNOR2_X1 U3678 ( .A(n2896), .B(n2897), .ZN(n2894) );
  XNOR2_X1 U3679 ( .A(n2895), .B(n2894), .ZN(n2870) );
  OAI22_X1 U3680 ( .A1(n3486), .A2(n4343), .B1(n4344), .B2(n2188), .ZN(n2865)
         );
  AOI211_X1 U3681 ( .C1(n2993), .C2(n3589), .A(n2866), .B(n2865), .ZN(n2869)
         );
  NAND2_X1 U3682 ( .A1(n3578), .A2(n2867), .ZN(n2868) );
  OAI211_X1 U3683 ( .C1(n2870), .C2(n3581), .A(n2869), .B(n2868), .ZN(U3224)
         );
  NAND4_X1 U3684 ( .A1(n2874), .A2(n2873), .A3(n2872), .A4(n2871), .ZN(n2875)
         );
  OR2_X1 U3685 ( .A1(n4507), .A2(n4334), .ZN(n4025) );
  NOR2_X2 U3686 ( .A1(n4025), .A2(n4559), .ZN(n4501) );
  OAI21_X1 U3687 ( .B1(n3015), .B2(n2882), .A(n2876), .ZN(n4540) );
  NAND2_X1 U3688 ( .A1(n2878), .A2(n2877), .ZN(n2884) );
  NAND2_X1 U3689 ( .A1(n2879), .A2(n4061), .ZN(n2881) );
  NAND2_X1 U3690 ( .A1(n2789), .A2(n4064), .ZN(n2880) );
  OAI211_X1 U3691 ( .C1(n4284), .C2(n2882), .A(n2881), .B(n2880), .ZN(n2883)
         );
  AOI21_X1 U3692 ( .B1(n2884), .B2(n4057), .A(n2883), .ZN(n2888) );
  AND2_X1 U3693 ( .A1(n2760), .A2(n2886), .ZN(n4543) );
  NAND2_X1 U3694 ( .A1(n4543), .A2(n3137), .ZN(n2887) );
  NAND2_X1 U3695 ( .A1(n2888), .A2(n2887), .ZN(n4541) );
  MUX2_X1 U3696 ( .A(n4541), .B(REG2_REG_1__SCAN_IN), .S(n4507), .Z(n2889) );
  INV_X1 U3697 ( .A(n2889), .ZN(n2891) );
  OR2_X1 U3698 ( .A1(n2728), .A2(n3822), .ZN(n2965) );
  OR2_X1 U3699 ( .A1(n4507), .A2(n2965), .ZN(n2950) );
  AOI22_X1 U3700 ( .A1(n4543), .A2(n4502), .B1(REG3_REG_1__SCAN_IN), .B2(n4497), .ZN(n2890) );
  OAI211_X1 U3701 ( .C1(n4006), .C2(n4540), .A(n2891), .B(n2890), .ZN(U3289)
         );
  INV_X1 U3702 ( .A(DATAO_REG_28__SCAN_IN), .ZN(n4098) );
  NAND2_X1 U3703 ( .A1(n3423), .A2(U4043), .ZN(n2892) );
  OAI21_X1 U3704 ( .B1(U4043), .B2(n4098), .A(n2892), .ZN(U3578) );
  INV_X1 U3705 ( .A(n2896), .ZN(n2898) );
  NAND2_X1 U3706 ( .A1(n2898), .A2(n2897), .ZN(n2899) );
  NAND2_X1 U3707 ( .A1(n2900), .A2(n2899), .ZN(n3025) );
  NAND2_X1 U3708 ( .A1(n3758), .A2(n2007), .ZN(n2902) );
  NAND2_X1 U3709 ( .A1(n2979), .A2(n2829), .ZN(n2901) );
  NAND2_X1 U3710 ( .A1(n2902), .A2(n2901), .ZN(n2903) );
  XNOR2_X1 U3711 ( .A(n2903), .B(n3425), .ZN(n2909) );
  INV_X1 U3712 ( .A(n2909), .ZN(n2907) );
  NAND2_X1 U3713 ( .A1(n3758), .A2(n3353), .ZN(n2905) );
  NAND2_X1 U3714 ( .A1(n2979), .A2(n2007), .ZN(n2904) );
  NAND2_X1 U3715 ( .A1(n2905), .A2(n2904), .ZN(n2908) );
  INV_X1 U3716 ( .A(n2908), .ZN(n2906) );
  NAND2_X1 U3717 ( .A1(n2907), .A2(n2906), .ZN(n3029) );
  INV_X1 U3718 ( .A(n3029), .ZN(n2910) );
  AND2_X1 U3719 ( .A1(n2909), .A2(n2908), .ZN(n3026) );
  NOR2_X1 U3720 ( .A1(n2910), .A2(n3026), .ZN(n2911) );
  XNOR2_X1 U3721 ( .A(n3025), .B(n2911), .ZN(n2917) );
  NOR2_X1 U3722 ( .A1(STATE_REG_SCAN_IN), .A2(n2912), .ZN(n4391) );
  OAI22_X1 U3723 ( .A1(n2913), .A2(n4343), .B1(n4344), .B2(n3078), .ZN(n2914)
         );
  AOI211_X1 U3724 ( .C1(n2979), .C2(n3589), .A(n4391), .B(n2914), .ZN(n2916)
         );
  NAND2_X1 U3725 ( .A1(n3578), .A2(n3018), .ZN(n2915) );
  OAI211_X1 U3726 ( .C1(n2917), .C2(n3581), .A(n2916), .B(n2915), .ZN(U3236)
         );
  XNOR2_X1 U3727 ( .A(n2918), .B(n3595), .ZN(n4546) );
  OAI21_X1 U3728 ( .B1(n3595), .B2(n2920), .A(n2919), .ZN(n2923) );
  AOI22_X1 U3729 ( .A1(n3760), .A2(n4064), .B1(n4277), .B2(n2926), .ZN(n2921)
         );
  OAI21_X1 U3730 ( .B1(n3487), .B2(n4018), .A(n2921), .ZN(n2922) );
  AOI21_X1 U3731 ( .B1(n2923), .B2(n4057), .A(n2922), .ZN(n2924) );
  OAI21_X1 U3732 ( .B1(n4546), .B2(n3212), .A(n2924), .ZN(n4547) );
  NAND2_X1 U3733 ( .A1(n4547), .A2(n4027), .ZN(n2930) );
  AOI21_X1 U3734 ( .B1(n2926), .B2(n2925), .A(n2932), .ZN(n4549) );
  OAI22_X1 U3735 ( .A1(n4027), .A2(n2927), .B1(REG3_REG_3__SCAN_IN), .B2(n3950), .ZN(n2928) );
  AOI21_X1 U3736 ( .B1(n4549), .B2(n4501), .A(n2928), .ZN(n2929) );
  OAI211_X1 U3737 ( .C1(n4546), .C2(n2950), .A(n2930), .B(n2929), .ZN(U3287)
         );
  OAI211_X1 U3738 ( .C1(n2932), .C2(n2931), .A(n2998), .B(n4574), .ZN(n4551)
         );
  NOR2_X1 U3739 ( .A1(n4551), .A2(n4334), .ZN(n2944) );
  XNOR2_X1 U3740 ( .A(n3597), .B(n2934), .ZN(n2942) );
  NAND2_X1 U3741 ( .A1(n2936), .A2(n3597), .ZN(n2937) );
  NAND2_X1 U3742 ( .A1(n2935), .A2(n2937), .ZN(n2946) );
  AOI22_X1 U3743 ( .A1(n3761), .A2(n4061), .B1(n2938), .B2(n4277), .ZN(n2940)
         );
  NAND2_X1 U3744 ( .A1(n3759), .A2(n4064), .ZN(n2939) );
  OAI211_X1 U3745 ( .C1(n2946), .C2(n3212), .A(n2940), .B(n2939), .ZN(n2941)
         );
  AOI21_X1 U3746 ( .B1(n2942), .B2(n4057), .A(n2941), .ZN(n2943) );
  INV_X1 U3747 ( .A(n2943), .ZN(n4552) );
  AOI211_X1 U3748 ( .C1(n4497), .C2(n2945), .A(n2944), .B(n4552), .ZN(n2948)
         );
  INV_X1 U3749 ( .A(n2946), .ZN(n4555) );
  AOI22_X1 U3750 ( .A1(n4555), .A2(n4502), .B1(REG2_REG_4__SCAN_IN), .B2(n4363), .ZN(n2947) );
  OAI21_X1 U3751 ( .B1(n2948), .B2(n4363), .A(n2947), .ZN(U3286) );
  OR2_X1 U3752 ( .A1(n4507), .A2(n4284), .ZN(n4056) );
  INV_X1 U3753 ( .A(n4056), .ZN(n3911) );
  AOI22_X1 U3754 ( .A1(n3911), .A2(n3459), .B1(REG3_REG_2__SCAN_IN), .B2(n4497), .ZN(n2949) );
  OAI21_X1 U3755 ( .B1(n2951), .B2(n2950), .A(n2949), .ZN(n2954) );
  MUX2_X1 U3756 ( .A(n2952), .B(REG2_REG_2__SCAN_IN), .S(n4507), .Z(n2953) );
  AOI211_X1 U3757 ( .C1(n4501), .C2(n2955), .A(n2954), .B(n2953), .ZN(n2956)
         );
  INV_X1 U3758 ( .A(n2956), .ZN(U3288) );
  XOR2_X1 U3759 ( .A(n3627), .B(n2957), .Z(n2960) );
  OAI22_X1 U3760 ( .A1(n3097), .A2(n3994), .B1(n3064), .B2(n4284), .ZN(n2958)
         );
  AOI21_X1 U3761 ( .B1(n4061), .B2(n3758), .A(n2958), .ZN(n2959) );
  OAI21_X1 U3762 ( .B1(n2960), .B2(n3998), .A(n2959), .ZN(n4565) );
  INV_X1 U3763 ( .A(n4565), .ZN(n2971) );
  INV_X1 U3764 ( .A(n4025), .ZN(n3008) );
  OAI21_X1 U3765 ( .B1(n2981), .B2(n3064), .A(n4574), .ZN(n2961) );
  NOR2_X1 U3766 ( .A1(n2961), .A2(n3074), .ZN(n4566) );
  INV_X1 U3767 ( .A(n3071), .ZN(n2962) );
  OAI22_X1 U3768 ( .A1(n4027), .A2(n2686), .B1(n2962), .B2(n3950), .ZN(n2969)
         );
  INV_X1 U3769 ( .A(n2963), .ZN(n2967) );
  AND2_X1 U3770 ( .A1(n2964), .A2(n3627), .ZN(n4564) );
  AND2_X1 U3771 ( .A1(n3212), .A2(n2965), .ZN(n2966) );
  NOR3_X1 U3772 ( .A1(n2967), .A2(n4564), .A3(n4070), .ZN(n2968) );
  AOI211_X1 U3773 ( .C1(n3008), .C2(n4566), .A(n2969), .B(n2968), .ZN(n2970)
         );
  OAI21_X1 U3774 ( .B1(n4507), .B2(n2971), .A(n2970), .ZN(U3283) );
  INV_X1 U3775 ( .A(REG0_REG_6__SCAN_IN), .ZN(n2985) );
  AND2_X1 U3776 ( .A1(n3656), .A2(n3667), .ZN(n3594) );
  XNOR2_X1 U3777 ( .A(n2972), .B(n3594), .ZN(n3022) );
  INV_X1 U3778 ( .A(n3022), .ZN(n2978) );
  XOR2_X1 U3779 ( .A(n3594), .B(n2973), .Z(n2976) );
  OAI22_X1 U3780 ( .A1(n3078), .A2(n3994), .B1(n4284), .B2(n2187), .ZN(n2974)
         );
  AOI21_X1 U3781 ( .B1(n4061), .B2(n3759), .A(n2974), .ZN(n2975) );
  OAI21_X1 U3782 ( .B1(n2976), .B2(n3998), .A(n2975), .ZN(n2977) );
  AOI21_X1 U3783 ( .B1(n3137), .B2(n3022), .A(n2977), .ZN(n3024) );
  OAI21_X1 U3784 ( .B1(n4545), .B2(n2978), .A(n3024), .ZN(n2986) );
  NAND2_X1 U3785 ( .A1(n2986), .A2(n4577), .ZN(n2984) );
  AND2_X1 U3786 ( .A1(n2999), .A2(n2979), .ZN(n2980) );
  NOR2_X1 U3787 ( .A1(n2981), .A2(n2980), .ZN(n3017) );
  NAND2_X1 U3788 ( .A1(n3017), .A2(n2982), .ZN(n2983) );
  OAI211_X1 U3789 ( .C1(n4577), .C2(n2985), .A(n2984), .B(n2983), .ZN(U3479)
         );
  INV_X1 U3790 ( .A(REG1_REG_6__SCAN_IN), .ZN(n2990) );
  NAND2_X1 U3791 ( .A1(n2986), .A2(n4588), .ZN(n2989) );
  NAND2_X1 U3792 ( .A1(n3017), .A2(n2987), .ZN(n2988) );
  OAI211_X1 U3793 ( .C1(n4588), .C2(n2990), .A(n2989), .B(n2988), .ZN(U3524)
         );
  INV_X1 U3794 ( .A(n2991), .ZN(n3652) );
  NAND2_X1 U3795 ( .A1(n3652), .A2(n3665), .ZN(n3622) );
  XNOR2_X1 U3796 ( .A(n2992), .B(n3622), .ZN(n2996) );
  AOI22_X1 U3797 ( .A1(n3758), .A2(n4064), .B1(n2993), .B2(n4277), .ZN(n2994)
         );
  OAI21_X1 U3798 ( .B1(n3486), .B2(n4018), .A(n2994), .ZN(n2995) );
  AOI21_X1 U3799 ( .B1(n2996), .B2(n4057), .A(n2995), .ZN(n4557) );
  XOR2_X1 U3800 ( .A(n2997), .B(n3622), .Z(n4562) );
  INV_X1 U3801 ( .A(n2998), .ZN(n3001) );
  OAI21_X1 U3802 ( .B1(n3001), .B2(n3000), .A(n2999), .ZN(n4558) );
  NOR2_X1 U3803 ( .A1(n4558), .A2(n4006), .ZN(n3004) );
  OAI22_X1 U3804 ( .A1(n4027), .A2(n2683), .B1(n3002), .B2(n3950), .ZN(n3003)
         );
  AOI211_X1 U3805 ( .C1(n4562), .C2(n3979), .A(n3004), .B(n3003), .ZN(n3005)
         );
  OAI21_X1 U3806 ( .B1(n4507), .B2(n4557), .A(n3005), .ZN(U3285) );
  INV_X1 U3807 ( .A(n3006), .ZN(n3007) );
  AOI21_X1 U3808 ( .B1(n3008), .B2(n3007), .A(n3911), .ZN(n3016) );
  INV_X1 U3809 ( .A(n3625), .ZN(n3013) );
  AOI22_X1 U3810 ( .A1(n3009), .A2(n4027), .B1(REG3_REG_0__SCAN_IN), .B2(n4497), .ZN(n3010) );
  OAI21_X1 U3811 ( .B1(n3011), .B2(n4027), .A(n3010), .ZN(n3012) );
  AOI21_X1 U3812 ( .B1(n4502), .B2(n3013), .A(n3012), .ZN(n3014) );
  OAI21_X1 U3813 ( .B1(n3016), .B2(n3015), .A(n3014), .ZN(U3290) );
  INV_X1 U3814 ( .A(n3017), .ZN(n3020) );
  INV_X1 U3815 ( .A(n4027), .ZN(n4363) );
  AOI22_X1 U3816 ( .A1(n4363), .A2(REG2_REG_6__SCAN_IN), .B1(n3018), .B2(n4497), .ZN(n3019) );
  OAI21_X1 U3817 ( .B1(n3020), .B2(n4006), .A(n3019), .ZN(n3021) );
  AOI21_X1 U3818 ( .B1(n3022), .B2(n4502), .A(n3021), .ZN(n3023) );
  OAI21_X1 U3819 ( .B1(n3024), .B2(n4363), .A(n3023), .ZN(U3284) );
  INV_X1 U3820 ( .A(n3025), .ZN(n3028) );
  INV_X1 U3821 ( .A(n3026), .ZN(n3027) );
  NAND2_X1 U3822 ( .A1(n3046), .A2(n2007), .ZN(n3031) );
  NAND2_X1 U3823 ( .A1(n3033), .A2(n2829), .ZN(n3030) );
  NAND2_X1 U3824 ( .A1(n3031), .A2(n3030), .ZN(n3032) );
  XNOR2_X1 U3825 ( .A(n3032), .B(n2860), .ZN(n3035) );
  AOI22_X1 U3826 ( .A1(n3046), .A2(n2005), .B1(n3033), .B2(n2007), .ZN(n3036)
         );
  XNOR2_X1 U3827 ( .A(n3035), .B(n3036), .ZN(n3068) );
  INV_X1 U3828 ( .A(n3035), .ZN(n3038) );
  INV_X1 U3829 ( .A(n3036), .ZN(n3037) );
  NAND2_X1 U3830 ( .A1(n3038), .A2(n3037), .ZN(n3039) );
  NAND2_X1 U3831 ( .A1(n3757), .A2(n2005), .ZN(n3041) );
  OR2_X1 U3832 ( .A1(n3077), .A2(n2862), .ZN(n3040) );
  NAND2_X1 U3833 ( .A1(n3041), .A2(n3040), .ZN(n3092) );
  NAND2_X1 U3834 ( .A1(n3757), .A2(n2007), .ZN(n3043) );
  OR2_X1 U3835 ( .A1(n3077), .A2(n3427), .ZN(n3042) );
  NAND2_X1 U3836 ( .A1(n3043), .A2(n3042), .ZN(n3044) );
  XNOR2_X1 U3837 ( .A(n3044), .B(n3425), .ZN(n3091) );
  XOR2_X1 U3838 ( .A(n3092), .B(n3091), .Z(n3045) );
  XNOR2_X1 U3839 ( .A(n3093), .B(n3045), .ZN(n3050) );
  AOI22_X1 U3840 ( .A1(n3476), .A2(n3046), .B1(n3475), .B2(n3756), .ZN(n3047)
         );
  NAND2_X1 U3841 ( .A1(REG3_REG_8__SCAN_IN), .A2(U3149), .ZN(n4395) );
  OAI211_X1 U3842 ( .C1(n4349), .C2(n3077), .A(n3047), .B(n4395), .ZN(n3048)
         );
  AOI21_X1 U3843 ( .B1(n4498), .B2(n3578), .A(n3048), .ZN(n3049) );
  OAI21_X1 U3844 ( .B1(n3050), .B2(n3581), .A(n3049), .ZN(U3218) );
  INV_X1 U3845 ( .A(n3663), .ZN(n3669) );
  NAND2_X1 U3846 ( .A1(n3669), .A2(n3661), .ZN(n3599) );
  XNOR2_X1 U3847 ( .A(n3051), .B(n3599), .ZN(n4570) );
  XOR2_X1 U3848 ( .A(n3599), .B(n3052), .Z(n3056) );
  OAI22_X1 U3849 ( .A1(n3181), .A2(n3994), .B1(n4284), .B2(n3053), .ZN(n3054)
         );
  AOI21_X1 U3850 ( .B1(n4061), .B2(n3757), .A(n3054), .ZN(n3055) );
  OAI21_X1 U3851 ( .B1(n3056), .B2(n3998), .A(n3055), .ZN(n4571) );
  NAND2_X1 U3852 ( .A1(n4571), .A2(n4027), .ZN(n3061) );
  AOI21_X1 U3853 ( .B1(n3100), .B2(n3073), .A(n2052), .ZN(n4573) );
  INV_X1 U3854 ( .A(n3101), .ZN(n3057) );
  OAI22_X1 U3855 ( .A1(n4027), .A2(n3058), .B1(n3057), .B2(n3950), .ZN(n3059)
         );
  AOI21_X1 U3856 ( .B1(n4573), .B2(n4501), .A(n3059), .ZN(n3060) );
  OAI211_X1 U3857 ( .C1(n4070), .C2(n4570), .A(n3061), .B(n3060), .ZN(U3281)
         );
  AOI22_X1 U3858 ( .A1(n3475), .A2(n3757), .B1(n3476), .B2(n3758), .ZN(n3063)
         );
  OAI211_X1 U3859 ( .C1(n4349), .C2(n3064), .A(n3063), .B(n3062), .ZN(n3070)
         );
  INV_X1 U3860 ( .A(n3065), .ZN(n3066) );
  AOI211_X1 U3861 ( .C1(n3068), .C2(n3067), .A(n3581), .B(n3066), .ZN(n3069)
         );
  AOI211_X1 U3862 ( .C1(n3071), .C2(n3578), .A(n3070), .B(n3069), .ZN(n3072)
         );
  INV_X1 U3863 ( .A(n3072), .ZN(U3210) );
  OAI21_X1 U3864 ( .B1(n3074), .B2(n3077), .A(n3073), .ZN(n4499) );
  INV_X1 U3865 ( .A(REG0_REG_8__SCAN_IN), .ZN(n3084) );
  NAND2_X1 U3866 ( .A1(n3660), .A2(n3668), .ZN(n3598) );
  XOR2_X1 U3867 ( .A(n3075), .B(n3598), .Z(n4503) );
  XOR2_X1 U3868 ( .A(n3598), .B(n3076), .Z(n3081) );
  OAI22_X1 U3869 ( .A1(n3078), .A2(n4018), .B1(n4284), .B2(n3077), .ZN(n3079)
         );
  AOI21_X1 U3870 ( .B1(n4064), .B2(n3756), .A(n3079), .ZN(n3080) );
  OAI21_X1 U3871 ( .B1(n3081), .B2(n3998), .A(n3080), .ZN(n3082) );
  AOI21_X1 U3872 ( .B1(n3137), .B2(n4503), .A(n3082), .ZN(n4506) );
  INV_X1 U3873 ( .A(n4506), .ZN(n3083) );
  AOI21_X1 U3874 ( .B1(n4554), .B2(n4503), .A(n3083), .ZN(n3086) );
  MUX2_X1 U3875 ( .A(n3084), .B(n3086), .S(n4577), .Z(n3085) );
  OAI21_X1 U3876 ( .B1(n4499), .B2(n4332), .A(n3085), .ZN(U3483) );
  MUX2_X1 U3877 ( .A(n4394), .B(n3086), .S(n4588), .Z(n3087) );
  OAI21_X1 U3878 ( .B1(n4499), .B2(n4289), .A(n3087), .ZN(U3526) );
  NAND2_X1 U3879 ( .A1(n3756), .A2(n2007), .ZN(n3089) );
  NAND2_X1 U3880 ( .A1(n3100), .A2(n2829), .ZN(n3088) );
  NAND2_X1 U3881 ( .A1(n3089), .A2(n3088), .ZN(n3090) );
  XNOR2_X1 U3882 ( .A(n3090), .B(n2860), .ZN(n3106) );
  AOI22_X1 U3883 ( .A1(n3756), .A2(n3353), .B1(n3100), .B2(n2007), .ZN(n3105)
         );
  XNOR2_X1 U3884 ( .A(n3106), .B(n3105), .ZN(n3096) );
  INV_X1 U3885 ( .A(n3112), .ZN(n3094) );
  AOI21_X1 U3886 ( .B1(n3096), .B2(n3095), .A(n3094), .ZN(n3104) );
  OAI22_X1 U3887 ( .A1(n3097), .A2(n4343), .B1(n4344), .B2(n3181), .ZN(n3098)
         );
  AOI211_X1 U3888 ( .C1(n3100), .C2(n3589), .A(n3099), .B(n3098), .ZN(n3103)
         );
  NAND2_X1 U3889 ( .A1(n3578), .A2(n3101), .ZN(n3102) );
  OAI211_X1 U3890 ( .C1(n3104), .C2(n3581), .A(n3103), .B(n3102), .ZN(U3228)
         );
  NAND2_X1 U3891 ( .A1(n3106), .A2(n3105), .ZN(n3110) );
  AND2_X1 U3892 ( .A1(n3112), .A2(n3110), .ZN(n3114) );
  NAND2_X1 U3893 ( .A1(n3154), .A2(n2007), .ZN(n3108) );
  NAND2_X1 U3894 ( .A1(n3118), .A2(n2829), .ZN(n3107) );
  NAND2_X1 U3895 ( .A1(n3108), .A2(n3107), .ZN(n3109) );
  XNOR2_X1 U3896 ( .A(n3109), .B(n3425), .ZN(n3176) );
  AOI22_X1 U3897 ( .A1(n3154), .A2(n2005), .B1(n3118), .B2(n2007), .ZN(n3174)
         );
  XNOR2_X1 U3898 ( .A(n3176), .B(n3174), .ZN(n3113) );
  AND2_X1 U3899 ( .A1(n3113), .A2(n3110), .ZN(n3111) );
  OAI211_X1 U3900 ( .C1(n3114), .C2(n3113), .A(n4357), .B(n3178), .ZN(n3120)
         );
  INV_X1 U3901 ( .A(REG3_REG_10__SCAN_IN), .ZN(n4182) );
  NOR2_X1 U3902 ( .A1(STATE_REG_SCAN_IN), .A2(n4182), .ZN(n4405) );
  OAI22_X1 U3903 ( .A1(n3116), .A2(n4343), .B1(n4344), .B2(n3115), .ZN(n3117)
         );
  AOI211_X1 U3904 ( .C1(n3118), .C2(n3589), .A(n4405), .B(n3117), .ZN(n3119)
         );
  OAI211_X1 U3905 ( .C1(n4362), .C2(n3121), .A(n3120), .B(n3119), .ZN(U3214)
         );
  INV_X1 U3906 ( .A(n3122), .ZN(n3123) );
  AOI21_X1 U3907 ( .B1(n3152), .B2(n3124), .A(n3123), .ZN(n3206) );
  NAND2_X1 U3908 ( .A1(n3205), .A2(n3203), .ZN(n3619) );
  XNOR2_X1 U3909 ( .A(n3206), .B(n3619), .ZN(n3125) );
  NAND2_X1 U3910 ( .A1(n3125), .A2(n4057), .ZN(n3127) );
  AOI22_X1 U3911 ( .A1(n4061), .A2(n3755), .B1(n3753), .B2(n4064), .ZN(n3126)
         );
  XNOR2_X1 U3912 ( .A(n3128), .B(n3619), .ZN(n3254) );
  OR2_X1 U3913 ( .A1(n3160), .A2(n3257), .ZN(n3129) );
  NAND2_X1 U3914 ( .A1(n3214), .A2(n3129), .ZN(n3263) );
  AOI22_X1 U3915 ( .A1(n4507), .A2(REG2_REG_12__SCAN_IN), .B1(n3199), .B2(
        n4497), .ZN(n3132) );
  NAND2_X1 U3916 ( .A1(n3911), .A2(n3130), .ZN(n3131) );
  OAI211_X1 U3917 ( .C1(n3263), .C2(n4006), .A(n3132), .B(n3131), .ZN(n3133)
         );
  AOI21_X1 U3918 ( .B1(n3254), .B2(n3979), .A(n3133), .ZN(n3134) );
  OAI21_X1 U3919 ( .B1(n3256), .B2(n4363), .A(n3134), .ZN(U3278) );
  INV_X1 U3920 ( .A(n3163), .ZN(n3135) );
  OAI21_X1 U3921 ( .B1(n2052), .B2(n3142), .A(n3135), .ZN(n4491) );
  NAND2_X1 U3922 ( .A1(n3671), .A2(n3676), .ZN(n3620) );
  XNOR2_X1 U3923 ( .A(n3136), .B(n3620), .ZN(n4493) );
  NAND2_X1 U3924 ( .A1(n4493), .A2(n3137), .ZN(n3146) );
  INV_X1 U3925 ( .A(n3620), .ZN(n3138) );
  XNOR2_X1 U3926 ( .A(n3139), .B(n3138), .ZN(n3144) );
  NAND2_X1 U3927 ( .A1(n3755), .A2(n4064), .ZN(n3141) );
  NAND2_X1 U3928 ( .A1(n3756), .A2(n4061), .ZN(n3140) );
  OAI211_X1 U3929 ( .C1(n4284), .C2(n3142), .A(n3141), .B(n3140), .ZN(n3143)
         );
  AOI21_X1 U3930 ( .B1(n3144), .B2(n4057), .A(n3143), .ZN(n3145) );
  AND2_X1 U3931 ( .A1(n3146), .A2(n3145), .ZN(n4496) );
  NAND2_X1 U3932 ( .A1(n4493), .A2(n4554), .ZN(n3147) );
  AND2_X1 U3933 ( .A1(n4496), .A2(n3147), .ZN(n3150) );
  INV_X1 U3934 ( .A(REG0_REG_10__SCAN_IN), .ZN(n3148) );
  MUX2_X1 U3935 ( .A(n3150), .B(n3148), .S(n4575), .Z(n3149) );
  OAI21_X1 U3936 ( .B1(n4491), .B2(n4332), .A(n3149), .ZN(U3487) );
  INV_X1 U3937 ( .A(REG1_REG_10__SCAN_IN), .ZN(n4404) );
  MUX2_X1 U3938 ( .A(n4404), .B(n3150), .S(n4588), .Z(n3151) );
  OAI21_X1 U3939 ( .B1(n4491), .B2(n4289), .A(n3151), .ZN(U3528) );
  XNOR2_X1 U3940 ( .A(n3152), .B(n3628), .ZN(n3158) );
  AOI21_X1 U3941 ( .B1(n3628), .B2(n3153), .A(n2040), .ZN(n3159) );
  AOI22_X1 U3942 ( .A1(n3754), .A2(n4064), .B1(n3183), .B2(n4277), .ZN(n3156)
         );
  NAND2_X1 U3943 ( .A1(n3154), .A2(n4061), .ZN(n3155) );
  OAI211_X1 U3944 ( .C1(n3159), .C2(n3212), .A(n3156), .B(n3155), .ZN(n3157)
         );
  AOI21_X1 U3945 ( .B1(n3158), .B2(n4057), .A(n3157), .ZN(n3293) );
  INV_X1 U3946 ( .A(n3159), .ZN(n3295) );
  INV_X1 U3947 ( .A(n3160), .ZN(n3161) );
  OAI21_X1 U3948 ( .B1(n3163), .B2(n3162), .A(n3161), .ZN(n3300) );
  AOI22_X1 U3949 ( .A1(n4363), .A2(REG2_REG_11__SCAN_IN), .B1(n3184), .B2(
        n4497), .ZN(n3164) );
  OAI21_X1 U3950 ( .B1(n3300), .B2(n4006), .A(n3164), .ZN(n3165) );
  AOI21_X1 U3951 ( .B1(n3295), .B2(n4502), .A(n3165), .ZN(n3166) );
  OAI21_X1 U3952 ( .B1(n3293), .B2(n4363), .A(n3166), .ZN(U3279) );
  NAND2_X1 U3953 ( .A1(n3755), .A2(n2007), .ZN(n3168) );
  NAND2_X1 U3954 ( .A1(n3183), .A2(n2829), .ZN(n3167) );
  NAND2_X1 U3955 ( .A1(n3168), .A2(n3167), .ZN(n3169) );
  XNOR2_X1 U3956 ( .A(n3169), .B(n2860), .ZN(n3173) );
  INV_X1 U3957 ( .A(n3173), .ZN(n3171) );
  AOI22_X1 U3958 ( .A1(n3755), .A2(n2005), .B1(n3183), .B2(n2007), .ZN(n3172)
         );
  INV_X1 U3959 ( .A(n3172), .ZN(n3170) );
  NAND2_X1 U3960 ( .A1(n3171), .A2(n3170), .ZN(n3190) );
  NAND2_X1 U3961 ( .A1(n3173), .A2(n3172), .ZN(n3188) );
  NAND2_X1 U3962 ( .A1(n3190), .A2(n3188), .ZN(n3179) );
  INV_X1 U3963 ( .A(n3174), .ZN(n3175) );
  NAND2_X1 U3964 ( .A1(n3176), .A2(n3175), .ZN(n3177) );
  XOR2_X1 U3965 ( .A(n3179), .B(n3189), .Z(n3187) );
  INV_X1 U3966 ( .A(REG3_REG_11__SCAN_IN), .ZN(n3180) );
  NOR2_X1 U3967 ( .A1(STATE_REG_SCAN_IN), .A2(n3180), .ZN(n4413) );
  OAI22_X1 U3968 ( .A1(n3323), .A2(n4344), .B1(n4343), .B2(n3181), .ZN(n3182)
         );
  AOI211_X1 U3969 ( .C1(n3183), .C2(n3589), .A(n4413), .B(n3182), .ZN(n3186)
         );
  NAND2_X1 U3970 ( .A1(n3578), .A2(n3184), .ZN(n3185) );
  OAI211_X1 U3971 ( .C1(n3187), .C2(n3581), .A(n3186), .B(n3185), .ZN(U3233)
         );
  NAND2_X1 U3972 ( .A1(n3754), .A2(n2007), .ZN(n3192) );
  OR2_X1 U3973 ( .A1(n3257), .A2(n3427), .ZN(n3191) );
  NAND2_X1 U3974 ( .A1(n3192), .A2(n3191), .ZN(n3193) );
  XNOR2_X1 U3975 ( .A(n3193), .B(n3425), .ZN(n3317) );
  NAND2_X1 U3976 ( .A1(n3754), .A2(n3353), .ZN(n3195) );
  OR2_X1 U3977 ( .A1(n3257), .A2(n2862), .ZN(n3194) );
  NAND2_X1 U3978 ( .A1(n3195), .A2(n3194), .ZN(n3316) );
  INV_X1 U3979 ( .A(n3316), .ZN(n3271) );
  XNOR2_X1 U3980 ( .A(n3317), .B(n3271), .ZN(n3196) );
  XNOR2_X1 U3981 ( .A(n3279), .B(n3196), .ZN(n3201) );
  AOI22_X1 U3982 ( .A1(n3476), .A2(n3755), .B1(n3475), .B2(n3753), .ZN(n3197)
         );
  NAND2_X1 U3983 ( .A1(REG3_REG_12__SCAN_IN), .A2(U3149), .ZN(n4423) );
  OAI211_X1 U3984 ( .C1(n4349), .C2(n3257), .A(n3197), .B(n4423), .ZN(n3198)
         );
  AOI21_X1 U3985 ( .B1(n3199), .B2(n3578), .A(n3198), .ZN(n3200) );
  OAI21_X1 U3986 ( .B1(n3201), .B2(n3581), .A(n3200), .ZN(U3221) );
  XNOR2_X1 U3987 ( .A(n3753), .B(n3267), .ZN(n3631) );
  XOR2_X1 U3988 ( .A(n3631), .B(n3202), .Z(n3213) );
  INV_X1 U3989 ( .A(n3203), .ZN(n3204) );
  AOI21_X1 U3990 ( .B1(n3206), .B2(n3205), .A(n3204), .ZN(n3207) );
  XOR2_X1 U3991 ( .A(n3631), .B(n3207), .Z(n3210) );
  AOI22_X1 U3992 ( .A1(n3283), .A2(n4064), .B1(n3326), .B2(n4277), .ZN(n3208)
         );
  OAI21_X1 U3993 ( .B1(n3323), .B2(n4018), .A(n3208), .ZN(n3209) );
  AOI21_X1 U3994 ( .B1(n3210), .B2(n4057), .A(n3209), .ZN(n3211) );
  OAI21_X1 U3995 ( .B1(n3213), .B2(n3212), .A(n3211), .ZN(n3331) );
  INV_X1 U3996 ( .A(n3331), .ZN(n3219) );
  INV_X1 U3997 ( .A(n3213), .ZN(n3332) );
  INV_X1 U3998 ( .A(n3214), .ZN(n3215) );
  OAI21_X1 U3999 ( .B1(n3215), .B2(n3267), .A(n3247), .ZN(n3337) );
  AOI22_X1 U4000 ( .A1(n4363), .A2(REG2_REG_13__SCAN_IN), .B1(n3327), .B2(
        n4497), .ZN(n3216) );
  OAI21_X1 U4001 ( .B1(n3337), .B2(n4006), .A(n3216), .ZN(n3217) );
  AOI21_X1 U4002 ( .B1(n3332), .B2(n4502), .A(n3217), .ZN(n3218) );
  OAI21_X1 U4003 ( .B1(n3219), .B2(n4363), .A(n3218), .ZN(U3277) );
  NAND2_X1 U4004 ( .A1(n3235), .A2(REG2_REG_11__SCAN_IN), .ZN(n3225) );
  INV_X1 U4005 ( .A(n3235), .ZN(n4531) );
  AOI22_X1 U4006 ( .A1(n3235), .A2(REG2_REG_11__SCAN_IN), .B1(n2378), .B2(
        n4531), .ZN(n4417) );
  OAI21_X1 U4007 ( .B1(n3058), .B2(n3221), .A(n3220), .ZN(n3223) );
  NAND2_X1 U4008 ( .A1(n3222), .A2(n3223), .ZN(n3224) );
  INV_X1 U4009 ( .A(n3222), .ZN(n4533) );
  XNOR2_X1 U4010 ( .A(n4533), .B(n3223), .ZN(n4408) );
  NAND2_X1 U4011 ( .A1(REG2_REG_10__SCAN_IN), .A2(n4408), .ZN(n4407) );
  NAND2_X1 U4012 ( .A1(n3224), .A2(n4407), .ZN(n4416) );
  NAND2_X1 U4013 ( .A1(n3226), .A2(n3227), .ZN(n3228) );
  NAND2_X1 U4014 ( .A1(n3228), .A2(n4426), .ZN(n3811) );
  NOR2_X1 U4015 ( .A1(n3244), .A2(n2267), .ZN(n3810) );
  AOI21_X1 U4016 ( .B1(n2267), .B2(n3244), .A(n3810), .ZN(n3230) );
  AOI21_X1 U4017 ( .B1(n3230), .B2(n3811), .A(n4479), .ZN(n3229) );
  OAI21_X1 U4018 ( .B1(n3811), .B2(n3230), .A(n3229), .ZN(n3243) );
  NOR2_X1 U4019 ( .A1(STATE_REG_SCAN_IN), .A2(n3231), .ZN(n3325) );
  INV_X1 U4020 ( .A(REG1_REG_12__SCAN_IN), .ZN(n4422) );
  NOR2_X1 U4021 ( .A1(n3233), .A2(n4533), .ZN(n3234) );
  INV_X1 U4022 ( .A(REG1_REG_11__SCAN_IN), .ZN(n3298) );
  AOI22_X1 U4023 ( .A1(n3235), .A2(n3298), .B1(REG1_REG_11__SCAN_IN), .B2(
        n4531), .ZN(n4412) );
  XNOR2_X1 U4024 ( .A(n3236), .B(n4529), .ZN(n4421) );
  NAND2_X1 U4025 ( .A1(n3809), .A2(REG1_REG_13__SCAN_IN), .ZN(n3796) );
  INV_X1 U4026 ( .A(REG1_REG_13__SCAN_IN), .ZN(n4197) );
  NAND2_X1 U4027 ( .A1(n3244), .A2(n4197), .ZN(n3237) );
  NAND2_X1 U4028 ( .A1(n3796), .A2(n3237), .ZN(n3239) );
  INV_X1 U4029 ( .A(n3797), .ZN(n3238) );
  AOI211_X1 U4030 ( .C1(n3240), .C2(n3239), .A(n3238), .B(n4476), .ZN(n3241)
         );
  AOI211_X1 U4031 ( .C1(n4462), .C2(ADDR_REG_13__SCAN_IN), .A(n3325), .B(n3241), .ZN(n3242) );
  OAI211_X1 U4032 ( .C1(n4475), .C2(n3244), .A(n3243), .B(n3242), .ZN(U3253)
         );
  XNOR2_X1 U4033 ( .A(n3719), .B(n2205), .ZN(n3245) );
  AOI222_X1 U4034 ( .A1(n4057), .A2(n3245), .B1(n3753), .B2(n4061), .C1(n4062), 
        .C2(n4064), .ZN(n4283) );
  OAI21_X1 U4035 ( .B1(n2051), .B2(n3621), .A(n3246), .ZN(n4287) );
  NAND2_X1 U4036 ( .A1(n4287), .A2(n3979), .ZN(n3253) );
  INV_X1 U4037 ( .A(n3247), .ZN(n3248) );
  OAI21_X1 U4038 ( .B1(n3248), .B2(n4285), .A(n3302), .ZN(n4333) );
  INV_X1 U4039 ( .A(n4333), .ZN(n3251) );
  AOI22_X1 U4040 ( .A1(n4363), .A2(REG2_REG_14__SCAN_IN), .B1(n3290), .B2(
        n4497), .ZN(n3249) );
  OAI21_X1 U4041 ( .B1(n4056), .B2(n4285), .A(n3249), .ZN(n3250) );
  AOI21_X1 U4042 ( .B1(n3251), .B2(n4501), .A(n3250), .ZN(n3252) );
  OAI211_X1 U40430 ( .C1(n4507), .C2(n4283), .A(n3253), .B(n3252), .ZN(U3276)
         );
  NAND2_X1 U4044 ( .A1(n3254), .A2(n4561), .ZN(n3255) );
  OAI211_X1 U4045 ( .C1(n4284), .C2(n3257), .A(n3256), .B(n3255), .ZN(n3260)
         );
  MUX2_X1 U4046 ( .A(REG0_REG_12__SCAN_IN), .B(n3260), .S(n4577), .Z(n3258) );
  INV_X1 U4047 ( .A(n3258), .ZN(n3259) );
  OAI21_X1 U4048 ( .B1(n3263), .B2(n4332), .A(n3259), .ZN(U3491) );
  MUX2_X1 U4049 ( .A(REG1_REG_12__SCAN_IN), .B(n3260), .S(n4588), .Z(n3261) );
  INV_X1 U4050 ( .A(n3261), .ZN(n3262) );
  OAI21_X1 U4051 ( .B1(n4289), .B2(n3263), .A(n3262), .ZN(U3530) );
  NAND2_X1 U4052 ( .A1(n3753), .A2(n2007), .ZN(n3265) );
  OR2_X1 U4053 ( .A1(n3267), .A2(n3427), .ZN(n3264) );
  NAND2_X1 U4054 ( .A1(n3265), .A2(n3264), .ZN(n3266) );
  XNOR2_X1 U4055 ( .A(n3266), .B(n3425), .ZN(n3272) );
  NAND2_X1 U4056 ( .A1(n3753), .A2(n2005), .ZN(n3269) );
  OR2_X1 U4057 ( .A1(n3267), .A2(n2862), .ZN(n3268) );
  NAND2_X1 U4058 ( .A1(n3269), .A2(n3268), .ZN(n3273) );
  NAND2_X1 U4059 ( .A1(n3272), .A2(n3273), .ZN(n3315) );
  NAND2_X1 U4060 ( .A1(n3317), .A2(n3316), .ZN(n3270) );
  NAND2_X1 U4061 ( .A1(n3315), .A2(n3270), .ZN(n3278) );
  INV_X1 U4062 ( .A(n3317), .ZN(n3319) );
  NAND3_X1 U4063 ( .A1(n3315), .A2(n3271), .A3(n3319), .ZN(n3276) );
  INV_X1 U4064 ( .A(n3272), .ZN(n3275) );
  INV_X1 U4065 ( .A(n3273), .ZN(n3274) );
  NAND2_X1 U4066 ( .A1(n3275), .A2(n3274), .ZN(n3314) );
  NAND2_X1 U4067 ( .A1(n3283), .A2(n2007), .ZN(n3281) );
  NAND2_X1 U4068 ( .A1(n3284), .A2(n2829), .ZN(n3280) );
  NAND2_X1 U4069 ( .A1(n3281), .A2(n3280), .ZN(n3282) );
  XNOR2_X1 U4070 ( .A(n3282), .B(n2860), .ZN(n3338) );
  INV_X1 U4071 ( .A(n3338), .ZN(n3342) );
  NAND2_X1 U4072 ( .A1(n3283), .A2(n2005), .ZN(n3286) );
  NAND2_X1 U4073 ( .A1(n3284), .A2(n2007), .ZN(n3285) );
  NAND2_X1 U4074 ( .A1(n3286), .A2(n3285), .ZN(n3339) );
  XNOR2_X1 U4075 ( .A(n3342), .B(n3339), .ZN(n3287) );
  XNOR2_X1 U4076 ( .A(n3341), .B(n3287), .ZN(n3292) );
  AOI22_X1 U4077 ( .A1(n3475), .A2(n4062), .B1(n3476), .B2(n3753), .ZN(n3288)
         );
  NAND2_X1 U4078 ( .A1(REG3_REG_14__SCAN_IN), .A2(U3149), .ZN(n4438) );
  OAI211_X1 U4079 ( .C1(n4349), .C2(n4285), .A(n3288), .B(n4438), .ZN(n3289)
         );
  AOI21_X1 U4080 ( .B1(n3290), .B2(n3578), .A(n3289), .ZN(n3291) );
  OAI21_X1 U4081 ( .B1(n3292), .B2(n3581), .A(n3291), .ZN(U3212) );
  INV_X1 U4082 ( .A(REG0_REG_11__SCAN_IN), .ZN(n4131) );
  INV_X1 U4083 ( .A(n3293), .ZN(n3294) );
  AOI21_X1 U4084 ( .B1(n4554), .B2(n3295), .A(n3294), .ZN(n3297) );
  MUX2_X1 U4085 ( .A(n4131), .B(n3297), .S(n4577), .Z(n3296) );
  OAI21_X1 U4086 ( .B1(n3300), .B2(n4332), .A(n3296), .ZN(U3489) );
  MUX2_X1 U4087 ( .A(n3298), .B(n3297), .S(n4588), .Z(n3299) );
  OAI21_X1 U4088 ( .B1(n4289), .B2(n3300), .A(n3299), .ZN(U3529) );
  XNOR2_X1 U4089 ( .A(n3301), .B(n2076), .ZN(n4282) );
  AOI21_X1 U4090 ( .B1(n4278), .B2(n3302), .A(n4050), .ZN(n4279) );
  AOI22_X1 U4091 ( .A1(n4363), .A2(REG2_REG_15__SCAN_IN), .B1(n3303), .B2(
        n4497), .ZN(n3304) );
  OAI21_X1 U4092 ( .B1(n4056), .B2(n3305), .A(n3304), .ZN(n3312) );
  AOI21_X1 U4093 ( .B1(n3307), .B2(n3306), .A(n3998), .ZN(n3310) );
  OAI22_X1 U4094 ( .A1(n3587), .A2(n4018), .B1(n3586), .B2(n3994), .ZN(n3308)
         );
  AOI21_X1 U4095 ( .B1(n3310), .B2(n3309), .A(n3308), .ZN(n4281) );
  NOR2_X1 U4096 ( .A1(n4281), .A2(n4363), .ZN(n3311) );
  AOI211_X1 U4097 ( .C1(n4279), .C2(n4501), .A(n3312), .B(n3311), .ZN(n3313)
         );
  OAI21_X1 U4098 ( .B1(n4282), .B2(n4070), .A(n3313), .ZN(U3275) );
  NAND2_X1 U4099 ( .A1(n3315), .A2(n3314), .ZN(n3322) );
  INV_X1 U4100 ( .A(n3279), .ZN(n3320) );
  OAI21_X1 U4101 ( .B1(n3279), .B2(n3317), .A(n3316), .ZN(n3318) );
  OAI21_X1 U4102 ( .B1(n3320), .B2(n3319), .A(n3318), .ZN(n3321) );
  XOR2_X1 U4103 ( .A(n3322), .B(n3321), .Z(n3330) );
  OAI22_X1 U4104 ( .A1(n3323), .A2(n4343), .B1(n4344), .B2(n3587), .ZN(n3324)
         );
  AOI211_X1 U4105 ( .C1(n3326), .C2(n3589), .A(n3325), .B(n3324), .ZN(n3329)
         );
  NAND2_X1 U4106 ( .A1(n3578), .A2(n3327), .ZN(n3328) );
  OAI211_X1 U4107 ( .C1(n3330), .C2(n3581), .A(n3329), .B(n3328), .ZN(U3231)
         );
  INV_X1 U4108 ( .A(REG0_REG_13__SCAN_IN), .ZN(n3333) );
  AOI21_X1 U4109 ( .B1(n4554), .B2(n3332), .A(n3331), .ZN(n3335) );
  MUX2_X1 U4110 ( .A(n3333), .B(n3335), .S(n4577), .Z(n3334) );
  OAI21_X1 U4111 ( .B1(n3337), .B2(n4332), .A(n3334), .ZN(U3493) );
  MUX2_X1 U4112 ( .A(n4197), .B(n3335), .S(n4588), .Z(n3336) );
  OAI21_X1 U4113 ( .B1(n4289), .B2(n3337), .A(n3336), .ZN(U3531) );
  NAND2_X1 U4114 ( .A1(n3341), .A2(n3338), .ZN(n3340) );
  NAND2_X1 U4115 ( .A1(n3340), .A2(n3339), .ZN(n3345) );
  INV_X1 U4116 ( .A(n3341), .ZN(n3343) );
  NAND2_X1 U4117 ( .A1(n3343), .A2(n3342), .ZN(n3344) );
  NAND2_X1 U4118 ( .A1(n3345), .A2(n3344), .ZN(n3352) );
  NAND2_X1 U4119 ( .A1(n4062), .A2(n2007), .ZN(n3347) );
  NAND2_X1 U4120 ( .A1(n4278), .A2(n2829), .ZN(n3346) );
  NAND2_X1 U4121 ( .A1(n3347), .A2(n3346), .ZN(n3348) );
  XNOR2_X1 U4122 ( .A(n3348), .B(n3425), .ZN(n3351) );
  NAND2_X1 U4123 ( .A1(n4062), .A2(n2005), .ZN(n3350) );
  NAND2_X1 U4124 ( .A1(n4278), .A2(n2007), .ZN(n3349) );
  AND2_X1 U4125 ( .A1(n3350), .A2(n3349), .ZN(n4354) );
  INV_X1 U4126 ( .A(n3353), .ZN(n3424) );
  OAI22_X1 U4127 ( .A1(n3586), .A2(n3424), .B1(n4348), .B2(n2862), .ZN(n3357)
         );
  NAND2_X1 U4128 ( .A1(n4034), .A2(n2007), .ZN(n3355) );
  NAND2_X1 U4129 ( .A1(n4272), .A2(n2829), .ZN(n3354) );
  NAND2_X1 U4130 ( .A1(n3355), .A2(n3354), .ZN(n3356) );
  XNOR2_X1 U4131 ( .A(n3356), .B(n3425), .ZN(n3358) );
  XOR2_X1 U4132 ( .A(n3357), .B(n3358), .Z(n4356) );
  NAND2_X1 U4133 ( .A1(n4063), .A2(n2007), .ZN(n3360) );
  OR2_X1 U4134 ( .A1(n4038), .A2(n3427), .ZN(n3359) );
  NAND2_X1 U4135 ( .A1(n3360), .A2(n3359), .ZN(n3361) );
  XNOR2_X1 U4136 ( .A(n3361), .B(n3425), .ZN(n3526) );
  NAND2_X1 U4137 ( .A1(n4063), .A2(n3353), .ZN(n3363) );
  OR2_X1 U4138 ( .A1(n4038), .A2(n2862), .ZN(n3362) );
  NAND2_X1 U4139 ( .A1(n3363), .A2(n3362), .ZN(n3525) );
  INV_X1 U4140 ( .A(n3526), .ZN(n3365) );
  INV_X1 U4141 ( .A(n3525), .ZN(n3364) );
  NAND2_X1 U4142 ( .A1(n4035), .A2(n2007), .ZN(n3367) );
  NAND2_X1 U4143 ( .A1(n4015), .A2(n2829), .ZN(n3366) );
  NAND2_X1 U4144 ( .A1(n3367), .A2(n3366), .ZN(n3368) );
  XNOR2_X1 U4145 ( .A(n3368), .B(n2860), .ZN(n3370) );
  AOI22_X1 U4146 ( .A1(n4035), .A2(n3353), .B1(n4015), .B2(n2007), .ZN(n3369)
         );
  NOR2_X1 U4147 ( .A1(n3370), .A2(n3369), .ZN(n3562) );
  NAND2_X1 U4148 ( .A1(n3370), .A2(n3369), .ZN(n3560) );
  OAI21_X1 U4149 ( .B1(n3564), .B2(n3562), .A(n3560), .ZN(n3494) );
  OAI22_X1 U4150 ( .A1(n3565), .A2(n3424), .B1(n4002), .B2(n2862), .ZN(n3375)
         );
  NAND2_X1 U4151 ( .A1(n4016), .A2(n2007), .ZN(n3372) );
  NAND2_X1 U4152 ( .A1(n3607), .A2(n2829), .ZN(n3371) );
  NAND2_X1 U4153 ( .A1(n3372), .A2(n3371), .ZN(n3373) );
  XNOR2_X1 U4154 ( .A(n3373), .B(n3425), .ZN(n3374) );
  XOR2_X1 U4155 ( .A(n3375), .B(n3374), .Z(n3496) );
  NAND2_X1 U4156 ( .A1(n3494), .A2(n3496), .ZN(n3495) );
  NAND2_X1 U4157 ( .A1(n3495), .A2(n3378), .ZN(n3506) );
  NAND2_X1 U4158 ( .A1(n3966), .A2(n2007), .ZN(n3380) );
  OR2_X1 U4159 ( .A1(n3427), .A2(n4256), .ZN(n3379) );
  NAND2_X1 U4160 ( .A1(n3380), .A2(n3379), .ZN(n3381) );
  XNOR2_X1 U4161 ( .A(n3381), .B(n2860), .ZN(n3384) );
  NOR2_X1 U4162 ( .A1(n4256), .A2(n2862), .ZN(n3382) );
  AOI21_X1 U4163 ( .B1(n3966), .B2(n2005), .A(n3382), .ZN(n3383) );
  OR2_X1 U4164 ( .A1(n3384), .A2(n3383), .ZN(n3544) );
  NAND2_X1 U4165 ( .A1(n3506), .A2(n3544), .ZN(n3543) );
  NAND2_X1 U4166 ( .A1(n3384), .A2(n3383), .ZN(n3546) );
  OAI22_X1 U4167 ( .A1(n3974), .A2(n2862), .B1(n3963), .B2(n3427), .ZN(n3385)
         );
  XNOR2_X1 U4168 ( .A(n3385), .B(n3425), .ZN(n3389) );
  OR2_X1 U4169 ( .A1(n3974), .A2(n3424), .ZN(n3387) );
  NAND2_X1 U4170 ( .A1(n4250), .A2(n2007), .ZN(n3386) );
  NAND2_X1 U4171 ( .A1(n3387), .A2(n3386), .ZN(n3388) );
  NOR2_X1 U4172 ( .A1(n3389), .A2(n3388), .ZN(n3503) );
  NAND2_X1 U4173 ( .A1(n3389), .A2(n3388), .ZN(n3504) );
  NAND2_X1 U4174 ( .A1(n3967), .A2(n2007), .ZN(n3391) );
  OR2_X1 U4175 ( .A1(n3427), .A2(n3947), .ZN(n3390) );
  NAND2_X1 U4176 ( .A1(n3391), .A2(n3390), .ZN(n3392) );
  XNOR2_X1 U4177 ( .A(n3392), .B(n3425), .ZN(n3394) );
  OAI22_X1 U4178 ( .A1(n3926), .A2(n3424), .B1(n3947), .B2(n2862), .ZN(n3393)
         );
  XNOR2_X1 U4179 ( .A(n3394), .B(n3393), .ZN(n3554) );
  NOR2_X1 U4180 ( .A1(n3394), .A2(n3393), .ZN(n3473) );
  NAND2_X1 U4181 ( .A1(n3944), .A2(n2007), .ZN(n3396) );
  OR2_X1 U4182 ( .A1(n3427), .A2(n3933), .ZN(n3395) );
  NAND2_X1 U4183 ( .A1(n3396), .A2(n3395), .ZN(n3397) );
  XNOR2_X1 U4184 ( .A(n3397), .B(n2860), .ZN(n3400) );
  NOR2_X1 U4185 ( .A1(n3933), .A2(n2862), .ZN(n3398) );
  AOI21_X1 U4186 ( .B1(n3944), .B2(n2005), .A(n3398), .ZN(n3399) );
  XNOR2_X1 U4187 ( .A(n3400), .B(n3399), .ZN(n3472) );
  NAND2_X1 U4188 ( .A1(n3928), .A2(n2005), .ZN(n3402) );
  OR2_X1 U4189 ( .A1(n2862), .A2(n4236), .ZN(n3401) );
  NAND2_X1 U4190 ( .A1(n3402), .A2(n3401), .ZN(n3404) );
  AOI22_X1 U4191 ( .A1(n3928), .A2(n2007), .B1(n3910), .B2(n2829), .ZN(n3403)
         );
  XNOR2_X1 U4192 ( .A(n3403), .B(n3425), .ZN(n3535) );
  NAND2_X1 U4193 ( .A1(n3898), .A2(n2007), .ZN(n3406) );
  OR2_X1 U4194 ( .A1(n3427), .A2(n3888), .ZN(n3405) );
  NAND2_X1 U4195 ( .A1(n3406), .A2(n3405), .ZN(n3407) );
  XNOR2_X1 U4196 ( .A(n3407), .B(n2860), .ZN(n3410) );
  NOR2_X1 U4197 ( .A1(n3888), .A2(n2862), .ZN(n3408) );
  AOI21_X1 U4198 ( .B1(n3898), .B2(n3353), .A(n3408), .ZN(n3409) );
  NAND2_X1 U4199 ( .A1(n3410), .A2(n3409), .ZN(n3516) );
  NOR2_X1 U4200 ( .A1(n3410), .A2(n3409), .ZN(n3517) );
  NAND2_X1 U4201 ( .A1(n3883), .A2(n2007), .ZN(n3412) );
  OR2_X1 U4202 ( .A1(n3427), .A2(n3872), .ZN(n3411) );
  NAND2_X1 U4203 ( .A1(n3412), .A2(n3411), .ZN(n3413) );
  XNOR2_X1 U4204 ( .A(n3413), .B(n2860), .ZN(n3416) );
  NOR2_X1 U4205 ( .A1(n3872), .A2(n2862), .ZN(n3414) );
  AOI21_X1 U4206 ( .B1(n3883), .B2(n2005), .A(n3414), .ZN(n3415) );
  OR2_X1 U4207 ( .A1(n3416), .A2(n3415), .ZN(n3571) );
  AND2_X1 U4208 ( .A1(n3416), .A2(n3415), .ZN(n3570) );
  AOI21_X1 U4209 ( .B1(n3574), .B2(n3571), .A(n3570), .ZN(n3465) );
  OAI22_X1 U4210 ( .A1(n3575), .A2(n2862), .B1(n4087), .B2(n3427), .ZN(n3417)
         );
  XNOR2_X1 U4211 ( .A(n3417), .B(n2860), .ZN(n3420) );
  OR2_X1 U4212 ( .A1(n3575), .A2(n3424), .ZN(n3419) );
  NAND2_X1 U4213 ( .A1(n3855), .A2(n2007), .ZN(n3418) );
  NAND2_X1 U4214 ( .A1(n3419), .A2(n3418), .ZN(n3422) );
  XNOR2_X1 U4215 ( .A(n3420), .B(n3422), .ZN(n3464) );
  INV_X1 U4216 ( .A(n3420), .ZN(n3421) );
  AOI22_X1 U4217 ( .A1(n3465), .A2(n3464), .B1(n3422), .B2(n3421), .ZN(n3431)
         );
  OAI22_X1 U4218 ( .A1(n3853), .A2(n3424), .B1(n3836), .B2(n2862), .ZN(n3426)
         );
  XNOR2_X1 U4219 ( .A(n3426), .B(n3425), .ZN(n3429) );
  OAI22_X1 U4220 ( .A1(n3853), .A2(n2862), .B1(n3836), .B2(n3427), .ZN(n3428)
         );
  XNOR2_X1 U4221 ( .A(n3429), .B(n3428), .ZN(n3430) );
  XNOR2_X1 U4222 ( .A(n3431), .B(n3430), .ZN(n3437) );
  INV_X1 U4223 ( .A(n3439), .ZN(n3435) );
  INV_X1 U4224 ( .A(REG3_REG_28__SCAN_IN), .ZN(n3432) );
  OAI22_X1 U4225 ( .A1(n4349), .A2(n3836), .B1(STATE_REG_SCAN_IN), .B2(n3432), 
        .ZN(n3434) );
  OAI22_X1 U4226 ( .A1(n3575), .A2(n4343), .B1(n3702), .B2(n4344), .ZN(n3433)
         );
  AOI211_X1 U4227 ( .C1(n3435), .C2(n3578), .A(n3434), .B(n3433), .ZN(n3436)
         );
  OAI21_X1 U4228 ( .B1(n3437), .B2(n3581), .A(n3436), .ZN(U3217) );
  OAI22_X1 U4229 ( .A1(n3439), .A2(n3950), .B1(n3438), .B2(n4027), .ZN(n3440)
         );
  AOI21_X1 U4230 ( .B1(n3441), .B2(n3911), .A(n3440), .ZN(n3442) );
  OAI21_X1 U4231 ( .B1(n3443), .B2(n4006), .A(n3442), .ZN(n3444) );
  AOI21_X1 U4232 ( .B1(n3445), .B2(n4027), .A(n3444), .ZN(n3446) );
  OAI21_X1 U4233 ( .B1(n3447), .B2(n4070), .A(n3446), .ZN(U3262) );
  NAND3_X1 U4234 ( .A1(n3449), .A2(IR_REG_31__SCAN_IN), .A3(STATE_REG_SCAN_IN), 
        .ZN(n3451) );
  INV_X1 U4235 ( .A(DATAI_31_), .ZN(n3450) );
  OAI22_X1 U4236 ( .A1(n3448), .A2(n3451), .B1(STATE_REG_SCAN_IN), .B2(n3450), 
        .ZN(U3321) );
  NOR2_X1 U4237 ( .A1(n3452), .A2(n2593), .ZN(n3453) );
  AOI22_X1 U4238 ( .A1(n4517), .A2(n3454), .B1(n3453), .B2(n2591), .ZN(U3458)
         );
  INV_X1 U4239 ( .A(n3456), .ZN(n3457) );
  AOI21_X1 U4240 ( .B1(n3455), .B2(n3458), .A(n3457), .ZN(n3463) );
  AOI22_X1 U4241 ( .A1(n3475), .A2(n3761), .B1(n3589), .B2(n3459), .ZN(n3462)
         );
  AOI22_X1 U4242 ( .A1(REG3_REG_2__SCAN_IN), .A2(n3460), .B1(n3476), .B2(n3763), .ZN(n3461) );
  OAI211_X1 U4243 ( .C1(n3463), .C2(n3581), .A(n3462), .B(n3461), .ZN(U3234)
         );
  XNOR2_X1 U4244 ( .A(n3465), .B(n3464), .ZN(n3470) );
  OAI22_X1 U4245 ( .A1(n4349), .A2(n4087), .B1(STATE_REG_SCAN_IN), .B2(n3466), 
        .ZN(n3468) );
  OAI22_X1 U4246 ( .A1(n3853), .A2(n4344), .B1(n3852), .B2(n4343), .ZN(n3467)
         );
  AOI211_X1 U4247 ( .C1(n3854), .C2(n3578), .A(n3468), .B(n3467), .ZN(n3469)
         );
  OAI21_X1 U4248 ( .B1(n3470), .B2(n3581), .A(n3469), .ZN(U3211) );
  OAI21_X1 U4249 ( .B1(n3471), .B2(n3473), .A(n3472), .ZN(n3474) );
  NAND3_X1 U4250 ( .A1(n2158), .A2(n4357), .A3(n3474), .ZN(n3481) );
  AOI22_X1 U4251 ( .A1(n3589), .A2(n3605), .B1(REG3_REG_23__SCAN_IN), .B2(
        U3149), .ZN(n3480) );
  AOI22_X1 U4252 ( .A1(n3476), .A2(n3967), .B1(n3475), .B2(n3928), .ZN(n3479)
         );
  INV_X1 U4253 ( .A(n3934), .ZN(n3477) );
  NAND2_X1 U4254 ( .A1(n3578), .A2(n3477), .ZN(n3478) );
  NAND4_X1 U4255 ( .A1(n3481), .A2(n3480), .A3(n3479), .A4(n3478), .ZN(U3213)
         );
  OAI21_X1 U4256 ( .B1(n3483), .B2(n3482), .A(n2840), .ZN(n3484) );
  NAND2_X1 U4257 ( .A1(n3484), .A2(n4357), .ZN(n3493) );
  OAI22_X1 U4258 ( .A1(n4344), .A2(n3486), .B1(n4349), .B2(n3485), .ZN(n3489)
         );
  NOR2_X1 U4259 ( .A1(n4343), .A2(n3487), .ZN(n3488) );
  NOR2_X1 U4260 ( .A1(n3489), .A2(n3488), .ZN(n3492) );
  MUX2_X1 U4261 ( .A(STATE_REG_SCAN_IN), .B(n4362), .S(n3490), .Z(n3491) );
  NAND3_X1 U4262 ( .A1(n3493), .A2(n3492), .A3(n3491), .ZN(U3215) );
  OAI21_X1 U4263 ( .B1(n3496), .B2(n3494), .A(n3495), .ZN(n3497) );
  NAND2_X1 U4264 ( .A1(n3497), .A2(n4357), .ZN(n3501) );
  NAND2_X1 U4265 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n3821) );
  INV_X1 U4266 ( .A(n3821), .ZN(n3499) );
  OAI22_X1 U4267 ( .A1(n3529), .A2(n4343), .B1(n4344), .B2(n3995), .ZN(n3498)
         );
  AOI211_X1 U4268 ( .C1(n3607), .C2(n3589), .A(n3499), .B(n3498), .ZN(n3500)
         );
  OAI211_X1 U4269 ( .C1(n4362), .C2(n3502), .A(n3501), .B(n3500), .ZN(U3216)
         );
  INV_X1 U4270 ( .A(n3503), .ZN(n3505) );
  NAND2_X1 U4271 ( .A1(n3505), .A2(n3504), .ZN(n3509) );
  INV_X1 U4272 ( .A(n3546), .ZN(n3507) );
  OAI211_X1 U4273 ( .C1(n3506), .C2(n3507), .A(n3544), .B(n3509), .ZN(n3508)
         );
  OAI211_X1 U4274 ( .C1(n3510), .C2(n3509), .A(n4357), .B(n3508), .ZN(n3515)
         );
  OAI22_X1 U4275 ( .A1(n4349), .A2(n3963), .B1(STATE_REG_SCAN_IN), .B2(n3511), 
        .ZN(n3513) );
  OAI22_X1 U4276 ( .A1(n3926), .A2(n4344), .B1(n4343), .B2(n3995), .ZN(n3512)
         );
  AOI211_X1 U4277 ( .C1(n3961), .C2(n3578), .A(n3513), .B(n3512), .ZN(n3514)
         );
  NAND2_X1 U4278 ( .A1(n3515), .A2(n3514), .ZN(U3220) );
  NOR2_X1 U4279 ( .A1(n3517), .A2(n2148), .ZN(n3518) );
  XNOR2_X1 U4280 ( .A(n3519), .B(n3518), .ZN(n3524) );
  OAI22_X1 U4281 ( .A1(n4349), .A2(n3888), .B1(STATE_REG_SCAN_IN), .B2(n4096), 
        .ZN(n3522) );
  INV_X1 U4282 ( .A(n3928), .ZN(n3520) );
  OAI22_X1 U4283 ( .A1(n3852), .A2(n4344), .B1(n3520), .B2(n4343), .ZN(n3521)
         );
  AOI211_X1 U4284 ( .C1(n3889), .C2(n3578), .A(n3522), .B(n3521), .ZN(n3523)
         );
  OAI21_X1 U4285 ( .B1(n3524), .B2(n3581), .A(n3523), .ZN(U3222) );
  XNOR2_X1 U4286 ( .A(n3526), .B(n3525), .ZN(n3527) );
  XNOR2_X1 U4287 ( .A(n3528), .B(n3527), .ZN(n3533) );
  INV_X1 U4288 ( .A(REG3_REG_17__SCAN_IN), .ZN(n4181) );
  NOR2_X1 U4289 ( .A1(STATE_REG_SCAN_IN), .A2(n4181), .ZN(n4461) );
  OAI22_X1 U4290 ( .A1(n3586), .A2(n4343), .B1(n4344), .B2(n3529), .ZN(n3530)
         );
  AOI211_X1 U4291 ( .C1(n4042), .C2(n3589), .A(n4461), .B(n3530), .ZN(n3532)
         );
  NAND2_X1 U4292 ( .A1(n3578), .A2(n4041), .ZN(n3531) );
  OAI211_X1 U4293 ( .C1(n3533), .C2(n3581), .A(n3532), .B(n3531), .ZN(U3225)
         );
  NAND2_X1 U4294 ( .A1(n2016), .A2(n3534), .ZN(n3536) );
  XNOR2_X1 U4295 ( .A(n3536), .B(n3535), .ZN(n3542) );
  INV_X1 U4296 ( .A(n3905), .ZN(n3540) );
  OAI22_X1 U4297 ( .A1(n4349), .A2(n4236), .B1(STATE_REG_SCAN_IN), .B2(n3537), 
        .ZN(n3539) );
  OAI22_X1 U4298 ( .A1(n3865), .A2(n4344), .B1(n3900), .B2(n4343), .ZN(n3538)
         );
  AOI211_X1 U4299 ( .C1(n3540), .C2(n3578), .A(n3539), .B(n3538), .ZN(n3541)
         );
  OAI21_X1 U4300 ( .B1(n3542), .B2(n3581), .A(n3541), .ZN(U3226) );
  INV_X1 U4301 ( .A(n3543), .ZN(n3547) );
  AOI21_X1 U4302 ( .B1(n3544), .B2(n3546), .A(n3506), .ZN(n3545) );
  AOI21_X1 U4303 ( .B1(n3547), .B2(n3546), .A(n3545), .ZN(n3552) );
  INV_X1 U4304 ( .A(REG3_REG_20__SCAN_IN), .ZN(n3548) );
  OAI22_X1 U4305 ( .A1(n4349), .A2(n4256), .B1(STATE_REG_SCAN_IN), .B2(n3548), 
        .ZN(n3550) );
  OAI22_X1 U4306 ( .A1(n3565), .A2(n4343), .B1(n4344), .B2(n3974), .ZN(n3549)
         );
  AOI211_X1 U4307 ( .C1(n3980), .C2(n3578), .A(n3550), .B(n3549), .ZN(n3551)
         );
  OAI21_X1 U4308 ( .B1(n3552), .B2(n3581), .A(n3551), .ZN(U3230) );
  AOI21_X1 U4309 ( .B1(n3554), .B2(n3553), .A(n3471), .ZN(n3559) );
  INV_X1 U4310 ( .A(n3951), .ZN(n3557) );
  OAI22_X1 U4311 ( .A1(n4349), .A2(n3947), .B1(STATE_REG_SCAN_IN), .B2(n4196), 
        .ZN(n3556) );
  OAI22_X1 U4312 ( .A1(n3900), .A2(n4344), .B1(n4343), .B2(n3974), .ZN(n3555)
         );
  AOI211_X1 U4313 ( .C1(n3557), .C2(n3578), .A(n3556), .B(n3555), .ZN(n3558)
         );
  OAI21_X1 U4314 ( .B1(n3559), .B2(n3581), .A(n3558), .ZN(U3232) );
  INV_X1 U4315 ( .A(n3560), .ZN(n3561) );
  NOR2_X1 U4316 ( .A1(n3562), .A2(n3561), .ZN(n3563) );
  XNOR2_X1 U4317 ( .A(n3564), .B(n3563), .ZN(n3569) );
  NOR2_X1 U4318 ( .A1(STATE_REG_SCAN_IN), .A2(n4202), .ZN(n4486) );
  OAI22_X1 U4319 ( .A1(n3565), .A2(n4344), .B1(n4343), .B2(n4345), .ZN(n3566)
         );
  AOI211_X1 U4320 ( .C1(n4015), .C2(n3589), .A(n4486), .B(n3566), .ZN(n3568)
         );
  NAND2_X1 U4321 ( .A1(n3578), .A2(n4023), .ZN(n3567) );
  OAI211_X1 U4322 ( .C1(n3569), .C2(n3581), .A(n3568), .B(n3567), .ZN(U3235)
         );
  INV_X1 U4323 ( .A(n3570), .ZN(n3572) );
  NAND2_X1 U4324 ( .A1(n3572), .A2(n3571), .ZN(n3573) );
  XNOR2_X1 U4325 ( .A(n3574), .B(n3573), .ZN(n3582) );
  INV_X1 U4326 ( .A(n3874), .ZN(n3579) );
  OAI22_X1 U4327 ( .A1(n4349), .A2(n3872), .B1(STATE_REG_SCAN_IN), .B2(n4094), 
        .ZN(n3577) );
  OAI22_X1 U4328 ( .A1(n3575), .A2(n4344), .B1(n3865), .B2(n4343), .ZN(n3576)
         );
  AOI211_X1 U4329 ( .C1(n3579), .C2(n3578), .A(n3577), .B(n3576), .ZN(n3580)
         );
  OAI21_X1 U4330 ( .B1(n3582), .B2(n3581), .A(n3580), .ZN(U3237) );
  INV_X1 U4331 ( .A(n4353), .ZN(n3583) );
  NOR2_X1 U4332 ( .A1(n4352), .A2(n3583), .ZN(n3584) );
  XNOR2_X1 U4333 ( .A(n3584), .B(n4354), .ZN(n3585) );
  NAND2_X1 U4334 ( .A1(n3585), .A2(n4357), .ZN(n3591) );
  AND2_X1 U4335 ( .A1(U3149), .A2(REG3_REG_15__SCAN_IN), .ZN(n4445) );
  OAI22_X1 U4336 ( .A1(n3587), .A2(n4343), .B1(n4344), .B2(n3586), .ZN(n3588)
         );
  AOI211_X1 U4337 ( .C1(n4278), .C2(n3589), .A(n4445), .B(n3588), .ZN(n3590)
         );
  OAI211_X1 U4338 ( .C1(n4362), .C2(n3592), .A(n3591), .B(n3590), .ZN(U3238)
         );
  INV_X1 U4339 ( .A(n3942), .ZN(n3593) );
  NAND2_X1 U4340 ( .A1(n3593), .A2(n4059), .ZN(n3601) );
  NAND4_X1 U4341 ( .A1(n3597), .A2(n3596), .A3(n3595), .A4(n3594), .ZN(n3600)
         );
  NOR4_X1 U4342 ( .A1(n3601), .A2(n3600), .A3(n3599), .A4(n3598), .ZN(n3626)
         );
  NOR2_X1 U4343 ( .A1(n3602), .A2(n2027), .ZN(n3863) );
  NOR2_X1 U4344 ( .A1(n3862), .A2(n3694), .ZN(n3880) );
  INV_X1 U4345 ( .A(n3603), .ZN(n3693) );
  OR2_X1 U4346 ( .A1(n3693), .A2(n3604), .ZN(n3903) );
  INV_X1 U4347 ( .A(n3903), .ZN(n3896) );
  XNOR2_X1 U4348 ( .A(n3944), .B(n3605), .ZN(n3925) );
  NAND4_X1 U4349 ( .A1(n3863), .A2(n3880), .A3(n3896), .A4(n3925), .ZN(n3618)
         );
  INV_X1 U4350 ( .A(n3606), .ZN(n3922) );
  NOR2_X1 U4351 ( .A1(n3692), .A2(n3922), .ZN(n3964) );
  XNOR2_X1 U4352 ( .A(n4016), .B(n3607), .ZN(n3992) );
  INV_X1 U4353 ( .A(n3988), .ZN(n3608) );
  AND2_X1 U4354 ( .A1(n3608), .A2(n3987), .ZN(n4031) );
  XNOR2_X1 U4355 ( .A(n3966), .B(n3609), .ZN(n3977) );
  NAND4_X1 U4356 ( .A1(n3964), .A2(n3992), .A3(n4031), .A4(n3977), .ZN(n3617)
         );
  NAND2_X1 U4357 ( .A1(n2462), .A2(DATAI_29_), .ZN(n4083) );
  XNOR2_X1 U4358 ( .A(n3702), .B(n4083), .ZN(n3839) );
  AND2_X1 U4359 ( .A1(n2462), .A2(DATAI_30_), .ZN(n4080) );
  NAND2_X1 U4360 ( .A1(n3610), .A2(REG1_REG_31__SCAN_IN), .ZN(n3615) );
  NAND2_X1 U4361 ( .A1(n3611), .A2(REG0_REG_31__SCAN_IN), .ZN(n3614) );
  INV_X1 U4362 ( .A(REG2_REG_31__SCAN_IN), .ZN(n3612) );
  OR2_X1 U4363 ( .A1(n2008), .A2(n3612), .ZN(n3613) );
  AND3_X1 U4364 ( .A1(n3615), .A2(n3614), .A3(n3613), .ZN(n4073) );
  NAND2_X1 U4365 ( .A1(n2462), .A2(DATAI_31_), .ZN(n4071) );
  INV_X1 U4366 ( .A(n4071), .ZN(n4074) );
  NOR2_X1 U4367 ( .A1(n4073), .A2(n4074), .ZN(n3707) );
  AOI21_X1 U4368 ( .B1(n3833), .B2(n4080), .A(n3707), .ZN(n3700) );
  NOR2_X1 U4369 ( .A1(n3833), .A2(n4080), .ZN(n3737) );
  AOI21_X1 U4370 ( .B1(n4073), .B2(n4074), .A(n3737), .ZN(n3706) );
  NAND4_X1 U4371 ( .A1(n3839), .A2(n3837), .A3(n3700), .A4(n3706), .ZN(n3616)
         );
  NOR4_X1 U4372 ( .A1(n4014), .A2(n3622), .A3(n3621), .A4(n3620), .ZN(n3623)
         );
  NAND4_X1 U4373 ( .A1(n3626), .A2(n3625), .A3(n3624), .A4(n3623), .ZN(n3632)
         );
  NAND4_X1 U4374 ( .A1(n3629), .A2(n2076), .A3(n3628), .A4(n3627), .ZN(n3630)
         );
  NOR2_X1 U4375 ( .A1(n3633), .A2(n3643), .ZN(n3710) );
  NAND2_X1 U4376 ( .A1(n3635), .A2(n3634), .ZN(n3664) );
  NAND2_X1 U4377 ( .A1(n3664), .A2(n3636), .ZN(n3717) );
  NAND2_X1 U4378 ( .A1(n3637), .A2(n3636), .ZN(n3718) );
  INV_X1 U4379 ( .A(n3718), .ZN(n3638) );
  NAND2_X1 U4380 ( .A1(n3639), .A2(n3638), .ZN(n3682) );
  OAI211_X1 U4381 ( .C1(n2084), .C2(n3643), .A(n3642), .B(n3641), .ZN(n3645)
         );
  NAND3_X1 U4382 ( .A1(n3645), .A2(n3644), .A3(n2545), .ZN(n3648) );
  NAND3_X1 U4383 ( .A1(n3648), .A2(n3647), .A3(n3646), .ZN(n3651) );
  NAND3_X1 U4384 ( .A1(n3651), .A2(n3650), .A3(n3649), .ZN(n3654) );
  NAND4_X1 U4385 ( .A1(n3654), .A2(n3653), .A3(n3652), .A4(n3667), .ZN(n3657)
         );
  INV_X1 U4386 ( .A(n3655), .ZN(n3666) );
  AOI21_X1 U4387 ( .B1(n3657), .B2(n3656), .A(n3666), .ZN(n3659) );
  OAI21_X1 U4388 ( .B1(n3659), .B2(n3658), .A(n3668), .ZN(n3662) );
  NAND3_X1 U4389 ( .A1(n3662), .A2(n3661), .A3(n3660), .ZN(n3675) );
  NOR2_X1 U4390 ( .A1(n3664), .A2(n3663), .ZN(n3674) );
  NOR2_X1 U4391 ( .A1(n3666), .A2(n3665), .ZN(n3670) );
  NAND4_X1 U4392 ( .A1(n3670), .A2(n3669), .A3(n3668), .A4(n3667), .ZN(n3672)
         );
  NAND2_X1 U4393 ( .A1(n3672), .A2(n3671), .ZN(n3673) );
  AOI22_X1 U4394 ( .A1(n3675), .A2(n3674), .B1(n3717), .B2(n3673), .ZN(n3680)
         );
  INV_X1 U4395 ( .A(n3676), .ZN(n3678) );
  NOR4_X1 U4396 ( .A1(n3680), .A2(n3679), .A3(n3678), .A4(n3677), .ZN(n3681)
         );
  AOI21_X1 U4397 ( .B1(n3717), .B2(n3682), .A(n3681), .ZN(n3684) );
  INV_X1 U4398 ( .A(n3683), .ZN(n3720) );
  OAI21_X1 U4399 ( .B1(n3684), .B2(n3720), .A(n3722), .ZN(n3688) );
  INV_X1 U4400 ( .A(n3685), .ZN(n3686) );
  AOI21_X1 U4401 ( .B1(n3688), .B2(n3687), .A(n3686), .ZN(n3690) );
  AOI221_X1 U4402 ( .B1(n3692), .B2(n3691), .C1(n3690), .C2(n3691), .A(n3689), 
        .ZN(n3696) );
  NOR2_X1 U4403 ( .A1(n3694), .A2(n3693), .ZN(n3716) );
  OAI21_X1 U4404 ( .B1(n3696), .B2(n3695), .A(n3716), .ZN(n3698) );
  INV_X1 U4405 ( .A(n4083), .ZN(n3703) );
  OAI21_X1 U4406 ( .B1(n3703), .B2(n3702), .A(n3828), .ZN(n3704) );
  OR2_X1 U4407 ( .A1(n3704), .A2(n2027), .ZN(n3711) );
  AOI211_X1 U4408 ( .C1(n3727), .C2(n3698), .A(n3697), .B(n3711), .ZN(n3708)
         );
  INV_X1 U4409 ( .A(n3699), .ZN(n3827) );
  NOR2_X1 U4410 ( .A1(n3827), .A2(n3732), .ZN(n3705) );
  INV_X1 U4411 ( .A(n3700), .ZN(n3701) );
  AOI21_X1 U4412 ( .B1(n3703), .B2(n3702), .A(n3701), .ZN(n3715) );
  OAI21_X1 U4413 ( .B1(n3705), .B2(n3704), .A(n3715), .ZN(n3712) );
  OAI22_X1 U4414 ( .A1(n3708), .A2(n3712), .B1(n3707), .B2(n3706), .ZN(n3709)
         );
  MUX2_X1 U4415 ( .A(n3710), .B(n3709), .S(n2576), .Z(n3742) );
  INV_X1 U4416 ( .A(n3711), .ZN(n3714) );
  INV_X1 U4417 ( .A(n3850), .ZN(n3713) );
  AOI21_X1 U4418 ( .B1(n3714), .B2(n3713), .A(n3712), .ZN(n3736) );
  INV_X1 U4419 ( .A(n3715), .ZN(n3733) );
  INV_X1 U4420 ( .A(n3716), .ZN(n3730) );
  OAI21_X1 U4421 ( .B1(n3719), .B2(n3718), .A(n3717), .ZN(n3721) );
  AOI21_X1 U4422 ( .B1(n3722), .B2(n3721), .A(n3720), .ZN(n3726) );
  INV_X1 U4423 ( .A(n3723), .ZN(n3724) );
  OAI21_X1 U4424 ( .B1(n3726), .B2(n3725), .A(n3724), .ZN(n3728) );
  OAI221_X1 U4425 ( .B1(n3730), .B2(n3729), .C1(n3730), .C2(n3728), .A(n3727), 
        .ZN(n3731) );
  NOR4_X1 U4426 ( .A1(n3733), .A2(n3827), .A3(n3732), .A4(n3731), .ZN(n3735)
         );
  INV_X1 U4427 ( .A(n4073), .ZN(n3751) );
  INV_X1 U4428 ( .A(n4080), .ZN(n3734) );
  OAI22_X1 U4429 ( .A1(n3736), .A2(n3735), .B1(n3751), .B2(n3734), .ZN(n3740)
         );
  OAI21_X1 U4430 ( .B1(n3737), .B2(n4073), .A(n4074), .ZN(n3739) );
  AOI21_X1 U4431 ( .B1(n3740), .B2(n3739), .A(n3738), .ZN(n3741) );
  NOR2_X1 U4432 ( .A1(n3742), .A2(n3741), .ZN(n3743) );
  XNOR2_X1 U4433 ( .A(n3743), .B(n4334), .ZN(n3750) );
  NAND2_X1 U4434 ( .A1(n3745), .A2(n3744), .ZN(n3746) );
  OAI211_X1 U4435 ( .C1(n3747), .C2(n3749), .A(n3746), .B(B_REG_SCAN_IN), .ZN(
        n3748) );
  OAI21_X1 U4436 ( .B1(n3750), .B2(n3749), .A(n3748), .ZN(U3239) );
  MUX2_X1 U4437 ( .A(n3751), .B(DATAO_REG_31__SCAN_IN), .S(n3762), .Z(U3581)
         );
  MUX2_X1 U4438 ( .A(DATAO_REG_27__SCAN_IN), .B(n3867), .S(n3775), .Z(U3577)
         );
  MUX2_X1 U4439 ( .A(DATAO_REG_26__SCAN_IN), .B(n3883), .S(n3775), .Z(U3576)
         );
  MUX2_X1 U4440 ( .A(n3898), .B(DATAO_REG_25__SCAN_IN), .S(n3762), .Z(U3575)
         );
  MUX2_X1 U4441 ( .A(n3928), .B(DATAO_REG_24__SCAN_IN), .S(n3762), .Z(U3574)
         );
  MUX2_X1 U4442 ( .A(n3944), .B(DATAO_REG_23__SCAN_IN), .S(n3762), .Z(U3573)
         );
  MUX2_X1 U4443 ( .A(DATAO_REG_22__SCAN_IN), .B(n3967), .S(n3775), .Z(U3572)
         );
  MUX2_X1 U4444 ( .A(DATAO_REG_21__SCAN_IN), .B(n3752), .S(n3775), .Z(U3571)
         );
  MUX2_X1 U4445 ( .A(n4016), .B(DATAO_REG_19__SCAN_IN), .S(n3762), .Z(U3569)
         );
  MUX2_X1 U4446 ( .A(n4035), .B(DATAO_REG_18__SCAN_IN), .S(n3762), .Z(U3568)
         );
  MUX2_X1 U4447 ( .A(n4063), .B(DATAO_REG_17__SCAN_IN), .S(n3762), .Z(U3567)
         );
  MUX2_X1 U4448 ( .A(n4034), .B(DATAO_REG_16__SCAN_IN), .S(n3762), .Z(U3566)
         );
  MUX2_X1 U4449 ( .A(n3753), .B(DATAO_REG_13__SCAN_IN), .S(n3762), .Z(U3563)
         );
  MUX2_X1 U4450 ( .A(n3754), .B(DATAO_REG_12__SCAN_IN), .S(n3762), .Z(U3562)
         );
  MUX2_X1 U4451 ( .A(n3755), .B(DATAO_REG_11__SCAN_IN), .S(n3762), .Z(U3561)
         );
  MUX2_X1 U4452 ( .A(n3756), .B(DATAO_REG_9__SCAN_IN), .S(n3762), .Z(U3559) );
  MUX2_X1 U4453 ( .A(n3757), .B(DATAO_REG_8__SCAN_IN), .S(n3762), .Z(U3558) );
  MUX2_X1 U4454 ( .A(n3758), .B(DATAO_REG_6__SCAN_IN), .S(n3762), .Z(U3556) );
  MUX2_X1 U4455 ( .A(n3759), .B(DATAO_REG_5__SCAN_IN), .S(n3762), .Z(U3555) );
  MUX2_X1 U4456 ( .A(n3760), .B(DATAO_REG_4__SCAN_IN), .S(n3762), .Z(U3554) );
  MUX2_X1 U4457 ( .A(n3761), .B(DATAO_REG_3__SCAN_IN), .S(n3762), .Z(U3553) );
  MUX2_X1 U4458 ( .A(n2789), .B(DATAO_REG_2__SCAN_IN), .S(n3762), .Z(U3552) );
  MUX2_X1 U4459 ( .A(n3763), .B(DATAO_REG_1__SCAN_IN), .S(n3762), .Z(U3551) );
  AOI22_X1 U4460 ( .A1(n4462), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n3770) );
  OAI211_X1 U4461 ( .C1(n3765), .C2(n3764), .A(n4470), .B(n3787), .ZN(n3769)
         );
  OAI211_X1 U4462 ( .C1(n3774), .C2(n3766), .A(n4472), .B(n3779), .ZN(n3768)
         );
  NAND2_X1 U4463 ( .A1(n4484), .A2(n4339), .ZN(n3767) );
  NAND4_X1 U4464 ( .A1(n3770), .A2(n3769), .A3(n3768), .A4(n3767), .ZN(U3241)
         );
  NAND2_X1 U4465 ( .A1(n3771), .A2(n3832), .ZN(n3773) );
  OAI211_X1 U4466 ( .C1(n3774), .C2(n3832), .A(n3773), .B(n3772), .ZN(n3776)
         );
  OAI211_X1 U4467 ( .C1(IR_REG_0__SCAN_IN), .C2(n3777), .A(n3776), .B(n3775), 
        .ZN(n4382) );
  AOI22_X1 U4468 ( .A1(ADDR_REG_2__SCAN_IN), .A2(n4462), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n3793) );
  MUX2_X1 U4469 ( .A(n2668), .B(REG2_REG_2__SCAN_IN), .S(n4338), .Z(n3780) );
  NAND3_X1 U4470 ( .A1(n3780), .A2(n3779), .A3(n3778), .ZN(n3782) );
  NAND3_X1 U4471 ( .A1(n4472), .A2(n3782), .A3(n3781), .ZN(n3784) );
  NAND2_X1 U4472 ( .A1(n4484), .A2(n4338), .ZN(n3783) );
  AND2_X1 U4473 ( .A1(n3784), .A2(n3783), .ZN(n3792) );
  MUX2_X1 U4474 ( .A(n3785), .B(REG1_REG_2__SCAN_IN), .S(n4338), .Z(n3788) );
  NAND3_X1 U4475 ( .A1(n3788), .A2(n3787), .A3(n3786), .ZN(n3789) );
  NAND3_X1 U4476 ( .A1(n4470), .A2(n3790), .A3(n3789), .ZN(n3791) );
  NAND4_X1 U4477 ( .A1(n4382), .A2(n3793), .A3(n3792), .A4(n3791), .ZN(U3242)
         );
  INV_X1 U4478 ( .A(REG1_REG_18__SCAN_IN), .ZN(n3794) );
  INV_X1 U4479 ( .A(n4483), .ZN(n4521) );
  AOI22_X1 U4480 ( .A1(n4483), .A2(n3794), .B1(REG1_REG_18__SCAN_IN), .B2(
        n4521), .ZN(n4477) );
  INV_X1 U4481 ( .A(REG1_REG_17__SCAN_IN), .ZN(n3795) );
  AOI22_X1 U4482 ( .A1(n3817), .A2(REG1_REG_17__SCAN_IN), .B1(n3795), .B2(
        n4522), .ZN(n4468) );
  NOR2_X1 U4483 ( .A1(n3799), .A2(n3798), .ZN(n3800) );
  INV_X1 U4484 ( .A(REG1_REG_14__SCAN_IN), .ZN(n4432) );
  INV_X1 U4485 ( .A(n3814), .ZN(n4526) );
  INV_X1 U4486 ( .A(REG1_REG_15__SCAN_IN), .ZN(n3801) );
  AOI22_X1 U4487 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4526), .B1(n3814), .B2(
        n3801), .ZN(n4447) );
  NAND2_X1 U4488 ( .A1(n3803), .A2(n4524), .ZN(n3804) );
  INV_X1 U4489 ( .A(REG1_REG_16__SCAN_IN), .ZN(n4455) );
  NAND2_X1 U4490 ( .A1(n4456), .A2(n4455), .ZN(n4454) );
  NAND2_X1 U4491 ( .A1(n3804), .A2(n4454), .ZN(n4467) );
  XNOR2_X1 U4492 ( .A(n4334), .B(REG1_REG_19__SCAN_IN), .ZN(n3805) );
  XNOR2_X1 U4493 ( .A(n3806), .B(n3805), .ZN(n3826) );
  NAND2_X1 U4494 ( .A1(n4483), .A2(REG2_REG_18__SCAN_IN), .ZN(n3807) );
  OAI21_X1 U4495 ( .B1(n4483), .B2(REG2_REG_18__SCAN_IN), .A(n3807), .ZN(n4482) );
  NOR2_X1 U4496 ( .A1(n3817), .A2(REG2_REG_17__SCAN_IN), .ZN(n3808) );
  AOI21_X1 U4497 ( .B1(REG2_REG_17__SCAN_IN), .B2(n3817), .A(n3808), .ZN(n4465) );
  NOR2_X1 U4498 ( .A1(n3798), .A2(n3812), .ZN(n3813) );
  XOR2_X1 U4499 ( .A(n4437), .B(n3812), .Z(n4434) );
  NOR2_X1 U4500 ( .A1(n2261), .A2(n4434), .ZN(n4433) );
  AOI22_X1 U4501 ( .A1(REG2_REG_15__SCAN_IN), .A2(n4526), .B1(n3814), .B2(
        n2406), .ZN(n4442) );
  NAND2_X1 U4502 ( .A1(n3815), .A2(n4524), .ZN(n3816) );
  NAND2_X1 U4503 ( .A1(n4453), .A2(n2417), .ZN(n4452) );
  NAND2_X1 U4504 ( .A1(n3816), .A2(n4452), .ZN(n4464) );
  NAND2_X1 U4505 ( .A1(n4465), .A2(n4464), .ZN(n4463) );
  OAI21_X1 U4506 ( .B1(n3817), .B2(REG2_REG_17__SCAN_IN), .A(n4463), .ZN(n4481) );
  NOR2_X1 U4507 ( .A1(n4482), .A2(n4481), .ZN(n4480) );
  AOI21_X1 U4508 ( .B1(REG2_REG_18__SCAN_IN), .B2(n4483), .A(n4480), .ZN(n3819) );
  MUX2_X1 U4509 ( .A(REG2_REG_19__SCAN_IN), .B(n2452), .S(n4334), .Z(n3818) );
  XNOR2_X1 U4510 ( .A(n3819), .B(n3818), .ZN(n3824) );
  NAND2_X1 U4511 ( .A1(n4462), .A2(ADDR_REG_19__SCAN_IN), .ZN(n3820) );
  OAI211_X1 U4512 ( .C1(n4475), .C2(n3822), .A(n3821), .B(n3820), .ZN(n3823)
         );
  AOI21_X1 U4513 ( .B1(n3824), .B2(n4472), .A(n3823), .ZN(n3825) );
  OAI21_X1 U4514 ( .B1(n3826), .B2(n4476), .A(n3825), .ZN(U3259) );
  AOI21_X1 U4515 ( .B1(n3829), .B2(n3828), .A(n3827), .ZN(n3830) );
  XNOR2_X1 U4516 ( .A(n3830), .B(n3839), .ZN(n3834) );
  INV_X1 U4517 ( .A(B_REG_SCAN_IN), .ZN(n3831) );
  OAI21_X1 U4518 ( .B1(n3832), .B2(n3831), .A(n4064), .ZN(n4072) );
  OAI222_X1 U4519 ( .A1(n4018), .A2(n3853), .B1(n3834), .B2(n3998), .C1(n4072), 
        .C2(n3833), .ZN(n4085) );
  AOI21_X1 U4520 ( .B1(n3835), .B2(n4497), .A(n4085), .ZN(n3847) );
  OAI22_X1 U4521 ( .A1(n3838), .A2(n3837), .B1(n3853), .B2(n3836), .ZN(n3840)
         );
  XNOR2_X1 U4522 ( .A(n3840), .B(n3839), .ZN(n4082) );
  NAND2_X1 U4523 ( .A1(n4082), .A2(n3979), .ZN(n3846) );
  INV_X1 U4524 ( .A(n4084), .ZN(n3844) );
  OAI22_X1 U4525 ( .A1(n4083), .A2(n4056), .B1(n4027), .B2(n3842), .ZN(n3843)
         );
  AOI21_X1 U4526 ( .B1(n3844), .B2(n4501), .A(n3843), .ZN(n3845) );
  OAI211_X1 U4527 ( .C1(n4507), .C2(n3847), .A(n3846), .B(n3845), .ZN(U3354)
         );
  XNOR2_X1 U4528 ( .A(n3848), .B(n3850), .ZN(n4091) );
  INV_X1 U4529 ( .A(n4091), .ZN(n3860) );
  XOR2_X1 U4530 ( .A(n3850), .B(n3849), .Z(n3851) );
  OAI222_X1 U4531 ( .A1(n3994), .A2(n3853), .B1(n4018), .B2(n3852), .C1(n3998), 
        .C2(n3851), .ZN(n4090) );
  XNOR2_X1 U4532 ( .A(n3870), .B(n4087), .ZN(n4088) );
  AOI22_X1 U4533 ( .A1(n3854), .A2(n4497), .B1(REG2_REG_27__SCAN_IN), .B2(
        n4363), .ZN(n3857) );
  NAND2_X1 U4534 ( .A1(n3911), .A2(n3855), .ZN(n3856) );
  OAI211_X1 U4535 ( .C1(n4088), .C2(n4006), .A(n3857), .B(n3856), .ZN(n3858)
         );
  AOI21_X1 U4536 ( .B1(n4090), .B2(n4027), .A(n3858), .ZN(n3859) );
  OAI21_X1 U4537 ( .B1(n3860), .B2(n4070), .A(n3859), .ZN(U3263) );
  XNOR2_X1 U4538 ( .A(n3861), .B(n3863), .ZN(n4228) );
  INV_X1 U4539 ( .A(n4228), .ZN(n3878) );
  NOR2_X1 U4540 ( .A1(n2036), .A2(n3862), .ZN(n3864) );
  XNOR2_X1 U4541 ( .A(n3864), .B(n3863), .ZN(n3869) );
  OAI22_X1 U4542 ( .A1(n3865), .A2(n4018), .B1(n3872), .B2(n4284), .ZN(n3866)
         );
  AOI21_X1 U4543 ( .B1(n3867), .B2(n4064), .A(n3866), .ZN(n3868) );
  OAI21_X1 U4544 ( .B1(n3869), .B2(n3998), .A(n3868), .ZN(n4227) );
  INV_X1 U4545 ( .A(n3870), .ZN(n3871) );
  OAI21_X1 U4546 ( .B1(n2097), .B2(n3872), .A(n3871), .ZN(n4302) );
  NOR2_X1 U4547 ( .A1(n4302), .A2(n4006), .ZN(n3876) );
  OAI22_X1 U4548 ( .A1(n3874), .A2(n3950), .B1(n3873), .B2(n4027), .ZN(n3875)
         );
  AOI211_X1 U4549 ( .C1(n4227), .C2(n4027), .A(n3876), .B(n3875), .ZN(n3877)
         );
  OAI21_X1 U4550 ( .B1(n3878), .B2(n4070), .A(n3877), .ZN(U3264) );
  XNOR2_X1 U4551 ( .A(n3879), .B(n3880), .ZN(n4232) );
  INV_X1 U4552 ( .A(n4232), .ZN(n3893) );
  XNOR2_X1 U4553 ( .A(n3881), .B(n3880), .ZN(n3886) );
  AOI22_X1 U4554 ( .A1(n3928), .A2(n4061), .B1(n3882), .B2(n4277), .ZN(n3885)
         );
  NAND2_X1 U4555 ( .A1(n3883), .A2(n4064), .ZN(n3884) );
  OAI211_X1 U4556 ( .C1(n3886), .C2(n3998), .A(n3885), .B(n3884), .ZN(n4231)
         );
  OAI21_X1 U4557 ( .B1(n2094), .B2(n3888), .A(n3887), .ZN(n4306) );
  AOI22_X1 U4558 ( .A1(n3889), .A2(n4497), .B1(n4363), .B2(
        REG2_REG_25__SCAN_IN), .ZN(n3890) );
  OAI21_X1 U4559 ( .B1(n4306), .B2(n4006), .A(n3890), .ZN(n3891) );
  AOI21_X1 U4560 ( .B1(n4231), .B2(n4027), .A(n3891), .ZN(n3892) );
  OAI21_X1 U4561 ( .B1(n3893), .B2(n4070), .A(n3892), .ZN(U3265) );
  OR2_X1 U4562 ( .A1(n3895), .A2(n3894), .ZN(n3897) );
  XNOR2_X1 U4563 ( .A(n3897), .B(n3896), .ZN(n3902) );
  NAND2_X1 U4564 ( .A1(n3898), .A2(n4064), .ZN(n3899) );
  OAI21_X1 U4565 ( .B1(n3900), .B2(n4018), .A(n3899), .ZN(n3901) );
  AOI21_X1 U4566 ( .B1(n3902), .B2(n4057), .A(n3901), .ZN(n4235) );
  XNOR2_X1 U4567 ( .A(n3904), .B(n3903), .ZN(n4238) );
  NAND2_X1 U4568 ( .A1(n4238), .A2(n3979), .ZN(n3913) );
  OAI22_X1 U4569 ( .A1(n4027), .A2(n3906), .B1(n3905), .B2(n3950), .ZN(n3909)
         );
  OAI21_X1 U4570 ( .B1(n3931), .B2(n4236), .A(n3907), .ZN(n4310) );
  NOR2_X1 U4571 ( .A1(n4310), .A2(n4006), .ZN(n3908) );
  AOI211_X1 U4572 ( .C1(n3911), .C2(n3910), .A(n3909), .B(n3908), .ZN(n3912)
         );
  OAI211_X1 U4573 ( .C1(n4507), .C2(n4235), .A(n3913), .B(n3912), .ZN(U3266)
         );
  XNOR2_X1 U4574 ( .A(n3914), .B(n3925), .ZN(n4242) );
  INV_X1 U4575 ( .A(n4242), .ZN(n3939) );
  INV_X1 U4576 ( .A(n3915), .ZN(n3916) );
  NAND2_X1 U4577 ( .A1(n3918), .A2(n3917), .ZN(n3972) );
  NAND2_X1 U4578 ( .A1(n3972), .A2(n3919), .ZN(n3921) );
  NAND2_X1 U4579 ( .A1(n3921), .A2(n3920), .ZN(n3965) );
  AOI21_X1 U4580 ( .B1(n3965), .B2(n3964), .A(n3922), .ZN(n3943) );
  OAI21_X1 U4581 ( .B1(n3943), .B2(n3942), .A(n3923), .ZN(n3924) );
  XOR2_X1 U4582 ( .A(n3925), .B(n3924), .Z(n3930) );
  OAI22_X1 U4583 ( .A1(n3926), .A2(n4018), .B1(n4284), .B2(n3933), .ZN(n3927)
         );
  AOI21_X1 U4584 ( .B1(n4064), .B2(n3928), .A(n3927), .ZN(n3929) );
  OAI21_X1 U4585 ( .B1(n3930), .B2(n3998), .A(n3929), .ZN(n4241) );
  INV_X1 U4586 ( .A(n3931), .ZN(n3932) );
  OAI21_X1 U4587 ( .B1(n2096), .B2(n3933), .A(n3932), .ZN(n4314) );
  NOR2_X1 U4588 ( .A1(n4314), .A2(n4006), .ZN(n3937) );
  OAI22_X1 U4589 ( .A1(n4027), .A2(n3935), .B1(n3934), .B2(n3950), .ZN(n3936)
         );
  AOI211_X1 U4590 ( .C1(n4241), .C2(n4027), .A(n3937), .B(n3936), .ZN(n3938)
         );
  OAI21_X1 U4591 ( .B1(n3939), .B2(n4070), .A(n3938), .ZN(U3267) );
  OAI21_X1 U4592 ( .B1(n3941), .B2(n3942), .A(n3940), .ZN(n4249) );
  XNOR2_X1 U4593 ( .A(n3943), .B(n3942), .ZN(n3949) );
  NAND2_X1 U4594 ( .A1(n3944), .A2(n4064), .ZN(n3946) );
  OR2_X1 U4595 ( .A1(n3974), .A2(n4018), .ZN(n3945) );
  OAI211_X1 U4596 ( .C1(n4284), .C2(n3947), .A(n3946), .B(n3945), .ZN(n3948)
         );
  AOI21_X1 U4597 ( .B1(n3949), .B2(n4057), .A(n3948), .ZN(n4248) );
  NOR2_X1 U4598 ( .A1(n3951), .A2(n3950), .ZN(n3952) );
  AOI21_X1 U4599 ( .B1(n4363), .B2(REG2_REG_22__SCAN_IN), .A(n3952), .ZN(n3955) );
  NAND2_X1 U4600 ( .A1(n3959), .A2(n3953), .ZN(n4245) );
  NAND3_X1 U4601 ( .A1(n4246), .A2(n4501), .A3(n4245), .ZN(n3954) );
  OAI211_X1 U4602 ( .C1(n4248), .C2(n4363), .A(n3955), .B(n3954), .ZN(n3956)
         );
  INV_X1 U4603 ( .A(n3956), .ZN(n3957) );
  OAI21_X1 U4604 ( .B1(n4249), .B2(n4070), .A(n3957), .ZN(U3268) );
  XNOR2_X1 U4605 ( .A(n3958), .B(n3964), .ZN(n4254) );
  INV_X1 U4606 ( .A(n3959), .ZN(n3960) );
  AOI21_X1 U4607 ( .B1(n4250), .B2(n2009), .A(n3960), .ZN(n4251) );
  AOI22_X1 U4608 ( .A1(n4507), .A2(REG2_REG_21__SCAN_IN), .B1(n3961), .B2(
        n4497), .ZN(n3962) );
  OAI21_X1 U4609 ( .B1(n4056), .B2(n3963), .A(n3962), .ZN(n3970) );
  XNOR2_X1 U4610 ( .A(n3965), .B(n3964), .ZN(n3968) );
  AOI222_X1 U4611 ( .A1(n4057), .A2(n3968), .B1(n3967), .B2(n4064), .C1(n3966), 
        .C2(n4061), .ZN(n4253) );
  NOR2_X1 U4612 ( .A1(n4253), .A2(n4363), .ZN(n3969) );
  AOI211_X1 U4613 ( .C1(n4251), .C2(n4501), .A(n3970), .B(n3969), .ZN(n3971)
         );
  OAI21_X1 U4614 ( .B1(n4254), .B2(n4070), .A(n3971), .ZN(U3269) );
  XNOR2_X1 U4615 ( .A(n3972), .B(n3977), .ZN(n3976) );
  NAND2_X1 U4616 ( .A1(n4016), .A2(n4061), .ZN(n3973) );
  OAI21_X1 U4617 ( .B1(n3974), .B2(n3994), .A(n3973), .ZN(n3975) );
  AOI21_X1 U4618 ( .B1(n3976), .B2(n4057), .A(n3975), .ZN(n4255) );
  XNOR2_X1 U4619 ( .A(n3978), .B(n3977), .ZN(n4258) );
  NAND2_X1 U4620 ( .A1(n4258), .A2(n3979), .ZN(n3985) );
  OAI21_X1 U4621 ( .B1(n4000), .B2(n4256), .A(n2009), .ZN(n4320) );
  INV_X1 U4622 ( .A(n4320), .ZN(n3983) );
  AOI22_X1 U4623 ( .A1(n4507), .A2(REG2_REG_20__SCAN_IN), .B1(n3980), .B2(
        n4497), .ZN(n3981) );
  OAI21_X1 U4624 ( .B1(n4056), .B2(n4256), .A(n3981), .ZN(n3982) );
  AOI21_X1 U4625 ( .B1(n3983), .B2(n4501), .A(n3982), .ZN(n3984) );
  OAI211_X1 U4626 ( .C1(n4507), .C2(n4255), .A(n3985), .B(n3984), .ZN(U3270)
         );
  XOR2_X1 U4627 ( .A(n3992), .B(n3986), .Z(n4262) );
  INV_X1 U4628 ( .A(n4262), .ZN(n4009) );
  OAI21_X1 U4629 ( .B1(n4033), .B2(n3988), .A(n3987), .ZN(n4013) );
  INV_X1 U4630 ( .A(n3989), .ZN(n3991) );
  OAI21_X1 U4631 ( .B1(n4013), .B2(n3991), .A(n3990), .ZN(n3993) );
  XNOR2_X1 U4632 ( .A(n3993), .B(n3992), .ZN(n3999) );
  OAI22_X1 U4633 ( .A1(n3995), .A2(n3994), .B1(n4284), .B2(n4002), .ZN(n3996)
         );
  AOI21_X1 U4634 ( .B1(n4061), .B2(n4035), .A(n3996), .ZN(n3997) );
  OAI21_X1 U4635 ( .B1(n3999), .B2(n3998), .A(n3997), .ZN(n4261) );
  INV_X1 U4636 ( .A(n4000), .ZN(n4001) );
  OAI21_X1 U4637 ( .B1(n4003), .B2(n4002), .A(n4001), .ZN(n4324) );
  AOI22_X1 U4638 ( .A1(n4507), .A2(REG2_REG_19__SCAN_IN), .B1(n4004), .B2(
        n4497), .ZN(n4005) );
  OAI21_X1 U4639 ( .B1(n4324), .B2(n4006), .A(n4005), .ZN(n4007) );
  AOI21_X1 U4640 ( .B1(n4261), .B2(n4027), .A(n4007), .ZN(n4008) );
  OAI21_X1 U4641 ( .B1(n4009), .B2(n4070), .A(n4008), .ZN(U3271) );
  OAI21_X1 U4642 ( .B1(n4011), .B2(n4014), .A(n4010), .ZN(n4012) );
  INV_X1 U4643 ( .A(n4012), .ZN(n4267) );
  XOR2_X1 U4644 ( .A(n4014), .B(n4013), .Z(n4020) );
  AOI22_X1 U4645 ( .A1(n4016), .A2(n4064), .B1(n4015), .B2(n4277), .ZN(n4017)
         );
  OAI21_X1 U4646 ( .B1(n4345), .B2(n4018), .A(n4017), .ZN(n4019) );
  AOI21_X1 U4647 ( .B1(n4020), .B2(n4057), .A(n4019), .ZN(n4266) );
  INV_X1 U4648 ( .A(n4266), .ZN(n4028) );
  XNOR2_X1 U4649 ( .A(n2048), .B(n4021), .ZN(n4022) );
  NAND2_X1 U4650 ( .A1(n4022), .A2(n4574), .ZN(n4265) );
  AOI22_X1 U4651 ( .A1(n4507), .A2(REG2_REG_18__SCAN_IN), .B1(n4023), .B2(
        n4497), .ZN(n4024) );
  OAI21_X1 U4652 ( .B1(n4265), .B2(n4025), .A(n4024), .ZN(n4026) );
  AOI21_X1 U4653 ( .B1(n4028), .B2(n4027), .A(n4026), .ZN(n4029) );
  OAI21_X1 U4654 ( .B1(n4267), .B2(n4070), .A(n4029), .ZN(U3272) );
  XOR2_X1 U4655 ( .A(n4031), .B(n4030), .Z(n4271) );
  INV_X1 U4656 ( .A(n4031), .ZN(n4032) );
  XNOR2_X1 U4657 ( .A(n4033), .B(n4032), .ZN(n4040) );
  NAND2_X1 U4658 ( .A1(n4034), .A2(n4061), .ZN(n4037) );
  NAND2_X1 U4659 ( .A1(n4035), .A2(n4064), .ZN(n4036) );
  OAI211_X1 U4660 ( .C1(n4284), .C2(n4038), .A(n4037), .B(n4036), .ZN(n4039)
         );
  AOI21_X1 U4661 ( .B1(n4040), .B2(n4057), .A(n4039), .ZN(n4270) );
  AOI22_X1 U4662 ( .A1(n4363), .A2(REG2_REG_17__SCAN_IN), .B1(n4041), .B2(
        n4497), .ZN(n4044) );
  NAND2_X1 U4663 ( .A1(n4051), .A2(n4042), .ZN(n4268) );
  NAND3_X1 U4664 ( .A1(n2048), .A2(n4501), .A3(n4268), .ZN(n4043) );
  OAI211_X1 U4665 ( .C1(n4270), .C2(n4363), .A(n4044), .B(n4043), .ZN(n4045)
         );
  INV_X1 U4666 ( .A(n4045), .ZN(n4046) );
  OAI21_X1 U4667 ( .B1(n4271), .B2(n4070), .A(n4046), .ZN(U3273) );
  OAI21_X1 U4668 ( .B1(n4049), .B2(n4048), .A(n4047), .ZN(n4276) );
  INV_X1 U4669 ( .A(n4050), .ZN(n4053) );
  INV_X1 U4670 ( .A(n4051), .ZN(n4052) );
  AOI21_X1 U4671 ( .B1(n4272), .B2(n4053), .A(n4052), .ZN(n4273) );
  AOI22_X1 U4672 ( .A1(n4507), .A2(REG2_REG_16__SCAN_IN), .B1(n4054), .B2(
        n4497), .ZN(n4055) );
  OAI21_X1 U4673 ( .B1(n4056), .B2(n4348), .A(n4055), .ZN(n4068) );
  OAI211_X1 U4674 ( .C1(n4060), .C2(n4059), .A(n4058), .B(n4057), .ZN(n4066)
         );
  AOI22_X1 U4675 ( .A1(n4064), .A2(n4063), .B1(n4062), .B2(n4061), .ZN(n4065)
         );
  AND2_X1 U4676 ( .A1(n4066), .A2(n4065), .ZN(n4275) );
  NOR2_X1 U4677 ( .A1(n4275), .A2(n4363), .ZN(n4067) );
  AOI211_X1 U4678 ( .C1(n4273), .C2(n4501), .A(n4068), .B(n4067), .ZN(n4069)
         );
  OAI21_X1 U4679 ( .B1(n4276), .B2(n4070), .A(n4069), .ZN(U3274) );
  XOR2_X1 U4680 ( .A(n4071), .B(n4077), .Z(n4364) );
  INV_X1 U4681 ( .A(n4364), .ZN(n4292) );
  INV_X1 U4682 ( .A(REG1_REG_31__SCAN_IN), .ZN(n4075) );
  NOR2_X1 U4683 ( .A1(n4073), .A2(n4072), .ZN(n4079) );
  AOI21_X1 U4684 ( .B1(n4074), .B2(n4277), .A(n4079), .ZN(n4366) );
  MUX2_X1 U4685 ( .A(n4075), .B(n4366), .S(n4588), .Z(n4076) );
  OAI21_X1 U4686 ( .B1(n4292), .B2(n4289), .A(n4076), .ZN(U3549) );
  AOI21_X1 U4687 ( .B1(n4080), .B2(n4078), .A(n4077), .ZN(n4367) );
  INV_X1 U4688 ( .A(n4367), .ZN(n4295) );
  INV_X1 U4689 ( .A(REG1_REG_30__SCAN_IN), .ZN(n4145) );
  AOI21_X1 U4690 ( .B1(n4080), .B2(n4277), .A(n4079), .ZN(n4369) );
  MUX2_X1 U4691 ( .A(n4145), .B(n4369), .S(n4588), .Z(n4081) );
  OAI21_X1 U4692 ( .B1(n4295), .B2(n4289), .A(n4081), .ZN(U3548) );
  NAND2_X1 U4693 ( .A1(n4082), .A2(n4561), .ZN(n4086) );
  MUX2_X1 U4694 ( .A(REG1_REG_29__SCAN_IN), .B(n4296), .S(n4588), .Z(U3547) );
  OAI22_X1 U4695 ( .A1(n4088), .A2(n4559), .B1(n4087), .B2(n4284), .ZN(n4089)
         );
  NOR2_X1 U4696 ( .A1(n4588), .A2(REG1_REG_27__SCAN_IN), .ZN(n4092) );
  AOI21_X1 U4697 ( .B1(n4298), .B2(n4588), .A(n4092), .ZN(n4226) );
  AOI22_X1 U4698 ( .A1(n4094), .A2(keyinput34), .B1(keyinput52), .B2(n4202), 
        .ZN(n4093) );
  OAI221_X1 U4699 ( .B1(n4094), .B2(keyinput34), .C1(n4202), .C2(keyinput52), 
        .A(n4093), .ZN(n4161) );
  AOI22_X1 U4700 ( .A1(n4196), .A2(keyinput58), .B1(n4096), .B2(keyinput63), 
        .ZN(n4095) );
  OAI221_X1 U4701 ( .B1(n4196), .B2(keyinput58), .C1(n4096), .C2(keyinput63), 
        .A(n4095), .ZN(n4160) );
  OAI22_X1 U4702 ( .A1(n4099), .A2(keyinput12), .B1(n4098), .B2(keyinput19), 
        .ZN(n4097) );
  AOI221_X1 U4703 ( .B1(n4099), .B2(keyinput12), .C1(keyinput19), .C2(n4098), 
        .A(n4097), .ZN(n4114) );
  XOR2_X1 U4704 ( .A(keyinput11), .B(DATAO_REG_7__SCAN_IN), .Z(n4110) );
  AOI22_X1 U4705 ( .A1(n3842), .A2(keyinput53), .B1(keyinput7), .B2(n4101), 
        .ZN(n4100) );
  OAI221_X1 U4706 ( .B1(n3842), .B2(keyinput53), .C1(n4101), .C2(keyinput7), 
        .A(n4100), .ZN(n4109) );
  INV_X1 U4707 ( .A(ADDR_REG_18__SCAN_IN), .ZN(n4489) );
  AOI22_X1 U4708 ( .A1(n2513), .A2(keyinput24), .B1(keyinput37), .B2(n4489), 
        .ZN(n4102) );
  OAI221_X1 U4709 ( .B1(n2513), .B2(keyinput24), .C1(n4489), .C2(keyinput37), 
        .A(n4102), .ZN(n4108) );
  XNOR2_X1 U4710 ( .A(keyinput33), .B(ADDR_REG_3__SCAN_IN), .ZN(n4105) );
  XOR2_X1 U4711 ( .A(keyinput43), .B(DATAO_REG_0__SCAN_IN), .Z(n4103) );
  AOI21_X1 U4712 ( .B1(keyinput54), .B2(n4106), .A(n4103), .ZN(n4104) );
  OAI211_X1 U4713 ( .C1(keyinput54), .C2(n4106), .A(n4105), .B(n4104), .ZN(
        n4107) );
  NOR4_X1 U4714 ( .A1(n4110), .A2(n4109), .A3(n4108), .A4(n4107), .ZN(n4113)
         );
  XNOR2_X1 U4715 ( .A(keyinput56), .B(DATAO_REG_15__SCAN_IN), .ZN(n4112) );
  XNOR2_X1 U4716 ( .A(keyinput20), .B(DATAO_REG_14__SCAN_IN), .ZN(n4111) );
  NAND4_X1 U4717 ( .A1(n4114), .A2(n4113), .A3(n4112), .A4(n4111), .ZN(n4159)
         );
  INV_X1 U4718 ( .A(D_REG_29__SCAN_IN), .ZN(n4509) );
  INV_X1 U4719 ( .A(D_REG_28__SCAN_IN), .ZN(n4510) );
  AOI22_X1 U4720 ( .A1(n4509), .A2(keyinput25), .B1(n4510), .B2(keyinput57), 
        .ZN(n4115) );
  OAI221_X1 U4721 ( .B1(n4509), .B2(keyinput25), .C1(n4510), .C2(keyinput57), 
        .A(n4115), .ZN(n4118) );
  XNOR2_X1 U4722 ( .A(n4201), .B(keyinput14), .ZN(n4117) );
  INV_X1 U4723 ( .A(D_REG_3__SCAN_IN), .ZN(n4515) );
  XNOR2_X1 U4724 ( .A(n4515), .B(keyinput62), .ZN(n4116) );
  OR3_X1 U4725 ( .A1(n4118), .A2(n4117), .A3(n4116), .ZN(n4123) );
  INV_X1 U4726 ( .A(D_REG_10__SCAN_IN), .ZN(n4512) );
  INV_X1 U4727 ( .A(D_REG_19__SCAN_IN), .ZN(n4511) );
  AOI22_X1 U4728 ( .A1(n4512), .A2(keyinput36), .B1(n4511), .B2(keyinput47), 
        .ZN(n4119) );
  OAI221_X1 U4729 ( .B1(n4512), .B2(keyinput36), .C1(n4511), .C2(keyinput47), 
        .A(n4119), .ZN(n4122) );
  INV_X1 U4730 ( .A(D_REG_5__SCAN_IN), .ZN(n4514) );
  INV_X1 U4731 ( .A(D_REG_6__SCAN_IN), .ZN(n4513) );
  AOI22_X1 U4732 ( .A1(n4514), .A2(keyinput10), .B1(n4513), .B2(keyinput41), 
        .ZN(n4120) );
  OAI221_X1 U4733 ( .B1(n4514), .B2(keyinput10), .C1(n4513), .C2(keyinput41), 
        .A(n4120), .ZN(n4121) );
  NOR3_X1 U4734 ( .A1(n4123), .A2(n4122), .A3(n4121), .ZN(n4157) );
  INV_X1 U4735 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4125) );
  INV_X1 U4736 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4322) );
  AOI22_X1 U4737 ( .A1(n4125), .A2(keyinput39), .B1(keyinput0), .B2(n4322), 
        .ZN(n4124) );
  OAI221_X1 U4738 ( .B1(n4125), .B2(keyinput39), .C1(n4322), .C2(keyinput0), 
        .A(n4124), .ZN(n4129) );
  INV_X1 U4739 ( .A(REG0_REG_15__SCAN_IN), .ZN(n4203) );
  INV_X1 U4740 ( .A(REG0_REG_14__SCAN_IN), .ZN(n4330) );
  AOI22_X1 U4741 ( .A1(n4203), .A2(keyinput61), .B1(n4330), .B2(keyinput60), 
        .ZN(n4126) );
  OAI221_X1 U4742 ( .B1(n4203), .B2(keyinput61), .C1(n4330), .C2(keyinput60), 
        .A(n4126), .ZN(n4128) );
  INV_X1 U4743 ( .A(REG0_REG_2__SCAN_IN), .ZN(n4213) );
  XNOR2_X1 U4744 ( .A(n4213), .B(keyinput18), .ZN(n4127) );
  OR3_X1 U4745 ( .A1(n4129), .A2(n4128), .A3(n4127), .ZN(n4134) );
  INV_X1 U4746 ( .A(REG0_REG_9__SCAN_IN), .ZN(n4576) );
  AOI22_X1 U4747 ( .A1(n4131), .A2(keyinput50), .B1(keyinput16), .B2(n4576), 
        .ZN(n4130) );
  OAI221_X1 U4748 ( .B1(n4131), .B2(keyinput50), .C1(n4576), .C2(keyinput16), 
        .A(n4130), .ZN(n4133) );
  INV_X1 U4749 ( .A(D_REG_30__SCAN_IN), .ZN(n4508) );
  XNOR2_X1 U4750 ( .A(n4508), .B(keyinput31), .ZN(n4132) );
  NOR3_X1 U4751 ( .A1(n4134), .A2(n4133), .A3(n4132), .ZN(n4156) );
  INV_X1 U4752 ( .A(REG0_REG_22__SCAN_IN), .ZN(n4136) );
  INV_X1 U4753 ( .A(REG0_REG_31__SCAN_IN), .ZN(n4290) );
  AOI22_X1 U4754 ( .A1(n4136), .A2(keyinput27), .B1(keyinput26), .B2(n4290), 
        .ZN(n4135) );
  OAI221_X1 U4755 ( .B1(n4136), .B2(keyinput27), .C1(n4290), .C2(keyinput26), 
        .A(n4135), .ZN(n4143) );
  INV_X1 U4756 ( .A(REG1_REG_7__SCAN_IN), .ZN(n4584) );
  AOI22_X1 U4757 ( .A1(n4584), .A2(keyinput30), .B1(n4582), .B2(keyinput28), 
        .ZN(n4137) );
  OAI221_X1 U4758 ( .B1(n4584), .B2(keyinput30), .C1(n4582), .C2(keyinput28), 
        .A(n4137), .ZN(n4142) );
  AOI22_X1 U4759 ( .A1(n2808), .A2(keyinput17), .B1(keyinput22), .B2(n4394), 
        .ZN(n4138) );
  OAI221_X1 U4760 ( .B1(n2808), .B2(keyinput17), .C1(n4394), .C2(keyinput22), 
        .A(n4138), .ZN(n4141) );
  INV_X1 U4761 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4263) );
  AOI22_X1 U4762 ( .A1(n4263), .A2(keyinput46), .B1(keyinput15), .B2(n4197), 
        .ZN(n4139) );
  OAI221_X1 U4763 ( .B1(n4263), .B2(keyinput46), .C1(n4197), .C2(keyinput15), 
        .A(n4139), .ZN(n4140) );
  NOR4_X1 U4764 ( .A1(n4143), .A2(n4142), .A3(n4141), .A4(n4140), .ZN(n4155)
         );
  INV_X1 U4765 ( .A(REG1_REG_28__SCAN_IN), .ZN(n4190) );
  AOI22_X1 U4766 ( .A1(n4145), .A2(keyinput23), .B1(n4190), .B2(keyinput48), 
        .ZN(n4144) );
  OAI221_X1 U4767 ( .B1(n4145), .B2(keyinput23), .C1(n4190), .C2(keyinput48), 
        .A(n4144), .ZN(n4153) );
  AOI22_X1 U4768 ( .A1(n4211), .A2(keyinput3), .B1(keyinput9), .B2(n2686), 
        .ZN(n4146) );
  OAI221_X1 U4769 ( .B1(n4211), .B2(keyinput3), .C1(n2686), .C2(keyinput9), 
        .A(n4146), .ZN(n4152) );
  AOI22_X1 U4770 ( .A1(n2390), .A2(keyinput6), .B1(keyinput2), .B2(n2406), 
        .ZN(n4147) );
  OAI221_X1 U4771 ( .B1(n2390), .B2(keyinput6), .C1(n2406), .C2(keyinput2), 
        .A(n4147), .ZN(n4151) );
  INV_X1 U4772 ( .A(REG2_REG_25__SCAN_IN), .ZN(n4149) );
  AOI22_X1 U4773 ( .A1(n4149), .A2(keyinput13), .B1(keyinput32), .B2(n2452), 
        .ZN(n4148) );
  OAI221_X1 U4774 ( .B1(n4149), .B2(keyinput13), .C1(n2452), .C2(keyinput32), 
        .A(n4148), .ZN(n4150) );
  NOR4_X1 U4775 ( .A1(n4153), .A2(n4152), .A3(n4151), .A4(n4150), .ZN(n4154)
         );
  NAND4_X1 U4776 ( .A1(n4157), .A2(n4156), .A3(n4155), .A4(n4154), .ZN(n4158)
         );
  NOR4_X1 U4777 ( .A1(n4161), .A2(n4160), .A3(n4159), .A4(n4158), .ZN(n4189)
         );
  XOR2_X1 U4778 ( .A(REG3_REG_4__SCAN_IN), .B(keyinput35), .Z(n4166) );
  XOR2_X1 U4779 ( .A(DATAI_4_), .B(keyinput45), .Z(n4165) );
  XOR2_X1 U4780 ( .A(IR_REG_0__SCAN_IN), .B(keyinput8), .Z(n4164) );
  XNOR2_X1 U4781 ( .A(n4162), .B(keyinput42), .ZN(n4163) );
  NOR4_X1 U4782 ( .A1(n4166), .A2(n4165), .A3(n4164), .A4(n4163), .ZN(n4179)
         );
  XOR2_X1 U4783 ( .A(n2422), .B(keyinput38), .Z(n4178) );
  INV_X1 U4784 ( .A(IR_REG_18__SCAN_IN), .ZN(n4167) );
  XOR2_X1 U4785 ( .A(n4167), .B(keyinput51), .Z(n4177) );
  INV_X1 U4786 ( .A(DATAI_15_), .ZN(n4525) );
  INV_X1 U4787 ( .A(DATAI_18_), .ZN(n4520) );
  AOI22_X1 U4788 ( .A1(n4525), .A2(keyinput4), .B1(n4520), .B2(keyinput55), 
        .ZN(n4168) );
  OAI221_X1 U4789 ( .B1(n4525), .B2(keyinput4), .C1(n4520), .C2(keyinput55), 
        .A(n4168), .ZN(n4175) );
  XOR2_X1 U4790 ( .A(n4214), .B(keyinput21), .Z(n4173) );
  XOR2_X1 U4791 ( .A(n4169), .B(keyinput44), .Z(n4172) );
  XNOR2_X1 U4792 ( .A(IR_REG_17__SCAN_IN), .B(keyinput29), .ZN(n4171) );
  XNOR2_X1 U4793 ( .A(IR_REG_20__SCAN_IN), .B(keyinput5), .ZN(n4170) );
  NAND4_X1 U4794 ( .A1(n4173), .A2(n4172), .A3(n4171), .A4(n4170), .ZN(n4174)
         );
  NOR2_X1 U4795 ( .A1(n4175), .A2(n4174), .ZN(n4176) );
  NAND4_X1 U4796 ( .A1(n4179), .A2(n4178), .A3(n4177), .A4(n4176), .ZN(n4187)
         );
  AOI22_X1 U4797 ( .A1(n4182), .A2(keyinput1), .B1(n4181), .B2(keyinput59), 
        .ZN(n4180) );
  OAI221_X1 U4798 ( .B1(n4182), .B2(keyinput1), .C1(n4181), .C2(keyinput59), 
        .A(n4180), .ZN(n4186) );
  INV_X1 U4799 ( .A(DATAI_28_), .ZN(n4340) );
  AOI22_X1 U4800 ( .A1(n4184), .A2(keyinput40), .B1(n4340), .B2(keyinput49), 
        .ZN(n4183) );
  OAI221_X1 U4801 ( .B1(n4184), .B2(keyinput40), .C1(n4340), .C2(keyinput49), 
        .A(n4183), .ZN(n4185) );
  NOR3_X1 U4802 ( .A1(n4187), .A2(n4186), .A3(n4185), .ZN(n4188) );
  NAND2_X1 U4803 ( .A1(n4189), .A2(n4188), .ZN(n4224) );
  NAND4_X1 U4804 ( .A1(REG2_REG_29__SCAN_IN), .A2(DATAO_REG_14__SCAN_IN), .A3(
        ADDR_REG_7__SCAN_IN), .A4(ADDR_REG_18__SCAN_IN), .ZN(n4195) );
  NAND3_X1 U4805 ( .A1(DATAO_REG_10__SCAN_IN), .A2(ADDR_REG_3__SCAN_IN), .A3(
        DATAO_REG_0__SCAN_IN), .ZN(n4194) );
  NOR3_X1 U4806 ( .A1(DATAI_28_), .A2(REG1_REG_30__SCAN_IN), .A3(n4190), .ZN(
        n4192) );
  NOR3_X1 U4807 ( .A1(DATAO_REG_20__SCAN_IN), .A2(DATAO_REG_28__SCAN_IN), .A3(
        n4290), .ZN(n4191) );
  NAND4_X1 U4808 ( .A1(REG0_REG_22__SCAN_IN), .A2(DATAO_REG_15__SCAN_IN), .A3(
        n4192), .A4(n4191), .ZN(n4193) );
  NOR4_X1 U4809 ( .A1(DATAO_REG_7__SCAN_IN), .A2(n4195), .A3(n4194), .A4(n4193), .ZN(n4222) );
  NOR4_X1 U4810 ( .A1(REG3_REG_26__SCAN_IN), .A2(REG3_REG_25__SCAN_IN), .A3(
        REG2_REG_27__SCAN_IN), .A4(n4196), .ZN(n4200) );
  NOR3_X1 U4811 ( .A1(DATAI_27_), .A2(REG2_REG_25__SCAN_IN), .A3(
        REG1_REG_19__SCAN_IN), .ZN(n4199) );
  NOR4_X1 U4812 ( .A1(REG0_REG_19__SCAN_IN), .A2(DATAI_18_), .A3(n2452), .A4(
        n4197), .ZN(n4198) );
  NAND4_X1 U4813 ( .A1(REG0_REG_21__SCAN_IN), .A2(n4200), .A3(n4199), .A4(
        n4198), .ZN(n4219) );
  NAND4_X1 U4814 ( .A1(D_REG_10__SCAN_IN), .A2(D_REG_29__SCAN_IN), .A3(
        D_REG_30__SCAN_IN), .A4(D_REG_5__SCAN_IN), .ZN(n4218) );
  NAND4_X1 U4815 ( .A1(n2242), .A2(n4201), .A3(IR_REG_2__SCAN_IN), .A4(
        IR_REG_5__SCAN_IN), .ZN(n4212) );
  NAND4_X1 U4816 ( .A1(REG3_REG_17__SCAN_IN), .A2(REG3_REG_10__SCAN_IN), .A3(
        REG3_REG_4__SCAN_IN), .A4(n4202), .ZN(n4205) );
  NAND4_X1 U4817 ( .A1(REG0_REG_14__SCAN_IN), .A2(REG2_REG_15__SCAN_IN), .A3(
        DATAI_15_), .A4(n4203), .ZN(n4204) );
  NOR2_X1 U4818 ( .A1(n4205), .A2(n4204), .ZN(n4209) );
  NOR4_X1 U4819 ( .A1(REG0_REG_11__SCAN_IN), .A2(REG1_REG_9__SCAN_IN), .A3(
        REG0_REG_9__SCAN_IN), .A4(n4394), .ZN(n4208) );
  NOR3_X1 U4820 ( .A1(IR_REG_15__SCAN_IN), .A2(IR_REG_20__SCAN_IN), .A3(n2132), 
        .ZN(n4207) );
  AND3_X1 U4821 ( .A1(REG2_REG_7__SCAN_IN), .A2(REG2_REG_12__SCAN_IN), .A3(
        n4584), .ZN(n4206) );
  NAND4_X1 U4822 ( .A1(n4209), .A2(n4208), .A3(n4207), .A4(n4206), .ZN(n4210)
         );
  OR4_X1 U4823 ( .A1(n4212), .A2(n4211), .A3(IR_REG_18__SCAN_IN), .A4(n4210), 
        .ZN(n4217) );
  INV_X1 U4824 ( .A(DATAI_4_), .ZN(n4215) );
  NAND4_X1 U4825 ( .A1(n4215), .A2(n4214), .A3(n4213), .A4(REG1_REG_5__SCAN_IN), .ZN(n4216) );
  NOR4_X1 U4826 ( .A1(n4219), .A2(n4218), .A3(n4217), .A4(n4216), .ZN(n4220)
         );
  NAND3_X1 U4827 ( .A1(n4222), .A2(n4221), .A3(n4220), .ZN(n4223) );
  XNOR2_X1 U4828 ( .A(n4224), .B(n4223), .ZN(n4225) );
  XNOR2_X1 U4829 ( .A(n4226), .B(n4225), .ZN(U3545) );
  INV_X1 U4830 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4229) );
  AOI21_X1 U4831 ( .B1(n4228), .B2(n4561), .A(n4227), .ZN(n4299) );
  MUX2_X1 U4832 ( .A(n4229), .B(n4299), .S(n4588), .Z(n4230) );
  OAI21_X1 U4833 ( .B1(n4289), .B2(n4302), .A(n4230), .ZN(U3544) );
  INV_X1 U4834 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4233) );
  AOI21_X1 U4835 ( .B1(n4232), .B2(n4561), .A(n4231), .ZN(n4303) );
  MUX2_X1 U4836 ( .A(n4233), .B(n4303), .S(n4588), .Z(n4234) );
  OAI21_X1 U4837 ( .B1(n4289), .B2(n4306), .A(n4234), .ZN(U3543) );
  INV_X1 U4838 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4239) );
  OAI21_X1 U4839 ( .B1(n4236), .B2(n4284), .A(n4235), .ZN(n4237) );
  AOI21_X1 U4840 ( .B1(n4238), .B2(n4561), .A(n4237), .ZN(n4307) );
  MUX2_X1 U4841 ( .A(n4239), .B(n4307), .S(n4588), .Z(n4240) );
  OAI21_X1 U4842 ( .B1(n4289), .B2(n4310), .A(n4240), .ZN(U3542) );
  INV_X1 U4843 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4243) );
  AOI21_X1 U4844 ( .B1(n4242), .B2(n4561), .A(n4241), .ZN(n4311) );
  MUX2_X1 U4845 ( .A(n4243), .B(n4311), .S(n4588), .Z(n4244) );
  OAI21_X1 U4846 ( .B1(n4289), .B2(n4314), .A(n4244), .ZN(U3541) );
  NAND3_X1 U4847 ( .A1(n4246), .A2(n4574), .A3(n4245), .ZN(n4247) );
  OAI211_X1 U4848 ( .C1(n4249), .C2(n4569), .A(n4248), .B(n4247), .ZN(n4315)
         );
  MUX2_X1 U4849 ( .A(REG1_REG_22__SCAN_IN), .B(n4315), .S(n4588), .Z(U3540) );
  AOI22_X1 U4850 ( .A1(n4251), .A2(n4574), .B1(n4250), .B2(n4277), .ZN(n4252)
         );
  OAI211_X1 U4851 ( .C1(n4254), .C2(n4569), .A(n4253), .B(n4252), .ZN(n4316)
         );
  MUX2_X1 U4852 ( .A(REG1_REG_21__SCAN_IN), .B(n4316), .S(n4588), .Z(U3539) );
  INV_X1 U4853 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4259) );
  OAI21_X1 U4854 ( .B1(n4256), .B2(n4284), .A(n4255), .ZN(n4257) );
  AOI21_X1 U4855 ( .B1(n4258), .B2(n4561), .A(n4257), .ZN(n4317) );
  MUX2_X1 U4856 ( .A(n4259), .B(n4317), .S(n4588), .Z(n4260) );
  OAI21_X1 U4857 ( .B1(n4289), .B2(n4320), .A(n4260), .ZN(U3538) );
  AOI21_X1 U4858 ( .B1(n4262), .B2(n4561), .A(n4261), .ZN(n4321) );
  MUX2_X1 U4859 ( .A(n4263), .B(n4321), .S(n4588), .Z(n4264) );
  OAI21_X1 U4860 ( .B1(n4289), .B2(n4324), .A(n4264), .ZN(U3537) );
  OAI211_X1 U4861 ( .C1(n4267), .C2(n4569), .A(n4266), .B(n4265), .ZN(n4325)
         );
  MUX2_X1 U4862 ( .A(REG1_REG_18__SCAN_IN), .B(n4325), .S(n4588), .Z(U3536) );
  NAND3_X1 U4863 ( .A1(n2048), .A2(n4574), .A3(n4268), .ZN(n4269) );
  OAI211_X1 U4864 ( .C1(n4271), .C2(n4569), .A(n4270), .B(n4269), .ZN(n4326)
         );
  MUX2_X1 U4865 ( .A(REG1_REG_17__SCAN_IN), .B(n4326), .S(n4588), .Z(U3535) );
  AOI22_X1 U4866 ( .A1(n4273), .A2(n4574), .B1(n4272), .B2(n4277), .ZN(n4274)
         );
  OAI211_X1 U4867 ( .C1(n4276), .C2(n4569), .A(n4275), .B(n4274), .ZN(n4327)
         );
  MUX2_X1 U4868 ( .A(REG1_REG_16__SCAN_IN), .B(n4327), .S(n4588), .Z(U3534) );
  AOI22_X1 U4869 ( .A1(n4279), .A2(n4574), .B1(n4278), .B2(n4277), .ZN(n4280)
         );
  OAI211_X1 U4870 ( .C1(n4282), .C2(n4569), .A(n4281), .B(n4280), .ZN(n4328)
         );
  MUX2_X1 U4871 ( .A(REG1_REG_15__SCAN_IN), .B(n4328), .S(n4588), .Z(U3533) );
  OAI21_X1 U4872 ( .B1(n4285), .B2(n4284), .A(n4283), .ZN(n4286) );
  AOI21_X1 U4873 ( .B1(n4287), .B2(n4561), .A(n4286), .ZN(n4329) );
  MUX2_X1 U4874 ( .A(n4432), .B(n4329), .S(n4588), .Z(n4288) );
  OAI21_X1 U4875 ( .B1(n4289), .B2(n4333), .A(n4288), .ZN(U3532) );
  MUX2_X1 U4876 ( .A(n4290), .B(n4366), .S(n4577), .Z(n4291) );
  OAI21_X1 U4877 ( .B1(n4292), .B2(n4332), .A(n4291), .ZN(U3517) );
  INV_X1 U4878 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4293) );
  MUX2_X1 U4879 ( .A(n4293), .B(n4369), .S(n4577), .Z(n4294) );
  OAI21_X1 U4880 ( .B1(n4295), .B2(n4332), .A(n4294), .ZN(U3516) );
  MUX2_X1 U4881 ( .A(REG0_REG_29__SCAN_IN), .B(n4296), .S(n4577), .Z(U3515) );
  NAND2_X1 U4882 ( .A1(n4575), .A2(REG0_REG_27__SCAN_IN), .ZN(n4297) );
  OAI21_X1 U4883 ( .B1(n4298), .B2(n4575), .A(n4297), .ZN(U3513) );
  INV_X1 U4884 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4300) );
  MUX2_X1 U4885 ( .A(n4300), .B(n4299), .S(n4577), .Z(n4301) );
  OAI21_X1 U4886 ( .B1(n4302), .B2(n4332), .A(n4301), .ZN(U3512) );
  INV_X1 U4887 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4304) );
  MUX2_X1 U4888 ( .A(n4304), .B(n4303), .S(n4577), .Z(n4305) );
  OAI21_X1 U4889 ( .B1(n4306), .B2(n4332), .A(n4305), .ZN(U3511) );
  INV_X1 U4890 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4308) );
  MUX2_X1 U4891 ( .A(n4308), .B(n4307), .S(n4577), .Z(n4309) );
  OAI21_X1 U4892 ( .B1(n4310), .B2(n4332), .A(n4309), .ZN(U3510) );
  INV_X1 U4893 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4312) );
  MUX2_X1 U4894 ( .A(n4312), .B(n4311), .S(n4577), .Z(n4313) );
  OAI21_X1 U4895 ( .B1(n4314), .B2(n4332), .A(n4313), .ZN(U3509) );
  MUX2_X1 U4896 ( .A(REG0_REG_22__SCAN_IN), .B(n4315), .S(n4577), .Z(U3508) );
  MUX2_X1 U4897 ( .A(REG0_REG_21__SCAN_IN), .B(n4316), .S(n4577), .Z(U3507) );
  INV_X1 U4898 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4318) );
  MUX2_X1 U4899 ( .A(n4318), .B(n4317), .S(n4577), .Z(n4319) );
  OAI21_X1 U4900 ( .B1(n4320), .B2(n4332), .A(n4319), .ZN(U3506) );
  MUX2_X1 U4901 ( .A(n4322), .B(n4321), .S(n4577), .Z(n4323) );
  OAI21_X1 U4902 ( .B1(n4324), .B2(n4332), .A(n4323), .ZN(U3505) );
  MUX2_X1 U4903 ( .A(REG0_REG_18__SCAN_IN), .B(n4325), .S(n4577), .Z(U3503) );
  MUX2_X1 U4904 ( .A(REG0_REG_17__SCAN_IN), .B(n4326), .S(n4577), .Z(U3501) );
  MUX2_X1 U4905 ( .A(REG0_REG_16__SCAN_IN), .B(n4327), .S(n4577), .Z(U3499) );
  MUX2_X1 U4906 ( .A(REG0_REG_15__SCAN_IN), .B(n4328), .S(n4577), .Z(U3497) );
  MUX2_X1 U4907 ( .A(n4330), .B(n4329), .S(n4577), .Z(n4331) );
  OAI21_X1 U4908 ( .B1(n4333), .B2(n4332), .A(n4331), .ZN(U3495) );
  MUX2_X1 U4909 ( .A(n4334), .B(DATAI_19_), .S(U3149), .Z(U3333) );
  MUX2_X1 U4910 ( .A(n4335), .B(DATAI_9_), .S(U3149), .Z(U3343) );
  MUX2_X1 U4911 ( .A(n4336), .B(DATAI_7_), .S(U3149), .Z(U3345) );
  MUX2_X1 U4912 ( .A(DATAI_4_), .B(n4377), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U4913 ( .A(n4337), .B(DATAI_3_), .S(U3149), .Z(U3349) );
  MUX2_X1 U4914 ( .A(n4338), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  MUX2_X1 U4915 ( .A(n4339), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  AOI22_X1 U4916 ( .A1(STATE_REG_SCAN_IN), .A2(n4341), .B1(n4340), .B2(U3149), 
        .ZN(U3324) );
  OAI22_X1 U4917 ( .A1(n4345), .A2(n4344), .B1(n4343), .B2(n4342), .ZN(n4351)
         );
  INV_X1 U4918 ( .A(REG3_REG_16__SCAN_IN), .ZN(n4346) );
  NOR2_X1 U4919 ( .A1(STATE_REG_SCAN_IN), .A2(n4346), .ZN(n4451) );
  INV_X1 U4920 ( .A(n4451), .ZN(n4347) );
  OAI21_X1 U4921 ( .B1(n4349), .B2(n4348), .A(n4347), .ZN(n4350) );
  NOR2_X1 U4922 ( .A1(n4351), .A2(n4350), .ZN(n4360) );
  AOI21_X1 U4923 ( .B1(n4354), .B2(n4353), .A(n4352), .ZN(n4355) );
  XOR2_X1 U4924 ( .A(n4356), .B(n4355), .Z(n4358) );
  NAND2_X1 U4925 ( .A1(n4358), .A2(n4357), .ZN(n4359) );
  OAI211_X1 U4926 ( .C1(n4362), .C2(n4361), .A(n4360), .B(n4359), .ZN(U3223)
         );
  AOI22_X1 U4927 ( .A1(n4364), .A2(n4501), .B1(n4363), .B2(
        REG2_REG_31__SCAN_IN), .ZN(n4365) );
  OAI21_X1 U4928 ( .B1(n4507), .B2(n4366), .A(n4365), .ZN(U3260) );
  AOI22_X1 U4929 ( .A1(n4367), .A2(n4501), .B1(REG2_REG_30__SCAN_IN), .B2(
        n4363), .ZN(n4368) );
  OAI21_X1 U4930 ( .B1(n4507), .B2(n4369), .A(n4368), .ZN(U3261) );
  INV_X1 U4931 ( .A(n4370), .ZN(n4371) );
  AOI21_X1 U4932 ( .B1(n4462), .B2(ADDR_REG_4__SCAN_IN), .A(n4371), .ZN(n4381)
         );
  XNOR2_X1 U4933 ( .A(n4372), .B(REG2_REG_4__SCAN_IN), .ZN(n4373) );
  NAND2_X1 U4934 ( .A1(n4472), .A2(n4373), .ZN(n4380) );
  INV_X1 U4935 ( .A(REG1_REG_4__SCAN_IN), .ZN(n4374) );
  XNOR2_X1 U4936 ( .A(n4375), .B(n4374), .ZN(n4376) );
  NAND2_X1 U4937 ( .A1(n4470), .A2(n4376), .ZN(n4379) );
  NAND2_X1 U4938 ( .A1(n4484), .A2(n4377), .ZN(n4378) );
  AND4_X1 U4939 ( .A1(n4381), .A2(n4380), .A3(n4379), .A4(n4378), .ZN(n4383)
         );
  NAND2_X1 U4940 ( .A1(n4383), .A2(n4382), .ZN(U3244) );
  OAI211_X1 U4941 ( .C1(REG1_REG_6__SCAN_IN), .C2(n4385), .A(n4470), .B(n4384), 
        .ZN(n4389) );
  OAI211_X1 U4942 ( .C1(REG2_REG_6__SCAN_IN), .C2(n4387), .A(n4472), .B(n4386), 
        .ZN(n4388) );
  OAI211_X1 U4943 ( .C1(n4475), .C2(n4536), .A(n4389), .B(n4388), .ZN(n4390)
         );
  AOI211_X1 U4944 ( .C1(n4462), .C2(ADDR_REG_6__SCAN_IN), .A(n4391), .B(n4390), 
        .ZN(n4392) );
  INV_X1 U4945 ( .A(n4392), .ZN(U3246) );
  AOI211_X1 U4946 ( .C1(n4394), .C2(n4393), .A(n2050), .B(n4476), .ZN(n4397)
         );
  INV_X1 U4947 ( .A(n4395), .ZN(n4396) );
  AOI211_X1 U4948 ( .C1(n4462), .C2(ADDR_REG_8__SCAN_IN), .A(n4397), .B(n4396), 
        .ZN(n4401) );
  OAI211_X1 U4949 ( .C1(REG2_REG_8__SCAN_IN), .C2(n4399), .A(n4472), .B(n4398), 
        .ZN(n4400) );
  OAI211_X1 U4950 ( .C1(n4475), .C2(n4534), .A(n4401), .B(n4400), .ZN(U3248)
         );
  AOI211_X1 U4951 ( .C1(n4404), .C2(n4403), .A(n4402), .B(n4476), .ZN(n4406)
         );
  AOI211_X1 U4952 ( .C1(n4462), .C2(ADDR_REG_10__SCAN_IN), .A(n4406), .B(n4405), .ZN(n4410) );
  OAI211_X1 U4953 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4408), .A(n4472), .B(n4407), .ZN(n4409) );
  OAI211_X1 U4954 ( .C1(n4475), .C2(n4533), .A(n4410), .B(n4409), .ZN(U3250)
         );
  AOI211_X1 U4955 ( .C1(n2049), .C2(n4412), .A(n4411), .B(n4476), .ZN(n4414)
         );
  AOI211_X1 U4956 ( .C1(n4462), .C2(ADDR_REG_11__SCAN_IN), .A(n4414), .B(n4413), .ZN(n4419) );
  OAI211_X1 U4957 ( .C1(n4417), .C2(n4416), .A(n4472), .B(n4415), .ZN(n4418)
         );
  OAI211_X1 U4958 ( .C1(n4475), .C2(n4531), .A(n4419), .B(n4418), .ZN(U3251)
         );
  AOI211_X1 U4959 ( .C1(n4422), .C2(n4421), .A(n4420), .B(n4476), .ZN(n4425)
         );
  INV_X1 U4960 ( .A(n4423), .ZN(n4424) );
  AOI211_X1 U4961 ( .C1(n4462), .C2(ADDR_REG_12__SCAN_IN), .A(n4425), .B(n4424), .ZN(n4429) );
  OAI211_X1 U4962 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4427), .A(n4472), .B(n4426), .ZN(n4428) );
  OAI211_X1 U4963 ( .C1(n4475), .C2(n4529), .A(n4429), .B(n4428), .ZN(U3252)
         );
  NAND2_X1 U4964 ( .A1(ADDR_REG_14__SCAN_IN), .A2(n4462), .ZN(n4440) );
  AOI211_X1 U4965 ( .C1(n4432), .C2(n4431), .A(n4430), .B(n4476), .ZN(n4436)
         );
  AOI211_X1 U4966 ( .C1(n2261), .C2(n4434), .A(n4433), .B(n4479), .ZN(n4435)
         );
  AOI211_X1 U4967 ( .C1(n4484), .C2(n4437), .A(n4436), .B(n4435), .ZN(n4439)
         );
  NAND3_X1 U4968 ( .A1(n4440), .A2(n4439), .A3(n4438), .ZN(U3254) );
  AOI211_X1 U4969 ( .C1(n4443), .C2(n4442), .A(n4441), .B(n4479), .ZN(n4444)
         );
  AOI211_X1 U4970 ( .C1(n4462), .C2(ADDR_REG_15__SCAN_IN), .A(n4445), .B(n4444), .ZN(n4450) );
  AOI21_X1 U4971 ( .B1(n4447), .B2(n2046), .A(n4446), .ZN(n4448) );
  NAND2_X1 U4972 ( .A1(n4470), .A2(n4448), .ZN(n4449) );
  OAI211_X1 U4973 ( .C1(n4475), .C2(n4526), .A(n4450), .B(n4449), .ZN(U3255)
         );
  AOI21_X1 U4974 ( .B1(n4462), .B2(ADDR_REG_16__SCAN_IN), .A(n4451), .ZN(n4460) );
  OAI21_X1 U4975 ( .B1(n4453), .B2(n2417), .A(n4452), .ZN(n4458) );
  OAI21_X1 U4976 ( .B1(n4456), .B2(n4455), .A(n4454), .ZN(n4457) );
  AOI22_X1 U4977 ( .A1(n4472), .A2(n4458), .B1(n4470), .B2(n4457), .ZN(n4459)
         );
  OAI211_X1 U4978 ( .C1(n4524), .C2(n4475), .A(n4460), .B(n4459), .ZN(U3256)
         );
  AOI21_X1 U4979 ( .B1(n4462), .B2(ADDR_REG_17__SCAN_IN), .A(n4461), .ZN(n4474) );
  OAI21_X1 U4980 ( .B1(n4465), .B2(n4464), .A(n4463), .ZN(n4471) );
  OAI21_X1 U4981 ( .B1(n4468), .B2(n4467), .A(n4466), .ZN(n4469) );
  AOI22_X1 U4982 ( .A1(n4472), .A2(n4471), .B1(n4470), .B2(n4469), .ZN(n4473)
         );
  OAI211_X1 U4983 ( .C1(n4522), .C2(n4475), .A(n4474), .B(n4473), .ZN(U3257)
         );
  AOI21_X1 U4984 ( .B1(n4478), .B2(n4477), .A(n4476), .ZN(n4485) );
  INV_X1 U4985 ( .A(n4486), .ZN(n4487) );
  AOI22_X1 U4986 ( .A1(n4490), .A2(n4497), .B1(REG2_REG_10__SCAN_IN), .B2(
        n4507), .ZN(n4495) );
  INV_X1 U4987 ( .A(n4491), .ZN(n4492) );
  AOI22_X1 U4988 ( .A1(n4493), .A2(n4502), .B1(n4501), .B2(n4492), .ZN(n4494)
         );
  OAI211_X1 U4989 ( .C1(n4507), .C2(n4496), .A(n4495), .B(n4494), .ZN(U3280)
         );
  AOI22_X1 U4990 ( .A1(n4498), .A2(n4497), .B1(REG2_REG_8__SCAN_IN), .B2(n4507), .ZN(n4505) );
  INV_X1 U4991 ( .A(n4499), .ZN(n4500) );
  AOI22_X1 U4992 ( .A1(n4503), .A2(n4502), .B1(n4501), .B2(n4500), .ZN(n4504)
         );
  OAI211_X1 U4993 ( .C1(n4507), .C2(n4506), .A(n4505), .B(n4504), .ZN(U3282)
         );
  AND2_X1 U4994 ( .A1(D_REG_31__SCAN_IN), .A2(n4517), .ZN(U3291) );
  NOR2_X1 U4995 ( .A1(n4516), .A2(n4508), .ZN(U3292) );
  NOR2_X1 U4996 ( .A1(n4516), .A2(n4509), .ZN(U3293) );
  NOR2_X1 U4997 ( .A1(n4516), .A2(n4510), .ZN(U3294) );
  AND2_X1 U4998 ( .A1(D_REG_27__SCAN_IN), .A2(n4517), .ZN(U3295) );
  AND2_X1 U4999 ( .A1(D_REG_26__SCAN_IN), .A2(n4517), .ZN(U3296) );
  AND2_X1 U5000 ( .A1(D_REG_25__SCAN_IN), .A2(n4517), .ZN(U3297) );
  AND2_X1 U5001 ( .A1(D_REG_24__SCAN_IN), .A2(n4517), .ZN(U3298) );
  AND2_X1 U5002 ( .A1(D_REG_23__SCAN_IN), .A2(n4517), .ZN(U3299) );
  AND2_X1 U5003 ( .A1(D_REG_22__SCAN_IN), .A2(n4517), .ZN(U3300) );
  AND2_X1 U5004 ( .A1(D_REG_21__SCAN_IN), .A2(n4517), .ZN(U3301) );
  AND2_X1 U5005 ( .A1(D_REG_20__SCAN_IN), .A2(n4517), .ZN(U3302) );
  NOR2_X1 U5006 ( .A1(n4516), .A2(n4511), .ZN(U3303) );
  AND2_X1 U5007 ( .A1(D_REG_18__SCAN_IN), .A2(n4517), .ZN(U3304) );
  AND2_X1 U5008 ( .A1(D_REG_17__SCAN_IN), .A2(n4517), .ZN(U3305) );
  AND2_X1 U5009 ( .A1(D_REG_16__SCAN_IN), .A2(n4517), .ZN(U3306) );
  AND2_X1 U5010 ( .A1(D_REG_15__SCAN_IN), .A2(n4517), .ZN(U3307) );
  AND2_X1 U5011 ( .A1(D_REG_14__SCAN_IN), .A2(n4517), .ZN(U3308) );
  AND2_X1 U5012 ( .A1(D_REG_13__SCAN_IN), .A2(n4517), .ZN(U3309) );
  AND2_X1 U5013 ( .A1(D_REG_12__SCAN_IN), .A2(n4517), .ZN(U3310) );
  AND2_X1 U5014 ( .A1(D_REG_11__SCAN_IN), .A2(n4517), .ZN(U3311) );
  NOR2_X1 U5015 ( .A1(n4516), .A2(n4512), .ZN(U3312) );
  AND2_X1 U5016 ( .A1(D_REG_9__SCAN_IN), .A2(n4517), .ZN(U3313) );
  AND2_X1 U5017 ( .A1(D_REG_8__SCAN_IN), .A2(n4517), .ZN(U3314) );
  AND2_X1 U5018 ( .A1(D_REG_7__SCAN_IN), .A2(n4517), .ZN(U3315) );
  NOR2_X1 U5019 ( .A1(n4516), .A2(n4513), .ZN(U3316) );
  NOR2_X1 U5020 ( .A1(n4516), .A2(n4514), .ZN(U3317) );
  AND2_X1 U5021 ( .A1(D_REG_4__SCAN_IN), .A2(n4517), .ZN(U3318) );
  NOR2_X1 U5022 ( .A1(n4516), .A2(n4515), .ZN(U3319) );
  AND2_X1 U5023 ( .A1(D_REG_2__SCAN_IN), .A2(n4517), .ZN(U3320) );
  INV_X1 U5024 ( .A(DATAI_23_), .ZN(n4519) );
  AOI21_X1 U5025 ( .B1(U3149), .B2(n4519), .A(n4518), .ZN(U3329) );
  AOI22_X1 U5026 ( .A1(STATE_REG_SCAN_IN), .A2(n4521), .B1(n4520), .B2(U3149), 
        .ZN(U3334) );
  AOI22_X1 U5027 ( .A1(STATE_REG_SCAN_IN), .A2(n4522), .B1(n2437), .B2(U3149), 
        .ZN(U3335) );
  INV_X1 U5028 ( .A(DATAI_16_), .ZN(n4523) );
  AOI22_X1 U5029 ( .A1(STATE_REG_SCAN_IN), .A2(n4524), .B1(n4523), .B2(U3149), 
        .ZN(U3336) );
  AOI22_X1 U5030 ( .A1(STATE_REG_SCAN_IN), .A2(n4526), .B1(n4525), .B2(U3149), 
        .ZN(U3337) );
  INV_X1 U5031 ( .A(DATAI_14_), .ZN(n4527) );
  AOI22_X1 U5032 ( .A1(STATE_REG_SCAN_IN), .A2(n3798), .B1(n4527), .B2(U3149), 
        .ZN(U3338) );
  AOI22_X1 U5033 ( .A1(STATE_REG_SCAN_IN), .A2(n4529), .B1(n4528), .B2(U3149), 
        .ZN(U3340) );
  INV_X1 U5034 ( .A(DATAI_11_), .ZN(n4530) );
  AOI22_X1 U5035 ( .A1(STATE_REG_SCAN_IN), .A2(n4531), .B1(n4530), .B2(U3149), 
        .ZN(U3341) );
  INV_X1 U5036 ( .A(DATAI_10_), .ZN(n4532) );
  AOI22_X1 U5037 ( .A1(STATE_REG_SCAN_IN), .A2(n4533), .B1(n4532), .B2(U3149), 
        .ZN(U3342) );
  AOI22_X1 U5038 ( .A1(STATE_REG_SCAN_IN), .A2(n4534), .B1(n4214), .B2(U3149), 
        .ZN(U3344) );
  INV_X1 U5039 ( .A(DATAI_6_), .ZN(n4535) );
  AOI22_X1 U5040 ( .A1(STATE_REG_SCAN_IN), .A2(n4536), .B1(n4535), .B2(U3149), 
        .ZN(U3346) );
  INV_X1 U5041 ( .A(DATAI_0_), .ZN(n4537) );
  AOI22_X1 U5042 ( .A1(STATE_REG_SCAN_IN), .A2(n2132), .B1(n4537), .B2(U3149), 
        .ZN(U3352) );
  INV_X1 U5043 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4538) );
  AOI22_X1 U5044 ( .A1(n4577), .A2(n4539), .B1(n4538), .B2(n4575), .ZN(U3467)
         );
  NOR2_X1 U5045 ( .A1(n4540), .A2(n4559), .ZN(n4542) );
  AOI211_X1 U5046 ( .C1(n4543), .C2(n4554), .A(n4542), .B(n4541), .ZN(n4578)
         );
  INV_X1 U5047 ( .A(REG0_REG_1__SCAN_IN), .ZN(n4544) );
  AOI22_X1 U5048 ( .A1(n4577), .A2(n4578), .B1(n4544), .B2(n4575), .ZN(U3469)
         );
  NOR2_X1 U5049 ( .A1(n4546), .A2(n4545), .ZN(n4548) );
  AOI211_X1 U5050 ( .C1(n4574), .C2(n4549), .A(n4548), .B(n4547), .ZN(n4580)
         );
  INV_X1 U5051 ( .A(REG0_REG_3__SCAN_IN), .ZN(n4550) );
  AOI22_X1 U5052 ( .A1(n4577), .A2(n4580), .B1(n4550), .B2(n4575), .ZN(U3473)
         );
  INV_X1 U5053 ( .A(n4551), .ZN(n4553) );
  AOI211_X1 U5054 ( .C1(n4555), .C2(n4554), .A(n4553), .B(n4552), .ZN(n4581)
         );
  INV_X1 U5055 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4556) );
  AOI22_X1 U5056 ( .A1(n4577), .A2(n4581), .B1(n4556), .B2(n4575), .ZN(U3475)
         );
  OAI21_X1 U5057 ( .B1(n4559), .B2(n4558), .A(n4557), .ZN(n4560) );
  AOI21_X1 U5058 ( .B1(n4562), .B2(n4561), .A(n4560), .ZN(n4583) );
  INV_X1 U5059 ( .A(REG0_REG_5__SCAN_IN), .ZN(n4563) );
  AOI22_X1 U5060 ( .A1(n4577), .A2(n4583), .B1(n4563), .B2(n4575), .ZN(U3477)
         );
  NOR2_X1 U5061 ( .A1(n4564), .A2(n4569), .ZN(n4567) );
  AOI211_X1 U5062 ( .C1(n4567), .C2(n2963), .A(n4566), .B(n4565), .ZN(n4585)
         );
  INV_X1 U5063 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4568) );
  AOI22_X1 U5064 ( .A1(n4577), .A2(n4585), .B1(n4568), .B2(n4575), .ZN(U3481)
         );
  NOR2_X1 U5065 ( .A1(n4570), .A2(n4569), .ZN(n4572) );
  AOI211_X1 U5066 ( .C1(n4574), .C2(n4573), .A(n4572), .B(n4571), .ZN(n4587)
         );
  AOI22_X1 U5067 ( .A1(n4577), .A2(n4587), .B1(n4576), .B2(n4575), .ZN(U3485)
         );
  AOI22_X1 U5068 ( .A1(n4588), .A2(n4578), .B1(n2663), .B2(n4586), .ZN(U3519)
         );
  INV_X1 U5069 ( .A(REG1_REG_3__SCAN_IN), .ZN(n4579) );
  AOI22_X1 U5070 ( .A1(n4588), .A2(n4580), .B1(n4579), .B2(n4586), .ZN(U3521)
         );
  AOI22_X1 U5071 ( .A1(n4588), .A2(n4581), .B1(n4374), .B2(n4586), .ZN(U3522)
         );
  AOI22_X1 U5072 ( .A1(n4588), .A2(n4583), .B1(n4582), .B2(n4586), .ZN(U3523)
         );
  AOI22_X1 U5073 ( .A1(n4588), .A2(n4585), .B1(n4584), .B2(n4586), .ZN(U3525)
         );
  AOI22_X1 U5074 ( .A1(n4588), .A2(n4587), .B1(n2808), .B2(n4586), .ZN(U3527)
         );
  INV_X4 U2258 ( .A(n2003), .ZN(n2007) );
  CLKBUF_X1 U2324 ( .A(n2284), .Z(n3611) );
endmodule

