

module b17_C_2inp_gates_syn ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, 
        DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, 
        DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, 
        DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, 
        DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, 
        DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, 
        READY1, READY2, P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN, 
        P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN, 
        P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN, 
        P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN, 
        P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN, 
        P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN, 
        P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN, 
        P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN, 
        P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN, 
        P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN, 
        P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN, 
        P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN, 
        P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN, 
        P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN, 
        P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN, 
        P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN, 
        P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN, 
        P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, 
        P1_REIP_REG_6__SCAN_IN, P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, 
        P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, 
        P1_REIP_REG_0__SCAN_IN, P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, 
        P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, 
        P1_EBX_REG_26__SCAN_IN, P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, 
        P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, 
        P1_EBX_REG_20__SCAN_IN, P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, 
        P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, 
        P1_EBX_REG_14__SCAN_IN, P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, 
        P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, 
        P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, 
        P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, 
        P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, 
        P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, 
        P1_EAX_REG_28__SCAN_IN, P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, 
        P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, 
        P1_EAX_REG_22__SCAN_IN, P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, 
        P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, 
        P1_EAX_REG_16__SCAN_IN, P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, 
        P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, 
        P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, 
        P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, 
        P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, 
        P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, U355, 
        U356, U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, 
        U369, U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, 
        U352, U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, 
        U240, U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, 
        U228, U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, 
        U216, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, 
        U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, 
        U274, U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, 
        U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, 
        P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, 
        P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, 
        P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, 
        P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, 
        P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, 
        P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, 
        P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, 
        P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, 
        P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, 
        P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, 
        P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, 
        P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, 
        P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, 
        P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, 
        P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, 
        P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, 
        P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, 
        P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, 
        P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, 
        P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, 
        P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, 
        P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, 
        P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, 
        P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, 
        P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, 
        P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, 
        P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, 
        P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, 
        P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, 
        P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, 
        P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, 
        P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, 
        P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, 
        P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, 
        P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, 
        P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, 
        P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, 
        P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, 
        P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, 
        P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, 
        P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, 
        P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, 
        P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, 
        P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, 
        P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, 
        P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, 
        P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, 
        P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, 
        P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, 
        P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, 
        P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, 
        P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, 
        P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, 
        P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, 
        P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, 
        P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, 
        P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, 
        P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, 
        P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, 
        P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, 
        P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, 
        P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, 
        P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, 
        P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, 
        P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, 
        P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, 
        P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, 
        P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, 
        P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, 
        P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, 
        P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, 
        P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, 
        P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, 
        P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, 
        P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, 
        P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, 
        P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, 
        P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, 
        P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, 
        P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, 
        P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, 
        P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, 
        P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, 
        P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, 
        P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, 
        P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, 
        P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, 
        P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, 
        P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, 
        P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, 
        P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, 
        P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, 
        P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, 
        P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, 
        P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, 
        P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, 
        P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, 
        P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, 
        P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, 
        P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, 
        P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, 
        P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, 
        P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, 
        P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, 
        P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, 
        P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, 
        P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, 
        P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, 
        P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, 
        P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, 
        P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, 
        P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, 
        P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, 
        P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, 
        P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, 
        P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, 
        P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, 
        P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, 
        P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, 
        P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, 
        P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, 
        P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, 
        P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, 
        P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, 
        P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, 
        P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, 
        P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, 
        P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, 
        P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, 
        P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, 
        P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, 
        P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, 
        P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, 
        P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, 
        P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, 
        P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, 
        P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, 
        P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, 
        P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, 
        P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, 
        P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, 
        P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, 
        P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, 
        P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, 
        P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, 
        P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, 
        P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, 
        P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, 
        P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, 
        P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, 
        P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, 
        P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, 
        P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, 
        P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, 
        P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, 
        P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, 
        P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, 
        P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, 
        P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, 
        P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, 
        P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, 
        P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, 
        P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, 
        P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, 
        P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, 
        P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, 
        P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, 
        P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, 
        P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, 
        P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, 
        P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, 
        P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, 
        P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, 
        P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, 
        P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, 
        P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, 
        P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, 
        P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, 
        P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, 
        P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, 
        P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, 
        P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, 
        P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, 
        P1_U2803, P1_U2802, P1_U3487, P1_U2801, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput0, keyinput1, keyinput2,
         keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8,
         keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9718, n9719,
         n9720, n9721, n9722, n9723, n9724, n9726, n9727, n9729, n9730, n9731,
         n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741,
         n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751,
         n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761,
         n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771,
         n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781,
         n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791,
         n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801,
         n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811,
         n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821,
         n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831,
         n9832, n9833, n9834, n9835, n9836, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9880, n9881, n9882, n9883,
         n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893,
         n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903,
         n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913,
         n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923,
         n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933,
         n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943,
         n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953,
         n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963,
         n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973,
         n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983,
         n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993,
         n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002,
         n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010,
         n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018,
         n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026,
         n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034,
         n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042,
         n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050,
         n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058,
         n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066,
         n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074,
         n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082,
         n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090,
         n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098,
         n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106,
         n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114,
         n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122,
         n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130,
         n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138,
         n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146,
         n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154,
         n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162,
         n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170,
         n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178,
         n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186,
         n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194,
         n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202,
         n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210,
         n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218,
         n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226,
         n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234,
         n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242,
         n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250,
         n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258,
         n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266,
         n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274,
         n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282,
         n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290,
         n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298,
         n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306,
         n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314,
         n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322,
         n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330,
         n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338,
         n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346,
         n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354,
         n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10363,
         n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371,
         n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379,
         n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387,
         n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395,
         n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403,
         n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411,
         n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419,
         n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427,
         n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435,
         n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443,
         n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451,
         n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459,
         n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467,
         n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475,
         n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483,
         n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491,
         n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499,
         n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507,
         n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515,
         n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523,
         n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531,
         n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539,
         n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547,
         n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555,
         n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563,
         n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571,
         n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579,
         n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587,
         n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595,
         n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603,
         n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611,
         n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619,
         n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627,
         n10628, n10629, n10630, n10631, n10632, n10633, n10634, n10635,
         n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643,
         n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651,
         n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659,
         n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667,
         n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675,
         n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683,
         n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691,
         n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699,
         n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707,
         n10708, n10709, n10710, n10711, n10712, n10713, n10714, n10715,
         n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723,
         n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731,
         n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739,
         n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747,
         n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755,
         n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763,
         n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771,
         n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779,
         n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787,
         n10788, n10789, n10790, n10791, n10792, n10793, n10794, n10795,
         n10796, n10797, n10798, n10799, n10800, n10801, n10802, n10803,
         n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811,
         n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819,
         n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827,
         n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835,
         n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843,
         n10844, n10845, n10846, n10847, n10848, n10849, n10850, n10851,
         n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859,
         n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867,
         n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875,
         n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883,
         n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891,
         n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899,
         n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907,
         n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915,
         n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923,
         n10924, n10925, n10926, n10927, n10928, n10929, n10930, n10931,
         n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939,
         n10940, n10941, n10942, n10943, n10944, n10945, n10946, n10947,
         n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955,
         n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963,
         n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971,
         n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979,
         n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987,
         n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995,
         n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003,
         n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11011,
         n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019,
         n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027,
         n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035,
         n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043,
         n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051,
         n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059,
         n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067,
         n11068, n11069, n11070, n11071, n11072, n11073, n11074, n11075,
         n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083,
         n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091,
         n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099,
         n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107,
         n11108, n11109, n11110, n11111, n11112, n11113, n11114, n11115,
         n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123,
         n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131,
         n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139,
         n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147,
         n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155,
         n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163,
         n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171,
         n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179,
         n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187,
         n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195,
         n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203,
         n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211,
         n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219,
         n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227,
         n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235,
         n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243,
         n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251,
         n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259,
         n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267,
         n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275,
         n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283,
         n11284, n11285, n11286, n11287, n11288, n11289, n11290, n11291,
         n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299,
         n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307,
         n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315,
         n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323,
         n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331,
         n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339,
         n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347,
         n11348, n11349, n11350, n11351, n11352, n11353, n11354, n11355,
         n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363,
         n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371,
         n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379,
         n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387,
         n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395,
         n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403,
         n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411,
         n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419,
         n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427,
         n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435,
         n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443,
         n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451,
         n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459,
         n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467,
         n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475,
         n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483,
         n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491,
         n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499,
         n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507,
         n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515,
         n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523,
         n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531,
         n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539,
         n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547,
         n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555,
         n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563,
         n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571,
         n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579,
         n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587,
         n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11595,
         n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603,
         n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611,
         n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619,
         n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627,
         n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635,
         n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643,
         n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651,
         n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659,
         n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667,
         n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675,
         n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683,
         n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691,
         n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699,
         n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707,
         n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715,
         n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723,
         n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731,
         n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739,
         n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747,
         n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755,
         n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11763,
         n11764, n11765, n11766, n11767, n11768, n11769, n11770, n11771,
         n11772, n11773, n11774, n11775, n11776, n11777, n11778, n11779,
         n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787,
         n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795,
         n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803,
         n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811,
         n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819,
         n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827,
         n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835,
         n11836, n11837, n11838, n11839, n11840, n11841, n11842, n11843,
         n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851,
         n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859,
         n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867,
         n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875,
         n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883,
         n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891,
         n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899,
         n11900, n11901, n11902, n11903, n11904, n11905, n11906, n11907,
         n11908, n11909, n11910, n11911, n11912, n11913, n11914, n11915,
         n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923,
         n11924, n11925, n11926, n11927, n11928, n11929, n11930, n11931,
         n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939,
         n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947,
         n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955,
         n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963,
         n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971,
         n11972, n11973, n11974, n11975, n11976, n11977, n11978, n11979,
         n11980, n11981, n11982, n11983, n11984, n11985, n11986, n11987,
         n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995,
         n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003,
         n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011,
         n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019,
         n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027,
         n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035,
         n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043,
         n12044, n12045, n12046, n12047, n12048, n12049, n12050, n12051,
         n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12059,
         n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067,
         n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12075,
         n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083,
         n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091,
         n12092, n12093, n12094, n12095, n12096, n12097, n12098, n12099,
         n12100, n12101, n12102, n12103, n12104, n12105, n12106, n12107,
         n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115,
         n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123,
         n12124, n12125, n12126, n12127, n12128, n12129, n12130, n12131,
         n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139,
         n12140, n12141, n12142, n12143, n12144, n12145, n12146, n12147,
         n12148, n12149, n12150, n12151, n12152, n12153, n12154, n12155,
         n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163,
         n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12171,
         n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179,
         n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187,
         n12188, n12189, n12190, n12191, n12192, n12193, n12194, n12195,
         n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203,
         n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211,
         n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219,
         n12220, n12221, n12222, n12223, n12224, n12225, n12226, n12227,
         n12228, n12229, n12230, n12231, n12232, n12233, n12234, n12235,
         n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243,
         n12244, n12245, n12246, n12247, n12248, n12249, n12250, n12251,
         n12252, n12253, n12254, n12255, n12256, n12257, n12258, n12259,
         n12260, n12261, n12262, n12263, n12264, n12265, n12266, n12267,
         n12268, n12269, n12270, n12271, n12272, n12273, n12274, n12275,
         n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283,
         n12284, n12285, n12286, n12287, n12288, n12289, n12290, n12291,
         n12292, n12293, n12294, n12295, n12296, n12297, n12298, n12299,
         n12300, n12301, n12302, n12303, n12304, n12305, n12306, n12307,
         n12308, n12309, n12310, n12311, n12312, n12313, n12314, n12315,
         n12316, n12317, n12318, n12319, n12320, n12321, n12322, n12323,
         n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331,
         n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12339,
         n12340, n12341, n12342, n12343, n12344, n12345, n12346, n12347,
         n12348, n12349, n12350, n12351, n12352, n12353, n12354, n12355,
         n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363,
         n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371,
         n12372, n12373, n12374, n12375, n12376, n12377, n12378, n12379,
         n12380, n12381, n12382, n12383, n12384, n12385, n12386, n12387,
         n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395,
         n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403,
         n12404, n12405, n12406, n12407, n12408, n12409, n12410, n12411,
         n12412, n12413, n12414, n12415, n12416, n12417, n12418, n12419,
         n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427,
         n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435,
         n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12443,
         n12444, n12445, n12446, n12447, n12448, n12449, n12450, n12451,
         n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459,
         n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467,
         n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475,
         n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483,
         n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491,
         n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499,
         n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507,
         n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515,
         n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523,
         n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531,
         n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539,
         n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547,
         n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555,
         n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563,
         n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571,
         n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579,
         n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587,
         n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595,
         n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603,
         n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611,
         n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619,
         n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627,
         n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635,
         n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643,
         n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651,
         n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659,
         n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667,
         n12668, n12669, n12670, n12671, n12672, n12673, n12674, n12675,
         n12676, n12677, n12678, n12679, n12680, n12681, n12682, n12683,
         n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691,
         n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699,
         n12702, n12703, n12704, n12705, n12706, n12707, n12708, n12709,
         n12710, n12711, n12712, n12713, n12714, n12715, n12716, n12717,
         n12718, n12719, n12720, n12721, n12722, n12723, n12724, n12725,
         n12726, n12727, n12728, n12729, n12730, n12731, n12732, n12733,
         n12734, n12735, n12736, n12737, n12738, n12739, n12740, n12741,
         n12742, n12743, n12744, n12745, n12746, n12747, n12748, n12749,
         n12750, n12751, n12752, n12753, n12754, n12755, n12756, n12757,
         n12758, n12759, n12760, n12761, n12762, n12763, n12764, n12765,
         n12766, n12767, n12768, n12769, n12770, n12771, n12772, n12773,
         n12774, n12775, n12776, n12777, n12778, n12779, n12780, n12781,
         n12782, n12783, n12784, n12785, n12786, n12787, n12788, n12789,
         n12790, n12791, n12792, n12793, n12794, n12795, n12796, n12797,
         n12798, n12799, n12800, n12801, n12802, n12803, n12804, n12805,
         n12806, n12807, n12808, n12809, n12810, n12811, n12812, n12813,
         n12814, n12815, n12816, n12817, n12818, n12819, n12820, n12821,
         n12822, n12823, n12824, n12825, n12826, n12827, n12828, n12829,
         n12830, n12831, n12832, n12833, n12834, n12835, n12836, n12837,
         n12838, n12839, n12840, n12841, n12842, n12843, n12844, n12845,
         n12846, n12847, n12848, n12849, n12850, n12851, n12852, n12853,
         n12854, n12855, n12856, n12857, n12858, n12859, n12860, n12861,
         n12862, n12863, n12864, n12865, n12866, n12867, n12868, n12869,
         n12870, n12871, n12872, n12873, n12874, n12875, n12876, n12877,
         n12878, n12879, n12880, n12881, n12882, n12883, n12884, n12885,
         n12886, n12887, n12888, n12889, n12890, n12891, n12892, n12893,
         n12894, n12895, n12896, n12897, n12898, n12899, n12900, n12901,
         n12902, n12903, n12904, n12905, n12906, n12907, n12908, n12909,
         n12910, n12911, n12912, n12913, n12914, n12915, n12916, n12917,
         n12918, n12919, n12920, n12921, n12922, n12923, n12924, n12925,
         n12926, n12927, n12928, n12929, n12930, n12931, n12932, n12933,
         n12934, n12935, n12936, n12937, n12938, n12939, n12940, n12941,
         n12942, n12943, n12944, n12945, n12946, n12947, n12948, n12949,
         n12950, n12951, n12952, n12953, n12954, n12955, n12956, n12957,
         n12958, n12959, n12960, n12961, n12962, n12963, n12964, n12965,
         n12966, n12967, n12968, n12969, n12970, n12971, n12972, n12973,
         n12974, n12975, n12976, n12977, n12978, n12979, n12980, n12981,
         n12982, n12983, n12984, n12985, n12986, n12987, n12988, n12989,
         n12990, n12991, n12992, n12993, n12994, n12995, n12996, n12997,
         n12998, n12999, n13000, n13001, n13002, n13003, n13004, n13005,
         n13006, n13007, n13008, n13009, n13010, n13011, n13012, n13013,
         n13014, n13015, n13016, n13017, n13018, n13019, n13020, n13021,
         n13022, n13023, n13024, n13025, n13026, n13027, n13028, n13029,
         n13030, n13031, n13032, n13033, n13034, n13035, n13036, n13037,
         n13038, n13039, n13040, n13041, n13042, n13043, n13044, n13045,
         n13046, n13047, n13048, n13049, n13050, n13051, n13052, n13053,
         n13054, n13055, n13056, n13057, n13058, n13059, n13060, n13061,
         n13062, n13063, n13064, n13065, n13066, n13067, n13068, n13069,
         n13070, n13071, n13072, n13073, n13074, n13075, n13076, n13077,
         n13078, n13079, n13080, n13081, n13082, n13083, n13084, n13085,
         n13086, n13087, n13088, n13089, n13090, n13091, n13092, n13093,
         n13094, n13095, n13096, n13097, n13098, n13099, n13100, n13101,
         n13102, n13103, n13104, n13105, n13106, n13107, n13108, n13109,
         n13110, n13111, n13112, n13113, n13114, n13115, n13116, n13117,
         n13118, n13119, n13120, n13121, n13122, n13123, n13124, n13125,
         n13126, n13127, n13128, n13129, n13130, n13131, n13132, n13133,
         n13134, n13135, n13136, n13137, n13138, n13139, n13140, n13141,
         n13142, n13143, n13144, n13145, n13146, n13147, n13148, n13149,
         n13150, n13151, n13152, n13153, n13154, n13155, n13156, n13157,
         n13158, n13159, n13160, n13161, n13162, n13163, n13164, n13165,
         n13166, n13167, n13168, n13169, n13170, n13171, n13172, n13173,
         n13174, n13175, n13176, n13177, n13178, n13179, n13180, n13181,
         n13182, n13183, n13184, n13185, n13186, n13187, n13188, n13189,
         n13190, n13191, n13192, n13193, n13194, n13195, n13196, n13197,
         n13198, n13199, n13200, n13201, n13202, n13203, n13204, n13205,
         n13206, n13207, n13208, n13209, n13210, n13211, n13212, n13213,
         n13214, n13215, n13216, n13217, n13218, n13219, n13220, n13221,
         n13222, n13223, n13224, n13225, n13226, n13227, n13228, n13229,
         n13230, n13231, n13232, n13233, n13234, n13235, n13236, n13237,
         n13238, n13239, n13240, n13241, n13242, n13243, n13244, n13245,
         n13246, n13247, n13248, n13249, n13250, n13251, n13252, n13253,
         n13254, n13255, n13256, n13257, n13258, n13259, n13260, n13261,
         n13262, n13263, n13264, n13265, n13266, n13267, n13268, n13269,
         n13270, n13271, n13272, n13273, n13274, n13275, n13276, n13277,
         n13278, n13279, n13280, n13281, n13282, n13283, n13284, n13285,
         n13286, n13287, n13288, n13289, n13290, n13291, n13292, n13293,
         n13294, n13295, n13296, n13297, n13298, n13299, n13300, n13301,
         n13302, n13303, n13304, n13305, n13306, n13307, n13308, n13309,
         n13310, n13311, n13312, n13313, n13314, n13315, n13316, n13317,
         n13318, n13319, n13320, n13321, n13322, n13323, n13324, n13325,
         n13326, n13327, n13328, n13329, n13330, n13331, n13332, n13333,
         n13334, n13335, n13336, n13337, n13338, n13339, n13340, n13341,
         n13342, n13343, n13344, n13345, n13346, n13347, n13348, n13349,
         n13350, n13351, n13352, n13353, n13354, n13355, n13356, n13357,
         n13358, n13359, n13360, n13361, n13362, n13363, n13364, n13365,
         n13366, n13367, n13368, n13369, n13370, n13371, n13372, n13373,
         n13374, n13375, n13376, n13377, n13378, n13379, n13380, n13381,
         n13382, n13383, n13384, n13385, n13386, n13387, n13388, n13389,
         n13390, n13391, n13392, n13393, n13394, n13395, n13396, n13397,
         n13398, n13399, n13400, n13401, n13402, n13403, n13404, n13405,
         n13406, n13407, n13408, n13409, n13410, n13411, n13412, n13413,
         n13414, n13415, n13416, n13417, n13418, n13419, n13420, n13421,
         n13422, n13423, n13424, n13425, n13426, n13427, n13428, n13429,
         n13430, n13431, n13432, n13433, n13434, n13435, n13436, n13437,
         n13438, n13439, n13440, n13441, n13442, n13443, n13444, n13445,
         n13446, n13447, n13448, n13449, n13450, n13451, n13452, n13453,
         n13454, n13455, n13456, n13457, n13458, n13459, n13460, n13461,
         n13462, n13463, n13464, n13465, n13466, n13467, n13468, n13469,
         n13470, n13471, n13472, n13473, n13474, n13475, n13476, n13477,
         n13478, n13479, n13480, n13481, n13482, n13483, n13484, n13485,
         n13486, n13487, n13488, n13489, n13490, n13491, n13492, n13493,
         n13494, n13495, n13496, n13497, n13498, n13499, n13500, n13501,
         n13502, n13503, n13504, n13505, n13506, n13507, n13508, n13509,
         n13510, n13511, n13512, n13513, n13514, n13515, n13516, n13517,
         n13518, n13519, n13520, n13521, n13522, n13523, n13524, n13525,
         n13526, n13527, n13528, n13529, n13530, n13531, n13532, n13533,
         n13534, n13535, n13536, n13537, n13538, n13539, n13540, n13541,
         n13542, n13543, n13544, n13545, n13546, n13547, n13548, n13549,
         n13550, n13551, n13552, n13553, n13554, n13555, n13556, n13557,
         n13558, n13559, n13560, n13561, n13562, n13563, n13564, n13565,
         n13566, n13567, n13568, n13569, n13570, n13571, n13572, n13573,
         n13574, n13575, n13576, n13577, n13578, n13579, n13580, n13581,
         n13582, n13583, n13584, n13585, n13586, n13587, n13588, n13589,
         n13590, n13591, n13592, n13593, n13594, n13595, n13596, n13597,
         n13598, n13599, n13600, n13601, n13602, n13603, n13604, n13605,
         n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613,
         n13614, n13615, n13616, n13617, n13618, n13619, n13620, n13621,
         n13622, n13623, n13624, n13625, n13626, n13627, n13628, n13629,
         n13630, n13631, n13632, n13633, n13634, n13635, n13636, n13637,
         n13638, n13639, n13640, n13641, n13642, n13643, n13644, n13645,
         n13646, n13647, n13648, n13649, n13650, n13651, n13652, n13653,
         n13654, n13655, n13656, n13657, n13658, n13659, n13660, n13661,
         n13662, n13663, n13664, n13665, n13666, n13667, n13668, n13669,
         n13670, n13671, n13672, n13673, n13674, n13675, n13676, n13677,
         n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685,
         n13686, n13687, n13688, n13689, n13690, n13691, n13692, n13693,
         n13694, n13695, n13696, n13697, n13698, n13699, n13700, n13701,
         n13702, n13703, n13704, n13705, n13706, n13707, n13708, n13709,
         n13710, n13711, n13712, n13713, n13714, n13715, n13716, n13717,
         n13718, n13719, n13720, n13721, n13722, n13723, n13724, n13725,
         n13726, n13727, n13728, n13729, n13730, n13731, n13732, n13733,
         n13734, n13735, n13736, n13737, n13738, n13739, n13740, n13741,
         n13742, n13743, n13744, n13745, n13746, n13747, n13748, n13749,
         n13750, n13751, n13752, n13753, n13754, n13755, n13756, n13757,
         n13758, n13759, n13760, n13761, n13762, n13763, n13764, n13765,
         n13766, n13767, n13768, n13769, n13770, n13771, n13772, n13773,
         n13774, n13775, n13776, n13777, n13778, n13779, n13780, n13781,
         n13782, n13783, n13784, n13785, n13786, n13787, n13788, n13789,
         n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797,
         n13798, n13799, n13800, n13801, n13802, n13803, n13804, n13805,
         n13806, n13807, n13808, n13809, n13810, n13811, n13812, n13813,
         n13814, n13815, n13816, n13817, n13818, n13819, n13820, n13821,
         n13822, n13823, n13824, n13825, n13826, n13827, n13828, n13829,
         n13830, n13831, n13832, n13833, n13834, n13835, n13836, n13837,
         n13838, n13839, n13840, n13841, n13842, n13843, n13844, n13845,
         n13846, n13847, n13848, n13849, n13850, n13851, n13852, n13853,
         n13854, n13855, n13856, n13857, n13858, n13859, n13860, n13861,
         n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869,
         n13870, n13871, n13872, n13873, n13874, n13875, n13876, n13877,
         n13878, n13879, n13880, n13881, n13882, n13883, n13884, n13885,
         n13886, n13887, n13888, n13889, n13890, n13891, n13892, n13893,
         n13894, n13895, n13896, n13897, n13898, n13899, n13900, n13901,
         n13902, n13903, n13904, n13905, n13906, n13907, n13908, n13909,
         n13910, n13911, n13912, n13913, n13914, n13915, n13916, n13917,
         n13918, n13919, n13920, n13921, n13922, n13923, n13924, n13925,
         n13926, n13927, n13928, n13929, n13930, n13931, n13932, n13933,
         n13934, n13935, n13936, n13937, n13938, n13939, n13940, n13941,
         n13942, n13943, n13944, n13945, n13946, n13947, n13948, n13949,
         n13950, n13951, n13952, n13953, n13954, n13955, n13956, n13957,
         n13958, n13959, n13960, n13961, n13962, n13963, n13964, n13965,
         n13966, n13967, n13968, n13969, n13970, n13971, n13972, n13973,
         n13974, n13975, n13976, n13977, n13978, n13979, n13980, n13981,
         n13982, n13983, n13984, n13985, n13986, n13987, n13988, n13989,
         n13990, n13991, n13992, n13993, n13994, n13995, n13996, n13997,
         n13998, n13999, n14000, n14001, n14002, n14003, n14004, n14005,
         n14006, n14007, n14008, n14009, n14010, n14011, n14012, n14013,
         n14014, n14015, n14016, n14017, n14018, n14019, n14020, n14021,
         n14022, n14023, n14024, n14025, n14026, n14027, n14028, n14029,
         n14030, n14031, n14032, n14033, n14034, n14035, n14036, n14037,
         n14038, n14039, n14040, n14041, n14042, n14043, n14044, n14045,
         n14046, n14047, n14048, n14049, n14050, n14051, n14052, n14053,
         n14054, n14055, n14056, n14057, n14058, n14059, n14060, n14061,
         n14062, n14063, n14064, n14065, n14066, n14067, n14068, n14069,
         n14070, n14071, n14072, n14073, n14074, n14075, n14076, n14077,
         n14078, n14079, n14080, n14081, n14082, n14083, n14084, n14085,
         n14086, n14087, n14088, n14089, n14090, n14091, n14092, n14093,
         n14094, n14095, n14096, n14097, n14098, n14099, n14100, n14101,
         n14102, n14103, n14104, n14105, n14106, n14107, n14108, n14109,
         n14110, n14111, n14112, n14113, n14114, n14115, n14116, n14117,
         n14118, n14119, n14120, n14121, n14122, n14123, n14124, n14125,
         n14126, n14127, n14128, n14129, n14130, n14131, n14132, n14133,
         n14134, n14135, n14136, n14137, n14138, n14139, n14140, n14141,
         n14142, n14143, n14144, n14145, n14146, n14147, n14148, n14149,
         n14150, n14151, n14152, n14153, n14154, n14155, n14156, n14157,
         n14158, n14159, n14160, n14161, n14162, n14163, n14164, n14165,
         n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173,
         n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14181,
         n14182, n14183, n14184, n14185, n14186, n14187, n14188, n14189,
         n14190, n14191, n14192, n14193, n14194, n14195, n14196, n14197,
         n14198, n14199, n14200, n14201, n14202, n14203, n14204, n14205,
         n14206, n14207, n14208, n14209, n14210, n14211, n14212, n14213,
         n14214, n14215, n14216, n14217, n14218, n14219, n14220, n14221,
         n14222, n14223, n14224, n14225, n14226, n14227, n14228, n14229,
         n14230, n14231, n14232, n14233, n14234, n14235, n14236, n14237,
         n14238, n14239, n14240, n14241, n14242, n14243, n14244, n14245,
         n14246, n14247, n14248, n14249, n14250, n14251, n14252, n14253,
         n14254, n14255, n14256, n14257, n14258, n14259, n14260, n14261,
         n14262, n14263, n14264, n14265, n14266, n14267, n14268, n14269,
         n14270, n14271, n14272, n14273, n14274, n14275, n14276, n14277,
         n14278, n14279, n14280, n14281, n14282, n14283, n14284, n14285,
         n14286, n14287, n14288, n14289, n14290, n14291, n14292, n14293,
         n14294, n14295, n14296, n14297, n14298, n14299, n14300, n14301,
         n14302, n14303, n14304, n14305, n14306, n14307, n14308, n14309,
         n14310, n14311, n14312, n14313, n14314, n14315, n14316, n14317,
         n14318, n14319, n14320, n14321, n14322, n14323, n14324, n14325,
         n14326, n14327, n14328, n14329, n14330, n14331, n14332, n14333,
         n14334, n14335, n14336, n14337, n14338, n14339, n14340, n14341,
         n14342, n14343, n14344, n14345, n14346, n14347, n14348, n14349,
         n14350, n14351, n14352, n14353, n14354, n14355, n14356, n14357,
         n14358, n14359, n14360, n14361, n14362, n14363, n14364, n14365,
         n14366, n14367, n14368, n14369, n14370, n14371, n14372, n14373,
         n14374, n14375, n14376, n14377, n14378, n14379, n14380, n14381,
         n14382, n14383, n14384, n14385, n14386, n14387, n14388, n14389,
         n14390, n14391, n14392, n14393, n14394, n14395, n14396, n14397,
         n14398, n14399, n14400, n14401, n14402, n14403, n14404, n14405,
         n14406, n14407, n14408, n14409, n14410, n14411, n14412, n14413,
         n14414, n14415, n14416, n14417, n14418, n14419, n14420, n14421,
         n14422, n14423, n14424, n14425, n14426, n14427, n14428, n14429,
         n14430, n14431, n14432, n14433, n14434, n14435, n14436, n14437,
         n14438, n14439, n14440, n14441, n14442, n14443, n14444, n14445,
         n14446, n14447, n14448, n14449, n14450, n14451, n14452, n14453,
         n14454, n14455, n14456, n14457, n14458, n14459, n14460, n14461,
         n14462, n14463, n14464, n14465, n14466, n14467, n14468, n14469,
         n14470, n14471, n14472, n14473, n14474, n14475, n14476, n14477,
         n14478, n14479, n14480, n14481, n14482, n14483, n14484, n14485,
         n14486, n14487, n14488, n14489, n14490, n14491, n14492, n14493,
         n14494, n14495, n14496, n14497, n14498, n14499, n14500, n14501,
         n14502, n14503, n14504, n14505, n14506, n14507, n14508, n14509,
         n14510, n14511, n14512, n14513, n14514, n14515, n14516, n14517,
         n14518, n14519, n14520, n14521, n14522, n14523, n14524, n14525,
         n14526, n14527, n14528, n14529, n14530, n14531, n14532, n14533,
         n14534, n14535, n14536, n14537, n14538, n14539, n14540, n14541,
         n14542, n14543, n14544, n14545, n14546, n14547, n14548, n14549,
         n14550, n14551, n14552, n14553, n14554, n14555, n14556, n14557,
         n14558, n14559, n14560, n14561, n14562, n14563, n14564, n14565,
         n14566, n14567, n14568, n14569, n14570, n14571, n14572, n14573,
         n14574, n14575, n14576, n14577, n14578, n14579, n14580, n14581,
         n14582, n14583, n14584, n14585, n14586, n14587, n14588, n14589,
         n14590, n14591, n14592, n14593, n14594, n14595, n14596, n14597,
         n14598, n14599, n14600, n14601, n14602, n14603, n14604, n14605,
         n14606, n14607, n14608, n14609, n14610, n14611, n14612, n14613,
         n14614, n14615, n14616, n14617, n14618, n14619, n14620, n14621,
         n14622, n14623, n14624, n14625, n14626, n14627, n14628, n14629,
         n14630, n14631, n14632, n14633, n14634, n14635, n14636, n14637,
         n14638, n14639, n14640, n14641, n14642, n14643, n14644, n14645,
         n14646, n14647, n14648, n14649, n14650, n14651, n14652, n14653,
         n14654, n14655, n14656, n14657, n14658, n14659, n14660, n14661,
         n14662, n14663, n14664, n14665, n14666, n14667, n14668, n14669,
         n14670, n14671, n14672, n14673, n14674, n14675, n14676, n14677,
         n14678, n14679, n14680, n14681, n14682, n14683, n14684, n14685,
         n14686, n14687, n14688, n14689, n14690, n14691, n14692, n14693,
         n14694, n14695, n14696, n14697, n14698, n14699, n14700, n14701,
         n14702, n14703, n14704, n14705, n14706, n14707, n14708, n14709,
         n14710, n14711, n14712, n14713, n14714, n14715, n14716, n14717,
         n14718, n14719, n14720, n14721, n14722, n14723, n14724, n14725,
         n14726, n14727, n14728, n14729, n14730, n14731, n14732, n14733,
         n14734, n14735, n14736, n14737, n14738, n14739, n14740, n14741,
         n14742, n14743, n14744, n14745, n14746, n14747, n14748, n14749,
         n14750, n14751, n14752, n14753, n14754, n14755, n14756, n14757,
         n14758, n14759, n14760, n14761, n14762, n14763, n14764, n14765,
         n14766, n14767, n14768, n14769, n14770, n14771, n14772, n14773,
         n14774, n14775, n14776, n14777, n14778, n14779, n14780, n14781,
         n14782, n14783, n14784, n14785, n14786, n14787, n14788, n14789,
         n14790, n14791, n14792, n14793, n14794, n14795, n14796, n14797,
         n14798, n14799, n14800, n14801, n14802, n14803, n14804, n14805,
         n14806, n14807, n14808, n14809, n14810, n14811, n14812, n14813,
         n14814, n14815, n14816, n14817, n14818, n14819, n14820, n14821,
         n14822, n14823, n14824, n14825, n14826, n14827, n14828, n14829,
         n14830, n14831, n14832, n14833, n14834, n14835, n14836, n14837,
         n14838, n14839, n14840, n14841, n14842, n14843, n14844, n14845,
         n14846, n14847, n14848, n14849, n14850, n14851, n14852, n14853,
         n14854, n14855, n14856, n14857, n14858, n14859, n14860, n14861,
         n14862, n14863, n14864, n14865, n14866, n14867, n14868, n14869,
         n14870, n14871, n14872, n14873, n14874, n14875, n14876, n14877,
         n14878, n14879, n14880, n14881, n14882, n14883, n14884, n14885,
         n14886, n14887, n14888, n14889, n14890, n14891, n14892, n14893,
         n14894, n14895, n14896, n14897, n14898, n14899, n14900, n14901,
         n14902, n14903, n14904, n14905, n14906, n14907, n14908, n14909,
         n14910, n14911, n14912, n14913, n14914, n14915, n14916, n14917,
         n14918, n14919, n14920, n14921, n14922, n14923, n14924, n14925,
         n14926, n14927, n14928, n14929, n14930, n14931, n14932, n14933,
         n14934, n14935, n14936, n14937, n14938, n14939, n14940, n14941,
         n14942, n14943, n14944, n14945, n14946, n14947, n14948, n14949,
         n14950, n14951, n14952, n14953, n14954, n14955, n14956, n14957,
         n14958, n14959, n14960, n14961, n14962, n14963, n14964, n14965,
         n14966, n14967, n14968, n14969, n14970, n14971, n14972, n14973,
         n14974, n14975, n14976, n14977, n14978, n14979, n14980, n14981,
         n14982, n14983, n14984, n14985, n14986, n14987, n14988, n14989,
         n14990, n14991, n14992, n14993, n14994, n14995, n14996, n14997,
         n14998, n14999, n15000, n15001, n15002, n15003, n15004, n15005,
         n15006, n15007, n15008, n15009, n15010, n15011, n15012, n15013,
         n15014, n15015, n15016, n15017, n15018, n15019, n15020, n15021,
         n15022, n15023, n15024, n15025, n15026, n15027, n15028, n15029,
         n15030, n15031, n15032, n15033, n15034, n15035, n15036, n15037,
         n15038, n15039, n15040, n15041, n15042, n15043, n15044, n15045,
         n15046, n15047, n15048, n15049, n15050, n15051, n15052, n15053,
         n15054, n15055, n15056, n15057, n15058, n15059, n15060, n15061,
         n15062, n15063, n15064, n15065, n15066, n15067, n15068, n15069,
         n15070, n15071, n15072, n15073, n15074, n15075, n15076, n15077,
         n15078, n15079, n15080, n15081, n15082, n15083, n15084, n15085,
         n15086, n15087, n15088, n15089, n15090, n15091, n15092, n15093,
         n15094, n15095, n15096, n15097, n15098, n15099, n15100, n15101,
         n15102, n15103, n15104, n15105, n15106, n15107, n15108, n15109,
         n15110, n15111, n15112, n15113, n15114, n15115, n15116, n15117,
         n15118, n15119, n15120, n15121, n15122, n15123, n15124, n15125,
         n15126, n15127, n15128, n15129, n15130, n15131, n15132, n15133,
         n15134, n15135, n15136, n15137, n15138, n15139, n15140, n15141,
         n15142, n15143, n15144, n15145, n15146, n15147, n15148, n15149,
         n15150, n15151, n15152, n15153, n15154, n15155, n15156, n15157,
         n15158, n15159, n15160, n15161, n15162, n15163, n15164, n15165,
         n15166, n15167, n15168, n15169, n15170, n15171, n15172, n15173,
         n15174, n15175, n15176, n15177, n15178, n15179, n15180, n15181,
         n15182, n15183, n15184, n15185, n15186, n15187, n15188, n15189,
         n15190, n15191, n15192, n15193, n15194, n15195, n15196, n15197,
         n15198, n15199, n15200, n15201, n15202, n15203, n15204, n15205,
         n15206, n15207, n15208, n15209, n15210, n15211, n15212, n15213,
         n15214, n15215, n15216, n15217, n15218, n15219, n15220, n15221,
         n15222, n15223, n15224, n15225, n15226, n15227, n15228, n15229,
         n15230, n15231, n15232, n15233, n15234, n15235, n15236, n15237,
         n15238, n15239, n15240, n15241, n15242, n15243, n15244, n15245,
         n15246, n15247, n15248, n15249, n15250, n15251, n15252, n15253,
         n15254, n15255, n15256, n15257, n15258, n15259, n15260, n15261,
         n15262, n15263, n15264, n15265, n15266, n15267, n15268, n15269,
         n15270, n15271, n15272, n15273, n15274, n15275, n15276, n15277,
         n15278, n15279, n15280, n15281, n15282, n15283, n15284, n15285,
         n15286, n15287, n15288, n15289, n15290, n15291, n15292, n15293,
         n15294, n15295, n15296, n15297, n15298, n15299, n15300, n15301,
         n15302, n15303, n15304, n15305, n15306, n15307, n15308, n15309,
         n15310, n15311, n15312, n15313, n15314, n15315, n15316, n15317,
         n15318, n15319, n15320, n15321, n15322, n15323, n15324, n15325,
         n15326, n15327, n15328, n15329, n15330, n15331, n15332, n15333,
         n15334, n15335, n15336, n15337, n15338, n15339, n15340, n15341,
         n15342, n15343, n15344, n15345, n15346, n15347, n15348, n15349,
         n15350, n15351, n15352, n15353, n15354, n15355, n15356, n15357,
         n15358, n15359, n15360, n15361, n15362, n15363, n15364, n15365,
         n15366, n15367, n15368, n15369, n15370, n15371, n15372, n15373,
         n15374, n15375, n15376, n15377, n15378, n15379, n15380, n15381,
         n15382, n15383, n15384, n15385, n15386, n15387, n15388, n15389,
         n15390, n15391, n15392, n15393, n15394, n15395, n15396, n15397,
         n15398, n15399, n15400, n15401, n15402, n15403, n15404, n15405,
         n15406, n15407, n15408, n15409, n15410, n15411, n15412, n15413,
         n15414, n15415, n15416, n15417, n15418, n15419, n15420, n15421,
         n15422, n15423, n15424, n15425, n15426, n15427, n15428, n15429,
         n15430, n15431, n15432, n15433, n15434, n15435, n15436, n15437,
         n15438, n15439, n15440, n15441, n15442, n15443, n15444, n15445,
         n15446, n15447, n15448, n15449, n15450, n15451, n15452, n15453,
         n15454, n15455, n15456, n15457, n15458, n15459, n15460, n15461,
         n15462, n15463, n15464, n15465, n15466, n15467, n15468, n15469,
         n15470, n15471, n15472, n15473, n15474, n15475, n15476, n15477,
         n15478, n15479, n15480, n15481, n15482, n15483, n15484, n15485,
         n15486, n15487, n15488, n15489, n15490, n15491, n15492, n15493,
         n15494, n15495, n15496, n15497, n15498, n15499, n15500, n15501,
         n15502, n15503, n15504, n15505, n15506, n15507, n15508, n15509,
         n15510, n15511, n15512, n15513, n15514, n15515, n15516, n15517,
         n15518, n15519, n15520, n15521, n15522, n15523, n15524, n15525,
         n15526, n15527, n15528, n15529, n15530, n15531, n15532, n15533,
         n15534, n15535, n15536, n15537, n15538, n15539, n15540, n15541,
         n15542, n15543, n15544, n15545, n15546, n15547, n15548, n15549,
         n15550, n15551, n15552, n15553, n15554, n15555, n15556, n15557,
         n15558, n15559, n15560, n15561, n15562, n15563, n15564, n15565,
         n15566, n15567, n15568, n15569, n15570, n15571, n15572, n15573,
         n15574, n15575, n15576, n15577, n15578, n15579, n15580, n15581,
         n15582, n15583, n15584, n15585, n15586, n15587, n15588, n15589,
         n15590, n15591, n15592, n15593, n15594, n15595, n15596, n15597,
         n15598, n15599, n15600, n15601, n15602, n15603, n15604, n15605,
         n15606, n15607, n15608, n15609, n15610, n15611, n15612, n15613,
         n15614, n15615, n15616, n15617, n15618, n15619, n15620, n15621,
         n15622, n15623, n15624, n15625, n15626, n15627, n15628, n15629,
         n15630, n15631, n15632, n15633, n15634, n15635, n15636, n15637,
         n15638, n15639, n15640, n15641, n15642, n15643, n15644, n15645,
         n15646, n15647, n15648, n15649, n15650, n15651, n15652, n15653,
         n15654, n15655, n15656, n15657, n15658, n15659, n15660, n15661,
         n15662, n15663, n15664, n15665, n15666, n15667, n15668, n15669,
         n15670, n15671, n15672, n15673, n15674, n15675, n15676, n15677,
         n15678, n15679, n15680, n15681, n15682, n15683, n15684, n15685,
         n15686, n15687, n15688, n15689, n15690, n15691, n15692, n15693,
         n15694, n15695, n15696, n15697, n15698, n15699, n15700, n15701,
         n15702, n15703, n15704, n15705, n15706, n15707, n15708, n15709,
         n15710, n15711, n15712, n15713, n15714, n15715, n15716, n15717,
         n15718, n15719, n15720, n15721, n15722, n15723, n15724, n15725,
         n15726, n15727, n15728, n15729, n15730, n15731, n15732, n15733,
         n15734, n15735, n15736, n15737, n15738, n15739, n15740, n15741,
         n15742, n15743, n15744, n15745, n15746, n15747, n15748, n15749,
         n15750, n15751, n15752, n15753, n15754, n15755, n15756, n15757,
         n15758, n15759, n15760, n15761, n15762, n15763, n15764, n15765,
         n15766, n15767, n15768, n15769, n15770, n15771, n15772, n15773,
         n15774, n15775, n15776, n15777, n15778, n15779, n15780, n15781,
         n15782, n15783, n15784, n15785, n15786, n15787, n15788, n15789,
         n15790, n15791, n15792, n15793, n15794, n15795, n15796, n15797,
         n15798, n15799, n15800, n15801, n15802, n15803, n15804, n15805,
         n15806, n15807, n15808, n15809, n15810, n15811, n15812, n15813,
         n15814, n15815, n15816, n15817, n15818, n15819, n15820, n15821,
         n15822, n15823, n15824, n15825, n15826, n15827, n15828, n15829,
         n15830, n15831, n15832, n15833, n15834, n15835, n15836, n15837,
         n15838, n15839, n15840, n15841, n15842, n15843, n15844, n15845,
         n15846, n15847, n15848, n15849, n15850, n15851, n15852, n15853,
         n15854, n15855, n15856, n15857, n15858, n15859, n15860, n15861,
         n15862, n15863, n15864, n15865, n15866, n15867, n15868, n15869,
         n15870, n15871, n15872, n15873, n15874, n15875, n15876, n15877,
         n15878, n15879, n15880, n15881, n15882, n15883, n15884, n15885,
         n15886, n15887, n15888, n15889, n15890, n15891, n15892, n15893,
         n15894, n15895, n15896, n15897, n15898, n15899, n15900, n15901,
         n15902, n15903, n15904, n15905, n15906, n15907, n15908, n15909,
         n15910, n15911, n15912, n15913, n15914, n15915, n15916, n15917,
         n15918, n15919, n15920, n15921, n15922, n15923, n15924, n15925,
         n15926, n15927, n15928, n15929, n15930, n15931, n15932, n15933,
         n15934, n15935, n15936, n15937, n15938, n15939, n15940, n15941,
         n15942, n15943, n15944, n15945, n15946, n15947, n15948, n15949,
         n15950, n15951, n15952, n15953, n15954, n15955, n15956, n15957,
         n15958, n15959, n15960, n15961, n15962, n15963, n15964, n15965,
         n15966, n15967, n15968, n15969, n15970, n15971, n15972, n15973,
         n15974, n15975, n15976, n15977, n15978, n15979, n15980, n15981,
         n15982, n15983, n15984, n15985, n15986, n15987, n15988, n15989,
         n15990, n15991, n15992, n15993, n15994, n15995, n15996, n15997,
         n15998, n15999, n16000, n16001, n16002, n16003, n16004, n16005,
         n16006, n16007, n16008, n16009, n16010, n16011, n16012, n16013,
         n16014, n16015, n16016, n16017, n16018, n16019, n16020, n16021,
         n16022, n16023, n16024, n16025, n16026, n16027, n16028, n16029,
         n16030, n16031, n16032, n16033, n16034, n16035, n16036, n16037,
         n16038, n16039, n16040, n16041, n16042, n16043, n16044, n16045,
         n16046, n16047, n16048, n16049, n16050, n16051, n16052, n16053,
         n16054, n16055, n16056, n16057, n16058, n16059, n16060, n16061,
         n16062, n16063, n16064, n16065, n16066, n16067, n16068, n16069,
         n16070, n16071, n16072, n16073, n16074, n16075, n16076, n16077,
         n16078, n16079, n16080, n16081, n16082, n16083, n16084, n16085,
         n16086, n16087, n16088, n16089, n16090, n16091, n16092, n16093,
         n16094, n16095, n16096, n16097, n16098, n16099, n16100, n16101,
         n16102, n16103, n16104, n16105, n16106, n16107, n16108, n16109,
         n16110, n16111, n16112, n16113, n16114, n16115, n16116, n16117,
         n16118, n16119, n16120, n16121, n16122, n16123, n16124, n16125,
         n16126, n16127, n16128, n16129, n16130, n16131, n16132, n16133,
         n16134, n16135, n16136, n16137, n16138, n16139, n16140, n16141,
         n16142, n16143, n16144, n16145, n16146, n16147, n16148, n16149,
         n16150, n16151, n16152, n16153, n16154, n16155, n16156, n16157,
         n16158, n16159, n16160, n16161, n16162, n16163, n16164, n16165,
         n16166, n16167, n16168, n16169, n16170, n16171, n16172, n16173,
         n16174, n16175, n16176, n16177, n16178, n16179, n16180, n16181,
         n16182, n16183, n16184, n16185, n16186, n16187, n16188, n16189,
         n16190, n16191, n16192, n16193, n16194, n16195, n16196, n16197,
         n16198, n16199, n16200, n16201, n16202, n16203, n16204, n16205,
         n16206, n16207, n16208, n16209, n16210, n16211, n16212, n16213,
         n16214, n16215, n16216, n16217, n16218, n16219, n16220, n16221,
         n16222, n16223, n16224, n16225, n16226, n16227, n16228, n16229,
         n16230, n16231, n16232, n16233, n16234, n16235, n16236, n16237,
         n16238, n16239, n16240, n16241, n16242, n16243, n16244, n16245,
         n16246, n16247, n16248, n16249, n16250, n16251, n16252, n16253,
         n16254, n16255, n16256, n16257, n16258, n16259, n16260, n16261,
         n16262, n16263, n16264, n16265, n16266, n16267, n16268, n16269,
         n16270, n16271, n16272, n16273, n16274, n16275, n16276, n16277,
         n16278, n16279, n16280, n16281, n16282, n16283, n16284, n16285,
         n16286, n16287, n16288, n16289, n16290, n16291, n16292, n16293,
         n16294, n16295, n16296, n16297, n16298, n16299, n16300, n16301,
         n16302, n16303, n16304, n16305, n16306, n16307, n16308, n16309,
         n16310, n16311, n16312, n16313, n16314, n16315, n16316, n16317,
         n16318, n16319, n16320, n16321, n16322, n16323, n16324, n16325,
         n16326, n16327, n16328, n16329, n16330, n16331, n16332, n16333,
         n16334, n16335, n16336, n16337, n16338, n16339, n16340, n16341,
         n16342, n16343, n16344, n16345, n16346, n16347, n16348, n16349,
         n16350, n16351, n16352, n16353, n16354, n16355, n16356, n16357,
         n16358, n16359, n16360, n16361, n16362, n16363, n16364, n16365,
         n16366, n16367, n16368, n16369, n16370, n16371, n16372, n16373,
         n16374, n16375, n16376, n16377, n16378, n16379, n16380, n16381,
         n16382, n16383, n16384, n16385, n16386, n16387, n16388, n16389,
         n16390, n16391, n16392, n16393, n16394, n16395, n16396, n16397,
         n16398, n16399, n16400, n16401, n16402, n16403, n16404, n16405,
         n16406, n16407, n16408, n16409, n16410, n16411, n16412, n16413,
         n16414, n16415, n16416, n16417, n16418, n16419, n16420, n16421,
         n16422, n16423, n16424, n16425, n16426, n16427, n16428, n16429,
         n16430, n16431, n16432, n16433, n16434, n16435, n16436, n16437,
         n16438, n16439, n16440, n16441, n16442, n16443, n16444, n16445,
         n16446, n16447, n16448, n16449, n16450, n16451, n16452, n16453,
         n16454, n16455, n16456, n16457, n16458, n16459, n16460, n16461,
         n16462, n16463, n16464, n16465, n16466, n16467, n16468, n16469,
         n16470, n16471, n16472, n16473, n16474, n16475, n16476, n16477,
         n16478, n16479, n16480, n16481, n16482, n16483, n16484, n16485,
         n16486, n16487, n16488, n16489, n16490, n16491, n16492, n16493,
         n16494, n16495, n16496, n16497, n16498, n16499, n16500, n16501,
         n16502, n16503, n16504, n16505, n16506, n16507, n16508, n16509,
         n16510, n16511, n16512, n16513, n16514, n16515, n16516, n16517,
         n16518, n16519, n16520, n16521, n16522, n16523, n16524, n16525,
         n16526, n16527, n16528, n16529, n16530, n16531, n16532, n16533,
         n16534, n16535, n16536, n16537, n16538, n16539, n16540, n16541,
         n16542, n16543, n16544, n16545, n16546, n16547, n16548, n16549,
         n16550, n16551, n16552, n16553, n16554, n16555, n16556, n16557,
         n16558, n16559, n16560, n16561, n16562, n16563, n16564, n16565,
         n16566, n16567, n16568, n16569, n16570, n16571, n16572, n16573,
         n16574, n16575, n16576, n16577, n16578, n16579, n16580, n16581,
         n16582, n16583, n16584, n16585, n16586, n16587, n16588, n16589,
         n16590, n16591, n16592, n16593, n16594, n16595, n16596, n16597,
         n16598, n16599, n16600, n16601, n16602, n16603, n16604, n16605,
         n16606, n16607, n16608, n16609, n16610, n16611, n16612, n16613,
         n16614, n16615, n16616, n16617, n16618, n16619, n16620, n16621,
         n16622, n16623, n16624, n16625, n16626, n16627, n16628, n16629,
         n16630, n16631, n16632, n16633, n16634, n16635, n16636, n16637,
         n16638, n16639, n16640, n16641, n16642, n16643, n16644, n16645,
         n16646, n16647, n16648, n16649, n16650, n16651, n16652, n16653,
         n16654, n16655, n16656, n16657, n16658, n16659, n16660, n16661,
         n16662, n16663, n16664, n16665, n16666, n16667, n16668, n16669,
         n16670, n16671, n16672, n16673, n16674, n16675, n16676, n16677,
         n16678, n16679, n16680, n16681, n16682, n16683, n16684, n16685,
         n16686, n16687, n16688, n16689, n16690, n16691, n16692, n16693,
         n16694, n16695, n16696, n16697, n16698, n16699, n16700, n16701,
         n16702, n16703, n16704, n16705, n16706, n16707, n16708, n16709,
         n16710, n16711, n16712, n16713, n16714, n16715, n16716, n16717,
         n16718, n16719, n16720, n16721, n16722, n16723, n16724, n16725,
         n16726, n16727, n16728, n16729, n16730, n16731, n16732, n16733,
         n16734, n16735, n16736, n16737, n16738, n16739, n16740, n16741,
         n16742, n16743, n16744, n16745, n16746, n16747, n16748, n16749,
         n16750, n16751, n16752, n16753, n16754, n16755, n16756, n16757,
         n16758, n16759, n16760, n16761, n16762, n16763, n16764, n16765,
         n16766, n16767, n16768, n16769, n16770, n16771, n16772, n16773,
         n16774, n16775, n16776, n16777, n16778, n16779, n16780, n16781,
         n16782, n16783, n16784, n16785, n16786, n16787, n16788, n16789,
         n16790, n16791, n16792, n16793, n16794, n16795, n16796, n16797,
         n16798, n16799, n16800, n16801, n16802, n16803, n16804, n16805,
         n16806, n16807, n16808, n16809, n16810, n16811, n16812, n16813,
         n16814, n16815, n16816, n16817, n16818, n16819, n16820, n16821,
         n16822, n16823, n16824, n16825, n16826, n16827, n16828, n16829,
         n16830, n16831, n16832, n16833, n16834, n16835, n16836, n16837,
         n16838, n16839, n16840, n16841, n16842, n16843, n16844, n16845,
         n16846, n16847, n16848, n16849, n16850, n16851, n16852, n16853,
         n16854, n16855, n16856, n16857, n16858, n16859, n16860, n16861,
         n16862, n16863, n16864, n16865, n16866, n16867, n16868, n16869,
         n16870, n16871, n16872, n16873, n16874, n16875, n16876, n16877,
         n16878, n16879, n16880, n16881, n16882, n16883, n16884, n16885,
         n16886, n16887, n16888, n16889, n16890, n16891, n16892, n16893,
         n16894, n16895, n16896, n16897, n16898, n16899, n16900, n16901,
         n16902, n16903, n16904, n16905, n16906, n16907, n16908, n16909,
         n16910, n16911, n16912, n16913, n16914, n16915, n16916, n16917,
         n16918, n16919, n16920, n16921, n16922, n16923, n16924, n16925,
         n16926, n16927, n16928, n16929, n16930, n16931, n16932, n16933,
         n16934, n16935, n16936, n16937, n16938, n16939, n16940, n16941,
         n16942, n16943, n16944, n16945, n16946, n16947, n16948, n16949,
         n16950, n16951, n16952, n16953, n16954, n16955, n16956, n16957,
         n16958, n16959, n16960, n16961, n16962, n16963, n16964, n16965,
         n16966, n16967, n16968, n16969, n16970, n16971, n16972, n16973,
         n16974, n16975, n16976, n16977, n16978, n16979, n16980, n16981,
         n16982, n16983, n16984, n16985, n16986, n16987, n16988, n16989,
         n16990, n16991, n16992, n16993, n16994, n16995, n16996, n16997,
         n16998, n16999, n17000, n17001, n17002, n17003, n17004, n17005,
         n17006, n17007, n17008, n17009, n17010, n17011, n17012, n17013,
         n17014, n17015, n17016, n17017, n17018, n17019, n17020, n17021,
         n17022, n17023, n17024, n17025, n17026, n17027, n17028, n17029,
         n17030, n17031, n17032, n17033, n17034, n17035, n17036, n17037,
         n17038, n17039, n17040, n17041, n17042, n17043, n17044, n17045,
         n17046, n17047, n17048, n17049, n17050, n17051, n17052, n17053,
         n17054, n17055, n17056, n17057, n17058, n17059, n17060, n17061,
         n17062, n17063, n17064, n17065, n17066, n17067, n17068, n17069,
         n17070, n17071, n17072, n17073, n17074, n17075, n17076, n17077,
         n17078, n17079, n17080, n17081, n17082, n17083, n17084, n17085,
         n17086, n17087, n17088, n17089, n17090, n17091, n17092, n17093,
         n17094, n17095, n17096, n17097, n17098, n17099, n17100, n17101,
         n17102, n17103, n17104, n17105, n17106, n17107, n17108, n17109,
         n17110, n17111, n17112, n17113, n17114, n17115, n17116, n17117,
         n17118, n17119, n17120, n17121, n17122, n17123, n17124, n17125,
         n17126, n17127, n17128, n17129, n17130, n17131, n17132, n17133,
         n17134, n17135, n17136, n17137, n17138, n17139, n17140, n17141,
         n17142, n17143, n17144, n17145, n17146, n17147, n17148, n17149,
         n17150, n17151, n17152, n17153, n17154, n17155, n17156, n17157,
         n17158, n17159, n17160, n17161, n17162, n17163, n17164, n17165,
         n17166, n17167, n17168, n17169, n17170, n17171, n17172, n17173,
         n17174, n17175, n17176, n17177, n17178, n17179, n17180, n17181,
         n17182, n17183, n17184, n17185, n17186, n17187, n17188, n17189,
         n17190, n17191, n17192, n17193, n17194, n17195, n17196, n17197,
         n17198, n17199, n17200, n17201, n17202, n17203, n17204, n17205,
         n17206, n17207, n17208, n17209, n17210, n17211, n17212, n17213,
         n17214, n17215, n17216, n17217, n17218, n17219, n17220, n17221,
         n17222, n17223, n17224, n17225, n17226, n17227, n17228, n17229,
         n17230, n17231, n17232, n17233, n17234, n17235, n17236, n17237,
         n17238, n17239, n17240, n17241, n17242, n17243, n17244, n17245,
         n17246, n17247, n17248, n17249, n17250, n17251, n17252, n17253,
         n17254, n17255, n17256, n17257, n17258, n17259, n17260, n17261,
         n17262, n17263, n17264, n17265, n17266, n17267, n17268, n17269,
         n17270, n17271, n17272, n17273, n17274, n17275, n17276, n17277,
         n17278, n17279, n17280, n17281, n17282, n17283, n17284, n17285,
         n17286, n17287, n17288, n17289, n17290, n17291, n17292, n17293,
         n17294, n17295, n17296, n17297, n17298, n17299, n17300, n17301,
         n17302, n17303, n17304, n17305, n17306, n17307, n17308, n17309,
         n17310, n17311, n17312, n17313, n17314, n17315, n17316, n17317,
         n17318, n17319, n17320, n17321, n17322, n17323, n17324, n17325,
         n17326, n17327, n17328, n17329, n17330, n17331, n17332, n17333,
         n17334, n17335, n17336, n17337, n17338, n17339, n17340, n17341,
         n17342, n17343, n17344, n17345, n17346, n17347, n17348, n17349,
         n17350, n17351, n17352, n17353, n17354, n17355, n17356, n17357,
         n17358, n17359, n17360, n17361, n17362, n17363, n17364, n17365,
         n17366, n17367, n17368, n17369, n17370, n17371, n17372, n17373,
         n17374, n17375, n17376, n17377, n17378, n17379, n17380, n17381,
         n17382, n17383, n17384, n17385, n17386, n17387, n17388, n17389,
         n17390, n17391, n17392, n17393, n17394, n17395, n17396, n17397,
         n17398, n17399, n17400, n17401, n17402, n17403, n17404, n17405,
         n17406, n17407, n17408, n17409, n17410, n17411, n17412, n17413,
         n17414, n17415, n17416, n17417, n17418, n17419, n17420, n17421,
         n17422, n17423, n17424, n17425, n17426, n17427, n17428, n17429,
         n17430, n17431, n17432, n17433, n17434, n17435, n17436, n17437,
         n17438, n17439, n17440, n17441, n17442, n17443, n17444, n17445,
         n17446, n17447, n17448, n17449, n17450, n17451, n17452, n17453,
         n17454, n17455, n17456, n17457, n17458, n17459, n17460, n17461,
         n17462, n17463, n17464, n17465, n17466, n17467, n17468, n17469,
         n17470, n17471, n17472, n17473, n17474, n17475, n17476, n17477,
         n17478, n17479, n17480, n17481, n17482, n17483, n17484, n17485,
         n17486, n17487, n17488, n17489, n17490, n17491, n17492, n17493,
         n17494, n17495, n17496, n17497, n17498, n17499, n17500, n17501,
         n17502, n17503, n17504, n17505, n17506, n17507, n17508, n17509,
         n17510, n17511, n17512, n17513, n17514, n17515, n17516, n17517,
         n17518, n17519, n17520, n17521, n17522, n17523, n17524, n17525,
         n17526, n17527, n17528, n17529, n17530, n17531, n17532, n17533,
         n17534, n17535, n17536, n17537, n17538, n17539, n17540, n17541,
         n17542, n17543, n17544, n17545, n17546, n17547, n17548, n17549,
         n17550, n17551, n17552, n17553, n17554, n17555, n17556, n17557,
         n17558, n17559, n17560, n17561, n17562, n17563, n17564, n17565,
         n17566, n17567, n17568, n17569, n17570, n17571, n17572, n17573,
         n17574, n17575, n17576, n17577, n17578, n17579, n17580, n17581,
         n17582, n17583, n17584, n17585, n17586, n17587, n17588, n17589,
         n17590, n17591, n17592, n17593, n17594, n17595, n17596, n17597,
         n17598, n17599, n17600, n17601, n17602, n17603, n17604, n17605,
         n17606, n17607, n17608, n17609, n17610, n17611, n17612, n17613,
         n17614, n17615, n17616, n17617, n17618, n17619, n17620, n17621,
         n17622, n17623, n17624, n17625, n17626, n17627, n17628, n17629,
         n17630, n17631, n17632, n17633, n17634, n17635, n17636, n17637,
         n17638, n17639, n17640, n17641, n17642, n17643, n17644, n17645,
         n17646, n17647, n17648, n17649, n17650, n17651, n17652, n17653,
         n17654, n17655, n17656, n17657, n17658, n17659, n17660, n17661,
         n17662, n17663, n17664, n17665, n17666, n17667, n17668, n17669,
         n17670, n17671, n17672, n17673, n17674, n17675, n17676, n17677,
         n17678, n17679, n17680, n17681, n17682, n17683, n17684, n17685,
         n17686, n17687, n17688, n17689, n17690, n17691, n17692, n17693,
         n17694, n17695, n17696, n17697, n17698, n17699, n17700, n17701,
         n17702, n17703, n17704, n17705, n17706, n17707, n17708, n17709,
         n17710, n17711, n17712, n17713, n17714, n17715, n17716, n17717,
         n17718, n17719, n17720, n17721, n17722, n17723, n17724, n17725,
         n17726, n17727, n17728, n17729, n17730, n17731, n17732, n17733,
         n17734, n17735, n17736, n17737, n17738, n17739, n17740, n17741,
         n17742, n17743, n17744, n17745, n17746, n17747, n17748, n17749,
         n17750, n17751, n17752, n17753, n17754, n17755, n17756, n17757,
         n17758, n17759, n17760, n17761, n17762, n17763, n17764, n17765,
         n17766, n17767, n17768, n17769, n17770, n17771, n17772, n17773,
         n17774, n17775, n17776, n17777, n17778, n17779, n17780, n17781,
         n17782, n17783, n17784, n17785, n17786, n17787, n17788, n17789,
         n17790, n17791, n17792, n17793, n17794, n17795, n17796, n17797,
         n17798, n17799, n17800, n17801, n17802, n17803, n17804, n17805,
         n17806, n17807, n17808, n17809, n17810, n17811, n17812, n17813,
         n17814, n17815, n17816, n17817, n17818, n17819, n17820, n17821,
         n17822, n17823, n17824, n17825, n17826, n17827, n17828, n17829,
         n17830, n17831, n17832, n17833, n17834, n17835, n17836, n17837,
         n17838, n17839, n17840, n17841, n17842, n17843, n17844, n17845,
         n17846, n17847, n17848, n17849, n17850, n17851, n17852, n17853,
         n17854, n17855, n17856, n17857, n17858, n17859, n17860, n17861,
         n17862, n17863, n17864, n17865, n17866, n17867, n17868, n17869,
         n17870, n17871, n17872, n17873, n17874, n17875, n17876, n17877,
         n17878, n17879, n17880, n17881, n17882, n17883, n17884, n17885,
         n17886, n17887, n17888, n17889, n17890, n17891, n17892, n17893,
         n17894, n17895, n17896, n17897, n17898, n17899, n17900, n17901,
         n17902, n17903, n17904, n17905, n17906, n17907, n17908, n17909,
         n17910, n17911, n17912, n17913, n17914, n17915, n17916, n17917,
         n17918, n17919, n17920, n17921, n17922, n17923, n17924, n17925,
         n17926, n17927, n17928, n17929, n17930, n17931, n17932, n17933,
         n17934, n17935, n17936, n17937, n17938, n17939, n17940, n17941,
         n17942, n17943, n17944, n17945, n17946, n17947, n17948, n17949,
         n17950, n17951, n17952, n17953, n17954, n17955, n17956, n17957,
         n17958, n17959, n17960, n17961, n17962, n17963, n17964, n17965,
         n17966, n17967, n17968, n17969, n17970, n17971, n17972, n17973,
         n17974, n17975, n17976, n17977, n17978, n17979, n17980, n17981,
         n17982, n17983, n17984, n17985, n17986, n17987, n17988, n17989,
         n17990, n17991, n17992, n17993, n17994, n17995, n17996, n17997,
         n17998, n17999, n18000, n18001, n18002, n18003, n18004, n18005,
         n18006, n18007, n18008, n18009, n18010, n18011, n18012, n18013,
         n18014, n18015, n18016, n18017, n18018, n18019, n18020, n18021,
         n18022, n18023, n18024, n18025, n18026, n18027, n18028, n18029,
         n18030, n18031, n18032, n18033, n18034, n18035, n18036, n18037,
         n18038, n18039, n18040, n18041, n18042, n18043, n18044, n18045,
         n18046, n18047, n18048, n18049, n18050, n18051, n18052, n18053,
         n18054, n18055, n18056, n18057, n18058, n18059, n18060, n18061,
         n18062, n18063, n18064, n18065, n18066, n18067, n18068, n18069,
         n18070, n18071, n18072, n18073, n18074, n18075, n18076, n18077,
         n18078, n18079, n18080, n18081, n18082, n18083, n18084, n18085,
         n18086, n18087, n18088, n18089, n18090, n18091, n18092, n18093,
         n18094, n18095, n18096, n18097, n18098, n18099, n18100, n18101,
         n18102, n18103, n18104, n18105, n18106, n18107, n18108, n18109,
         n18110, n18111, n18112, n18113, n18114, n18115, n18116, n18117,
         n18118, n18119, n18120, n18121, n18122, n18123, n18124, n18125,
         n18126, n18127, n18128, n18129, n18130, n18131, n18132, n18133,
         n18134, n18135, n18136, n18137, n18138, n18139, n18140, n18141,
         n18142, n18143, n18144, n18145, n18146, n18147, n18148, n18149,
         n18150, n18151, n18152, n18153, n18154, n18155, n18156, n18157,
         n18158, n18159, n18160, n18161, n18162, n18163, n18164, n18165,
         n18166, n18167, n18168, n18169, n18170, n18171, n18172, n18173,
         n18174, n18175, n18176, n18177, n18178, n18179, n18180, n18181,
         n18182, n18183, n18184, n18185, n18186, n18187, n18188, n18189,
         n18190, n18191, n18192, n18193, n18194, n18195, n18196, n18197,
         n18198, n18199, n18200, n18201, n18202, n18203, n18204, n18205,
         n18206, n18207, n18208, n18209, n18210, n18211, n18212, n18213,
         n18214, n18215, n18216, n18217, n18218, n18219, n18220, n18221,
         n18222, n18223, n18224, n18225, n18226, n18227, n18228, n18229,
         n18230, n18231, n18232, n18233, n18234, n18235, n18236, n18237,
         n18238, n18239, n18240, n18241, n18242, n18243, n18244, n18245,
         n18246, n18247, n18248, n18249, n18250, n18251, n18252, n18253,
         n18254, n18255, n18256, n18257, n18258, n18259, n18260, n18261,
         n18262, n18263, n18264, n18265, n18266, n18267, n18268, n18269,
         n18270, n18271, n18272, n18273, n18274, n18275, n18276, n18277,
         n18278, n18279, n18280, n18281, n18282, n18283, n18284, n18285,
         n18286, n18287, n18288, n18289, n18290, n18291, n18292, n18293,
         n18294, n18295, n18296, n18297, n18298, n18299, n18300, n18301,
         n18302, n18303, n18304, n18305, n18306, n18307, n18308, n18309,
         n18310, n18311, n18312, n18313, n18314, n18315, n18316, n18317,
         n18318, n18319, n18320, n18321, n18322, n18323, n18324, n18325,
         n18326, n18327, n18328, n18329, n18330, n18331, n18332, n18333,
         n18334, n18335, n18336, n18337, n18338, n18339, n18340, n18341,
         n18342, n18343, n18344, n18345, n18346, n18347, n18348, n18349,
         n18350, n18351, n18352, n18353, n18354, n18355, n18356, n18357,
         n18358, n18359, n18360, n18361, n18362, n18363, n18364, n18365,
         n18366, n18367, n18368, n18369, n18370, n18371, n18372, n18373,
         n18374, n18375, n18376, n18377, n18378, n18379, n18380, n18381,
         n18382, n18383, n18384, n18385, n18386, n18387, n18388, n18389,
         n18390, n18391, n18392, n18393, n18394, n18395, n18396, n18397,
         n18398, n18399, n18400, n18401, n18402, n18403, n18404, n18405,
         n18406, n18407, n18408, n18409, n18410, n18411, n18412, n18413,
         n18414, n18415, n18416, n18417, n18418, n18419, n18420, n18421,
         n18422, n18423, n18424, n18425, n18426, n18427, n18428, n18429,
         n18430, n18431, n18432, n18433, n18434, n18435, n18436, n18437,
         n18438, n18439, n18440, n18441, n18442, n18443, n18444, n18445,
         n18446, n18447, n18448, n18449, n18450, n18451, n18452, n18453,
         n18454, n18455, n18456, n18457, n18458, n18459, n18460, n18461,
         n18462, n18463, n18464, n18465, n18466, n18467, n18468, n18469,
         n18470, n18471, n18472, n18473, n18474, n18475, n18476, n18477,
         n18478, n18479, n18480, n18481, n18482, n18483, n18484, n18485,
         n18486, n18487, n18488, n18489, n18490, n18491, n18492, n18493,
         n18494, n18495, n18496, n18497, n18498, n18499, n18500, n18501,
         n18502, n18503, n18504, n18505, n18506, n18507, n18508, n18509,
         n18510, n18511, n18512, n18513, n18514, n18515, n18516, n18517,
         n18518, n18519, n18520, n18521, n18522, n18523, n18524, n18525,
         n18526, n18527, n18528, n18529, n18530, n18531, n18532, n18533,
         n18534, n18535, n18536, n18537, n18538, n18539, n18540, n18541,
         n18542, n18543, n18544, n18545, n18546, n18547, n18548, n18549,
         n18550, n18551, n18552, n18553, n18554, n18555, n18556, n18557,
         n18558, n18559, n18560, n18561, n18562, n18563, n18564, n18565,
         n18566, n18567, n18568, n18569, n18570, n18571, n18572, n18573,
         n18574, n18575, n18576, n18577, n18578, n18579, n18580, n18581,
         n18582, n18583, n18584, n18585, n18586, n18587, n18588, n18589,
         n18590, n18591, n18592, n18593, n18594, n18595, n18596, n18597,
         n18598, n18599, n18600, n18601, n18602, n18603, n18604, n18605,
         n18606, n18607, n18608, n18609, n18610, n18611, n18612, n18613,
         n18614, n18615, n18616, n18617, n18618, n18619, n18620, n18621,
         n18622, n18623, n18624, n18625, n18626, n18627, n18628, n18629,
         n18630, n18631, n18632, n18633, n18634, n18635, n18636, n18637,
         n18638, n18639, n18640, n18641, n18642, n18643, n18644, n18645,
         n18646, n18647, n18648, n18649, n18650, n18651, n18652, n18653,
         n18654, n18655, n18656, n18657, n18658, n18659, n18660, n18661,
         n18662, n18663, n18664, n18665, n18666, n18667, n18668, n18669,
         n18670, n18671, n18672, n18673, n18674, n18675, n18676, n18677,
         n18678, n18679, n18680, n18681, n18682, n18683, n18684, n18685,
         n18686, n18687, n18688, n18689, n18690, n18691, n18692, n18693,
         n18694, n18695, n18696, n18697, n18698, n18699, n18700, n18701,
         n18702, n18703, n18704, n18705, n18706, n18707, n18708, n18709,
         n18710, n18711, n18712, n18713, n18714, n18715, n18716, n18717,
         n18718, n18719, n18720, n18721, n18722, n18723, n18724, n18725,
         n18726, n18727, n18728, n18729, n18730, n18731, n18732, n18733,
         n18734, n18735, n18736, n18737, n18738, n18739, n18740, n18741,
         n18742, n18743, n18744, n18745, n18746, n18747, n18748, n18749,
         n18750, n18751, n18752, n18753, n18754, n18755, n18756, n18757,
         n18758, n18759, n18760, n18761, n18762, n18763, n18764, n18765,
         n18766, n18767, n18768, n18769, n18770, n18771, n18772, n18773,
         n18774, n18775, n18776, n18777, n18778, n18779, n18780, n18781,
         n18782, n18783, n18784, n18785, n18786, n18787, n18788, n18789,
         n18790, n18791, n18792, n18793, n18794, n18795, n18796, n18797,
         n18798, n18799, n18800, n18801, n18802, n18803, n18804, n18805,
         n18806, n18807, n18808, n18809, n18810, n18811, n18812, n18813,
         n18814, n18815, n18816, n18817, n18818, n18819, n18820, n18821,
         n18822, n18823, n18824, n18825, n18826, n18827, n18828, n18829,
         n18830, n18831, n18832, n18833, n18834, n18835, n18836, n18837,
         n18838, n18839, n18840, n18841, n18842, n18843, n18844, n18845,
         n18846, n18847, n18848, n18849, n18850, n18851, n18852, n18853,
         n18854, n18855, n18856, n18857, n18858, n18859, n18860, n18861,
         n18862, n18863, n18864, n18865, n18866, n18867, n18868, n18869,
         n18870, n18871, n18872, n18873, n18874, n18875, n18876, n18877,
         n18878, n18879, n18880, n18881, n18882, n18883, n18884, n18885,
         n18886, n18887, n18888, n18889, n18890, n18891, n18892, n18893,
         n18894, n18895, n18896, n18897, n18898, n18899, n18900, n18901,
         n18902, n18903, n18904, n18905, n18906, n18907, n18908, n18909,
         n18910, n18911, n18912, n18913, n18914, n18915, n18916, n18917,
         n18918, n18919, n18920, n18921, n18922, n18923, n18924, n18925,
         n18926, n18927, n18928, n18929, n18930, n18931, n18932, n18933,
         n18934, n18935, n18936, n18937, n18938, n18939, n18940, n18941,
         n18942, n18943, n18944, n18945, n18946, n18947, n18948, n18949,
         n18950, n18951, n18952, n18953, n18954, n18955, n18956, n18957,
         n18958, n18959, n18960, n18961, n18962, n18963, n18964, n18965,
         n18966, n18967, n18968, n18969, n18970, n18971, n18972, n18973,
         n18974, n18975, n18976, n18977, n18978, n18979, n18980, n18981,
         n18982, n18983, n18984, n18985, n18986, n18987, n18988, n18989,
         n18990, n18991, n18992, n18993, n18994, n18995, n18996, n18997,
         n18998, n18999, n19000, n19001, n19002, n19003, n19004, n19005,
         n19006, n19007, n19008, n19009, n19010, n19011, n19012, n19013,
         n19014, n19015, n19016, n19017, n19018, n19019, n19020, n19021,
         n19022, n19023, n19024, n19025, n19026, n19027, n19028, n19029,
         n19030, n19031, n19032, n19033, n19034, n19035, n19036, n19037,
         n19038, n19039, n19040, n19041, n19042, n19043, n19044, n19045,
         n19046, n19047, n19048, n19049, n19050, n19051, n19052, n19053,
         n19054, n19055, n19056, n19057, n19058, n19059, n19060, n19061,
         n19062, n19063, n19064, n19065, n19066, n19067, n19068, n19069,
         n19070, n19071, n19072, n19073, n19074, n19075, n19076, n19077,
         n19078, n19079, n19080, n19081, n19082, n19083, n19084, n19085,
         n19086, n19087, n19088, n19089, n19090, n19091, n19092, n19093,
         n19094, n19095, n19096, n19097, n19098, n19099, n19100, n19101,
         n19102, n19103, n19104, n19105, n19106, n19107, n19108, n19109,
         n19110, n19111, n19112, n19113, n19114, n19115, n19116, n19117,
         n19118, n19119, n19120, n19121, n19122, n19123, n19124, n19125,
         n19126, n19127, n19128, n19129, n19130, n19131, n19132, n19133,
         n19134, n19135, n19136, n19137, n19138, n19139, n19140, n19141,
         n19142, n19143, n19144, n19145, n19146, n19147, n19148, n19149,
         n19150, n19151, n19152, n19153, n19154, n19155, n19156, n19157,
         n19158, n19159, n19160, n19161, n19162, n19163, n19164, n19165,
         n19166, n19167, n19168, n19169, n19170, n19171, n19172, n19173,
         n19174, n19175, n19176, n19177, n19178, n19179, n19180, n19181,
         n19182, n19183, n19184, n19185, n19186, n19187, n19188, n19189,
         n19190, n19191, n19192, n19193, n19194, n19195, n19196, n19197,
         n19198, n19199, n19200, n19201, n19202, n19203, n19204, n19205,
         n19206, n19207, n19208, n19209, n19210, n19211, n19212, n19213,
         n19214, n19215, n19216, n19217, n19218, n19219, n19220, n19221,
         n19222, n19223, n19224, n19225, n19226, n19227, n19228, n19229,
         n19230, n19231, n19232, n19233, n19234, n19235, n19236, n19237,
         n19238, n19239, n19240, n19241, n19242, n19243, n19244, n19245,
         n19246, n19247, n19248, n19249, n19250, n19251, n19252, n19253,
         n19254, n19255, n19256, n19257, n19258, n19259, n19260, n19261,
         n19262, n19263, n19264, n19265, n19266, n19267, n19268, n19269,
         n19270, n19271, n19272, n19273, n19274, n19275, n19276, n19277,
         n19278, n19279, n19280, n19281, n19282, n19283, n19284, n19285,
         n19286, n19287, n19288, n19289, n19290, n19291, n19292, n19293,
         n19294, n19295, n19296, n19297, n19298, n19299, n19300, n19301,
         n19302, n19303, n19304, n19305, n19306, n19307, n19308, n19309,
         n19310, n19311, n19312, n19313, n19314, n19315, n19316, n19317,
         n19318, n19319, n19320, n19321, n19322, n19323, n19324, n19325,
         n19326, n19327, n19328, n19329, n19330, n19331, n19332, n19333,
         n19334, n19335, n19336, n19337, n19338, n19339, n19340, n19341,
         n19342, n19343, n19344, n19345, n19346, n19347, n19348, n19349,
         n19350, n19351, n19352, n19353, n19354, n19355, n19356, n19357,
         n19358, n19359, n19360, n19361, n19362, n19363, n19364, n19365,
         n19366, n19367, n19368, n19369, n19370, n19371, n19372, n19373,
         n19374, n19375, n19376, n19377, n19378, n19379, n19380, n19381,
         n19382, n19383, n19384, n19385, n19386, n19387, n19388, n19389,
         n19390, n19391, n19392, n19393, n19394, n19395, n19396, n19397,
         n19398, n19399, n19400, n19401, n19402, n19403, n19404, n19405,
         n19406, n19407, n19408, n19409, n19410, n19411, n19412, n19413,
         n19414, n19415, n19416, n19417, n19418, n19419, n19420, n19421,
         n19422, n19423, n19424, n19425, n19426, n19427, n19428, n19429,
         n19430, n19431, n19432, n19433, n19434, n19435, n19436, n19437,
         n19438, n19439, n19440, n19441, n19442, n19443, n19444, n19445,
         n19446, n19447, n19448, n19449, n19450, n19451, n19452, n19453,
         n19454, n19455, n19456, n19457, n19458, n19459, n19460, n19461,
         n19462, n19463, n19464, n19465, n19466, n19467, n19468, n19469,
         n19470, n19471, n19472, n19473, n19474, n19475, n19476, n19477,
         n19478, n19479, n19480, n19481, n19482, n19483, n19484, n19485,
         n19486, n19487, n19488, n19489, n19490, n19491, n19492, n19493,
         n19494, n19495, n19496, n19497, n19498, n19499, n19500, n19501,
         n19502, n19503, n19504, n19505, n19506, n19507, n19508, n19509,
         n19510, n19511, n19512, n19513, n19514, n19515, n19516, n19517,
         n19518, n19519, n19520, n19521, n19522, n19523, n19524, n19525,
         n19526, n19527, n19528, n19529, n19530, n19531, n19532, n19533,
         n19534, n19535, n19536, n19537, n19538, n19539, n19540, n19541,
         n19542, n19543, n19544, n19545, n19546, n19547, n19548, n19549,
         n19550, n19551, n19552, n19553, n19554, n19555, n19556, n19557,
         n19558, n19559, n19560, n19561, n19562, n19563, n19564, n19565,
         n19566, n19567, n19568, n19569, n19570, n19571, n19572, n19573,
         n19574, n19575, n19576, n19577, n19578, n19579, n19580, n19581,
         n19582, n19583, n19584, n19585, n19586, n19587, n19588, n19589,
         n19590, n19591, n19592, n19593, n19594, n19595, n19596, n19597,
         n19598, n19599, n19600, n19601, n19602, n19603, n19604, n19605,
         n19606, n19607, n19608, n19609, n19610, n19611, n19612, n19613,
         n19614, n19615, n19616, n19617, n19618, n19619, n19620, n19621,
         n19622, n19623, n19624, n19625, n19626, n19627, n19628, n19629,
         n19630, n19631, n19632, n19633, n19634, n19635, n19636, n19637,
         n19638, n19639, n19640, n19641, n19642, n19643, n19644, n19645,
         n19646, n19647, n19648, n19649, n19650, n19651, n19652, n19653,
         n19654, n19655, n19656, n19657, n19658, n19659, n19660, n19661,
         n19662, n19663, n19664, n19665, n19666, n19667, n19668, n19669,
         n19670, n19671, n19672, n19673, n19674, n19675, n19676, n19677,
         n19678, n19679, n19680, n19681, n19682, n19683, n19684, n19685,
         n19686, n19687, n19688, n19689, n19690, n19691, n19692, n19693,
         n19694, n19695, n19696, n19697, n19698, n19699, n19700, n19701,
         n19702, n19703, n19704, n19705, n19706, n19707, n19708, n19709,
         n19710, n19711, n19712, n19713, n19714, n19715, n19716, n19717,
         n19718, n19719, n19720, n19721, n19722, n19723, n19724, n19725,
         n19726, n19727, n19728, n19729, n19730, n19731, n19732, n19733,
         n19734, n19735, n19736, n19737, n19738, n19739, n19740, n19741,
         n19742, n19743, n19744, n19745, n19746, n19747, n19748, n19749,
         n19750, n19751, n19752, n19753, n19754, n19755, n19756, n19757,
         n19758, n19759, n19760, n19761, n19762, n19763, n19764, n19765,
         n19766, n19767, n19768, n19769, n19770, n19771, n19772, n19773,
         n19774, n19775, n19776, n19777, n19778, n19779, n19780, n19781,
         n19782, n19783, n19784, n19785, n19786, n19787, n19788, n19789,
         n19790, n19791, n19792, n19793, n19794, n19795, n19796, n19797,
         n19798, n19799, n19800, n19801, n19802, n19803, n19804, n19805,
         n19806, n19807, n19808, n19809, n19810, n19811, n19812, n19813,
         n19814, n19815, n19816, n19817, n19818, n19819, n19820, n19821,
         n19822, n19823, n19824, n19825, n19826, n19827, n19828, n19829,
         n19830, n19831, n19832, n19833, n19834, n19835, n19836, n19837,
         n19838, n19839, n19840, n19841, n19842, n19843, n19844, n19845,
         n19846, n19847, n19848, n19849, n19850, n19851, n19852, n19853,
         n19854, n19855, n19856, n19857, n19858, n19859, n19860, n19861,
         n19862, n19863, n19864, n19865, n19866, n19867, n19868, n19869,
         n19870, n19871, n19872, n19873, n19874, n19875, n19876, n19877,
         n19878, n19879, n19880, n19881, n19882, n19883, n19884, n19885,
         n19886, n19887, n19888, n19889, n19890, n19891, n19892, n19893,
         n19894, n19895, n19896, n19897, n19898, n19899, n19900, n19901,
         n19902, n19903, n19904, n19905, n19906, n19907, n19908, n19909,
         n19910, n19911, n19912, n19913, n19914, n19915, n19916, n19917,
         n19918, n19919, n19920, n19921, n19922, n19923, n19924, n19925,
         n19926, n19927, n19928, n19929, n19930, n19931, n19932, n19933,
         n19934, n19935, n19936, n19937, n19938, n19939, n19940, n19941,
         n19942, n19943, n19944, n19945, n19946, n19947, n19948, n19949,
         n19950, n19951, n19952, n19953, n19954, n19955, n19956, n19957,
         n19958, n19959, n19960, n19961, n19962, n19963, n19964, n19965,
         n19966, n19967, n19968, n19969, n19970, n19971, n19972, n19973,
         n19974, n19975, n19976, n19977, n19978, n19979, n19980, n19981,
         n19982, n19983, n19984, n19985, n19986, n19987, n19988, n19989,
         n19990, n19991, n19992, n19993, n19994, n19995, n19996, n19997,
         n19998, n19999, n20000, n20001, n20002, n20003, n20004, n20005,
         n20006, n20007, n20008, n20009, n20010, n20011, n20012, n20013,
         n20014, n20015, n20016, n20017, n20018, n20019, n20020, n20021,
         n20022, n20023, n20024, n20025, n20026, n20027, n20028, n20029,
         n20030, n20031, n20032, n20033, n20034, n20035, n20036, n20037,
         n20038, n20039, n20040, n20041, n20042, n20043, n20044, n20045,
         n20046, n20047, n20048, n20049, n20050, n20051, n20052, n20053,
         n20054, n20055, n20056, n20057, n20058, n20059, n20060, n20061,
         n20062, n20063, n20064, n20065, n20066, n20067, n20068, n20069,
         n20070, n20071, n20072, n20073, n20074, n20075, n20076, n20077,
         n20078, n20079, n20080, n20081, n20082, n20083, n20084, n20085,
         n20086, n20087, n20088, n20089, n20090, n20091, n20092, n20093,
         n20094, n20095, n20096, n20097, n20098, n20099, n20100, n20101,
         n20102, n20103, n20104, n20105, n20106, n20107, n20108, n20109,
         n20110, n20111, n20112, n20113, n20114, n20115, n20116, n20117,
         n20118, n20119, n20120, n20121, n20122, n20123, n20124, n20125,
         n20126, n20127, n20128, n20129, n20130, n20131, n20132, n20133,
         n20134, n20135, n20136, n20137, n20138, n20139, n20140, n20141,
         n20142, n20143, n20144, n20145, n20146, n20147, n20148, n20149,
         n20150, n20151, n20152, n20153, n20154, n20155, n20156, n20157,
         n20158, n20159, n20160, n20161, n20162, n20163, n20164, n20165,
         n20166, n20167, n20168, n20169, n20170, n20171, n20172, n20173,
         n20174, n20175, n20176, n20177, n20178, n20179, n20180, n20181,
         n20182, n20183, n20184, n20185, n20186, n20187, n20188, n20189,
         n20190, n20191, n20192, n20193, n20194, n20195, n20196, n20197,
         n20198, n20199, n20200, n20201, n20202, n20203, n20204, n20205,
         n20206, n20207, n20208, n20209, n20210, n20211, n20212, n20213,
         n20214, n20215, n20216, n20217, n20218, n20219, n20220, n20221,
         n20222, n20223, n20224, n20225, n20226, n20227, n20228, n20229,
         n20230, n20231, n20232, n20233, n20234, n20235, n20236, n20237,
         n20238, n20239, n20240, n20241, n20242, n20243, n20244, n20245,
         n20246, n20247, n20248, n20249, n20250, n20251, n20252, n20253,
         n20254, n20255, n20256, n20257, n20258, n20259, n20260, n20261,
         n20262, n20263, n20264, n20265, n20266, n20267, n20268, n20269,
         n20270, n20271, n20272, n20273, n20274, n20275, n20276, n20277,
         n20278, n20279, n20280, n20281, n20282, n20283, n20284, n20285,
         n20286, n20287, n20288, n20289, n20290, n20291, n20292, n20293,
         n20294, n20295, n20296, n20297, n20298, n20299, n20300, n20301,
         n20302, n20303, n20304, n20305, n20306, n20307, n20308, n20309,
         n20310, n20311, n20312, n20313, n20314, n20315, n20316, n20317,
         n20318, n20319, n20320, n20321, n20322, n20323, n20324, n20325,
         n20326, n20327, n20328, n20329, n20330, n20331, n20332, n20333,
         n20334, n20335, n20336, n20337, n20338, n20339, n20340, n20341,
         n20342, n20343, n20344, n20345, n20346, n20347, n20348, n20349,
         n20350, n20351, n20352, n20353, n20354, n20355, n20356, n20357,
         n20358, n20359, n20360, n20361, n20362, n20363, n20364, n20365,
         n20366, n20367, n20368, n20369, n20370, n20371, n20372, n20373,
         n20374, n20375, n20376, n20377, n20378, n20379, n20380, n20381,
         n20382, n20383, n20384, n20385, n20386, n20387, n20388, n20389,
         n20390, n20391, n20392, n20393, n20394, n20395, n20396, n20397,
         n20398, n20399, n20400, n20401, n20402, n20403, n20404, n20405,
         n20406, n20407, n20408, n20409, n20410, n20411, n20412, n20413,
         n20414, n20415, n20416, n20417, n20418, n20419, n20420, n20421,
         n20422, n20423, n20424, n20425, n20426, n20427, n20428, n20429,
         n20430, n20431, n20432, n20433, n20434, n20435, n20436, n20437,
         n20438, n20439, n20440, n20441, n20442, n20443, n20444, n20445,
         n20446, n20447, n20448, n20449, n20450, n20451, n20452, n20453,
         n20454, n20455, n20456, n20457, n20458, n20459, n20460, n20461,
         n20462, n20463, n20464, n20465, n20466, n20467, n20468, n20469,
         n20470, n20471, n20472, n20473, n20474, n20475, n20476, n20477,
         n20478, n20479, n20480, n20481, n20482, n20483, n20484, n20485,
         n20486, n20487, n20488, n20489, n20490, n20491, n20492, n20493,
         n20494, n20495, n20496, n20497, n20498, n20499, n20500, n20501,
         n20502, n20503, n20504, n20505, n20506, n20507, n20508, n20509,
         n20510, n20511, n20512, n20513, n20514, n20515, n20516, n20517,
         n20518, n20519, n20520, n20521, n20522, n20523, n20524, n20525,
         n20526, n20527, n20528, n20529, n20530, n20531, n20532, n20533,
         n20534, n20535, n20536, n20537, n20538, n20539, n20540, n20541,
         n20542, n20543, n20544, n20545, n20546, n20547, n20548, n20549,
         n20550, n20551, n20552, n20553, n20554, n20555, n20556, n20557,
         n20558, n20559, n20560, n20561, n20562, n20563, n20564, n20565,
         n20566, n20567, n20568, n20569, n20570, n20571, n20572, n20573,
         n20574, n20575, n20576, n20577, n20578, n20579, n20580, n20581,
         n20582, n20583, n20584, n20585, n20586, n20587, n20588, n20589,
         n20590, n20591, n20592, n20593, n20594, n20595, n20596, n20597,
         n20598, n20599, n20600, n20601, n20602, n20603, n20604, n20605,
         n20606, n20607, n20608, n20609, n20610, n20611, n20612, n20613,
         n20614, n20615, n20616, n20617, n20618, n20619, n20620, n20621,
         n20622, n20623, n20624, n20625, n20626, n20627, n20628, n20629,
         n20630, n20631, n20632, n20633, n20634, n20635, n20636, n20637,
         n20638, n20639, n20640, n20641, n20642, n20643, n20644, n20645,
         n20646, n20647, n20648, n20649, n20650, n20651, n20652, n20653,
         n20654, n20655, n20656, n20657, n20658, n20659, n20660, n20661,
         n20662, n20663, n20664, n20665, n20666, n20667, n20668, n20669,
         n20670, n20671, n20672, n20673, n20674, n20675, n20676, n20677,
         n20678, n20679, n20680, n20681, n20682, n20683, n20684, n20685,
         n20686, n20687, n20688, n20689, n20690, n20691, n20692, n20693,
         n20694, n20695, n20696, n20697, n20698, n20699, n20700, n20701,
         n20702, n20703, n20704, n20705, n20706, n20707, n20708, n20709,
         n20710, n20711, n20712, n20713, n20714, n20715, n20716, n20717,
         n20718, n20719, n20720, n20721, n20722, n20723, n20724, n20725,
         n20726, n20727, n20728, n20729, n20730, n20731, n20732, n20733,
         n20734, n20735, n20736, n20737, n20738, n20739, n20740, n20741,
         n20742, n20743, n20744, n20745, n20746, n20747, n20748, n20749,
         n20750, n20751, n20752, n20753, n20754, n20755, n20756, n20757,
         n20758, n20759, n20760, n20761, n20762, n20763, n20764, n20765,
         n20766, n20767, n20768, n20769, n20770, n20771, n20772, n20773,
         n20774, n20775, n20776, n20777, n20778, n20779, n20780, n20781,
         n20782, n20783, n20784, n20785, n20786, n20787, n20788, n20789,
         n20790, n20791, n20792, n20793, n20794, n20795, n20796, n20797,
         n20798, n20799, n20800, n20801, n20802, n20803, n20804, n20805,
         n20806, n20807, n20808, n20809, n20810, n20811, n20812, n20813,
         n20814, n20815, n20816, n20817, n20818, n20819, n20820, n20821,
         n20822, n20823, n20824, n20825, n20826, n20827, n20828, n20829,
         n20830, n20831, n20832, n20833, n20834, n20835, n20836, n20837,
         n20838, n20839, n20840, n20841, n20842, n20843, n20844, n20845,
         n20846, n20847, n20848, n20849, n20850, n20851, n20852, n20853,
         n20854, n20855, n20856, n20857, n20858, n20859, n20860, n20861,
         n20862, n20863, n20864, n20865, n20866, n20867, n20868, n20869,
         n20870, n20871, n20872, n20873, n20874, n20875, n20876, n20877,
         n20878, n20879, n20880, n20881, n20882, n20883, n20884, n20885,
         n20886, n20887, n20888, n20889, n20890, n20891, n20892, n20893,
         n20894, n20895, n20896, n20897, n20898, n20899, n20900, n20901,
         n20902, n20903, n20904, n20905, n20906, n20907, n20908, n20909,
         n20910, n20911, n20912, n20913, n20914, n20915, n20916, n20917,
         n20918, n20919, n20920, n20921, n20922, n20923, n20924, n20925,
         n20926, n20927, n20928, n20929, n20930, n20931, n20932, n20933,
         n20934, n20935, n20936, n20937, n20938, n20939, n20940, n20941,
         n20942, n20943, n20944, n20945, n20946, n20947, n20948, n20949,
         n20950, n20951, n20952, n20953, n20954, n20955, n20956, n20957,
         n20958, n20959, n20960, n20961, n20962, n20963, n20964, n20965,
         n20966, n20967, n20968, n20969, n20970, n20971, n20972, n20973,
         n20974, n20975, n20976, n20977, n20978, n20979, n20980, n20981,
         n20982, n20983, n20984, n20985, n20986, n20987, n20988, n20989,
         n20990, n20991, n20992, n20993, n20994, n20995, n20996, n20997,
         n20998, n20999, n21000, n21001, n21002, n21003, n21004, n21005,
         n21006, n21007, n21008, n21009, n21010, n21011, n21012, n21013,
         n21014, n21015, n21016, n21017, n21018, n21019, n21020, n21021,
         n21022, n21023, n21024, n21025, n21026, n21027, n21028, n21029,
         n21030, n21031, n21032, n21033, n21034, n21035, n21036, n21037,
         n21038, n21039, n21040, n21041, n21042, n21043, n21044, n21045,
         n21046, n21047, n21048, n21049, n21050, n21051, n21052, n21053,
         n21054, n21055, n21056, n21057, n21058, n21059, n21060, n21061,
         n21062, n21063, n21064, n21065, n21066, n21067, n21068, n21069,
         n21070, n21071, n21072, n21073, n21074, n21075, n21076, n21077,
         n21078, n21079, n21080, n21081, n21082, n21083, n21084, n21085,
         n21086, n21087, n21088, n21089, n21090, n21091, n21092, n21093,
         n21094, n21095, n21096, n21097, n21098, n21099, n21100, n21101,
         n21102, n21103, n21104, n21105, n21106, n21107, n21108, n21109,
         n21110, n21111, n21112, n21113, n21114, n21115, n21116, n21117,
         n21118, n21119, n21120, n21121, n21122, n21123, n21124, n21125,
         n21126, n21127, n21128, n21129, n21130, n21131, n21132, n21133,
         n21134, n21135, n21136, n21137, n21138, n21139, n21140, n21141,
         n21142, n21143, n21144, n21145, n21146, n21147, n21148, n21149,
         n21150, n21151, n21152, n21153, n21154, n21155, n21156, n21157,
         n21158, n21159, n21160, n21161, n21162, n21163, n21164, n21165,
         n21166, n21167, n21168, n21169, n21170, n21171, n21172, n21173,
         n21174, n21175, n21176, n21177, n21178, n21179, n21180, n21181,
         n21182, n21183, n21184, n21185, n21186, n21187, n21188, n21189,
         n21190, n21191, n21192, n21193, n21194, n21195, n21196, n21197,
         n21198, n21199, n21200, n21201, n21202, n21203, n21204, n21205,
         n21206, n21207, n21208, n21209, n21210, n21211, n21212, n21213,
         n21214, n21215, n21216, n21217, n21218, n21219, n21220, n21221,
         n21222, n21223, n21224, n21225, n21226, n21227, n21228, n21229,
         n21230, n21231, n21232, n21233, n21234, n21235, n21236, n21237,
         n21238, n21239, n21240, n21241, n21242, n21243, n21244, n21245,
         n21246, n21247, n21248, n21249, n21250, n21251, n21252, n21253,
         n21254, n21255, n21256, n21257, n21258, n21259, n21260, n21261,
         n21262, n21263, n21264, n21265, n21266, n21267, n21268, n21269,
         n21270, n21271, n21272, n21273, n21274, n21275, n21276, n21277,
         n21278, n21279, n21280, n21281, n21282, n21283, n21284, n21285,
         n21286, n21287, n21288, n21289, n21290, n21291, n21292, n21293,
         n21294, n21295, n21296, n21297, n21298, n21299, n21300, n21301,
         n21302, n21303, n21304, n21305, n21306, n21307, n21308, n21309,
         n21310, n21311, n21312, n21313, n21314, n21315, n21316, n21317,
         n21318, n21319, n21320, n21321, n21322, n21323, n21324, n21325,
         n21326, n21327, n21328, n21329, n21330, n21331, n21332, n21333,
         n21334, n21335, n21336, n21337, n21338, n21339, n21340, n21341,
         n21342, n21343, n21344, n21345, n21346, n21347, n21348, n21349,
         n21350, n21351, n21352, n21353, n21354, n21355, n21356, n21357,
         n21358, n21359, n21360, n21361, n21362, n21363, n21364, n21365,
         n21366, n21367, n21368, n21369, n21370, n21371, n21372, n21373,
         n21374, n21375, n21376, n21377, n21378, n21379, n21380, n21381,
         n21382, n21383, n21384, n21385, n21386, n21387, n21388, n21389,
         n21390, n21391, n21392, n21393, n21394, n21395, n21396, n21397,
         n21398, n21399, n21400, n21401, n21402, n21403, n21404, n21405,
         n21406, n21407, n21408, n21409, n21410, n21411, n21412, n21413,
         n21414, n21415, n21416, n21417, n21418, n21419, n21420, n21421,
         n21422, n21423, n21424, n21425, n21426, n21427, n21428, n21429,
         n21430, n21431, n21432, n21433, n21434, n21435, n21436, n21437,
         n21438, n21439, n21440, n21441, n21442, n21443, n21444, n21445,
         n21446, n21447, n21448, n21449, n21450, n21451, n21452, n21453,
         n21454, n21455, n21456, n21457, n21458, n21459, n21460, n21461,
         n21462, n21463, n21464, n21465, n21466, n21467, n21468, n21469,
         n21470, n21471, n21472, n21473, n21474, n21475, n21476, n21477,
         n21478, n21479, n21480, n21481, n21482, n21483, n21484, n21485,
         n21486, n21487, n21488, n21489, n21490, n21491, n21492, n21493,
         n21494, n21495, n21496, n21497, n21498, n21499, n21500, n21501,
         n21502, n21503, n21504, n21505, n21506, n21507, n21508, n21509,
         n21510, n21511, n21512, n21513, n21514, n21515, n21516, n21517,
         n21518, n21519, n21520, n21521, n21522, n21523, n21524, n21525,
         n21526, n21527, n21528, n21529, n21530, n21531, n21532, n21533,
         n21534, n21535, n21536, n21537, n21538, n21539, n21540, n21541,
         n21542, n21543, n21544, n21545, n21546, n21547, n21548, n21549,
         n21550, n21551, n21552, n21553, n21554, n21555, n21556, n21557,
         n21558, n21559, n21560, n21561, n21562, n21563, n21564, n21565,
         n21566, n21567, n21568, n21569, n21570, n21571, n21572, n21573,
         n21574, n21575, n21576, n21577, n21578, n21579, n21580, n21581,
         n21582, n21583, n21584, n21585, n21586, n21587, n21588, n21589,
         n21590, n21591, n21592, n21593, n21594, n21595, n21596, n21597,
         n21598, n21599, n21600, n21601, n21602, n21603, n21604, n21605,
         n21606, n21607, n21608, n21609, n21610, n21611, n21612, n21613,
         n21614, n21615, n21616, n21617, n21618, n21619, n21620, n21621,
         n21622, n21623, n21624, n21625, n21626, n21627, n21628, n21629,
         n21630, n21631, n21632, n21633, n21634, n21635, n21636, n21637,
         n21638, n21639, n21640, n21641, n21642, n21643, n21644, n21645,
         n21646, n21647, n21648, n21649, n21650, n21651, n21652, n21653,
         n21654, n21655, n21656, n21657, n21658, n21659, n21660, n21661,
         n21662, n21663, n21664, n21665, n21666, n21667, n21668, n21669,
         n21670, n21671, n21672, n21673, n21674, n21675, n21676, n21677,
         n21678, n21679, n21680, n21681, n21682, n21683, n21684, n21685,
         n21686, n21687, n21688, n21689, n21690, n21691, n21692, n21693,
         n21694, n21695, n21696, n21697, n21698, n21699, n21700, n21701,
         n21702, n21703, n21704, n21705, n21706, n21707, n21708, n21709,
         n21710, n21711, n21712, n21713, n21714, n21715, n21716, n21717,
         n21718, n21719, n21720, n21721, n21722, n21723, n21724, n21725,
         n21726, n21727, n21728, n21729, n21730, n21731, n21732, n21733,
         n21734, n21735, n21736, n21737, n21738, n21739, n21740, n21741,
         n21742, n21743, n21744, n21745, n21746, n21747, n21748, n21749,
         n21750, n21751, n21752, n21753, n21754, n21755, n21756, n21757,
         n21758, n21759, n21760, n21761, n21762, n21763, n21764, n21765,
         n21766, n21767, n21768, n21769, n21770, n21771, n21772, n21773,
         n21774, n21775, n21776, n21777, n21778, n21779, n21780, n21781,
         n21782, n21783, n21784, n21785, n21786, n21787, n21788, n21789,
         n21790, n21791, n21792, n21793, n21794, n21795, n21796, n21797,
         n21798, n21799, n21800, n21801, n21802, n21803, n21804, n21805,
         n21806, n21807, n21808, n21809, n21810, n21811, n21812, n21813,
         n21814, n21815, n21816, n21817, n21818, n21819, n21820, n21821,
         n21822, n21823, n21824, n21825, n21826, n21827, n21828, n21829,
         n21830, n21831, n21832, n21833, n21834, n21835, n21836, n21837,
         n21838, n21839, n21840, n21841, n21842, n21843, n21844, n21845,
         n21846, n21847, n21848, n21849, n21850, n21851, n21852, n21853,
         n21854, n21855, n21856, n21857, n21858, n21859, n21860, n21861,
         n21862, n21863, n21864, n21865, n21866, n21867, n21868, n21869,
         n21870, n21871, n21872, n21873, n21874, n21875, n21876, n21877,
         n21878, n21879, n21880, n21881, n21882, n21883, n21884, n21885,
         n21886, n21887, n21888, n21889, n21890, n21891, n21892, n21893,
         n21894, n21895, n21896, n21897, n21898, n21899, n21900, n21901,
         n21902, n21903, n21904, n21905, n21906, n21907, n21908, n21909,
         n21910, n21911, n21912, n21913, n21914, n21915, n21916, n21917,
         n21918, n21919, n21920, n21921, n21922, n21923, n21924, n21925,
         n21926, n21927, n21928, n21929, n21930, n21931, n21932, n21933,
         n21934, n21935, n21936, n21937, n21938, n21939, n21940, n21941,
         n21942, n21943, n21944, n21945, n21946, n21947, n21948, n21949,
         n21950, n21951, n21952, n21953, n21954, n21955, n21956, n21957,
         n21958, n21959, n21960, n21961, n21962, n21963, n21964, n21965,
         n21966, n21967, n21968, n21969, n21970, n21971, n21972, n21973,
         n21974, n21975, n21976, n21977, n21978, n21979, n21980, n21981,
         n21982, n21983, n21984, n21985, n21986, n21987, n21988, n21989,
         n21990, n21991, n21992, n21993, n21994, n21995, n21996, n21997,
         n21998, n21999, n22000, n22001, n22002, n22003, n22004, n22005,
         n22006, n22007, n22008, n22009, n22010, n22011, n22012, n22013,
         n22014, n22015, n22016, n22017, n22018, n22019, n22020, n22021,
         n22022, n22023, n22024, n22025, n22026, n22027, n22028, n22029,
         n22030, n22031, n22032, n22033, n22034, n22035, n22036, n22037,
         n22038, n22039, n22040, n22041, n22042, n22043, n22044, n22045,
         n22046, n22047, n22048, n22049, n22050, n22051, n22052, n22053,
         n22054, n22055, n22056, n22057, n22058, n22059, n22060, n22061,
         n22062, n22063, n22064, n22065, n22066, n22067, n22068, n22069,
         n22070, n22071, n22072, n22073, n22074, n22075, n22076, n22077,
         n22078, n22079, n22080, n22081, n22082, n22083, n22084, n22085,
         n22086, n22087, n22088, n22089, n22090, n22091, n22092, n22093,
         n22094, n22095, n22096, n22097, n22098, n22099, n22100, n22101,
         n22102, n22103, n22104, n22105, n22106, n22107, n22108, n22109,
         n22110, n22111, n22112, n22113, n22114, n22115, n22116, n22117,
         n22118, n22119, n22120, n22121, n22122, n22123, n22124, n22125,
         n22126, n22127, n22128, n22129, n22130, n22131, n22132, n22133,
         n22134, n22135, n22136, n22137, n22138, n22139, n22140, n22141,
         n22142, n22143, n22144, n22145, n22146, n22147, n22148, n22149,
         n22150, n22151, n22152, n22153, n22154, n22155, n22156, n22157,
         n22158, n22159, n22160, n22161, n22162, n22163, n22164, n22165,
         n22166, n22167, n22168, n22169, n22170, n22171, n22172, n22173,
         n22174, n22175, n22176, n22177, n22178, n22179, n22180, n22181,
         n22182, n22183, n22184, n22185, n22186, n22187, n22188, n22189,
         n22190, n22191, n22192, n22193, n22194, n22195, n22196, n22197,
         n22198, n22199, n22200, n22201, n22202, n22203, n22204, n22205,
         n22206, n22207, n22208, n22209, n22210, n22211, n22212, n22213,
         n22214, n22215, n22216, n22217, n22218, n22219, n22220, n22221,
         n22222, n22223, n22224, n22225, n22226, n22227, n22228, n22229,
         n22230, n22231, n22232, n22233, n22234, n22235, n22236;

  NOR2_X2 U11151 ( .A1(n20843), .A2(n21111), .ZN(n20869) );
  AND2_X1 U11152 ( .A1(n14208), .A2(n14065), .ZN(n20671) );
  NAND3_X1 U11153 ( .A1(n9998), .A2(n10516), .A3(n11046), .ZN(n17730) );
  AOI21_X1 U11154 ( .B1(n9798), .B2(n20013), .A(n18857), .ZN(n20190) );
  NAND2_X1 U11155 ( .A1(n10302), .A2(n10303), .ZN(n17629) );
  XNOR2_X1 U11156 ( .A(n12519), .B(n9930), .ZN(n15888) );
  CLKBUF_X2 U11157 ( .A(n10780), .Z(n14477) );
  INV_X1 U11158 ( .A(n12335), .ZN(n13244) );
  BUF_X1 U11159 ( .A(n20440), .Z(n9722) );
  INV_X1 U11160 ( .A(n15300), .ZN(n21906) );
  INV_X1 U11161 ( .A(n11880), .ZN(n17561) );
  INV_X1 U11162 ( .A(n10660), .ZN(n18627) );
  NOR2_X1 U11163 ( .A1(n13935), .A2(n15091), .ZN(n13851) );
  AND2_X2 U11164 ( .A1(n14123), .A2(n10700), .ZN(n10732) );
  NAND2_X1 U11165 ( .A1(n11814), .A2(n20146), .ZN(n9783) );
  AND4_X1 U11166 ( .A1(n12266), .A2(n12265), .A3(n12264), .A4(n12263), .ZN(
        n12283) );
  NAND4_X1 U11167 ( .A1(n12204), .A2(n12203), .A3(n12202), .A4(n12201), .ZN(
        n12307) );
  AND2_X1 U11168 ( .A1(n10700), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n9729) );
  INV_X1 U11169 ( .A(n12259), .ZN(n13079) );
  INV_X1 U11170 ( .A(n12342), .ZN(n12741) );
  AND2_X2 U11171 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10700) );
  NAND2_X2 U11172 ( .A1(n13873), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12259) );
  CLKBUF_X1 U11173 ( .A(n18255), .Z(n9707) );
  NOR2_X1 U11174 ( .A1(n12005), .A2(n12004), .ZN(n18255) );
  CLKBUF_X1 U11175 ( .A(n20254), .Z(n9708) );
  NOR2_X1 U11176 ( .A1(n13629), .A2(n11713), .ZN(n20254) );
  INV_X1 U11177 ( .A(n13093), .ZN(n12392) );
  NAND2_X1 U11178 ( .A1(n12624), .A2(n12623), .ZN(n12658) );
  NAND2_X1 U11179 ( .A1(n10878), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n14497) );
  INV_X1 U11180 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10710) );
  AND2_X2 U11181 ( .A1(n10446), .A2(n12123), .ZN(n13075) );
  INV_X1 U11182 ( .A(n12654), .ZN(n12624) );
  CLKBUF_X2 U11183 ( .A(n11161), .Z(n11699) );
  AND2_X1 U11184 ( .A1(n10874), .A2(n10873), .ZN(n10875) );
  NAND2_X1 U11185 ( .A1(n10963), .A2(n10964), .ZN(n9942) );
  OAI21_X1 U11186 ( .B1(n17127), .B2(n12027), .A(n13776), .ZN(n17152) );
  INV_X1 U11187 ( .A(n17547), .ZN(n18616) );
  INV_X1 U11189 ( .A(n15545), .ZN(n10100) );
  NOR2_X1 U11190 ( .A1(n15556), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15543) );
  CLKBUF_X2 U11191 ( .A(n11160), .Z(n11243) );
  CLKBUF_X2 U11192 ( .A(n11471), .Z(n9737) );
  CLKBUF_X2 U11193 ( .A(n11472), .Z(n11689) );
  INV_X2 U11194 ( .A(n10322), .ZN(n13512) );
  NAND2_X1 U11195 ( .A1(n10321), .A2(n10319), .ZN(n11467) );
  NAND2_X1 U11196 ( .A1(n11049), .A2(n11351), .ZN(n10521) );
  NOR2_X1 U11197 ( .A1(n10981), .A2(n17744), .ZN(n20784) );
  INV_X2 U11199 ( .A(n12288), .ZN(n21334) );
  INV_X2 U11201 ( .A(n20376), .ZN(n9969) );
  NAND2_X1 U11202 ( .A1(n11456), .A2(n16523), .ZN(n12017) );
  OAI21_X1 U11203 ( .B1(n16703), .B2(n16690), .A(n16689), .ZN(n9960) );
  NOR3_X2 U11204 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n18267) );
  INV_X2 U11205 ( .A(n18615), .ZN(n14232) );
  AND2_X1 U11206 ( .A1(n17271), .A2(n19259), .ZN(n18942) );
  OR2_X1 U11207 ( .A1(n21910), .A2(n13528), .ZN(n21170) );
  OAI21_X1 U11208 ( .B1(n15896), .B2(n12881), .A(n12699), .ZN(n15180) );
  AND2_X1 U11210 ( .A1(n10065), .A2(n11150), .ZN(n16772) );
  AND2_X1 U11211 ( .A1(n10226), .A2(n10227), .ZN(n16541) );
  AND2_X1 U11212 ( .A1(n20457), .A2(n21111), .ZN(n20502) );
  NOR2_X1 U11213 ( .A1(n20671), .A2(n20373), .ZN(n20506) );
  INV_X1 U11214 ( .A(n20547), .ZN(n20570) );
  OAI21_X1 U11215 ( .B1(n20679), .B2(n20682), .A(n20941), .ZN(n20709) );
  OAI21_X1 U11216 ( .B1(n20757), .B2(n20773), .A(n20941), .ZN(n20776) );
  AND2_X1 U11217 ( .A1(n20935), .A2(n20779), .ZN(n20995) );
  NAND2_X1 U11218 ( .A1(n10166), .A2(n9813), .ZN(n19147) );
  INV_X1 U11219 ( .A(n21212), .ZN(n17648) );
  AND2_X1 U11220 ( .A1(n13941), .A2(n14788), .ZN(n15194) );
  OR2_X1 U11221 ( .A1(n17609), .A2(n21146), .ZN(n21153) );
  AOI211_X1 U11222 ( .C1(n17741), .C2(n16857), .A(n16856), .B(n16855), .ZN(
        n16858) );
  OR2_X1 U11223 ( .A1(n21091), .A2(n21111), .ZN(n20670) );
  NAND2_X1 U11224 ( .A1(n20836), .A2(n21111), .ZN(n20933) );
  NAND2_X1 U11225 ( .A1(n20935), .A2(n20873), .ZN(n20999) );
  INV_X1 U11226 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n21106) );
  OR2_X1 U11227 ( .A1(n19239), .A2(n19188), .ZN(n19105) );
  INV_X1 U11228 ( .A(n19128), .ZN(n19118) );
  NAND2_X1 U11229 ( .A1(n19147), .A2(n19327), .ZN(n19079) );
  OR2_X1 U11230 ( .A1(n14715), .A2(n17082), .ZN(n9709) );
  OR2_X1 U11231 ( .A1(n20884), .A2(n11053), .ZN(n9710) );
  OR2_X1 U11232 ( .A1(n10066), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9711) );
  INV_X1 U11233 ( .A(n11911), .ZN(n11861) );
  NOR2_X2 U11234 ( .A1(n14147), .A2(n10565), .ZN(n14359) );
  NOR2_X2 U11235 ( .A1(n14843), .A2(n14825), .ZN(n14824) );
  OR2_X1 U11236 ( .A1(n10986), .A2(n13778), .ZN(n11002) );
  AND2_X1 U11237 ( .A1(n10986), .A2(n13790), .ZN(n10975) );
  NOR2_X2 U11238 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n18258), .ZN(n18235) );
  NAND2_X1 U11239 ( .A1(n10878), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n9712) );
  NOR2_X2 U11240 ( .A1(n18522), .A2(n18521), .ZN(n18520) );
  NAND2_X1 U11241 ( .A1(n12300), .A2(n12288), .ZN(n13385) );
  NAND2_X2 U11242 ( .A1(n9956), .A2(n9955), .ZN(n10966) );
  AOI221_X1 U11243 ( .B1(n18657), .B2(n18670), .C1(n18765), .C2(n18670), .A(
        P3_EBX_REG_2__SCAN_IN), .ZN(n18659) );
  NAND2_X1 U11244 ( .A1(n19532), .A2(n18765), .ZN(n11975) );
  NOR2_X4 U11245 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10394) );
  AND2_X1 U11246 ( .A1(n10700), .A2(n10750), .ZN(n9714) );
  NOR2_X2 U11249 ( .A1(n9727), .A2(n10194), .ZN(n20888) );
  NAND2_X2 U11250 ( .A1(n11140), .A2(n11139), .ZN(n11143) );
  OAI21_X2 U11251 ( .B1(n15105), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n12414), 
        .ZN(n10455) );
  INV_X2 U11253 ( .A(n22236), .ZN(n9718) );
  NOR2_X1 U11254 ( .A1(n11001), .A2(n17733), .ZN(n20449) );
  AND2_X1 U11255 ( .A1(n10693), .A2(n10710), .ZN(n9719) );
  AND2_X1 U11256 ( .A1(n10693), .A2(n10710), .ZN(n9720) );
  NAND2_X1 U11257 ( .A1(n10229), .A2(n10230), .ZN(n10405) );
  AND2_X1 U11258 ( .A1(n10196), .A2(n10195), .ZN(n9967) );
  NAND2_X1 U11259 ( .A1(n16054), .A2(n9864), .ZN(n15998) );
  INV_X2 U11260 ( .A(n21174), .ZN(n21263) );
  INV_X2 U11261 ( .A(n11346), .ZN(n10020) );
  NAND2_X1 U11262 ( .A1(n14271), .A2(n10146), .ZN(n14366) );
  INV_X1 U11263 ( .A(n20671), .ZN(n21090) );
  INV_X1 U11264 ( .A(n11351), .ZN(n9721) );
  NAND2_X1 U11265 ( .A1(n10396), .A2(n10395), .ZN(n9998) );
  INV_X4 U11266 ( .A(n15554), .ZN(n15545) );
  OR2_X2 U11267 ( .A1(n10194), .A2(n11002), .ZN(n11050) );
  INV_X1 U11268 ( .A(n19235), .ZN(n10167) );
  OR2_X1 U11269 ( .A1(n17146), .A2(n10990), .ZN(n10981) );
  AND2_X1 U11270 ( .A1(n10987), .A2(n17146), .ZN(n20580) );
  OR2_X1 U11271 ( .A1(n17930), .A2(n19535), .ZN(n19239) );
  NOR2_X1 U11272 ( .A1(n18083), .A2(n18504), .ZN(n18461) );
  INV_X1 U11273 ( .A(n10975), .ZN(n9727) );
  OR2_X1 U11274 ( .A1(n12402), .A2(n12401), .ZN(n12415) );
  NAND2_X1 U11275 ( .A1(n13817), .A2(n17793), .ZN(n20303) );
  AND2_X1 U11276 ( .A1(n10965), .A2(n10967), .ZN(n10397) );
  OAI211_X1 U11277 ( .C1(n10957), .C2(n11040), .A(n10945), .B(n10944), .ZN(
        n10951) );
  NAND2_X1 U11278 ( .A1(n12048), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10957) );
  CLKBUF_X1 U11279 ( .A(n11705), .Z(n17779) );
  CLKBUF_X1 U11280 ( .A(n9737), .Z(n11688) );
  NAND2_X2 U11281 ( .A1(n9970), .A2(n9969), .ZN(n10926) );
  CLKBUF_X3 U11283 ( .A(n13383), .Z(n13937) );
  OR2_X1 U11284 ( .A1(n11894), .A2(n11893), .ZN(n18680) );
  AND2_X2 U11285 ( .A1(n21361), .A2(n12672), .ZN(n13857) );
  NOR2_X1 U11286 ( .A1(n14109), .A2(n14108), .ZN(n17287) );
  NAND2_X1 U11287 ( .A1(n10006), .A2(n9790), .ZN(n17296) );
  NAND4_X2 U11288 ( .A1(n11860), .A2(n11859), .A3(n11858), .A4(n11857), .ZN(
        n18765) );
  AND2_X1 U11289 ( .A1(n13350), .A2(n12297), .ZN(n12301) );
  AND4_X1 U11290 ( .A1(n20400), .A2(n13819), .A3(n20415), .A4(n12056), .ZN(
        n10907) );
  NAND2_X2 U11291 ( .A1(n21334), .A2(n12289), .ZN(n15091) );
  NAND2_X1 U11292 ( .A1(n21334), .A2(n15303), .ZN(n15094) );
  AND2_X1 U11293 ( .A1(n15303), .A2(n12288), .ZN(n13383) );
  BUF_X2 U11294 ( .A(n12298), .Z(n15303) );
  INV_X1 U11295 ( .A(n12297), .ZN(n12300) );
  INV_X2 U11296 ( .A(n12293), .ZN(n12296) );
  INV_X1 U11297 ( .A(n10875), .ZN(n10894) );
  INV_X4 U11298 ( .A(n9718), .ZN(n18591) );
  INV_X2 U11299 ( .A(n9718), .ZN(n18413) );
  BUF_X2 U11300 ( .A(n11066), .Z(n14493) );
  INV_X4 U11301 ( .A(n18611), .ZN(n18586) );
  CLKBUF_X2 U11302 ( .A(n12944), .Z(n13061) );
  CLKBUF_X2 U11303 ( .A(n13079), .Z(n13056) );
  INV_X4 U11304 ( .A(n18599), .ZN(n18628) );
  CLKBUF_X2 U11305 ( .A(n12364), .Z(n13255) );
  CLKBUF_X2 U11306 ( .A(n12267), .Z(n13254) );
  INV_X4 U11307 ( .A(n18585), .ZN(n18613) );
  NAND2_X2 U11308 ( .A1(n13870), .A2(n12112), .ZN(n12381) );
  AND2_X2 U11309 ( .A1(n12128), .A2(n12123), .ZN(n13125) );
  NAND2_X1 U11310 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n21915), .ZN(n21876) );
  INV_X2 U11311 ( .A(n17561), .ZN(n9723) );
  AND2_X2 U11312 ( .A1(n14123), .A2(n10703), .ZN(n10781) );
  INV_X4 U11313 ( .A(n18556), .ZN(n9724) );
  CLKBUF_X2 U11314 ( .A(n9785), .Z(n13256) );
  INV_X4 U11315 ( .A(n9783), .ZN(n9726) );
  AND2_X2 U11316 ( .A1(n12121), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10192) );
  AND2_X1 U11317 ( .A1(n17149), .A2(n10701), .ZN(n10813) );
  INV_X4 U11319 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14126) );
  NOR2_X1 U11320 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20880) );
  XNOR2_X1 U11321 ( .A(n10232), .B(n9860), .ZN(n16891) );
  XOR2_X1 U11322 ( .A(n12017), .B(n9799), .Z(n9832) );
  XNOR2_X1 U11323 ( .A(n10456), .B(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15626) );
  AOI21_X1 U11324 ( .B1(n10127), .B2(n10126), .A(n10123), .ZN(n16599) );
  AOI21_X1 U11325 ( .B1(n14722), .B2(n20357), .A(n14721), .ZN(n14723) );
  NOR2_X1 U11326 ( .A1(n16580), .A2(n9818), .ZN(n16835) );
  NOR2_X1 U11327 ( .A1(n16616), .A2(n12102), .ZN(n10232) );
  AOI21_X1 U11328 ( .B1(n14730), .B2(n11150), .A(n13522), .ZN(n14735) );
  OR2_X1 U11329 ( .A1(n16879), .A2(n16762), .ZN(n10682) );
  OAI21_X1 U11330 ( .B1(n16798), .B2(n16737), .A(n9939), .ZN(n9938) );
  AND2_X1 U11331 ( .A1(n14759), .A2(n14758), .ZN(n16907) );
  XNOR2_X1 U11332 ( .A(n9959), .B(n13523), .ZN(n14715) );
  NAND2_X1 U11333 ( .A1(n10493), .A2(n10491), .ZN(n15386) );
  AOI21_X1 U11334 ( .B1(n14762), .B2(n9807), .A(n10557), .ZN(n16603) );
  OAI21_X1 U11335 ( .B1(n10004), .B2(n9778), .A(n16864), .ZN(n10003) );
  NOR2_X1 U11336 ( .A1(n10004), .A2(n9778), .ZN(n16617) );
  XNOR2_X1 U11337 ( .A(n16542), .B(n9940), .ZN(n16798) );
  AND2_X1 U11338 ( .A1(n9988), .A2(n15388), .ZN(n9987) );
  NAND2_X1 U11339 ( .A1(n13522), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9959) );
  NAND2_X1 U11340 ( .A1(n10034), .A2(n9862), .ZN(n14762) );
  OAI211_X1 U11341 ( .C1(n10227), .C2(n16551), .A(n16550), .B(n10157), .ZN(
        n16542) );
  AND3_X1 U11342 ( .A1(n9965), .A2(n9847), .A3(n9964), .ZN(n16911) );
  NAND2_X1 U11343 ( .A1(n16673), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n16674) );
  NAND2_X1 U11344 ( .A1(n10176), .A2(n10175), .ZN(n15402) );
  NAND2_X1 U11345 ( .A1(n10177), .A2(n15554), .ZN(n15422) );
  NAND2_X1 U11346 ( .A1(n15423), .A2(n15383), .ZN(n15415) );
  NAND2_X1 U11347 ( .A1(n10047), .A2(n10046), .ZN(n10227) );
  NAND2_X1 U11348 ( .A1(n12603), .A2(n10498), .ZN(n10493) );
  OAI21_X1 U11349 ( .B1(n9801), .B2(n16576), .A(n16577), .ZN(n16570) );
  AOI21_X1 U11350 ( .B1(n16725), .B2(n16723), .A(n16688), .ZN(n16717) );
  NAND2_X1 U11351 ( .A1(n12602), .A2(n10441), .ZN(n12603) );
  OAI21_X1 U11352 ( .B1(n10405), .B2(n9833), .A(n10235), .ZN(n16649) );
  OR2_X1 U11353 ( .A1(n14602), .A2(n14601), .ZN(n14606) );
  CLKBUF_X1 U11354 ( .A(n14821), .Z(n14822) );
  NAND2_X1 U11355 ( .A1(n9984), .A2(n9983), .ZN(n15556) );
  NAND2_X1 U11356 ( .A1(n9994), .A2(n9995), .ZN(n15462) );
  OR2_X1 U11357 ( .A1(n11703), .A2(n11255), .ZN(n16310) );
  XNOR2_X1 U11358 ( .A(n13514), .B(n13513), .ZN(n15927) );
  NAND2_X1 U11359 ( .A1(n9985), .A2(n15562), .ZN(n9984) );
  NAND2_X1 U11360 ( .A1(n13514), .A2(n11704), .ZN(n14741) );
  NAND2_X1 U11361 ( .A1(n9918), .A2(n10097), .ZN(n12602) );
  OAI21_X1 U11362 ( .B1(n16404), .B2(n16487), .A(n16403), .ZN(n10585) );
  INV_X1 U11363 ( .A(n15467), .ZN(n15514) );
  AOI211_X1 U11364 ( .C1(n16490), .C2(BUF2_REG_28__SCAN_IN), .A(n16408), .B(
        n16407), .ZN(n16409) );
  AND2_X1 U11365 ( .A1(n11253), .A2(n11254), .ZN(n11703) );
  CLKBUF_X1 U11366 ( .A(n11253), .Z(n15957) );
  AND2_X1 U11367 ( .A1(n10196), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10345) );
  NAND2_X1 U11368 ( .A1(n10170), .A2(n12594), .ZN(n15467) );
  NOR3_X1 U11369 ( .A1(n15998), .A2(n15958), .A3(n10535), .ZN(n11253) );
  NOR2_X1 U11370 ( .A1(n15998), .A2(n15999), .ZN(n15983) );
  NAND2_X1 U11371 ( .A1(n15955), .A2(n15954), .ZN(n16770) );
  OR2_X1 U11372 ( .A1(n15998), .A2(n10534), .ZN(n10533) );
  XNOR2_X1 U11373 ( .A(n11352), .B(n22168), .ZN(n9961) );
  NAND3_X1 U11374 ( .A1(n10021), .A2(n10016), .A3(n11342), .ZN(n17065) );
  CLKBUF_X1 U11375 ( .A(n14931), .Z(n14932) );
  AOI21_X1 U11376 ( .B1(n17662), .B2(n17664), .A(n17663), .ZN(n17657) );
  NAND2_X1 U11377 ( .A1(n16685), .A2(n10673), .ZN(n10140) );
  NAND2_X1 U11378 ( .A1(n16352), .A2(n10603), .ZN(n10147) );
  NAND2_X1 U11379 ( .A1(n10186), .A2(n10184), .ZN(n17067) );
  NOR2_X2 U11380 ( .A1(n12104), .A2(n16073), .ZN(n16054) );
  AND2_X1 U11381 ( .A1(n14381), .A2(n9877), .ZN(n16356) );
  NAND2_X1 U11382 ( .A1(n20713), .A2(n21111), .ZN(n20758) );
  NAND2_X1 U11383 ( .A1(n17333), .A2(n17269), .ZN(n17334) );
  NAND2_X1 U11384 ( .A1(n9721), .A2(n10198), .ZN(n11141) );
  AND2_X1 U11385 ( .A1(n10114), .A2(n10112), .ZN(n10443) );
  AND2_X1 U11386 ( .A1(n20506), .A2(n21099), .ZN(n20457) );
  AND2_X1 U11387 ( .A1(n12587), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17663) );
  NAND2_X1 U11388 ( .A1(n18968), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n18956) );
  AND2_X1 U11389 ( .A1(n20935), .A2(n21099), .ZN(n20836) );
  NAND2_X1 U11390 ( .A1(n20671), .A2(n21100), .ZN(n21092) );
  NOR2_X1 U11391 ( .A1(n16749), .A2(n11452), .ZN(n11347) );
  AND2_X1 U11392 ( .A1(n20671), .A2(n20373), .ZN(n20935) );
  NAND2_X1 U11393 ( .A1(n9941), .A2(n11120), .ZN(n16749) );
  AND2_X1 U11394 ( .A1(n14114), .A2(n15181), .ZN(n10275) );
  INV_X1 U11395 ( .A(n21100), .ZN(n20373) );
  NAND2_X1 U11396 ( .A1(n9980), .A2(n22186), .ZN(n18957) );
  OR2_X1 U11397 ( .A1(n14063), .A2(n14064), .ZN(n14065) );
  AND3_X1 U11398 ( .A1(n10044), .A2(n10042), .A3(n10043), .ZN(n10040) );
  AND2_X1 U11399 ( .A1(n11431), .A2(n11433), .ZN(n16036) );
  OR2_X1 U11400 ( .A1(n15554), .A2(n12599), .ZN(n15468) );
  AND2_X1 U11401 ( .A1(n14210), .A2(n10145), .ZN(n14064) );
  OR2_X1 U11402 ( .A1(n14211), .A2(n14062), .ZN(n10145) );
  AND2_X1 U11403 ( .A1(n14049), .A2(n14048), .ZN(n14051) );
  NAND3_X1 U11404 ( .A1(n12513), .A2(n9923), .A3(n9921), .ZN(n12581) );
  NAND2_X1 U11405 ( .A1(n10440), .A2(n12513), .ZN(n12548) );
  OAI21_X1 U11406 ( .B1(n11050), .B2(n11051), .A(n9909), .ZN(n11055) );
  CLKBUF_X1 U11407 ( .A(n15888), .Z(n21330) );
  AOI22_X1 U11408 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20449), .B1(
        n20543), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11004) );
  NAND2_X1 U11409 ( .A1(n10013), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17313) );
  NOR2_X1 U11410 ( .A1(n10182), .A2(n10991), .ZN(n20641) );
  AND2_X1 U11411 ( .A1(n19450), .A2(n19185), .ZN(n19187) );
  BUF_X2 U11412 ( .A(n10991), .Z(n17733) );
  NAND2_X1 U11413 ( .A1(n20023), .A2(n20179), .ZN(n17930) );
  INV_X1 U11414 ( .A(n13801), .ZN(n17104) );
  INV_X1 U11415 ( .A(n13364), .ZN(n13493) );
  NAND2_X1 U11416 ( .A1(n10437), .A2(n12468), .ZN(n15893) );
  NAND2_X1 U11417 ( .A1(n10269), .A2(n12538), .ZN(n13828) );
  NAND2_X1 U11418 ( .A1(n17736), .A2(n13773), .ZN(n20368) );
  AND2_X1 U11419 ( .A1(n13337), .A2(n14788), .ZN(n13364) );
  XNOR2_X1 U11420 ( .A(n17308), .B(n10387), .ZN(n19199) );
  AND2_X1 U11421 ( .A1(n17255), .A2(n9846), .ZN(n17257) );
  AND2_X1 U11422 ( .A1(n10525), .A2(n14338), .ZN(n10524) );
  NAND3_X1 U11423 ( .A1(n10956), .A2(n10955), .A3(n10968), .ZN(n11157) );
  XNOR2_X1 U11424 ( .A(n12445), .B(n21470), .ZN(n13864) );
  OAI221_X1 U11425 ( .B1(n18259), .B2(n9707), .C1(n18183), .C2(n9707), .A(
        P3_EBX_REG_9__SCAN_IN), .ZN(n18181) );
  NAND2_X2 U11426 ( .A1(n15930), .A2(n11724), .ZN(n20271) );
  NOR2_X1 U11427 ( .A1(n11180), .A2(n14281), .ZN(n10525) );
  NOR2_X2 U11428 ( .A1(n19978), .A2(n19986), .ZN(n19488) );
  AND2_X1 U11429 ( .A1(n14701), .A2(n9843), .ZN(n16225) );
  OR2_X1 U11430 ( .A1(n14135), .A2(n13816), .ZN(n13817) );
  NAND2_X1 U11431 ( .A1(n10369), .A2(n10368), .ZN(n19986) );
  INV_X2 U11432 ( .A(n18853), .ZN(n18850) );
  NAND2_X1 U11433 ( .A1(n9942), .A2(n10397), .ZN(n10956) );
  INV_X1 U11434 ( .A(n19349), .ZN(n19978) );
  OR2_X1 U11435 ( .A1(n12446), .A2(n12717), .ZN(n12421) );
  INV_X2 U11436 ( .A(n13716), .ZN(n20348) );
  INV_X2 U11437 ( .A(n18900), .ZN(n18919) );
  AND2_X1 U11438 ( .A1(n11178), .A2(n11177), .ZN(n14259) );
  NAND2_X1 U11439 ( .A1(n10633), .A2(n9915), .ZN(n11360) );
  NAND2_X1 U11440 ( .A1(n16282), .A2(n11485), .ZN(n11493) );
  OR2_X1 U11441 ( .A1(n14022), .A2(n13979), .ZN(n10349) );
  NOR2_X1 U11442 ( .A1(n14188), .A2(n14176), .ZN(n14022) );
  NAND2_X1 U11443 ( .A1(n17359), .A2(n17301), .ZN(n19233) );
  AND2_X1 U11444 ( .A1(n11330), .A2(n11329), .ZN(n11319) );
  OAI21_X1 U11445 ( .B1(n11291), .B2(n11288), .A(n11290), .ZN(n11330) );
  OR2_X2 U11446 ( .A1(n17407), .A2(n18802), .ZN(n19185) );
  AND2_X1 U11447 ( .A1(n12041), .A2(n10923), .ZN(n11161) );
  AND2_X1 U11448 ( .A1(n10628), .A2(n11267), .ZN(n11291) );
  NOR4_X2 U11449 ( .A1(n19532), .A2(n14026), .A3(n18680), .A4(n11968), .ZN(
        n17919) );
  AND2_X1 U11450 ( .A1(n13815), .A2(n9971), .ZN(n10936) );
  CLKBUF_X1 U11451 ( .A(n10927), .Z(n11712) );
  AND2_X1 U11452 ( .A1(n10661), .A2(n13614), .ZN(n11705) );
  AND4_X1 U11453 ( .A1(n11499), .A2(n11498), .A3(n11497), .A4(n11496), .ZN(
        n16254) );
  AND2_X1 U11454 ( .A1(n13400), .A2(n12302), .ZN(n13346) );
  NAND2_X1 U11455 ( .A1(n18765), .A2(n11965), .ZN(n14026) );
  CLKBUF_X1 U11456 ( .A(n13400), .Z(n13485) );
  NAND2_X1 U11457 ( .A1(n9750), .A2(n9812), .ZN(n9957) );
  AND2_X1 U11458 ( .A1(n12063), .A2(n17165), .ZN(n13814) );
  AND2_X1 U11459 ( .A1(n10918), .A2(n10908), .ZN(n9999) );
  AND2_X1 U11460 ( .A1(n10933), .A2(n9952), .ZN(n10064) );
  AND2_X2 U11461 ( .A1(n10909), .A2(n10907), .ZN(n12041) );
  NAND2_X1 U11462 ( .A1(n11288), .A2(n11289), .ZN(n11290) );
  AND2_X1 U11463 ( .A1(n17295), .A2(n17278), .ZN(n17226) );
  OR2_X1 U11464 ( .A1(n10746), .A2(n10747), .ZN(n11486) );
  NAND2_X1 U11465 ( .A1(n12289), .A2(n12288), .ZN(n15300) );
  CLKBUF_X2 U11466 ( .A(n9970), .Z(n9736) );
  AND3_X1 U11467 ( .A1(n11879), .A2(n11878), .A3(n11877), .ZN(n19543) );
  CLKBUF_X1 U11468 ( .A(n12303), .Z(n13860) );
  NAND2_X1 U11469 ( .A1(n12300), .A2(n13350), .ZN(n12313) );
  CLKBUF_X1 U11470 ( .A(n12307), .Z(n13852) );
  INV_X1 U11471 ( .A(n10894), .ZN(n11462) );
  INV_X2 U11472 ( .A(n10902), .ZN(n20400) );
  NAND2_X1 U11473 ( .A1(n10211), .A2(n10210), .ZN(n11479) );
  BUF_X1 U11474 ( .A(n10902), .Z(n12040) );
  AND2_X1 U11475 ( .A1(n10287), .A2(n14172), .ZN(n9977) );
  NOR2_X1 U11476 ( .A1(n17879), .A2(n17836), .ZN(n17880) );
  AND4_X1 U11477 ( .A1(n11865), .A2(n11864), .A3(n11863), .A4(n11862), .ZN(
        n11879) );
  INV_X1 U11478 ( .A(n10900), .ZN(n13779) );
  BUF_X2 U11479 ( .A(n20376), .Z(n9731) );
  INV_X1 U11480 ( .A(n20415), .ZN(n10908) );
  NOR2_X1 U11481 ( .A1(n19066), .A2(n19072), .ZN(n19053) );
  NAND2_X1 U11482 ( .A1(n9907), .A2(n9905), .ZN(n10902) );
  NAND2_X1 U11483 ( .A1(n10843), .A2(n10842), .ZN(n12056) );
  NAND4_X2 U11484 ( .A1(n12161), .A2(n12160), .A3(n12159), .A4(n12158), .ZN(
        n12672) );
  NAND4_X1 U11485 ( .A1(n12257), .A2(n12256), .A3(n12255), .A4(n12254), .ZN(
        n12298) );
  NAND4_X2 U11486 ( .A1(n12181), .A2(n12180), .A3(n12179), .A4(n12178), .ZN(
        n12293) );
  AND4_X1 U11487 ( .A1(n12245), .A2(n12244), .A3(n12243), .A4(n12242), .ZN(
        n12256) );
  AND4_X1 U11488 ( .A1(n12230), .A2(n12229), .A3(n12228), .A4(n12227), .ZN(
        n12236) );
  AND4_X1 U11489 ( .A1(n12146), .A2(n12145), .A3(n12144), .A4(n12143), .ZN(
        n12161) );
  AND4_X1 U11490 ( .A1(n12191), .A2(n12190), .A3(n12189), .A4(n12188), .ZN(
        n12203) );
  AND4_X1 U11491 ( .A1(n12196), .A2(n12195), .A3(n12194), .A4(n12193), .ZN(
        n12202) );
  AND4_X1 U11492 ( .A1(n12166), .A2(n12165), .A3(n12164), .A4(n12163), .ZN(
        n12181) );
  NAND2_X1 U11493 ( .A1(n10857), .A2(n10856), .ZN(n10900) );
  NAND4_X1 U11494 ( .A1(n10841), .A2(n10840), .A3(n10839), .A4(n10838), .ZN(
        n10910) );
  AND4_X1 U11495 ( .A1(n12221), .A2(n12220), .A3(n12219), .A4(n12218), .ZN(
        n12222) );
  AND4_X1 U11496 ( .A1(n12170), .A2(n12169), .A3(n12168), .A4(n12167), .ZN(
        n12180) );
  AND4_X1 U11497 ( .A1(n12253), .A2(n12252), .A3(n12251), .A4(n12250), .ZN(
        n12254) );
  AND4_X1 U11498 ( .A1(n12249), .A2(n12248), .A3(n12247), .A4(n12246), .ZN(
        n12255) );
  AND4_X1 U11499 ( .A1(n12279), .A2(n12278), .A3(n12277), .A4(n12276), .ZN(
        n12280) );
  AND3_X1 U11500 ( .A1(n12275), .A2(n12274), .A3(n12273), .ZN(n12281) );
  AND4_X1 U11501 ( .A1(n12127), .A2(n12126), .A3(n12125), .A4(n12124), .ZN(
        n12140) );
  AOI22_X1 U11502 ( .A1(n12549), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12186), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12120) );
  AND4_X1 U11503 ( .A1(n12154), .A2(n12153), .A3(n12152), .A4(n12151), .ZN(
        n12159) );
  AND4_X1 U11504 ( .A1(n12150), .A2(n12149), .A3(n12148), .A4(n12147), .ZN(
        n12160) );
  AND4_X1 U11505 ( .A1(n12200), .A2(n12199), .A3(n12198), .A4(n12197), .ZN(
        n12201) );
  NAND2_X2 U11506 ( .A1(n21140), .A2(n21030), .ZN(n21080) );
  AND2_X1 U11507 ( .A1(n14666), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11066) );
  INV_X2 U11508 ( .A(n17904), .ZN(U215) );
  AND3_X1 U11509 ( .A1(n10726), .A2(n10725), .A3(n10724), .ZN(n10729) );
  AND2_X2 U11510 ( .A1(n11823), .A2(n18270), .ZN(n18585) );
  INV_X2 U11511 ( .A(n17913), .ZN(n17915) );
  NAND2_X1 U11512 ( .A1(n11823), .A2(n14031), .ZN(n18556) );
  NAND2_X2 U11513 ( .A1(n11829), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n18611) );
  NAND2_X2 U11514 ( .A1(n11814), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n18599) );
  CLKBUF_X3 U11515 ( .A(n10828), .Z(n14646) );
  NAND2_X2 U11516 ( .A1(n12128), .A2(n10192), .ZN(n12379) );
  OR3_X2 U11517 ( .A1(n20140), .A2(P3_STATE2_REG_0__SCAN_IN), .A3(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n14191) );
  AND2_X2 U11518 ( .A1(n10868), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10877) );
  AND2_X2 U11519 ( .A1(n10693), .A2(n10710), .ZN(n14664) );
  AND2_X1 U11520 ( .A1(n14126), .A2(n10224), .ZN(n14123) );
  AND3_X1 U11521 ( .A1(n20157), .A2(n17459), .A3(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11829) );
  AND2_X2 U11522 ( .A1(n10394), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n9730) );
  AND3_X1 U11523 ( .A1(n10260), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A3(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11814) );
  AND2_X2 U11524 ( .A1(n15871), .A2(n10446), .ZN(n9785) );
  NAND2_X2 U11525 ( .A1(n13870), .A2(n12113), .ZN(n12261) );
  AND2_X2 U11526 ( .A1(n10394), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10828) );
  AND2_X1 U11527 ( .A1(n12114), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12129) );
  AND3_X2 U11528 ( .A1(n10224), .A2(n10586), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10865) );
  AND2_X1 U11529 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n18270) );
  INV_X2 U11530 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n12682) );
  NOR2_X1 U11531 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n19995) );
  AND2_X1 U11532 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12123) );
  NOR2_X1 U11533 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12113) );
  NOR2_X2 U11534 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10446) );
  AND2_X1 U11535 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12134) );
  NOR2_X1 U11536 ( .A1(n11467), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n11471) );
  NAND2_X1 U11537 ( .A1(n18270), .A2(n11819), .ZN(n11880) );
  NAND2_X1 U11538 ( .A1(n9969), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10922) );
  AND2_X2 U11539 ( .A1(n10700), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10866) );
  AND2_X2 U11540 ( .A1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n12692), .ZN(
        n12686) );
  INV_X4 U11541 ( .A(n11937), .ZN(n17550) );
  AND2_X1 U11542 ( .A1(n11829), .A2(n20146), .ZN(n11937) );
  XNOR2_X2 U11543 ( .A(n12543), .B(n15752), .ZN(n14072) );
  NAND2_X2 U11544 ( .A1(n12542), .A2(n12541), .ZN(n12543) );
  XNOR2_X2 U11545 ( .A(n12409), .B(n12417), .ZN(n21438) );
  AND2_X2 U11546 ( .A1(n14126), .A2(n10868), .ZN(n14503) );
  OAI21_X1 U11547 ( .B1(n10957), .B2(n17751), .A(n9824), .ZN(n11159) );
  AND4_X1 U11548 ( .A1(n11026), .A2(n11025), .A3(n11024), .A4(n11023), .ZN(
        n11034) );
  NAND2_X1 U11549 ( .A1(n10926), .A2(n10919), .ZN(n11256) );
  INV_X1 U11550 ( .A(n10926), .ZN(n10927) );
  NOR2_X2 U11551 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n18063), .ZN(n18046) );
  NAND2_X1 U11552 ( .A1(n10486), .A2(n10485), .ZN(n20376) );
  AND2_X1 U11553 ( .A1(n10693), .A2(n10710), .ZN(n9732) );
  AND2_X1 U11554 ( .A1(n10693), .A2(n10710), .ZN(n9733) );
  XNOR2_X1 U11555 ( .A(n12532), .B(n12533), .ZN(n13825) );
  NAND2_X1 U11556 ( .A1(n14041), .A2(n13801), .ZN(n10194) );
  NOR2_X2 U11557 ( .A1(n9781), .A2(n10576), .ZN(n15952) );
  OR2_X2 U11558 ( .A1(n15996), .A2(n15997), .ZN(n9781) );
  AND2_X1 U11559 ( .A1(n16596), .A2(n20357), .ZN(n10127) );
  NAND2_X1 U11560 ( .A1(n10318), .A2(n9898), .ZN(n16596) );
  INV_X1 U11561 ( .A(n9736), .ZN(n10898) );
  NOR2_X2 U11562 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n18039), .ZN(n18025) );
  NOR2_X2 U11563 ( .A1(n11003), .A2(n11002), .ZN(n20543) );
  NAND2_X1 U11564 ( .A1(n17146), .A2(n17104), .ZN(n11003) );
  NAND2_X1 U11565 ( .A1(n10921), .A2(n13814), .ZN(n10941) );
  INV_X1 U11566 ( .A(n11467), .ZN(n9970) );
  AND2_X1 U11567 ( .A1(n14646), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10780) );
  OR2_X1 U11568 ( .A1(n11351), .A2(n11350), .ZN(n10398) );
  XNOR2_X2 U11569 ( .A(n10969), .B(n10685), .ZN(n10974) );
  NOR2_X2 U11570 ( .A1(n14005), .A2(n14086), .ZN(n14085) );
  NOR2_X2 U11571 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n17998), .ZN(n17985) );
  NOR2_X2 U11572 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n17977), .ZN(n17963) );
  NOR2_X2 U11573 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n18212), .ZN(n18183) );
  AND2_X1 U11574 ( .A1(n13784), .A2(n9831), .ZN(n9738) );
  AND2_X1 U11575 ( .A1(n13784), .A2(n9831), .ZN(n9739) );
  AND2_X4 U11576 ( .A1(n13784), .A2(n9831), .ZN(n11465) );
  INV_X2 U11577 ( .A(n11465), .ZN(n11475) );
  NAND2_X1 U11578 ( .A1(n16729), .A2(n11143), .ZN(n10196) );
  NAND2_X1 U11579 ( .A1(n9920), .A2(n10438), .ZN(n10440) );
  NAND2_X1 U11580 ( .A1(n13864), .A2(n9748), .ZN(n9920) );
  INV_X1 U11581 ( .A(n10517), .ZN(n10396) );
  INV_X1 U11582 ( .A(n10906), .ZN(n10909) );
  NAND2_X1 U11583 ( .A1(n10159), .A2(n16561), .ZN(n10226) );
  NAND2_X1 U11584 ( .A1(n13778), .A2(n14056), .ZN(n10597) );
  NAND2_X1 U11585 ( .A1(n21170), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15095) );
  INV_X1 U11586 ( .A(n10960), .ZN(n9953) );
  INV_X1 U11587 ( .A(n10231), .ZN(n9954) );
  OAI211_X1 U11588 ( .C1(n10957), .C2(n17130), .A(n10929), .B(n10928), .ZN(
        n10231) );
  NOR2_X1 U11589 ( .A1(n17006), .A2(n14753), .ZN(n10195) );
  NAND2_X1 U11590 ( .A1(n16649), .A2(n16646), .ZN(n10034) );
  NAND2_X1 U11591 ( .A1(n16673), .A2(n10002), .ZN(n16605) );
  AND2_X1 U11592 ( .A1(n9899), .A2(n10489), .ZN(n10002) );
  NOR2_X1 U11593 ( .A1(n22065), .A2(n16864), .ZN(n10346) );
  NAND2_X1 U11594 ( .A1(n10890), .A2(n17793), .ZN(n13626) );
  OAI21_X1 U11595 ( .B1(n12318), .B2(n12287), .A(n21334), .ZN(n12314) );
  AOI22_X1 U11596 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20611), .B1(
        n20543), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11026) );
  NOR2_X1 U11597 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n12111), .ZN(
        n12112) );
  CLKBUF_X1 U11598 ( .A(n12343), .Z(n12365) );
  AND2_X1 U11599 ( .A1(n12408), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12417) );
  NAND2_X1 U11600 ( .A1(n12288), .A2(n12293), .ZN(n12612) );
  NAND2_X1 U11601 ( .A1(n11052), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n10118) );
  NAND2_X1 U11602 ( .A1(n10903), .A2(n10907), .ZN(n10905) );
  NAND2_X1 U11603 ( .A1(n11256), .A2(n10908), .ZN(n10930) );
  AOI21_X1 U11604 ( .B1(n20002), .B2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n11984), .ZN(n11990) );
  OAI22_X1 U11605 ( .A1(n20157), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(
        n20011), .B2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11989) );
  NAND2_X1 U11606 ( .A1(n13977), .A2(n18680), .ZN(n11974) );
  INV_X1 U11607 ( .A(n19555), .ZN(n13977) );
  INV_X1 U11608 ( .A(n19543), .ZN(n11965) );
  NOR2_X1 U11609 ( .A1(n14931), .A2(n9883), .ZN(n14919) );
  NAND2_X1 U11610 ( .A1(n12755), .A2(n10277), .ZN(n14931) );
  NOR2_X1 U11611 ( .A1(n10651), .A2(n10278), .ZN(n10277) );
  NAND2_X1 U11612 ( .A1(n10652), .A2(n14943), .ZN(n10651) );
  INV_X1 U11613 ( .A(n10279), .ZN(n10278) );
  INV_X1 U11614 ( .A(n15149), .ZN(n10643) );
  NAND2_X1 U11615 ( .A1(n12568), .A2(n9989), .ZN(n12670) );
  NAND2_X1 U11616 ( .A1(n12548), .A2(n12566), .ZN(n9989) );
  INV_X1 U11617 ( .A(n13349), .ZN(n13384) );
  NAND2_X1 U11618 ( .A1(n9997), .A2(n10638), .ZN(n12607) );
  AOI21_X1 U11619 ( .B1(n9740), .B2(n12604), .A(n9802), .ZN(n10638) );
  NAND2_X1 U11620 ( .A1(n9992), .A2(n10178), .ZN(n15383) );
  NAND2_X1 U11621 ( .A1(n9994), .A2(n9993), .ZN(n9992) );
  AND2_X1 U11622 ( .A1(n9995), .A2(n10100), .ZN(n9993) );
  AND2_X1 U11623 ( .A1(n10442), .A2(n10099), .ZN(n10098) );
  AND2_X1 U11624 ( .A1(n10683), .A2(n9900), .ZN(n10442) );
  AND2_X1 U11625 ( .A1(n10683), .A2(n9996), .ZN(n9995) );
  NAND2_X1 U11626 ( .A1(n15545), .A2(n9893), .ZN(n9996) );
  OAI21_X1 U11627 ( .B1(n10443), .B2(n15545), .A(n15514), .ZN(n9994) );
  INV_X1 U11628 ( .A(n9924), .ZN(n9923) );
  NAND2_X1 U11629 ( .A1(n9922), .A2(n10438), .ZN(n9921) );
  OAI21_X1 U11630 ( .B1(n9925), .B2(n9748), .A(n9829), .ZN(n9924) );
  NAND2_X1 U11631 ( .A1(n10086), .A2(n10085), .ZN(n10091) );
  NOR2_X1 U11632 ( .A1(n10088), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10085) );
  OR2_X1 U11633 ( .A1(n13338), .A2(n15091), .ZN(n13885) );
  NAND2_X1 U11634 ( .A1(n12453), .A2(n12452), .ZN(n21470) );
  OR2_X1 U11635 ( .A1(n12446), .A2(n12697), .ZN(n12453) );
  NOR2_X1 U11636 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n21333), .ZN(n21336) );
  NAND2_X2 U11637 ( .A1(n10306), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12654) );
  INV_X1 U11638 ( .A(n12612), .ZN(n10306) );
  OAI211_X1 U11639 ( .C1(n11393), .C2(n10217), .A(n10621), .B(n9912), .ZN(
        n11362) );
  NAND2_X1 U11640 ( .A1(n9913), .A2(n11372), .ZN(n10621) );
  NAND2_X1 U11641 ( .A1(n9913), .A2(n10216), .ZN(n9912) );
  CLKBUF_X1 U11642 ( .A(n11157), .Z(n11158) );
  INV_X1 U11643 ( .A(n15999), .ZN(n10537) );
  INV_X1 U11644 ( .A(n16014), .ZN(n10538) );
  AND2_X1 U11645 ( .A1(n9858), .A2(n10582), .ZN(n10581) );
  INV_X1 U11646 ( .A(n16025), .ZN(n10582) );
  NAND2_X1 U11647 ( .A1(n10569), .A2(n10684), .ZN(n10568) );
  INV_X1 U11648 ( .A(n14327), .ZN(n10569) );
  INV_X1 U11649 ( .A(n14007), .ZN(n11571) );
  NAND2_X1 U11650 ( .A1(n9949), .A2(n10519), .ZN(n16750) );
  AND2_X1 U11651 ( .A1(n17060), .A2(n10520), .ZN(n9949) );
  NAND2_X2 U11652 ( .A1(n10023), .A2(n10396), .ZN(n11351) );
  AOI21_X1 U11653 ( .B1(n9973), .B2(n19195), .A(n9808), .ZN(n9972) );
  INV_X1 U11654 ( .A(n19195), .ZN(n9974) );
  NAND2_X1 U11655 ( .A1(n19204), .A2(n17306), .ZN(n17308) );
  NOR2_X1 U11656 ( .A1(n11953), .A2(n11952), .ZN(n11964) );
  NAND2_X1 U11657 ( .A1(n10291), .A2(n19185), .ZN(n17262) );
  OR2_X1 U11658 ( .A1(n19161), .A2(n9889), .ZN(n10291) );
  NAND2_X1 U11659 ( .A1(n10249), .A2(n14179), .ZN(n10248) );
  INV_X1 U11660 ( .A(n14175), .ZN(n10249) );
  AND2_X1 U11661 ( .A1(n12298), .A2(n12297), .ZN(n13349) );
  NOR2_X1 U11662 ( .A1(n13348), .A2(n13347), .ZN(n13934) );
  OR3_X1 U11663 ( .A1(n14789), .A2(n10658), .A3(n14823), .ZN(n10654) );
  INV_X1 U11664 ( .A(n14809), .ZN(n10658) );
  NAND2_X1 U11665 ( .A1(n10509), .A2(n10508), .ZN(n10507) );
  NOR2_X1 U11666 ( .A1(n10510), .A2(n14825), .ZN(n10508) );
  INV_X1 U11667 ( .A(n14841), .ZN(n10509) );
  NAND2_X1 U11668 ( .A1(n15402), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10268) );
  NAND2_X1 U11669 ( .A1(n9917), .A2(n15545), .ZN(n15423) );
  NAND2_X1 U11670 ( .A1(n12602), .A2(n9891), .ZN(n9917) );
  INV_X1 U11671 ( .A(n11743), .ZN(n11749) );
  NAND2_X1 U11672 ( .A1(n10940), .A2(n10939), .ZN(n10964) );
  AND2_X1 U11673 ( .A1(n9859), .A2(n9861), .ZN(n10146) );
  NAND2_X1 U11674 ( .A1(n10152), .A2(n10150), .ZN(n16398) );
  NAND2_X1 U11675 ( .A1(n14607), .A2(n10151), .ZN(n10150) );
  NAND2_X1 U11676 ( .A1(n16317), .A2(n10610), .ZN(n10152) );
  INV_X1 U11677 ( .A(n10614), .ZN(n10151) );
  NAND2_X1 U11678 ( .A1(n11764), .A2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11769) );
  INV_X1 U11679 ( .A(n10236), .ZN(n10235) );
  NOR2_X2 U11680 ( .A1(n15955), .A2(n14726), .ZN(n14725) );
  NAND2_X1 U11681 ( .A1(n10155), .A2(n9826), .ZN(n11456) );
  NOR2_X1 U11682 ( .A1(n14730), .A2(n22042), .ZN(n10523) );
  NAND2_X1 U11683 ( .A1(n10405), .A2(n9784), .ZN(n10047) );
  OAI21_X1 U11684 ( .B1(n9827), .B2(n10140), .A(n10401), .ZN(n10404) );
  NAND2_X1 U11685 ( .A1(n16054), .A2(n9868), .ZN(n16055) );
  OAI21_X1 U11686 ( .B1(n10560), .B2(n10559), .A(n10558), .ZN(n10557) );
  INV_X1 U11687 ( .A(n16588), .ZN(n10559) );
  NAND2_X1 U11688 ( .A1(n10233), .A2(n10560), .ZN(n16616) );
  NAND2_X1 U11689 ( .A1(n14762), .A2(n10561), .ZN(n10233) );
  INV_X1 U11690 ( .A(n16675), .ZN(n10556) );
  NAND2_X1 U11691 ( .A1(n9967), .A2(n10240), .ZN(n9962) );
  NAND2_X1 U11692 ( .A1(n17098), .A2(n17097), .ZN(n10519) );
  NAND4_X1 U11693 ( .A1(n11697), .A2(n10941), .A3(n10063), .A4(n13614), .ZN(
        n12048) );
  AND2_X1 U11694 ( .A1(n12047), .A2(n17793), .ZN(n12092) );
  AND4_X1 U11695 ( .A1(n14136), .A2(n17768), .A3(n12044), .A4(n12043), .ZN(
        n12045) );
  AOI21_X1 U11696 ( .B1(n13778), .B2(n10587), .A(n9835), .ZN(n10590) );
  NOR2_X1 U11697 ( .A1(n10596), .A2(n10588), .ZN(n10587) );
  AND2_X1 U11698 ( .A1(n11282), .A2(n21132), .ZN(n20941) );
  AND2_X1 U11699 ( .A1(n9981), .A2(n9979), .ZN(n17333) );
  AOI21_X1 U11700 ( .B1(n18957), .B2(n19185), .A(n9867), .ZN(n9979) );
  NAND2_X1 U11701 ( .A1(n18958), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n9981) );
  NOR2_X1 U11702 ( .A1(n19329), .A2(n10388), .ZN(n19281) );
  AND2_X1 U11703 ( .A1(n19444), .A2(n9886), .ZN(n10388) );
  NOR2_X1 U11704 ( .A1(n11981), .A2(n14027), .ZN(n14025) );
  AND2_X1 U11705 ( .A1(n20048), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n20179) );
  AOI21_X1 U11706 ( .B1(n10203), .B2(n16893), .A(n9743), .ZN(n10201) );
  INV_X1 U11707 ( .A(n19188), .ZN(n18802) );
  NAND2_X1 U11708 ( .A1(n20509), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n10036) );
  INV_X1 U11709 ( .A(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13100) );
  AOI21_X1 U11710 ( .B1(n12306), .B2(n12297), .A(n12305), .ZN(n12312) );
  NAND2_X1 U11711 ( .A1(n12310), .A2(n12309), .ZN(n12311) );
  NAND2_X1 U11712 ( .A1(n12667), .A2(n12296), .ZN(n13331) );
  INV_X1 U11713 ( .A(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12470) );
  AOI21_X1 U11714 ( .B1(n9719), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10320) );
  NAND2_X1 U11715 ( .A1(n10868), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n10311) );
  OAI22_X1 U11716 ( .A1(n9783), .A2(n18454), .B1(n18599), .B2(n22105), .ZN(
        n10353) );
  AND2_X1 U11717 ( .A1(n12649), .A2(n12648), .ZN(n12653) );
  INV_X1 U11718 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12121) );
  AND2_X1 U11719 ( .A1(n12565), .A2(n12564), .ZN(n12567) );
  INV_X2 U11720 ( .A(n12379), .ZN(n13279) );
  NAND2_X1 U11721 ( .A1(n10144), .A2(n12502), .ZN(n12568) );
  AND2_X1 U11722 ( .A1(n15468), .A2(n9932), .ZN(n10683) );
  OR2_X1 U11723 ( .A1(n12575), .A2(n12574), .ZN(n12584) );
  AND2_X1 U11724 ( .A1(n12671), .A2(n12295), .ZN(n12320) );
  INV_X1 U11725 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12406) );
  INV_X1 U11726 ( .A(n12041), .ZN(n11721) );
  INV_X1 U11727 ( .A(n10057), .ZN(n10056) );
  OAI21_X1 U11728 ( .B1(n10020), .B2(n10058), .A(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n10057) );
  NOR2_X1 U11729 ( .A1(n14012), .A2(n13977), .ZN(n11970) );
  NAND2_X1 U11730 ( .A1(n17296), .A2(n17295), .ZN(n17292) );
  NOR2_X1 U11731 ( .A1(n10504), .A2(n10506), .ZN(n10503) );
  INV_X1 U11732 ( .A(n15050), .ZN(n10506) );
  INV_X1 U11733 ( .A(n10505), .ZN(n10504) );
  OR2_X1 U11734 ( .A1(n13346), .A2(n13345), .ZN(n13348) );
  NAND2_X1 U11735 ( .A1(n12287), .A2(n21361), .ZN(n13935) );
  INV_X1 U11736 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12697) );
  OR2_X1 U11737 ( .A1(n14963), .A2(n14974), .ZN(n10653) );
  INV_X1 U11738 ( .A(n13264), .ZN(n13299) );
  AND2_X1 U11739 ( .A1(n13872), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13264) );
  AND2_X1 U11740 ( .A1(n12933), .A2(n9742), .ZN(n10279) );
  NOR2_X1 U11741 ( .A1(n12932), .A2(n14990), .ZN(n12933) );
  XNOR2_X1 U11742 ( .A(n12581), .B(n12572), .ZN(n12729) );
  INV_X1 U11743 ( .A(n14945), .ZN(n10512) );
  NOR2_X1 U11744 ( .A1(n10515), .A2(n10514), .ZN(n10513) );
  INV_X1 U11745 ( .A(n14960), .ZN(n10514) );
  INV_X1 U11746 ( .A(n14982), .ZN(n10515) );
  NOR2_X1 U11747 ( .A1(n10081), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10080) );
  INV_X1 U11748 ( .A(n12517), .ZN(n10081) );
  OAI21_X1 U11749 ( .B1(n15896), .B2(n10084), .A(n10082), .ZN(n10094) );
  NAND2_X1 U11750 ( .A1(n12623), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10084) );
  INV_X1 U11751 ( .A(n10083), .ZN(n10082) );
  OAI21_X1 U11752 ( .B1(n12517), .B2(n15569), .A(n10095), .ZN(n10083) );
  INV_X1 U11753 ( .A(n12690), .ZN(n10087) );
  NAND2_X1 U11754 ( .A1(n14793), .A2(n13937), .ZN(n13471) );
  OR2_X1 U11755 ( .A1(n12371), .A2(n12370), .ZN(n12534) );
  OAI211_X1 U11756 ( .C1(n12654), .C2(n12762), .A(n12400), .B(n12399), .ZN(
        n12401) );
  OAI21_X1 U11757 ( .B1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n12418), .A(
        n12417), .ZN(n12422) );
  INV_X1 U11758 ( .A(n17600), .ZN(n15877) );
  AND3_X2 U11759 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13873) );
  CLKBUF_X1 U11760 ( .A(n13851), .Z(n13865) );
  NAND2_X1 U11761 ( .A1(n13864), .A2(n21908), .ZN(n10437) );
  INV_X1 U11762 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n21636) );
  NAND2_X1 U11763 ( .A1(n10904), .A2(n10905), .ZN(n12088) );
  NOR2_X1 U11764 ( .A1(n10219), .A2(n9800), .ZN(n10218) );
  INV_X1 U11765 ( .A(n10635), .ZN(n10219) );
  NOR2_X1 U11766 ( .A1(n10632), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n10631) );
  AND2_X1 U11767 ( .A1(n11354), .A2(n10629), .ZN(n11380) );
  NOR2_X1 U11768 ( .A1(n10630), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n10629) );
  INV_X1 U11769 ( .A(n10631), .ZN(n10630) );
  NAND2_X1 U11770 ( .A1(n10209), .A2(n10208), .ZN(n11329) );
  NAND2_X1 U11771 ( .A1(n11288), .A2(n11292), .ZN(n10208) );
  NAND2_X1 U11772 ( .A1(n11479), .A2(n11462), .ZN(n10209) );
  NOR2_X1 U11773 ( .A1(n10322), .A2(n14730), .ZN(n10340) );
  NAND2_X1 U11774 ( .A1(n10920), .A2(n10547), .ZN(n12061) );
  AND2_X1 U11775 ( .A1(n20440), .A2(n20415), .ZN(n10547) );
  INV_X1 U11776 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n10414) );
  AND2_X1 U11777 ( .A1(n10415), .A2(n10414), .ZN(n10412) );
  INV_X1 U11778 ( .A(n10415), .ZN(n10410) );
  NOR2_X1 U11779 ( .A1(n10322), .A2(n13517), .ZN(n10343) );
  AND2_X1 U11780 ( .A1(n11785), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11155) );
  AND2_X1 U11781 ( .A1(n11781), .A2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11785) );
  NOR2_X1 U11782 ( .A1(n10322), .A2(n22170), .ZN(n10334) );
  NAND2_X1 U11783 ( .A1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n10430) );
  OR2_X1 U11784 ( .A1(n10430), .A2(n10429), .ZN(n10428) );
  NAND2_X1 U11785 ( .A1(n10546), .A2(n14764), .ZN(n10545) );
  INV_X1 U11786 ( .A(n14353), .ZN(n10546) );
  NAND2_X1 U11787 ( .A1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n10435) );
  NOR2_X1 U11788 ( .A1(n10922), .A2(n10898), .ZN(n10923) );
  NOR2_X1 U11789 ( .A1(n10031), .A2(n10030), .ZN(n10029) );
  NAND2_X1 U11790 ( .A1(n10028), .A2(n10234), .ZN(n10027) );
  INV_X1 U11791 ( .A(n15972), .ZN(n10536) );
  NOR2_X1 U11792 ( .A1(n10322), .A2(n12070), .ZN(n10337) );
  NAND2_X1 U11793 ( .A1(n9803), .A2(n10032), .ZN(n10033) );
  INV_X1 U11794 ( .A(n16601), .ZN(n10032) );
  NOR2_X1 U11795 ( .A1(n16587), .A2(n16600), .ZN(n11405) );
  AND3_X1 U11796 ( .A1(n11399), .A2(n16590), .A3(n9764), .ZN(n11404) );
  NAND2_X1 U11797 ( .A1(n10626), .A2(n9791), .ZN(n10625) );
  NAND2_X1 U11798 ( .A1(n16576), .A2(n16577), .ZN(n10627) );
  INV_X1 U11799 ( .A(n16050), .ZN(n10583) );
  INV_X1 U11800 ( .A(n11426), .ZN(n10401) );
  NAND2_X1 U11801 ( .A1(n10544), .A2(n10543), .ZN(n10542) );
  INV_X1 U11802 ( .A(n16116), .ZN(n10543) );
  INV_X1 U11803 ( .A(n10545), .ZN(n10544) );
  NOR2_X1 U11804 ( .A1(n10322), .A2(n16667), .ZN(n10331) );
  NOR2_X1 U11805 ( .A1(n10531), .A2(n10530), .ZN(n10529) );
  INV_X1 U11806 ( .A(n14347), .ZN(n10530) );
  AND2_X1 U11807 ( .A1(n16190), .A2(n11452), .ZN(n11411) );
  NOR2_X1 U11808 ( .A1(n10322), .A2(n17025), .ZN(n10328) );
  NOR2_X1 U11809 ( .A1(n16749), .A2(n11346), .ZN(n10198) );
  INV_X1 U11810 ( .A(n16194), .ZN(n10575) );
  AND4_X1 U11811 ( .A1(n11125), .A2(n11124), .A3(n11123), .A4(n11122), .ZN(
        n11138) );
  AND4_X1 U11812 ( .A1(n11130), .A2(n11129), .A3(n11128), .A4(n11127), .ZN(
        n11137) );
  AOI21_X1 U11813 ( .B1(n11347), .B2(n11346), .A(n16221), .ZN(n11349) );
  INV_X1 U11814 ( .A(n14251), .ZN(n11172) );
  OR2_X1 U11815 ( .A1(n11118), .A2(n11117), .ZN(n11510) );
  AND2_X1 U11816 ( .A1(n11335), .A2(n10189), .ZN(n10188) );
  NAND2_X1 U11817 ( .A1(n16263), .A2(n11452), .ZN(n10189) );
  NAND2_X1 U11818 ( .A1(n10188), .A2(n10190), .ZN(n10185) );
  MUX2_X1 U11819 ( .A(n11296), .B(P2_EBX_REG_4__SCAN_IN), .S(n11288), .Z(
        n11334) );
  INV_X1 U11820 ( .A(n14047), .ZN(n10596) );
  NAND2_X1 U11821 ( .A1(n10932), .A2(n10895), .ZN(n10934) );
  AND3_X1 U11822 ( .A1(n12040), .A2(n20415), .A3(n13819), .ZN(n9952) );
  NOR2_X1 U11823 ( .A1(n11002), .A2(n17146), .ZN(n10999) );
  NAND2_X1 U11824 ( .A1(n17146), .A2(n10183), .ZN(n10182) );
  AND3_X1 U11825 ( .A1(n10829), .A2(n10831), .A3(n14126), .ZN(n10361) );
  AND3_X1 U11826 ( .A1(n17146), .A2(n10991), .A3(n10183), .ZN(n20940) );
  NOR2_X1 U11827 ( .A1(n21096), .A2(n22183), .ZN(n20936) );
  AND2_X1 U11828 ( .A1(n10802), .A2(n10801), .ZN(n11276) );
  OR2_X1 U11829 ( .A1(n10800), .A2(n10799), .ZN(n10802) );
  NAND2_X1 U11830 ( .A1(n19995), .A2(n11831), .ZN(n9786) );
  AND2_X1 U11831 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11831) );
  INV_X1 U11832 ( .A(n19097), .ZN(n10482) );
  NAND2_X1 U11833 ( .A1(n17350), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17255) );
  OR2_X1 U11834 ( .A1(n17242), .A2(n17209), .ZN(n17247) );
  NOR2_X1 U11835 ( .A1(n19086), .A2(n19062), .ZN(n17260) );
  NAND2_X1 U11836 ( .A1(n17279), .A2(n17226), .ZN(n17242) );
  NAND2_X1 U11837 ( .A1(n19232), .A2(n17302), .ZN(n17303) );
  XNOR2_X1 U11838 ( .A(n17242), .B(n17287), .ZN(n17239) );
  NAND2_X1 U11839 ( .A1(n19233), .A2(n19234), .ZN(n19232) );
  AND2_X1 U11840 ( .A1(n11992), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11994) );
  AND2_X1 U11841 ( .A1(n11982), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13970) );
  AOI21_X1 U11842 ( .B1(n11990), .B2(n11989), .A(n11988), .ZN(n14178) );
  INV_X1 U11843 ( .A(n11975), .ZN(n10373) );
  NOR2_X1 U11844 ( .A1(n11974), .A2(n11965), .ZN(n10372) );
  NOR2_X1 U11845 ( .A1(n10354), .A2(n10351), .ZN(n10350) );
  AND2_X1 U11846 ( .A1(n17625), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n14788) );
  OR3_X1 U11847 ( .A1(n17629), .A2(n14785), .A3(n21146), .ZN(n15302) );
  NAND2_X1 U11848 ( .A1(n13268), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13307) );
  NAND2_X1 U11849 ( .A1(n14807), .A2(n14809), .ZN(n14808) );
  NAND2_X1 U11850 ( .A1(n13167), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n13212) );
  CLKBUF_X1 U11851 ( .A(n14850), .Z(n14851) );
  NOR2_X1 U11852 ( .A1(n13047), .A2(n15432), .ZN(n10054) );
  NAND2_X1 U11853 ( .A1(n10054), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n13113) );
  NAND2_X1 U11854 ( .A1(n13002), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n13047) );
  NAND2_X1 U11855 ( .A1(n12956), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n13001) );
  OR2_X1 U11856 ( .A1(n15010), .A2(n15009), .ZN(n15045) );
  AND3_X1 U11857 ( .A1(n12775), .A2(n12774), .A3(n12773), .ZN(n15149) );
  AND2_X1 U11858 ( .A1(n15168), .A2(n15157), .ZN(n10272) );
  NAND2_X1 U11859 ( .A1(n12706), .A2(n12705), .ZN(n13933) );
  NAND2_X1 U11860 ( .A1(n13933), .A2(n13932), .ZN(n14115) );
  OR2_X1 U11861 ( .A1(n17629), .A2(n13339), .ZN(n17609) );
  AND2_X1 U11862 ( .A1(n13477), .A2(n13476), .ZN(n14825) );
  NOR2_X1 U11863 ( .A1(n10107), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10106) );
  INV_X1 U11864 ( .A(n15392), .ZN(n10107) );
  INV_X1 U11865 ( .A(n15373), .ZN(n10110) );
  NOR2_X1 U11866 ( .A1(n15392), .A2(n9902), .ZN(n10109) );
  OR2_X1 U11867 ( .A1(n14840), .A2(n14841), .ZN(n14843) );
  NAND2_X1 U11868 ( .A1(n15423), .A2(n9756), .ZN(n10102) );
  NAND2_X1 U11869 ( .A1(n10501), .A2(n10500), .ZN(n10499) );
  NOR2_X1 U11870 ( .A1(n10502), .A2(n14881), .ZN(n10501) );
  INV_X1 U11871 ( .A(n14897), .ZN(n10500) );
  NAND2_X1 U11872 ( .A1(n15651), .A2(n13372), .ZN(n15635) );
  AOI21_X1 U11873 ( .B1(n10178), .B2(n15545), .A(n15545), .ZN(n10175) );
  AND2_X1 U11874 ( .A1(n10100), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10266) );
  AND2_X1 U11875 ( .A1(n15461), .A2(n10458), .ZN(n10457) );
  INV_X1 U11876 ( .A(n15647), .ZN(n10458) );
  AND2_X1 U11877 ( .A1(n15694), .A2(n13370), .ZN(n15670) );
  NOR2_X1 U11878 ( .A1(n14933), .A2(n14926), .ZN(n14928) );
  NAND2_X1 U11879 ( .A1(n15467), .A2(n10098), .ZN(n10097) );
  NAND2_X1 U11880 ( .A1(n9919), .A2(n9817), .ZN(n9918) );
  INV_X1 U11881 ( .A(n10443), .ZN(n9919) );
  NAND2_X1 U11882 ( .A1(n15467), .A2(n9932), .ZN(n15478) );
  NOR2_X1 U11883 ( .A1(n12597), .A2(n12596), .ZN(n12598) );
  XNOR2_X1 U11884 ( .A(n15554), .B(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15518) );
  NAND2_X1 U11885 ( .A1(n15835), .A2(n15834), .ZN(n9986) );
  AND2_X1 U11886 ( .A1(n15764), .A2(n15682), .ZN(n15816) );
  OR2_X1 U11887 ( .A1(n13312), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15837) );
  XNOR2_X1 U11888 ( .A(n12539), .B(n13828), .ZN(n13910) );
  OR2_X1 U11889 ( .A1(n15884), .A2(n21332), .ZN(n21469) );
  INV_X1 U11890 ( .A(n21584), .ZN(n21667) );
  NOR2_X1 U11891 ( .A1(n21477), .A2(n21476), .ZN(n21781) );
  NOR2_X1 U11892 ( .A1(n13896), .A2(n21701), .ZN(n21806) );
  INV_X1 U11893 ( .A(n21502), .ZN(n21728) );
  INV_X1 U11894 ( .A(n21523), .ZN(n21775) );
  AND2_X1 U11895 ( .A1(n21330), .A2(n15893), .ZN(n21776) );
  AND2_X1 U11896 ( .A1(n15884), .A2(n21332), .ZN(n21666) );
  NOR2_X2 U11897 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n21819) );
  INV_X1 U11898 ( .A(n21336), .ZN(n21476) );
  INV_X1 U11899 ( .A(n10304), .ZN(n10303) );
  NAND2_X1 U11900 ( .A1(n13321), .A2(n12664), .ZN(n12665) );
  NAND2_X1 U11901 ( .A1(n9834), .A2(n10301), .ZN(n10302) );
  INV_X1 U11902 ( .A(n9782), .ZN(n10301) );
  AND2_X1 U11903 ( .A1(n21871), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n17625) );
  NAND2_X1 U11904 ( .A1(n13502), .A2(n11439), .ZN(n11440) );
  NAND2_X1 U11905 ( .A1(n11429), .A2(n11436), .ZN(n11371) );
  NAND2_X1 U11906 ( .A1(n11362), .A2(n11306), .ZN(n11368) );
  OR2_X1 U11907 ( .A1(n11398), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n11402) );
  NAND2_X1 U11908 ( .A1(n11393), .A2(n11436), .ZN(n11382) );
  NAND2_X1 U11909 ( .A1(n11354), .A2(n10631), .ZN(n11384) );
  NOR2_X2 U11910 ( .A1(n11360), .A2(n11358), .ZN(n11354) );
  NOR2_X1 U11911 ( .A1(n17723), .A2(n10419), .ZN(n10418) );
  INV_X1 U11912 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10419) );
  INV_X1 U11913 ( .A(n20240), .ZN(n20260) );
  AND2_X1 U11914 ( .A1(n14270), .A2(n9866), .ZN(n10606) );
  OR2_X1 U11915 ( .A1(n11532), .A2(n11531), .ZN(n14335) );
  NOR2_X1 U11916 ( .A1(n13779), .A2(n21132), .ZN(n13799) );
  INV_X1 U11917 ( .A(n14607), .ZN(n16312) );
  NOR2_X1 U11918 ( .A1(n9781), .A2(n15986), .ZN(n15968) );
  INV_X1 U11919 ( .A(n16352), .ZN(n14456) );
  NOR2_X1 U11920 ( .A1(n14512), .A2(n16353), .ZN(n10605) );
  NOR2_X1 U11921 ( .A1(n20303), .A2(n13820), .ZN(n14677) );
  AND2_X1 U11922 ( .A1(n11732), .A2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11759) );
  OR2_X1 U11923 ( .A1(n16139), .A2(n11413), .ZN(n16646) );
  INV_X1 U11924 ( .A(n11755), .ZN(n11153) );
  NAND2_X1 U11925 ( .A1(n10528), .A2(n11159), .ZN(n10527) );
  NOR2_X1 U11926 ( .A1(n13499), .A2(n10050), .ZN(n10270) );
  INV_X1 U11927 ( .A(n13504), .ZN(n10215) );
  NAND2_X1 U11928 ( .A1(n10577), .A2(n15970), .ZN(n10576) );
  INV_X1 U11929 ( .A(n15986), .ZN(n10577) );
  NAND2_X1 U11930 ( .A1(n15952), .A2(n15953), .ZN(n15955) );
  NAND2_X1 U11931 ( .A1(n10066), .A2(n9746), .ZN(n11150) );
  AND2_X1 U11932 ( .A1(n11443), .A2(n10137), .ZN(n10131) );
  OAI211_X1 U11933 ( .C1(n16541), .C2(n10134), .A(n10133), .B(n10130), .ZN(
        n16534) );
  AOI21_X1 U11934 ( .B1(n10135), .B2(n10225), .A(n9916), .ZN(n10133) );
  INV_X1 U11935 ( .A(n10135), .ZN(n10134) );
  NAND2_X1 U11936 ( .A1(n16541), .A2(n10132), .ZN(n10130) );
  NAND2_X1 U11937 ( .A1(n10537), .A2(n15984), .ZN(n10534) );
  NOR2_X1 U11938 ( .A1(n16596), .A2(n16841), .ZN(n16580) );
  NAND2_X1 U11939 ( .A1(n10571), .A2(n16083), .ZN(n10570) );
  INV_X1 U11940 ( .A(n10573), .ZN(n10571) );
  AND2_X1 U11941 ( .A1(n11663), .A2(n11662), .ZN(n16119) );
  INV_X1 U11942 ( .A(n16663), .ZN(n10553) );
  AND3_X1 U11943 ( .A1(n11641), .A2(n11640), .A3(n11639), .ZN(n14327) );
  NOR2_X1 U11944 ( .A1(n16674), .A2(n16667), .ZN(n16666) );
  AND3_X1 U11945 ( .A1(n11589), .A2(n11588), .A3(n11587), .ZN(n14086) );
  AND3_X1 U11946 ( .A1(n11570), .A2(n11569), .A3(n11568), .ZN(n14007) );
  OR2_X1 U11947 ( .A1(n11411), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n16701) );
  NAND2_X1 U11948 ( .A1(n16717), .A2(n16714), .ZN(n16703) );
  OR2_X1 U11949 ( .A1(n11412), .A2(n17006), .ZN(n16715) );
  NAND2_X1 U11950 ( .A1(n16728), .A2(n11143), .ZN(n10122) );
  INV_X1 U11951 ( .A(n16729), .ZN(n10239) );
  NAND2_X1 U11952 ( .A1(n11314), .A2(n11313), .ZN(n10141) );
  NAND2_X1 U11953 ( .A1(n17067), .A2(n17065), .ZN(n11343) );
  NOR2_X1 U11954 ( .A1(n10905), .A2(n10876), .ZN(n17777) );
  CLKBUF_X1 U11955 ( .A(n16750), .Z(n16751) );
  INV_X1 U11956 ( .A(n10364), .ZN(n17059) );
  NOR2_X1 U11957 ( .A1(n10905), .A2(n10926), .ZN(n21118) );
  NAND2_X1 U11958 ( .A1(n17730), .A2(n11048), .ZN(n10067) );
  NAND2_X1 U11959 ( .A1(n10597), .A2(n10593), .ZN(n10592) );
  NOR2_X1 U11960 ( .A1(n21092), .A2(n20672), .ZN(n20713) );
  AND2_X1 U11961 ( .A1(n20672), .A2(n20673), .ZN(n20873) );
  AND2_X1 U11962 ( .A1(n20672), .A2(n21111), .ZN(n20779) );
  AND2_X1 U11963 ( .A1(n20370), .A2(n20369), .ZN(n20437) );
  INV_X1 U11964 ( .A(n20941), .ZN(n20811) );
  INV_X1 U11965 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n20945) );
  NAND2_X1 U11966 ( .A1(n10377), .A2(n17172), .ZN(n20023) );
  NOR2_X1 U11967 ( .A1(n17954), .A2(n17955), .ZN(n17953) );
  OR2_X1 U11968 ( .A1(n18044), .A2(n18227), .ZN(n10068) );
  NAND2_X1 U11969 ( .A1(n10068), .A2(n11806), .ZN(n18033) );
  NAND2_X1 U11970 ( .A1(n18670), .A2(n13981), .ZN(n18640) );
  AND2_X1 U11971 ( .A1(n18648), .A2(n10677), .ZN(n13981) );
  AND2_X1 U11972 ( .A1(n10259), .A2(P3_EAX_REG_16__SCAN_IN), .ZN(n10258) );
  NOR2_X1 U11973 ( .A1(n14164), .A2(n10288), .ZN(n10287) );
  INV_X1 U11974 ( .A(n14173), .ZN(n10288) );
  AOI22_X1 U11975 ( .A1(n17547), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n18585), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10459) );
  AOI22_X1 U11976 ( .A1(n18390), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_13__0__SCAN_IN), .B2(n18403), .ZN(n10008) );
  AOI21_X1 U11977 ( .B1(n20013), .B2(n10665), .A(n14010), .ZN(n14091) );
  OR2_X1 U11978 ( .A1(n18858), .A2(n19535), .ZN(n10665) );
  NAND2_X1 U11979 ( .A1(n19555), .A2(n18680), .ZN(n14110) );
  NOR2_X1 U11980 ( .A1(n10476), .A2(n10473), .ZN(n10472) );
  NAND2_X1 U11981 ( .A1(n10474), .A2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10473) );
  INV_X1 U11982 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n18134) );
  INV_X1 U11983 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n18145) );
  OR2_X1 U11984 ( .A1(n10079), .A2(n10484), .ZN(n19096) );
  NAND2_X1 U11985 ( .A1(n19198), .A2(n17309), .ZN(n17347) );
  OR2_X1 U11986 ( .A1(n17347), .A2(n17348), .ZN(n10013) );
  NAND2_X1 U11987 ( .A1(n19199), .A2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n19198) );
  AOI22_X1 U11988 ( .A1(n18628), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n9726), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11961) );
  AND2_X1 U11989 ( .A1(n17319), .A2(n10012), .ZN(n17325) );
  NOR2_X1 U11990 ( .A1(n17824), .A2(n17391), .ZN(n10009) );
  NOR2_X1 U11991 ( .A1(n17592), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n17632) );
  NOR2_X1 U11992 ( .A1(n17593), .A2(n17825), .ZN(n17633) );
  NAND2_X1 U11993 ( .A1(n18957), .A2(n17268), .ZN(n18958) );
  OAI21_X1 U11994 ( .B1(n17262), .B2(n10450), .A(n10448), .ZN(n10447) );
  NOR2_X1 U11995 ( .A1(n10449), .A2(n9806), .ZN(n10448) );
  OR2_X1 U11996 ( .A1(n19161), .A2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n19162) );
  NAND2_X1 U11997 ( .A1(n19990), .A2(n14025), .ZN(n20013) );
  AND3_X1 U11998 ( .A1(n11838), .A2(n11837), .A3(n11836), .ZN(n19532) );
  AND4_X1 U11999 ( .A1(n11818), .A2(n11817), .A3(n11816), .A4(n11815), .ZN(
        n11838) );
  NOR2_X1 U12000 ( .A1(n11835), .A2(n11834), .ZN(n11836) );
  CLKBUF_X2 U12001 ( .A(n13349), .Z(n13740) );
  INV_X1 U12002 ( .A(n14788), .ZN(n21146) );
  INV_X1 U12003 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n21905) );
  INV_X1 U12004 ( .A(n21233), .ZN(n21253) );
  AND2_X1 U12005 ( .A1(n13541), .A2(n13529), .ZN(n21259) );
  OR2_X1 U12006 ( .A1(n21212), .A2(n15092), .ZN(n21265) );
  NAND2_X1 U12007 ( .A1(n10657), .A2(n13304), .ZN(n10656) );
  XNOR2_X1 U12008 ( .A(n13307), .B(n13306), .ZN(n15361) );
  NAND2_X1 U12009 ( .A1(n14808), .A2(n14789), .ZN(n10280) );
  OR2_X1 U12010 ( .A1(n15389), .A2(n17671), .ZN(n9988) );
  INV_X1 U12011 ( .A(n17676), .ZN(n17661) );
  XNOR2_X1 U12012 ( .A(n13488), .B(n13487), .ZN(n14364) );
  XNOR2_X1 U12013 ( .A(n9990), .B(n12611), .ZN(n13495) );
  NAND2_X1 U12014 ( .A1(n9991), .A2(n12610), .ZN(n9990) );
  NAND2_X1 U12015 ( .A1(n12608), .A2(n12609), .ZN(n9991) );
  NOR3_X1 U12016 ( .A1(n15595), .A2(n15357), .A3(n10297), .ZN(n15587) );
  AND2_X1 U12017 ( .A1(n17681), .A2(n15367), .ZN(n10297) );
  NAND2_X1 U12018 ( .A1(n10445), .A2(n10444), .ZN(n15358) );
  NAND2_X1 U12019 ( .A1(n15356), .A2(n10100), .ZN(n10444) );
  OAI21_X1 U12020 ( .B1(n15386), .B2(n9903), .A(n15545), .ZN(n10445) );
  XNOR2_X1 U12021 ( .A(n10172), .B(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15607) );
  NAND2_X1 U12022 ( .A1(n10174), .A2(n10173), .ZN(n10172) );
  NAND2_X1 U12023 ( .A1(n15387), .A2(n10100), .ZN(n10174) );
  NAND2_X1 U12024 ( .A1(n15386), .A2(n15545), .ZN(n10173) );
  XNOR2_X1 U12025 ( .A(n9933), .B(n15617), .ZN(n15625) );
  NAND2_X1 U12026 ( .A1(n9935), .A2(n9934), .ZN(n9933) );
  OAI21_X1 U12027 ( .B1(n15415), .B2(n15391), .A(n15545), .ZN(n9934) );
  INV_X1 U12028 ( .A(n9936), .ZN(n9935) );
  OR2_X1 U12029 ( .A1(n13493), .A2(n13492), .ZN(n15839) );
  OR2_X1 U12030 ( .A1(n13493), .A2(n13342), .ZN(n15864) );
  CLKBUF_X1 U12031 ( .A(n15105), .Z(n21702) );
  NAND2_X1 U12032 ( .A1(n20348), .A2(n11698), .ZN(n20276) );
  INV_X1 U12034 ( .A(n9942), .ZN(n10971) );
  INV_X1 U12035 ( .A(n20276), .ZN(n20244) );
  NOR2_X1 U12036 ( .A1(n20250), .A2(n21006), .ZN(n16299) );
  NOR2_X2 U12037 ( .A1(n13629), .A2(n11708), .ZN(n20242) );
  AND2_X1 U12038 ( .A1(n10619), .A2(n10609), .ZN(n10608) );
  NAND2_X1 U12039 ( .A1(n10617), .A2(n16314), .ZN(n10609) );
  NAND2_X1 U12040 ( .A1(n16317), .A2(n10607), .ZN(n10612) );
  AND2_X1 U12041 ( .A1(n9776), .A2(n16319), .ZN(n10607) );
  INV_X1 U12042 ( .A(n16398), .ZN(n10620) );
  NAND2_X1 U12043 ( .A1(n16317), .A2(n16319), .ZN(n16318) );
  NOR2_X1 U12044 ( .A1(n16398), .A2(n9772), .ZN(n10149) );
  NAND2_X1 U12045 ( .A1(n9711), .A2(n16544), .ZN(n16795) );
  NAND2_X1 U12046 ( .A1(n16598), .A2(n20370), .ZN(n10125) );
  INV_X1 U12047 ( .A(n16597), .ZN(n10124) );
  INV_X1 U12048 ( .A(n16622), .ZN(n10207) );
  NAND2_X1 U12049 ( .A1(n9968), .A2(n11143), .ZN(n9965) );
  NAND2_X1 U12050 ( .A1(n9966), .A2(n11143), .ZN(n9964) );
  NAND2_X1 U12051 ( .A1(n13626), .A2(n11151), .ZN(n17736) );
  INV_X1 U12052 ( .A(n17736), .ZN(n20356) );
  XNOR2_X1 U12053 ( .A(n13522), .B(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14736) );
  INV_X1 U12054 ( .A(n12087), .ZN(n9951) );
  XNOR2_X1 U12055 ( .A(n10051), .B(n12019), .ZN(n14745) );
  INV_X1 U12056 ( .A(n10049), .ZN(n10048) );
  NAND2_X1 U12057 ( .A1(n16397), .A2(n17741), .ZN(n10408) );
  INV_X1 U12058 ( .A(n14734), .ZN(n10579) );
  OAI21_X1 U12059 ( .B1(n16310), .B2(n17745), .A(n14733), .ZN(n14734) );
  INV_X1 U12060 ( .A(n16543), .ZN(n9940) );
  NAND2_X1 U12061 ( .A1(n10159), .A2(n9863), .ZN(n10157) );
  INV_X1 U12062 ( .A(n16795), .ZN(n10169) );
  AND2_X1 U12063 ( .A1(n16797), .A2(n17741), .ZN(n10367) );
  XNOR2_X1 U12064 ( .A(n16603), .B(n16602), .ZN(n16878) );
  NAND2_X1 U12065 ( .A1(n16605), .A2(n10003), .ZN(n16879) );
  AOI21_X1 U12066 ( .B1(n14762), .B2(n10564), .A(n10563), .ZN(n16614) );
  OAI21_X1 U12067 ( .B1(n16678), .B2(n10556), .A(n16676), .ZN(n16665) );
  INV_X1 U12068 ( .A(n17745), .ZN(n17076) );
  INV_X1 U12069 ( .A(n17741), .ZN(n17105) );
  NAND2_X1 U12070 ( .A1(n12092), .A2(n12049), .ZN(n17745) );
  INV_X1 U12071 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n22183) );
  INV_X1 U12072 ( .A(n20952), .ZN(n20877) );
  INV_X1 U12073 ( .A(n20951), .ZN(n20894) );
  INV_X1 U12074 ( .A(n20966), .ZN(n20901) );
  INV_X1 U12075 ( .A(n20972), .ZN(n20906) );
  INV_X1 U12076 ( .A(n21922), .ZN(n20914) );
  INV_X1 U12077 ( .A(n20986), .ZN(n20921) );
  INV_X1 U12078 ( .A(n20994), .ZN(n20927) );
  AOI211_X1 U12079 ( .C1(n17954), .C2(n17955), .A(n17953), .B(n20051), .ZN(
        n10070) );
  NAND2_X1 U12080 ( .A1(n17959), .A2(n20125), .ZN(n10074) );
  OR2_X1 U12081 ( .A1(n17961), .A2(n20125), .ZN(n10073) );
  NOR2_X1 U12082 ( .A1(n18481), .A2(n10357), .ZN(n18445) );
  INV_X1 U12083 ( .A(n18765), .ZN(n19561) );
  AND2_X1 U12084 ( .A1(n18670), .A2(n18765), .ZN(n18667) );
  AOI21_X1 U12085 ( .B1(n18685), .B2(n10245), .A(n10244), .ZN(n10243) );
  INV_X1 U12086 ( .A(P3_EAX_REG_31__SCAN_IN), .ZN(n10244) );
  OR2_X1 U12087 ( .A1(n18724), .A2(P3_EAX_REG_30__SCAN_IN), .ZN(n10245) );
  NOR2_X1 U12088 ( .A1(n18700), .A2(n18679), .ZN(n10242) );
  NOR2_X1 U12089 ( .A1(n18716), .A2(n18873), .ZN(n18715) );
  NAND2_X1 U12090 ( .A1(n10383), .A2(n10381), .ZN(n10380) );
  INV_X1 U12091 ( .A(n17815), .ZN(n10383) );
  NAND2_X1 U12092 ( .A1(n10382), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10381) );
  NOR2_X2 U12093 ( .A1(n19194), .A2(n20044), .ZN(n19128) );
  OR2_X1 U12094 ( .A1(n19239), .A2(n18802), .ZN(n19150) );
  NAND3_X1 U12095 ( .A1(n17225), .A2(n17224), .A3(n17223), .ZN(n19188) );
  AND4_X1 U12096 ( .A1(n17218), .A2(n17217), .A3(n17216), .A4(n17215), .ZN(
        n17224) );
  AND4_X1 U12097 ( .A1(n17214), .A2(n17213), .A3(n17212), .A4(n17211), .ZN(
        n17225) );
  INV_X1 U12098 ( .A(n10391), .ZN(n10390) );
  OAI21_X1 U12099 ( .B1(n19293), .B2(n19287), .A(n19288), .ZN(n10391) );
  AOI211_X1 U12100 ( .C1(n19430), .C2(n19286), .A(n19285), .B(n10393), .ZN(
        n10392) );
  NOR2_X1 U12101 ( .A1(n20019), .A2(n19297), .ZN(n10393) );
  NOR2_X1 U12102 ( .A1(n19305), .A2(n19284), .ZN(n19296) );
  NOR2_X2 U12103 ( .A1(n19505), .A2(n18802), .ZN(n19455) );
  AND2_X1 U12104 ( .A1(n14190), .A2(n20179), .ZN(n19457) );
  NAND2_X1 U12105 ( .A1(n13344), .A2(n13890), .ZN(n12310) );
  NAND2_X1 U12106 ( .A1(n10117), .A2(n9710), .ZN(n11054) );
  NAND2_X1 U12107 ( .A1(n11052), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n10117) );
  NAND2_X1 U12108 ( .A1(n20543), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n9909) );
  NAND2_X1 U12109 ( .A1(n20784), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n10038) );
  NAND2_X1 U12110 ( .A1(n20449), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n10037) );
  NAND2_X1 U12111 ( .A1(n20718), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n10039) );
  AND2_X1 U12112 ( .A1(n10864), .A2(n10863), .ZN(n10872) );
  NAND2_X1 U12113 ( .A1(n14458), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n10860) );
  AOI21_X1 U12114 ( .B1(n14664), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10858) );
  INV_X1 U12115 ( .A(n13125), .ZN(n12332) );
  INV_X1 U12116 ( .A(n12508), .ZN(n10490) );
  OR2_X1 U12117 ( .A1(n12440), .A2(n12439), .ZN(n12503) );
  INV_X1 U12118 ( .A(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12488) );
  INV_X1 U12119 ( .A(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13119) );
  INV_X1 U12120 ( .A(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13121) );
  INV_X1 U12121 ( .A(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13135) );
  INV_X1 U12122 ( .A(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12936) );
  OR2_X1 U12123 ( .A1(n12342), .A2(n12187), .ZN(n12190) );
  XNOR2_X1 U12124 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n10796) );
  OAI21_X1 U12125 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n20157), .A(
        n11985), .ZN(n11986) );
  AND2_X1 U12126 ( .A1(n21729), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12634) );
  INV_X1 U12127 ( .A(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12800) );
  INV_X1 U12128 ( .A(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12260) );
  INV_X1 U12129 ( .A(n10653), .ZN(n10652) );
  CLKBUF_X1 U12130 ( .A(n13175), .Z(n13221) );
  BUF_X1 U12131 ( .A(n12379), .Z(n13250) );
  INV_X1 U12132 ( .A(n13379), .ZN(n10639) );
  NAND2_X1 U12133 ( .A1(n17663), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12588) );
  NAND2_X1 U12134 ( .A1(n10439), .A2(n10490), .ZN(n10438) );
  INV_X1 U12135 ( .A(n12468), .ZN(n10439) );
  OR2_X1 U12136 ( .A1(n12563), .A2(n12562), .ZN(n12573) );
  OR2_X1 U12137 ( .A1(n12483), .A2(n12482), .ZN(n12510) );
  INV_X1 U12139 ( .A(n13344), .ZN(n12668) );
  NOR2_X1 U12140 ( .A1(n13945), .A2(n10263), .ZN(n10262) );
  AND3_X1 U12141 ( .A1(n12330), .A2(n12329), .A3(n12328), .ZN(n12410) );
  INV_X1 U12142 ( .A(n12442), .ZN(n9927) );
  CLKBUF_X1 U12143 ( .A(n12318), .Z(n12319) );
  BUF_X1 U12144 ( .A(n12419), .Z(n12446) );
  NAND2_X1 U12145 ( .A1(n12612), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12626) );
  AOI21_X1 U12146 ( .B1(n21636), .B2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n12653), .ZN(n12662) );
  OAI211_X1 U12147 ( .C1(n12333), .C2(n13120), .A(n12239), .B(n12238), .ZN(
        n12240) );
  NOR2_X1 U12148 ( .A1(n10637), .A2(n10636), .ZN(n10635) );
  INV_X1 U12149 ( .A(n10678), .ZN(n10637) );
  CLKBUF_X1 U12150 ( .A(n14666), .Z(n14632) );
  NOR2_X1 U12151 ( .A1(n10417), .A2(n10416), .ZN(n10415) );
  NAND2_X1 U12152 ( .A1(n10518), .A2(n11036), .ZN(n10517) );
  NAND2_X1 U12153 ( .A1(n10312), .A2(n10311), .ZN(n10309) );
  AOI22_X1 U12154 ( .A1(n10865), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n10828), .ZN(n10712) );
  AND2_X1 U12155 ( .A1(n10403), .A2(n16813), .ZN(n10028) );
  AND4_X1 U12156 ( .A1(n11134), .A2(n11133), .A3(n11132), .A4(n11131), .ZN(
        n11136) );
  NAND2_X1 U12157 ( .A1(n10119), .A2(n16749), .ZN(n11350) );
  AND2_X1 U12158 ( .A1(n10120), .A2(n9872), .ZN(n10119) );
  INV_X1 U12159 ( .A(n20940), .ZN(n11091) );
  INV_X1 U12160 ( .A(n10866), .ZN(n14659) );
  AOI22_X1 U12161 ( .A1(n14458), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9720), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10818) );
  AND2_X1 U12162 ( .A1(n10749), .A2(n10748), .ZN(n10752) );
  OR2_X1 U12163 ( .A1(n11258), .A2(n10880), .ZN(n10749) );
  OR2_X1 U12164 ( .A1(n10800), .A2(n10801), .ZN(n10883) );
  INV_X1 U12165 ( .A(n17246), .ZN(n9973) );
  XNOR2_X1 U12166 ( .A(n17289), .B(n18811), .ZN(n17290) );
  INV_X1 U12167 ( .A(n11906), .ZN(n10354) );
  NAND2_X1 U12168 ( .A1(n11904), .A2(n10352), .ZN(n10351) );
  NOR2_X1 U12169 ( .A1(n11898), .A2(n10353), .ZN(n10352) );
  NOR2_X1 U12170 ( .A1(n15082), .A2(n15064), .ZN(n10505) );
  INV_X1 U12171 ( .A(n12261), .ZN(n13155) );
  INV_X1 U12172 ( .A(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13284) );
  NAND2_X1 U12173 ( .A1(n13075), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n12276) );
  OR2_X1 U12174 ( .A1(n10645), .A2(n10646), .ZN(n10644) );
  INV_X1 U12175 ( .A(n14867), .ZN(n10645) );
  NAND2_X1 U12176 ( .A1(n10648), .A2(n10647), .ZN(n10646) );
  INV_X1 U12177 ( .A(n10649), .ZN(n10648) );
  INV_X1 U12178 ( .A(n14880), .ZN(n10647) );
  NAND2_X1 U12179 ( .A1(n14891), .A2(n10650), .ZN(n10649) );
  INV_X1 U12180 ( .A(n14907), .ZN(n10650) );
  OR2_X1 U12181 ( .A1(n15009), .A2(n12931), .ZN(n14990) );
  INV_X1 U12182 ( .A(n15007), .ZN(n15042) );
  NOR2_X1 U12183 ( .A1(n14989), .A2(n15042), .ZN(n15043) );
  AND2_X1 U12184 ( .A1(n12682), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n13303) );
  INV_X1 U12185 ( .A(n15163), .ZN(n10274) );
  NOR2_X1 U12186 ( .A1(n12604), .A2(n10496), .ZN(n10495) );
  NAND2_X1 U12187 ( .A1(n13379), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10496) );
  INV_X1 U12188 ( .A(n14815), .ZN(n10510) );
  NOR2_X1 U12189 ( .A1(n10100), .A2(n12604), .ZN(n10498) );
  AND2_X1 U12190 ( .A1(n9902), .A2(n9891), .ZN(n10441) );
  INV_X1 U12191 ( .A(n14864), .ZN(n10502) );
  AND2_X1 U12192 ( .A1(n10179), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10178) );
  OR2_X1 U12193 ( .A1(n9755), .A2(n15545), .ZN(n10179) );
  NOR2_X1 U12194 ( .A1(n15481), .A2(n10113), .ZN(n10112) );
  INV_X1 U12195 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n10113) );
  OR2_X1 U12196 ( .A1(n15554), .A2(n12601), .ZN(n9932) );
  OR2_X1 U12197 ( .A1(n13338), .A2(n12668), .ZN(n13339) );
  AND2_X1 U12198 ( .A1(n12354), .A2(n12353), .ZN(n12582) );
  INV_X1 U12199 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13092) );
  INV_X1 U12200 ( .A(n12582), .ZN(n12579) );
  XNOR2_X1 U12201 ( .A(n12412), .B(n12410), .ZN(n12708) );
  OR2_X1 U12202 ( .A1(n12398), .A2(n12397), .ZN(n12528) );
  INV_X1 U12203 ( .A(n12403), .ZN(n9931) );
  INV_X1 U12204 ( .A(n12304), .ZN(n12294) );
  OR2_X1 U12205 ( .A1(n12342), .A2(n12212), .ZN(n12215) );
  AND4_X1 U12206 ( .A1(n12174), .A2(n12173), .A3(n12172), .A4(n12171), .ZN(
        n12179) );
  INV_X1 U12207 ( .A(n12307), .ZN(n12671) );
  AOI21_X1 U12208 ( .B1(n21907), .B2(n15878), .A(n15916), .ZN(n21333) );
  INV_X1 U12209 ( .A(n12626), .ZN(n12664) );
  AOI221_X1 U12210 ( .B1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n12662), 
        .C1(n15872), .C2(n12662), .A(n12661), .ZN(n13321) );
  NOR2_X1 U12211 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n21326), .ZN(
        n12661) );
  AOI21_X1 U12212 ( .B1(n10299), .B2(n12643), .A(n9828), .ZN(n10298) );
  AND2_X1 U12213 ( .A1(n11288), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n11448) );
  NOR2_X1 U12214 ( .A1(n11449), .A2(n11448), .ZN(n11710) );
  NOR2_X1 U12215 ( .A1(n11783), .A2(n11782), .ZN(n11781) );
  AND2_X1 U12216 ( .A1(n11446), .A2(n11436), .ZN(n13502) );
  AND2_X1 U12217 ( .A1(n11298), .A2(n11344), .ZN(n9915) );
  MUX2_X1 U12218 ( .A(n11294), .B(n11293), .S(n11288), .Z(n11318) );
  NAND2_X1 U12219 ( .A1(n9945), .A2(n9958), .ZN(n9944) );
  AND2_X1 U12220 ( .A1(n12063), .A2(n10927), .ZN(n9971) );
  CLKBUF_X1 U12221 ( .A(n14565), .Z(n14631) );
  CLKBUF_X1 U12222 ( .A(n14457), .Z(n14665) );
  INV_X1 U12223 ( .A(n14657), .ZN(n14650) );
  NAND2_X1 U12224 ( .A1(n16307), .A2(n10615), .ZN(n10614) );
  NOR2_X1 U12225 ( .A1(n10614), .A2(n10611), .ZN(n10610) );
  INV_X1 U12226 ( .A(n16319), .ZN(n10611) );
  XNOR2_X1 U12227 ( .A(n16337), .B(n14576), .ZN(n16322) );
  AND2_X1 U12228 ( .A1(n14380), .A2(n10599), .ZN(n10598) );
  INV_X1 U12229 ( .A(n16372), .ZN(n10599) );
  AND2_X1 U12230 ( .A1(n13799), .A2(n9736), .ZN(n14599) );
  INV_X1 U12231 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n11782) );
  NAND2_X1 U12232 ( .A1(n10425), .A2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11783) );
  NOR2_X1 U12233 ( .A1(n11771), .A2(n16017), .ZN(n10425) );
  NOR2_X1 U12234 ( .A1(n11769), .A2(n11768), .ZN(n11767) );
  INV_X1 U12235 ( .A(n16039), .ZN(n10539) );
  AOI21_X1 U12236 ( .B1(n10555), .B2(n10552), .A(n10551), .ZN(n10550) );
  INV_X1 U12237 ( .A(n16654), .ZN(n10551) );
  NAND2_X1 U12238 ( .A1(n12097), .A2(n12096), .ZN(n10237) );
  NAND2_X1 U12239 ( .A1(n10552), .A2(n16655), .ZN(n10548) );
  INV_X1 U12240 ( .A(n12096), .ZN(n10238) );
  AND2_X1 U12241 ( .A1(n11443), .A2(n16524), .ZN(n10132) );
  NOR2_X1 U12242 ( .A1(n10136), .A2(n16524), .ZN(n10135) );
  INV_X1 U12243 ( .A(n16523), .ZN(n10136) );
  NOR2_X1 U12244 ( .A1(n16523), .A2(n10137), .ZN(n9916) );
  AND2_X1 U12245 ( .A1(n11148), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10522) );
  NOR2_X1 U12246 ( .A1(n16849), .A2(n11147), .ZN(n11148) );
  INV_X1 U12247 ( .A(n10033), .ZN(n11425) );
  INV_X1 U12248 ( .A(n16587), .ZN(n10558) );
  NAND2_X1 U12249 ( .A1(n11664), .A2(n10574), .ZN(n10573) );
  INV_X1 U12250 ( .A(n16100), .ZN(n10574) );
  NAND2_X1 U12251 ( .A1(n16612), .A2(n10563), .ZN(n10560) );
  NOR2_X1 U12252 ( .A1(n12101), .A2(n10562), .ZN(n10561) );
  INV_X1 U12253 ( .A(n10564), .ZN(n10562) );
  NAND2_X1 U12254 ( .A1(n11192), .A2(n10532), .ZN(n10531) );
  INV_X1 U12255 ( .A(n16154), .ZN(n10532) );
  AND2_X1 U12256 ( .A1(n11395), .A2(n16955), .ZN(n12098) );
  NAND2_X1 U12257 ( .A1(n16750), .A2(n9947), .ZN(n10062) );
  NAND2_X1 U12258 ( .A1(n9948), .A2(n11141), .ZN(n9947) );
  INV_X1 U12259 ( .A(n14217), .ZN(n10528) );
  NAND2_X1 U12260 ( .A1(n10118), .A2(n9822), .ZN(n11084) );
  AND2_X1 U12261 ( .A1(n11467), .A2(n9969), .ZN(n12029) );
  NAND2_X1 U12262 ( .A1(n11312), .A2(n17073), .ZN(n17060) );
  NAND2_X1 U12263 ( .A1(n11346), .A2(n11340), .ZN(n10022) );
  INV_X1 U12264 ( .A(n9878), .ZN(n10019) );
  NAND2_X1 U12265 ( .A1(n10020), .A2(n10025), .ZN(n10024) );
  INV_X1 U12266 ( .A(n11340), .ZN(n10025) );
  NAND2_X1 U12267 ( .A1(n11346), .A2(n9878), .ZN(n10026) );
  OR2_X1 U12268 ( .A1(n11079), .A2(n11078), .ZN(n11505) );
  NAND2_X1 U12269 ( .A1(n10187), .A2(n16263), .ZN(n17084) );
  NAND2_X1 U12270 ( .A1(n11316), .A2(n11300), .ZN(n10187) );
  INV_X1 U12271 ( .A(n11013), .ZN(n10210) );
  NOR2_X1 U12272 ( .A1(n11021), .A2(n10212), .ZN(n10211) );
  NOR2_X1 U12273 ( .A1(n10906), .A2(n9969), .ZN(n10931) );
  NOR2_X1 U12274 ( .A1(n10709), .A2(n10708), .ZN(n11464) );
  OR2_X1 U12275 ( .A1(n10699), .A2(n10698), .ZN(n10709) );
  NAND2_X1 U12276 ( .A1(n13780), .A2(n21106), .ZN(n14059) );
  AND2_X1 U12277 ( .A1(n14599), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n14047) );
  AND2_X1 U12278 ( .A1(n14599), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n14062) );
  INV_X1 U12279 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n21982) );
  INV_X1 U12280 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20837) );
  AOI21_X1 U12281 ( .B1(n14664), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10725) );
  NAND2_X1 U12282 ( .A1(n14458), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n10718) );
  NAND2_X1 U12283 ( .A1(n9908), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9907) );
  NAND2_X1 U12284 ( .A1(n9906), .A2(n14126), .ZN(n9905) );
  NAND2_X1 U12285 ( .A1(n10913), .A2(n14126), .ZN(n10843) );
  NAND2_X1 U12286 ( .A1(n10910), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10842) );
  AND2_X1 U12287 ( .A1(n10851), .A2(n10850), .ZN(n10855) );
  NAND2_X1 U12288 ( .A1(n9714), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n10851) );
  AND2_X1 U12289 ( .A1(n10845), .A2(n10844), .ZN(n10849) );
  NAND2_X1 U12290 ( .A1(n14458), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n10844) );
  NAND2_X1 U12291 ( .A1(n10883), .A2(n10882), .ZN(n11272) );
  INV_X1 U12292 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n17770) );
  NAND2_X1 U12293 ( .A1(n19539), .A2(n11970), .ZN(n11968) );
  NOR2_X1 U12294 ( .A1(n10375), .A2(n14188), .ZN(n10374) );
  INV_X1 U12295 ( .A(n10376), .ZN(n10375) );
  NAND2_X1 U12296 ( .A1(n10247), .A2(n14179), .ZN(n17929) );
  INV_X1 U12297 ( .A(n11981), .ZN(n10247) );
  NOR2_X1 U12298 ( .A1(n18108), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n18094) );
  NOR2_X1 U12299 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11824) );
  NAND2_X1 U12300 ( .A1(n19995), .A2(n11830), .ZN(n18466) );
  NOR2_X1 U12301 ( .A1(n17459), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11830) );
  AND2_X1 U12302 ( .A1(n20157), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11823) );
  AND2_X1 U12303 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11819) );
  AND2_X1 U12304 ( .A1(n20146), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11812) );
  INV_X1 U12306 ( .A(n18998), .ZN(n10474) );
  NOR2_X1 U12307 ( .A1(n19444), .A2(n20171), .ZN(n10376) );
  NOR2_X1 U12308 ( .A1(n17261), .A2(n10450), .ZN(n10449) );
  NAND2_X1 U12309 ( .A1(n17255), .A2(n17254), .ZN(n9978) );
  NAND2_X1 U12310 ( .A1(n9885), .A2(n10290), .ZN(n10289) );
  AND2_X1 U12311 ( .A1(n19138), .A2(n10463), .ZN(n10462) );
  XNOR2_X1 U12312 ( .A(n17290), .B(n19511), .ZN(n19234) );
  NOR2_X1 U12313 ( .A1(n11979), .A2(n11978), .ZN(n14016) );
  OR2_X1 U12314 ( .A1(n11977), .A2(n11976), .ZN(n11978) );
  OR3_X1 U12315 ( .A1(n14026), .A2(n14189), .A3(n13978), .ZN(n14176) );
  NOR2_X1 U12316 ( .A1(n19997), .A2(n20146), .ZN(n17576) );
  NOR2_X1 U12317 ( .A1(n20171), .A2(n18858), .ZN(n18856) );
  NAND2_X1 U12318 ( .A1(n15911), .A2(n21908), .ZN(n13312) );
  OR2_X1 U12319 ( .A1(n15459), .A2(n13302), .ZN(n12981) );
  AND2_X1 U12320 ( .A1(n13435), .A2(n13434), .ZN(n15050) );
  AND2_X1 U12321 ( .A1(n13431), .A2(n10503), .ZN(n15052) );
  OR2_X1 U12322 ( .A1(n15291), .A2(n13860), .ZN(n14748) );
  INV_X1 U12323 ( .A(n10654), .ZN(n10657) );
  AOI21_X1 U12324 ( .B1(n15364), .B2(n13267), .A(n13266), .ZN(n14809) );
  AND2_X1 U12325 ( .A1(n13166), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n13167) );
  NOR2_X1 U12326 ( .A1(n13113), .A2(n15416), .ZN(n13114) );
  NAND2_X1 U12327 ( .A1(n13114), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n13165) );
  CLKBUF_X1 U12328 ( .A(n14905), .Z(n14906) );
  NOR2_X1 U12329 ( .A1(n13001), .A2(n10055), .ZN(n13002) );
  OR2_X1 U12330 ( .A1(n15447), .A2(n13302), .ZN(n13027) );
  CLKBUF_X1 U12331 ( .A(n14919), .Z(n14920) );
  AND2_X1 U12332 ( .A1(n12955), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n12956) );
  AND2_X1 U12333 ( .A1(n12818), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12796) );
  NAND2_X1 U12334 ( .A1(n12796), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12954) );
  NOR2_X1 U12335 ( .A1(n12841), .A2(n12840), .ZN(n12818) );
  NAND2_X1 U12336 ( .A1(n10053), .A2(n10052), .ZN(n12841) );
  NOR2_X1 U12337 ( .A1(n15049), .A2(n15069), .ZN(n10052) );
  INV_X1 U12338 ( .A(n12911), .ZN(n10053) );
  INV_X1 U12339 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n15049) );
  INV_X1 U12340 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n15069) );
  NAND2_X1 U12341 ( .A1(n12907), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n12911) );
  NOR2_X1 U12342 ( .A1(n12795), .A2(n15550), .ZN(n12907) );
  OR2_X1 U12343 ( .A1(n12776), .A2(n15557), .ZN(n12795) );
  NAND2_X1 U12344 ( .A1(n12771), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12776) );
  NAND2_X1 U12345 ( .A1(n9884), .A2(n10643), .ZN(n10641) );
  NAND2_X1 U12346 ( .A1(n12686), .A2(n9823), .ZN(n12730) );
  AND2_X1 U12347 ( .A1(n12686), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12724) );
  INV_X1 U12348 ( .A(n12678), .ZN(n12679) );
  NOR2_X1 U12349 ( .A1(n12691), .A2(n21254), .ZN(n12692) );
  OR2_X1 U12350 ( .A1(n13836), .A2(n13837), .ZN(n13838) );
  INV_X1 U12351 ( .A(n13937), .ZN(n14786) );
  OR2_X1 U12352 ( .A1(n14814), .A2(n14793), .ZN(n13484) );
  NAND2_X1 U12353 ( .A1(n14814), .A2(n14794), .ZN(n13483) );
  NAND2_X1 U12354 ( .A1(n15369), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12609) );
  INV_X1 U12355 ( .A(n12607), .ZN(n15369) );
  AND2_X1 U12356 ( .A1(n13464), .A2(n13463), .ZN(n14881) );
  NAND2_X1 U12357 ( .A1(n14994), .A2(n9865), .ZN(n14933) );
  INV_X1 U12358 ( .A(n14935), .ZN(n10511) );
  NAND2_X1 U12359 ( .A1(n14994), .A2(n9855), .ZN(n14947) );
  AND2_X1 U12360 ( .A1(n15714), .A2(n15703), .ZN(n15706) );
  AND2_X1 U12361 ( .A1(n10114), .A2(n10111), .ZN(n10115) );
  INV_X1 U12362 ( .A(n15481), .ZN(n10111) );
  OR2_X1 U12363 ( .A1(n15014), .A2(n15015), .ZN(n15017) );
  AND2_X1 U12364 ( .A1(n13444), .A2(n13443), .ZN(n14995) );
  NAND2_X1 U12365 ( .A1(n13364), .A2(n13359), .ZN(n15764) );
  NAND2_X1 U12366 ( .A1(n13431), .A2(n13430), .ZN(n15084) );
  AND2_X1 U12367 ( .A1(n13365), .A2(n15814), .ZN(n15840) );
  CLKBUF_X1 U12368 ( .A(n15514), .Z(n15542) );
  OR2_X1 U12369 ( .A1(n15564), .A2(n15561), .ZN(n9983) );
  NAND2_X1 U12370 ( .A1(n15564), .A2(n15561), .ZN(n9985) );
  NAND2_X1 U12371 ( .A1(n13409), .A2(n10674), .ZN(n15172) );
  NAND2_X1 U12372 ( .A1(n10096), .A2(n10094), .ZN(n10093) );
  OR2_X1 U12373 ( .A1(n13493), .A2(n15908), .ZN(n15682) );
  OR2_X1 U12374 ( .A1(n13364), .A2(n17697), .ZN(n10292) );
  NAND2_X1 U12375 ( .A1(n13825), .A2(n13826), .ZN(n10269) );
  INV_X1 U12376 ( .A(n10292), .ZN(n15766) );
  AND2_X1 U12377 ( .A1(n13364), .A2(n13934), .ZN(n15851) );
  OR2_X1 U12378 ( .A1(n15764), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10293) );
  CLKBUF_X1 U12379 ( .A(n12708), .Z(n12709) );
  NOR2_X1 U12380 ( .A1(n12424), .A2(n12423), .ZN(n12425) );
  NAND2_X1 U12381 ( .A1(n12426), .A2(n12422), .ZN(n10104) );
  OR2_X1 U12382 ( .A1(n15896), .A2(n21330), .ZN(n21584) );
  INV_X1 U12383 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13945) );
  AND2_X1 U12385 ( .A1(n13893), .A2(n13892), .ZN(n17600) );
  NAND2_X1 U12386 ( .A1(n21331), .A2(n15896), .ZN(n21436) );
  OR2_X1 U12387 ( .A1(n21440), .A2(n21815), .ZN(n21444) );
  INV_X1 U12388 ( .A(n21370), .ZN(n21371) );
  OR3_X1 U12389 ( .A1(n21704), .A2(P1_STATE2_REG_0__SCAN_IN), .A3(n21333), 
        .ZN(n21374) );
  NAND2_X1 U12390 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n15878) );
  XNOR2_X1 U12391 ( .A(n15923), .B(P1_STATE_REG_1__SCAN_IN), .ZN(n13322) );
  CLKBUF_X1 U12392 ( .A(n11256), .Z(n11257) );
  AND2_X1 U12393 ( .A1(n12020), .A2(n11278), .ZN(n17774) );
  AND2_X1 U12394 ( .A1(n12090), .A2(n12089), .ZN(n17776) );
  AND2_X1 U12395 ( .A1(n11693), .A2(n11692), .ZN(n14726) );
  NAND2_X1 U12396 ( .A1(n10223), .A2(n10222), .ZN(n11446) );
  NOR2_X1 U12397 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(P2_EBX_REG_25__SCAN_IN), 
        .ZN(n10222) );
  INV_X1 U12398 ( .A(n11438), .ZN(n10223) );
  NAND2_X1 U12399 ( .A1(n11437), .A2(n11444), .ZN(n11449) );
  INV_X1 U12400 ( .A(n13502), .ZN(n11437) );
  INV_X1 U12401 ( .A(n16609), .ZN(n10431) );
  NAND2_X1 U12402 ( .A1(n10434), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n11740) );
  INV_X1 U12403 ( .A(n11737), .ZN(n10434) );
  NOR2_X1 U12404 ( .A1(n11737), .A2(n10435), .ZN(n11756) );
  NOR2_X1 U12405 ( .A1(n12036), .A2(n11722), .ZN(n13632) );
  INV_X1 U12406 ( .A(n20269), .ZN(n20256) );
  NOR2_X1 U12407 ( .A1(n20233), .A2(n21006), .ZN(n16174) );
  NAND2_X1 U12408 ( .A1(n13629), .A2(n11719), .ZN(n20269) );
  NAND2_X1 U12409 ( .A1(n11251), .A2(n10339), .ZN(n11254) );
  NOR2_X1 U12410 ( .A1(n10341), .A2(n10340), .ZN(n10339) );
  INV_X1 U12411 ( .A(n11252), .ZN(n10341) );
  AND2_X1 U12412 ( .A1(n11240), .A2(n11239), .ZN(n15999) );
  AND2_X1 U12413 ( .A1(n11214), .A2(n11213), .ZN(n16116) );
  INV_X1 U12414 ( .A(n10936), .ZN(n13776) );
  NAND2_X1 U12415 ( .A1(n13512), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10323) );
  CLKBUF_X1 U12416 ( .A(n16322), .Z(n16323) );
  CLKBUF_X1 U12417 ( .A(n16356), .Z(n16357) );
  INV_X1 U12418 ( .A(n11476), .ZN(n13818) );
  NAND2_X1 U12419 ( .A1(n16281), .A2(n16280), .ZN(n16282) );
  INV_X1 U12420 ( .A(n13614), .ZN(n14134) );
  NAND2_X1 U12421 ( .A1(n10410), .A2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n10409) );
  NAND2_X1 U12422 ( .A1(n11155), .A2(n10412), .ZN(n10411) );
  OR2_X1 U12423 ( .A1(n11155), .A2(n10414), .ZN(n10413) );
  INV_X1 U12424 ( .A(n11243), .ZN(n13510) );
  NAND2_X1 U12425 ( .A1(n11700), .A2(n10342), .ZN(n11702) );
  NOR2_X1 U12426 ( .A1(n10344), .A2(n10343), .ZN(n10342) );
  INV_X1 U12427 ( .A(n11701), .ZN(n10344) );
  NAND2_X1 U12428 ( .A1(n11703), .A2(n11702), .ZN(n13514) );
  INV_X1 U12429 ( .A(n10425), .ZN(n11776) );
  NOR2_X1 U12430 ( .A1(n10335), .A2(n10334), .ZN(n10333) );
  INV_X1 U12431 ( .A(n11233), .ZN(n10335) );
  INV_X1 U12432 ( .A(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n11768) );
  NAND2_X1 U12433 ( .A1(n10427), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n10426) );
  INV_X1 U12434 ( .A(n10428), .ZN(n10427) );
  NAND2_X1 U12435 ( .A1(n13512), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n10326) );
  AND2_X1 U12436 ( .A1(n9892), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10488) );
  INV_X1 U12437 ( .A(n10307), .ZN(n9966) );
  NOR2_X1 U12438 ( .A1(n12103), .A2(n16955), .ZN(n10489) );
  NAND2_X1 U12439 ( .A1(n11759), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11758) );
  NAND2_X1 U12440 ( .A1(n13512), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10325) );
  NAND2_X1 U12441 ( .A1(n10433), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10432) );
  INV_X1 U12442 ( .A(n10435), .ZN(n10433) );
  AND2_X1 U12443 ( .A1(n11208), .A2(n11207), .ZN(n14353) );
  NAND2_X1 U12444 ( .A1(n11749), .A2(n9820), .ZN(n11755) );
  AND2_X1 U12445 ( .A1(n11749), .A2(n9762), .ZN(n11753) );
  NAND2_X1 U12446 ( .A1(n13512), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10324) );
  AND2_X1 U12447 ( .A1(n11749), .A2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11751) );
  NAND2_X1 U12448 ( .A1(n11749), .A2(n9749), .ZN(n11748) );
  AND2_X1 U12449 ( .A1(n10422), .A2(n10421), .ZN(n11745) );
  NOR2_X1 U12450 ( .A1(n11746), .A2(n10423), .ZN(n10422) );
  NOR2_X1 U12451 ( .A1(n17737), .A2(n17723), .ZN(n10421) );
  INV_X1 U12452 ( .A(n11746), .ZN(n10424) );
  NAND2_X1 U12453 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n11746) );
  OAI21_X1 U12454 ( .B1(n16523), .B2(n10050), .A(n13496), .ZN(n10049) );
  INV_X1 U12455 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14730) );
  AND2_X1 U12456 ( .A1(n10625), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n10623) );
  NAND2_X1 U12457 ( .A1(n10140), .A2(n10401), .ZN(n10138) );
  INV_X1 U12458 ( .A(n16561), .ZN(n10158) );
  NOR2_X1 U12459 ( .A1(n11455), .A2(n11441), .ZN(n16543) );
  NAND2_X1 U12460 ( .A1(n11241), .A2(n10336), .ZN(n15984) );
  NOR2_X1 U12461 ( .A1(n10338), .A2(n10337), .ZN(n10336) );
  INV_X1 U12462 ( .A(n11242), .ZN(n10338) );
  AND2_X1 U12463 ( .A1(n11683), .A2(n11682), .ZN(n15997) );
  AND2_X1 U12464 ( .A1(n10581), .A2(n16010), .ZN(n10580) );
  INV_X1 U12465 ( .A(n10140), .ZN(n10230) );
  NAND2_X1 U12466 ( .A1(n16756), .A2(n11361), .ZN(n10229) );
  AND2_X1 U12467 ( .A1(n11678), .A2(n11677), .ZN(n16025) );
  AND2_X1 U12468 ( .A1(n11674), .A2(n10581), .ZN(n16027) );
  NAND2_X1 U12469 ( .A1(n11674), .A2(n9858), .ZN(n16048) );
  NAND2_X1 U12470 ( .A1(n11407), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n16591) );
  CLKBUF_X1 U12471 ( .A(n16056), .Z(n16057) );
  AND2_X1 U12472 ( .A1(n11423), .A2(n16860), .ZN(n16600) );
  AND2_X1 U12473 ( .A1(n11424), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n16601) );
  NAND2_X1 U12474 ( .A1(n10541), .A2(n11218), .ZN(n10540) );
  INV_X1 U12475 ( .A(n10542), .ZN(n10541) );
  AND2_X1 U12476 ( .A1(n16624), .A2(n12100), .ZN(n10564) );
  INV_X1 U12477 ( .A(n16625), .ZN(n10563) );
  INV_X1 U12478 ( .A(n14766), .ZN(n10572) );
  OR2_X1 U12479 ( .A1(n16978), .A2(n14755), .ZN(n16926) );
  NAND2_X1 U12480 ( .A1(n10566), .A2(n14360), .ZN(n10565) );
  INV_X1 U12481 ( .A(n10568), .ZN(n10566) );
  AND2_X1 U12482 ( .A1(n11202), .A2(n11201), .ZN(n14317) );
  NAND2_X1 U12483 ( .A1(n11197), .A2(n10330), .ZN(n14347) );
  NOR2_X1 U12484 ( .A1(n10332), .A2(n10331), .ZN(n10330) );
  INV_X1 U12485 ( .A(n11198), .ZN(n10332) );
  INV_X1 U12486 ( .A(n14278), .ZN(n11187) );
  INV_X1 U12487 ( .A(n14275), .ZN(n11188) );
  NOR2_X1 U12488 ( .A1(n17023), .A2(n12081), .ZN(n16989) );
  INV_X1 U12489 ( .A(n13920), .ZN(n11553) );
  NAND2_X1 U12490 ( .A1(n11173), .A2(n10327), .ZN(n16196) );
  NOR2_X1 U12491 ( .A1(n10329), .A2(n10328), .ZN(n10327) );
  INV_X1 U12492 ( .A(n11174), .ZN(n10329) );
  NAND2_X1 U12493 ( .A1(n10199), .A2(n17025), .ZN(n11142) );
  NAND2_X1 U12494 ( .A1(n10198), .A2(n10197), .ZN(n10199) );
  NOR2_X1 U12495 ( .A1(n11351), .A2(n11300), .ZN(n10197) );
  AND3_X1 U12496 ( .A1(n11535), .A2(n11534), .A3(n11533), .ZN(n16194) );
  XNOR2_X1 U12497 ( .A(n11141), .B(n11300), .ZN(n16739) );
  AND2_X1 U12498 ( .A1(n10185), .A2(n11339), .ZN(n10184) );
  INV_X1 U12499 ( .A(n20355), .ZN(n20217) );
  INV_X1 U12500 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n17130) );
  MUX2_X1 U12501 ( .A(n16103), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .S(
        P2_STATE2_REG_0__SCAN_IN), .Z(n20250) );
  INV_X1 U12502 ( .A(n20250), .ZN(n20233) );
  CLKBUF_X1 U12503 ( .A(n14127), .Z(n17150) );
  INV_X1 U12504 ( .A(n10919), .ZN(n17165) );
  NAND2_X1 U12505 ( .A1(n10064), .A2(n10903), .ZN(n17167) );
  INV_X1 U12506 ( .A(n20543), .ZN(n20546) );
  INV_X1 U12507 ( .A(n11050), .ZN(n20611) );
  INV_X1 U12508 ( .A(n21092), .ZN(n20780) );
  INV_X1 U12509 ( .A(n20836), .ZN(n20843) );
  INV_X1 U12510 ( .A(n11087), .ZN(n20839) );
  INV_X1 U12511 ( .A(n12056), .ZN(n10895) );
  NAND2_X2 U12512 ( .A1(n10360), .A2(n10359), .ZN(n20415) );
  NAND3_X1 U12513 ( .A1(n9793), .A2(n10826), .A3(n10827), .ZN(n10359) );
  NAND2_X1 U12514 ( .A1(n20941), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20441) );
  INV_X1 U12515 ( .A(n20888), .ZN(n20884) );
  INV_X1 U12516 ( .A(n20880), .ZN(n20883) );
  OR2_X1 U12517 ( .A1(n20940), .A2(n20939), .ZN(n20948) );
  NOR2_X1 U12518 ( .A1(n11261), .A2(n11272), .ZN(n10885) );
  NOR2_X1 U12519 ( .A1(n11276), .A2(n10884), .ZN(n17778) );
  AND2_X1 U12520 ( .A1(n11263), .A2(n10885), .ZN(n10884) );
  CLKBUF_X1 U12521 ( .A(n11697), .Z(n17795) );
  NAND2_X1 U12522 ( .A1(n12022), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n14120) );
  NOR2_X1 U12523 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n17796) );
  NAND2_X1 U12524 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n21133) );
  INV_X1 U12525 ( .A(n17929), .ZN(n17918) );
  NOR2_X1 U12526 ( .A1(n17982), .A2(n18227), .ZN(n17974) );
  AND2_X1 U12527 ( .A1(n18004), .A2(n17277), .ZN(n17994) );
  NOR2_X1 U12528 ( .A1(n17994), .A2(n17995), .ZN(n17993) );
  NOR2_X1 U12529 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n18018), .ZN(n18003) );
  NOR2_X1 U12530 ( .A1(n18023), .A2(n18227), .ZN(n18013) );
  NOR2_X1 U12531 ( .A1(n18013), .A2(n18014), .ZN(n18012) );
  NAND2_X1 U12532 ( .A1(n17277), .A2(n10480), .ZN(n10479) );
  NAND2_X1 U12533 ( .A1(n18054), .A2(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n10480) );
  NOR2_X1 U12534 ( .A1(n18068), .A2(n19041), .ZN(n18054) );
  NAND2_X1 U12535 ( .A1(n18094), .A2(n19025), .ZN(n18068) );
  INV_X1 U12536 ( .A(n18098), .ZN(n18099) );
  NOR2_X1 U12537 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n18130), .ZN(n18119) );
  NOR2_X1 U12538 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n18156), .ZN(n18140) );
  NOR2_X1 U12539 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n18166), .ZN(n18165) );
  NOR3_X1 U12540 ( .A1(n18481), .A2(n10357), .A3(n10355), .ZN(n17558) );
  NAND2_X1 U12541 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(P3_EBX_REG_19__SCAN_IN), 
        .ZN(n10357) );
  AND2_X1 U12542 ( .A1(n9777), .A2(P3_EAX_REG_25__SCAN_IN), .ZN(n10255) );
  NAND2_X1 U12543 ( .A1(n11812), .A2(n18270), .ZN(n18551) );
  NAND2_X2 U12544 ( .A1(n14031), .A2(n11819), .ZN(n10660) );
  NOR2_X1 U12545 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11813) );
  OR2_X1 U12546 ( .A1(n17191), .A2(n17190), .ZN(n17279) );
  OAI21_X1 U12547 ( .B1(n14030), .B2(n18856), .A(n20170), .ZN(n18816) );
  INV_X1 U12548 ( .A(n17919), .ZN(n18858) );
  NAND2_X1 U12549 ( .A1(n17823), .A2(n17821), .ZN(n10382) );
  AND2_X1 U12550 ( .A1(n11795), .A2(n10468), .ZN(n11802) );
  AND2_X1 U12551 ( .A1(n9773), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n10468) );
  NOR2_X1 U12552 ( .A1(n18925), .A2(n10470), .ZN(n10469) );
  NAND2_X1 U12553 ( .A1(n11795), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n18924) );
  NAND2_X1 U12554 ( .A1(n10477), .A2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n10476) );
  INV_X1 U12555 ( .A(n19027), .ZN(n10477) );
  NOR2_X1 U12556 ( .A1(n19112), .A2(n19071), .ZN(n19069) );
  INV_X1 U12557 ( .A(n19112), .ZN(n18116) );
  AND2_X1 U12558 ( .A1(n11794), .A2(n9797), .ZN(n10481) );
  OR2_X1 U12559 ( .A1(n18184), .A2(n19097), .ZN(n19112) );
  INV_X1 U12560 ( .A(n19105), .ZN(n19145) );
  NAND2_X1 U12561 ( .A1(n18171), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18184) );
  NOR2_X1 U12562 ( .A1(n22084), .A2(n10077), .ZN(n10076) );
  NAND2_X1 U12563 ( .A1(n10075), .A2(n10078), .ZN(n19193) );
  NOR2_X1 U12564 ( .A1(n22149), .A2(n10077), .ZN(n10075) );
  INV_X1 U12565 ( .A(n17307), .ZN(n10387) );
  NAND2_X1 U12566 ( .A1(n18942), .A2(n9976), .ZN(n17592) );
  NOR2_X1 U12567 ( .A1(n19063), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n9976) );
  INV_X1 U12568 ( .A(n18942), .ZN(n17409) );
  NAND2_X1 U12569 ( .A1(n17334), .A2(n10285), .ZN(n17408) );
  NOR2_X1 U12570 ( .A1(n10286), .A2(n19259), .ZN(n10285) );
  OR2_X1 U12571 ( .A1(n17247), .A2(n17283), .ZN(n17407) );
  AND2_X1 U12572 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17372) );
  INV_X1 U12573 ( .A(n17434), .ZN(n9980) );
  AND2_X1 U12574 ( .A1(n19185), .A2(n17266), .ZN(n19043) );
  NAND2_X1 U12575 ( .A1(n19371), .A2(n10389), .ZN(n19329) );
  OR2_X1 U12576 ( .A1(n19366), .A2(n19452), .ZN(n10389) );
  AND2_X1 U12577 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n19354), .ZN(
        n19327) );
  OR2_X1 U12578 ( .A1(n19161), .A2(n10289), .ZN(n19102) );
  INV_X1 U12579 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n19101) );
  NAND2_X1 U12580 ( .A1(n10461), .A2(n10462), .ZN(n19125) );
  INV_X1 U12581 ( .A(n19162), .ZN(n10461) );
  INV_X1 U12582 ( .A(n19975), .ZN(n10368) );
  OR2_X1 U12583 ( .A1(n10371), .A2(n10370), .ZN(n10369) );
  INV_X1 U12584 ( .A(n19976), .ZN(n10370) );
  INV_X1 U12585 ( .A(n19080), .ZN(n19415) );
  NAND2_X1 U12586 ( .A1(n19219), .A2(n17305), .ZN(n19205) );
  NAND2_X1 U12587 ( .A1(n19205), .A2(n19206), .ZN(n19204) );
  XNOR2_X1 U12588 ( .A(n17303), .B(n10160), .ZN(n19220) );
  INV_X1 U12589 ( .A(n17304), .ZN(n10160) );
  NAND2_X1 U12590 ( .A1(n19220), .A2(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n19219) );
  AND2_X1 U12591 ( .A1(n11996), .A2(n11995), .ZN(n17927) );
  INV_X1 U12592 ( .A(n18256), .ZN(n19997) );
  NAND2_X1 U12593 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19611), .ZN(
        n19655) );
  AND4_X1 U12594 ( .A1(n11910), .A2(n11909), .A3(n11908), .A4(n11907), .ZN(
        n11925) );
  AND4_X1 U12595 ( .A1(n11929), .A2(n11928), .A3(n11927), .A4(n11926), .ZN(
        n11944) );
  NAND2_X1 U12596 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20002), .ZN(
        n19752) );
  NAND2_X1 U12597 ( .A1(n20002), .A2(n11982), .ZN(n20007) );
  NAND2_X1 U12598 ( .A1(n20175), .A2(n19530), .ZN(n19565) );
  AND4_X1 U12599 ( .A1(n13571), .A2(n13570), .A3(n13569), .A4(n21032), .ZN(
        n13572) );
  NAND2_X1 U12600 ( .A1(n12682), .A2(n21871), .ZN(n21907) );
  INV_X1 U12601 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n21194) );
  INV_X1 U12602 ( .A(n21256), .ZN(n21223) );
  AND2_X1 U12603 ( .A1(n14799), .A2(n14798), .ZN(n21174) );
  OR2_X1 U12604 ( .A1(n21251), .A2(n21249), .ZN(n21217) );
  INV_X1 U12605 ( .A(n15195), .ZN(n15145) );
  INV_X1 U12606 ( .A(n15194), .ZN(n15174) );
  AND2_X1 U12607 ( .A1(n15194), .A2(n21373), .ZN(n15175) );
  INV_X1 U12608 ( .A(n15145), .ZN(n15187) );
  INV_X1 U12609 ( .A(n15175), .ZN(n15192) );
  NAND2_X1 U12610 ( .A1(n10280), .A2(n9747), .ZN(n15202) );
  AND2_X1 U12611 ( .A1(n15296), .A2(n13857), .ZN(n15272) );
  OR2_X1 U12612 ( .A1(n14748), .A2(n21329), .ZN(n15274) );
  INV_X1 U12613 ( .A(n15274), .ZN(n15280) );
  NOR2_X2 U12614 ( .A1(n14748), .A2(n21327), .ZN(n15281) );
  AND2_X1 U12615 ( .A1(n13856), .A2(n14788), .ZN(n15296) );
  OAI21_X1 U12616 ( .B1(n17629), .B2(n13855), .A(n13854), .ZN(n13856) );
  AND2_X1 U12617 ( .A1(n13888), .A2(n13853), .ZN(n13854) );
  INV_X1 U12618 ( .A(n15292), .ZN(n15298) );
  NAND2_X1 U12619 ( .A1(n21301), .A2(n21281), .ZN(n21285) );
  AND2_X1 U12620 ( .A1(n13950), .A2(n17621), .ZN(n21283) );
  OR3_X1 U12621 ( .A1(n17629), .A2(n21146), .A3(n15908), .ZN(n13949) );
  INV_X2 U12622 ( .A(n15354), .ZN(n21322) );
  NOR2_X2 U12623 ( .A1(n21321), .A2(n12289), .ZN(n21311) );
  OAI21_X1 U12624 ( .B1(n14807), .B2(n14809), .A(n14808), .ZN(n15372) );
  INV_X1 U12625 ( .A(n13268), .ZN(n13237) );
  INV_X1 U12626 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n15416) );
  INV_X1 U12627 ( .A(n10054), .ZN(n13048) );
  OAI21_X1 U12628 ( .B1(n15029), .B2(n15028), .A(n15027), .ZN(n15511) );
  INV_X1 U12629 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n15550) );
  NAND2_X1 U12630 ( .A1(n14817), .A2(n14816), .ZN(n15598) );
  OAI211_X1 U12631 ( .C1(n15415), .C2(n9902), .A(n10108), .B(n10105), .ZN(
        n15374) );
  NOR2_X1 U12632 ( .A1(n10110), .A2(n10109), .ZN(n10108) );
  NAND2_X1 U12633 ( .A1(n10101), .A2(n10193), .ZN(n10456) );
  NAND2_X1 U12634 ( .A1(n10102), .A2(n15545), .ZN(n10101) );
  OAI21_X1 U12635 ( .B1(n10268), .B2(n15403), .A(n10100), .ZN(n10193) );
  OR2_X1 U12636 ( .A1(n15635), .A2(n13374), .ZN(n15630) );
  OR2_X1 U12637 ( .A1(n15793), .A2(n15768), .ZN(n15637) );
  NAND2_X1 U12638 ( .A1(n15402), .A2(n10266), .ZN(n10267) );
  AND2_X1 U12639 ( .A1(n15670), .A2(n13371), .ZN(n15651) );
  NAND2_X1 U12640 ( .A1(n12602), .A2(n15677), .ZN(n15435) );
  INV_X1 U12641 ( .A(n12602), .ZN(n15444) );
  NAND2_X1 U12642 ( .A1(n12598), .A2(n15518), .ZN(n15505) );
  INV_X1 U12643 ( .A(n15837), .ZN(n17697) );
  INV_X1 U12644 ( .A(n15864), .ZN(n17700) );
  INV_X1 U12645 ( .A(n10096), .ZN(n15571) );
  NAND2_X1 U12646 ( .A1(n15771), .A2(n15816), .ZN(n17681) );
  AND2_X1 U12647 ( .A1(n10293), .A2(n10292), .ZN(n15814) );
  INV_X1 U12648 ( .A(n10293), .ZN(n15765) );
  INV_X1 U12649 ( .A(n21819), .ZN(n21810) );
  INV_X1 U12651 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n21586) );
  AND2_X1 U12652 ( .A1(n15895), .A2(n21819), .ZN(n21815) );
  CLKBUF_X1 U12653 ( .A(n13864), .Z(n21585) );
  INV_X1 U12654 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n21326) );
  OAI21_X1 U12655 ( .B1(n15879), .B2(n17715), .A(n21476), .ZN(n21325) );
  NOR2_X1 U12656 ( .A1(n17629), .A2(n21704), .ZN(n15916) );
  INV_X1 U12657 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n15872) );
  NOR2_X1 U12658 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n15911) );
  OAI22_X1 U12659 ( .A1(n21346), .A2(n21345), .B1(n21642), .B2(n21472), .ZN(
        n21377) );
  OAI211_X1 U12660 ( .C1(n21344), .C2(n12682), .A(n21639), .B(n21340), .ZN(
        n21378) );
  OAI22_X1 U12661 ( .A1(n21413), .A2(n21412), .B1(n21642), .B2(n21530), .ZN(
        n21431) );
  INV_X1 U12662 ( .A(n21428), .ZN(n21430) );
  INV_X1 U12663 ( .A(n21461), .ZN(n21463) );
  OAI221_X1 U12664 ( .B1(n10676), .B2(n21704), .C1(n10676), .C2(n21478), .A(
        n21781), .ZN(n21495) );
  OAI21_X1 U12665 ( .B1(n21773), .B2(n21472), .A(n21471), .ZN(n21493) );
  OAI22_X1 U12666 ( .A1(n21532), .A2(n21531), .B1(n21530), .B2(n21773), .ZN(
        n21549) );
  INV_X1 U12667 ( .A(n21583), .ZN(n21574) );
  OAI211_X1 U12668 ( .C1(n10679), .C2(n21704), .A(n21639), .B(n21591), .ZN(
        n21608) );
  INV_X1 U12669 ( .A(n21577), .ZN(n21607) );
  OAI22_X1 U12670 ( .A1(n21644), .A2(n21643), .B1(n21642), .B2(n21774), .ZN(
        n21661) );
  OAI211_X1 U12671 ( .C1(n21644), .C2(n21641), .A(n21640), .B(n21639), .ZN(
        n21662) );
  INV_X1 U12672 ( .A(n21696), .ZN(n21687) );
  OAI211_X1 U12673 ( .C1(n10675), .C2(n21704), .A(n21781), .B(n21703), .ZN(
        n21724) );
  AND2_X1 U12674 ( .A1(n21776), .A2(n21697), .ZN(n21767) );
  OAI211_X1 U12675 ( .C1(n21797), .C2(n21782), .A(n21781), .B(n21780), .ZN(
        n21800) );
  OAI21_X1 U12676 ( .B1(n21774), .B2(n21773), .A(n21772), .ZN(n21798) );
  NAND2_X1 U12677 ( .A1(n21776), .A2(n21775), .ZN(n21869) );
  AND2_X1 U12678 ( .A1(n21776), .A2(n21666), .ZN(n21865) );
  NAND2_X1 U12679 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n21912) );
  INV_X1 U12680 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n21871) );
  INV_X1 U12681 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n21908) );
  INV_X1 U12682 ( .A(n21912), .ZN(n17713) );
  AND2_X1 U12683 ( .A1(n21143), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n21915) );
  INV_X1 U12684 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n21116) );
  INV_X1 U12685 ( .A(n11715), .ZN(n11716) );
  OAI21_X1 U12686 ( .B1(n14741), .B2(n20277), .A(n11714), .ZN(n11715) );
  NAND2_X1 U12687 ( .A1(n12018), .A2(n9708), .ZN(n11714) );
  NAND2_X1 U12688 ( .A1(n9914), .A2(n16342), .ZN(n11438) );
  INV_X1 U12689 ( .A(n11431), .ZN(n9914) );
  NAND2_X1 U12690 ( .A1(n11371), .A2(n10220), .ZN(n11431) );
  NOR2_X1 U12691 ( .A1(n11432), .A2(n10221), .ZN(n10220) );
  AND2_X1 U12692 ( .A1(n11427), .A2(n11430), .ZN(n16046) );
  AND2_X1 U12693 ( .A1(n11366), .A2(n11368), .ZN(n16085) );
  INV_X1 U12694 ( .A(n11364), .ZN(n16113) );
  AND2_X1 U12695 ( .A1(n11374), .A2(n11373), .ZN(n16128) );
  AOI21_X1 U12696 ( .B1(n11398), .B2(n11400), .A(n9913), .ZN(n11401) );
  NAND2_X1 U12697 ( .A1(n11397), .A2(n11396), .ZN(n10634) );
  INV_X1 U12698 ( .A(n16299), .ZN(n16261) );
  AND2_X1 U12699 ( .A1(n11436), .A2(n10154), .ZN(n11386) );
  NAND2_X1 U12700 ( .A1(n11384), .A2(n11383), .ZN(n10154) );
  NAND2_X1 U12701 ( .A1(n10633), .A2(n11298), .ZN(n11345) );
  INV_X1 U12702 ( .A(n9708), .ZN(n20273) );
  INV_X1 U12703 ( .A(n10964), .ZN(n10487) );
  INV_X1 U12704 ( .A(n16174), .ZN(n16302) );
  OR2_X1 U12705 ( .A1(n11638), .A2(n11637), .ZN(n14323) );
  OR2_X1 U12706 ( .A1(n11621), .A2(n11620), .ZN(n14345) );
  OR2_X1 U12707 ( .A1(n11603), .A2(n11602), .ZN(n16382) );
  OR2_X1 U12708 ( .A1(n11567), .A2(n11566), .ZN(n14319) );
  OR2_X1 U12709 ( .A1(n11549), .A2(n11548), .ZN(n14336) );
  OR2_X1 U12710 ( .A1(n13800), .A2(n13786), .ZN(n20673) );
  NAND2_X1 U12711 ( .A1(n10600), .A2(n10603), .ZN(n16339) );
  NAND2_X1 U12712 ( .A1(n14456), .A2(n10605), .ZN(n10600) );
  AND2_X1 U12713 ( .A1(n14677), .A2(n14329), .ZN(n16490) );
  NAND2_X1 U12714 ( .A1(n14677), .A2(n20369), .ZN(n16495) );
  AND2_X1 U12715 ( .A1(n16487), .A2(n20298), .ZN(n20283) );
  AND2_X1 U12716 ( .A1(n16519), .A2(n9722), .ZN(n20304) );
  AND2_X1 U12717 ( .A1(n16481), .A2(n13821), .ZN(n20311) );
  INV_X1 U12718 ( .A(n13746), .ZN(n20313) );
  INV_X1 U12719 ( .A(n20347), .ZN(n20340) );
  INV_X1 U12720 ( .A(n21125), .ZN(n20344) );
  NAND2_X1 U12721 ( .A1(n20343), .A2(n21125), .ZN(n20347) );
  NOR2_X2 U12722 ( .A1(n13633), .A2(n9735), .ZN(n20350) );
  NAND2_X1 U12723 ( .A1(n16673), .A2(n9896), .ZN(n16627) );
  INV_X1 U12724 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17723) );
  INV_X1 U12725 ( .A(n16730), .ZN(n20355) );
  NAND2_X1 U12726 ( .A1(n10526), .A2(n11159), .ZN(n14218) );
  OAI211_X1 U12727 ( .C1(n13498), .C2(n10215), .A(n10214), .B(n10213), .ZN(
        n14724) );
  AOI21_X1 U12728 ( .B1(n16534), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n10128), .ZN(n16527) );
  NAND2_X1 U12729 ( .A1(n10129), .A2(n9796), .ZN(n10128) );
  NAND2_X1 U12730 ( .A1(n17738), .A2(n10316), .ZN(n10315) );
  NAND2_X1 U12731 ( .A1(n16849), .A2(n16848), .ZN(n10316) );
  NAND2_X1 U12732 ( .A1(n16911), .A2(n17738), .ZN(n16914) );
  NAND2_X1 U12733 ( .A1(n16673), .A2(n9892), .ZN(n16643) );
  OR2_X1 U12734 ( .A1(n16938), .A2(n14761), .ZN(n16892) );
  NAND2_X1 U12735 ( .A1(n10549), .A2(n10552), .ZN(n16657) );
  NAND2_X1 U12736 ( .A1(n16678), .A2(n10554), .ZN(n10549) );
  XNOR2_X1 U12737 ( .A(n9960), .B(n16693), .ZN(n16984) );
  CLKBUF_X1 U12738 ( .A(n16726), .Z(n16727) );
  XNOR2_X1 U12739 ( .A(n9961), .B(n16756), .ZN(n17056) );
  NAND2_X1 U12740 ( .A1(n16754), .A2(n10365), .ZN(n16755) );
  AND2_X1 U12741 ( .A1(n17064), .A2(n17063), .ZN(n17720) );
  AND2_X1 U12742 ( .A1(n10519), .A2(n10520), .ZN(n17062) );
  NAND2_X1 U12743 ( .A1(n14701), .A2(n11494), .ZN(n16255) );
  NAND2_X1 U12744 ( .A1(n14751), .A2(n14756), .ZN(n17111) );
  INV_X1 U12745 ( .A(n13778), .ZN(n13790) );
  INV_X1 U12746 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n21114) );
  INV_X1 U12747 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n21096) );
  NAND2_X1 U12748 ( .A1(n21090), .A2(n20613), .ZN(n21091) );
  INV_X1 U12749 ( .A(n20673), .ZN(n21111) );
  NAND2_X1 U12750 ( .A1(n10595), .A2(n10592), .ZN(n13805) );
  INV_X1 U12751 ( .A(n10589), .ZN(n10595) );
  AND2_X1 U12752 ( .A1(n20448), .A2(n21114), .ZN(n20442) );
  OAI21_X1 U12753 ( .B1(n20515), .B2(n20514), .A(n20513), .ZN(n20536) );
  INV_X1 U12754 ( .A(n20531), .ZN(n20540) );
  NOR2_X1 U12755 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20582), .ZN(
        n20568) );
  INV_X1 U12756 ( .A(n20620), .ZN(n20635) );
  INV_X1 U12757 ( .A(n20670), .ZN(n20662) );
  INV_X1 U12758 ( .A(n20706), .ZN(n20666) );
  INV_X1 U12759 ( .A(n20655), .ZN(n20667) );
  AND2_X1 U12760 ( .A1(n20647), .A2(n20646), .ZN(n20665) );
  OAI21_X1 U12761 ( .B1(n20721), .B2(n20717), .A(n20716), .ZN(n20746) );
  OAI21_X1 U12762 ( .B1(n20781), .B2(n20751), .A(n20750), .ZN(n20774) );
  NOR2_X1 U12763 ( .A1(n20812), .A2(n20810), .ZN(n20831) );
  NAND2_X1 U12764 ( .A1(n20392), .A2(n20391), .ZN(n20848) );
  NAND2_X1 U12765 ( .A1(n20399), .A2(n20398), .ZN(n20851) );
  NAND2_X1 U12766 ( .A1(n20407), .A2(n20406), .ZN(n20854) );
  NAND2_X1 U12767 ( .A1(n20414), .A2(n20413), .ZN(n20857) );
  NAND2_X1 U12768 ( .A1(n20422), .A2(n20421), .ZN(n20860) );
  NAND2_X1 U12769 ( .A1(n20430), .A2(n20429), .ZN(n20863) );
  NAND2_X1 U12770 ( .A1(n20439), .A2(n20438), .ZN(n20868) );
  NAND2_X1 U12771 ( .A1(n20375), .A2(n20374), .ZN(n20952) );
  NAND2_X1 U12772 ( .A1(n20372), .A2(n20371), .ZN(n20951) );
  INV_X1 U12773 ( .A(n20876), .ZN(n20949) );
  INV_X1 U12774 ( .A(n20895), .ZN(n20957) );
  INV_X1 U12775 ( .A(n20848), .ZN(n20963) );
  NAND2_X1 U12776 ( .A1(n20397), .A2(n20396), .ZN(n20966) );
  INV_X1 U12777 ( .A(n20900), .ZN(n20964) );
  INV_X1 U12778 ( .A(n20851), .ZN(n20969) );
  NAND2_X1 U12779 ( .A1(n20405), .A2(n20404), .ZN(n20972) );
  INV_X1 U12780 ( .A(n20854), .ZN(n20975) );
  NAND2_X1 U12781 ( .A1(n20412), .A2(n20411), .ZN(n21922) );
  INV_X1 U12782 ( .A(n20910), .ZN(n21919) );
  NAND2_X1 U12783 ( .A1(n20420), .A2(n20419), .ZN(n20980) );
  INV_X1 U12784 ( .A(n20915), .ZN(n20978) );
  INV_X1 U12785 ( .A(n20860), .ZN(n20983) );
  NAND2_X1 U12786 ( .A1(n20428), .A2(n20427), .ZN(n20986) );
  INV_X1 U12787 ( .A(n20863), .ZN(n20989) );
  INV_X1 U12788 ( .A(n20938), .ZN(n20991) );
  NAND2_X1 U12789 ( .A1(n20435), .A2(n20434), .ZN(n20994) );
  INV_X1 U12790 ( .A(n20959), .ZN(n20996) );
  INV_X1 U12791 ( .A(n20926), .ZN(n20990) );
  INV_X1 U12792 ( .A(n20868), .ZN(n21000) );
  INV_X1 U12793 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n21132) );
  NOR2_X1 U12794 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n21135) );
  AOI211_X1 U12795 ( .C1(P2_STATE_REG_1__SCAN_IN), .C2(P2_STATE_REG_2__SCAN_IN), .A(P2_STATE_REG_0__SCAN_IN), .B(n21013), .ZN(n21129) );
  INV_X1 U12796 ( .A(P2_BE_N_REG_3__SCAN_IN), .ZN(n22104) );
  NAND2_X1 U12797 ( .A1(READY22_REG_SCAN_IN), .A2(READY2), .ZN(n20181) );
  INV_X1 U12798 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n20175) );
  OR2_X1 U12799 ( .A1(n17950), .A2(n17949), .ZN(n10670) );
  INV_X1 U12800 ( .A(n17952), .ZN(n10465) );
  NOR2_X1 U12801 ( .A1(n17993), .A2(n18227), .ZN(n17983) );
  NOR2_X1 U12802 ( .A1(n17983), .A2(n17984), .ZN(n17982) );
  AND2_X1 U12803 ( .A1(n18009), .A2(n11999), .ZN(n17988) );
  NOR2_X1 U12804 ( .A1(n18012), .A2(n18227), .ZN(n18006) );
  NOR2_X1 U12805 ( .A1(n18024), .A2(n18997), .ZN(n18023) );
  AND2_X1 U12806 ( .A1(n18033), .A2(n17277), .ZN(n18024) );
  INV_X1 U12807 ( .A(n10068), .ZN(n18035) );
  AND2_X1 U12808 ( .A1(n10479), .A2(n10478), .ZN(n18044) );
  INV_X1 U12809 ( .A(n19018), .ZN(n10478) );
  INV_X1 U12810 ( .A(n10479), .ZN(n18045) );
  NOR2_X1 U12811 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n18081), .ZN(n18072) );
  NOR2_X1 U12812 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n18106), .ZN(n18092) );
  INV_X1 U12813 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n18633) );
  INV_X1 U12814 ( .A(n18259), .ZN(n18295) );
  INV_X1 U12815 ( .A(n18288), .ZN(n18252) );
  NOR2_X2 U12816 ( .A1(n20138), .A2(n18298), .ZN(n18288) );
  NAND4_X1 U12817 ( .A1(n14191), .A2(n20177), .A3(n20051), .A4(n20041), .ZN(
        n18242) );
  NOR2_X1 U12818 ( .A1(n18002), .A2(n18352), .ZN(n18357) );
  AND2_X1 U12819 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(n18388), .ZN(n18367) );
  NOR2_X1 U12820 ( .A1(n18358), .A2(n18409), .ZN(n18388) );
  NOR2_X1 U12821 ( .A1(n18640), .A2(n10347), .ZN(n17462) );
  NAND2_X1 U12822 ( .A1(n10348), .A2(P3_EBX_REG_11__SCAN_IN), .ZN(n10347) );
  INV_X1 U12823 ( .A(n18581), .ZN(n10348) );
  INV_X2 U12824 ( .A(n18667), .ZN(n18661) );
  AND2_X1 U12825 ( .A1(n10349), .A2(n9876), .ZN(n18670) );
  NOR2_X1 U12826 ( .A1(n22041), .A2(n18701), .ZN(n18696) );
  NAND2_X1 U12827 ( .A1(n18715), .A2(n10254), .ZN(n18701) );
  AND2_X1 U12828 ( .A1(n10255), .A2(P3_EAX_REG_26__SCAN_IN), .ZN(n10254) );
  NAND2_X1 U12829 ( .A1(n18715), .A2(n19561), .ZN(n18709) );
  NAND2_X1 U12830 ( .A1(n18715), .A2(n9777), .ZN(n18710) );
  AND2_X1 U12831 ( .A1(n18676), .A2(n9887), .ZN(n18677) );
  NOR2_X1 U12832 ( .A1(n18725), .A2(n18723), .ZN(n10257) );
  INV_X1 U12833 ( .A(n18760), .ZN(n18748) );
  AND2_X1 U12834 ( .A1(n18675), .A2(P3_EAX_REG_15__SCAN_IN), .ZN(n10259) );
  NAND2_X1 U12835 ( .A1(n18676), .A2(n10258), .ZN(n18757) );
  AND4_X1 U12836 ( .A1(n11856), .A2(n11855), .A3(n11854), .A4(n11853), .ZN(
        n11857) );
  AND4_X1 U12837 ( .A1(n11845), .A2(n11844), .A3(n11843), .A4(n11842), .ZN(
        n11860) );
  NAND2_X1 U12838 ( .A1(n18676), .A2(n18675), .ZN(n18761) );
  NAND2_X1 U12839 ( .A1(n10252), .A2(n10250), .ZN(n18797) );
  NOR2_X1 U12840 ( .A1(n18671), .A2(n10251), .ZN(n10250) );
  INV_X1 U12841 ( .A(n18672), .ZN(n10252) );
  NOR2_X1 U12842 ( .A1(n18895), .A2(n14093), .ZN(n18805) );
  INV_X1 U12843 ( .A(n17279), .ZN(n18811) );
  INV_X1 U12844 ( .A(n18785), .ZN(n18812) );
  AND2_X1 U12845 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n14223), .ZN(n18809) );
  NAND2_X2 U12846 ( .A1(n10005), .A2(n9977), .ZN(n17295) );
  NOR2_X1 U12847 ( .A1(n9825), .A2(n9759), .ZN(n10005) );
  NAND2_X1 U12848 ( .A1(n14246), .A2(P3_EAX_REG_1__SCAN_IN), .ZN(n18672) );
  NOR2_X1 U12849 ( .A1(n14159), .A2(n10007), .ZN(n10006) );
  OR2_X1 U12850 ( .A1(n14091), .A2(n14090), .ZN(n14092) );
  INV_X1 U12851 ( .A(n10349), .ZN(n14089) );
  INV_X1 U12852 ( .A(n18815), .ZN(n18796) );
  NOR2_X1 U12853 ( .A1(n18857), .A2(n18816), .ZN(n18843) );
  INV_X1 U12854 ( .A(n18843), .ZN(n18855) );
  INV_X1 U12855 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n22041) );
  NOR2_X1 U12856 ( .A1(n18857), .A2(n20035), .ZN(n18900) );
  NAND2_X1 U12857 ( .A1(n17379), .A2(n17817), .ZN(n10385) );
  OR2_X1 U12858 ( .A1(n17432), .A2(n19150), .ZN(n10164) );
  INV_X1 U12859 ( .A(n17344), .ZN(n10163) );
  NOR3_X1 U12860 ( .A1(n11801), .A2(n10476), .A3(n18998), .ZN(n18981) );
  INV_X1 U12861 ( .A(n18975), .ZN(n18989) );
  OR2_X1 U12862 ( .A1(n19079), .A2(n19295), .ZN(n19037) );
  NOR2_X1 U12863 ( .A1(n18145), .A2(n18134), .ZN(n19098) );
  NAND2_X1 U12864 ( .A1(n19080), .A2(n10167), .ZN(n10166) );
  INV_X1 U12865 ( .A(n10013), .ZN(n17346) );
  INV_X1 U12866 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n22084) );
  NAND2_X1 U12867 ( .A1(n9975), .A2(n17246), .ZN(n19196) );
  NOR2_X1 U12868 ( .A1(n18244), .A2(n22149), .ZN(n19208) );
  INV_X1 U12869 ( .A(n19207), .ZN(n19231) );
  INV_X1 U12870 ( .A(n19882), .ZN(n19921) );
  INV_X1 U12871 ( .A(n19215), .ZN(n19248) );
  NAND2_X1 U12872 ( .A1(n19207), .A2(n19218), .ZN(n19194) );
  OAI21_X1 U12873 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n20178), .A(n17930), 
        .ZN(n19207) );
  NAND2_X1 U12874 ( .A1(n20175), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n19068) );
  INV_X1 U12875 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n20044) );
  NOR2_X1 U12876 ( .A1(n17387), .A2(n10010), .ZN(n17393) );
  NOR2_X1 U12877 ( .A1(n17325), .A2(n10011), .ZN(n10010) );
  AND2_X1 U12878 ( .A1(n10284), .A2(n10282), .ZN(n17396) );
  NAND2_X1 U12879 ( .A1(n19488), .A2(n20019), .ZN(n19355) );
  NAND2_X1 U12880 ( .A1(n19279), .A2(n19416), .ZN(n19371) );
  INV_X1 U12881 ( .A(n19986), .ZN(n19424) );
  NOR2_X1 U12882 ( .A1(n19162), .A2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n19136) );
  NOR2_X1 U12883 ( .A1(n19403), .A2(n19517), .ZN(n19437) );
  NAND2_X1 U12884 ( .A1(n10454), .A2(n17238), .ZN(n19223) );
  NAND2_X1 U12885 ( .A1(n19238), .A2(n17236), .ZN(n10454) );
  INV_X1 U12886 ( .A(n19457), .ZN(n19517) );
  INV_X1 U12887 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n20022) );
  INV_X1 U12888 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n18236) );
  NAND2_X1 U12889 ( .A1(n14024), .A2(n14023), .ZN(n20155) );
  INV_X1 U12890 ( .A(n20179), .ZN(n20042) );
  NOR2_X1 U12891 ( .A1(n20175), .A2(P3_STATE2_REG_1__SCAN_IN), .ZN(n20048) );
  INV_X1 U12892 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n20138) );
  NAND2_X1 U12893 ( .A1(n20073), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n20185) );
  AND2_X2 U12894 ( .A1(n13562), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n21327)
         );
  INV_X1 U12895 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n21032) );
  OAI21_X1 U12896 ( .B1(n14364), .B2(n17647), .A(n13547), .ZN(n13548) );
  AND4_X1 U12897 ( .A1(n15111), .A2(n15110), .A3(n15109), .A4(n15108), .ZN(
        n15112) );
  AOI21_X1 U12898 ( .B1(n9753), .B2(n10280), .A(n15362), .ZN(n15363) );
  NAND2_X1 U12899 ( .A1(n10171), .A2(n9987), .ZN(P1_U2972) );
  NAND2_X1 U12900 ( .A1(n15607), .A2(n12669), .ZN(n10171) );
  OAI21_X1 U12901 ( .B1(n15625), .B2(n21153), .A(n15398), .ZN(P1_U2973) );
  AND2_X1 U12902 ( .A1(n13494), .A2(n9805), .ZN(n10142) );
  OAI21_X1 U12903 ( .B1(n15590), .B2(n15864), .A(n10294), .ZN(P1_U3001) );
  NOR3_X1 U12904 ( .A1(n10296), .A2(n15588), .A3(n10295), .ZN(n10294) );
  NOR2_X1 U12905 ( .A1(n15586), .A2(n15587), .ZN(n10296) );
  AND2_X1 U12906 ( .A1(n15589), .A2(n17698), .ZN(n10295) );
  AOI211_X1 U12907 ( .C1(n15949), .C2(n9708), .A(n15948), .B(n15947), .ZN(
        n15950) );
  NAND2_X1 U12908 ( .A1(n10620), .A2(n10618), .ZN(n16309) );
  NAND2_X1 U12909 ( .A1(n10613), .A2(n10612), .ZN(n10618) );
  NAND2_X1 U12910 ( .A1(n10148), .A2(n10584), .ZN(P2_U2890) );
  NAND2_X1 U12911 ( .A1(n10153), .A2(n10149), .ZN(n10148) );
  NAND2_X1 U12912 ( .A1(n10616), .A2(n16318), .ZN(n10153) );
  OAI21_X1 U12913 ( .B1(n16795), .B2(n16762), .A(n9937), .ZN(P2_U2988) );
  INV_X1 U12914 ( .A(n9938), .ZN(n9937) );
  INV_X1 U12915 ( .A(n16549), .ZN(n9939) );
  NAND2_X1 U12916 ( .A1(n16835), .A2(n20357), .ZN(n16586) );
  NAND2_X1 U12917 ( .A1(n10125), .A2(n10124), .ZN(n10123) );
  NAND2_X1 U12918 ( .A1(n10317), .A2(n16848), .ZN(n10126) );
  NAND2_X1 U12919 ( .A1(n16611), .A2(n10116), .ZN(P2_U2994) );
  NAND2_X1 U12920 ( .A1(n10205), .A2(n10202), .ZN(n16623) );
  INV_X1 U12921 ( .A(n9911), .ZN(n9910) );
  OAI21_X1 U12922 ( .B1(n16963), .B2(n16737), .A(n16671), .ZN(n9911) );
  INV_X1 U12923 ( .A(n9950), .ZN(n12094) );
  OAI21_X1 U12924 ( .B1(n14736), .B2(n17082), .A(n9951), .ZN(n9950) );
  NAND2_X1 U12925 ( .A1(n14735), .A2(n17738), .ZN(n10578) );
  NAND2_X1 U12926 ( .A1(n9832), .A2(n17748), .ZN(n10406) );
  OAI211_X1 U12927 ( .C1(n16798), .C2(n17101), .A(n10168), .B(n10366), .ZN(
        P2_U3020) );
  NOR2_X1 U12928 ( .A1(n16796), .A2(n10367), .ZN(n10366) );
  NAND2_X1 U12929 ( .A1(n10169), .A2(n17738), .ZN(n10168) );
  INV_X1 U12930 ( .A(n16879), .ZN(n16889) );
  OAI21_X1 U12931 ( .B1(n10467), .B2(n20051), .A(n10464), .ZN(P3_U2641) );
  XNOR2_X1 U12932 ( .A(n17946), .B(n17947), .ZN(n10467) );
  NOR3_X1 U12933 ( .A1(n10466), .A2(n10670), .A3(n10465), .ZN(n10464) );
  NOR2_X1 U12934 ( .A1(n17956), .A2(P3_EBX_REG_30__SCAN_IN), .ZN(n10466) );
  NAND2_X1 U12935 ( .A1(n10071), .A2(n10069), .ZN(P3_U2642) );
  NOR2_X1 U12936 ( .A1(n17958), .A2(n10072), .ZN(n10071) );
  INV_X1 U12937 ( .A(n10070), .ZN(n10069) );
  NOR2_X1 U12938 ( .A1(n18481), .A2(n18462), .ZN(n18429) );
  NAND2_X1 U12939 ( .A1(n10246), .A2(n10241), .ZN(P3_U2704) );
  NAND2_X1 U12940 ( .A1(n18678), .A2(P3_EAX_REG_30__SCAN_IN), .ZN(n10246) );
  NOR2_X1 U12941 ( .A1(n10243), .A2(n10242), .ZN(n10241) );
  NAND2_X1 U12942 ( .A1(n17816), .A2(n19172), .ZN(n10386) );
  NOR2_X1 U12943 ( .A1(n19250), .A2(n10385), .ZN(n10384) );
  NAND2_X1 U12944 ( .A1(n10165), .A2(n10161), .ZN(P3_U2804) );
  AOI21_X1 U12945 ( .B1(n18946), .B2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n10162), .ZN(n10161) );
  NAND2_X1 U12946 ( .A1(n18975), .A2(n9745), .ZN(n10165) );
  NAND2_X1 U12947 ( .A1(n10164), .A2(n10163), .ZN(n10162) );
  AOI21_X1 U12948 ( .B1(n19296), .B2(n10392), .A(n10390), .ZN(n19289) );
  NAND2_X1 U12949 ( .A1(n17836), .A2(U214), .ZN(U212) );
  INV_X2 U12950 ( .A(n12298), .ZN(n12289) );
  OR2_X1 U12951 ( .A1(n15554), .A2(n12606), .ZN(n9740) );
  NOR2_X1 U12952 ( .A1(n15998), .A2(n10535), .ZN(n15956) );
  AND2_X1 U12953 ( .A1(n16054), .A2(n9770), .ZN(n9741) );
  AND2_X1 U12954 ( .A1(n9884), .A2(n9758), .ZN(n9742) );
  AND2_X1 U12955 ( .A1(n10207), .A2(n16762), .ZN(n9743) );
  AND2_X1 U12956 ( .A1(n11159), .A2(n14252), .ZN(n9744) );
  INV_X1 U12957 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n22099) );
  AND3_X1 U12958 ( .A1(n19264), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        n17269), .ZN(n9745) );
  AND2_X1 U12959 ( .A1(n9780), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n9746) );
  OR2_X1 U12960 ( .A1(n14821), .A2(n10654), .ZN(n9747) );
  NAND2_X1 U12961 ( .A1(n14271), .A2(n14270), .ZN(n14321) );
  NOR3_X1 U12962 ( .A1(n14904), .A2(n14897), .A3(n14881), .ZN(n14863) );
  NAND2_X1 U12963 ( .A1(n14381), .A2(n14380), .ZN(n16371) );
  NAND2_X1 U12964 ( .A1(n10567), .A2(n10684), .ZN(n14264) );
  OR2_X1 U12965 ( .A1(n14905), .A2(n10649), .ZN(n14879) );
  OR2_X1 U12966 ( .A1(n14973), .A2(n14974), .ZN(n14962) );
  NAND2_X1 U12967 ( .A1(n14050), .A2(n14051), .ZN(n14055) );
  AND2_X1 U12968 ( .A1(n10490), .A2(n21908), .ZN(n9748) );
  AND2_X1 U12969 ( .A1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n9749) );
  NAND2_X1 U12970 ( .A1(n10572), .A2(n11664), .ZN(n16099) );
  NAND2_X1 U12971 ( .A1(n12755), .A2(n9884), .ZN(n15148) );
  NOR2_X1 U12972 ( .A1(n14315), .A2(n14353), .ZN(n14352) );
  OR2_X1 U12973 ( .A1(n15980), .A2(n11300), .ZN(n16524) );
  AND3_X1 U12974 ( .A1(n10933), .A2(n20400), .A3(n10892), .ZN(n9750) );
  AND2_X1 U12975 ( .A1(n14456), .A2(n14455), .ZN(n9751) );
  AND2_X1 U12976 ( .A1(n10674), .A2(n9811), .ZN(n9752) );
  AND2_X1 U12977 ( .A1(n9747), .A2(n21328), .ZN(n9753) );
  AND2_X1 U12978 ( .A1(n13810), .A2(n10575), .ZN(n9754) );
  AND2_X1 U12979 ( .A1(n10457), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n9755) );
  AND2_X1 U12980 ( .A1(n15383), .A2(n9904), .ZN(n9756) );
  AND2_X1 U12981 ( .A1(n9821), .A2(n17664), .ZN(n9757) );
  AND2_X1 U12982 ( .A1(n10643), .A2(n15140), .ZN(n9758) );
  NAND4_X1 U12983 ( .A1(n14168), .A2(n14167), .A3(n14166), .A4(n14165), .ZN(
        n9759) );
  AND2_X1 U12984 ( .A1(n11121), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n9760) );
  NAND2_X1 U12985 ( .A1(n16524), .A2(n16777), .ZN(n9761) );
  AND2_X1 U12986 ( .A1(n9749), .A2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n9762) );
  OR2_X1 U12987 ( .A1(n10657), .A2(n13304), .ZN(n9763) );
  AND3_X1 U12988 ( .A1(n16625), .A2(n14763), .A3(n9840), .ZN(n9764) );
  AND2_X1 U12989 ( .A1(n9752), .A2(n9810), .ZN(n9765) );
  INV_X1 U12990 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n22149) );
  AND2_X1 U12991 ( .A1(n10034), .A2(n16647), .ZN(n9766) );
  OR2_X1 U12992 ( .A1(n10400), .A2(n10033), .ZN(n10402) );
  INV_X1 U12993 ( .A(n10402), .ZN(n10403) );
  INV_X1 U12994 ( .A(n12755), .ZN(n10642) );
  AND2_X1 U12995 ( .A1(n10503), .A2(n15030), .ZN(n9767) );
  NOR2_X1 U12996 ( .A1(n10622), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n9768) );
  BUF_X2 U12997 ( .A(n10986), .Z(n10991) );
  INV_X1 U12998 ( .A(n10991), .ZN(n17744) );
  AND2_X1 U12999 ( .A1(n11500), .A2(n9882), .ZN(n9769) );
  NAND2_X1 U13000 ( .A1(n14271), .A2(n9859), .ZN(n14354) );
  NAND2_X1 U13001 ( .A1(n9870), .A2(n14701), .ZN(n16240) );
  OR2_X1 U13002 ( .A1(n16368), .A2(n9722), .ZN(n16388) );
  INV_X1 U13003 ( .A(n16388), .ZN(n10619) );
  AND2_X1 U13004 ( .A1(n9868), .A2(n10539), .ZN(n9770) );
  NAND2_X1 U13005 ( .A1(n13811), .A2(n9754), .ZN(n9771) );
  INV_X1 U13006 ( .A(n11355), .ZN(n10632) );
  INV_X1 U13007 ( .A(n11428), .ZN(n10221) );
  OR2_X1 U13008 ( .A1(n20298), .A2(n9869), .ZN(n9772) );
  AND2_X1 U13009 ( .A1(n15303), .A2(n12618), .ZN(n12623) );
  AND2_X1 U13010 ( .A1(n10469), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9773) );
  AND2_X1 U13011 ( .A1(n9770), .A2(n16024), .ZN(n9774) );
  AND2_X1 U13012 ( .A1(n10598), .A2(n16366), .ZN(n9775) );
  AND2_X1 U13013 ( .A1(n10619), .A2(n10615), .ZN(n9776) );
  AND2_X1 U13014 ( .A1(n19561), .A2(P3_EAX_REG_24__SCAN_IN), .ZN(n9777) );
  NAND2_X1 U13015 ( .A1(n16865), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n9778) );
  AND2_X1 U13016 ( .A1(n10522), .A2(n11149), .ZN(n9779) );
  AND2_X1 U13017 ( .A1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n9780) );
  AND2_X2 U13018 ( .A1(n14123), .A2(n10686), .ZN(n10733) );
  NAND2_X1 U13019 ( .A1(n12755), .A2(n9742), .ZN(n14989) );
  NAND2_X1 U13020 ( .A1(n19488), .A2(n10376), .ZN(n10378) );
  AND2_X2 U13021 ( .A1(n9733), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10764) );
  NAND2_X1 U13022 ( .A1(n16713), .A2(n10522), .ZN(n16553) );
  AND2_X1 U13023 ( .A1(n13321), .A2(n12663), .ZN(n9782) );
  AND2_X1 U13024 ( .A1(n15554), .A2(n15384), .ZN(n12604) );
  AND2_X1 U13025 ( .A1(n10156), .A2(n10625), .ZN(n9784) );
  OAI21_X1 U13026 ( .B1(n10455), .B2(n9931), .A(n12415), .ZN(n9930) );
  NAND2_X1 U13027 ( .A1(n11382), .A2(n11392), .ZN(n11391) );
  NAND2_X1 U13028 ( .A1(n15462), .A2(n15461), .ZN(n15441) );
  NOR2_X1 U13029 ( .A1(n14766), .A2(n10573), .ZN(n16082) );
  NAND2_X1 U13030 ( .A1(n11674), .A2(n11673), .ZN(n16047) );
  AND2_X1 U13031 ( .A1(n14381), .A2(n10598), .ZN(n9787) );
  INV_X1 U13032 ( .A(n12016), .ZN(n10050) );
  NOR2_X1 U13033 ( .A1(n14905), .A2(n10646), .ZN(n14866) );
  NOR2_X1 U13034 ( .A1(n14905), .A2(n14907), .ZN(n14890) );
  NAND2_X1 U13035 ( .A1(n16074), .A2(n16609), .ZN(n16060) );
  OR2_X1 U13036 ( .A1(n14904), .A2(n14897), .ZN(n9788) );
  NAND2_X1 U13037 ( .A1(n12755), .A2(n10279), .ZN(n14973) );
  INV_X1 U13038 ( .A(n14179), .ZN(n19539) );
  OR2_X1 U13039 ( .A1(n11801), .A2(n19027), .ZN(n9789) );
  NAND2_X1 U13040 ( .A1(n14064), .A2(n14063), .ZN(n14208) );
  AND4_X1 U13041 ( .A1(n14154), .A2(n14153), .A3(n14152), .A4(n14151), .ZN(
        n9790) );
  INV_X1 U13042 ( .A(n12267), .ZN(n12333) );
  AND2_X1 U13043 ( .A1(n14046), .A2(n14054), .ZN(n14050) );
  INV_X1 U13044 ( .A(n10371), .ZN(n19990) );
  OR3_X1 U13045 ( .A1(n17919), .A2(n14030), .A3(n9816), .ZN(n10371) );
  AND2_X1 U13046 ( .A1(n12485), .A2(n12484), .ZN(n12508) );
  NOR2_X1 U13047 ( .A1(n14766), .A2(n10570), .ZN(n16071) );
  OR3_X1 U13048 ( .A1(n11435), .A2(n11300), .A3(n22170), .ZN(n9791) );
  NAND2_X1 U13049 ( .A1(n12105), .A2(n12106), .ZN(n12104) );
  INV_X1 U13050 ( .A(n10990), .ZN(n10183) );
  NAND2_X1 U13051 ( .A1(n15177), .A2(n15168), .ZN(n15162) );
  OR2_X1 U13052 ( .A1(n14315), .A2(n10545), .ZN(n9792) );
  AND3_X1 U13053 ( .A1(n10824), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n10825), .ZN(n9793) );
  OR2_X1 U13054 ( .A1(n14315), .A2(n10542), .ZN(n9794) );
  OR3_X1 U13055 ( .A1(n18481), .A2(n10357), .A3(n10356), .ZN(n9795) );
  OR2_X1 U13056 ( .A1(n16523), .A2(n16524), .ZN(n9796) );
  NOR2_X1 U13057 ( .A1(n14840), .A2(n10507), .ZN(n14814) );
  AND2_X1 U13058 ( .A1(n10483), .A2(n10482), .ZN(n9797) );
  INV_X1 U13059 ( .A(n10253), .ZN(n14246) );
  NOR2_X1 U13060 ( .A1(n10642), .A2(n10641), .ZN(n15139) );
  NOR2_X1 U13061 ( .A1(n17919), .A2(n14030), .ZN(n9798) );
  AND2_X1 U13062 ( .A1(n10271), .A2(n15168), .ZN(n15156) );
  AND2_X1 U13063 ( .A1(n13496), .A2(n12016), .ZN(n9799) );
  OR2_X1 U13064 ( .A1(n17930), .A2(n20171), .ZN(n19235) );
  NAND2_X1 U13065 ( .A1(n11302), .A2(n11462), .ZN(n11436) );
  INV_X1 U13066 ( .A(n11436), .ZN(n9913) );
  AND2_X1 U13067 ( .A1(n11288), .A2(n11304), .ZN(n9800) );
  NAND2_X1 U13068 ( .A1(n11354), .A2(n11355), .ZN(n11353) );
  AND2_X1 U13069 ( .A1(n10404), .A2(n11425), .ZN(n9801) );
  AND2_X1 U13070 ( .A1(n15554), .A2(n10639), .ZN(n9802) );
  AND4_X1 U13071 ( .A1(n16591), .A2(n11422), .A3(n16588), .A4(n16612), .ZN(
        n9803) );
  NAND2_X1 U13072 ( .A1(n12415), .A2(n12403), .ZN(n9804) );
  NAND2_X1 U13073 ( .A1(n11204), .A2(n11203), .ZN(n14315) );
  NAND2_X2 U13074 ( .A1(n9963), .A2(n9962), .ZN(n16673) );
  NAND2_X1 U13075 ( .A1(n14055), .A2(n14054), .ZN(n14063) );
  AND2_X1 U13076 ( .A1(n16040), .A2(n16583), .ZN(n16028) );
  OR2_X1 U13077 ( .A1(n14364), .A2(n15839), .ZN(n9805) );
  NOR2_X1 U13078 ( .A1(n11746), .A2(n17737), .ZN(n10420) );
  AND2_X2 U13079 ( .A1(n14606), .A2(n14603), .ZN(n16317) );
  NOR2_X1 U13080 ( .A1(n19068), .A2(n19231), .ZN(n17326) );
  INV_X1 U13081 ( .A(n19444), .ZN(n20019) );
  NOR2_X1 U13082 ( .A1(n20189), .A2(n14176), .ZN(n19444) );
  AND3_X1 U13083 ( .A1(n18990), .A2(n18988), .A3(n19288), .ZN(n9806) );
  AND2_X1 U13084 ( .A1(n10561), .A2(n16588), .ZN(n9807) );
  INV_X1 U13085 ( .A(n15082), .ZN(n13430) );
  NAND2_X1 U13086 ( .A1(n10358), .A2(n10307), .ZN(n16728) );
  AND2_X1 U13087 ( .A1(n17249), .A2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n9808) );
  INV_X1 U13088 ( .A(n10014), .ZN(n10920) );
  NAND2_X1 U13089 ( .A1(n13779), .A2(n10894), .ZN(n10014) );
  INV_X1 U13090 ( .A(n10004), .ZN(n16653) );
  NAND2_X1 U13091 ( .A1(n16673), .A2(n10489), .ZN(n10004) );
  AND3_X1 U13092 ( .A1(n10714), .A2(n10715), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n9809) );
  AND2_X1 U13093 ( .A1(n15151), .A2(n15154), .ZN(n9810) );
  AND2_X1 U13094 ( .A1(n15159), .A2(n15165), .ZN(n9811) );
  AND2_X1 U13095 ( .A1(n10901), .A2(n13819), .ZN(n9812) );
  OR2_X1 U13096 ( .A1(n19105), .A2(n19144), .ZN(n9813) );
  INV_X1 U13097 ( .A(n10225), .ZN(n11443) );
  NAND2_X1 U13098 ( .A1(n16543), .A2(n16550), .ZN(n10225) );
  AND4_X1 U13099 ( .A1(n14097), .A2(n14096), .A3(n14095), .A4(n14094), .ZN(
        n9814) );
  AND3_X1 U13100 ( .A1(n10860), .A2(n10859), .A3(n10858), .ZN(n9815) );
  AND2_X1 U13101 ( .A1(n11967), .A2(n11966), .ZN(n9816) );
  AND2_X1 U13102 ( .A1(n10098), .A2(n10100), .ZN(n9817) );
  AND2_X1 U13103 ( .A1(n16596), .A2(n16841), .ZN(n9818) );
  AND2_X1 U13104 ( .A1(n11402), .A2(n11436), .ZN(n9819) );
  AND2_X1 U13105 ( .A1(n9762), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n9820) );
  OR2_X1 U13106 ( .A1(n15532), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n9821) );
  INV_X1 U13107 ( .A(n11143), .ZN(n10240) );
  INV_X1 U13108 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10224) );
  OR2_X1 U13109 ( .A1(n20884), .A2(n11083), .ZN(n9822) );
  AND2_X1 U13110 ( .A1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n9823) );
  AND2_X1 U13111 ( .A1(n10958), .A2(n10959), .ZN(n9824) );
  INV_X1 U13112 ( .A(n10484), .ZN(n10483) );
  NAND2_X1 U13113 ( .A1(n9836), .A2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10484) );
  NAND3_X1 U13114 ( .A1(n14161), .A2(n14160), .A3(n10459), .ZN(n9825) );
  OR2_X1 U13115 ( .A1(n11453), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n9826) );
  AND2_X1 U13116 ( .A1(n16756), .A2(n11361), .ZN(n9827) );
  AOI21_X1 U13117 ( .B1(n10556), .B2(n10554), .A(n10553), .ZN(n10552) );
  AND2_X1 U13118 ( .A1(n12654), .A2(n13318), .ZN(n9828) );
  NOR2_X1 U13119 ( .A1(n12567), .A2(n12566), .ZN(n9829) );
  INV_X1 U13120 ( .A(n14281), .ZN(n11171) );
  AND2_X1 U13121 ( .A1(n11170), .A2(n11169), .ZN(n14281) );
  OR3_X1 U13122 ( .A1(n11763), .A2(n11766), .A3(n10431), .ZN(n9830) );
  AND2_X1 U13123 ( .A1(n10894), .A2(n13819), .ZN(n9831) );
  OR2_X1 U13124 ( .A1(n10548), .A2(n10238), .ZN(n9833) );
  NAND2_X1 U13125 ( .A1(n16054), .A2(n9774), .ZN(n16012) );
  INV_X1 U13126 ( .A(n10555), .ZN(n10554) );
  NAND2_X1 U13127 ( .A1(n16676), .A2(n16662), .ZN(n10555) );
  AND2_X1 U13128 ( .A1(n12657), .A2(n12656), .ZN(n9834) );
  NOR2_X1 U13129 ( .A1(n10596), .A2(n13782), .ZN(n9835) );
  AND2_X1 U13130 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n9836) );
  NAND2_X1 U13131 ( .A1(n11421), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n16612) );
  INV_X1 U13132 ( .A(n19185), .ZN(n19063) );
  NOR2_X1 U13133 ( .A1(n14315), .A2(n10540), .ZN(n12105) );
  INV_X1 U13134 ( .A(n10217), .ZN(n10216) );
  NAND2_X1 U13135 ( .A1(n10218), .A2(n9768), .ZN(n10217) );
  OR3_X1 U13136 ( .A1(n12015), .A2(n12014), .A3(n12013), .ZN(P3_U2640) );
  AND2_X1 U13137 ( .A1(n14762), .A2(n12100), .ZN(n9838) );
  AND3_X1 U13138 ( .A1(n16714), .A2(n16722), .A3(n16741), .ZN(n9839) );
  AND3_X1 U13139 ( .A1(n16654), .A2(n16662), .A3(n16647), .ZN(n9840) );
  AND3_X1 U13140 ( .A1(n12589), .A2(n12588), .A3(n10436), .ZN(n9841) );
  AND2_X1 U13141 ( .A1(n9731), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9842) );
  INV_X1 U13142 ( .A(n10405), .ZN(n10234) );
  AND2_X1 U13143 ( .A1(n11494), .A2(n9769), .ZN(n9843) );
  INV_X1 U13144 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17737) );
  AND2_X1 U13145 ( .A1(n10215), .A2(n13498), .ZN(n9844) );
  AND2_X1 U13146 ( .A1(n10498), .A2(n13379), .ZN(n9845) );
  AND2_X1 U13147 ( .A1(n17254), .A2(n17256), .ZN(n9846) );
  INV_X1 U13148 ( .A(n16524), .ZN(n10137) );
  AND2_X1 U13149 ( .A1(n9967), .A2(n10488), .ZN(n9847) );
  INV_X1 U13150 ( .A(n19547), .ZN(n14012) );
  AND3_X1 U13151 ( .A1(n11925), .A2(n11924), .A3(n11923), .ZN(n19547) );
  AND2_X1 U13152 ( .A1(n9754), .A2(n11553), .ZN(n9848) );
  AND2_X1 U13153 ( .A1(n10303), .A2(n10305), .ZN(n9849) );
  NOR2_X1 U13154 ( .A1(n14973), .A2(n10653), .ZN(n9850) );
  NAND2_X1 U13155 ( .A1(n15554), .A2(n15758), .ZN(n9851) );
  INV_X1 U13156 ( .A(n10624), .ZN(n10400) );
  AND2_X1 U13157 ( .A1(n9791), .A2(n16577), .ZN(n10624) );
  INV_X1 U13158 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n20157) );
  INV_X1 U13159 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10260) );
  INV_X1 U13160 ( .A(n10204), .ZN(n10203) );
  NAND2_X1 U13161 ( .A1(n10207), .A2(n22065), .ZN(n10204) );
  NAND2_X1 U13162 ( .A1(n11143), .A2(n11142), .ZN(n16729) );
  INV_X1 U13163 ( .A(n12884), .ZN(n13232) );
  INV_X1 U13164 ( .A(n12342), .ZN(n13874) );
  INV_X2 U13165 ( .A(n21285), .ZN(n21298) );
  NAND2_X1 U13166 ( .A1(n11516), .A2(n11515), .ZN(n13811) );
  NAND2_X1 U13167 ( .A1(n11172), .A2(n11171), .ZN(n14258) );
  NAND2_X1 U13168 ( .A1(n11155), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11727) );
  NOR2_X1 U13169 ( .A1(n11158), .A2(n10527), .ZN(n14216) );
  NOR2_X1 U13170 ( .A1(n14147), .A2(n10568), .ZN(n14326) );
  AND2_X1 U13171 ( .A1(n14271), .A2(n10606), .ZN(n14322) );
  NAND2_X1 U13172 ( .A1(n13811), .A2(n13810), .ZN(n13809) );
  NAND2_X1 U13173 ( .A1(n14994), .A2(n10513), .ZN(n14944) );
  AND2_X1 U13174 ( .A1(n18715), .A2(n10255), .ZN(n9852) );
  OR2_X1 U13175 ( .A1(n11758), .A2(n11154), .ZN(n9853) );
  OR2_X1 U13176 ( .A1(n11758), .A2(n10430), .ZN(n9854) );
  NOR2_X1 U13177 ( .A1(n16344), .A2(n16343), .ZN(n10604) );
  NOR2_X1 U13178 ( .A1(n11737), .A2(n10432), .ZN(n11732) );
  AND2_X1 U13179 ( .A1(n13976), .A2(n13975), .ZN(n20020) );
  AND2_X1 U13180 ( .A1(n10513), .A2(n10512), .ZN(n9855) );
  OAI21_X1 U13181 ( .B1(n16139), .B2(n11300), .A(n16924), .ZN(n16647) );
  NAND2_X1 U13182 ( .A1(n10475), .A2(n10472), .ZN(n11799) );
  NOR2_X1 U13183 ( .A1(n14276), .A2(n10531), .ZN(n14346) );
  AND2_X1 U13184 ( .A1(n13431), .A2(n10505), .ZN(n9856) );
  AND2_X1 U13185 ( .A1(n14381), .A2(n9775), .ZN(n9857) );
  INV_X1 U13186 ( .A(n11372), .ZN(n10622) );
  INV_X1 U13187 ( .A(n11392), .ZN(n10636) );
  OAI211_X1 U13188 ( .C1(n11478), .C2(n11464), .A(n11487), .B(n11463), .ZN(
        n13791) );
  AND2_X1 U13189 ( .A1(n11673), .A2(n10583), .ZN(n9858) );
  AND2_X1 U13190 ( .A1(n10606), .A2(n14323), .ZN(n9859) );
  XNOR2_X1 U13191 ( .A(n12546), .B(n15756), .ZN(n15834) );
  NAND2_X1 U13192 ( .A1(n20250), .A2(n11763), .ZN(n16074) );
  NAND2_X1 U13193 ( .A1(n14092), .A2(n20179), .ZN(n10253) );
  NOR2_X1 U13194 ( .A1(n14904), .A2(n10499), .ZN(n14847) );
  AND2_X1 U13195 ( .A1(n14994), .A2(n14982), .ZN(n14959) );
  AND2_X1 U13196 ( .A1(n11172), .A2(n10525), .ZN(n14337) );
  NOR2_X1 U13197 ( .A1(n11799), .A2(n18953), .ZN(n11795) );
  AND2_X1 U13198 ( .A1(n16588), .A2(n12095), .ZN(n9860) );
  NAND2_X1 U13199 ( .A1(n21365), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12881) );
  INV_X1 U13200 ( .A(n12881), .ZN(n12930) );
  NOR2_X1 U13201 ( .A1(n11758), .A2(n10426), .ZN(n11764) );
  NOR2_X1 U13202 ( .A1(n11758), .A2(n10428), .ZN(n11728) );
  NAND2_X1 U13203 ( .A1(n14277), .A2(n11192), .ZN(n14309) );
  OR2_X1 U13204 ( .A1(n11654), .A2(n11653), .ZN(n9861) );
  AND2_X1 U13205 ( .A1(n16647), .A2(n14763), .ZN(n9862) );
  NOR2_X1 U13206 ( .A1(n16551), .A2(n10158), .ZN(n9863) );
  INV_X1 U13207 ( .A(n14147), .ZN(n10567) );
  INV_X1 U13208 ( .A(n19388), .ZN(n10011) );
  NAND2_X1 U13209 ( .A1(n9978), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n19086) );
  INV_X1 U13210 ( .A(n19086), .ZN(n10281) );
  AND2_X1 U13211 ( .A1(n9774), .A2(n10538), .ZN(n9864) );
  AND2_X1 U13212 ( .A1(n9855), .A2(n10511), .ZN(n9865) );
  AND4_X1 U13213 ( .A1(n16382), .A2(n14320), .A3(n14319), .A4(n14345), .ZN(
        n9866) );
  INV_X1 U13214 ( .A(n12512), .ZN(n10088) );
  INV_X1 U13215 ( .A(n10604), .ZN(n10603) );
  AND2_X1 U13216 ( .A1(n19063), .A2(n19263), .ZN(n9867) );
  NAND2_X1 U13217 ( .A1(n11232), .A2(n10333), .ZN(n16024) );
  AND2_X1 U13218 ( .A1(n11288), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n11432) );
  NAND2_X1 U13219 ( .A1(n11228), .A2(n11227), .ZN(n9868) );
  NOR2_X1 U13220 ( .A1(n16307), .A2(n10615), .ZN(n9869) );
  AND2_X1 U13221 ( .A1(n11494), .A2(n11500), .ZN(n9870) );
  NAND2_X1 U13222 ( .A1(n11037), .A2(n11022), .ZN(n9871) );
  NAND2_X1 U13223 ( .A1(n11153), .A2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11737) );
  INV_X1 U13224 ( .A(n10273), .ZN(n15177) );
  NAND2_X1 U13225 ( .A1(n12722), .A2(n10275), .ZN(n10273) );
  AND2_X1 U13226 ( .A1(n11300), .A2(n11080), .ZN(n9872) );
  NAND2_X1 U13227 ( .A1(n11188), .A2(n11187), .ZN(n14276) );
  INV_X1 U13228 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n11734) );
  AND2_X1 U13229 ( .A1(n9765), .A2(n13409), .ZN(n9873) );
  AND2_X1 U13230 ( .A1(n17167), .A2(n9731), .ZN(n9874) );
  AND2_X1 U13231 ( .A1(n18676), .A2(n10259), .ZN(n9875) );
  AND2_X1 U13232 ( .A1(n20171), .A2(n13980), .ZN(n9876) );
  INV_X1 U13233 ( .A(n16749), .ZN(n10058) );
  AND2_X1 U13234 ( .A1(n9775), .A2(n16362), .ZN(n9877) );
  OR2_X1 U13235 ( .A1(n11452), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n9878) );
  INV_X1 U13236 ( .A(n13267), .ZN(n13302) );
  INV_X1 U13237 ( .A(n13302), .ZN(n13526) );
  NOR2_X2 U13238 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n13267) );
  INV_X1 U13239 ( .A(n17320), .ZN(n10450) );
  INV_X1 U13240 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20002) );
  AND2_X1 U13241 ( .A1(n11795), .A2(n9773), .ZN(n9880) );
  AND2_X1 U13242 ( .A1(n13409), .A2(n9752), .ZN(n9881) );
  NAND2_X1 U13243 ( .A1(n12092), .A2(n21118), .ZN(n17101) );
  INV_X1 U13244 ( .A(n17101), .ZN(n17748) );
  NOR2_X1 U13245 ( .A1(n14075), .A2(n14074), .ZN(n14073) );
  NAND3_X1 U13246 ( .A1(n11504), .A2(n11503), .A3(n11502), .ZN(n9882) );
  INV_X1 U13247 ( .A(n16263), .ZN(n10190) );
  INV_X1 U13248 ( .A(n12331), .ZN(n13133) );
  BUF_X1 U13249 ( .A(n13384), .Z(n14793) );
  OR2_X1 U13250 ( .A1(n10775), .A2(n10774), .ZN(n11501) );
  INV_X1 U13251 ( .A(n11501), .ZN(n10121) );
  INV_X1 U13252 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n10429) );
  NAND2_X1 U13253 ( .A1(n13027), .A2(n13026), .ZN(n9883) );
  INV_X1 U13254 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n22107) );
  INV_X1 U13255 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n18164) );
  NAND2_X1 U13256 ( .A1(n12754), .A2(n12753), .ZN(n9884) );
  AND2_X1 U13257 ( .A1(n10462), .A2(n10460), .ZN(n9885) );
  OR2_X1 U13258 ( .A1(n19280), .A2(n19295), .ZN(n9886) );
  AND2_X1 U13259 ( .A1(n10258), .A2(n10257), .ZN(n9887) );
  OR2_X1 U13260 ( .A1(n11801), .A2(n10476), .ZN(n9888) );
  OR2_X1 U13261 ( .A1(n10289), .A2(n17258), .ZN(n9889) );
  INV_X1 U13262 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n10263) );
  INV_X1 U13263 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n10077) );
  INV_X1 U13264 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n10460) );
  INV_X1 U13265 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n10470) );
  NAND2_X1 U13266 ( .A1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n18244) );
  INV_X1 U13267 ( .A(n18244), .ZN(n10078) );
  INV_X1 U13268 ( .A(n20227), .ZN(n21006) );
  AND2_X1 U13269 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n17641), .ZN(n20227) );
  INV_X1 U13270 ( .A(n16314), .ZN(n10615) );
  AND2_X1 U13271 ( .A1(n18206), .A2(n9797), .ZN(n9890) );
  AND2_X1 U13272 ( .A1(n15677), .A2(n15672), .ZN(n9891) );
  AND2_X1 U13273 ( .A1(n10489), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n9892) );
  OR2_X1 U13274 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n9893) );
  AND2_X1 U13275 ( .A1(n18206), .A2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n9894) );
  AND2_X1 U13276 ( .A1(n11795), .A2(n10469), .ZN(n9895) );
  AND2_X1 U13277 ( .A1(n10489), .A2(n16865), .ZN(n9896) );
  AND2_X1 U13278 ( .A1(n13305), .A2(n21819), .ZN(n21328) );
  INV_X1 U13279 ( .A(n21328), .ZN(n17671) );
  AND2_X1 U13280 ( .A1(n10523), .A2(n9780), .ZN(n9897) );
  AND2_X1 U13281 ( .A1(n12082), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n9898) );
  AND2_X1 U13282 ( .A1(n21132), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n14056) );
  INV_X1 U13283 ( .A(n14056), .ZN(n10588) );
  INV_X1 U13284 ( .A(n12606), .ZN(n10640) );
  INV_X1 U13285 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16667) );
  INV_X1 U13286 ( .A(n14760), .ZN(n14753) );
  AND2_X1 U13287 ( .A1(n16865), .A2(n10346), .ZN(n9899) );
  NOR2_X1 U13288 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n9900) );
  AND2_X1 U13289 ( .A1(n9779), .A2(n9897), .ZN(n9901) );
  INV_X1 U13290 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n18920) );
  INV_X1 U13291 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n18877) );
  INV_X1 U13292 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n10356) );
  INV_X1 U13293 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n10290) );
  NOR2_X1 U13294 ( .A1(n20044), .A2(n20053), .ZN(n18280) );
  INV_X1 U13295 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n10256) );
  INV_X1 U13296 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n10463) );
  AND3_X1 U13297 ( .A1(n15390), .A2(n15650), .A3(n15617), .ZN(n9902) );
  INV_X1 U13298 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n10416) );
  INV_X1 U13299 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n22065) );
  INV_X1 U13300 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n10095) );
  INV_X1 U13301 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n10471) );
  INV_X1 U13302 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n10055) );
  OR2_X1 U13303 ( .A1(n10640), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9903) );
  INV_X1 U13304 ( .A(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n10423) );
  AND2_X1 U13305 ( .A1(n15403), .A2(n15650), .ZN(n9904) );
  INV_X1 U13306 ( .A(n18810), .ZN(n18784) );
  NAND2_X1 U13307 ( .A1(n18687), .A2(n18810), .ZN(n18685) );
  NOR2_X1 U13308 ( .A1(n22056), .A2(n19882), .ZN(n19895) );
  OR2_X1 U13309 ( .A1(n19565), .A2(n19830), .ZN(n19882) );
  NAND4_X1 U13310 ( .A1(n10808), .A2(n10806), .A3(n10805), .A4(n10807), .ZN(
        n9906) );
  NAND4_X1 U13311 ( .A1(n10812), .A2(n10810), .A3(n10809), .A4(n10811), .ZN(
        n9908) );
  NAND3_X1 U13312 ( .A1(n11721), .A2(n11277), .A3(n12088), .ZN(n9946) );
  NAND2_X1 U13313 ( .A1(n16672), .A2(n9910), .ZN(P2_U3001) );
  NOR2_X2 U13314 ( .A1(n11317), .A2(n11334), .ZN(n10633) );
  INV_X1 U13315 ( .A(n13864), .ZN(n9922) );
  INV_X1 U13316 ( .A(n10438), .ZN(n9925) );
  AND2_X2 U13317 ( .A1(n12520), .A2(n12518), .ZN(n12513) );
  OAI211_X1 U13318 ( .C1(n9929), .C2(n10103), .A(n9928), .B(n9926), .ZN(n12518) );
  INV_X1 U13319 ( .A(n9930), .ZN(n12520) );
  NAND2_X1 U13320 ( .A1(n12444), .A2(n9927), .ZN(n9926) );
  NAND3_X1 U13321 ( .A1(n10103), .A2(n12442), .A3(n9929), .ZN(n9928) );
  INV_X1 U13322 ( .A(n12444), .ZN(n9929) );
  OAI21_X1 U13323 ( .B1(n15415), .B2(n15545), .A(n15392), .ZN(n9936) );
  NAND3_X1 U13324 ( .A1(n11104), .A2(n10666), .A3(n11103), .ZN(n9941) );
  NAND2_X1 U13325 ( .A1(n10979), .A2(n9942), .ZN(n10970) );
  NAND3_X2 U13326 ( .A1(n9946), .A2(n9944), .A3(n9943), .ZN(n10960) );
  NAND3_X1 U13327 ( .A1(n9957), .A2(n9842), .A3(n17167), .ZN(n9943) );
  NAND3_X1 U13328 ( .A1(n10897), .A2(n9969), .A3(n10896), .ZN(n9945) );
  NAND2_X1 U13329 ( .A1(n12041), .A2(n9969), .ZN(n10661) );
  NAND2_X1 U13330 ( .A1(n10364), .A2(n10060), .ZN(n9948) );
  NAND2_X2 U13331 ( .A1(n10062), .A2(n11121), .ZN(n16738) );
  NAND3_X2 U13332 ( .A1(n10064), .A2(n9731), .A3(n10903), .ZN(n13614) );
  NAND2_X2 U13333 ( .A1(n9954), .A2(n9953), .ZN(n10963) );
  AND2_X2 U13334 ( .A1(n10966), .A2(n10965), .ZN(n10979) );
  NAND2_X1 U13335 ( .A1(n10950), .A2(n10951), .ZN(n10965) );
  INV_X1 U13336 ( .A(n10951), .ZN(n9955) );
  INV_X1 U13337 ( .A(n10950), .ZN(n9956) );
  NAND2_X1 U13338 ( .A1(n9957), .A2(n9874), .ZN(n12060) );
  AND2_X1 U13339 ( .A1(n12062), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9958) );
  AND2_X2 U13340 ( .A1(n16713), .A2(n9901), .ZN(n13522) );
  OAI21_X2 U13341 ( .B1(n16686), .B2(n9961), .A(n16685), .ZN(n16744) );
  INV_X1 U13342 ( .A(n10358), .ZN(n9968) );
  NAND3_X1 U13343 ( .A1(n10358), .A2(n9967), .A3(n10307), .ZN(n9963) );
  OAI21_X2 U13344 ( .B1(n9975), .B2(n9974), .A(n9972), .ZN(n17253) );
  NAND2_X1 U13345 ( .A1(n19211), .A2(n17244), .ZN(n9975) );
  NAND2_X2 U13346 ( .A1(n9982), .A2(n12517), .ZN(n15579) );
  NAND2_X1 U13347 ( .A1(n9982), .A2(n10080), .ZN(n10090) );
  OR2_X2 U13348 ( .A1(n15896), .A2(n13827), .ZN(n9982) );
  AND2_X2 U13349 ( .A1(n10272), .A2(n10271), .ZN(n12755) );
  NAND2_X2 U13350 ( .A1(n9986), .A2(n12547), .ZN(n17662) );
  OAI21_X1 U13351 ( .B1(n13495), .B2(n21153), .A(n13315), .ZN(P1_U2968) );
  NAND2_X4 U13352 ( .A1(n12581), .A2(n12580), .ZN(n15554) );
  NAND3_X1 U13353 ( .A1(n15383), .A2(n12605), .A3(n9740), .ZN(n9997) );
  NAND2_X1 U13354 ( .A1(n9998), .A2(n10121), .ZN(n11049) );
  AND2_X1 U13355 ( .A1(n9998), .A2(n10516), .ZN(n11316) );
  NAND3_X1 U13356 ( .A1(n11256), .A2(n9999), .A3(n10931), .ZN(n10063) );
  OAI211_X1 U13357 ( .C1(n10020), .C2(n10058), .A(n10001), .B(n10000), .ZN(
        n16752) );
  NAND2_X1 U13358 ( .A1(n11351), .A2(n16749), .ZN(n10000) );
  NAND3_X1 U13359 ( .A1(n10020), .A2(n9721), .A3(n10058), .ZN(n10001) );
  NAND3_X1 U13360 ( .A1(n10528), .A2(n9744), .A3(n10526), .ZN(n14251) );
  INV_X2 U13361 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n17459) );
  NAND3_X1 U13362 ( .A1(n14155), .A2(n14156), .A3(n10008), .ZN(n10007) );
  OR2_X2 U13363 ( .A1(n17357), .A2(n17356), .ZN(n17359) );
  NOR2_X1 U13364 ( .A1(n10009), .A2(n17317), .ZN(n10012) );
  NOR2_X2 U13365 ( .A1(n19279), .A2(n10450), .ZN(n18968) );
  NAND2_X2 U13366 ( .A1(n19080), .A2(n19327), .ZN(n19279) );
  NAND2_X2 U13367 ( .A1(n19176), .A2(n17315), .ZN(n19080) );
  NAND2_X1 U13368 ( .A1(n10015), .A2(n9844), .ZN(n10213) );
  NAND2_X1 U13369 ( .A1(n12017), .A2(n10270), .ZN(n10015) );
  NAND2_X1 U13370 ( .A1(n10017), .A2(n11351), .ZN(n10016) );
  NAND2_X1 U13371 ( .A1(n10022), .A2(n10018), .ZN(n10017) );
  NAND2_X1 U13372 ( .A1(n10020), .A2(n10019), .ZN(n10018) );
  NAND3_X1 U13373 ( .A1(n10024), .A2(n10026), .A3(n9721), .ZN(n10021) );
  NOR2_X2 U13374 ( .A1(n10180), .A2(n10121), .ZN(n10023) );
  NOR2_X1 U13375 ( .A1(n9784), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n10030) );
  NAND3_X1 U13376 ( .A1(n10029), .A2(n10226), .A3(n10027), .ZN(n10045) );
  NAND3_X1 U13377 ( .A1(n9761), .A2(n16550), .A3(n16543), .ZN(n10031) );
  INV_X1 U13378 ( .A(n10633), .ZN(n11310) );
  NAND2_X1 U13379 ( .A1(n13779), .A2(n10875), .ZN(n10892) );
  NAND2_X1 U13380 ( .A1(n10894), .A2(n10900), .ZN(n10906) );
  XNOR2_X1 U13381 ( .A(n10875), .B(n10900), .ZN(n12030) );
  NOR2_X1 U13382 ( .A1(n11060), .A2(n10035), .ZN(n10041) );
  NAND4_X1 U13383 ( .A1(n10039), .A2(n10038), .A3(n10037), .A4(n10036), .ZN(
        n10035) );
  INV_X1 U13384 ( .A(n11064), .ZN(n10042) );
  INV_X1 U13385 ( .A(n11061), .ZN(n10044) );
  INV_X1 U13386 ( .A(n11063), .ZN(n10043) );
  NAND3_X1 U13387 ( .A1(n10041), .A2(n11065), .A3(n10040), .ZN(n10120) );
  NAND2_X1 U13388 ( .A1(n10045), .A2(n10228), .ZN(n10155) );
  AOI21_X1 U13389 ( .B1(n9784), .B2(n10402), .A(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n10046) );
  OAI21_X1 U13390 ( .B1(n10405), .B2(n10402), .A(n9784), .ZN(n16563) );
  OAI21_X1 U13391 ( .B1(n11456), .B2(n10050), .A(n10048), .ZN(n10051) );
  NOR2_X2 U13392 ( .A1(n12730), .A2(n21194), .ZN(n12771) );
  NOR2_X2 U13393 ( .A1(n13215), .A2(n13214), .ZN(n13268) );
  OAI21_X1 U13394 ( .B1(n9721), .B2(n10058), .A(n10056), .ZN(n10060) );
  INV_X1 U13395 ( .A(n11312), .ZN(n10059) );
  XNOR2_X2 U13396 ( .A(n11351), .B(n11346), .ZN(n11312) );
  NAND2_X1 U13397 ( .A1(n10059), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10364) );
  NAND2_X2 U13398 ( .A1(n10061), .A2(n16739), .ZN(n10307) );
  NAND2_X1 U13399 ( .A1(n9760), .A2(n10062), .ZN(n10061) );
  NAND2_X2 U13400 ( .A1(n16738), .A2(n22145), .ZN(n10358) );
  AND2_X1 U13401 ( .A1(n16627), .A2(n22065), .ZN(n10206) );
  XNOR2_X2 U13402 ( .A(n10067), .B(n10521), .ZN(n17098) );
  NAND2_X1 U13403 ( .A1(n12041), .A2(n12029), .ZN(n11697) );
  AND2_X2 U13404 ( .A1(n10895), .A2(n20400), .ZN(n12063) );
  NAND3_X1 U13405 ( .A1(n10239), .A2(n10358), .A3(n10307), .ZN(n16726) );
  NAND2_X1 U13406 ( .A1(n16784), .A2(n22042), .ZN(n10065) );
  NAND2_X2 U13407 ( .A1(n10066), .A2(n9780), .ZN(n16784) );
  INV_X2 U13408 ( .A(n16556), .ZN(n10066) );
  NAND2_X2 U13409 ( .A1(n16713), .A2(n9779), .ZN(n16556) );
  NAND2_X2 U13410 ( .A1(n16726), .A2(n11143), .ZN(n16713) );
  NAND3_X1 U13411 ( .A1(n10074), .A2(n10073), .A3(n17960), .ZN(n10072) );
  NAND3_X1 U13412 ( .A1(n10078), .A2(n10076), .A3(
        P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n10079) );
  INV_X1 U13413 ( .A(n10079), .ZN(n18206) );
  NAND2_X1 U13414 ( .A1(n14071), .A2(n14072), .ZN(n10092) );
  NAND2_X1 U13415 ( .A1(n10086), .A2(n12512), .ZN(n10096) );
  NAND2_X1 U13416 ( .A1(n10087), .A2(n12623), .ZN(n10086) );
  XNOR2_X2 U13417 ( .A(n15893), .B(n12513), .ZN(n15896) );
  NAND3_X1 U13418 ( .A1(n10093), .A2(n10089), .A3(n12545), .ZN(n15835) );
  NAND3_X1 U13419 ( .A1(n15570), .A2(n10091), .A3(n10090), .ZN(n10089) );
  NAND2_X2 U13420 ( .A1(n10092), .A2(n12544), .ZN(n15570) );
  NAND2_X1 U13421 ( .A1(n15545), .A2(n9893), .ZN(n10099) );
  NAND3_X1 U13422 ( .A1(n12445), .A2(n10263), .A3(n12427), .ZN(n10103) );
  NAND2_X2 U13423 ( .A1(n10104), .A2(n12424), .ZN(n12445) );
  NAND2_X1 U13424 ( .A1(n15415), .A2(n10106), .ZN(n10105) );
  NAND2_X1 U13425 ( .A1(n15479), .A2(n15468), .ZN(n10114) );
  OAI21_X1 U13426 ( .B1(n15478), .B2(n15480), .A(n10115), .ZN(n15469) );
  OAI21_X1 U13427 ( .B1(n15606), .B2(n21153), .A(n15379), .ZN(P1_U2971) );
  OR2_X1 U13428 ( .A1(n16878), .A2(n16737), .ZN(n10116) );
  NAND2_X2 U13429 ( .A1(n10120), .A2(n11080), .ZN(n11346) );
  INV_X1 U13430 ( .A(n10180), .ZN(n10395) );
  NAND2_X2 U13431 ( .A1(n10122), .A2(n10345), .ZN(n16712) );
  NAND2_X1 U13432 ( .A1(n16541), .A2(n10131), .ZN(n10129) );
  NAND3_X1 U13433 ( .A1(n10139), .A2(n10403), .A3(n10138), .ZN(n10276) );
  NAND3_X1 U13434 ( .A1(n16756), .A2(n10401), .A3(n11361), .ZN(n10139) );
  NAND2_X2 U13435 ( .A1(n10141), .A2(n11343), .ZN(n16756) );
  OAI21_X1 U13436 ( .B1(n13495), .B2(n15864), .A(n10142), .ZN(P1_U3000) );
  NAND2_X1 U13437 ( .A1(n17662), .A2(n9757), .ZN(n10143) );
  NAND2_X1 U13438 ( .A1(n9841), .A2(n10143), .ZN(n10170) );
  OAI21_X2 U13439 ( .B1(n12670), .B2(n13827), .A(n12507), .ZN(n12546) );
  INV_X1 U13440 ( .A(n12548), .ZN(n10144) );
  NAND2_X1 U13441 ( .A1(n14208), .A2(n14207), .ZN(n14213) );
  NAND2_X1 U13442 ( .A1(n14211), .A2(n14062), .ZN(n14210) );
  INV_X1 U13443 ( .A(n14366), .ZN(n14381) );
  NAND2_X2 U13444 ( .A1(n10147), .A2(n10601), .ZN(n16337) );
  NAND3_X1 U13445 ( .A1(n16701), .A2(n16691), .A3(n9839), .ZN(n12097) );
  NAND3_X1 U13446 ( .A1(n11426), .A2(n11425), .A3(n10624), .ZN(n10156) );
  AND2_X2 U13447 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10693) );
  INV_X1 U13448 ( .A(n17313), .ZN(n17310) );
  NAND2_X1 U13449 ( .A1(n10276), .A2(n10623), .ZN(n10159) );
  INV_X1 U13450 ( .A(n10399), .ZN(n11352) );
  OR2_X1 U13451 ( .A1(n10399), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11361) );
  NAND2_X1 U13452 ( .A1(n10399), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n16685) );
  OAI21_X1 U13453 ( .B1(n10455), .B2(n12289), .A(n12531), .ZN(n12539) );
  NAND2_X1 U13454 ( .A1(n15462), .A2(n10178), .ZN(n10176) );
  NAND2_X1 U13455 ( .A1(n15462), .A2(n9755), .ZN(n10177) );
  NAND2_X1 U13456 ( .A1(n10517), .A2(n10180), .ZN(n10516) );
  OAI21_X2 U13457 ( .B1(n11009), .B2(n11008), .A(n9871), .ZN(n10180) );
  OAI21_X1 U13458 ( .B1(n11091), .B2(n10992), .A(n10181), .ZN(n10993) );
  NAND4_X1 U13459 ( .A1(n17744), .A2(n17146), .A3(
        P2_INSTQUEUE_REG_7__1__SCAN_IN), .A4(n10183), .ZN(n10181) );
  NAND3_X1 U13460 ( .A1(n17730), .A2(n11048), .A3(n10521), .ZN(n10520) );
  NAND2_X1 U13461 ( .A1(n11316), .A2(n10188), .ZN(n10186) );
  NAND2_X1 U13462 ( .A1(n10191), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12419) );
  NAND2_X1 U13463 ( .A1(n10191), .A2(n10262), .ZN(n10261) );
  NAND4_X1 U13464 ( .A1(n12407), .A2(n12315), .A3(n12314), .A4(n12316), .ZN(
        n10191) );
  AND2_X2 U13465 ( .A1(n10192), .A2(n12134), .ZN(n12391) );
  AND2_X2 U13466 ( .A1(n10192), .A2(n10446), .ZN(n12331) );
  AND2_X4 U13467 ( .A1(n12122), .A2(n10192), .ZN(n12390) );
  NAND2_X1 U13468 ( .A1(n14061), .A2(n14060), .ZN(n14211) );
  NAND2_X2 U13469 ( .A1(n16356), .A2(n16358), .ZN(n16352) );
  OAI211_X1 U13470 ( .C1(n14724), .C2(n17101), .A(n13524), .B(n9709), .ZN(
        P2_U3015) );
  NAND2_X1 U13471 ( .A1(n16617), .A2(n10207), .ZN(n10205) );
  INV_X1 U13472 ( .A(n10200), .ZN(n10202) );
  OAI21_X1 U13473 ( .B1(n16653), .B2(n10204), .A(n10201), .ZN(n10200) );
  NOR2_X1 U13474 ( .A1(n16617), .A2(n10206), .ZN(n16904) );
  NAND3_X1 U13475 ( .A1(n11014), .A2(n11015), .A3(n11016), .ZN(n10212) );
  NAND3_X1 U13476 ( .A1(n12017), .A2(n10270), .A3(n13504), .ZN(n10214) );
  NAND2_X1 U13477 ( .A1(n11382), .A2(n10218), .ZN(n11398) );
  NAND2_X1 U13478 ( .A1(n11382), .A2(n10635), .ZN(n11378) );
  NAND2_X1 U13479 ( .A1(n11371), .A2(n11428), .ZN(n11427) );
  AND2_X2 U13480 ( .A1(n10394), .A2(n14123), .ZN(n14504) );
  INV_X1 U13481 ( .A(n11454), .ZN(n10228) );
  INV_X1 U13482 ( .A(n11316), .ZN(n11315) );
  OAI21_X1 U13483 ( .B1(n10234), .B2(n12097), .A(n12096), .ZN(n16678) );
  OAI22_X1 U13484 ( .A1(n10548), .A2(n10237), .B1(n10550), .B2(n12099), .ZN(
        n10236) );
  NOR2_X1 U13485 ( .A1(n10248), .A2(n11981), .ZN(n14030) );
  NAND3_X1 U13486 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(P3_EAX_REG_0__SCAN_IN), 
        .A3(P3_EAX_REG_6__SCAN_IN), .ZN(n10251) );
  AND2_X2 U13487 ( .A1(n17459), .A2(n10260), .ZN(n14031) );
  NAND2_X1 U13488 ( .A1(n10261), .A2(n12317), .ZN(n12412) );
  NAND2_X1 U13489 ( .A1(n12708), .A2(n21908), .ZN(n12374) );
  NAND2_X1 U13490 ( .A1(n10264), .A2(n10267), .ZN(n15407) );
  NAND3_X1 U13491 ( .A1(n10268), .A2(n15545), .A3(n10265), .ZN(n10264) );
  INV_X1 U13492 ( .A(n15415), .ZN(n10265) );
  AND3_X2 U13493 ( .A1(n12722), .A2(n10274), .A3(n10275), .ZN(n10271) );
  NAND2_X1 U13494 ( .A1(n15893), .A2(n12513), .ZN(n12514) );
  NOR2_X1 U13495 ( .A1(n10281), .A2(n17257), .ZN(n19450) );
  OAI21_X1 U13496 ( .B1(n10283), .B2(n17272), .A(n17274), .ZN(n10282) );
  NOR2_X1 U13497 ( .A1(n17633), .A2(n19185), .ZN(n17272) );
  NOR2_X1 U13498 ( .A1(n17273), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10283) );
  NAND2_X1 U13499 ( .A1(n17276), .A2(n17275), .ZN(n10284) );
  NAND2_X1 U13500 ( .A1(n17334), .A2(n17270), .ZN(n17271) );
  INV_X1 U13501 ( .A(n17270), .ZN(n10286) );
  NAND2_X1 U13502 ( .A1(n17294), .A2(n17299), .ZN(n17228) );
  OR2_X1 U13503 ( .A1(n17295), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17299) );
  INV_X1 U13504 ( .A(n12638), .ZN(n10299) );
  NAND2_X1 U13505 ( .A1(n10300), .A2(n10298), .ZN(n12652) );
  NAND3_X1 U13506 ( .A1(n12632), .A2(n12631), .A3(n12643), .ZN(n10300) );
  NAND2_X1 U13507 ( .A1(n10302), .A2(n9849), .ZN(n13328) );
  OAI21_X1 U13508 ( .B1(n9782), .B2(n12660), .A(n12665), .ZN(n10304) );
  INV_X1 U13509 ( .A(n13327), .ZN(n10305) );
  NOR2_X2 U13510 ( .A1(n15630), .A2(n15617), .ZN(n15616) );
  NAND3_X1 U13511 ( .A1(n10712), .A2(n10713), .A3(n10308), .ZN(n10319) );
  NOR2_X1 U13512 ( .A1(n10310), .A2(n10309), .ZN(n10308) );
  NAND2_X1 U13513 ( .A1(n10313), .A2(n10320), .ZN(n10310) );
  NAND2_X1 U13514 ( .A1(n14458), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n10313) );
  NAND2_X1 U13515 ( .A1(n14457), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n10312) );
  OR2_X1 U13516 ( .A1(n16712), .A2(n16849), .ZN(n10317) );
  AOI21_X1 U13517 ( .B1(n16712), .B2(n16848), .A(n10315), .ZN(n10314) );
  INV_X1 U13518 ( .A(n16712), .ZN(n10318) );
  AND2_X2 U13519 ( .A1(n16596), .A2(n10314), .ZN(n16855) );
  INV_X1 U13520 ( .A(n10317), .ZN(n16604) );
  NAND3_X1 U13521 ( .A1(n9809), .A2(n10716), .A3(n10717), .ZN(n10321) );
  CLKBUF_X1 U13522 ( .A(n10957), .Z(n10322) );
  NAND3_X1 U13523 ( .A1(n11166), .A2(n11165), .A3(n10323), .ZN(n14252) );
  NAND3_X1 U13524 ( .A1(n11182), .A2(n11181), .A3(n10324), .ZN(n14338) );
  NAND3_X1 U13525 ( .A1(n11210), .A2(n11209), .A3(n10325), .ZN(n14764) );
  NAND3_X1 U13526 ( .A1(n11220), .A2(n11219), .A3(n10326), .ZN(n12106) );
  AOI21_X1 U13527 ( .B1(n16605), .B2(n16860), .A(n16604), .ZN(n16876) );
  NAND4_X1 U13528 ( .A1(n11902), .A2(n10350), .A3(n11903), .A4(n11905), .ZN(
        n14179) );
  NAND4_X1 U13529 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(P3_EBX_REG_23__SCAN_IN), 
        .A3(P3_EBX_REG_22__SCAN_IN), .A4(P3_EBX_REG_24__SCAN_IN), .ZN(n10355)
         );
  NAND3_X1 U13530 ( .A1(n10832), .A2(n10361), .A3(n10830), .ZN(n10360) );
  INV_X1 U13531 ( .A(n20415), .ZN(n10891) );
  NOR2_X1 U13533 ( .A1(n17059), .A2(n10363), .ZN(n17061) );
  INV_X1 U13534 ( .A(n17060), .ZN(n10363) );
  NAND2_X1 U13535 ( .A1(n16751), .A2(n10364), .ZN(n16753) );
  NAND2_X1 U13536 ( .A1(n17059), .A2(n16749), .ZN(n10365) );
  NAND3_X1 U13537 ( .A1(n19547), .A2(n10373), .A3(n10372), .ZN(n11981) );
  INV_X4 U13538 ( .A(n18525), .ZN(n18390) );
  NAND2_X2 U13539 ( .A1(n11812), .A2(n14031), .ZN(n18525) );
  INV_X2 U13540 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n20146) );
  NAND2_X1 U13541 ( .A1(n19488), .A2(n10374), .ZN(n10377) );
  INV_X1 U13542 ( .A(n10378), .ZN(n19416) );
  NAND2_X1 U13543 ( .A1(n10386), .A2(n10379), .ZN(P3_U2800) );
  AOI21_X1 U13544 ( .B1(n18975), .B2(n10384), .A(n10380), .ZN(n10379) );
  INV_X2 U13545 ( .A(n18551), .ZN(n18597) );
  NOR2_X1 U13546 ( .A1(n10394), .A2(n10700), .ZN(n17138) );
  NAND3_X1 U13547 ( .A1(n10398), .A2(n11349), .A3(n11348), .ZN(n10399) );
  NAND3_X1 U13548 ( .A1(n10578), .A2(n10407), .A3(n10406), .ZN(P2_U3017) );
  AND2_X1 U13549 ( .A1(n10579), .A2(n10408), .ZN(n10407) );
  NAND3_X1 U13550 ( .A1(n10413), .A2(n10411), .A3(n10409), .ZN(n16103) );
  INV_X1 U13551 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n10417) );
  NAND3_X1 U13552 ( .A1(n10420), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A3(
        n10418), .ZN(n11743) );
  NAND3_X1 U13553 ( .A1(n10424), .A2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n11747) );
  NAND2_X1 U13554 ( .A1(n20250), .A2(n9830), .ZN(n16040) );
  INV_X1 U13555 ( .A(n12590), .ZN(n10436) );
  AND2_X2 U13556 ( .A1(n12129), .A2(n10446), .ZN(n12267) );
  NAND2_X1 U13557 ( .A1(n17262), .A2(n17261), .ZN(n19064) );
  NAND2_X1 U13558 ( .A1(n19020), .A2(n10447), .ZN(n17434) );
  NAND2_X1 U13559 ( .A1(n10451), .A2(n19224), .ZN(n10452) );
  INV_X1 U13560 ( .A(n17238), .ZN(n10451) );
  NAND3_X1 U13561 ( .A1(n10453), .A2(n17241), .A3(n10452), .ZN(n19211) );
  NAND3_X1 U13562 ( .A1(n19238), .A2(n19224), .A3(n17236), .ZN(n10453) );
  NAND2_X1 U13563 ( .A1(n12426), .A2(n21381), .ZN(n15105) );
  OR2_X2 U13564 ( .A1(n21438), .A2(n12413), .ZN(n12426) );
  NAND2_X1 U13565 ( .A1(n15462), .A2(n10457), .ZN(n15436) );
  AND2_X4 U13566 ( .A1(n18270), .A2(n11824), .ZN(n17547) );
  INV_X1 U13567 ( .A(n11801), .ZN(n10475) );
  INV_X2 U13568 ( .A(n17277), .ZN(n18227) );
  NAND2_X1 U13569 ( .A1(n10481), .A2(n18206), .ZN(n19066) );
  NAND3_X1 U13570 ( .A1(n10729), .A2(n10727), .A3(n10728), .ZN(n10485) );
  NAND4_X1 U13571 ( .A1(n10723), .A2(n10721), .A3(n10722), .A4(n10720), .ZN(
        n10486) );
  XNOR2_X2 U13572 ( .A(n10963), .B(n10487), .ZN(n13778) );
  NAND2_X1 U13573 ( .A1(n12445), .A2(n12427), .ZN(n13896) );
  NAND3_X1 U13574 ( .A1(n9851), .A2(n12598), .A3(n15518), .ZN(n15479) );
  NAND2_X1 U13575 ( .A1(n15422), .A2(n10492), .ZN(n10491) );
  NAND2_X1 U13576 ( .A1(n12603), .A2(n9845), .ZN(n10497) );
  NAND2_X1 U13577 ( .A1(n12603), .A2(n15545), .ZN(n12605) );
  NOR2_X1 U13578 ( .A1(n12604), .A2(n15424), .ZN(n10492) );
  NAND2_X1 U13579 ( .A1(n10497), .A2(n10494), .ZN(n15355) );
  NAND2_X1 U13580 ( .A1(n15422), .A2(n10495), .ZN(n10494) );
  NAND2_X1 U13581 ( .A1(n13431), .A2(n9767), .ZN(n15014) );
  NAND3_X1 U13582 ( .A1(n9765), .A2(n15142), .A3(n13409), .ZN(n15081) );
  INV_X1 U13583 ( .A(n14814), .ZN(n14817) );
  NOR2_X2 U13584 ( .A1(n11003), .A2(n9727), .ZN(n11052) );
  NAND4_X1 U13585 ( .A1(n11034), .A2(n11033), .A3(n11031), .A4(n11032), .ZN(
        n10518) );
  NAND2_X1 U13586 ( .A1(n11172), .A2(n10524), .ZN(n14275) );
  INV_X1 U13587 ( .A(n11158), .ZN(n10526) );
  NAND2_X1 U13588 ( .A1(n14277), .A2(n10529), .ZN(n14316) );
  NAND3_X1 U13589 ( .A1(n10537), .A2(n15984), .A3(n10536), .ZN(n10535) );
  NAND2_X1 U13590 ( .A1(n13811), .A2(n9848), .ZN(n13919) );
  NAND2_X1 U13591 ( .A1(n11674), .A2(n10580), .ZN(n15996) );
  INV_X1 U13592 ( .A(n10868), .ZN(n14657) );
  AND3_X4 U13593 ( .A1(n10702), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10868) );
  INV_X2 U13594 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10702) );
  INV_X1 U13595 ( .A(n10585), .ZN(n10584) );
  INV_X1 U13596 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10586) );
  INV_X1 U13597 ( .A(n13804), .ZN(n10591) );
  AOI21_X1 U13598 ( .B1(n10597), .B2(n13782), .A(n10596), .ZN(n10589) );
  NAND3_X1 U13599 ( .A1(n10591), .A2(n10590), .A3(n10592), .ZN(n14049) );
  NAND2_X1 U13600 ( .A1(n10597), .A2(n13782), .ZN(n13800) );
  NOR2_X1 U13601 ( .A1(n10594), .A2(n14047), .ZN(n10593) );
  INV_X1 U13602 ( .A(n13782), .ZN(n10594) );
  INV_X1 U13603 ( .A(n10602), .ZN(n10601) );
  OAI21_X1 U13604 ( .B1(n10605), .B2(n10604), .A(n16338), .ZN(n10602) );
  OR2_X2 U13605 ( .A1(n14213), .A2(n14212), .ZN(n14271) );
  OAI21_X1 U13606 ( .B1(n14607), .B2(n16307), .A(n10608), .ZN(n10613) );
  AND2_X1 U13607 ( .A1(n16312), .A2(n10617), .ZN(n10616) );
  INV_X1 U13608 ( .A(n16307), .ZN(n10617) );
  NAND2_X1 U13609 ( .A1(n16569), .A2(n10627), .ZN(n10626) );
  OAI21_X1 U13610 ( .B1(n10746), .B2(n10747), .A(n10927), .ZN(n10628) );
  AOI22_X1 U13611 ( .A1(n10877), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n14503), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10744) );
  NAND2_X1 U13612 ( .A1(n10634), .A2(n11398), .ZN(n16139) );
  OR2_X2 U13613 ( .A1(n14905), .A2(n10644), .ZN(n14850) );
  OAI211_X1 U13614 ( .C1(n14821), .C2(n10656), .A(n10655), .B(n9763), .ZN(
        n14747) );
  NAND2_X1 U13615 ( .A1(n14821), .A2(n10659), .ZN(n10655) );
  NOR2_X2 U13616 ( .A1(n14821), .A2(n14823), .ZN(n14807) );
  INV_X1 U13617 ( .A(n13304), .ZN(n10659) );
  INV_X1 U13618 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10701) );
  INV_X2 U13619 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10750) );
  BUF_X2 U13620 ( .A(n10813), .Z(n10867) );
  NAND2_X1 U13621 ( .A1(n16227), .A2(n11511), .ZN(n13822) );
  INV_X1 U13622 ( .A(n15170), .ZN(n13409) );
  NOR2_X1 U13623 ( .A1(n16337), .A2(n14576), .ZN(n16324) );
  INV_X1 U13624 ( .A(n15081), .ZN(n13431) );
  NOR2_X1 U13625 ( .A1(n10930), .A2(n9722), .ZN(n10935) );
  NOR2_X1 U13626 ( .A1(n15598), .A2(n17647), .ZN(n14818) );
  INV_X1 U13627 ( .A(n14316), .ZN(n11204) );
  OAI21_X2 U13628 ( .B1(n14050), .B2(n14051), .A(n14055), .ZN(n21100) );
  NAND2_X1 U13629 ( .A1(n11319), .A2(n11318), .ZN(n11317) );
  AND2_X1 U13630 ( .A1(n11402), .A2(n11401), .ZN(n20220) );
  INV_X1 U13631 ( .A(n12061), .ZN(n13815) );
  INV_X1 U13632 ( .A(n13548), .ZN(n13549) );
  OAI21_X1 U13633 ( .B1(n15927), .B2(n20363), .A(n14720), .ZN(n14721) );
  CLKBUF_X1 U13634 ( .A(n12671), .Z(n21365) );
  OAI211_X1 U13635 ( .C1(n11373), .C2(n11288), .A(n11365), .B(n11363), .ZN(
        n11364) );
  NAND2_X1 U13636 ( .A1(n11373), .A2(n10669), .ZN(n11363) );
  NAND2_X1 U13637 ( .A1(n13324), .A2(n13383), .ZN(n13847) );
  CLKBUF_X1 U13638 ( .A(n13332), .Z(n14777) );
  NAND2_X1 U13639 ( .A1(n12320), .A2(n12294), .ZN(n12306) );
  NAND2_X1 U13640 ( .A1(n11467), .A2(n9731), .ZN(n10919) );
  OR2_X1 U13641 ( .A1(n13175), .A2(n12258), .ZN(n12266) );
  OR2_X1 U13642 ( .A1(n13175), .A2(n13119), .ZN(n12253) );
  OR2_X1 U13643 ( .A1(n13175), .A2(n12162), .ZN(n12163) );
  INV_X1 U13644 ( .A(n13175), .ZN(n12343) );
  XNOR2_X2 U13645 ( .A(n13508), .B(n13507), .ZN(n16394) );
  AND2_X1 U13646 ( .A1(n16324), .A2(n16327), .ZN(n14580) );
  AND2_X4 U13647 ( .A1(n12115), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12128) );
  INV_X1 U13648 ( .A(n17070), .ZN(n14751) );
  AND2_X1 U13649 ( .A1(n12092), .A2(n17775), .ZN(n17070) );
  INV_X1 U13650 ( .A(n17082), .ZN(n17738) );
  INV_X1 U13651 ( .A(n13819), .ZN(n20440) );
  AND2_X1 U13652 ( .A1(n20250), .A2(n16270), .ZN(n10662) );
  NAND2_X1 U13653 ( .A1(n15988), .A2(n16548), .ZN(n15973) );
  INV_X1 U13654 ( .A(n10922), .ZN(n11277) );
  AND3_X1 U13655 ( .A1(n12905), .A2(n12904), .A3(n12903), .ZN(n10663) );
  NOR2_X1 U13656 ( .A1(n21338), .A2(n21585), .ZN(n10664) );
  INV_X1 U13657 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n19165) );
  AND4_X1 U13658 ( .A1(n11102), .A2(n11101), .A3(n11100), .A4(n11099), .ZN(
        n10666) );
  AND2_X1 U13659 ( .A1(n11717), .A2(n11716), .ZN(n10667) );
  XNOR2_X1 U13660 ( .A(n15928), .B(n15937), .ZN(n10668) );
  AND2_X1 U13661 ( .A1(n11288), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n10669) );
  INV_X1 U13662 ( .A(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n11738) );
  INV_X1 U13663 ( .A(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n18610) );
  NOR2_X1 U13664 ( .A1(n17796), .A2(n20945), .ZN(n10671) );
  AND2_X1 U13665 ( .A1(n17296), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10672) );
  AND2_X1 U13666 ( .A1(n20941), .A2(n11283), .ZN(n20370) );
  AND2_X1 U13667 ( .A1(n16723), .A2(n16742), .ZN(n10673) );
  INV_X1 U13668 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16942) );
  NOR2_X1 U13669 ( .A1(n15184), .A2(n15171), .ZN(n10674) );
  NOR2_X1 U13670 ( .A1(n21698), .A2(n21807), .ZN(n10675) );
  NOR2_X1 U13671 ( .A1(n21698), .A2(n21524), .ZN(n10676) );
  INV_X1 U13672 ( .A(n16788), .ZN(n11149) );
  AND2_X1 U13673 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(P3_EBX_REG_4__SCAN_IN), 
        .ZN(n10677) );
  INV_X1 U13674 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n21959) );
  INV_X1 U13675 ( .A(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n19755) );
  INV_X1 U13676 ( .A(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n19758) );
  INV_X1 U13677 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n11305) );
  INV_X1 U13678 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12611) );
  NAND2_X1 U13679 ( .A1(n15554), .A2(n15798), .ZN(n15517) );
  INV_X1 U13680 ( .A(n15517), .ZN(n12596) );
  INV_X1 U13681 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n21011) );
  NAND2_X1 U13682 ( .A1(n11288), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n10678) );
  INV_X1 U13683 ( .A(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12762) );
  INV_X1 U13684 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n11301) );
  INV_X1 U13685 ( .A(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11951) );
  NOR2_X1 U13686 ( .A1(n21698), .A2(n21668), .ZN(n10679) );
  INV_X1 U13687 ( .A(n16550), .ZN(n11442) );
  INV_X1 U13688 ( .A(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n22105) );
  AND3_X1 U13689 ( .A1(n12018), .A2(n11452), .A3(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n10680) );
  INV_X1 U13690 ( .A(n19004), .ZN(n11806) );
  INV_X1 U13691 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n11154) );
  INV_X1 U13692 ( .A(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n21977) );
  AND2_X1 U13693 ( .A1(n20240), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10681) );
  INV_X1 U13694 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n15751) );
  INV_X1 U13695 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16695) );
  INV_X1 U13696 ( .A(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n18476) );
  INV_X1 U13697 ( .A(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n21980) );
  INV_X2 U13698 ( .A(n20185), .ZN(n20184) );
  INV_X1 U13699 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n17256) );
  INV_X1 U13700 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n21704) );
  NOR2_X2 U13701 ( .A1(n21916), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n13612) );
  OR2_X1 U13702 ( .A1(n13626), .A2(n9736), .ZN(n16762) );
  INV_X1 U13703 ( .A(n16762), .ZN(n20357) );
  INV_X1 U13704 ( .A(n16737), .ZN(n11457) );
  AND2_X1 U13705 ( .A1(n13777), .A2(n17793), .ZN(n16363) );
  INV_X1 U13706 ( .A(n16363), .ZN(n16386) );
  INV_X2 U13707 ( .A(n21141), .ZN(n21140) );
  NAND2_X2 U13708 ( .A1(n13574), .A2(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n14329)
         );
  NAND3_X1 U13709 ( .A1(n11624), .A2(n11623), .A3(n11622), .ZN(n10684) );
  INV_X1 U13710 ( .A(n15296), .ZN(n15291) );
  NAND2_X2 U13711 ( .A1(n15296), .A2(n13859), .ZN(n15299) );
  AND2_X1 U13712 ( .A1(n10968), .A2(n10967), .ZN(n10685) );
  INV_X1 U13713 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n11279) );
  INV_X1 U13714 ( .A(n13082), .ZN(n13245) );
  NAND2_X1 U13715 ( .A1(n12308), .A2(n13350), .ZN(n12309) );
  NOR2_X1 U13716 ( .A1(n12327), .A2(n13346), .ZN(n12315) );
  INV_X1 U13717 ( .A(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13172) );
  AOI21_X1 U13718 ( .B1(n9732), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A(
        n14126), .ZN(n10864) );
  AND2_X1 U13719 ( .A1(n12025), .A2(n13819), .ZN(n10893) );
  NAND2_X1 U13720 ( .A1(n10900), .A2(n20415), .ZN(n10901) );
  OAI22_X1 U13721 ( .A1(n12379), .A2(n12983), .B1(n13175), .B2(n13172), .ZN(
        n12226) );
  INV_X1 U13722 ( .A(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12867) );
  INV_X1 U13723 ( .A(n12391), .ZN(n13082) );
  OR2_X1 U13724 ( .A1(n12500), .A2(n12499), .ZN(n12505) );
  INV_X1 U13725 ( .A(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12184) );
  AOI21_X1 U13726 ( .B1(n9732), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10850) );
  AOI21_X1 U13727 ( .B1(n9732), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A(
        n14126), .ZN(n10845) );
  NOR2_X1 U13728 ( .A1(n12226), .A2(n12225), .ZN(n12230) );
  INV_X1 U13729 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12717) );
  AND4_X1 U13730 ( .A1(n12339), .A2(n12338), .A3(n12337), .A4(n12336), .ZN(
        n12354) );
  NOR2_X1 U13731 ( .A1(n12293), .A2(n21908), .ZN(n12441) );
  OR2_X1 U13732 ( .A1(n13175), .A2(n12192), .ZN(n12196) );
  NOR2_X1 U13733 ( .A1(n10793), .A2(n10792), .ZN(n10794) );
  NAND2_X1 U13734 ( .A1(n14458), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n10724) );
  INV_X1 U13735 ( .A(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n18448) );
  AND4_X1 U13736 ( .A1(n12234), .A2(n12233), .A3(n12232), .A4(n12231), .ZN(
        n12235) );
  INV_X1 U13737 ( .A(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13120) );
  OR4_X1 U13738 ( .A1(n13139), .A2(n13138), .A3(n13137), .A4(n13136), .ZN(
        n13145) );
  NOR2_X1 U13739 ( .A1(n12672), .A2(n12682), .ZN(n12723) );
  NOR2_X1 U13740 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12606) );
  INV_X1 U13741 ( .A(n15516), .ZN(n12597) );
  OR2_X1 U13742 ( .A1(n13175), .A2(n12116), .ZN(n12117) );
  AND2_X1 U13743 ( .A1(n14599), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n14044) );
  INV_X1 U13744 ( .A(n14655), .ZN(n14633) );
  OR2_X1 U13745 ( .A1(n11179), .A2(n14259), .ZN(n11180) );
  INV_X1 U13746 ( .A(n16059), .ZN(n11673) );
  AND2_X1 U13747 ( .A1(n10719), .A2(n10718), .ZN(n10723) );
  INV_X1 U13748 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n11982) );
  INV_X1 U13749 ( .A(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n18612) );
  INV_X1 U13750 ( .A(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n18527) );
  OR2_X1 U13751 ( .A1(n12379), .A2(n12142), .ZN(n12143) );
  OR2_X1 U13752 ( .A1(n12379), .A2(n12800), .ZN(n12264) );
  OR2_X1 U13753 ( .A1(n12379), .A2(n12936), .ZN(n12242) );
  INV_X1 U13754 ( .A(n12954), .ZN(n12955) );
  INV_X1 U13755 ( .A(n12723), .ZN(n12884) );
  INV_X1 U13756 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n21254) );
  OR2_X1 U13757 ( .A1(n15907), .A2(n12289), .ZN(n13347) );
  OAI211_X1 U13758 ( .C1(n12654), .C2(n13092), .A(n12376), .B(n12375), .ZN(
        n12533) );
  OR2_X1 U13760 ( .A1(n12467), .A2(n12466), .ZN(n12516) );
  INV_X1 U13761 ( .A(n11505), .ZN(n11297) );
  NOR2_X1 U13762 ( .A1(n20883), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n13781) );
  INV_X1 U13763 ( .A(n14659), .ZN(n17147) );
  OR2_X1 U13764 ( .A1(n14492), .A2(n14491), .ZN(n14538) );
  INV_X1 U13765 ( .A(n11710), .ZN(n11451) );
  INV_X1 U13766 ( .A(n11514), .ZN(n11300) );
  NAND2_X1 U13767 ( .A1(n11705), .A2(n10941), .ZN(n14127) );
  OR2_X2 U13768 ( .A1(n17146), .A2(n10985), .ZN(n11001) );
  INV_X1 U13769 ( .A(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n22079) );
  INV_X1 U13770 ( .A(n18963), .ZN(n11809) );
  INV_X1 U13771 ( .A(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17478) );
  INV_X1 U13772 ( .A(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13982) );
  INV_X1 U13773 ( .A(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n18447) );
  INV_X1 U13774 ( .A(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n18454) );
  INV_X1 U13775 ( .A(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n17507) );
  AOI21_X1 U13776 ( .B1(n19521), .B2(n20174), .A(n20151), .ZN(n17173) );
  NAND2_X1 U13777 ( .A1(n12307), .A2(n12672), .ZN(n12303) );
  AND4_X1 U13778 ( .A1(n12271), .A2(n12270), .A3(n12269), .A4(n12268), .ZN(
        n12282) );
  INV_X1 U13779 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n12840) );
  OAI21_X2 U13780 ( .B1(n12690), .B2(n12881), .A(n12689), .ZN(n15181) );
  AND2_X1 U13781 ( .A1(n12579), .A2(n12623), .ZN(n12580) );
  OAI211_X1 U13782 ( .C1(n11368), .C2(P2_EBX_REG_20__SCAN_IN), .A(n11288), .B(
        P2_EBX_REG_21__SCAN_IN), .ZN(n11369) );
  INV_X1 U13783 ( .A(n16097), .ZN(n11218) );
  AND2_X1 U13784 ( .A1(n20217), .A2(n11718), .ZN(n11719) );
  INV_X1 U13785 ( .A(n14317), .ZN(n11203) );
  INV_X1 U13786 ( .A(n14310), .ZN(n11192) );
  AOI21_X1 U13787 ( .B1(n14059), .B2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n13781), .ZN(n13782) );
  INV_X1 U13788 ( .A(n14606), .ZN(n14607) );
  AND2_X1 U13789 ( .A1(n14476), .A2(n14475), .ZN(n14535) );
  AND2_X1 U13790 ( .A1(n11666), .A2(n11665), .ZN(n16100) );
  NAND2_X1 U13791 ( .A1(n13573), .A2(n13572), .ZN(n13574) );
  OAI21_X1 U13792 ( .B1(n14718), .B2(n20368), .A(n14717), .ZN(n14719) );
  INV_X1 U13793 ( .A(n10979), .ZN(n10980) );
  INV_X1 U13794 ( .A(n13496), .ZN(n13497) );
  AND2_X1 U13795 ( .A1(n11685), .A2(n11684), .ZN(n15986) );
  AND2_X1 U13796 ( .A1(n11452), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11139) );
  INV_X1 U13797 ( .A(n17774), .ZN(n12022) );
  AND2_X1 U13798 ( .A1(n20370), .A2(n14329), .ZN(n20436) );
  NOR2_X1 U13799 ( .A1(n18252), .A2(n17332), .ZN(n12009) );
  NOR2_X1 U13800 ( .A1(n20034), .A2(n12005), .ZN(n18272) );
  AND2_X1 U13801 ( .A1(n17337), .A2(n17264), .ZN(n18978) );
  AND2_X1 U13802 ( .A1(n19010), .A2(n19286), .ZN(n18990) );
  INV_X1 U13803 ( .A(n20020), .ZN(n14188) );
  INV_X1 U13804 ( .A(n17173), .ZN(n19530) );
  NAND2_X1 U13805 ( .A1(n21170), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n14797) );
  NAND2_X1 U13806 ( .A1(n13541), .A2(n13540), .ZN(n21256) );
  AND2_X1 U13807 ( .A1(n13446), .A2(n13445), .ZN(n14982) );
  INV_X1 U13808 ( .A(n15272), .ZN(n15278) );
  INV_X1 U13809 ( .A(n13860), .ZN(n13858) );
  AND2_X1 U13810 ( .A1(n15300), .A2(n17713), .ZN(n15301) );
  INV_X1 U13811 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n15432) );
  AND2_X1 U13812 ( .A1(n12930), .A2(n12929), .ZN(n15077) );
  INV_X1 U13813 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n15557) );
  AND2_X1 U13814 ( .A1(n13468), .A2(n13467), .ZN(n14864) );
  INV_X1 U13815 ( .A(n21702), .ZN(n21778) );
  OR2_X1 U13816 ( .A1(n21343), .A2(n12682), .ZN(n21642) );
  INV_X1 U13817 ( .A(n9734), .ZN(n21332) );
  INV_X1 U13818 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21808) );
  NAND2_X1 U13819 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21804) );
  AOI21_X1 U13820 ( .B1(n15941), .B2(n15943), .A(n20233), .ZN(n15937) );
  INV_X1 U13821 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n20259) );
  NAND2_X1 U13822 ( .A1(n13632), .A2(n21133), .ZN(n13633) );
  NOR2_X1 U13823 ( .A1(n10680), .A2(n13497), .ZN(n13498) );
  AND2_X1 U13824 ( .A1(n11247), .A2(n11246), .ZN(n15972) );
  AND2_X1 U13825 ( .A1(n11672), .A2(n11671), .ZN(n16059) );
  NAND2_X1 U13826 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n12103) );
  AND2_X1 U13827 ( .A1(n17007), .A2(n12072), .ZN(n16993) );
  AND3_X1 U13828 ( .A1(n11552), .A2(n11551), .A3(n11550), .ZN(n13920) );
  INV_X1 U13829 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n22145) );
  INV_X1 U13830 ( .A(n11464), .ZN(n13769) );
  NAND2_X1 U13831 ( .A1(n14120), .A2(n11281), .ZN(n11282) );
  INV_X1 U13832 ( .A(n20614), .ZN(n20604) );
  OR3_X1 U13833 ( .A1(n20641), .A2(n20681), .A3(n20945), .ZN(n20647) );
  OR2_X1 U13834 ( .A1(n20784), .A2(n20783), .ZN(n20790) );
  INV_X1 U13835 ( .A(n20887), .ZN(n20925) );
  OR2_X1 U13836 ( .A1(n20441), .A2(n9735), .ZN(n20895) );
  OR2_X1 U13837 ( .A1(n20441), .A2(n11288), .ZN(n20915) );
  OR2_X1 U13838 ( .A1(n20441), .A2(n9722), .ZN(n20926) );
  OR2_X1 U13839 ( .A1(n11259), .A2(n10886), .ZN(n10887) );
  INV_X1 U13840 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n21021) );
  INV_X1 U13841 ( .A(n18222), .ZN(n18205) );
  NAND2_X1 U13842 ( .A1(n20190), .A2(n18818), .ZN(n12005) );
  INV_X1 U13843 ( .A(n18272), .ZN(n18291) );
  INV_X1 U13844 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n18462) );
  NOR2_X1 U13845 ( .A1(n19532), .A2(n20042), .ZN(n13980) );
  NOR2_X1 U13846 ( .A1(n18674), .A2(n18673), .ZN(n18675) );
  INV_X1 U13847 ( .A(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n18393) );
  NOR2_X1 U13848 ( .A1(n19104), .A2(n19377), .ZN(n19366) );
  INV_X1 U13849 ( .A(n19122), .ZN(n19379) );
  INV_X1 U13850 ( .A(n17326), .ZN(n18996) );
  AND4_X1 U13851 ( .A1(n11957), .A2(n11956), .A3(n11955), .A4(n11954), .ZN(
        n11963) );
  NOR2_X1 U13852 ( .A1(n19362), .A2(n19101), .ZN(n19354) );
  INV_X1 U13853 ( .A(n19430), .ZN(n19422) );
  INV_X1 U13854 ( .A(n17398), .ZN(n20015) );
  NOR2_X1 U13855 ( .A1(n20002), .A2(n20011), .ZN(n19681) );
  NOR2_X2 U13856 ( .A1(n14799), .A2(n14797), .ZN(n21212) );
  AND2_X1 U13857 ( .A1(n13541), .A2(n13539), .ZN(n21251) );
  AND2_X1 U13858 ( .A1(n21170), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n21233) );
  INV_X1 U13859 ( .A(n12672), .ZN(n21373) );
  NOR2_X1 U13860 ( .A1(n15291), .A2(n12672), .ZN(n14746) );
  OR2_X1 U13861 ( .A1(n13861), .A2(n15272), .ZN(n15292) );
  INV_X1 U13862 ( .A(n15352), .ZN(n15346) );
  OR2_X1 U13863 ( .A1(n15302), .A2(n15301), .ZN(n21321) );
  AND2_X1 U13864 ( .A1(n10642), .A2(n15158), .ZN(n21200) );
  INV_X1 U13865 ( .A(n17670), .ZN(n15576) );
  AND2_X1 U13866 ( .A1(n15714), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15740) );
  NOR3_X1 U13867 ( .A1(n15861), .A2(n15854), .A3(n15756), .ZN(n17699) );
  OR2_X1 U13868 ( .A1(n17685), .A2(n15755), .ZN(n15855) );
  INV_X1 U13869 ( .A(n15839), .ZN(n17698) );
  INV_X1 U13870 ( .A(n21339), .ZN(n21375) );
  OR2_X1 U13871 ( .A1(n15884), .A2(n9734), .ZN(n21502) );
  INV_X1 U13872 ( .A(n21446), .ZN(n21464) );
  INV_X1 U13873 ( .A(n21468), .ZN(n21494) );
  INV_X1 U13874 ( .A(n21553), .ZN(n21541) );
  INV_X1 U13875 ( .A(n21526), .ZN(n21548) );
  AND2_X1 U13876 ( .A1(n21330), .A2(n15894), .ZN(n21561) );
  INV_X1 U13877 ( .A(n21469), .ZN(n21697) );
  INV_X1 U13878 ( .A(n21665), .ZN(n21655) );
  OAI22_X1 U13879 ( .A1(n21708), .A2(n21707), .B1(n21773), .B2(n21706), .ZN(
        n21723) );
  INV_X1 U13880 ( .A(n21847), .ZN(n21752) );
  INV_X1 U13881 ( .A(n21869), .ZN(n21799) );
  INV_X1 U13882 ( .A(n21369), .ZN(n21372) );
  INV_X1 U13883 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n15923) );
  INV_X1 U13884 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n21143) );
  OR2_X1 U13885 ( .A1(n11586), .A2(n11585), .ZN(n14320) );
  INV_X1 U13886 ( .A(n14329), .ZN(n20369) );
  OR2_X1 U13887 ( .A1(n14510), .A2(n14509), .ZN(n16349) );
  OR2_X1 U13888 ( .A1(n14427), .A2(n14426), .ZN(n16362) );
  AND2_X1 U13889 ( .A1(n16240), .A2(n16256), .ZN(n20288) );
  OAI21_X1 U13890 ( .B1(n14141), .B2(n13717), .A(n13716), .ZN(n13718) );
  OAI21_X1 U13891 ( .B1(n14741), .B2(n20363), .A(n14740), .ZN(n14742) );
  AOI21_X1 U13892 ( .B1(n16914), .B2(n16913), .A(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16915) );
  AND2_X1 U13893 ( .A1(n12092), .A2(n12091), .ZN(n17741) );
  INV_X1 U13894 ( .A(n17111), .ZN(n17071) );
  NAND2_X1 U13895 ( .A1(n14049), .A2(n13806), .ZN(n20672) );
  OAI21_X1 U13896 ( .B1(n20386), .B2(n20385), .A(n20384), .ZN(n20444) );
  INV_X1 U13897 ( .A(n20452), .ZN(n20472) );
  AND2_X1 U13898 ( .A1(n20506), .A2(n20873), .ZN(n20531) );
  OAI21_X1 U13899 ( .B1(n20551), .B2(n20545), .A(n20544), .ZN(n20569) );
  OAI21_X1 U13900 ( .B1(n20583), .B2(n20582), .A(n20581), .ZN(n20607) );
  OAI21_X1 U13901 ( .B1(n20639), .B2(n20751), .A(n20612), .ZN(n20634) );
  INV_X1 U13902 ( .A(n20678), .ZN(n20681) );
  NAND2_X1 U13903 ( .A1(n20684), .A2(n20683), .ZN(n20708) );
  OAI21_X1 U13904 ( .B1(n20721), .B2(n20720), .A(n20719), .ZN(n20745) );
  INV_X1 U13905 ( .A(n20758), .ZN(n20775) );
  AND2_X1 U13906 ( .A1(n20790), .A2(n20786), .ZN(n21921) );
  OAI21_X1 U13907 ( .B1(n20830), .B2(n21106), .A(n20815), .ZN(n20832) );
  OAI21_X1 U13908 ( .B1(n20891), .B2(n20890), .A(n20889), .ZN(n20929) );
  NAND2_X1 U13909 ( .A1(n20390), .A2(n20389), .ZN(n20960) );
  INV_X1 U13910 ( .A(n20905), .ZN(n20970) );
  INV_X1 U13911 ( .A(n20920), .ZN(n20984) );
  AND3_X1 U13912 ( .A1(n11279), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n17793) );
  NOR2_X1 U13913 ( .A1(n11279), .A2(n20945), .ZN(n14142) );
  INV_X1 U13914 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n21030) );
  NOR2_X1 U13915 ( .A1(n18099), .A2(n11998), .ZN(n18009) );
  INV_X1 U13916 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n18389) );
  NOR2_X1 U13917 ( .A1(n22146), .A2(n18118), .ZN(n18098) );
  INV_X1 U13918 ( .A(n18242), .ZN(n18298) );
  INV_X1 U13919 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n18358) );
  INV_X1 U13920 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n18191) );
  INV_X1 U13921 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n18641) );
  NOR3_X1 U13922 ( .A1(n18765), .A2(n18757), .A3(n18723), .ZN(n18744) );
  NOR2_X1 U13923 ( .A1(n18908), .A2(n18791), .ZN(n18783) );
  NAND2_X1 U13924 ( .A1(n18765), .A2(n14246), .ZN(n18810) );
  INV_X1 U13925 ( .A(n19532), .ZN(n18818) );
  NAND2_X1 U13926 ( .A1(n20179), .A2(n17927), .ZN(n18857) );
  INV_X2 U13927 ( .A(n18902), .ZN(n18917) );
  INV_X1 U13928 ( .A(n19150), .ZN(n19172) );
  INV_X1 U13929 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n22088) );
  AND2_X1 U13930 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n19331) );
  INV_X1 U13931 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n19138) );
  INV_X1 U13932 ( .A(n19512), .ZN(n19473) );
  NAND2_X1 U13933 ( .A1(n19457), .A2(n20015), .ZN(n19505) );
  AND2_X1 U13934 ( .A1(n19416), .A2(n19457), .ZN(n19388) );
  NAND2_X1 U13935 ( .A1(n20044), .A2(n20138), .ZN(n20140) );
  INV_X1 U13936 ( .A(n20039), .ZN(n20151) );
  INV_X1 U13937 ( .A(n19611), .ZN(n19567) );
  NAND2_X1 U13938 ( .A1(n20021), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n19656) );
  CLKBUF_X1 U13939 ( .A(n19792), .Z(n19785) );
  INV_X1 U13940 ( .A(n19937), .ZN(n19808) );
  INV_X1 U13941 ( .A(n19963), .ZN(n19872) );
  NOR2_X1 U13942 ( .A1(n20002), .A2(n19778), .ZN(n19803) );
  INV_X1 U13943 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n20187) );
  OAI21_X1 U13944 ( .B1(P3_STATE_REG_1__SCAN_IN), .B2(n20059), .A(n20116), 
        .ZN(n20170) );
  INV_X1 U13945 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n20066) );
  INV_X1 U13946 ( .A(P1_M_IO_N_REG_SCAN_IN), .ZN(n22167) );
  INV_X1 U13947 ( .A(U212), .ZN(n17876) );
  NOR2_X1 U13948 ( .A1(n21144), .A2(n21143), .ZN(n21151) );
  INV_X1 U13949 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n22052) );
  INV_X1 U13950 ( .A(n21259), .ZN(n17647) );
  INV_X1 U13951 ( .A(n21265), .ZN(n21225) );
  OR2_X1 U13952 ( .A1(n15174), .A2(n21373), .ZN(n15195) );
  NAND2_X1 U13953 ( .A1(n21283), .A2(n12288), .ZN(n21270) );
  NAND2_X1 U13954 ( .A1(n21908), .A2(n17710), .ZN(n21281) );
  INV_X1 U13955 ( .A(n21283), .ZN(n21301) );
  INV_X1 U13956 ( .A(n21321), .ZN(n15352) );
  OR2_X1 U13957 ( .A1(n21321), .A2(n15303), .ZN(n15354) );
  NAND2_X1 U13958 ( .A1(n17676), .A2(n13841), .ZN(n17670) );
  NAND2_X1 U13959 ( .A1(n21153), .A2(n13309), .ZN(n17676) );
  INV_X1 U13960 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n21729) );
  AOI21_X1 U13961 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n21908), .A(n13924), 
        .ZN(n13947) );
  OR2_X1 U13962 ( .A1(n21436), .A2(n21469), .ZN(n21401) );
  OR2_X1 U13963 ( .A1(n21436), .A2(n21502), .ZN(n21428) );
  OR2_X1 U13964 ( .A1(n21436), .A2(n21523), .ZN(n21461) );
  OR2_X1 U13965 ( .A1(n21436), .A2(n21435), .ZN(n21468) );
  NAND2_X1 U13966 ( .A1(n21561), .A2(n21697), .ZN(n21522) );
  NAND2_X1 U13967 ( .A1(n21561), .A2(n21775), .ZN(n21583) );
  NAND2_X1 U13968 ( .A1(n21667), .A2(n21697), .ZN(n21634) );
  NAND2_X1 U13969 ( .A1(n21667), .A2(n21728), .ZN(n21665) );
  NAND2_X1 U13970 ( .A1(n21667), .A2(n21775), .ZN(n21696) );
  NAND2_X1 U13971 ( .A1(n21667), .A2(n21666), .ZN(n21727) );
  AOI22_X1 U13972 ( .A1(DATAI_20_), .A2(n21371), .B1(BUF1_REG_20__SCAN_IN), 
        .B2(n21372), .ZN(n21755) );
  NAND2_X1 U13973 ( .A1(n21776), .A2(n21728), .ZN(n21803) );
  AOI22_X1 U13974 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n21372), .B1(DATAI_24_), 
        .B2(n21371), .ZN(n21823) );
  AOI22_X1 U13975 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n21372), .B1(DATAI_29_), 
        .B2(n21371), .ZN(n21853) );
  INV_X1 U13976 ( .A(n21895), .ZN(n21875) );
  NAND2_X1 U13977 ( .A1(n13322), .A2(n21143), .ZN(n15925) );
  INV_X1 U13978 ( .A(P1_ADDRESS_REG_3__SCAN_IN), .ZN(n13613) );
  OR2_X1 U13979 ( .A1(n13813), .A2(n13625), .ZN(n13629) );
  INV_X1 U13980 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n20842) );
  NAND2_X1 U13981 ( .A1(n10668), .A2(n20227), .ZN(n11792) );
  INV_X1 U13982 ( .A(n20271), .ZN(n20231) );
  INV_X1 U13983 ( .A(n20242), .ZN(n20277) );
  INV_X1 U13984 ( .A(n16363), .ZN(n16368) );
  INV_X1 U13985 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n16342) );
  INV_X1 U13986 ( .A(n20672), .ZN(n21099) );
  INV_X1 U13987 ( .A(n20304), .ZN(n16487) );
  INV_X1 U13988 ( .A(n20303), .ZN(n16519) );
  AND2_X1 U13989 ( .A1(n13667), .A2(n13666), .ZN(n20393) );
  OR2_X1 U13990 ( .A1(n20343), .A2(n10922), .ZN(n13746) );
  NAND2_X1 U13991 ( .A1(n13718), .A2(n21129), .ZN(n20343) );
  OR2_X1 U13992 ( .A1(n17795), .A2(n13615), .ZN(n13716) );
  AOI21_X1 U13993 ( .B1(n16880), .B2(n20370), .A(n12109), .ZN(n12110) );
  OR2_X1 U13994 ( .A1(n13626), .A2(n9735), .ZN(n16737) );
  NAND2_X1 U13995 ( .A1(n14681), .A2(n17741), .ZN(n12093) );
  AOI211_X1 U13996 ( .C1(n17741), .C2(n16917), .A(n16916), .B(n16915), .ZN(
        n16918) );
  NAND2_X1 U13997 ( .A1(n12092), .A2(n17777), .ZN(n17082) );
  INV_X1 U13998 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n17751) );
  AOI21_X1 U13999 ( .B1(n17771), .B2(n17793), .A(n14144), .ZN(n17168) );
  NAND2_X2 U14000 ( .A1(n20457), .A2(n20673), .ZN(n20477) );
  NAND2_X1 U14001 ( .A1(n20506), .A2(n20779), .ZN(n20547) );
  NAND2_X1 U14002 ( .A1(n21090), .A2(n20541), .ZN(n20605) );
  NAND2_X1 U14003 ( .A1(n21090), .A2(n20575), .ZN(n20620) );
  AND2_X1 U14004 ( .A1(n20644), .A2(n20643), .ZN(n20655) );
  OR2_X1 U14005 ( .A1(n21091), .A2(n20673), .ZN(n20706) );
  NAND2_X1 U14006 ( .A1(n20713), .A2(n20673), .ZN(n20743) );
  NAND2_X1 U14007 ( .A1(n20780), .A2(n20873), .ZN(n21927) );
  NAND2_X1 U14008 ( .A1(n20780), .A2(n20779), .ZN(n20835) );
  INV_X1 U14009 ( .A(n20980), .ZN(n20916) );
  INV_X1 U14010 ( .A(n20960), .ZN(n20899) );
  AND2_X1 U14011 ( .A1(n20944), .A2(n20943), .ZN(n20959) );
  INV_X1 U14012 ( .A(n20857), .ZN(n21928) );
  INV_X1 U14013 ( .A(n21085), .ZN(n21009) );
  INV_X1 U14014 ( .A(HOLD), .ZN(n21020) );
  INV_X1 U14015 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n17926) );
  INV_X1 U14016 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n18002) );
  INV_X1 U14017 ( .A(n9707), .ZN(n18290) );
  INV_X1 U14018 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n18301) );
  INV_X1 U14019 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n18644) );
  INV_X1 U14020 ( .A(BUF2_REG_27__SCAN_IN), .ZN(n22056) );
  NAND2_X1 U14021 ( .A1(n19551), .A2(n18784), .ZN(n18760) );
  NOR2_X1 U14022 ( .A1(n22098), .A2(n18774), .ZN(n18777) );
  NOR2_X1 U14023 ( .A1(n17208), .A2(n17207), .ZN(n18806) );
  INV_X1 U14024 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n18817) );
  NAND2_X1 U14025 ( .A1(n18843), .A2(n18818), .ZN(n18834) );
  NAND2_X1 U14026 ( .A1(n18854), .A2(n18855), .ZN(n18853) );
  INV_X1 U14027 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n18873) );
  INV_X1 U14028 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n18875) );
  INV_X1 U14029 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n18887) );
  AOI211_X1 U14030 ( .C1(n20171), .C2(n20172), .A(n18858), .B(n18857), .ZN(
        n18902) );
  INV_X1 U14031 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n18988) );
  INV_X1 U14032 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n19319) );
  INV_X1 U14033 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n19377) );
  NAND2_X1 U14034 ( .A1(n19517), .A2(n14191), .ZN(n19512) );
  INV_X1 U14035 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20011) );
  INV_X1 U14036 ( .A(n20155), .ZN(n20158) );
  INV_X1 U14037 ( .A(n19910), .ZN(n19880) );
  INV_X1 U14038 ( .A(n19618), .ZN(n19631) );
  INV_X1 U14039 ( .A(n19645), .ZN(n19654) );
  INV_X1 U14040 ( .A(n19671), .ZN(n19680) );
  INV_X1 U14041 ( .A(n19692), .ZN(n19705) );
  INV_X1 U14042 ( .A(n19720), .ZN(n19727) );
  INV_X1 U14043 ( .A(n19740), .ZN(n19750) );
  INV_X1 U14044 ( .A(n19820), .ZN(n19828) );
  NAND2_X1 U14045 ( .A1(n19921), .A2(BUF2_REG_22__SCAN_IN), .ZN(n19875) );
  NAND2_X1 U14046 ( .A1(n19921), .A2(BUF2_REG_19__SCAN_IN), .ZN(n19898) );
  NAND2_X1 U14047 ( .A1(n19921), .A2(BUF2_REG_18__SCAN_IN), .ZN(n19937) );
  NAND2_X1 U14048 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n19921), .ZN(n19949) );
  INV_X1 U14049 ( .A(n18280), .ZN(n20051) );
  INV_X1 U14050 ( .A(n20136), .ZN(n20054) );
  INV_X1 U14051 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n20073) );
  INV_X1 U14052 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n22085) );
  INV_X1 U14053 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n20113) );
  NAND2_X1 U14054 ( .A1(n20184), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n20130) );
  NOR2_X1 U14055 ( .A1(n14329), .A2(n13575), .ZN(n17836) );
  INV_X1 U14056 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n22011) );
  INV_X1 U14057 ( .A(n17880), .ZN(n17878) );
  OAI211_X1 U14058 ( .C1(n16891), .C2(n16737), .A(n10682), .B(n12110), .ZN(
        P2_U2995) );
  AND2_X1 U14059 ( .A1(n10710), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10686) );
  AOI22_X1 U14060 ( .A1(n10732), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10733), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10692) );
  NAND2_X1 U14061 ( .A1(n10780), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n10691) );
  AND2_X2 U14062 ( .A1(n9730), .A2(n14126), .ZN(n10758) );
  NAND2_X1 U14063 ( .A1(n10758), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n10690) );
  INV_X1 U14064 ( .A(n10693), .ZN(n10687) );
  NOR2_X1 U14065 ( .A1(n10687), .A2(n14126), .ZN(n10878) );
  INV_X1 U14066 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10688) );
  OR2_X1 U14067 ( .A1(n9712), .A2(n10688), .ZN(n10689) );
  NAND4_X1 U14068 ( .A1(n10692), .A2(n10691), .A3(n10690), .A4(n10689), .ZN(
        n10699) );
  BUF_X1 U14069 ( .A(n10865), .Z(n14666) );
  NAND2_X1 U14070 ( .A1(n11066), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n10697) );
  BUF_X4 U14071 ( .A(n10813), .Z(n14565) );
  AND2_X2 U14072 ( .A1(n14565), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10759) );
  NAND2_X1 U14073 ( .A1(n10759), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n10696) );
  AND2_X2 U14074 ( .A1(n9733), .A2(n14126), .ZN(n14416) );
  NAND2_X1 U14075 ( .A1(n14416), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n10695) );
  NAND2_X1 U14076 ( .A1(n10764), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n10694) );
  NAND4_X1 U14077 ( .A1(n10697), .A2(n10696), .A3(n10695), .A4(n10694), .ZN(
        n10698) );
  AND2_X4 U14078 ( .A1(n10700), .A2(n10750), .ZN(n14458) );
  AND2_X2 U14079 ( .A1(n14458), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10769) );
  NAND2_X1 U14080 ( .A1(n10866), .A2(n14126), .ZN(n14125) );
  INV_X2 U14081 ( .A(n14125), .ZN(n14444) );
  AOI22_X1 U14082 ( .A1(n10769), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n14444), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10707) );
  AND3_X4 U14083 ( .A1(n10750), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(
        n10701), .ZN(n14457) );
  AND2_X2 U14084 ( .A1(n14457), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14486) );
  AOI22_X1 U14085 ( .A1(n14486), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10877), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10706) );
  AND2_X1 U14086 ( .A1(n10702), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10703) );
  AOI22_X1 U14087 ( .A1(n14504), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10781), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10705) );
  NAND2_X1 U14088 ( .A1(n14503), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n10704) );
  NAND4_X1 U14089 ( .A1(n10707), .A2(n10706), .A3(n10705), .A4(n10704), .ZN(
        n10708) );
  NAND2_X1 U14090 ( .A1(n21114), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10880) );
  NAND2_X1 U14091 ( .A1(n10710), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n10711) );
  NAND2_X1 U14092 ( .A1(n10880), .A2(n10711), .ZN(n11259) );
  INV_X1 U14093 ( .A(n11259), .ZN(n11264) );
  AOI22_X1 U14094 ( .A1(n14565), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n9729), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10713) );
  AOI22_X1 U14095 ( .A1(n14457), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10868), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10715) );
  AOI22_X1 U14096 ( .A1(n14458), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9720), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10714) );
  AOI22_X1 U14097 ( .A1(n14565), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n9729), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10717) );
  AOI22_X1 U14098 ( .A1(n10828), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10865), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10716) );
  AOI21_X1 U14099 ( .B1(n14664), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A(
        n14126), .ZN(n10719) );
  AOI22_X1 U14100 ( .A1(n14457), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10868), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10722) );
  AOI22_X1 U14101 ( .A1(n14565), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n9729), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10721) );
  AOI22_X1 U14102 ( .A1(n10828), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10865), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10720) );
  AOI22_X1 U14103 ( .A1(n14457), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10868), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10726) );
  AOI22_X1 U14104 ( .A1(n10828), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10865), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10728) );
  AOI22_X1 U14105 ( .A1(n14565), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n10866), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10727) );
  MUX2_X1 U14106 ( .A(n13769), .B(n11264), .S(n10926), .Z(n11323) );
  NAND2_X1 U14107 ( .A1(n20837), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10748) );
  NAND2_X1 U14108 ( .A1(n10702), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n10730) );
  NAND2_X1 U14109 ( .A1(n10748), .A2(n10730), .ZN(n11258) );
  INV_X1 U14110 ( .A(n11258), .ZN(n10731) );
  NAND2_X1 U14111 ( .A1(n11323), .A2(n10731), .ZN(n10757) );
  AOI22_X1 U14112 ( .A1(n11066), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10780), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10741) );
  AOI22_X1 U14113 ( .A1(n10758), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10759), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10740) );
  INV_X1 U14114 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10736) );
  NAND2_X1 U14115 ( .A1(n10732), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n10735) );
  NAND2_X1 U14116 ( .A1(n10733), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n10734) );
  OAI211_X1 U14117 ( .C1(n14497), .C2(n10736), .A(n10735), .B(n10734), .ZN(
        n10737) );
  INV_X1 U14118 ( .A(n10737), .ZN(n10739) );
  AOI22_X1 U14119 ( .A1(n10764), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n14444), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10738) );
  NAND4_X1 U14120 ( .A1(n10741), .A2(n10740), .A3(n10739), .A4(n10738), .ZN(
        n10747) );
  AOI22_X1 U14121 ( .A1(n10769), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n14416), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10745) );
  AOI22_X1 U14122 ( .A1(n14504), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n10781), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10743) );
  NAND2_X1 U14123 ( .A1(n14486), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n10742) );
  NAND4_X1 U14124 ( .A1(n10745), .A2(n10744), .A3(n10743), .A4(n10742), .ZN(
        n10746) );
  NAND2_X1 U14125 ( .A1(n22183), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10776) );
  NAND2_X1 U14126 ( .A1(n10750), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10751) );
  NAND2_X1 U14127 ( .A1(n10776), .A2(n10751), .ZN(n10753) );
  NAND2_X1 U14128 ( .A1(n10752), .A2(n10753), .ZN(n10756) );
  INV_X1 U14129 ( .A(n10752), .ZN(n10755) );
  INV_X1 U14130 ( .A(n10753), .ZN(n10754) );
  NAND2_X1 U14131 ( .A1(n10755), .A2(n10754), .ZN(n10777) );
  NAND2_X1 U14132 ( .A1(n10756), .A2(n10777), .ZN(n11261) );
  INV_X1 U14133 ( .A(n11261), .ZN(n11268) );
  NAND2_X1 U14134 ( .A1(n10926), .A2(n11268), .ZN(n11267) );
  NAND2_X1 U14135 ( .A1(n10757), .A2(n11291), .ZN(n10804) );
  AOI22_X1 U14136 ( .A1(n10758), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11066), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10768) );
  AOI22_X1 U14137 ( .A1(n10759), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10780), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10767) );
  INV_X1 U14138 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10762) );
  NAND2_X1 U14139 ( .A1(n10732), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n10761) );
  NAND2_X1 U14140 ( .A1(n10733), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n10760) );
  OAI211_X1 U14141 ( .C1(n14497), .C2(n10762), .A(n10761), .B(n10760), .ZN(
        n10763) );
  INV_X1 U14142 ( .A(n10763), .ZN(n10766) );
  AOI22_X1 U14143 ( .A1(n10764), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n14444), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10765) );
  NAND4_X1 U14144 ( .A1(n10768), .A2(n10767), .A3(n10766), .A4(n10765), .ZN(
        n10775) );
  AOI22_X1 U14145 ( .A1(n10769), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n14416), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10773) );
  AOI22_X1 U14146 ( .A1(n10877), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n14503), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10772) );
  AOI22_X1 U14147 ( .A1(n14504), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n10781), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10771) );
  NAND2_X1 U14148 ( .A1(n14486), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n10770) );
  NAND4_X1 U14149 ( .A1(n10773), .A2(n10772), .A3(n10771), .A4(n10770), .ZN(
        n10774) );
  NAND2_X1 U14150 ( .A1(n10777), .A2(n10776), .ZN(n10798) );
  NAND2_X1 U14151 ( .A1(n10798), .A2(n10796), .ZN(n10779) );
  NAND2_X1 U14152 ( .A1(n21096), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10778) );
  NAND2_X1 U14153 ( .A1(n10779), .A2(n10778), .ZN(n10800) );
  NAND2_X1 U14154 ( .A1(n17770), .A2(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(
        n10801) );
  MUX2_X1 U14155 ( .A(n11501), .B(n10883), .S(n10926), .Z(n11295) );
  AOI22_X1 U14156 ( .A1(n14493), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n14477), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10795) );
  AOI22_X1 U14157 ( .A1(n10769), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n14444), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10785) );
  AOI22_X1 U14158 ( .A1(n10877), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n14503), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10784) );
  AOI22_X1 U14159 ( .A1(n10781), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10733), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10783) );
  NAND2_X1 U14160 ( .A1(n14486), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n10782) );
  NAND4_X1 U14161 ( .A1(n10785), .A2(n10784), .A3(n10783), .A4(n10782), .ZN(
        n10793) );
  INV_X1 U14162 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11027) );
  NAND2_X1 U14163 ( .A1(n14504), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n10787) );
  NAND2_X1 U14164 ( .A1(n10732), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n10786) );
  OAI211_X1 U14165 ( .C1(n14497), .C2(n11027), .A(n10787), .B(n10786), .ZN(
        n10788) );
  INV_X1 U14166 ( .A(n10788), .ZN(n10791) );
  AOI22_X1 U14167 ( .A1(n14416), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n10764), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10790) );
  AOI22_X1 U14168 ( .A1(n10758), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10759), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10789) );
  NAND3_X1 U14169 ( .A1(n10791), .A2(n10790), .A3(n10789), .ZN(n10792) );
  NAND2_X1 U14170 ( .A1(n10795), .A2(n10794), .ZN(n11495) );
  INV_X1 U14171 ( .A(n10796), .ZN(n10797) );
  XNOR2_X1 U14172 ( .A(n10798), .B(n10797), .ZN(n10882) );
  MUX2_X1 U14173 ( .A(n11495), .B(n10882), .S(n10926), .Z(n11294) );
  AND2_X1 U14174 ( .A1(n11295), .A2(n11294), .ZN(n10803) );
  NOR2_X1 U14175 ( .A1(n17770), .A2(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(
        n10799) );
  AOI21_X1 U14176 ( .B1(n10804), .B2(n10803), .A(n11276), .ZN(n17781) );
  AOI22_X1 U14177 ( .A1(n9730), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n10865), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10808) );
  AOI22_X1 U14178 ( .A1(n14457), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10868), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10807) );
  AOI22_X1 U14179 ( .A1(n14565), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10866), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10806) );
  AOI22_X1 U14180 ( .A1(n14458), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n14664), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10805) );
  AOI22_X1 U14181 ( .A1(n9730), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10865), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10812) );
  AOI22_X1 U14182 ( .A1(n14457), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10868), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10811) );
  AOI22_X1 U14183 ( .A1(n14565), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n9714), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10810) );
  AOI22_X1 U14184 ( .A1(n9733), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9729), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10809) );
  AOI22_X1 U14185 ( .A1(n10867), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n10866), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10817) );
  AOI22_X1 U14186 ( .A1(n14457), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n10868), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10816) );
  AOI22_X1 U14187 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n10865), .B1(
        n10828), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10815) );
  AOI22_X1 U14188 ( .A1(n9714), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(n9733), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10814) );
  NAND4_X1 U14189 ( .A1(n10817), .A2(n10816), .A3(n10815), .A4(n10814), .ZN(
        n10914) );
  NAND2_X1 U14190 ( .A1(n10914), .A2(n14126), .ZN(n10823) );
  AOI22_X1 U14191 ( .A1(n10867), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n9729), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10821) );
  AOI22_X1 U14192 ( .A1(n14457), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10868), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10820) );
  AOI22_X1 U14193 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n10828), .B1(
        n10865), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10819) );
  NAND4_X1 U14194 ( .A1(n10821), .A2(n10820), .A3(n10819), .A4(n10818), .ZN(
        n10911) );
  NAND2_X1 U14195 ( .A1(n10911), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10822) );
  NAND2_X4 U14196 ( .A1(n10823), .A2(n10822), .ZN(n13819) );
  AOI22_X1 U14197 ( .A1(n14457), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10868), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10825) );
  AOI22_X1 U14198 ( .A1(n14458), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9732), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10824) );
  AOI22_X1 U14199 ( .A1(n14646), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10865), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10827) );
  AOI22_X1 U14200 ( .A1(n10867), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10866), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10826) );
  AOI22_X1 U14201 ( .A1(n9730), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n10865), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10832) );
  AOI22_X1 U14202 ( .A1(n14457), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n10868), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10831) );
  AOI22_X1 U14203 ( .A1(n10867), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n9729), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10830) );
  AOI22_X1 U14204 ( .A1(n9714), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n14664), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10829) );
  AOI22_X1 U14205 ( .A1(n14458), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n14664), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10834) );
  AOI22_X1 U14206 ( .A1(n14457), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10868), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10833) );
  AND2_X1 U14207 ( .A1(n10834), .A2(n10833), .ZN(n10837) );
  AOI22_X1 U14208 ( .A1(n9730), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n10865), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10836) );
  AOI22_X1 U14209 ( .A1(n14565), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n10866), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10835) );
  NAND3_X1 U14210 ( .A1(n10837), .A2(n10836), .A3(n10835), .ZN(n10913) );
  AOI22_X1 U14211 ( .A1(n9730), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10865), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10841) );
  AOI22_X1 U14212 ( .A1(n14457), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10868), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10840) );
  AOI22_X1 U14213 ( .A1(n10867), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10866), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10839) );
  AOI22_X1 U14214 ( .A1(n9714), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n14664), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10838) );
  AOI22_X1 U14215 ( .A1(n9730), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10865), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10848) );
  AOI22_X1 U14216 ( .A1(n14565), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n9729), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10847) );
  AOI22_X1 U14217 ( .A1(n14457), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10868), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10846) );
  NAND4_X1 U14218 ( .A1(n10849), .A2(n10848), .A3(n10847), .A4(n10846), .ZN(
        n10857) );
  AOI22_X1 U14219 ( .A1(n9730), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n10865), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10854) );
  AOI22_X1 U14220 ( .A1(n10867), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n10866), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10853) );
  AOI22_X1 U14221 ( .A1(n14457), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10868), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10852) );
  NAND4_X1 U14222 ( .A1(n10855), .A2(n10854), .A3(n10853), .A4(n10852), .ZN(
        n10856) );
  AOI22_X1 U14223 ( .A1(n14457), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10868), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10859) );
  AOI22_X1 U14224 ( .A1(n14565), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10866), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10862) );
  AOI22_X1 U14225 ( .A1(n9730), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10865), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10861) );
  NAND3_X1 U14226 ( .A1(n9815), .A2(n10862), .A3(n10861), .ZN(n10874) );
  NAND2_X1 U14227 ( .A1(n14458), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n10863) );
  AOI22_X1 U14228 ( .A1(n9730), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10865), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10871) );
  AOI22_X1 U14229 ( .A1(n10867), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10866), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10870) );
  AOI22_X1 U14230 ( .A1(n14457), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10868), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10869) );
  NAND4_X1 U14231 ( .A1(n10872), .A2(n10871), .A3(n10870), .A4(n10869), .ZN(
        n10873) );
  INV_X1 U14232 ( .A(n12029), .ZN(n10876) );
  NAND2_X1 U14233 ( .A1(n17781), .A2(n17777), .ZN(n17768) );
  INV_X1 U14234 ( .A(n10877), .ZN(n10879) );
  NOR2_X1 U14235 ( .A1(n10878), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n17163) );
  AOI21_X1 U14236 ( .B1(n10879), .B2(n17163), .A(P2_FLUSH_REG_SCAN_IN), .ZN(
        n21108) );
  INV_X1 U14237 ( .A(n10880), .ZN(n10881) );
  XNOR2_X1 U14238 ( .A(n11258), .B(n10881), .ZN(n11263) );
  INV_X1 U14239 ( .A(n10885), .ZN(n10886) );
  NAND2_X1 U14240 ( .A1(n17778), .A2(n10887), .ZN(n10888) );
  MUX2_X1 U14241 ( .A(n21108), .B(n10888), .S(n11279), .Z(n21119) );
  INV_X1 U14242 ( .A(n21119), .ZN(n12039) );
  NAND2_X1 U14243 ( .A1(n12039), .A2(n21118), .ZN(n10889) );
  NAND2_X1 U14244 ( .A1(n17768), .A2(n10889), .ZN(n10890) );
  NAND2_X1 U14245 ( .A1(n10875), .A2(n10900), .ZN(n10899) );
  NAND2_X1 U14246 ( .A1(n10899), .A2(n10891), .ZN(n12025) );
  NAND2_X1 U14247 ( .A1(n12030), .A2(n20415), .ZN(n12028) );
  NAND2_X1 U14248 ( .A1(n10893), .A2(n12028), .ZN(n12054) );
  NAND2_X1 U14249 ( .A1(n12054), .A2(n12056), .ZN(n10897) );
  NAND2_X1 U14250 ( .A1(n12061), .A2(n10895), .ZN(n10896) );
  NAND2_X1 U14251 ( .A1(n11476), .A2(n10898), .ZN(n12062) );
  NAND2_X1 U14252 ( .A1(n10899), .A2(n12056), .ZN(n10933) );
  INV_X1 U14253 ( .A(n10892), .ZN(n10903) );
  AND2_X1 U14254 ( .A1(n20400), .A2(n9736), .ZN(n10904) );
  INV_X1 U14255 ( .A(n10910), .ZN(n10912) );
  NAND3_X1 U14256 ( .A1(n10912), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n10911), .ZN(n10917) );
  INV_X1 U14257 ( .A(n10913), .ZN(n10915) );
  NAND3_X1 U14258 ( .A1(n10915), .A2(n14126), .A3(n10914), .ZN(n10916) );
  AOI21_X1 U14259 ( .B1(n10917), .B2(n10916), .A(n12040), .ZN(n10918) );
  NOR2_X1 U14260 ( .A1(n10014), .A2(n9722), .ZN(n10921) );
  INV_X1 U14261 ( .A(n17796), .ZN(n10937) );
  NAND2_X1 U14262 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n10924) );
  NAND2_X1 U14263 ( .A1(n10937), .A2(n10924), .ZN(n10925) );
  AOI21_X1 U14264 ( .B1(n11161), .B2(P2_REIP_REG_0__SCAN_IN), .A(n10925), .ZN(
        n10929) );
  AND2_X2 U14265 ( .A1(n10936), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11160) );
  NAND2_X1 U14266 ( .A1(n11160), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n10928) );
  INV_X1 U14267 ( .A(n10931), .ZN(n10932) );
  NAND3_X1 U14268 ( .A1(n10935), .A2(n10934), .A3(n10933), .ZN(n17127) );
  INV_X1 U14269 ( .A(n12063), .ZN(n12027) );
  NOR2_X1 U14270 ( .A1(n10937), .A2(n21114), .ZN(n10938) );
  AOI21_X1 U14271 ( .B1(n17152), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n10938), 
        .ZN(n10940) );
  NAND2_X1 U14272 ( .A1(n10960), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10939) );
  NAND2_X1 U14273 ( .A1(n10960), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10943) );
  AOI22_X1 U14274 ( .A1(n14127), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n17796), .ZN(n10942) );
  NAND2_X1 U14275 ( .A1(n10943), .A2(n10942), .ZN(n10950) );
  INV_X1 U14276 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n11040) );
  NAND2_X1 U14277 ( .A1(n11160), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(n10945) );
  AOI22_X1 U14278 ( .A1(n11161), .A2(P2_REIP_REG_1__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n10944) );
  NAND2_X1 U14279 ( .A1(n10960), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10947) );
  AOI21_X1 U14280 ( .B1(n21132), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n10946) );
  NAND2_X1 U14281 ( .A1(n10947), .A2(n10946), .ZN(n10954) );
  INV_X1 U14282 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n12077) );
  AOI22_X1 U14283 ( .A1(n11161), .A2(P2_REIP_REG_2__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10949) );
  NAND2_X1 U14284 ( .A1(n11160), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n10948) );
  OAI211_X1 U14285 ( .C1(n10957), .C2(n12077), .A(n10949), .B(n10948), .ZN(
        n10953) );
  NAND2_X1 U14286 ( .A1(n10954), .A2(n10953), .ZN(n10967) );
  INV_X1 U14287 ( .A(n10966), .ZN(n10952) );
  NAND2_X1 U14288 ( .A1(n10952), .A2(n10967), .ZN(n10955) );
  OR2_X1 U14289 ( .A1(n10954), .A2(n10953), .ZN(n10968) );
  AOI22_X1 U14290 ( .A1(n11161), .A2(P2_REIP_REG_3__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10959) );
  NAND2_X1 U14291 ( .A1(n11160), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n10958) );
  AOI22_X1 U14292 ( .A1(n10960), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n17796), .B2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n10961) );
  XNOR2_X1 U14293 ( .A(n11159), .B(n10961), .ZN(n10962) );
  XNOR2_X2 U14294 ( .A(n11157), .B(n10962), .ZN(n10986) );
  NAND2_X1 U14295 ( .A1(n10970), .A2(n10966), .ZN(n10969) );
  BUF_X2 U14296 ( .A(n10974), .Z(n14041) );
  INV_X1 U14297 ( .A(n14041), .ZN(n14714) );
  AND2_X2 U14298 ( .A1(n10975), .A2(n14714), .ZN(n11000) );
  NAND2_X1 U14299 ( .A1(n10980), .A2(n10971), .ZN(n10972) );
  NAND2_X2 U14300 ( .A1(n10973), .A2(n10972), .ZN(n13801) );
  NAND2_X2 U14301 ( .A1(n11000), .A2(n13801), .ZN(n20754) );
  INV_X1 U14302 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n14521) );
  NAND2_X1 U14303 ( .A1(n20888), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n10977) );
  BUF_X4 U14304 ( .A(n10974), .Z(n17146) );
  NAND2_X1 U14305 ( .A1(n11052), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n10976) );
  OAI211_X1 U14306 ( .C1(n20754), .C2(n14521), .A(n10977), .B(n10976), .ZN(
        n10978) );
  INV_X1 U14307 ( .A(n10978), .ZN(n10998) );
  NAND2_X1 U14308 ( .A1(n13778), .A2(n10979), .ZN(n10990) );
  NAND2_X1 U14309 ( .A1(n10980), .A2(n13778), .ZN(n10985) );
  NOR2_X2 U14310 ( .A1(n11001), .A2(n17744), .ZN(n20718) );
  AOI22_X1 U14311 ( .A1(n20784), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n20718), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10997) );
  NOR2_X2 U14312 ( .A1(n10981), .A2(n17733), .ZN(n20509) );
  INV_X1 U14313 ( .A(n10985), .ZN(n10982) );
  NAND3_X1 U14314 ( .A1(n17146), .A2(n10982), .A3(n10991), .ZN(n11087) );
  INV_X1 U14315 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10983) );
  OAI21_X1 U14316 ( .B1(n11087), .B2(n10983), .A(n9736), .ZN(n10984) );
  AOI21_X1 U14317 ( .B1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n20509), .A(
        n10984), .ZN(n10996) );
  INV_X1 U14318 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10989) );
  NOR2_X1 U14319 ( .A1(n10986), .A2(n10985), .ZN(n10987) );
  INV_X1 U14320 ( .A(n20580), .ZN(n11086) );
  INV_X1 U14321 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10988) );
  OAI22_X1 U14322 ( .A1(n11050), .A2(n10989), .B1(n11086), .B2(n10988), .ZN(
        n10994) );
  INV_X1 U14323 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10992) );
  NOR2_X1 U14324 ( .A1(n10994), .A2(n10993), .ZN(n10995) );
  NAND4_X1 U14325 ( .A1(n10998), .A2(n10997), .A3(n10996), .A4(n10995), .ZN(
        n11009) );
  NAND2_X1 U14326 ( .A1(n10999), .A2(n13801), .ZN(n20481) );
  INV_X1 U14327 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n14514) );
  OR2_X1 U14328 ( .A1(n20481), .A2(n14514), .ZN(n11007) );
  NAND2_X1 U14329 ( .A1(n10999), .A2(n17104), .ZN(n20382) );
  INV_X1 U14330 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11012) );
  OR2_X1 U14331 ( .A1(n20382), .A2(n11012), .ZN(n11006) );
  NAND2_X2 U14332 ( .A1(n11000), .A2(n17104), .ZN(n11097) );
  INV_X1 U14333 ( .A(n11097), .ZN(n20676) );
  NAND2_X1 U14334 ( .A1(n20676), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11005) );
  NAND4_X1 U14335 ( .A1(n11007), .A2(n11006), .A3(n11005), .A4(n11004), .ZN(
        n11008) );
  AOI22_X1 U14336 ( .A1(n10758), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11066), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11016) );
  AOI22_X1 U14337 ( .A1(n10759), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10780), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11015) );
  NAND2_X1 U14338 ( .A1(n14504), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11011) );
  NAND2_X1 U14339 ( .A1(n10732), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n11010) );
  OAI211_X1 U14340 ( .C1(n14497), .C2(n11012), .A(n11011), .B(n11010), .ZN(
        n11013) );
  AOI22_X1 U14341 ( .A1(n14416), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n10764), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11014) );
  AOI22_X1 U14342 ( .A1(n10769), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n14444), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11020) );
  AOI22_X1 U14343 ( .A1(n14486), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n14503), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11019) );
  AOI22_X1 U14344 ( .A1(n10781), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n10733), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11018) );
  NAND2_X1 U14345 ( .A1(n10877), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n11017) );
  NAND4_X1 U14346 ( .A1(n11020), .A2(n11019), .A3(n11018), .A4(n11017), .ZN(
        n11021) );
  NAND3_X1 U14347 ( .A1(n13769), .A2(n9735), .A3(n11479), .ZN(n11037) );
  INV_X1 U14348 ( .A(n11486), .ZN(n11022) );
  AOI22_X1 U14349 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n11052), .B1(
        n20888), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11025) );
  AOI22_X1 U14350 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20580), .B1(
        n20641), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11024) );
  AOI22_X1 U14351 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20839), .B1(
        n20940), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11023) );
  INV_X1 U14352 ( .A(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n14559) );
  OAI22_X1 U14353 ( .A1(n14559), .A2(n20481), .B1(n20382), .B2(n11027), .ZN(
        n11030) );
  INV_X1 U14354 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11028) );
  INV_X1 U14355 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n14567) );
  OAI22_X1 U14356 ( .A1(n11028), .A2(n11097), .B1(n20754), .B2(n14567), .ZN(
        n11029) );
  NOR2_X1 U14357 ( .A1(n11030), .A2(n11029), .ZN(n11033) );
  AOI22_X1 U14358 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20784), .B1(
        n20449), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11032) );
  AOI22_X1 U14359 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20509), .B1(
        n20718), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11031) );
  INV_X1 U14360 ( .A(n11495), .ZN(n11035) );
  NAND2_X1 U14361 ( .A1(n11035), .A2(n9735), .ZN(n11036) );
  XNOR2_X1 U14362 ( .A(n11486), .B(n11037), .ZN(n11043) );
  XNOR2_X1 U14363 ( .A(n11043), .B(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n14686) );
  INV_X1 U14364 ( .A(n11479), .ZN(n11038) );
  NOR3_X1 U14365 ( .A1(n11038), .A2(n17130), .A3(n13769), .ZN(n11042) );
  NAND2_X1 U14366 ( .A1(n11464), .A2(n17130), .ZN(n11039) );
  XNOR2_X1 U14367 ( .A(n11039), .B(n11479), .ZN(n13761) );
  NOR2_X1 U14368 ( .A1(n11040), .A2(n13761), .ZN(n11041) );
  OR2_X1 U14369 ( .A1(n11042), .A2(n11041), .ZN(n14685) );
  NAND2_X1 U14370 ( .A1(n14686), .A2(n14685), .ZN(n14688) );
  INV_X1 U14371 ( .A(n11043), .ZN(n11044) );
  NAND2_X1 U14372 ( .A1(n11044), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11045) );
  NAND2_X1 U14373 ( .A1(n14688), .A2(n11045), .ZN(n11047) );
  XNOR2_X1 U14374 ( .A(n11047), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n17732) );
  INV_X1 U14375 ( .A(n17732), .ZN(n11046) );
  NAND2_X1 U14376 ( .A1(n11047), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11048) );
  INV_X1 U14377 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n17097) );
  INV_X1 U14378 ( .A(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11051) );
  INV_X1 U14379 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11053) );
  NOR2_X1 U14380 ( .A1(n11055), .A2(n11054), .ZN(n11065) );
  INV_X1 U14381 ( .A(n20641), .ZN(n11092) );
  INV_X1 U14382 ( .A(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11057) );
  INV_X1 U14383 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11056) );
  OAI22_X1 U14384 ( .A1(n11092), .A2(n11057), .B1(n11091), .B2(n11056), .ZN(
        n11061) );
  INV_X1 U14385 ( .A(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11059) );
  INV_X1 U14386 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11058) );
  OAI22_X1 U14387 ( .A1(n11086), .A2(n11059), .B1(n11087), .B2(n11058), .ZN(
        n11060) );
  INV_X1 U14388 ( .A(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n14609) );
  INV_X1 U14389 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11062) );
  OAI22_X1 U14390 ( .A1(n14609), .A2(n20481), .B1(n11097), .B2(n11062), .ZN(
        n11063) );
  INV_X1 U14391 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n14616) );
  INV_X1 U14392 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n14283) );
  OAI22_X1 U14393 ( .A1(n14616), .A2(n20754), .B1(n20382), .B2(n14283), .ZN(
        n11064) );
  AOI22_X1 U14394 ( .A1(n10758), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n14493), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11073) );
  AOI22_X1 U14395 ( .A1(n10759), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n14477), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11072) );
  NAND2_X1 U14396 ( .A1(n10732), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n11068) );
  NAND2_X1 U14397 ( .A1(n10733), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n11067) );
  OAI211_X1 U14398 ( .C1(n14497), .C2(n14283), .A(n11068), .B(n11067), .ZN(
        n11069) );
  INV_X1 U14399 ( .A(n11069), .ZN(n11071) );
  AOI22_X1 U14400 ( .A1(n10764), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n14444), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11070) );
  NAND4_X1 U14401 ( .A1(n11073), .A2(n11072), .A3(n11071), .A4(n11070), .ZN(
        n11079) );
  AOI22_X1 U14402 ( .A1(n10769), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n14416), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11077) );
  AOI22_X1 U14403 ( .A1(n10877), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n14503), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11076) );
  AOI22_X1 U14404 ( .A1(n14504), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10781), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11075) );
  NAND2_X1 U14405 ( .A1(n14486), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n11074) );
  NAND4_X1 U14406 ( .A1(n11077), .A2(n11076), .A3(n11075), .A4(n11074), .ZN(
        n11078) );
  NAND2_X1 U14407 ( .A1(n11297), .A2(n9735), .ZN(n11080) );
  INV_X1 U14408 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n17073) );
  INV_X1 U14409 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11082) );
  INV_X1 U14410 ( .A(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11081) );
  OAI22_X1 U14411 ( .A1(n11082), .A2(n11050), .B1(n20546), .B2(n11081), .ZN(
        n11085) );
  INV_X1 U14412 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11083) );
  NOR2_X1 U14413 ( .A1(n11085), .A2(n11084), .ZN(n11104) );
  INV_X1 U14414 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11089) );
  INV_X1 U14415 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11088) );
  OAI22_X1 U14416 ( .A1(n11086), .A2(n11089), .B1(n11087), .B2(n11088), .ZN(
        n11094) );
  INV_X1 U14417 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n14625) );
  INV_X1 U14418 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11090) );
  OAI22_X1 U14419 ( .A1(n11092), .A2(n14625), .B1(n11091), .B2(n11090), .ZN(
        n11093) );
  NOR2_X1 U14420 ( .A1(n11094), .A2(n11093), .ZN(n11103) );
  AOI22_X1 U14421 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20509), .B1(
        n20718), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11102) );
  INV_X1 U14422 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11107) );
  INV_X1 U14423 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n14635) );
  OAI22_X1 U14424 ( .A1(n11107), .A2(n20382), .B1(n20754), .B2(n14635), .ZN(
        n11095) );
  INV_X1 U14425 ( .A(n11095), .ZN(n11101) );
  INV_X1 U14426 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n14496) );
  INV_X1 U14427 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11096) );
  OAI22_X1 U14428 ( .A1(n14496), .A2(n20481), .B1(n11097), .B2(n11096), .ZN(
        n11098) );
  INV_X1 U14429 ( .A(n11098), .ZN(n11100) );
  AOI22_X1 U14430 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20784), .B1(
        n20449), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11099) );
  AOI22_X1 U14431 ( .A1(n10758), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n14493), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11112) );
  AOI22_X1 U14432 ( .A1(n10759), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n14477), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11111) );
  NAND2_X1 U14433 ( .A1(n10732), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n11106) );
  NAND2_X1 U14434 ( .A1(n10733), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n11105) );
  OAI211_X1 U14435 ( .C1(n14497), .C2(n11107), .A(n11106), .B(n11105), .ZN(
        n11108) );
  INV_X1 U14436 ( .A(n11108), .ZN(n11110) );
  AOI22_X1 U14437 ( .A1(n10764), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n14444), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11109) );
  NAND4_X1 U14438 ( .A1(n11112), .A2(n11111), .A3(n11110), .A4(n11109), .ZN(
        n11118) );
  AOI22_X1 U14439 ( .A1(n10769), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n14416), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11116) );
  AOI22_X1 U14440 ( .A1(n10877), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n14503), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11115) );
  AOI22_X1 U14441 ( .A1(n14504), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n10781), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11114) );
  NAND2_X1 U14442 ( .A1(n14486), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n11113) );
  NAND4_X1 U14443 ( .A1(n11116), .A2(n11115), .A3(n11114), .A4(n11113), .ZN(
        n11117) );
  INV_X1 U14444 ( .A(n11510), .ZN(n11119) );
  NAND2_X1 U14445 ( .A1(n11119), .A2(n9735), .ZN(n11120) );
  INV_X1 U14446 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n22168) );
  NAND2_X1 U14447 ( .A1(n16752), .A2(n22168), .ZN(n11121) );
  AOI22_X1 U14448 ( .A1(n14504), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n10781), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11125) );
  NAND2_X1 U14449 ( .A1(n10877), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n11124) );
  NAND2_X1 U14450 ( .A1(n14503), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n11123) );
  NAND2_X1 U14451 ( .A1(n14486), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n11122) );
  AOI22_X1 U14452 ( .A1(n10732), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n10733), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11130) );
  NAND2_X1 U14453 ( .A1(n10758), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n11129) );
  NAND2_X1 U14454 ( .A1(n14493), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n11128) );
  INV_X1 U14455 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11126) );
  OR2_X1 U14456 ( .A1(n14497), .A2(n11126), .ZN(n11127) );
  NAND2_X1 U14457 ( .A1(n10759), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n11134) );
  NAND2_X1 U14458 ( .A1(n14477), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n11133) );
  NAND2_X1 U14459 ( .A1(n10764), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n11132) );
  NAND2_X1 U14460 ( .A1(n14444), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n11131) );
  AOI22_X1 U14461 ( .A1(n10769), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n14416), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11135) );
  NAND4_X1 U14462 ( .A1(n11138), .A2(n11137), .A3(n11136), .A4(n11135), .ZN(
        n11514) );
  INV_X1 U14463 ( .A(n11141), .ZN(n11140) );
  INV_X1 U14464 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n17025) );
  AND2_X1 U14465 ( .A1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16912) );
  NAND2_X1 U14466 ( .A1(n16912), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n16893) );
  NAND2_X1 U14467 ( .A1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n11144) );
  NOR2_X1 U14468 ( .A1(n16893), .A2(n11144), .ZN(n16861) );
  AND2_X1 U14469 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n16936) );
  NAND2_X1 U14470 ( .A1(n16936), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n14761) );
  AND2_X1 U14471 ( .A1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n14760) );
  NAND2_X1 U14472 ( .A1(n14760), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11145) );
  NOR2_X1 U14473 ( .A1(n14761), .A2(n11145), .ZN(n11146) );
  NAND2_X1 U14474 ( .A1(n16861), .A2(n11146), .ZN(n16849) );
  NAND3_X1 U14475 ( .A1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n11147) );
  NAND2_X1 U14476 ( .A1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n16788) );
  NOR2_X1 U14477 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n21086) );
  OR2_X1 U14478 ( .A1(n20880), .A2(n21086), .ZN(n21110) );
  NAND2_X1 U14479 ( .A1(n21110), .A2(n21132), .ZN(n11151) );
  NAND2_X1 U14480 ( .A1(n20842), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n11152) );
  NAND2_X1 U14481 ( .A1(n10588), .A2(n11152), .ZN(n13773) );
  NAND2_X1 U14482 ( .A1(n11767), .A2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11771) );
  INV_X1 U14483 ( .A(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n16017) );
  INV_X1 U14484 ( .A(n11155), .ZN(n11791) );
  NAND2_X1 U14485 ( .A1(n11791), .A2(n10416), .ZN(n11156) );
  NAND2_X1 U14486 ( .A1(n11727), .A2(n11156), .ZN(n15943) );
  INV_X1 U14487 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n14221) );
  NAND2_X1 U14488 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n11163) );
  NAND2_X1 U14489 ( .A1(n11699), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n11162) );
  OAI211_X1 U14490 ( .C1(n13510), .C2(n14221), .A(n11163), .B(n11162), .ZN(
        n11164) );
  AOI21_X1 U14491 ( .B1(n13512), .B2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(
        n11164), .ZN(n14217) );
  AOI22_X1 U14492 ( .A1(n11699), .A2(P2_REIP_REG_5__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11166) );
  NAND2_X1 U14493 ( .A1(n11243), .A2(P2_EBX_REG_5__SCAN_IN), .ZN(n11165) );
  NAND2_X1 U14494 ( .A1(n13512), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11170) );
  AOI22_X1 U14495 ( .A1(n11699), .A2(P2_REIP_REG_6__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11168) );
  NAND2_X1 U14496 ( .A1(n11243), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n11167) );
  AND2_X1 U14497 ( .A1(n11168), .A2(n11167), .ZN(n11169) );
  AOI22_X1 U14498 ( .A1(n11699), .A2(P2_REIP_REG_8__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11174) );
  NAND2_X1 U14499 ( .A1(n11243), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n11173) );
  INV_X1 U14500 ( .A(n16196), .ZN(n11179) );
  NAND2_X1 U14501 ( .A1(n13512), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11178) );
  AOI22_X1 U14502 ( .A1(n11699), .A2(P2_REIP_REG_7__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11176) );
  NAND2_X1 U14503 ( .A1(n11243), .A2(P2_EBX_REG_7__SCAN_IN), .ZN(n11175) );
  AND2_X1 U14504 ( .A1(n11176), .A2(n11175), .ZN(n11177) );
  INV_X1 U14505 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n17006) );
  AOI22_X1 U14506 ( .A1(n11699), .A2(P2_REIP_REG_9__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11182) );
  NAND2_X1 U14507 ( .A1(n11243), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n11181) );
  INV_X1 U14508 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n11185) );
  NAND2_X1 U14509 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n11184) );
  NAND2_X1 U14510 ( .A1(n11699), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n11183) );
  OAI211_X1 U14511 ( .C1(n13510), .C2(n11185), .A(n11184), .B(n11183), .ZN(
        n11186) );
  AOI21_X1 U14512 ( .B1(n13512), .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n11186), .ZN(n14278) );
  NAND2_X1 U14513 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n11190) );
  NAND2_X1 U14514 ( .A1(n11699), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n11189) );
  OAI211_X1 U14515 ( .C1(n13510), .C2(n21982), .A(n11190), .B(n11189), .ZN(
        n11191) );
  AOI21_X1 U14516 ( .B1(n13512), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n11191), .ZN(n14310) );
  INV_X1 U14517 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n11195) );
  NAND2_X1 U14518 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n11194) );
  NAND2_X1 U14519 ( .A1(n11699), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n11193) );
  OAI211_X1 U14520 ( .C1(n13510), .C2(n11195), .A(n11194), .B(n11193), .ZN(
        n11196) );
  AOI21_X1 U14521 ( .B1(n13512), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n11196), .ZN(n16154) );
  AOI22_X1 U14522 ( .A1(n11699), .A2(P2_REIP_REG_13__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n11198) );
  NAND2_X1 U14523 ( .A1(n11243), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n11197) );
  NAND2_X1 U14524 ( .A1(n13512), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11202) );
  AOI22_X1 U14525 ( .A1(n11699), .A2(P2_REIP_REG_14__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n11200) );
  NAND2_X1 U14526 ( .A1(n11243), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n11199) );
  AND2_X1 U14527 ( .A1(n11200), .A2(n11199), .ZN(n11201) );
  NAND2_X1 U14528 ( .A1(n13512), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11208) );
  AOI22_X1 U14529 ( .A1(n11699), .A2(P2_REIP_REG_15__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), 
        .ZN(n11206) );
  NAND2_X1 U14530 ( .A1(n11243), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n11205) );
  AND2_X1 U14531 ( .A1(n11206), .A2(n11205), .ZN(n11207) );
  INV_X1 U14532 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n14773) );
  AOI22_X1 U14533 ( .A1(n11699), .A2(P2_REIP_REG_16__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), 
        .ZN(n11210) );
  NAND2_X1 U14534 ( .A1(n11243), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n11209) );
  NAND2_X1 U14535 ( .A1(n13512), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n11214) );
  AOI22_X1 U14536 ( .A1(n11699), .A2(P2_REIP_REG_17__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), 
        .ZN(n11212) );
  NAND2_X1 U14537 ( .A1(n11243), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n11211) );
  AND2_X1 U14538 ( .A1(n11212), .A2(n11211), .ZN(n11213) );
  INV_X1 U14539 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n16369) );
  NAND2_X1 U14540 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n11216) );
  NAND2_X1 U14541 ( .A1(n11699), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n11215) );
  OAI211_X1 U14542 ( .C1(n13510), .C2(n16369), .A(n11216), .B(n11215), .ZN(
        n11217) );
  AOI21_X1 U14543 ( .B1(n13512), .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n11217), .ZN(n16097) );
  INV_X1 U14544 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n16864) );
  AOI22_X1 U14545 ( .A1(n11699), .A2(P2_REIP_REG_19__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), 
        .ZN(n11220) );
  NAND2_X1 U14546 ( .A1(n11243), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n11219) );
  INV_X1 U14547 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n11223) );
  NAND2_X1 U14548 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n11222) );
  NAND2_X1 U14549 ( .A1(n11699), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n11221) );
  OAI211_X1 U14550 ( .C1(n13510), .C2(n11223), .A(n11222), .B(n11221), .ZN(
        n11224) );
  AOI21_X1 U14551 ( .B1(n13512), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n11224), .ZN(n16073) );
  NAND2_X1 U14552 ( .A1(n13512), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11228) );
  AOI22_X1 U14553 ( .A1(n11699), .A2(P2_REIP_REG_21__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), 
        .ZN(n11226) );
  NAND2_X1 U14554 ( .A1(n11243), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n11225) );
  AND2_X1 U14555 ( .A1(n11226), .A2(n11225), .ZN(n11227) );
  INV_X1 U14556 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n16041) );
  NAND2_X1 U14557 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n11230) );
  NAND2_X1 U14558 ( .A1(n11699), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n11229) );
  OAI211_X1 U14559 ( .C1(n13510), .C2(n16041), .A(n11230), .B(n11229), .ZN(
        n11231) );
  AOI21_X1 U14560 ( .B1(n13512), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n11231), .ZN(n16039) );
  INV_X1 U14561 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n22170) );
  AOI22_X1 U14562 ( .A1(n11699), .A2(P2_REIP_REG_23__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), 
        .ZN(n11233) );
  NAND2_X1 U14563 ( .A1(n11243), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n11232) );
  NAND2_X1 U14564 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n11235) );
  NAND2_X1 U14565 ( .A1(n11699), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n11234) );
  OAI211_X1 U14566 ( .C1(n13510), .C2(n16342), .A(n11235), .B(n11234), .ZN(
        n11236) );
  AOI21_X1 U14567 ( .B1(n13512), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n11236), .ZN(n16014) );
  NAND2_X1 U14568 ( .A1(n13512), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11240) );
  AOI22_X1 U14569 ( .A1(n11699), .A2(P2_REIP_REG_25__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), 
        .ZN(n11238) );
  NAND2_X1 U14570 ( .A1(n11243), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n11237) );
  AND2_X1 U14571 ( .A1(n11238), .A2(n11237), .ZN(n11239) );
  INV_X1 U14572 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n12070) );
  AOI22_X1 U14573 ( .A1(n11699), .A2(P2_REIP_REG_26__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), 
        .ZN(n11242) );
  NAND2_X1 U14574 ( .A1(n11243), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n11241) );
  NAND2_X1 U14575 ( .A1(n13512), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11247) );
  AOI22_X1 U14576 ( .A1(n11699), .A2(P2_REIP_REG_27__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), 
        .ZN(n11245) );
  NAND2_X1 U14577 ( .A1(n11243), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n11244) );
  AND2_X1 U14578 ( .A1(n11245), .A2(n11244), .ZN(n11246) );
  INV_X1 U14579 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n15961) );
  NAND2_X1 U14580 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n11249) );
  NAND2_X1 U14581 ( .A1(n11699), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n11248) );
  OAI211_X1 U14582 ( .C1(n13510), .C2(n15961), .A(n11249), .B(n11248), .ZN(
        n11250) );
  AOI21_X1 U14583 ( .B1(n13512), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n11250), .ZN(n15958) );
  AOI22_X1 U14584 ( .A1(n11699), .A2(P2_REIP_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n11252) );
  NAND2_X1 U14585 ( .A1(n11243), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n11251) );
  NOR2_X1 U14586 ( .A1(n15957), .A2(n11254), .ZN(n11255) );
  INV_X1 U14587 ( .A(n16310), .ZN(n11284) );
  NOR2_X1 U14588 ( .A1(n11259), .A2(n11258), .ZN(n11260) );
  AOI21_X1 U14589 ( .B1(n10926), .B2(n11261), .A(n11260), .ZN(n11262) );
  NAND2_X1 U14590 ( .A1(n11257), .A2(n11262), .ZN(n11266) );
  OAI211_X1 U14591 ( .C1(n9736), .C2(n11264), .A(n9731), .B(n11263), .ZN(
        n11265) );
  NAND2_X1 U14592 ( .A1(n11266), .A2(n11265), .ZN(n11271) );
  INV_X1 U14593 ( .A(n11272), .ZN(n11270) );
  OAI211_X1 U14594 ( .C1(n11268), .C2(n10922), .A(n11267), .B(n9736), .ZN(
        n11269) );
  NAND3_X1 U14595 ( .A1(n11271), .A2(n11270), .A3(n11269), .ZN(n11274) );
  AOI21_X1 U14596 ( .B1(n11712), .B2(n11272), .A(n11276), .ZN(n11273) );
  NAND2_X1 U14597 ( .A1(n11274), .A2(n11273), .ZN(n11275) );
  MUX2_X1 U14598 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B(n11275), .S(
        P2_STATE2_REG_0__SCAN_IN), .Z(n12020) );
  NAND2_X1 U14599 ( .A1(n11277), .A2(n11276), .ZN(n11278) );
  INV_X1 U14600 ( .A(n21135), .ZN(n11280) );
  INV_X1 U14601 ( .A(n14142), .ZN(n21107) );
  NAND2_X1 U14602 ( .A1(n11280), .A2(n21107), .ZN(n11281) );
  NAND2_X1 U14603 ( .A1(n20880), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n21098) );
  INV_X1 U14604 ( .A(n21098), .ZN(n11283) );
  NAND2_X1 U14605 ( .A1(n11284), .A2(n20370), .ZN(n11286) );
  NAND2_X1 U14606 ( .A1(n17796), .A2(n20880), .ZN(n16730) );
  INV_X1 U14607 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n21076) );
  NOR2_X1 U14608 ( .A1(n16730), .A2(n21076), .ZN(n14732) );
  AOI21_X1 U14609 ( .B1(n20356), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n14732), .ZN(n11285) );
  OAI211_X1 U14610 ( .C1(n20368), .C2(n15943), .A(n11286), .B(n11285), .ZN(
        n11287) );
  AOI21_X1 U14611 ( .B1(n20357), .B2(n14735), .A(n11287), .ZN(n11459) );
  INV_X4 U14612 ( .A(n11462), .ZN(n11288) );
  INV_X1 U14613 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n11289) );
  NOR2_X1 U14614 ( .A1(P2_EBX_REG_1__SCAN_IN), .A2(P2_EBX_REG_0__SCAN_IN), 
        .ZN(n11292) );
  INV_X1 U14615 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n11293) );
  INV_X1 U14616 ( .A(n11295), .ZN(n11296) );
  MUX2_X1 U14617 ( .A(n11297), .B(P2_EBX_REG_5__SCAN_IN), .S(n11288), .Z(
        n11311) );
  INV_X1 U14618 ( .A(n11311), .ZN(n11298) );
  INV_X1 U14619 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n11299) );
  MUX2_X1 U14620 ( .A(n11510), .B(n11299), .S(n11288), .Z(n11344) );
  MUX2_X1 U14621 ( .A(n11300), .B(P2_EBX_REG_7__SCAN_IN), .S(n11288), .Z(
        n11358) );
  NAND2_X1 U14622 ( .A1(n11288), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n11355) );
  NAND2_X1 U14623 ( .A1(n11380), .A2(n21982), .ZN(n11393) );
  INV_X1 U14624 ( .A(n11360), .ZN(n11302) );
  NAND2_X1 U14625 ( .A1(n11288), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n11392) );
  INV_X1 U14626 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n11303) );
  INV_X1 U14627 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n14358) );
  NAND2_X1 U14628 ( .A1(n11303), .A2(n14358), .ZN(n11304) );
  NAND2_X1 U14629 ( .A1(n11288), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n11372) );
  OAI21_X1 U14630 ( .B1(P2_EBX_REG_19__SCAN_IN), .B2(P2_EBX_REG_18__SCAN_IN), 
        .A(n11288), .ZN(n11306) );
  INV_X1 U14631 ( .A(n11368), .ZN(n11308) );
  NOR2_X1 U14632 ( .A1(P2_EBX_REG_20__SCAN_IN), .A2(P2_EBX_REG_21__SCAN_IN), 
        .ZN(n11307) );
  NAND2_X1 U14633 ( .A1(n11308), .A2(n11307), .ZN(n11429) );
  NAND2_X1 U14634 ( .A1(n11288), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n11428) );
  NAND2_X1 U14635 ( .A1(n11288), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n11444) );
  NAND2_X1 U14636 ( .A1(n11288), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n11709) );
  XNOR2_X1 U14637 ( .A(n11710), .B(n11709), .ZN(n11309) );
  INV_X1 U14638 ( .A(n11309), .ZN(n15949) );
  NAND3_X1 U14639 ( .A1(n15949), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n11452), .ZN(n13496) );
  OAI21_X1 U14640 ( .B1(n11309), .B2(n11300), .A(n14730), .ZN(n12016) );
  XNOR2_X1 U14641 ( .A(n11310), .B(n11311), .ZN(n16237) );
  NAND2_X1 U14642 ( .A1(n11312), .A2(n16237), .ZN(n11314) );
  AOI21_X1 U14643 ( .B1(n16237), .B2(n11452), .A(n17073), .ZN(n11313) );
  INV_X1 U14644 ( .A(n11318), .ZN(n11321) );
  INV_X1 U14645 ( .A(n11319), .ZN(n11320) );
  NAND2_X1 U14646 ( .A1(n11321), .A2(n11320), .ZN(n11322) );
  NAND2_X1 U14647 ( .A1(n11317), .A2(n11322), .ZN(n16263) );
  MUX2_X1 U14648 ( .A(n11323), .B(P2_EBX_REG_0__SCAN_IN), .S(n11288), .Z(
        n16298) );
  NAND2_X1 U14649 ( .A1(n16298), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13770) );
  INV_X1 U14650 ( .A(n11329), .ZN(n11325) );
  NAND3_X1 U14651 ( .A1(n11288), .A2(P2_EBX_REG_0__SCAN_IN), .A3(
        P2_EBX_REG_1__SCAN_IN), .ZN(n11324) );
  NAND2_X1 U14652 ( .A1(n11325), .A2(n11324), .ZN(n16289) );
  INV_X1 U14653 ( .A(n16289), .ZN(n11326) );
  XNOR2_X1 U14654 ( .A(n13770), .B(n11326), .ZN(n13766) );
  NAND2_X1 U14655 ( .A1(n13766), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17113) );
  INV_X1 U14656 ( .A(n13770), .ZN(n11327) );
  NAND2_X1 U14657 ( .A1(n11327), .A2(n11326), .ZN(n11328) );
  NAND2_X1 U14658 ( .A1(n17113), .A2(n11328), .ZN(n11332) );
  XNOR2_X1 U14659 ( .A(n11330), .B(n11329), .ZN(n16275) );
  XNOR2_X1 U14660 ( .A(n11332), .B(n16275), .ZN(n14693) );
  NAND2_X1 U14661 ( .A1(n14693), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n14711) );
  INV_X1 U14662 ( .A(n16275), .ZN(n11331) );
  NAND2_X1 U14663 ( .A1(n11332), .A2(n11331), .ZN(n11333) );
  AND2_X1 U14664 ( .A1(n14711), .A2(n11333), .ZN(n17086) );
  XNOR2_X1 U14665 ( .A(n11317), .B(n11334), .ZN(n17088) );
  AND2_X1 U14666 ( .A1(n17088), .A2(n17097), .ZN(n11336) );
  AOI21_X1 U14667 ( .B1(n17086), .B2(n17751), .A(n11336), .ZN(n11335) );
  INV_X1 U14668 ( .A(n17086), .ZN(n17728) );
  INV_X1 U14669 ( .A(n11336), .ZN(n11337) );
  AND2_X1 U14670 ( .A1(n11337), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11338) );
  INV_X1 U14671 ( .A(n17088), .ZN(n16250) );
  AOI22_X1 U14672 ( .A1(n17728), .A2(n11338), .B1(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n16250), .ZN(n11339) );
  AND2_X1 U14673 ( .A1(n16237), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11340) );
  OAI21_X1 U14674 ( .B1(n11300), .B2(n17073), .A(n16237), .ZN(n11341) );
  OAI21_X1 U14675 ( .B1(n16237), .B2(n17073), .A(n11341), .ZN(n11342) );
  INV_X2 U14676 ( .A(n11300), .ZN(n11452) );
  XNOR2_X1 U14677 ( .A(n11345), .B(n11344), .ZN(n16221) );
  NAND2_X1 U14678 ( .A1(n11351), .A2(n11347), .ZN(n11348) );
  INV_X1 U14679 ( .A(n11354), .ZN(n11356) );
  NAND2_X1 U14680 ( .A1(n11356), .A2(n10632), .ZN(n11357) );
  NAND2_X1 U14681 ( .A1(n11353), .A2(n11357), .ZN(n16208) );
  NOR2_X1 U14682 ( .A1(n16208), .A2(n11300), .ZN(n11389) );
  NAND2_X1 U14683 ( .A1(n11389), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16723) );
  INV_X1 U14684 ( .A(n11358), .ZN(n11359) );
  XNOR2_X1 U14685 ( .A(n11360), .B(n11359), .ZN(n11388) );
  NAND2_X1 U14686 ( .A1(n11388), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16742) );
  INV_X1 U14687 ( .A(n11362), .ZN(n11373) );
  NAND2_X1 U14688 ( .A1(n11362), .A2(n16369), .ZN(n11365) );
  NAND2_X1 U14689 ( .A1(n16113), .A2(n11452), .ZN(n11420) );
  NAND2_X1 U14690 ( .A1(n11420), .A2(n22065), .ZN(n16615) );
  NAND3_X1 U14691 ( .A1(n11365), .A2(n11288), .A3(P2_EBX_REG_19__SCAN_IN), 
        .ZN(n11366) );
  NAND2_X1 U14692 ( .A1(n16085), .A2(n11452), .ZN(n11418) );
  NAND2_X1 U14693 ( .A1(n11418), .A2(n16864), .ZN(n12095) );
  NAND2_X1 U14694 ( .A1(n16615), .A2(n12095), .ZN(n16587) );
  NAND2_X1 U14695 ( .A1(n11288), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n11367) );
  XNOR2_X1 U14696 ( .A(n11368), .B(n11367), .ZN(n16079) );
  NAND2_X1 U14697 ( .A1(n16079), .A2(n11452), .ZN(n11423) );
  INV_X1 U14698 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n16860) );
  INV_X1 U14699 ( .A(n11369), .ZN(n11370) );
  NOR2_X1 U14700 ( .A1(n11371), .A2(n11370), .ZN(n16068) );
  NAND2_X1 U14701 ( .A1(n16068), .A2(n11452), .ZN(n11406) );
  INV_X1 U14702 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n16848) );
  NAND2_X1 U14703 ( .A1(n11406), .A2(n16848), .ZN(n16590) );
  NAND2_X1 U14704 ( .A1(n9819), .A2(n10622), .ZN(n11374) );
  NAND2_X1 U14705 ( .A1(n16128), .A2(n11452), .ZN(n11376) );
  INV_X1 U14706 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n11375) );
  NAND2_X1 U14707 ( .A1(n11376), .A2(n11375), .ZN(n16625) );
  NAND2_X1 U14708 ( .A1(n11288), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n11377) );
  MUX2_X1 U14709 ( .A(n11288), .B(n11377), .S(n11378), .Z(n11379) );
  OR2_X1 U14710 ( .A1(n11378), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n11397) );
  NAND2_X1 U14711 ( .A1(n11379), .A2(n11397), .ZN(n20237) );
  OR2_X1 U14712 ( .A1(n20237), .A2(n11300), .ZN(n11414) );
  NAND2_X1 U14713 ( .A1(n11414), .A2(n16942), .ZN(n16654) );
  INV_X1 U14714 ( .A(n11380), .ZN(n11385) );
  AND3_X1 U14715 ( .A1(n11385), .A2(n11288), .A3(P2_EBX_REG_11__SCAN_IN), .ZN(
        n11381) );
  NOR2_X1 U14716 ( .A1(n11382), .A2(n11381), .ZN(n16179) );
  NAND2_X1 U14717 ( .A1(n16179), .A2(n11452), .ZN(n11410) );
  INV_X1 U14718 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n22118) );
  NAND2_X1 U14719 ( .A1(n11410), .A2(n22118), .ZN(n16691) );
  AND2_X1 U14720 ( .A1(n11288), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n11383) );
  AND2_X1 U14721 ( .A1(n11386), .A2(n11385), .ZN(n16190) );
  INV_X1 U14722 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16992) );
  NAND2_X1 U14723 ( .A1(n11288), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n11387) );
  XNOR2_X1 U14724 ( .A(n11353), .B(n11387), .ZN(n20255) );
  NAND2_X1 U14725 ( .A1(n20255), .A2(n11452), .ZN(n11412) );
  NAND2_X1 U14726 ( .A1(n11412), .A2(n17006), .ZN(n16714) );
  INV_X1 U14727 ( .A(n11388), .ZN(n20274) );
  NAND2_X1 U14728 ( .A1(n20274), .A2(n22145), .ZN(n16741) );
  INV_X1 U14729 ( .A(n11389), .ZN(n11390) );
  NAND2_X1 U14730 ( .A1(n11390), .A2(n17025), .ZN(n16722) );
  NAND2_X1 U14731 ( .A1(n11393), .A2(n10636), .ZN(n11394) );
  NAND2_X1 U14732 ( .A1(n11391), .A2(n11394), .ZN(n16165) );
  OR2_X1 U14733 ( .A1(n16165), .A2(n11300), .ZN(n11395) );
  INV_X1 U14734 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n16955) );
  NOR2_X1 U14735 ( .A1(n12097), .A2(n12098), .ZN(n11399) );
  AND2_X1 U14736 ( .A1(n11288), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n11396) );
  INV_X1 U14737 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16924) );
  XNOR2_X1 U14738 ( .A(n11391), .B(n10678), .ZN(n16142) );
  NAND2_X1 U14739 ( .A1(n16142), .A2(n11452), .ZN(n11416) );
  NAND2_X1 U14740 ( .A1(n11416), .A2(n16667), .ZN(n16662) );
  AND2_X1 U14741 ( .A1(n11288), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n11400) );
  NAND2_X1 U14742 ( .A1(n20220), .A2(n11452), .ZN(n11403) );
  XNOR2_X1 U14743 ( .A(n11403), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14763) );
  NAND2_X1 U14744 ( .A1(n11405), .A2(n11404), .ZN(n11426) );
  INV_X1 U14745 ( .A(n11406), .ZN(n11407) );
  AND2_X1 U14746 ( .A1(n11452), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n11408) );
  NAND2_X1 U14747 ( .A1(n16128), .A2(n11408), .ZN(n16624) );
  AND2_X1 U14748 ( .A1(n11452), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11409) );
  NAND2_X1 U14749 ( .A1(n20220), .A2(n11409), .ZN(n12100) );
  OR2_X1 U14750 ( .A1(n11410), .A2(n22118), .ZN(n16692) );
  NAND2_X1 U14751 ( .A1(n11411), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n16702) );
  AND2_X1 U14752 ( .A1(n16702), .A2(n16715), .ZN(n16689) );
  AND2_X1 U14753 ( .A1(n16692), .A2(n16689), .ZN(n12096) );
  NAND2_X1 U14754 ( .A1(n11452), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11413) );
  OR3_X1 U14755 ( .A1(n16165), .A2(n11300), .A3(n16955), .ZN(n16675) );
  AND4_X1 U14756 ( .A1(n12100), .A2(n12096), .A3(n16646), .A4(n16675), .ZN(
        n11417) );
  INV_X1 U14757 ( .A(n11414), .ZN(n11415) );
  NAND2_X1 U14758 ( .A1(n11415), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n16655) );
  OR2_X1 U14759 ( .A1(n11416), .A2(n16667), .ZN(n16663) );
  AND4_X1 U14760 ( .A1(n16624), .A2(n11417), .A3(n16655), .A4(n16663), .ZN(
        n11422) );
  INV_X1 U14761 ( .A(n11418), .ZN(n11419) );
  NAND2_X1 U14762 ( .A1(n11419), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n16588) );
  INV_X1 U14763 ( .A(n11420), .ZN(n11421) );
  INV_X1 U14764 ( .A(n11423), .ZN(n11424) );
  NAND2_X1 U14765 ( .A1(n11429), .A2(n10221), .ZN(n11430) );
  AOI21_X1 U14766 ( .B1(n16046), .B2(n11452), .A(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n16576) );
  NAND3_X1 U14767 ( .A1(n16046), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        n11452), .ZN(n16577) );
  NAND2_X1 U14768 ( .A1(n11427), .A2(n11432), .ZN(n11433) );
  NAND2_X1 U14769 ( .A1(n16036), .A2(n11452), .ZN(n11434) );
  XNOR2_X1 U14770 ( .A(n11434), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n16569) );
  INV_X1 U14771 ( .A(n16036), .ZN(n11435) );
  INV_X1 U14772 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n16813) );
  NAND2_X1 U14773 ( .A1(n11436), .A2(n11452), .ZN(n16561) );
  OAI211_X1 U14774 ( .C1(n11438), .C2(P2_EBX_REG_25__SCAN_IN), .A(
        P2_EBX_REG_26__SCAN_IN), .B(n11288), .ZN(n11439) );
  NOR3_X1 U14775 ( .A1(n11440), .A2(n11300), .A3(n12070), .ZN(n11455) );
  INV_X1 U14776 ( .A(n11440), .ZN(n15993) );
  AOI21_X1 U14777 ( .B1(n15993), .B2(n11452), .A(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n11441) );
  INV_X1 U14778 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n16554) );
  NAND2_X1 U14779 ( .A1(n16561), .A2(n16554), .ZN(n16550) );
  INV_X1 U14780 ( .A(n11444), .ZN(n11445) );
  NAND2_X1 U14781 ( .A1(n11446), .A2(n11445), .ZN(n11447) );
  NAND2_X1 U14782 ( .A1(n11449), .A2(n11447), .ZN(n15980) );
  INV_X1 U14783 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n16777) );
  INV_X1 U14784 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n22042) );
  NAND2_X1 U14785 ( .A1(n11449), .A2(n11448), .ZN(n11450) );
  AND2_X1 U14786 ( .A1(n11451), .A2(n11450), .ZN(n15960) );
  NAND2_X1 U14787 ( .A1(n15960), .A2(n11452), .ZN(n16525) );
  AOI21_X1 U14788 ( .B1(n22042), .B2(n16777), .A(n16525), .ZN(n11454) );
  INV_X1 U14789 ( .A(n16525), .ZN(n11453) );
  NOR2_X1 U14790 ( .A1(n16561), .A2(n16554), .ZN(n16551) );
  NOR2_X1 U14791 ( .A1(n11455), .A2(n16551), .ZN(n16523) );
  NAND2_X1 U14792 ( .A1(n9832), .A2(n11457), .ZN(n11458) );
  NAND2_X1 U14793 ( .A1(n11459), .A2(n11458), .ZN(P2_U2985) );
  NOR2_X1 U14794 ( .A1(n13819), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n11472) );
  AOI22_X1 U14795 ( .A1(n9737), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B1(
        n11689), .B2(P2_EAX_REG_30__SCAN_IN), .ZN(n11461) );
  AND2_X1 U14796 ( .A1(n11467), .A2(n21106), .ZN(n13784) );
  NAND2_X1 U14797 ( .A1(n11465), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n11460) );
  AND2_X1 U14798 ( .A1(n11461), .A2(n11460), .ZN(n11696) );
  NAND2_X1 U14799 ( .A1(n13784), .A2(n11462), .ZN(n11478) );
  NAND2_X1 U14800 ( .A1(n9737), .A2(n13818), .ZN(n11487) );
  MUX2_X1 U14801 ( .A(n13819), .B(n21114), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n11463) );
  NAND2_X1 U14802 ( .A1(n9738), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n11470) );
  NAND2_X1 U14803 ( .A1(n9722), .A2(P2_EAX_REG_0__SCAN_IN), .ZN(n11466) );
  OAI211_X1 U14804 ( .C1(n11467), .C2(n17130), .A(n11466), .B(n21106), .ZN(
        n11468) );
  INV_X1 U14805 ( .A(n11468), .ZN(n11469) );
  NAND2_X1 U14806 ( .A1(n11470), .A2(n11469), .ZN(n13792) );
  NAND2_X1 U14807 ( .A1(n13791), .A2(n13792), .ZN(n11484) );
  INV_X1 U14808 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n21031) );
  NAND2_X1 U14809 ( .A1(n9737), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11474) );
  NAND2_X1 U14810 ( .A1(n11472), .A2(P2_EAX_REG_1__SCAN_IN), .ZN(n11473) );
  OAI211_X2 U14811 ( .C1(n11475), .C2(n21031), .A(n11474), .B(n11473), .ZN(
        n11482) );
  XNOR2_X1 U14812 ( .A(n11484), .B(n11482), .ZN(n16281) );
  NAND2_X1 U14813 ( .A1(n11476), .A2(n13819), .ZN(n11477) );
  MUX2_X1 U14814 ( .A(n11477), .B(n20837), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n11481) );
  INV_X2 U14815 ( .A(n11478), .ZN(n11655) );
  NAND2_X1 U14816 ( .A1(n11655), .A2(n11479), .ZN(n11480) );
  AND2_X1 U14817 ( .A1(n11481), .A2(n11480), .ZN(n16280) );
  INV_X1 U14818 ( .A(n11482), .ZN(n11483) );
  NAND2_X1 U14819 ( .A1(n11484), .A2(n11483), .ZN(n11485) );
  NAND2_X1 U14820 ( .A1(n11655), .A2(n11486), .ZN(n11488) );
  OAI211_X1 U14821 ( .C1(n21106), .C2(n22183), .A(n11488), .B(n11487), .ZN(
        n11491) );
  XNOR2_X1 U14822 ( .A(n11493), .B(n11491), .ZN(n14699) );
  AOI22_X1 U14823 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n11688), .B1(
        n11689), .B2(P2_EAX_REG_2__SCAN_IN), .ZN(n11490) );
  NAND2_X1 U14824 ( .A1(n11465), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n11489) );
  AND2_X1 U14825 ( .A1(n11490), .A2(n11489), .ZN(n14698) );
  NAND2_X2 U14826 ( .A1(n14699), .A2(n14698), .ZN(n14701) );
  INV_X1 U14827 ( .A(n11491), .ZN(n11492) );
  NAND2_X1 U14828 ( .A1(n11493), .A2(n11492), .ZN(n11494) );
  AOI22_X1 U14829 ( .A1(n11688), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n11499) );
  NAND2_X1 U14830 ( .A1(n9739), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n11498) );
  NAND2_X1 U14831 ( .A1(n11655), .A2(n11495), .ZN(n11497) );
  NAND2_X1 U14832 ( .A1(n11689), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n11496) );
  INV_X1 U14833 ( .A(n16254), .ZN(n11500) );
  AOI22_X1 U14834 ( .A1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n11688), .B1(
        n11689), .B2(P2_EAX_REG_4__SCAN_IN), .ZN(n11504) );
  NAND2_X1 U14835 ( .A1(n11465), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n11503) );
  NAND2_X1 U14836 ( .A1(n11655), .A2(n11501), .ZN(n11502) );
  NAND2_X1 U14837 ( .A1(n11465), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n11509) );
  NAND2_X1 U14838 ( .A1(n11655), .A2(n11505), .ZN(n11508) );
  NAND2_X1 U14839 ( .A1(n11688), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11507) );
  NAND2_X1 U14840 ( .A1(n11689), .A2(P2_EAX_REG_5__SCAN_IN), .ZN(n11506) );
  NAND4_X1 U14841 ( .A1(n11509), .A2(n11508), .A3(n11507), .A4(n11506), .ZN(
        n16224) );
  NAND2_X1 U14842 ( .A1(n16225), .A2(n16224), .ZN(n16227) );
  NAND2_X1 U14843 ( .A1(n11655), .A2(n11510), .ZN(n11511) );
  INV_X1 U14844 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n21040) );
  NAND2_X1 U14845 ( .A1(n11688), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11513) );
  NAND2_X1 U14846 ( .A1(n11689), .A2(P2_EAX_REG_6__SCAN_IN), .ZN(n11512) );
  OAI211_X1 U14847 ( .C1(n11475), .C2(n21040), .A(n11513), .B(n11512), .ZN(
        n13823) );
  NAND2_X1 U14848 ( .A1(n13822), .A2(n13823), .ZN(n11516) );
  NAND2_X1 U14849 ( .A1(n11655), .A2(n11514), .ZN(n11515) );
  INV_X1 U14850 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n21042) );
  NAND2_X1 U14851 ( .A1(n11688), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11518) );
  NAND2_X1 U14852 ( .A1(n11689), .A2(P2_EAX_REG_7__SCAN_IN), .ZN(n11517) );
  OAI211_X1 U14853 ( .C1(n11475), .C2(n21042), .A(n11518), .B(n11517), .ZN(
        n13810) );
  AOI22_X1 U14854 ( .A1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n11688), .B1(
        n11689), .B2(P2_EAX_REG_8__SCAN_IN), .ZN(n11535) );
  AOI22_X1 U14855 ( .A1(n10758), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n14493), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11526) );
  AOI22_X1 U14856 ( .A1(n10759), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n14477), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11525) );
  INV_X1 U14857 ( .A(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11521) );
  NAND2_X1 U14858 ( .A1(n10732), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n11520) );
  NAND2_X1 U14859 ( .A1(n10733), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n11519) );
  OAI211_X1 U14860 ( .C1(n14497), .C2(n11521), .A(n11520), .B(n11519), .ZN(
        n11522) );
  INV_X1 U14861 ( .A(n11522), .ZN(n11524) );
  AOI22_X1 U14862 ( .A1(n10764), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n14444), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11523) );
  NAND4_X1 U14863 ( .A1(n11526), .A2(n11525), .A3(n11524), .A4(n11523), .ZN(
        n11532) );
  AOI22_X1 U14864 ( .A1(n10769), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n14416), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11530) );
  AOI22_X1 U14865 ( .A1(n14486), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10877), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11529) );
  AOI22_X1 U14866 ( .A1(n14504), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10781), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11528) );
  NAND2_X1 U14867 ( .A1(n14503), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n11527) );
  NAND4_X1 U14868 ( .A1(n11530), .A2(n11529), .A3(n11528), .A4(n11527), .ZN(
        n11531) );
  NAND2_X1 U14869 ( .A1(n11655), .A2(n14335), .ZN(n11534) );
  NAND2_X1 U14870 ( .A1(n11465), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n11533) );
  AOI22_X1 U14871 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n9737), .B1(
        n11689), .B2(P2_EAX_REG_9__SCAN_IN), .ZN(n11552) );
  AOI22_X1 U14872 ( .A1(n10758), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n14493), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11543) );
  AOI22_X1 U14873 ( .A1(n10759), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n14477), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11542) );
  INV_X1 U14874 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11538) );
  NAND2_X1 U14875 ( .A1(n10732), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n11537) );
  NAND2_X1 U14876 ( .A1(n10733), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n11536) );
  OAI211_X1 U14877 ( .C1(n14497), .C2(n11538), .A(n11537), .B(n11536), .ZN(
        n11539) );
  INV_X1 U14878 ( .A(n11539), .ZN(n11541) );
  AOI22_X1 U14879 ( .A1(n10764), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n14444), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11540) );
  NAND4_X1 U14880 ( .A1(n11543), .A2(n11542), .A3(n11541), .A4(n11540), .ZN(
        n11549) );
  AOI22_X1 U14881 ( .A1(n10769), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n14416), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11547) );
  AOI22_X1 U14882 ( .A1(n10877), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n14503), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11546) );
  AOI22_X1 U14883 ( .A1(n14504), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n10781), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11545) );
  NAND2_X1 U14884 ( .A1(n14486), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11544) );
  NAND4_X1 U14885 ( .A1(n11547), .A2(n11546), .A3(n11545), .A4(n11544), .ZN(
        n11548) );
  NAND2_X1 U14886 ( .A1(n11655), .A2(n14336), .ZN(n11551) );
  NAND2_X1 U14887 ( .A1(n11465), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n11550) );
  INV_X1 U14888 ( .A(n13919), .ZN(n11572) );
  AOI22_X1 U14889 ( .A1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n9737), .B1(
        n11689), .B2(P2_EAX_REG_10__SCAN_IN), .ZN(n11570) );
  AOI22_X1 U14890 ( .A1(n10758), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n14493), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11561) );
  AOI22_X1 U14891 ( .A1(n10759), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n14477), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11560) );
  INV_X1 U14892 ( .A(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11556) );
  NAND2_X1 U14893 ( .A1(n14504), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n11555) );
  NAND2_X1 U14894 ( .A1(n10732), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n11554) );
  OAI211_X1 U14895 ( .C1(n14497), .C2(n11556), .A(n11555), .B(n11554), .ZN(
        n11557) );
  INV_X1 U14896 ( .A(n11557), .ZN(n11559) );
  AOI22_X1 U14897 ( .A1(n10764), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n14444), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11558) );
  NAND4_X1 U14898 ( .A1(n11561), .A2(n11560), .A3(n11559), .A4(n11558), .ZN(
        n11567) );
  AOI22_X1 U14899 ( .A1(n10769), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n14416), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11565) );
  AOI22_X1 U14900 ( .A1(n10877), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n14503), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11564) );
  AOI22_X1 U14901 ( .A1(n10781), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n10733), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11563) );
  NAND2_X1 U14902 ( .A1(n14486), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n11562) );
  NAND4_X1 U14903 ( .A1(n11565), .A2(n11564), .A3(n11563), .A4(n11562), .ZN(
        n11566) );
  NAND2_X1 U14904 ( .A1(n11655), .A2(n14319), .ZN(n11569) );
  NAND2_X1 U14905 ( .A1(n11465), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n11568) );
  NAND2_X1 U14906 ( .A1(n11572), .A2(n11571), .ZN(n14005) );
  AOI22_X1 U14907 ( .A1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n9737), .B1(
        n11689), .B2(P2_EAX_REG_11__SCAN_IN), .ZN(n11589) );
  AOI22_X1 U14908 ( .A1(n10758), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n14493), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11580) );
  AOI22_X1 U14909 ( .A1(n10759), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n14477), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11579) );
  INV_X1 U14910 ( .A(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11575) );
  NAND2_X1 U14911 ( .A1(n10732), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n11574) );
  NAND2_X1 U14912 ( .A1(n10733), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n11573) );
  OAI211_X1 U14913 ( .C1(n14497), .C2(n11575), .A(n11574), .B(n11573), .ZN(
        n11576) );
  INV_X1 U14914 ( .A(n11576), .ZN(n11578) );
  AOI22_X1 U14915 ( .A1(n10764), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n14444), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11577) );
  NAND4_X1 U14916 ( .A1(n11580), .A2(n11579), .A3(n11578), .A4(n11577), .ZN(
        n11586) );
  AOI22_X1 U14917 ( .A1(n10769), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n14416), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11584) );
  AOI22_X1 U14918 ( .A1(n10877), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n14503), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11583) );
  AOI22_X1 U14919 ( .A1(n14504), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10781), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11582) );
  NAND2_X1 U14920 ( .A1(n14486), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n11581) );
  NAND4_X1 U14921 ( .A1(n11584), .A2(n11583), .A3(n11582), .A4(n11581), .ZN(
        n11585) );
  NAND2_X1 U14922 ( .A1(n11655), .A2(n14320), .ZN(n11588) );
  NAND2_X1 U14923 ( .A1(n11465), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n11587) );
  NAND2_X1 U14924 ( .A1(n11465), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n11607) );
  AOI22_X1 U14925 ( .A1(n10758), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n14477), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11597) );
  AOI22_X1 U14926 ( .A1(n14493), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10759), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11596) );
  INV_X1 U14927 ( .A(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11592) );
  NAND2_X1 U14928 ( .A1(n10732), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n11591) );
  NAND2_X1 U14929 ( .A1(n10733), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n11590) );
  OAI211_X1 U14930 ( .C1(n14497), .C2(n11592), .A(n11591), .B(n11590), .ZN(
        n11593) );
  INV_X1 U14931 ( .A(n11593), .ZN(n11595) );
  AOI22_X1 U14932 ( .A1(n10764), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n14444), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11594) );
  NAND4_X1 U14933 ( .A1(n11597), .A2(n11596), .A3(n11595), .A4(n11594), .ZN(
        n11603) );
  AOI22_X1 U14934 ( .A1(n10769), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n14416), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11601) );
  AOI22_X1 U14935 ( .A1(n10877), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n14503), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11600) );
  AOI22_X1 U14936 ( .A1(n14504), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n10781), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11599) );
  NAND2_X1 U14937 ( .A1(n14486), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n11598) );
  NAND4_X1 U14938 ( .A1(n11601), .A2(n11600), .A3(n11599), .A4(n11598), .ZN(
        n11602) );
  NAND2_X1 U14939 ( .A1(n11655), .A2(n16382), .ZN(n11606) );
  NAND2_X1 U14940 ( .A1(n11688), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n11605) );
  NAND2_X1 U14941 ( .A1(n11689), .A2(P2_EAX_REG_12__SCAN_IN), .ZN(n11604) );
  NAND4_X1 U14942 ( .A1(n11607), .A2(n11606), .A3(n11605), .A4(n11604), .ZN(
        n14148) );
  NAND2_X1 U14943 ( .A1(n14085), .A2(n14148), .ZN(n14147) );
  AOI22_X1 U14944 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n9737), .B1(
        n11689), .B2(P2_EAX_REG_13__SCAN_IN), .ZN(n11624) );
  AOI22_X1 U14945 ( .A1(n10758), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n14493), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11615) );
  AOI22_X1 U14946 ( .A1(n10759), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n14477), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11614) );
  INV_X1 U14947 ( .A(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11610) );
  NAND2_X1 U14948 ( .A1(n10732), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n11609) );
  NAND2_X1 U14949 ( .A1(n10733), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n11608) );
  OAI211_X1 U14950 ( .C1(n14497), .C2(n11610), .A(n11609), .B(n11608), .ZN(
        n11611) );
  INV_X1 U14951 ( .A(n11611), .ZN(n11613) );
  AOI22_X1 U14952 ( .A1(n10764), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n14444), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11612) );
  NAND4_X1 U14953 ( .A1(n11615), .A2(n11614), .A3(n11613), .A4(n11612), .ZN(
        n11621) );
  AOI22_X1 U14954 ( .A1(n10769), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n14416), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11619) );
  AOI22_X1 U14955 ( .A1(n10877), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n14503), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11618) );
  AOI22_X1 U14956 ( .A1(n14504), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10781), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11617) );
  NAND2_X1 U14957 ( .A1(n14486), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n11616) );
  NAND4_X1 U14958 ( .A1(n11619), .A2(n11618), .A3(n11617), .A4(n11616), .ZN(
        n11620) );
  NAND2_X1 U14959 ( .A1(n11655), .A2(n14345), .ZN(n11623) );
  NAND2_X1 U14960 ( .A1(n9739), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n11622) );
  AOI22_X1 U14961 ( .A1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n9737), .B1(
        n11689), .B2(P2_EAX_REG_14__SCAN_IN), .ZN(n11641) );
  AOI22_X1 U14962 ( .A1(n10758), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n14493), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11632) );
  AOI22_X1 U14963 ( .A1(n10759), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n14477), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11631) );
  INV_X1 U14964 ( .A(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11627) );
  NAND2_X1 U14965 ( .A1(n14504), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n11626) );
  NAND2_X1 U14966 ( .A1(n10732), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n11625) );
  OAI211_X1 U14967 ( .C1(n14497), .C2(n11627), .A(n11626), .B(n11625), .ZN(
        n11628) );
  INV_X1 U14968 ( .A(n11628), .ZN(n11630) );
  AOI22_X1 U14969 ( .A1(n10769), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10764), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11629) );
  NAND4_X1 U14970 ( .A1(n11632), .A2(n11631), .A3(n11630), .A4(n11629), .ZN(
        n11638) );
  AOI22_X1 U14971 ( .A1(n14416), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n14444), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11636) );
  AOI22_X1 U14972 ( .A1(n10877), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n14503), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11635) );
  AOI22_X1 U14973 ( .A1(n10781), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n10733), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11634) );
  NAND2_X1 U14974 ( .A1(n14486), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n11633) );
  NAND4_X1 U14975 ( .A1(n11636), .A2(n11635), .A3(n11634), .A4(n11633), .ZN(
        n11637) );
  NAND2_X1 U14976 ( .A1(n11655), .A2(n14323), .ZN(n11640) );
  NAND2_X1 U14977 ( .A1(n11465), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n11639) );
  NAND2_X1 U14978 ( .A1(n11465), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n11659) );
  AOI22_X1 U14979 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n10758), .B1(
        n14493), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11648) );
  AOI22_X1 U14980 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n14477), .B1(
        n10759), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11647) );
  INV_X1 U14981 ( .A(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n14656) );
  NAND2_X1 U14982 ( .A1(n10732), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n11643) );
  NAND2_X1 U14983 ( .A1(n10733), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n11642) );
  OAI211_X1 U14984 ( .C1(n14497), .C2(n14656), .A(n11643), .B(n11642), .ZN(
        n11644) );
  INV_X1 U14985 ( .A(n11644), .ZN(n11646) );
  AOI22_X1 U14986 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n14444), .B1(
        n10764), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11645) );
  NAND4_X1 U14987 ( .A1(n11648), .A2(n11647), .A3(n11646), .A4(n11645), .ZN(
        n11654) );
  AOI22_X1 U14988 ( .A1(n10769), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n14416), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11652) );
  AOI22_X1 U14989 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n14503), .B1(
        n10877), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11651) );
  AOI22_X1 U14990 ( .A1(n14504), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n10781), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11650) );
  NAND2_X1 U14991 ( .A1(n14486), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n11649) );
  NAND4_X1 U14992 ( .A1(n11652), .A2(n11651), .A3(n11650), .A4(n11649), .ZN(
        n11653) );
  NAND2_X1 U14993 ( .A1(n11655), .A2(n9861), .ZN(n11658) );
  NAND2_X1 U14994 ( .A1(n11688), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11657) );
  NAND2_X1 U14995 ( .A1(n11689), .A2(P2_EAX_REG_15__SCAN_IN), .ZN(n11656) );
  NAND4_X1 U14996 ( .A1(n11659), .A2(n11658), .A3(n11657), .A4(n11656), .ZN(
        n14360) );
  INV_X1 U14997 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n21056) );
  NAND2_X1 U14998 ( .A1(n11688), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11661) );
  NAND2_X1 U14999 ( .A1(n11689), .A2(P2_EAX_REG_16__SCAN_IN), .ZN(n11660) );
  OAI211_X1 U15000 ( .C1(n11475), .C2(n21056), .A(n11661), .B(n11660), .ZN(
        n14767) );
  NAND2_X1 U15001 ( .A1(n14359), .A2(n14767), .ZN(n14766) );
  AOI22_X1 U15002 ( .A1(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n9737), .B1(
        n11689), .B2(P2_EAX_REG_17__SCAN_IN), .ZN(n11663) );
  NAND2_X1 U15003 ( .A1(n9739), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n11662) );
  INV_X1 U15004 ( .A(n16119), .ZN(n11664) );
  AOI22_X1 U15005 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n9737), .B1(
        n11689), .B2(P2_EAX_REG_18__SCAN_IN), .ZN(n11666) );
  NAND2_X1 U15006 ( .A1(n9739), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n11665) );
  INV_X1 U15007 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n21061) );
  NAND2_X1 U15008 ( .A1(n9737), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11668) );
  NAND2_X1 U15009 ( .A1(n11689), .A2(P2_EAX_REG_19__SCAN_IN), .ZN(n11667) );
  OAI211_X1 U15010 ( .C1(n11475), .C2(n21061), .A(n11668), .B(n11667), .ZN(
        n16083) );
  INV_X1 U15011 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n16606) );
  NAND2_X1 U15012 ( .A1(n9737), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11670) );
  NAND2_X1 U15013 ( .A1(n11689), .A2(P2_EAX_REG_20__SCAN_IN), .ZN(n11669) );
  OAI211_X1 U15014 ( .C1(n11475), .C2(n16606), .A(n11670), .B(n11669), .ZN(
        n16072) );
  NAND2_X1 U15015 ( .A1(n16071), .A2(n16072), .ZN(n16056) );
  INV_X1 U15016 ( .A(n16056), .ZN(n11674) );
  AOI22_X1 U15017 ( .A1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n9737), .B1(
        n11689), .B2(P2_EAX_REG_21__SCAN_IN), .ZN(n11672) );
  NAND2_X1 U15018 ( .A1(n11465), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n11671) );
  AOI22_X1 U15019 ( .A1(n11688), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B1(
        n11689), .B2(P2_EAX_REG_22__SCAN_IN), .ZN(n11676) );
  NAND2_X1 U15020 ( .A1(n9739), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n11675) );
  AND2_X1 U15021 ( .A1(n11676), .A2(n11675), .ZN(n16050) );
  AOI22_X1 U15022 ( .A1(n9737), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B1(
        n11689), .B2(P2_EAX_REG_23__SCAN_IN), .ZN(n11678) );
  NAND2_X1 U15023 ( .A1(n11465), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n11677) );
  INV_X1 U15024 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n11681) );
  NAND2_X1 U15025 ( .A1(n9737), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11680) );
  NAND2_X1 U15026 ( .A1(n11689), .A2(P2_EAX_REG_24__SCAN_IN), .ZN(n11679) );
  OAI211_X1 U15027 ( .C1(n11475), .C2(n11681), .A(n11680), .B(n11679), .ZN(
        n16010) );
  AOI22_X1 U15028 ( .A1(n9737), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .B1(
        n11689), .B2(P2_EAX_REG_25__SCAN_IN), .ZN(n11683) );
  NAND2_X1 U15029 ( .A1(n9739), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n11682) );
  AOI22_X1 U15030 ( .A1(n9737), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .B1(
        n11689), .B2(P2_EAX_REG_26__SCAN_IN), .ZN(n11685) );
  NAND2_X1 U15031 ( .A1(n11465), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n11684) );
  INV_X1 U15032 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n21074) );
  NAND2_X1 U15033 ( .A1(n11688), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11687) );
  NAND2_X1 U15034 ( .A1(n11689), .A2(P2_EAX_REG_27__SCAN_IN), .ZN(n11686) );
  OAI211_X1 U15035 ( .C1(n11475), .C2(n21074), .A(n11687), .B(n11686), .ZN(
        n15970) );
  INV_X1 U15036 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n16528) );
  NAND2_X1 U15037 ( .A1(n11688), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11691) );
  NAND2_X1 U15038 ( .A1(n11689), .A2(P2_EAX_REG_28__SCAN_IN), .ZN(n11690) );
  OAI211_X1 U15039 ( .C1(n11475), .C2(n16528), .A(n11691), .B(n11690), .ZN(
        n15953) );
  AOI22_X1 U15040 ( .A1(n9737), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .B1(
        n11689), .B2(P2_EAX_REG_29__SCAN_IN), .ZN(n11693) );
  NAND2_X1 U15041 ( .A1(n9739), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n11692) );
  INV_X1 U15042 ( .A(n14725), .ZN(n11695) );
  INV_X1 U15043 ( .A(n11696), .ZN(n11694) );
  AND2_X2 U15044 ( .A1(n14725), .A2(n11694), .ZN(n13508) );
  AOI21_X2 U15045 ( .B1(n11696), .B2(n11695), .A(n13508), .ZN(n14681) );
  NAND2_X1 U15046 ( .A1(n17778), .A2(n17793), .ZN(n13615) );
  NAND2_X1 U15047 ( .A1(n21021), .A2(n21030), .ZN(n21025) );
  INV_X1 U15048 ( .A(n21025), .ZN(n21013) );
  NAND2_X1 U15049 ( .A1(n21129), .A2(n21133), .ZN(n13623) );
  OR2_X1 U15050 ( .A1(n13623), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n17794) );
  INV_X1 U15051 ( .A(n17794), .ZN(n11698) );
  NAND2_X1 U15052 ( .A1(n14681), .A2(n20244), .ZN(n11717) );
  INV_X1 U15053 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n13517) );
  AOI22_X1 U15054 ( .A1(n11699), .A2(P2_REIP_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n11701) );
  NAND2_X1 U15055 ( .A1(n11243), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n11700) );
  OR2_X1 U15056 ( .A1(n11703), .A2(n11702), .ZN(n11704) );
  INV_X1 U15057 ( .A(n17779), .ZN(n11706) );
  NAND2_X1 U15058 ( .A1(n11706), .A2(n17778), .ZN(n13813) );
  INV_X1 U15059 ( .A(n17793), .ZN(n13625) );
  NAND2_X1 U15060 ( .A1(n21133), .A2(n20842), .ZN(n11723) );
  INV_X1 U15061 ( .A(n11723), .ZN(n11707) );
  NAND2_X1 U15062 ( .A1(n11712), .A2(n11707), .ZN(n11708) );
  NAND2_X1 U15063 ( .A1(n11710), .A2(n11709), .ZN(n13500) );
  NAND2_X1 U15064 ( .A1(n11288), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n11711) );
  XNOR2_X1 U15065 ( .A(n13500), .B(n11711), .ZN(n12018) );
  NAND3_X1 U15066 ( .A1(n11712), .A2(P2_EBX_REG_31__SCAN_IN), .A3(n11723), 
        .ZN(n11713) );
  NOR3_X1 U15067 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(P2_STATEBS16_REG_SCAN_IN), .ZN(n17641) );
  NAND2_X1 U15068 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n20945), .ZN(n21003) );
  NOR3_X1 U15069 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n21106), .A3(n21003), 
        .ZN(n17792) );
  NOR2_X1 U15070 ( .A1(n20227), .A2(n17792), .ZN(n11718) );
  NAND2_X1 U15071 ( .A1(n20348), .A2(n17794), .ZN(n15930) );
  INV_X1 U15072 ( .A(n17778), .ZN(n11720) );
  OR2_X1 U15073 ( .A1(n11721), .A2(n11720), .ZN(n12036) );
  NAND2_X1 U15074 ( .A1(n9969), .A2(n17793), .ZN(n11722) );
  INV_X1 U15075 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n15931) );
  NAND3_X1 U15076 ( .A1(n13632), .A2(n15931), .A3(n11723), .ZN(n11724) );
  AOI22_X1 U15077 ( .A1(n20256), .A2(P2_REIP_REG_30__SCAN_IN), .B1(
        P2_EBX_REG_30__SCAN_IN), .B2(n20271), .ZN(n11725) );
  INV_X1 U15078 ( .A(n11725), .ZN(n11726) );
  AND2_X2 U15079 ( .A1(n20269), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20240) );
  NOR2_X1 U15080 ( .A1(n11726), .A2(n10681), .ZN(n11793) );
  XNOR2_X1 U15081 ( .A(n11727), .B(n10417), .ZN(n15928) );
  INV_X1 U15082 ( .A(n11728), .ZN(n11730) );
  NAND2_X1 U15083 ( .A1(n9854), .A2(n10429), .ZN(n11729) );
  NAND2_X1 U15084 ( .A1(n11730), .A2(n11729), .ZN(n16093) );
  NAND2_X1 U15085 ( .A1(n11154), .A2(n11758), .ZN(n11731) );
  NAND2_X1 U15086 ( .A1(n9853), .A2(n11731), .ZN(n16629) );
  NOR2_X1 U15087 ( .A1(n11732), .A2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11733) );
  OR2_X1 U15088 ( .A1(n11759), .A2(n11733), .ZN(n16645) );
  INV_X1 U15089 ( .A(n16645), .ZN(n16134) );
  INV_X1 U15090 ( .A(n11756), .ZN(n11736) );
  NAND2_X1 U15091 ( .A1(n11740), .A2(n11734), .ZN(n11735) );
  NAND2_X1 U15092 ( .A1(n11736), .A2(n11735), .ZN(n16669) );
  NAND2_X1 U15093 ( .A1(n11737), .A2(n11738), .ZN(n11739) );
  NAND2_X1 U15094 ( .A1(n11740), .A2(n11739), .ZN(n16679) );
  INV_X1 U15095 ( .A(n16679), .ZN(n16163) );
  NAND2_X1 U15096 ( .A1(n11755), .A2(n16695), .ZN(n11741) );
  AND2_X1 U15097 ( .A1(n11737), .A2(n11741), .ZN(n16697) );
  AND2_X1 U15098 ( .A1(n11748), .A2(n20259), .ZN(n11742) );
  NOR2_X1 U15099 ( .A1(n11753), .A2(n11742), .ZN(n20251) );
  OR2_X1 U15100 ( .A1(n11745), .A2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11744) );
  NAND2_X1 U15101 ( .A1(n11744), .A2(n11743), .ZN(n16757) );
  AOI21_X1 U15102 ( .B1(n17723), .B2(n11747), .A(n11745), .ZN(n17717) );
  AOI21_X1 U15103 ( .B1(n17737), .B2(n11746), .A(n10420), .ZN(n17724) );
  OAI21_X1 U15104 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n11746), .ZN(n14684) );
  MUX2_X1 U15105 ( .A(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .S(P2_STATE2_REG_0__SCAN_IN), .Z(
        n16294) );
  INV_X1 U15106 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n16286) );
  MUX2_X1 U15107 ( .A(n16286), .B(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .S(
        P2_STATE2_REG_0__SCAN_IN), .Z(n16284) );
  NOR2_X1 U15108 ( .A1(n16294), .A2(n16284), .ZN(n16269) );
  NAND2_X1 U15109 ( .A1(n14684), .A2(n16269), .ZN(n16262) );
  NOR2_X1 U15110 ( .A1(n17724), .A2(n16262), .ZN(n16243) );
  OAI21_X1 U15111 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n10420), .A(
        n11747), .ZN(n20367) );
  NAND2_X1 U15112 ( .A1(n16243), .A2(n20367), .ZN(n16229) );
  NOR2_X1 U15113 ( .A1(n17717), .A2(n16229), .ZN(n16214) );
  NAND2_X1 U15114 ( .A1(n16757), .A2(n16214), .ZN(n16199) );
  INV_X1 U15115 ( .A(n16199), .ZN(n11752) );
  OAI21_X1 U15116 ( .B1(n11751), .B2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n11748), .ZN(n16732) );
  NOR2_X1 U15117 ( .A1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n11749), .ZN(
        n11750) );
  NOR2_X1 U15118 ( .A1(n11751), .A2(n11750), .ZN(n20267) );
  INV_X1 U15119 ( .A(n20267), .ZN(n16200) );
  NAND3_X1 U15120 ( .A1(n11752), .A2(n16732), .A3(n16200), .ZN(n20249) );
  NOR2_X1 U15121 ( .A1(n20251), .A2(n20249), .ZN(n16183) );
  OR2_X1 U15122 ( .A1(n11753), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11754) );
  NAND2_X1 U15123 ( .A1(n11755), .A2(n11754), .ZN(n16707) );
  NAND2_X1 U15124 ( .A1(n16183), .A2(n16707), .ZN(n16171) );
  OR2_X1 U15125 ( .A1(n16697), .A2(n16171), .ZN(n16172) );
  NOR2_X1 U15126 ( .A1(n16163), .A2(n16172), .ZN(n16145) );
  AND2_X1 U15127 ( .A1(n16669), .A2(n16145), .ZN(n20232) );
  NOR2_X1 U15128 ( .A1(n11756), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11757) );
  OR2_X1 U15129 ( .A1(n11732), .A2(n11757), .ZN(n20234) );
  NAND2_X1 U15130 ( .A1(n20232), .A2(n20234), .ZN(n16133) );
  NOR2_X1 U15131 ( .A1(n16134), .A2(n16133), .ZN(n20221) );
  OAI21_X1 U15132 ( .B1(n11759), .B2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n11758), .ZN(n20223) );
  NAND2_X1 U15133 ( .A1(n20221), .A2(n20223), .ZN(n16121) );
  INV_X1 U15134 ( .A(n16121), .ZN(n11760) );
  AND2_X1 U15135 ( .A1(n16629), .A2(n11760), .ZN(n16102) );
  INV_X1 U15136 ( .A(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n11761) );
  NAND2_X1 U15137 ( .A1(n9853), .A2(n11761), .ZN(n11762) );
  NAND2_X1 U15138 ( .A1(n9854), .A2(n11762), .ZN(n16619) );
  AND2_X1 U15139 ( .A1(n16102), .A2(n16619), .ZN(n16087) );
  NAND2_X1 U15140 ( .A1(n16093), .A2(n16087), .ZN(n11763) );
  INV_X1 U15141 ( .A(n11764), .ZN(n11765) );
  OAI21_X1 U15142 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n11728), .A(
        n11765), .ZN(n16609) );
  OAI21_X1 U15143 ( .B1(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n11764), .A(
        n11769), .ZN(n16595) );
  INV_X1 U15144 ( .A(n16595), .ZN(n11766) );
  INV_X1 U15145 ( .A(n11767), .ZN(n11772) );
  NAND2_X1 U15146 ( .A1(n11769), .A2(n11768), .ZN(n11770) );
  NAND2_X1 U15147 ( .A1(n11772), .A2(n11770), .ZN(n16583) );
  INV_X1 U15148 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n16033) );
  NAND2_X1 U15149 ( .A1(n11772), .A2(n16033), .ZN(n11773) );
  NAND2_X1 U15150 ( .A1(n11771), .A2(n11773), .ZN(n16572) );
  NAND2_X1 U15151 ( .A1(n16028), .A2(n16572), .ZN(n11774) );
  NAND2_X1 U15152 ( .A1(n11774), .A2(n20250), .ZN(n16015) );
  NAND2_X1 U15153 ( .A1(n11771), .A2(n16017), .ZN(n11775) );
  NAND2_X1 U15154 ( .A1(n11776), .A2(n11775), .ZN(n16565) );
  NAND2_X1 U15155 ( .A1(n16015), .A2(n16565), .ZN(n16000) );
  INV_X1 U15156 ( .A(n16000), .ZN(n11779) );
  NAND2_X1 U15157 ( .A1(n11776), .A2(n22107), .ZN(n11777) );
  AND2_X1 U15158 ( .A1(n11783), .A2(n11777), .ZN(n16005) );
  INV_X1 U15159 ( .A(n16005), .ZN(n11778) );
  NAND2_X1 U15160 ( .A1(n11779), .A2(n11778), .ZN(n11780) );
  NAND2_X1 U15161 ( .A1(n11780), .A2(n20250), .ZN(n15988) );
  INV_X1 U15162 ( .A(n11781), .ZN(n11786) );
  NAND2_X1 U15163 ( .A1(n11783), .A2(n11782), .ZN(n11784) );
  NAND2_X1 U15164 ( .A1(n11786), .A2(n11784), .ZN(n16548) );
  INV_X1 U15165 ( .A(n11785), .ZN(n11789) );
  INV_X1 U15166 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n16536) );
  NAND2_X1 U15167 ( .A1(n11786), .A2(n16536), .ZN(n11787) );
  AND2_X1 U15168 ( .A1(n11789), .A2(n11787), .ZN(n15978) );
  OAI21_X1 U15169 ( .B1(n15973), .B2(n15978), .A(n20250), .ZN(n15959) );
  INV_X1 U15170 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n11788) );
  NAND2_X1 U15171 ( .A1(n11789), .A2(n11788), .ZN(n11790) );
  NAND2_X1 U15172 ( .A1(n11791), .A2(n11790), .ZN(n16531) );
  NAND2_X1 U15173 ( .A1(n15959), .A2(n16531), .ZN(n15944) );
  INV_X1 U15174 ( .A(n15944), .ZN(n15941) );
  NAND3_X1 U15175 ( .A1(n10667), .A2(n11793), .A3(n11792), .ZN(P2_U2825) );
  INV_X1 U15176 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n17948) );
  NAND2_X1 U15177 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n19097) );
  NAND2_X1 U15178 ( .A1(n19098), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n19071) );
  INV_X1 U15179 ( .A(n19071), .ZN(n11794) );
  NAND2_X1 U15180 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n19072) );
  NAND2_X1 U15181 ( .A1(n19053), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n11801) );
  NAND2_X1 U15182 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n19027) );
  NAND2_X1 U15183 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n18998) );
  NAND2_X1 U15184 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n18953) );
  NAND2_X1 U15185 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n18925) );
  XNOR2_X1 U15186 ( .A(n17948), .B(n11802), .ZN(n17947) );
  NAND2_X1 U15187 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n11795), .ZN(
        n17339) );
  NOR2_X1 U15188 ( .A1(n17339), .A2(n10470), .ZN(n11798) );
  INV_X1 U15189 ( .A(n11798), .ZN(n11797) );
  OR2_X1 U15190 ( .A1(n11797), .A2(n18925), .ZN(n17174) );
  AOI21_X1 U15191 ( .B1(n17174), .B2(n10471), .A(n11802), .ZN(n17955) );
  INV_X1 U15192 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n18943) );
  NOR2_X1 U15193 ( .A1(n11797), .A2(n18943), .ZN(n11796) );
  OAI21_X1 U15194 ( .B1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n11796), .A(
        n17174), .ZN(n18928) );
  INV_X1 U15195 ( .A(n18928), .ZN(n17966) );
  AOI21_X1 U15196 ( .B1(n11797), .B2(n18943), .A(n11796), .ZN(n18937) );
  AOI21_X1 U15197 ( .B1(n17339), .B2(n10470), .A(n11798), .ZN(n17984) );
  INV_X1 U15198 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n18966) );
  NOR3_X1 U15199 ( .A1(n18301), .A2(n11799), .A3(n18966), .ZN(n11807) );
  OAI21_X1 U15200 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n11807), .A(
        n17339), .ZN(n18955) );
  INV_X1 U15201 ( .A(n18955), .ZN(n17995) );
  NOR2_X1 U15202 ( .A1(n18301), .A2(n9789), .ZN(n18994) );
  NAND2_X1 U15203 ( .A1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n18994), .ZN(
        n11804) );
  NOR2_X1 U15204 ( .A1(n18998), .A2(n11804), .ZN(n18951) );
  OAI22_X1 U15205 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n18951), .B1(
        n18301), .B2(n11799), .ZN(n18984) );
  INV_X1 U15206 ( .A(n18984), .ZN(n18014) );
  INV_X1 U15207 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n18026) );
  INV_X1 U15208 ( .A(n11804), .ZN(n11805) );
  NAND2_X1 U15209 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n11805), .ZN(
        n11800) );
  AOI21_X1 U15210 ( .B1(n18026), .B2(n11800), .A(n18951), .ZN(n18997) );
  INV_X1 U15211 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n19016) );
  INV_X1 U15212 ( .A(n18994), .ZN(n18055) );
  AOI21_X1 U15213 ( .B1(n19016), .B2(n18055), .A(n11805), .ZN(n19018) );
  INV_X1 U15214 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n19041) );
  NOR2_X1 U15215 ( .A1(n18301), .A2(n11801), .ZN(n19025) );
  INV_X1 U15216 ( .A(n19096), .ZN(n18171) );
  NAND2_X1 U15217 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n19069), .ZN(
        n18108) );
  NAND2_X1 U15218 ( .A1(n11802), .A2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11803) );
  XNOR2_X2 U15219 ( .A(n11803), .B(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n17277) );
  INV_X1 U15220 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n19007) );
  AOI22_X1 U15221 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n11805), .B1(
        n11804), .B2(n19007), .ZN(n19004) );
  INV_X1 U15222 ( .A(n18006), .ZN(n11810) );
  OR2_X1 U15223 ( .A1(n18301), .A2(n11799), .ZN(n11808) );
  AOI21_X1 U15224 ( .B1(n18966), .B2(n11808), .A(n11807), .ZN(n18963) );
  NAND2_X1 U15225 ( .A1(n11810), .A2(n11809), .ZN(n18004) );
  NOR2_X1 U15226 ( .A1(n18937), .A2(n17974), .ZN(n17973) );
  NOR2_X1 U15227 ( .A1(n17973), .A2(n18227), .ZN(n17965) );
  NOR2_X1 U15228 ( .A1(n17966), .A2(n17965), .ZN(n17964) );
  NOR2_X1 U15229 ( .A1(n17964), .A2(n18227), .ZN(n17954) );
  NOR2_X1 U15230 ( .A1(n17953), .A2(n18227), .ZN(n17946) );
  NAND3_X1 U15231 ( .A1(n20175), .A2(n20187), .A3(n17926), .ZN(n20053) );
  NOR2_X1 U15232 ( .A1(n18227), .A2(n20051), .ZN(n18289) );
  INV_X1 U15233 ( .A(n18289), .ZN(n11811) );
  NOR3_X1 U15234 ( .A1(n17947), .A2(n17946), .A3(n11811), .ZN(n12015) );
  AOI22_X1 U15235 ( .A1(n18390), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n18403), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11818) );
  INV_X2 U15236 ( .A(n18551), .ZN(n18626) );
  AND2_X2 U15237 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n18256) );
  NAND2_X2 U15238 ( .A1(n18256), .A2(n11813), .ZN(n18615) );
  AOI22_X1 U15239 ( .A1(n18626), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n14232), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11817) );
  OR2_X1 U15240 ( .A1(n18599), .A2(n18612), .ZN(n11816) );
  NAND2_X1 U15241 ( .A1(n9726), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n11815) );
  NAND2_X1 U15242 ( .A1(n18591), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11821) );
  NAND2_X1 U15243 ( .A1(n18586), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11820) );
  OAI211_X1 U15244 ( .C1(n17478), .C2(n11880), .A(n11821), .B(n11820), .ZN(
        n11822) );
  INV_X1 U15245 ( .A(n11822), .ZN(n11837) );
  NAND2_X1 U15246 ( .A1(n18585), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11828) );
  NAND2_X1 U15247 ( .A1(n9724), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11827) );
  NAND2_X1 U15248 ( .A1(n17547), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11826) );
  AND2_X2 U15249 ( .A1(n14031), .A2(n11824), .ZN(n11911) );
  NAND2_X1 U15250 ( .A1(n11911), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11825) );
  NAND4_X1 U15251 ( .A1(n11828), .A2(n11827), .A3(n11826), .A4(n11825), .ZN(
        n11835) );
  INV_X1 U15252 ( .A(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n18609) );
  INV_X4 U15253 ( .A(n18466), .ZN(n18620) );
  NAND2_X1 U15254 ( .A1(n18620), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11833) );
  INV_X2 U15255 ( .A(n9786), .ZN(n18489) );
  NAND2_X1 U15256 ( .A1(n18489), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11832) );
  OAI211_X1 U15257 ( .C1(n17550), .C2(n18609), .A(n11833), .B(n11832), .ZN(
        n11834) );
  AOI22_X1 U15258 ( .A1(n18597), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11911), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11845) );
  INV_X1 U15259 ( .A(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11839) );
  OAI22_X1 U15260 ( .A1(n18613), .A2(n11839), .B1(n18615), .B2(n22079), .ZN(
        n11840) );
  INV_X1 U15261 ( .A(n11840), .ZN(n11844) );
  INV_X1 U15262 ( .A(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11841) );
  OR2_X1 U15263 ( .A1(n18599), .A2(n11841), .ZN(n11843) );
  NAND2_X1 U15264 ( .A1(n9726), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n11842) );
  INV_X1 U15265 ( .A(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11848) );
  NAND2_X1 U15266 ( .A1(n18591), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n11847) );
  NAND2_X1 U15267 ( .A1(n18627), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n11846) );
  OAI211_X1 U15268 ( .C1(n17550), .C2(n11848), .A(n11847), .B(n11846), .ZN(
        n11849) );
  INV_X1 U15269 ( .A(n11849), .ZN(n11859) );
  INV_X1 U15270 ( .A(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n19777) );
  NAND2_X1 U15271 ( .A1(n18620), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n11851) );
  NAND2_X1 U15272 ( .A1(n18586), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n11850) );
  OAI211_X1 U15273 ( .C1(n9786), .C2(n19777), .A(n11851), .B(n11850), .ZN(
        n11852) );
  INV_X1 U15274 ( .A(n11852), .ZN(n11858) );
  NAND2_X1 U15275 ( .A1(n18390), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n11856) );
  NAND2_X1 U15276 ( .A1(n17547), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n11855) );
  NAND2_X1 U15277 ( .A1(n9724), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n11854) );
  NAND2_X1 U15278 ( .A1(n17561), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n11853) );
  AOI22_X1 U15279 ( .A1(n11911), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n14232), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11865) );
  AOI22_X1 U15280 ( .A1(n18390), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17561), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11864) );
  INV_X1 U15281 ( .A(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n18575) );
  OR2_X1 U15282 ( .A1(n18599), .A2(n18575), .ZN(n11863) );
  NAND2_X1 U15283 ( .A1(n9726), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n11862) );
  INV_X1 U15284 ( .A(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17176) );
  NAND2_X1 U15285 ( .A1(n18591), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n11867) );
  NAND2_X1 U15286 ( .A1(n18586), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n11866) );
  OAI211_X1 U15287 ( .C1(n10660), .C2(n17176), .A(n11867), .B(n11866), .ZN(
        n11868) );
  INV_X1 U15288 ( .A(n11868), .ZN(n11878) );
  NAND2_X1 U15289 ( .A1(n18585), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n11872) );
  NAND2_X1 U15290 ( .A1(n9724), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n11871) );
  NAND2_X1 U15291 ( .A1(n17547), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n11870) );
  NAND2_X1 U15292 ( .A1(n18597), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n11869) );
  NAND4_X1 U15293 ( .A1(n11872), .A2(n11871), .A3(n11870), .A4(n11869), .ZN(
        n11876) );
  INV_X1 U15294 ( .A(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n18431) );
  NAND2_X1 U15295 ( .A1(n18620), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n11874) );
  NAND2_X1 U15296 ( .A1(n18489), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n11873) );
  OAI211_X1 U15297 ( .C1(n17550), .C2(n18431), .A(n11874), .B(n11873), .ZN(
        n11875) );
  NOR2_X1 U15298 ( .A1(n11876), .A2(n11875), .ZN(n11877) );
  INV_X1 U15299 ( .A(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n18394) );
  INV_X1 U15300 ( .A(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17542) );
  OAI22_X1 U15301 ( .A1(n18613), .A2(n18394), .B1(n18616), .B2(n17542), .ZN(
        n11882) );
  OAI22_X1 U15302 ( .A1(n18393), .A2(n18615), .B1(n11880), .B2(n17543), .ZN(
        n11881) );
  NOR2_X1 U15303 ( .A1(n11882), .A2(n11881), .ZN(n11889) );
  AOI22_X1 U15304 ( .A1(n18586), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11911), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11888) );
  INV_X1 U15305 ( .A(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n18395) );
  NAND2_X1 U15306 ( .A1(n18620), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n11884) );
  NAND2_X1 U15307 ( .A1(n18489), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n11883) );
  OAI211_X1 U15308 ( .C1(n17550), .C2(n18395), .A(n11884), .B(n11883), .ZN(
        n11885) );
  INV_X1 U15309 ( .A(n11885), .ZN(n11887) );
  NAND2_X1 U15310 ( .A1(n18591), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n11886) );
  NAND4_X1 U15311 ( .A1(n11889), .A2(n11888), .A3(n11887), .A4(n11886), .ZN(
        n11894) );
  AOI22_X1 U15312 ( .A1(n18628), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9726), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11892) );
  AOI22_X1 U15313 ( .A1(n18597), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n18390), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11891) );
  AOI22_X1 U15314 ( .A1(n9724), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n18403), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11890) );
  NAND3_X1 U15315 ( .A1(n11892), .A2(n11891), .A3(n11890), .ZN(n11893) );
  AOI22_X1 U15316 ( .A1(n9724), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n18620), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11906) );
  INV_X2 U15317 ( .A(n9786), .ZN(n18619) );
  AOI22_X1 U15318 ( .A1(n18626), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n18619), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11895) );
  OAI21_X1 U15319 ( .B1(n17550), .B2(n18447), .A(n11895), .ZN(n11896) );
  INV_X1 U15320 ( .A(n11896), .ZN(n11905) );
  INV_X1 U15321 ( .A(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11897) );
  OAI22_X1 U15322 ( .A1(n10660), .A2(n11897), .B1(n18615), .B2(n18448), .ZN(
        n11898) );
  INV_X1 U15323 ( .A(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13992) );
  OAI22_X1 U15324 ( .A1(n18525), .A2(n13992), .B1(n11880), .B2(n13982), .ZN(
        n11899) );
  INV_X1 U15325 ( .A(n11899), .ZN(n11904) );
  AOI22_X1 U15326 ( .A1(n11911), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17547), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11903) );
  INV_X1 U15327 ( .A(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11900) );
  INV_X1 U15328 ( .A(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n18449) );
  OAI22_X1 U15329 ( .A1(n18611), .A2(n11900), .B1(n18613), .B2(n18449), .ZN(
        n11901) );
  AOI21_X1 U15330 ( .B1(n18413), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A(
        n11901), .ZN(n11902) );
  AOI22_X1 U15331 ( .A1(n18390), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n18403), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11910) );
  AOI22_X1 U15332 ( .A1(n18626), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n14232), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11909) );
  INV_X1 U15333 ( .A(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n18411) );
  OR2_X1 U15334 ( .A1(n18599), .A2(n18411), .ZN(n11908) );
  NAND2_X1 U15335 ( .A1(n9726), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n11907) );
  INV_X1 U15336 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n18650) );
  NAND2_X1 U15337 ( .A1(n18591), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n11913) );
  NAND2_X1 U15338 ( .A1(n18586), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n11912) );
  OAI211_X1 U15339 ( .C1(n11861), .C2(n18650), .A(n11913), .B(n11912), .ZN(
        n11914) );
  INV_X1 U15340 ( .A(n11914), .ZN(n11924) );
  NAND2_X1 U15341 ( .A1(n18585), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n11918) );
  NAND2_X1 U15342 ( .A1(n9724), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n11917) );
  NAND2_X1 U15343 ( .A1(n17547), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n11916) );
  NAND2_X1 U15344 ( .A1(n17561), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n11915) );
  NAND4_X1 U15345 ( .A1(n11918), .A2(n11917), .A3(n11916), .A4(n11915), .ZN(
        n11922) );
  INV_X1 U15346 ( .A(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n18418) );
  NAND2_X1 U15347 ( .A1(n18620), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n11920) );
  NAND2_X1 U15348 ( .A1(n18489), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n11919) );
  OAI211_X1 U15349 ( .C1(n17550), .C2(n18418), .A(n11920), .B(n11919), .ZN(
        n11921) );
  NOR2_X1 U15350 ( .A1(n11922), .A2(n11921), .ZN(n11923) );
  AOI22_X1 U15351 ( .A1(n18390), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n18627), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11929) );
  AOI22_X1 U15352 ( .A1(n18597), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n14232), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11928) );
  OR2_X1 U15353 ( .A1(n18599), .A2(n18527), .ZN(n11927) );
  NAND2_X1 U15354 ( .A1(n9726), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n11926) );
  NAND2_X1 U15355 ( .A1(n18591), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n11931) );
  NAND2_X1 U15356 ( .A1(n18586), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n11930) );
  OAI211_X1 U15357 ( .C1(n11861), .C2(n18644), .A(n11931), .B(n11930), .ZN(
        n11932) );
  INV_X1 U15358 ( .A(n11932), .ZN(n11943) );
  NAND2_X1 U15359 ( .A1(n18585), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n11936) );
  NAND2_X1 U15360 ( .A1(n9724), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n11935) );
  NAND2_X1 U15361 ( .A1(n17547), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n11934) );
  NAND2_X1 U15362 ( .A1(n17561), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n11933) );
  NAND4_X1 U15363 ( .A1(n11936), .A2(n11935), .A3(n11934), .A4(n11933), .ZN(
        n11941) );
  INV_X1 U15364 ( .A(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n18369) );
  NAND2_X1 U15365 ( .A1(n18620), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n11939) );
  NAND2_X1 U15366 ( .A1(n18489), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n11938) );
  OAI211_X1 U15367 ( .C1(n17550), .C2(n18369), .A(n11939), .B(n11938), .ZN(
        n11940) );
  NOR2_X1 U15368 ( .A1(n11941), .A2(n11940), .ZN(n11942) );
  AND3_X2 U15369 ( .A1(n11944), .A2(n11943), .A3(n11942), .ZN(n19555) );
  NAND2_X1 U15370 ( .A1(n18585), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11948) );
  NAND2_X1 U15371 ( .A1(n17547), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11947) );
  NAND2_X1 U15372 ( .A1(n9724), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11946) );
  NAND2_X1 U15373 ( .A1(n11911), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11945) );
  NAND4_X1 U15374 ( .A1(n11948), .A2(n11947), .A3(n11946), .A4(n11945), .ZN(
        n11953) );
  NAND2_X1 U15375 ( .A1(n18620), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11950) );
  NAND2_X1 U15376 ( .A1(n18489), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11949) );
  OAI211_X1 U15377 ( .C1(n17550), .C2(n11951), .A(n11950), .B(n11949), .ZN(
        n11952) );
  NAND2_X1 U15378 ( .A1(n18597), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n11957) );
  NAND2_X1 U15379 ( .A1(n18390), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n11956) );
  NAND2_X1 U15380 ( .A1(n18627), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11955) );
  NAND2_X1 U15381 ( .A1(n17561), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11954) );
  NAND2_X1 U15382 ( .A1(n18591), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n11959) );
  NAND2_X1 U15383 ( .A1(n18586), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11958) );
  OAI211_X1 U15384 ( .C1(n17507), .C2(n18615), .A(n11959), .B(n11958), .ZN(
        n11960) );
  INV_X1 U15385 ( .A(n11960), .ZN(n11962) );
  NAND4_X4 U15386 ( .A1(n11964), .A2(n11963), .A3(n11962), .A4(n11961), .ZN(
        n20171) );
  NAND2_X1 U15387 ( .A1(n19532), .A2(n20171), .ZN(n14175) );
  NOR2_X1 U15388 ( .A1(n11965), .A2(n14179), .ZN(n19976) );
  NOR2_X1 U15389 ( .A1(n19555), .A2(n18680), .ZN(n14011) );
  NAND2_X1 U15390 ( .A1(n19976), .A2(n14011), .ZN(n13968) );
  INV_X1 U15391 ( .A(n13968), .ZN(n11967) );
  NOR2_X1 U15392 ( .A1(n20171), .A2(n11975), .ZN(n11966) );
  NAND2_X1 U15393 ( .A1(n18680), .A2(n19539), .ZN(n14189) );
  NAND2_X1 U15394 ( .A1(n19535), .A2(n18818), .ZN(n14174) );
  AOI21_X1 U15395 ( .B1(n18765), .B2(n14110), .A(n14174), .ZN(n14018) );
  AOI21_X1 U15396 ( .B1(n14189), .B2(n11968), .A(n14018), .ZN(n11980) );
  INV_X1 U15397 ( .A(n11974), .ZN(n11973) );
  NAND2_X1 U15398 ( .A1(n14175), .A2(n19539), .ZN(n14014) );
  INV_X1 U15399 ( .A(n14014), .ZN(n11972) );
  OAI21_X1 U15400 ( .B1(n14179), .B2(n18818), .A(n14110), .ZN(n11969) );
  OAI21_X1 U15401 ( .B1(n11973), .B2(n11970), .A(n11969), .ZN(n11971) );
  OAI21_X1 U15402 ( .B1(n11973), .B2(n11972), .A(n11971), .ZN(n11979) );
  AOI21_X1 U15403 ( .B1(n18765), .B2(n11974), .A(n19547), .ZN(n11977) );
  AND2_X1 U15404 ( .A1(n19543), .A2(n11975), .ZN(n11976) );
  OAI21_X1 U15405 ( .B1(n19543), .B2(n11980), .A(n14016), .ZN(n14027) );
  INV_X1 U15406 ( .A(n13970), .ZN(n11983) );
  MUX2_X1 U15407 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n20002), .S(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n13971) );
  NOR2_X1 U15408 ( .A1(n11983), .A2(n13971), .ZN(n11984) );
  OR2_X1 U15409 ( .A1(n11989), .A2(n11990), .ZN(n11985) );
  OAI22_X1 U15410 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n20022), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n11986), .ZN(n11993) );
  NOR2_X1 U15411 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n20022), .ZN(
        n11987) );
  NAND2_X1 U15412 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n11986), .ZN(
        n11992) );
  AOI22_X1 U15413 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n11993), .B1(
        n11987), .B2(n11992), .ZN(n13973) );
  OAI21_X1 U15414 ( .B1(n11990), .B2(n11989), .A(n13973), .ZN(n11988) );
  XNOR2_X1 U15415 ( .A(n13971), .B(n13970), .ZN(n11991) );
  NAND2_X1 U15416 ( .A1(n14178), .A2(n11991), .ZN(n11996) );
  OAI22_X1 U15417 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n18236), .B1(
        n11994), .B2(n11993), .ZN(n13974) );
  INV_X1 U15418 ( .A(n13974), .ZN(n11995) );
  NAND2_X1 U15419 ( .A1(n20171), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n12003) );
  AOI211_X4 U15420 ( .C1(n17926), .C2(n20181), .A(n12005), .B(n12003), .ZN(
        n18259) );
  INV_X1 U15421 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n18649) );
  NAND2_X1 U15422 ( .A1(n18267), .A2(n18649), .ZN(n18258) );
  NAND2_X1 U15423 ( .A1(n18235), .A2(n18641), .ZN(n18232) );
  NOR2_X1 U15424 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n18232), .ZN(n18215) );
  NAND2_X1 U15425 ( .A1(n18215), .A2(n18633), .ZN(n18212) );
  NAND2_X1 U15426 ( .A1(n18183), .A2(n18191), .ZN(n18166) );
  NAND2_X1 U15427 ( .A1(n18165), .A2(n18164), .ZN(n18156) );
  INV_X1 U15428 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n18131) );
  NAND2_X1 U15429 ( .A1(n18140), .A2(n18131), .ZN(n18130) );
  INV_X1 U15430 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n18522) );
  NAND2_X1 U15431 ( .A1(n18119), .A2(n18522), .ZN(n18106) );
  INV_X1 U15432 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n18083) );
  NAND2_X1 U15433 ( .A1(n18092), .A2(n18083), .ZN(n18081) );
  INV_X1 U15434 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n18064) );
  NAND2_X1 U15435 ( .A1(n18072), .A2(n18064), .ZN(n18063) );
  NAND2_X1 U15436 ( .A1(n18046), .A2(n18389), .ZN(n18039) );
  NAND2_X1 U15437 ( .A1(n18025), .A2(n22099), .ZN(n18018) );
  NAND2_X1 U15438 ( .A1(n18003), .A2(n18002), .ZN(n17998) );
  INV_X1 U15439 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n18346) );
  NAND2_X1 U15440 ( .A1(n17985), .A2(n18346), .ZN(n17977) );
  INV_X1 U15441 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n18338) );
  NAND2_X1 U15442 ( .A1(n17963), .A2(n18338), .ZN(n17945) );
  NOR2_X1 U15443 ( .A1(n18295), .A2(n17945), .ZN(n17951) );
  INV_X1 U15444 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n18304) );
  AND2_X1 U15445 ( .A1(n17951), .A2(n18304), .ZN(n12014) );
  INV_X1 U15446 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n20125) );
  NAND2_X1 U15447 ( .A1(P3_STATE_REG_2__SCAN_IN), .A2(n20073), .ZN(n20059) );
  NAND2_X2 U15448 ( .A1(n20184), .A2(n20066), .ZN(n20116) );
  OAI211_X1 U15449 ( .C1(n20171), .C2(n20170), .A(n20181), .B(n17926), .ZN(
        n20034) );
  INV_X1 U15450 ( .A(n20190), .ZN(n20177) );
  NAND2_X1 U15451 ( .A1(n20187), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n20046) );
  INV_X1 U15452 ( .A(n20046), .ZN(n19915) );
  NAND2_X1 U15453 ( .A1(n20048), .A2(n19915), .ZN(n20041) );
  NAND2_X1 U15454 ( .A1(n18291), .A2(n18242), .ZN(n18097) );
  NAND2_X1 U15455 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .ZN(n12000) );
  INV_X1 U15456 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n20117) );
  INV_X1 U15457 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n20114) );
  NOR2_X1 U15458 ( .A1(n20117), .A2(n20114), .ZN(n11999) );
  INV_X1 U15459 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n20105) );
  INV_X1 U15460 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n20102) );
  NAND2_X1 U15461 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(P3_REIP_REG_15__SCAN_IN), 
        .ZN(n18084) );
  NOR2_X1 U15462 ( .A1(n20102), .A2(n18084), .ZN(n18058) );
  NAND2_X1 U15463 ( .A1(P3_REIP_REG_18__SCAN_IN), .A2(n18058), .ZN(n18059) );
  NOR2_X1 U15464 ( .A1(n20105), .A2(n18059), .ZN(n18043) );
  NAND2_X1 U15465 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n18043), .ZN(n18022) );
  NAND2_X1 U15466 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(P3_REIP_REG_21__SCAN_IN), 
        .ZN(n18030) );
  OR3_X1 U15467 ( .A1(n20113), .A2(n18022), .A3(n18030), .ZN(n11998) );
  INV_X1 U15468 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n20095) );
  INV_X1 U15469 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n20091) );
  INV_X1 U15470 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n20077) );
  NAND2_X1 U15471 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .ZN(n18271) );
  NOR2_X1 U15472 ( .A1(n20077), .A2(n18271), .ZN(n18243) );
  NAND3_X1 U15473 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(P3_REIP_REG_4__SCAN_IN), 
        .A3(n18243), .ZN(n18174) );
  NAND3_X1 U15474 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(P3_REIP_REG_7__SCAN_IN), 
        .A3(P3_REIP_REG_6__SCAN_IN), .ZN(n18173) );
  NOR2_X1 U15475 ( .A1(n22085), .A2(n18173), .ZN(n18169) );
  NAND2_X1 U15476 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(n18169), .ZN(n18152) );
  NOR3_X1 U15477 ( .A1(n20091), .A2(n18174), .A3(n18152), .ZN(n18143) );
  NAND2_X1 U15478 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n18143), .ZN(n18128) );
  NOR2_X1 U15479 ( .A1(n20095), .A2(n18128), .ZN(n11997) );
  NAND3_X1 U15480 ( .A1(n11997), .A2(P3_REIP_REG_14__SCAN_IN), .A3(n18242), 
        .ZN(n18096) );
  OAI21_X1 U15481 ( .B1(n11998), .B2(n18096), .A(n18097), .ZN(n18015) );
  OAI221_X1 U15482 ( .B1(n18291), .B2(P3_REIP_REG_26__SCAN_IN), .C1(n18291), 
        .C2(n11999), .A(n18015), .ZN(n17981) );
  AOI221_X1 U15483 ( .B1(n20125), .B2(n18097), .C1(n12000), .C2(n18097), .A(
        n17981), .ZN(n17961) );
  INV_X1 U15484 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n22146) );
  NAND2_X1 U15485 ( .A1(n18272), .A2(n11997), .ZN(n18118) );
  NAND2_X1 U15486 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(n17988), .ZN(n17980) );
  NOR2_X1 U15487 ( .A1(n17980), .A2(n12000), .ZN(n17959) );
  NAND2_X1 U15488 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n17959), .ZN(n12006) );
  NOR2_X1 U15489 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n12006), .ZN(n17949) );
  INV_X1 U15490 ( .A(n17949), .ZN(n12001) );
  INV_X1 U15491 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n20127) );
  AOI21_X1 U15492 ( .B1(n17961), .B2(n12001), .A(n20127), .ZN(n12002) );
  INV_X1 U15493 ( .A(n12002), .ZN(n12012) );
  NAND2_X1 U15494 ( .A1(n20034), .A2(n12003), .ZN(n12004) );
  INV_X1 U15495 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n20129) );
  NOR3_X1 U15496 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n20129), .A3(n12006), 
        .ZN(n12007) );
  AOI21_X1 U15497 ( .B1(n9707), .B2(P3_EBX_REG_31__SCAN_IN), .A(n12007), .ZN(
        n12008) );
  INV_X1 U15498 ( .A(n12008), .ZN(n12010) );
  INV_X1 U15499 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n17332) );
  NOR2_X1 U15500 ( .A1(n12010), .A2(n12009), .ZN(n12011) );
  NAND2_X1 U15501 ( .A1(n12012), .A2(n12011), .ZN(n12013) );
  AOI21_X1 U15502 ( .B1(n12018), .B2(n11452), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n13499) );
  NOR2_X1 U15503 ( .A1(n10680), .A2(n13499), .ZN(n12019) );
  OR2_X1 U15504 ( .A1(n13623), .A2(n20400), .ZN(n12024) );
  NAND2_X1 U15505 ( .A1(n12020), .A2(n9731), .ZN(n12021) );
  NAND2_X1 U15506 ( .A1(n12021), .A2(n10908), .ZN(n12023) );
  NAND2_X1 U15507 ( .A1(n12022), .A2(n9736), .ZN(n14141) );
  MUX2_X1 U15508 ( .A(n12024), .B(n12023), .S(n14141), .Z(n12046) );
  NAND2_X1 U15509 ( .A1(n12025), .A2(n20400), .ZN(n12026) );
  NAND2_X1 U15510 ( .A1(n13614), .A2(n12026), .ZN(n12035) );
  AND2_X1 U15511 ( .A1(n12028), .A2(n12027), .ZN(n12034) );
  OAI21_X1 U15512 ( .B1(n12030), .B2(n9722), .A(n12029), .ZN(n12055) );
  NAND2_X1 U15513 ( .A1(n10908), .A2(n9735), .ZN(n12051) );
  NAND2_X1 U15514 ( .A1(n12051), .A2(n9731), .ZN(n12031) );
  NAND2_X1 U15515 ( .A1(n12031), .A2(n13819), .ZN(n12032) );
  NAND2_X1 U15516 ( .A1(n12032), .A2(n20400), .ZN(n12033) );
  NAND4_X1 U15517 ( .A1(n12035), .A2(n12034), .A3(n12055), .A4(n12033), .ZN(
        n12050) );
  NOR2_X1 U15518 ( .A1(n12036), .A2(n13623), .ZN(n12037) );
  NOR2_X1 U15519 ( .A1(n12050), .A2(n12037), .ZN(n14136) );
  INV_X1 U15520 ( .A(n10905), .ZN(n12038) );
  NAND3_X1 U15521 ( .A1(n12039), .A2(n12038), .A3(n9736), .ZN(n12044) );
  MUX2_X1 U15522 ( .A(n12041), .B(n12040), .S(n9735), .Z(n12042) );
  NAND3_X1 U15523 ( .A1(n12042), .A2(n17778), .A3(n21133), .ZN(n12043) );
  NAND2_X1 U15524 ( .A1(n12046), .A2(n12045), .ZN(n12047) );
  AND2_X1 U15525 ( .A1(n12048), .A2(n9735), .ZN(n12049) );
  INV_X1 U15526 ( .A(n12050), .ZN(n12053) );
  INV_X1 U15527 ( .A(n12051), .ZN(n12052) );
  NAND2_X1 U15528 ( .A1(n12053), .A2(n12052), .ZN(n14121) );
  INV_X1 U15529 ( .A(n14121), .ZN(n17775) );
  NAND2_X1 U15530 ( .A1(n12054), .A2(n9736), .ZN(n17126) );
  NAND2_X1 U15531 ( .A1(n17126), .A2(n12055), .ZN(n12057) );
  NAND2_X1 U15532 ( .A1(n12057), .A2(n12056), .ZN(n12067) );
  OAI22_X1 U15533 ( .A1(n11257), .A2(n20415), .B1(n9731), .B2(n20400), .ZN(
        n12058) );
  INV_X1 U15534 ( .A(n12058), .ZN(n12059) );
  AND2_X1 U15535 ( .A1(n12060), .A2(n12059), .ZN(n12066) );
  AND2_X1 U15536 ( .A1(n12061), .A2(n12062), .ZN(n12064) );
  INV_X1 U15537 ( .A(n11257), .ZN(n13630) );
  OAI21_X1 U15538 ( .B1(n12064), .B2(n13630), .A(n12063), .ZN(n12065) );
  AND3_X1 U15539 ( .A1(n12067), .A2(n12066), .A3(n12065), .ZN(n14124) );
  NAND2_X1 U15540 ( .A1(n14124), .A2(n13776), .ZN(n12068) );
  NAND2_X1 U15541 ( .A1(n12092), .A2(n12068), .ZN(n14756) );
  NAND3_X1 U15542 ( .A1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n13516) );
  NAND2_X1 U15543 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n17110) );
  INV_X1 U15544 ( .A(n17110), .ZN(n14696) );
  INV_X1 U15545 ( .A(n12092), .ZN(n12069) );
  NAND2_X1 U15546 ( .A1(n12069), .A2(n20217), .ZN(n17103) );
  OAI21_X1 U15547 ( .B1(n14756), .B2(n14696), .A(n17103), .ZN(n14709) );
  NOR2_X1 U15548 ( .A1(n14756), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n14697) );
  OR2_X1 U15549 ( .A1(n14709), .A2(n14697), .ZN(n17068) );
  INV_X1 U15550 ( .A(n17068), .ZN(n17021) );
  NAND2_X1 U15551 ( .A1(n17021), .A2(n17071), .ZN(n12074) );
  INV_X1 U15552 ( .A(n12074), .ZN(n12076) );
  NOR2_X1 U15553 ( .A1(n16788), .A2(n12070), .ZN(n12083) );
  NOR2_X1 U15554 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n14696), .ZN(
        n17069) );
  NAND3_X1 U15555 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n17026) );
  NOR2_X1 U15556 ( .A1(n17069), .A2(n17026), .ZN(n17016) );
  NAND4_X1 U15557 ( .A1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A4(n17016), .ZN(n17001) );
  AND2_X1 U15558 ( .A1(n17111), .A2(n17001), .ZN(n12071) );
  NOR2_X1 U15559 ( .A1(n12071), .A2(n17068), .ZN(n17007) );
  NAND2_X1 U15560 ( .A1(n17111), .A2(n17006), .ZN(n12072) );
  AOI21_X1 U15561 ( .B1(n17111), .B2(n16849), .A(n16848), .ZN(n12073) );
  NAND2_X1 U15562 ( .A1(n16993), .A2(n12073), .ZN(n16851) );
  NAND2_X1 U15563 ( .A1(n16851), .A2(n12074), .ZN(n16842) );
  INV_X1 U15564 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n16841) );
  OR2_X1 U15565 ( .A1(n22170), .A2(n16841), .ZN(n16824) );
  NAND2_X1 U15566 ( .A1(n12074), .A2(n16824), .ZN(n12075) );
  AND2_X1 U15567 ( .A1(n16842), .A2(n12075), .ZN(n16814) );
  OAI21_X1 U15568 ( .B1(n12076), .B2(n12083), .A(n16814), .ZN(n14727) );
  AOI21_X1 U15569 ( .B1(n17111), .B2(n13516), .A(n14727), .ZN(n13515) );
  INV_X1 U15570 ( .A(n13515), .ZN(n12085) );
  INV_X1 U15571 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n21078) );
  NOR2_X1 U15572 ( .A1(n16730), .A2(n21078), .ZN(n14737) );
  NOR2_X1 U15573 ( .A1(n12077), .A2(n17110), .ZN(n14703) );
  INV_X1 U15574 ( .A(n14703), .ZN(n12078) );
  NAND2_X1 U15575 ( .A1(n14751), .A2(n12078), .ZN(n12079) );
  NAND2_X1 U15576 ( .A1(n17111), .A2(n12079), .ZN(n17023) );
  INV_X1 U15577 ( .A(n17001), .ZN(n12080) );
  NAND2_X1 U15578 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n12080), .ZN(
        n12081) );
  INV_X1 U15579 ( .A(n16849), .ZN(n12082) );
  NAND3_X1 U15580 ( .A1(n16989), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        n12082), .ZN(n16823) );
  NOR2_X1 U15581 ( .A1(n16823), .A2(n16824), .ZN(n16789) );
  NAND2_X1 U15582 ( .A1(n16789), .A2(n12083), .ZN(n16764) );
  NOR3_X1 U15583 ( .A1(n16764), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n13516), .ZN(n12084) );
  AOI211_X1 U15584 ( .C1(n12085), .C2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n14737), .B(n12084), .ZN(n12086) );
  OAI21_X1 U15585 ( .B1(n14741), .B2(n17745), .A(n12086), .ZN(n12087) );
  INV_X1 U15586 ( .A(n17127), .ZN(n12090) );
  INV_X1 U15587 ( .A(n12088), .ZN(n12089) );
  INV_X1 U15588 ( .A(n17776), .ZN(n14122) );
  OAI21_X1 U15589 ( .B1(n9735), .B2(n17779), .A(n14122), .ZN(n12091) );
  OAI211_X1 U15590 ( .C1(n14745), .C2(n17101), .A(n12094), .B(n12093), .ZN(
        P2_U3016) );
  INV_X1 U15591 ( .A(n12098), .ZN(n16676) );
  INV_X1 U15592 ( .A(n16655), .ZN(n12099) );
  INV_X1 U15593 ( .A(n16612), .ZN(n12101) );
  INV_X1 U15594 ( .A(n16615), .ZN(n12102) );
  INV_X1 U15595 ( .A(n16893), .ZN(n16865) );
  OR2_X1 U15596 ( .A1(n12105), .A2(n12106), .ZN(n12107) );
  AND2_X1 U15597 ( .A1(n12104), .A2(n12107), .ZN(n16880) );
  NOR2_X1 U15598 ( .A1(n16730), .A2(n21061), .ZN(n16881) );
  AOI21_X1 U15599 ( .B1(n20356), .B2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n16881), .ZN(n12108) );
  OAI21_X1 U15600 ( .B1(n20368), .B2(n16093), .A(n12108), .ZN(n12109) );
  AND2_X2 U15601 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13870) );
  INV_X1 U15602 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12111) );
  INV_X1 U15603 ( .A(n12261), .ZN(n12186) );
  NAND2_X4 U15604 ( .A1(n13873), .A2(n12697), .ZN(n12342) );
  NAND2_X1 U15605 ( .A1(n12741), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n12119) );
  AND2_X2 U15606 ( .A1(n12697), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12122) );
  NOR2_X4 U15607 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15871) );
  AND2_X4 U15608 ( .A1(n12122), .A2(n15871), .ZN(n12944) );
  NAND2_X1 U15609 ( .A1(n12944), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n12118) );
  INV_X1 U15610 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12114) );
  INV_X1 U15611 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12115) );
  NAND2_X4 U15612 ( .A1(n12129), .A2(n12128), .ZN(n13175) );
  INV_X1 U15613 ( .A(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12116) );
  AND4_X2 U15614 ( .A1(n12120), .A2(n12119), .A3(n12118), .A4(n12117), .ZN(
        n12141) );
  NAND2_X1 U15615 ( .A1(n12390), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n12127) );
  NAND2_X1 U15616 ( .A1(n13125), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n12126) );
  NAND2_X1 U15617 ( .A1(n12391), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n12125) );
  NAND2_X1 U15618 ( .A1(n13075), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n12124) );
  NAND2_X1 U15619 ( .A1(n13279), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n12133) );
  AND2_X2 U15620 ( .A1(n12128), .A2(n15871), .ZN(n12364) );
  NAND2_X1 U15621 ( .A1(n12364), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n12132) );
  NAND2_X1 U15622 ( .A1(n12267), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n12131) );
  NAND2_X1 U15623 ( .A1(n9785), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n12130) );
  AND4_X2 U15624 ( .A1(n12133), .A2(n12132), .A3(n12131), .A4(n12130), .ZN(
        n12139) );
  NAND2_X1 U15625 ( .A1(n12331), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n12136) );
  AND2_X2 U15626 ( .A1(n15871), .A2(n12134), .ZN(n13089) );
  NAND2_X1 U15627 ( .A1(n13089), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n12135) );
  OAI211_X1 U15628 ( .C1(n12259), .C2(n12488), .A(n12136), .B(n12135), .ZN(
        n12137) );
  INV_X1 U15629 ( .A(n12137), .ZN(n12138) );
  NAND4_X4 U15630 ( .A1(n12141), .A2(n12140), .A3(n12139), .A4(n12138), .ZN(
        n12295) );
  AOI22_X1 U15631 ( .A1(n13240), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n13155), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12146) );
  NAND2_X1 U15632 ( .A1(n13079), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n12145) );
  NAND2_X1 U15633 ( .A1(n12343), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n12144) );
  INV_X1 U15634 ( .A(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12142) );
  NAND2_X1 U15635 ( .A1(n12390), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n12150) );
  NAND2_X1 U15636 ( .A1(n12364), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n12149) );
  NAND2_X1 U15637 ( .A1(n12944), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n12148) );
  NAND2_X1 U15638 ( .A1(n13075), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n12147) );
  NAND2_X1 U15639 ( .A1(n12331), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n12154) );
  NAND2_X1 U15640 ( .A1(n12267), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n12153) );
  NAND2_X1 U15641 ( .A1(n9785), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n12152) );
  NAND2_X1 U15642 ( .A1(n13089), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n12151) );
  NAND2_X1 U15643 ( .A1(n13125), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n12156) );
  NAND2_X1 U15644 ( .A1(n12391), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n12155) );
  OAI211_X1 U15645 ( .C1(n12342), .C2(n13284), .A(n12156), .B(n12155), .ZN(
        n12157) );
  INV_X1 U15646 ( .A(n12157), .ZN(n12158) );
  NAND2_X1 U15647 ( .A1(n13279), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n12166) );
  NAND2_X1 U15648 ( .A1(n13079), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n12165) );
  AOI22_X1 U15649 ( .A1(n13240), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12186), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12164) );
  INV_X1 U15650 ( .A(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12162) );
  NAND2_X1 U15651 ( .A1(n12390), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n12170) );
  NAND2_X1 U15652 ( .A1(n12364), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n12169) );
  NAND2_X1 U15653 ( .A1(n12944), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n12168) );
  NAND2_X1 U15654 ( .A1(n13075), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n12167) );
  NAND2_X1 U15655 ( .A1(n12331), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n12174) );
  NAND2_X1 U15656 ( .A1(n12267), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n12173) );
  NAND2_X1 U15657 ( .A1(n9785), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n12172) );
  NAND2_X1 U15658 ( .A1(n13089), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n12171) );
  NAND2_X1 U15659 ( .A1(n13125), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n12176) );
  NAND2_X1 U15660 ( .A1(n12391), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n12175) );
  OAI211_X1 U15661 ( .C1(n12342), .C2(n12470), .A(n12176), .B(n12175), .ZN(
        n12177) );
  INV_X1 U15662 ( .A(n12177), .ZN(n12178) );
  NAND2_X1 U15663 ( .A1(n12331), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n12183) );
  NAND2_X1 U15664 ( .A1(n13089), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n12182) );
  OAI211_X1 U15665 ( .C1(n12259), .C2(n12184), .A(n12183), .B(n12182), .ZN(
        n12185) );
  INV_X1 U15666 ( .A(n12185), .ZN(n12204) );
  AOI22_X1 U15667 ( .A1(n12549), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12186), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12191) );
  INV_X1 U15668 ( .A(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12187) );
  NAND2_X1 U15669 ( .A1(n13075), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n12189) );
  NAND2_X1 U15670 ( .A1(n12944), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n12188) );
  INV_X1 U15671 ( .A(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12192) );
  NAND2_X1 U15672 ( .A1(n13279), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n12195) );
  NAND2_X1 U15673 ( .A1(n12390), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n12194) );
  NAND2_X1 U15674 ( .A1(n12391), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n12193) );
  NAND2_X1 U15675 ( .A1(n12364), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n12200) );
  NAND2_X1 U15676 ( .A1(n13125), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n12199) );
  NAND2_X1 U15677 ( .A1(n12267), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n12198) );
  NAND2_X1 U15678 ( .A1(n9785), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n12197) );
  NOR2_X1 U15679 ( .A1(n12293), .A2(n12307), .ZN(n12237) );
  NAND2_X1 U15680 ( .A1(n12343), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n12211) );
  NAND2_X1 U15681 ( .A1(n13079), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n12210) );
  INV_X1 U15682 ( .A(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12206) );
  INV_X1 U15683 ( .A(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12205) );
  OAI22_X1 U15684 ( .A1(n12381), .A2(n12206), .B1(n12261), .B2(n12205), .ZN(
        n12207) );
  INV_X1 U15685 ( .A(n12207), .ZN(n12209) );
  INV_X1 U15686 ( .A(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12962) );
  OR2_X1 U15687 ( .A1(n12379), .A2(n12962), .ZN(n12208) );
  NAND4_X1 U15688 ( .A1(n12211), .A2(n12210), .A3(n12209), .A4(n12208), .ZN(
        n12217) );
  INV_X1 U15689 ( .A(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12212) );
  NAND2_X1 U15690 ( .A1(n13125), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n12214) );
  NAND2_X1 U15691 ( .A1(n12391), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n12213) );
  NAND3_X1 U15692 ( .A1(n12215), .A2(n12214), .A3(n12213), .ZN(n12216) );
  NOR2_X1 U15693 ( .A1(n12217), .A2(n12216), .ZN(n12223) );
  AOI22_X1 U15694 ( .A1(n12364), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12390), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12221) );
  AOI22_X1 U15695 ( .A1(n12944), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n13075), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12220) );
  AOI22_X1 U15696 ( .A1(n12267), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n9785), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12219) );
  AOI22_X1 U15697 ( .A1(n12331), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n13089), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12218) );
  AND2_X2 U15698 ( .A1(n12223), .A2(n12222), .ZN(n13350) );
  INV_X1 U15699 ( .A(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12983) );
  INV_X1 U15700 ( .A(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13174) );
  INV_X1 U15701 ( .A(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12224) );
  OAI22_X1 U15702 ( .A1(n12381), .A2(n13174), .B1(n12261), .B2(n12224), .ZN(
        n12225) );
  AOI22_X1 U15703 ( .A1(n13125), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12391), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12229) );
  NAND2_X1 U15704 ( .A1(n12741), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n12228) );
  NAND2_X1 U15705 ( .A1(n13079), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n12227) );
  AOI22_X1 U15706 ( .A1(n12267), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n9785), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12234) );
  AOI22_X1 U15707 ( .A1(n12944), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n13075), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12233) );
  AOI22_X1 U15708 ( .A1(n12364), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12390), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12232) );
  AOI22_X1 U15709 ( .A1(n12331), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n13089), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12231) );
  NAND2_X2 U15710 ( .A1(n12236), .A2(n12235), .ZN(n12297) );
  AND3_X2 U15711 ( .A1(n13857), .A2(n12237), .A3(n12301), .ZN(n13324) );
  NAND2_X1 U15712 ( .A1(n13079), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n12239) );
  NAND2_X1 U15713 ( .A1(n12331), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n12238) );
  INV_X1 U15714 ( .A(n12240), .ZN(n12257) );
  NAND2_X1 U15715 ( .A1(n12741), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n12245) );
  OAI22_X1 U15716 ( .A1(n12381), .A2(n13121), .B1(n12261), .B2(n13135), .ZN(
        n12241) );
  INV_X1 U15717 ( .A(n12241), .ZN(n12244) );
  NAND2_X1 U15718 ( .A1(n12944), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n12243) );
  NAND2_X1 U15719 ( .A1(n13125), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n12249) );
  NAND2_X1 U15720 ( .A1(n12390), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n12248) );
  NAND2_X1 U15721 ( .A1(n13089), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n12247) );
  NAND2_X1 U15722 ( .A1(n9785), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12246) );
  NAND2_X1 U15723 ( .A1(n12391), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n12252) );
  NAND2_X1 U15724 ( .A1(n13075), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n12251) );
  NAND2_X1 U15725 ( .A1(n12364), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n12250) );
  INV_X1 U15726 ( .A(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12258) );
  NAND2_X1 U15727 ( .A1(n13079), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n12265) );
  OAI22_X1 U15728 ( .A1(n12381), .A2(n13100), .B1(n12261), .B2(n12260), .ZN(
        n12262) );
  INV_X1 U15729 ( .A(n12262), .ZN(n12263) );
  NAND2_X1 U15730 ( .A1(n12331), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n12271) );
  NAND2_X1 U15731 ( .A1(n12267), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n12270) );
  NAND2_X1 U15732 ( .A1(n9785), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n12269) );
  NAND2_X1 U15733 ( .A1(n13089), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n12268) );
  INV_X1 U15734 ( .A(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12272) );
  OR2_X1 U15735 ( .A1(n12342), .A2(n12272), .ZN(n12275) );
  NAND2_X1 U15736 ( .A1(n13125), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n12274) );
  NAND2_X1 U15737 ( .A1(n12391), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n12273) );
  NAND2_X1 U15738 ( .A1(n12390), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n12279) );
  NAND2_X1 U15739 ( .A1(n12364), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n12278) );
  NAND2_X1 U15740 ( .A1(n12944), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n12277) );
  NAND4_X4 U15741 ( .A1(n12283), .A2(n12282), .A3(n12281), .A4(n12280), .ZN(
        n12288) );
  NAND2_X1 U15742 ( .A1(n12300), .A2(n12295), .ZN(n12284) );
  NOR2_X1 U15743 ( .A1(n12284), .A2(n12303), .ZN(n12286) );
  NOR3_X1 U15744 ( .A1(n12293), .A2(n12288), .A3(n13350), .ZN(n12285) );
  AND2_X1 U15745 ( .A1(n12286), .A2(n12285), .ZN(n13332) );
  NAND2_X1 U15746 ( .A1(n13332), .A2(n12289), .ZN(n13849) );
  AND2_X2 U15747 ( .A1(n13847), .A2(n13849), .ZN(n13340) );
  AND2_X2 U15748 ( .A1(n13324), .A2(n12288), .ZN(n13490) );
  NAND2_X1 U15749 ( .A1(n13490), .A2(n13322), .ZN(n12290) );
  INV_X1 U15750 ( .A(n12313), .ZN(n12287) );
  INV_X2 U15751 ( .A(n12295), .ZN(n21361) );
  NAND2_X1 U15752 ( .A1(n13851), .A2(n13858), .ZN(n13489) );
  AND3_X2 U15753 ( .A1(n13340), .A2(n12290), .A3(n13489), .ZN(n12407) );
  NAND2_X1 U15754 ( .A1(n12320), .A2(n12296), .ZN(n12292) );
  NAND2_X1 U15755 ( .A1(n21361), .A2(n12307), .ZN(n12291) );
  AND2_X1 U15756 ( .A1(n12291), .A2(n12672), .ZN(n12323) );
  NAND2_X1 U15757 ( .A1(n12292), .A2(n12323), .ZN(n13352) );
  INV_X1 U15758 ( .A(n13352), .ZN(n12667) );
  NAND2_X1 U15759 ( .A1(n12672), .A2(n12293), .ZN(n12304) );
  NAND2_X1 U15760 ( .A1(n13331), .A2(n15907), .ZN(n12316) );
  AND2_X2 U15761 ( .A1(n12296), .A2(n12295), .ZN(n13344) );
  NAND2_X1 U15762 ( .A1(n13344), .A2(n13349), .ZN(n13866) );
  INV_X1 U15763 ( .A(n13350), .ZN(n13890) );
  NAND2_X1 U15764 ( .A1(n13890), .A2(n12288), .ZN(n13343) );
  AND2_X1 U15765 ( .A1(n15094), .A2(n13343), .ZN(n12299) );
  OAI211_X1 U15766 ( .C1(n12296), .C2(n15300), .A(n13866), .B(n12299), .ZN(
        n12327) );
  NAND2_X1 U15767 ( .A1(n13385), .A2(n13384), .ZN(n13400) );
  INV_X1 U15768 ( .A(n12301), .ZN(n12302) );
  AND2_X1 U15769 ( .A1(n12304), .A2(n12303), .ZN(n12305) );
  NAND2_X1 U15770 ( .A1(n12295), .A2(n13852), .ZN(n12308) );
  NAND2_X1 U15771 ( .A1(n12312), .A2(n12311), .ZN(n12318) );
  MUX2_X1 U15772 ( .A(n13312), .B(n17625), .S(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Z(n12317) );
  INV_X1 U15773 ( .A(n12320), .ZN(n12321) );
  NAND3_X1 U15774 ( .A1(n15091), .A2(n12321), .A3(n12297), .ZN(n12322) );
  NAND2_X1 U15775 ( .A1(n12319), .A2(n12322), .ZN(n12330) );
  OR2_X1 U15776 ( .A1(n12313), .A2(n13852), .ZN(n13357) );
  INV_X1 U15777 ( .A(n12323), .ZN(n12324) );
  NAND2_X1 U15778 ( .A1(n12324), .A2(n21906), .ZN(n12325) );
  NAND4_X1 U15779 ( .A1(n13357), .A2(n12325), .A3(n15911), .A4(
        P1_STATE2_REG_0__SCAN_IN), .ZN(n12326) );
  NOR2_X1 U15780 ( .A1(n12327), .A2(n12326), .ZN(n12329) );
  NAND3_X1 U15781 ( .A1(n13331), .A2(n15907), .A3(n15303), .ZN(n12328) );
  AOI22_X1 U15782 ( .A1(n12390), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12331), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12339) );
  AOI22_X1 U15783 ( .A1(n13279), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12391), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12338) );
  INV_X2 U15784 ( .A(n12332), .ZN(n13275) );
  AOI22_X1 U15785 ( .A1(n13275), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12267), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12337) );
  INV_X1 U15786 ( .A(n12364), .ZN(n12334) );
  INV_X1 U15787 ( .A(n13075), .ZN(n12335) );
  AOI22_X1 U15788 ( .A1(n12364), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n13244), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12336) );
  INV_X1 U15789 ( .A(n12381), .ZN(n12549) );
  INV_X2 U15790 ( .A(n12549), .ZN(n13053) );
  INV_X1 U15791 ( .A(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12340) );
  INV_X1 U15792 ( .A(n13155), .ZN(n12356) );
  OAI22_X1 U15793 ( .A1(n13053), .A2(n12340), .B1(n12356), .B2(n13284), .ZN(
        n12341) );
  INV_X1 U15794 ( .A(n12341), .ZN(n12347) );
  NAND2_X1 U15795 ( .A1(n13874), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n12346) );
  NAND2_X1 U15796 ( .A1(n12944), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n12345) );
  NAND2_X1 U15797 ( .A1(n12365), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n12344) );
  NAND4_X1 U15798 ( .A1(n12347), .A2(n12346), .A3(n12345), .A4(n12344), .ZN(
        n12352) );
  NAND2_X1 U15799 ( .A1(n13056), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n12350) );
  NAND2_X1 U15800 ( .A1(n12392), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n12349) );
  NAND2_X1 U15801 ( .A1(n13256), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n12348) );
  NAND3_X1 U15802 ( .A1(n12350), .A2(n12349), .A3(n12348), .ZN(n12351) );
  NOR2_X1 U15803 ( .A1(n12352), .A2(n12351), .ZN(n12353) );
  NAND2_X1 U15804 ( .A1(n12944), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n12355) );
  OAI21_X1 U15805 ( .B1(n12379), .B2(n12258), .A(n12355), .ZN(n12359) );
  INV_X1 U15806 ( .A(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12357) );
  OAI22_X1 U15807 ( .A1(n12357), .A2(n12381), .B1(n12356), .B2(n12272), .ZN(
        n12358) );
  NOR2_X1 U15808 ( .A1(n12359), .A2(n12358), .ZN(n12363) );
  AOI22_X1 U15809 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n13275), .B1(
        n12391), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12362) );
  NAND2_X1 U15810 ( .A1(n13056), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n12361) );
  NAND2_X1 U15811 ( .A1(n13874), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n12360) );
  NAND4_X1 U15812 ( .A1(n12363), .A2(n12362), .A3(n12361), .A4(n12360), .ZN(
        n12371) );
  AOI22_X1 U15813 ( .A1(n12364), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12267), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12369) );
  AOI22_X1 U15814 ( .A1(n12365), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12392), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12368) );
  AOI22_X1 U15815 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n12331), .B1(
        n13256), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12367) );
  AOI22_X1 U15816 ( .A1(n12390), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n13244), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12366) );
  NAND4_X1 U15817 ( .A1(n12369), .A2(n12368), .A3(n12367), .A4(n12366), .ZN(
        n12370) );
  XNOR2_X1 U15818 ( .A(n12582), .B(n12534), .ZN(n12372) );
  NAND2_X1 U15819 ( .A1(n12372), .A2(n12441), .ZN(n12373) );
  NAND2_X1 U15820 ( .A1(n12374), .A2(n12373), .ZN(n12532) );
  AOI21_X1 U15821 ( .B1(n12296), .B2(n12579), .A(n21908), .ZN(n12376) );
  NAND2_X1 U15822 ( .A1(n21334), .A2(n12534), .ZN(n12375) );
  NAND2_X1 U15823 ( .A1(n12532), .A2(n12533), .ZN(n12378) );
  NAND2_X1 U15824 ( .A1(n12441), .A2(n12579), .ZN(n12377) );
  NAND2_X1 U15825 ( .A1(n12378), .A2(n12377), .ZN(n12402) );
  NOR2_X1 U15826 ( .A1(n12288), .A2(n21908), .ZN(n12443) );
  NAND2_X1 U15827 ( .A1(n13075), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n12380) );
  OAI21_X1 U15828 ( .B1(n13250), .B2(n13119), .A(n12380), .ZN(n12385) );
  INV_X1 U15829 ( .A(n12381), .ZN(n13240) );
  INV_X1 U15830 ( .A(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12383) );
  INV_X1 U15831 ( .A(n13155), .ZN(n12486) );
  INV_X1 U15832 ( .A(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12382) );
  OAI22_X1 U15833 ( .A1(n13053), .A2(n12383), .B1(n12486), .B2(n12382), .ZN(
        n12384) );
  NOR2_X1 U15834 ( .A1(n12385), .A2(n12384), .ZN(n12389) );
  INV_X2 U15835 ( .A(n13133), .ZN(n13274) );
  AOI22_X1 U15836 ( .A1(n13274), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12267), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12388) );
  NAND2_X1 U15837 ( .A1(n13056), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12387) );
  NAND2_X1 U15838 ( .A1(n12741), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n12386) );
  NAND4_X1 U15839 ( .A1(n12389), .A2(n12388), .A3(n12387), .A4(n12386), .ZN(
        n12398) );
  AOI22_X1 U15840 ( .A1(n12365), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12944), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12396) );
  INV_X1 U15841 ( .A(n12390), .ZN(n13285) );
  INV_X2 U15842 ( .A(n13285), .ZN(n13129) );
  AOI22_X1 U15843 ( .A1(n12364), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n13129), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12395) );
  AOI22_X1 U15844 ( .A1(n13275), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13245), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12394) );
  INV_X1 U15845 ( .A(n13256), .ZN(n13282) );
  AOI22_X1 U15846 ( .A1(n13256), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n12392), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12393) );
  NAND4_X1 U15847 ( .A1(n12396), .A2(n12395), .A3(n12394), .A4(n12393), .ZN(
        n12397) );
  NAND2_X1 U15848 ( .A1(n12443), .A2(n12528), .ZN(n12400) );
  NAND2_X1 U15849 ( .A1(n12441), .A2(n12582), .ZN(n12399) );
  NAND2_X1 U15850 ( .A1(n12402), .A2(n12401), .ZN(n12403) );
  NAND2_X1 U15851 ( .A1(n21729), .A2(n21808), .ZN(n21698) );
  NAND2_X1 U15852 ( .A1(n21698), .A2(n21804), .ZN(n21637) );
  OR2_X1 U15853 ( .A1(n17625), .A2(n21808), .ZN(n12416) );
  OAI21_X1 U15854 ( .B1(n13312), .B2(n21637), .A(n12416), .ZN(n12404) );
  INV_X1 U15855 ( .A(n12404), .ZN(n12405) );
  OAI21_X2 U15856 ( .B1(n12419), .B2(n12406), .A(n12405), .ZN(n12409) );
  INV_X1 U15857 ( .A(n12407), .ZN(n12408) );
  INV_X1 U15858 ( .A(n12410), .ZN(n12411) );
  NAND2_X1 U15859 ( .A1(n12412), .A2(n12411), .ZN(n12413) );
  NAND2_X1 U15860 ( .A1(n21438), .A2(n12413), .ZN(n21381) );
  NAND2_X1 U15861 ( .A1(n12441), .A2(n12528), .ZN(n12414) );
  INV_X1 U15862 ( .A(n12416), .ZN(n12418) );
  INV_X1 U15863 ( .A(n13312), .ZN(n12451) );
  XNOR2_X1 U15864 ( .A(n21804), .B(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n21343) );
  NAND2_X1 U15865 ( .A1(n12451), .A2(n21343), .ZN(n12420) );
  OAI211_X1 U15866 ( .C1(n17625), .C2(n21586), .A(n12421), .B(n12420), .ZN(
        n12424) );
  INV_X1 U15867 ( .A(n12422), .ZN(n12423) );
  NAND2_X1 U15868 ( .A1(n12426), .A2(n12425), .ZN(n12427) );
  INV_X1 U15869 ( .A(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12428) );
  INV_X1 U15870 ( .A(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n13151) );
  OAI22_X1 U15871 ( .A1(n13250), .A2(n12428), .B1(n13175), .B2(n13151), .ZN(
        n12430) );
  INV_X1 U15872 ( .A(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13148) );
  OAI22_X1 U15873 ( .A1(n13053), .A2(n13148), .B1(n12486), .B2(n12212), .ZN(
        n12429) );
  NOR2_X1 U15874 ( .A1(n12430), .A2(n12429), .ZN(n12434) );
  AOI22_X1 U15875 ( .A1(n13275), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13245), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12433) );
  NAND2_X1 U15876 ( .A1(n13874), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n12432) );
  NAND2_X1 U15877 ( .A1(n13056), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n12431) );
  NAND4_X1 U15878 ( .A1(n12434), .A2(n12433), .A3(n12432), .A4(n12431), .ZN(
        n12440) );
  AOI22_X1 U15879 ( .A1(n13255), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n13129), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12438) );
  AOI22_X1 U15880 ( .A1(n13061), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n13244), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12437) );
  AOI22_X1 U15881 ( .A1(n12267), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n13256), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12436) );
  AOI22_X1 U15882 ( .A1(n13274), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12392), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12435) );
  NAND4_X1 U15883 ( .A1(n12438), .A2(n12437), .A3(n12436), .A4(n12435), .ZN(
        n12439) );
  NAND2_X1 U15884 ( .A1(n12441), .A2(n12503), .ZN(n12442) );
  AOI22_X1 U15885 ( .A1(n12624), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12443), .B2(n12503), .ZN(n12444) );
  OAI21_X1 U15886 ( .B1(n21804), .B2(n21586), .A(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n12449) );
  INV_X1 U15887 ( .A(n21804), .ZN(n12448) );
  NAND2_X1 U15888 ( .A1(n21636), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n21524) );
  INV_X1 U15889 ( .A(n21524), .ZN(n12447) );
  NAND2_X1 U15890 ( .A1(n12448), .A2(n12447), .ZN(n21554) );
  NAND2_X1 U15891 ( .A1(n12449), .A2(n21554), .ZN(n21587) );
  INV_X1 U15892 ( .A(n17625), .ZN(n12450) );
  AOI22_X1 U15893 ( .A1(n12451), .A2(n21587), .B1(n12450), .B2(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n12452) );
  INV_X1 U15894 ( .A(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12914) );
  OAI22_X1 U15895 ( .A1(n13250), .A2(n13172), .B1(n13221), .B2(n12914), .ZN(
        n12457) );
  INV_X1 U15896 ( .A(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12455) );
  INV_X1 U15897 ( .A(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12454) );
  OAI22_X1 U15898 ( .A1(n13053), .A2(n12455), .B1(n12486), .B2(n12454), .ZN(
        n12456) );
  NOR2_X1 U15899 ( .A1(n12457), .A2(n12456), .ZN(n12461) );
  AOI22_X1 U15900 ( .A1(n13275), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13245), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12460) );
  NAND2_X1 U15901 ( .A1(n12741), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n12459) );
  NAND2_X1 U15902 ( .A1(n13056), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n12458) );
  NAND4_X1 U15903 ( .A1(n12461), .A2(n12460), .A3(n12459), .A4(n12458), .ZN(
        n12467) );
  AOI22_X1 U15904 ( .A1(n13255), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n13129), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12465) );
  AOI22_X1 U15905 ( .A1(n13061), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n13244), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12464) );
  AOI22_X1 U15906 ( .A1(n13254), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n13256), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12463) );
  AOI22_X1 U15907 ( .A1(n13274), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12392), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12462) );
  NAND4_X1 U15908 ( .A1(n12465), .A2(n12464), .A3(n12463), .A4(n12462), .ZN(
        n12466) );
  AOI22_X1 U15909 ( .A1(n12624), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12664), .B2(n12516), .ZN(n12468) );
  NAND2_X1 U15910 ( .A1(n12624), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n12485) );
  INV_X1 U15911 ( .A(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n13194) );
  NAND2_X1 U15912 ( .A1(n13075), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n12469) );
  OAI21_X1 U15913 ( .B1(n13194), .B2(n13175), .A(n12469), .ZN(n12473) );
  INV_X1 U15914 ( .A(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12471) );
  OAI22_X1 U15915 ( .A1(n13053), .A2(n12471), .B1(n12486), .B2(n12470), .ZN(
        n12472) );
  NOR2_X1 U15916 ( .A1(n12473), .A2(n12472), .ZN(n12477) );
  AOI22_X1 U15917 ( .A1(n13254), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n13256), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12476) );
  NAND2_X1 U15918 ( .A1(n13056), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n12475) );
  NAND2_X1 U15919 ( .A1(n13874), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n12474) );
  NAND4_X1 U15920 ( .A1(n12477), .A2(n12476), .A3(n12475), .A4(n12474), .ZN(
        n12483) );
  AOI22_X1 U15921 ( .A1(n13279), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12944), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12481) );
  AOI22_X1 U15922 ( .A1(n13255), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n13129), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12480) );
  AOI22_X1 U15923 ( .A1(n13275), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n13245), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12479) );
  AOI22_X1 U15924 ( .A1(n13274), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n12392), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12478) );
  NAND4_X1 U15925 ( .A1(n12481), .A2(n12480), .A3(n12479), .A4(n12478), .ZN(
        n12482) );
  NAND2_X1 U15926 ( .A1(n12664), .A2(n12510), .ZN(n12484) );
  INV_X1 U15927 ( .A(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12865) );
  OAI22_X1 U15928 ( .A1(n13250), .A2(n12116), .B1(n13175), .B2(n12865), .ZN(
        n12490) );
  INV_X1 U15929 ( .A(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12487) );
  OAI22_X1 U15930 ( .A1(n13053), .A2(n12488), .B1(n12486), .B2(n12487), .ZN(
        n12489) );
  NOR2_X1 U15931 ( .A1(n12490), .A2(n12489), .ZN(n12494) );
  AOI22_X1 U15932 ( .A1(n13275), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n13245), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12493) );
  NAND2_X1 U15933 ( .A1(n13874), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n12492) );
  NAND2_X1 U15934 ( .A1(n13056), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n12491) );
  NAND4_X1 U15935 ( .A1(n12494), .A2(n12493), .A3(n12492), .A4(n12491), .ZN(
        n12500) );
  AOI22_X1 U15936 ( .A1(n13255), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n13129), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12498) );
  AOI22_X1 U15937 ( .A1(n13061), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n13244), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12497) );
  AOI22_X1 U15938 ( .A1(n13254), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n13256), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12496) );
  INV_X1 U15939 ( .A(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n21979) );
  AOI22_X1 U15940 ( .A1(n13274), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12392), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12495) );
  NAND4_X1 U15941 ( .A1(n12498), .A2(n12497), .A3(n12496), .A4(n12495), .ZN(
        n12499) );
  NAND2_X1 U15942 ( .A1(n12664), .A2(n12505), .ZN(n12501) );
  OAI21_X1 U15943 ( .B1(n12654), .B2(n12867), .A(n12501), .ZN(n12502) );
  INV_X1 U15944 ( .A(n12502), .ZN(n12566) );
  INV_X1 U15945 ( .A(n12623), .ZN(n13827) );
  INV_X1 U15946 ( .A(n12503), .ZN(n12523) );
  NAND2_X1 U15947 ( .A1(n12534), .A2(n12528), .ZN(n12522) );
  NAND2_X1 U15948 ( .A1(n12523), .A2(n12522), .ZN(n12521) );
  NAND2_X1 U15949 ( .A1(n12521), .A2(n12516), .ZN(n12515) );
  INV_X1 U15950 ( .A(n12510), .ZN(n12504) );
  NOR2_X1 U15951 ( .A1(n12515), .A2(n12504), .ZN(n12506) );
  NAND2_X1 U15952 ( .A1(n12506), .A2(n12505), .ZN(n12575) );
  OAI211_X1 U15953 ( .C1(n12506), .C2(n12505), .A(n12575), .B(n21906), .ZN(
        n12507) );
  INV_X1 U15954 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n15756) );
  NAND2_X1 U15955 ( .A1(n12514), .A2(n12508), .ZN(n12509) );
  NAND2_X1 U15956 ( .A1(n12548), .A2(n12509), .ZN(n12690) );
  XNOR2_X1 U15957 ( .A(n12515), .B(n12510), .ZN(n12511) );
  NAND2_X1 U15958 ( .A1(n12511), .A2(n21906), .ZN(n12512) );
  OAI211_X1 U15959 ( .C1(n12516), .C2(n12521), .A(n12515), .B(n21906), .ZN(
        n12517) );
  NAND3_X1 U15960 ( .A1(n15579), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n12545) );
  BUF_X1 U15961 ( .A(n12518), .Z(n12519) );
  NAND2_X1 U15962 ( .A1(n15888), .A2(n12623), .ZN(n12527) );
  OAI21_X1 U15963 ( .B1(n12523), .B2(n12522), .A(n12521), .ZN(n12525) );
  NAND2_X1 U15964 ( .A1(n21334), .A2(n12297), .ZN(n12535) );
  INV_X1 U15965 ( .A(n12535), .ZN(n12524) );
  AOI21_X1 U15966 ( .B1(n12525), .B2(n21906), .A(n12524), .ZN(n12526) );
  NAND2_X1 U15967 ( .A1(n12527), .A2(n12526), .ZN(n14071) );
  XNOR2_X1 U15968 ( .A(n12528), .B(n12534), .ZN(n12529) );
  OAI211_X1 U15969 ( .C1(n12529), .C2(n15300), .A(n13350), .B(n12618), .ZN(
        n12530) );
  INV_X1 U15970 ( .A(n12530), .ZN(n12531) );
  OR2_X1 U15971 ( .A1(n15300), .A2(n12534), .ZN(n12536) );
  AND2_X1 U15972 ( .A1(n12536), .A2(n12535), .ZN(n13826) );
  NAND3_X1 U15973 ( .A1(n12536), .A2(n13827), .A3(n12535), .ZN(n12537) );
  AND2_X1 U15974 ( .A1(n12537), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12538) );
  NAND2_X1 U15975 ( .A1(n13910), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12542) );
  INV_X1 U15976 ( .A(n13828), .ZN(n12540) );
  NAND2_X1 U15977 ( .A1(n12540), .A2(n12539), .ZN(n12541) );
  INV_X1 U15978 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n15752) );
  NAND2_X1 U15979 ( .A1(n12543), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12544) );
  INV_X1 U15980 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n15569) );
  NAND2_X1 U15981 ( .A1(n12546), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12547) );
  NAND2_X1 U15982 ( .A1(n12624), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n12565) );
  NAND2_X1 U15983 ( .A1(n13129), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n12553) );
  NAND2_X1 U15984 ( .A1(n13061), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n12552) );
  NAND2_X1 U15985 ( .A1(n12549), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n12551) );
  NAND2_X1 U15986 ( .A1(n13155), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n12550) );
  AND4_X1 U15987 ( .A1(n12553), .A2(n12552), .A3(n12551), .A4(n12550), .ZN(
        n12557) );
  AOI22_X1 U15988 ( .A1(n13245), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n13256), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12556) );
  NAND2_X1 U15989 ( .A1(n13056), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n12555) );
  NAND2_X1 U15990 ( .A1(n12741), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n12554) );
  NAND4_X1 U15991 ( .A1(n12557), .A2(n12556), .A3(n12555), .A4(n12554), .ZN(
        n12563) );
  AOI22_X1 U15992 ( .A1(n12365), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n13274), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12561) );
  AOI22_X1 U15993 ( .A1(n13279), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n13244), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12560) );
  AOI22_X1 U15994 ( .A1(n13275), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13254), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12559) );
  AOI22_X1 U15995 ( .A1(n13255), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12392), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12558) );
  NAND4_X1 U15996 ( .A1(n12561), .A2(n12560), .A3(n12559), .A4(n12558), .ZN(
        n12562) );
  NAND2_X1 U15997 ( .A1(n12664), .A2(n12573), .ZN(n12564) );
  NAND2_X1 U15998 ( .A1(n12568), .A2(n12567), .ZN(n12728) );
  NAND3_X1 U15999 ( .A1(n12581), .A2(n12728), .A3(n12623), .ZN(n12571) );
  XNOR2_X1 U16000 ( .A(n12575), .B(n12573), .ZN(n12569) );
  NAND2_X1 U16001 ( .A1(n12569), .A2(n21906), .ZN(n12570) );
  NAND2_X1 U16002 ( .A1(n12571), .A2(n12570), .ZN(n12587) );
  OR2_X1 U16003 ( .A1(n12587), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17664) );
  INV_X1 U16004 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13081) );
  OAI22_X1 U16005 ( .A1(n12654), .A2(n13081), .B1(n12626), .B2(n12582), .ZN(
        n12572) );
  NAND2_X1 U16006 ( .A1(n12729), .A2(n12623), .ZN(n12578) );
  INV_X1 U16007 ( .A(n12573), .ZN(n12574) );
  XNOR2_X1 U16008 ( .A(n12584), .B(n12579), .ZN(n12576) );
  NAND2_X1 U16009 ( .A1(n12576), .A2(n21906), .ZN(n12577) );
  NAND2_X1 U16010 ( .A1(n12578), .A2(n12577), .ZN(n15532) );
  OR2_X1 U16011 ( .A1(n15300), .A2(n12582), .ZN(n12583) );
  NOR2_X1 U16012 ( .A1(n12584), .A2(n12583), .ZN(n12591) );
  NAND2_X1 U16013 ( .A1(n12591), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12586) );
  NOR2_X1 U16014 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n12585) );
  AOI21_X1 U16015 ( .B1(n15554), .B2(n12586), .A(n12585), .ZN(n12590) );
  OAI21_X1 U16016 ( .B1(n17663), .B2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n15532), .ZN(n12589) );
  INV_X1 U16017 ( .A(n12591), .ZN(n15533) );
  INV_X1 U16018 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n15561) );
  NAND2_X1 U16019 ( .A1(n15533), .A2(n15561), .ZN(n12592) );
  NAND2_X1 U16020 ( .A1(n12592), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12593) );
  NAND2_X1 U16021 ( .A1(n15554), .A2(n12593), .ZN(n12594) );
  NAND2_X1 U16022 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n12595) );
  NAND2_X1 U16023 ( .A1(n15554), .A2(n12595), .ZN(n15516) );
  INV_X1 U16024 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15798) );
  INV_X1 U16025 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15758) );
  INV_X1 U16026 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15504) );
  NAND2_X1 U16027 ( .A1(n15758), .A2(n15504), .ZN(n15495) );
  NOR2_X1 U16028 ( .A1(n15495), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12599) );
  XNOR2_X1 U16029 ( .A(n15554), .B(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15483) );
  INV_X1 U16030 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15739) );
  NAND2_X1 U16031 ( .A1(n15554), .A2(n15739), .ZN(n12600) );
  NAND2_X1 U16032 ( .A1(n15483), .A2(n12600), .ZN(n15481) );
  INV_X1 U16033 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15534) );
  INV_X1 U16034 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15807) );
  NAND2_X1 U16035 ( .A1(n15534), .A2(n15807), .ZN(n15515) );
  NOR2_X1 U16036 ( .A1(n15515), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12601) );
  XNOR2_X1 U16037 ( .A(n15554), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15461) );
  NAND2_X1 U16038 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15647) );
  INV_X1 U16039 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15672) );
  NOR2_X1 U16040 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15390) );
  INV_X1 U16041 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15650) );
  INV_X1 U16042 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15617) );
  AND2_X1 U16043 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n13373) );
  NAND3_X1 U16044 ( .A1(n13373), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15384) );
  AND2_X1 U16045 ( .A1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n13379) );
  INV_X1 U16046 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15367) );
  NAND2_X1 U16047 ( .A1(n12607), .A2(n15367), .ZN(n12608) );
  INV_X1 U16048 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15357) );
  MUX2_X1 U16049 ( .A(n15357), .B(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .S(
        n15554), .Z(n12610) );
  NAND2_X1 U16050 ( .A1(n12612), .A2(n15303), .ZN(n12613) );
  NAND2_X1 U16051 ( .A1(n12613), .A2(n12618), .ZN(n12614) );
  NAND2_X1 U16052 ( .A1(n12614), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12616) );
  NAND2_X1 U16053 ( .A1(n12616), .A2(n15303), .ZN(n12615) );
  XNOR2_X1 U16054 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n12633) );
  XNOR2_X1 U16055 ( .A(n12633), .B(n12634), .ZN(n13317) );
  NAND2_X1 U16056 ( .A1(n12615), .A2(n13317), .ZN(n12630) );
  INV_X1 U16057 ( .A(n13317), .ZN(n12617) );
  OAI21_X1 U16058 ( .B1(n12654), .B2(n12617), .A(n12616), .ZN(n12629) );
  NAND2_X1 U16059 ( .A1(n12289), .A2(n12618), .ZN(n12619) );
  AND2_X1 U16060 ( .A1(n15091), .A2(n12619), .ZN(n12640) );
  INV_X1 U16061 ( .A(n12634), .ZN(n12621) );
  NAND2_X1 U16062 ( .A1(n13945), .A2(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n12620) );
  NAND2_X1 U16063 ( .A1(n12621), .A2(n12620), .ZN(n12625) );
  INV_X1 U16064 ( .A(n12625), .ZN(n12622) );
  OAI211_X1 U16065 ( .C1(n21334), .C2(n12668), .A(n12640), .B(n12622), .ZN(
        n12628) );
  OAI21_X1 U16066 ( .B1(n12626), .B2(n12625), .A(n12658), .ZN(n12627) );
  OAI211_X1 U16067 ( .C1(n12630), .C2(n12629), .A(n12628), .B(n12627), .ZN(
        n12632) );
  NAND2_X1 U16068 ( .A1(n12630), .A2(n12629), .ZN(n12631) );
  NAND2_X1 U16069 ( .A1(n12634), .A2(n12633), .ZN(n12636) );
  NAND2_X1 U16070 ( .A1(n21808), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12635) );
  NAND2_X1 U16071 ( .A1(n12636), .A2(n12635), .ZN(n12645) );
  XNOR2_X1 U16072 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n12644) );
  XNOR2_X1 U16073 ( .A(n12645), .B(n12644), .ZN(n13316) );
  INV_X1 U16074 ( .A(n13316), .ZN(n12637) );
  NAND2_X1 U16075 ( .A1(n12664), .A2(n12637), .ZN(n12639) );
  OAI211_X1 U16076 ( .C1(n12637), .C2(n12654), .A(n12639), .B(n12640), .ZN(
        n12638) );
  INV_X1 U16077 ( .A(n12639), .ZN(n12642) );
  INV_X1 U16078 ( .A(n12640), .ZN(n12641) );
  NAND2_X1 U16079 ( .A1(n12642), .A2(n12641), .ZN(n12643) );
  NAND2_X1 U16080 ( .A1(n12645), .A2(n12644), .ZN(n12647) );
  NAND2_X1 U16081 ( .A1(n21586), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12646) );
  NAND2_X1 U16082 ( .A1(n12647), .A2(n12646), .ZN(n12649) );
  XNOR2_X1 U16083 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n12648) );
  NOR2_X1 U16084 ( .A1(n12649), .A2(n12648), .ZN(n12650) );
  OR2_X1 U16085 ( .A1(n12653), .A2(n12650), .ZN(n13318) );
  INV_X1 U16086 ( .A(n12658), .ZN(n12663) );
  NAND2_X1 U16087 ( .A1(n12663), .A2(n13318), .ZN(n12651) );
  NAND2_X1 U16088 ( .A1(n12652), .A2(n12651), .ZN(n12657) );
  NAND3_X1 U16089 ( .A1(n15872), .A2(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A3(
        n12662), .ZN(n13319) );
  INV_X1 U16090 ( .A(n13319), .ZN(n12655) );
  NAND2_X1 U16091 ( .A1(n12655), .A2(n12654), .ZN(n12656) );
  OAI22_X1 U16092 ( .A1(n12658), .A2(n13319), .B1(P1_STATE2_REG_0__SCAN_IN), 
        .B2(n15872), .ZN(n12659) );
  INV_X1 U16093 ( .A(n12659), .ZN(n12660) );
  NAND2_X1 U16094 ( .A1(n15907), .A2(n21334), .ZN(n12666) );
  NAND3_X1 U16095 ( .A1(n12667), .A2(n12301), .A3(n12666), .ZN(n13338) );
  INV_X1 U16096 ( .A(n21153), .ZN(n12669) );
  INV_X1 U16097 ( .A(n12670), .ZN(n12680) );
  INV_X1 U16098 ( .A(n13303), .ZN(n12733) );
  INV_X1 U16099 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17677) );
  NAND2_X1 U16100 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12691) );
  INV_X1 U16101 ( .A(n12724), .ZN(n12675) );
  INV_X1 U16102 ( .A(n12686), .ZN(n12673) );
  NAND2_X1 U16103 ( .A1(n12673), .A2(n17677), .ZN(n12674) );
  NAND2_X1 U16104 ( .A1(n12675), .A2(n12674), .ZN(n21218) );
  NAND2_X1 U16105 ( .A1(n21218), .A2(n13526), .ZN(n12676) );
  OAI21_X1 U16106 ( .B1(n12733), .B2(n17677), .A(n12676), .ZN(n12677) );
  AOI21_X1 U16107 ( .B1(n13232), .B2(P1_EAX_REG_5__SCAN_IN), .A(n12677), .ZN(
        n12678) );
  AOI21_X1 U16108 ( .B1(n12680), .B2(n12930), .A(n12679), .ZN(n12681) );
  INV_X1 U16109 ( .A(n12681), .ZN(n15168) );
  NAND2_X1 U16110 ( .A1(n13858), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12718) );
  OAI21_X1 U16111 ( .B1(n21905), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n12682), .ZN(n12684) );
  NAND2_X1 U16112 ( .A1(n12723), .A2(P1_EAX_REG_4__SCAN_IN), .ZN(n12683) );
  OAI211_X1 U16113 ( .C1(n12718), .C2(n15872), .A(n12684), .B(n12683), .ZN(
        n12688) );
  NOR2_X1 U16114 ( .A1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n12692), .ZN(
        n12685) );
  NOR2_X1 U16115 ( .A1(n12686), .A2(n12685), .ZN(n21231) );
  NAND2_X1 U16116 ( .A1(n21231), .A2(n13267), .ZN(n12687) );
  NAND2_X1 U16117 ( .A1(n12688), .A2(n12687), .ZN(n12689) );
  INV_X1 U16118 ( .A(n12691), .ZN(n12694) );
  INV_X1 U16119 ( .A(n12692), .ZN(n12693) );
  OAI21_X1 U16120 ( .B1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n12694), .A(
        n12693), .ZN(n21262) );
  AOI22_X1 U16121 ( .A1(n13526), .A2(n21262), .B1(n13303), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n12696) );
  NAND2_X1 U16122 ( .A1(n13232), .A2(P1_EAX_REG_3__SCAN_IN), .ZN(n12695) );
  OAI211_X1 U16123 ( .C1(n12718), .C2(n12697), .A(n12696), .B(n12695), .ZN(
        n12698) );
  INV_X1 U16124 ( .A(n12698), .ZN(n12699) );
  XNOR2_X2 U16125 ( .A(n9804), .B(n10455), .ZN(n15884) );
  NAND2_X1 U16126 ( .A1(n15884), .A2(n12930), .ZN(n12706) );
  AOI22_X1 U16127 ( .A1(n13232), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n12682), .ZN(n12704) );
  INV_X1 U16128 ( .A(n12718), .ZN(n12702) );
  NAND2_X1 U16129 ( .A1(n12702), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12703) );
  AND2_X1 U16130 ( .A1(n12704), .A2(n12703), .ZN(n12705) );
  NAND2_X1 U16131 ( .A1(n9734), .A2(n21365), .ZN(n12707) );
  NAND2_X1 U16132 ( .A1(n12707), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13836) );
  NAND2_X1 U16133 ( .A1(n12682), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12711) );
  NAND2_X1 U16134 ( .A1(n13232), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n12710) );
  OAI211_X1 U16135 ( .C1(n12718), .C2(n13945), .A(n12711), .B(n12710), .ZN(
        n12712) );
  AOI21_X1 U16136 ( .B1(n12709), .B2(n12930), .A(n12712), .ZN(n13837) );
  NAND2_X1 U16137 ( .A1(n13837), .A2(n13267), .ZN(n12713) );
  NAND2_X1 U16138 ( .A1(n13838), .A2(n12713), .ZN(n13932) );
  NAND2_X1 U16139 ( .A1(n13303), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n15178) );
  NAND2_X1 U16140 ( .A1(n14115), .A2(n15178), .ZN(n12714) );
  AND2_X1 U16141 ( .A1(n15180), .A2(n12714), .ZN(n12722) );
  NAND2_X1 U16142 ( .A1(n15888), .A2(n12930), .ZN(n12721) );
  XNOR2_X1 U16143 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n15104) );
  AOI21_X1 U16144 ( .B1(n13526), .B2(n15104), .A(n13303), .ZN(n12716) );
  NAND2_X1 U16145 ( .A1(n13232), .A2(P1_EAX_REG_2__SCAN_IN), .ZN(n12715) );
  OAI211_X1 U16146 ( .C1(n12718), .C2(n12717), .A(n12716), .B(n12715), .ZN(
        n12719) );
  INV_X1 U16147 ( .A(n12719), .ZN(n12720) );
  NAND2_X1 U16148 ( .A1(n12721), .A2(n12720), .ZN(n14114) );
  INV_X1 U16149 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n12726) );
  OAI21_X1 U16150 ( .B1(n12724), .B2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n12730), .ZN(n21206) );
  AOI22_X1 U16151 ( .A1(n21206), .A2(n13526), .B1(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n13303), .ZN(n12725) );
  OAI21_X1 U16152 ( .B1(n12884), .B2(n12726), .A(n12725), .ZN(n12727) );
  AOI21_X1 U16153 ( .B1(n12728), .B2(n12930), .A(n12727), .ZN(n15163) );
  NAND2_X1 U16154 ( .A1(n12729), .A2(n12930), .ZN(n12736) );
  AND2_X1 U16155 ( .A1(n12730), .A2(n21194), .ZN(n12731) );
  OR2_X1 U16156 ( .A1(n12731), .A2(n12771), .ZN(n21196) );
  NAND2_X1 U16157 ( .A1(n21196), .A2(n13267), .ZN(n12732) );
  OAI21_X1 U16158 ( .B1(n12733), .B2(n21194), .A(n12732), .ZN(n12734) );
  AOI21_X1 U16159 ( .B1(n13232), .B2(P1_EAX_REG_7__SCAN_IN), .A(n12734), .ZN(
        n12735) );
  NAND2_X1 U16160 ( .A1(n12736), .A2(n12735), .ZN(n15157) );
  AOI22_X1 U16161 ( .A1(n12723), .A2(P1_EAX_REG_8__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n13303), .ZN(n12754) );
  INV_X1 U16162 ( .A(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12799) );
  NAND2_X1 U16163 ( .A1(n13061), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n12737) );
  OAI21_X1 U16164 ( .B1(n13175), .B2(n12799), .A(n12737), .ZN(n12740) );
  INV_X1 U16165 ( .A(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12738) );
  OAI22_X1 U16166 ( .A1(n13092), .A2(n13053), .B1(n12356), .B2(n12738), .ZN(
        n12739) );
  NOR2_X1 U16167 ( .A1(n12740), .A2(n12739), .ZN(n12745) );
  AOI22_X1 U16168 ( .A1(n13245), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12392), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12744) );
  NAND2_X1 U16169 ( .A1(n13056), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n12743) );
  NAND2_X1 U16170 ( .A1(n12741), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n12742) );
  NAND4_X1 U16171 ( .A1(n12745), .A2(n12744), .A3(n12743), .A4(n12742), .ZN(
        n12751) );
  AOI22_X1 U16172 ( .A1(n13275), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n13274), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12749) );
  AOI22_X1 U16173 ( .A1(n13279), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n13244), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12748) );
  AOI22_X1 U16174 ( .A1(n13255), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n13254), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12747) );
  AOI22_X1 U16175 ( .A1(n13129), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n13256), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12746) );
  NAND4_X1 U16176 ( .A1(n12749), .A2(n12748), .A3(n12747), .A4(n12746), .ZN(
        n12750) );
  OR2_X1 U16177 ( .A1(n12751), .A2(n12750), .ZN(n12752) );
  XNOR2_X1 U16178 ( .A(n12771), .B(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n21186) );
  AOI22_X1 U16179 ( .A1(n12930), .A2(n12752), .B1(n13526), .B2(n21186), .ZN(
        n12753) );
  AOI22_X1 U16180 ( .A1(n12365), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13255), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12759) );
  AOI22_X1 U16181 ( .A1(n13129), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n13244), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12758) );
  AOI22_X1 U16182 ( .A1(n13275), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n13256), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12757) );
  AOI22_X1 U16183 ( .A1(n13254), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12392), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12756) );
  NAND4_X1 U16184 ( .A1(n12759), .A2(n12758), .A3(n12757), .A4(n12756), .ZN(
        n12770) );
  INV_X1 U16185 ( .A(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13128) );
  NAND2_X1 U16186 ( .A1(n13061), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n12760) );
  OAI21_X1 U16187 ( .B1(n13128), .B2(n13250), .A(n12760), .ZN(n12764) );
  INV_X1 U16188 ( .A(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12761) );
  OAI22_X1 U16189 ( .A1(n13053), .A2(n12762), .B1(n12356), .B2(n12761), .ZN(
        n12763) );
  NOR2_X1 U16190 ( .A1(n12764), .A2(n12763), .ZN(n12768) );
  AOI22_X1 U16191 ( .A1(n13274), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n13245), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12767) );
  NAND2_X1 U16192 ( .A1(n13056), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n12766) );
  NAND2_X1 U16193 ( .A1(n13874), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n12765) );
  NAND4_X1 U16194 ( .A1(n12768), .A2(n12767), .A3(n12766), .A4(n12765), .ZN(
        n12769) );
  OAI21_X1 U16195 ( .B1(n12770), .B2(n12769), .A(n12930), .ZN(n12775) );
  XOR2_X1 U16196 ( .A(n15557), .B(n12776), .Z(n21175) );
  INV_X1 U16197 ( .A(n21175), .ZN(n12772) );
  AOI22_X1 U16198 ( .A1(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n13303), .B1(
        n13526), .B2(n12772), .ZN(n12774) );
  NAND2_X1 U16199 ( .A1(n13232), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n12773) );
  XNOR2_X1 U16200 ( .A(n12795), .B(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n17642) );
  OR2_X1 U16201 ( .A1(n17642), .A2(n13302), .ZN(n12794) );
  NAND2_X1 U16202 ( .A1(n13232), .A2(P1_EAX_REG_10__SCAN_IN), .ZN(n12793) );
  AOI22_X1 U16203 ( .A1(n13255), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12944), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12780) );
  AOI22_X1 U16204 ( .A1(n13129), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n13244), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12779) );
  AOI22_X1 U16205 ( .A1(n13254), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n13256), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12778) );
  AOI22_X1 U16206 ( .A1(n13245), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12392), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12777) );
  NAND4_X1 U16207 ( .A1(n12780), .A2(n12779), .A3(n12778), .A4(n12777), .ZN(
        n12790) );
  INV_X1 U16208 ( .A(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12781) );
  OAI22_X1 U16209 ( .A1(n13250), .A2(n13151), .B1(n13221), .B2(n12781), .ZN(
        n12784) );
  INV_X1 U16210 ( .A(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13147) );
  INV_X1 U16211 ( .A(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12782) );
  OAI22_X1 U16212 ( .A1(n13053), .A2(n13147), .B1(n12486), .B2(n12782), .ZN(
        n12783) );
  NOR2_X1 U16213 ( .A1(n12784), .A2(n12783), .ZN(n12788) );
  AOI22_X1 U16214 ( .A1(n13275), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13274), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12787) );
  NAND2_X1 U16215 ( .A1(n13056), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n12786) );
  NAND2_X1 U16216 ( .A1(n13874), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n12785) );
  NAND4_X1 U16217 ( .A1(n12788), .A2(n12787), .A3(n12786), .A4(n12785), .ZN(
        n12789) );
  OAI21_X1 U16218 ( .B1(n12790), .B2(n12789), .A(n12930), .ZN(n12792) );
  NAND2_X1 U16219 ( .A1(n13303), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12791) );
  NAND4_X1 U16220 ( .A1(n12794), .A2(n12793), .A3(n12792), .A4(n12791), .ZN(
        n15140) );
  INV_X1 U16221 ( .A(n12796), .ZN(n12797) );
  INV_X1 U16222 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n15485) );
  NAND2_X1 U16223 ( .A1(n12797), .A2(n15485), .ZN(n12798) );
  AND2_X1 U16224 ( .A1(n12954), .A2(n12798), .ZN(n15489) );
  INV_X1 U16225 ( .A(n15907), .ZN(n13872) );
  INV_X1 U16226 ( .A(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n13094) );
  OAI22_X1 U16227 ( .A1(n12799), .A2(n13250), .B1(n13175), .B2(n13094), .ZN(
        n12803) );
  INV_X1 U16228 ( .A(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12801) );
  OAI22_X1 U16229 ( .A1(n12801), .A2(n13053), .B1(n12486), .B2(n12800), .ZN(
        n12802) );
  NOR2_X1 U16230 ( .A1(n12803), .A2(n12802), .ZN(n12807) );
  AOI22_X1 U16231 ( .A1(n13275), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n13274), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12806) );
  NAND2_X1 U16232 ( .A1(n13056), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n12805) );
  NAND2_X1 U16233 ( .A1(n13874), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n12804) );
  NAND4_X1 U16234 ( .A1(n12807), .A2(n12806), .A3(n12805), .A4(n12804), .ZN(
        n12813) );
  AOI22_X1 U16235 ( .A1(n13255), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n13129), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12811) );
  AOI22_X1 U16236 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n13245), .B1(
        n13244), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12810) );
  AOI22_X1 U16237 ( .A1(n13061), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n13256), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12809) );
  AOI22_X1 U16238 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n13254), .B1(
        n12392), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12808) );
  NAND4_X1 U16239 ( .A1(n12811), .A2(n12810), .A3(n12809), .A4(n12808), .ZN(
        n12812) );
  OR2_X1 U16240 ( .A1(n12813), .A2(n12812), .ZN(n12816) );
  INV_X1 U16241 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n15277) );
  NAND2_X1 U16242 ( .A1(n12682), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12814) );
  OAI211_X1 U16243 ( .C1(n12884), .C2(n15277), .A(n13302), .B(n12814), .ZN(
        n12815) );
  AOI21_X1 U16244 ( .B1(n13264), .B2(n12816), .A(n12815), .ZN(n12817) );
  AOI21_X1 U16245 ( .B1(n15489), .B2(n13526), .A(n12817), .ZN(n14992) );
  INV_X1 U16246 ( .A(n12818), .ZN(n12820) );
  INV_X1 U16247 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n12819) );
  XNOR2_X1 U16248 ( .A(n12820), .B(n12819), .ZN(n15492) );
  NAND2_X1 U16249 ( .A1(n15492), .A2(n13267), .ZN(n12839) );
  AOI22_X1 U16250 ( .A1(n13255), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n13274), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12824) );
  AOI22_X1 U16251 ( .A1(n13061), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n13245), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12823) );
  AOI22_X1 U16252 ( .A1(n13279), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n13244), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12822) );
  AOI22_X1 U16253 ( .A1(n13275), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12392), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12821) );
  NAND4_X1 U16254 ( .A1(n12824), .A2(n12823), .A3(n12822), .A4(n12821), .ZN(
        n12834) );
  INV_X1 U16255 ( .A(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n13287) );
  NAND2_X1 U16256 ( .A1(n13256), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n12825) );
  OAI21_X1 U16257 ( .B1(n13287), .B2(n13175), .A(n12825), .ZN(n12828) );
  INV_X1 U16258 ( .A(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12826) );
  OAI22_X1 U16259 ( .A1(n13053), .A2(n13081), .B1(n12356), .B2(n12826), .ZN(
        n12827) );
  NOR2_X1 U16260 ( .A1(n12828), .A2(n12827), .ZN(n12832) );
  AOI22_X1 U16261 ( .A1(n13129), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n13254), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12831) );
  NAND2_X1 U16262 ( .A1(n13874), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n12830) );
  NAND2_X1 U16263 ( .A1(n13056), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n12829) );
  NAND4_X1 U16264 ( .A1(n12832), .A2(n12831), .A3(n12830), .A4(n12829), .ZN(
        n12833) );
  OAI21_X1 U16265 ( .B1(n12834), .B2(n12833), .A(n12930), .ZN(n12837) );
  NAND2_X1 U16266 ( .A1(n12723), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n12836) );
  NAND2_X1 U16267 ( .A1(n13303), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12835) );
  AND3_X1 U16268 ( .A1(n12837), .A2(n12836), .A3(n12835), .ZN(n12838) );
  NAND2_X1 U16269 ( .A1(n12839), .A2(n12838), .ZN(n15013) );
  XNOR2_X1 U16270 ( .A(n12841), .B(n12840), .ZN(n15502) );
  NAND2_X1 U16271 ( .A1(n15502), .A2(n13267), .ZN(n12862) );
  AOI22_X1 U16272 ( .A1(n12365), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13255), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12845) );
  AOI22_X1 U16273 ( .A1(n13254), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n13244), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12844) );
  AOI22_X1 U16274 ( .A1(n13275), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n13256), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12843) );
  AOI22_X1 U16275 ( .A1(n13129), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12392), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12842) );
  NAND4_X1 U16276 ( .A1(n12845), .A2(n12844), .A3(n12843), .A4(n12842), .ZN(
        n12857) );
  INV_X1 U16277 ( .A(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12847) );
  NAND2_X1 U16278 ( .A1(n13061), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n12846) );
  OAI21_X1 U16279 ( .B1(n12847), .B2(n13250), .A(n12846), .ZN(n12851) );
  INV_X1 U16280 ( .A(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12849) );
  INV_X1 U16281 ( .A(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12848) );
  OAI22_X1 U16282 ( .A1(n13053), .A2(n12849), .B1(n12486), .B2(n12848), .ZN(
        n12850) );
  NOR2_X1 U16283 ( .A1(n12851), .A2(n12850), .ZN(n12855) );
  AOI22_X1 U16284 ( .A1(n13274), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n13245), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12854) );
  NAND2_X1 U16285 ( .A1(n13874), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n12853) );
  NAND2_X1 U16286 ( .A1(n13056), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n12852) );
  NAND4_X1 U16287 ( .A1(n12855), .A2(n12854), .A3(n12853), .A4(n12852), .ZN(
        n12856) );
  OAI21_X1 U16288 ( .B1(n12857), .B2(n12856), .A(n12930), .ZN(n12860) );
  NAND2_X1 U16289 ( .A1(n13232), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n12859) );
  NAND2_X1 U16290 ( .A1(n13303), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12858) );
  AND3_X1 U16291 ( .A1(n12860), .A2(n12859), .A3(n12858), .ZN(n12861) );
  NAND2_X1 U16292 ( .A1(n12862), .A2(n12861), .ZN(n15028) );
  NAND3_X1 U16293 ( .A1(n14992), .A2(n15013), .A3(n15028), .ZN(n12932) );
  OR2_X1 U16294 ( .A1(n12911), .A2(n15069), .ZN(n12863) );
  XNOR2_X1 U16295 ( .A(n12863), .B(n15049), .ZN(n15512) );
  NAND2_X1 U16296 ( .A1(n15512), .A2(n13267), .ZN(n12887) );
  INV_X1 U16297 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n22101) );
  NAND2_X1 U16298 ( .A1(n13061), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n12864) );
  OAI21_X1 U16299 ( .B1(n12865), .B2(n13250), .A(n12864), .ZN(n12869) );
  INV_X1 U16300 ( .A(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12866) );
  OAI22_X1 U16301 ( .A1(n13053), .A2(n12867), .B1(n12486), .B2(n12866), .ZN(
        n12868) );
  NOR2_X1 U16302 ( .A1(n12869), .A2(n12868), .ZN(n12873) );
  AOI22_X1 U16303 ( .A1(n13275), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13245), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12872) );
  NAND2_X1 U16304 ( .A1(n13874), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n12871) );
  NAND2_X1 U16305 ( .A1(n13056), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n12870) );
  NAND4_X1 U16306 ( .A1(n12873), .A2(n12872), .A3(n12871), .A4(n12870), .ZN(
        n12879) );
  AOI22_X1 U16307 ( .A1(n13129), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n13254), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12877) );
  AOI22_X1 U16308 ( .A1(n13255), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13274), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12876) );
  AOI22_X1 U16309 ( .A1(n12365), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n13256), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12875) );
  AOI22_X1 U16310 ( .A1(n13244), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12392), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12874) );
  NAND4_X1 U16311 ( .A1(n12877), .A2(n12876), .A3(n12875), .A4(n12874), .ZN(
        n12878) );
  NOR2_X1 U16312 ( .A1(n12879), .A2(n12878), .ZN(n12880) );
  OR2_X1 U16313 ( .A1(n12881), .A2(n12880), .ZN(n12883) );
  NAND2_X1 U16314 ( .A1(n13303), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n12882) );
  OAI211_X1 U16315 ( .C1(n12884), .C2(n22101), .A(n12883), .B(n12882), .ZN(
        n12885) );
  INV_X1 U16316 ( .A(n12885), .ZN(n12886) );
  NAND2_X1 U16317 ( .A1(n12887), .A2(n12886), .ZN(n15046) );
  XNOR2_X1 U16318 ( .A(n12911), .B(n15069), .ZN(n15524) );
  NAND2_X1 U16319 ( .A1(n15524), .A2(n13267), .ZN(n12906) );
  AOI22_X1 U16320 ( .A1(n13255), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n13245), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12891) );
  AOI22_X1 U16321 ( .A1(n12365), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12392), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12890) );
  AOI22_X1 U16322 ( .A1(n13129), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n13256), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12889) );
  AOI22_X1 U16323 ( .A1(n13254), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n13244), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12888) );
  NAND4_X1 U16324 ( .A1(n12891), .A2(n12890), .A3(n12889), .A4(n12888), .ZN(
        n12902) );
  NAND2_X1 U16325 ( .A1(n13061), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n12892) );
  OAI21_X1 U16326 ( .B1(n13194), .B2(n13250), .A(n12892), .ZN(n12896) );
  INV_X1 U16327 ( .A(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12894) );
  INV_X1 U16328 ( .A(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12893) );
  OAI22_X1 U16329 ( .A1(n13053), .A2(n12894), .B1(n12486), .B2(n12893), .ZN(
        n12895) );
  NOR2_X1 U16330 ( .A1(n12896), .A2(n12895), .ZN(n12900) );
  AOI22_X1 U16331 ( .A1(n13275), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n13274), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12899) );
  NAND2_X1 U16332 ( .A1(n13056), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n12898) );
  NAND2_X1 U16333 ( .A1(n13874), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n12897) );
  NAND4_X1 U16334 ( .A1(n12900), .A2(n12899), .A3(n12898), .A4(n12897), .ZN(
        n12901) );
  OAI21_X1 U16335 ( .B1(n12902), .B2(n12901), .A(n12930), .ZN(n12905) );
  NAND2_X1 U16336 ( .A1(n13232), .A2(P1_EAX_REG_12__SCAN_IN), .ZN(n12904) );
  NAND2_X1 U16337 ( .A1(n13303), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12903) );
  NAND2_X1 U16338 ( .A1(n12906), .A2(n10663), .ZN(n15044) );
  NAND2_X1 U16339 ( .A1(n15046), .A2(n15044), .ZN(n15009) );
  INV_X1 U16340 ( .A(n12907), .ZN(n12909) );
  INV_X1 U16341 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n12908) );
  NAND2_X1 U16342 ( .A1(n12909), .A2(n12908), .ZN(n12910) );
  NAND2_X1 U16343 ( .A1(n12911), .A2(n12910), .ZN(n15538) );
  NAND2_X1 U16344 ( .A1(n15538), .A2(n13267), .ZN(n12913) );
  AOI22_X1 U16345 ( .A1(n13232), .A2(P1_EAX_REG_11__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n13303), .ZN(n12912) );
  NAND2_X1 U16346 ( .A1(n12913), .A2(n12912), .ZN(n15007) );
  INV_X1 U16347 ( .A(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12982) );
  OAI22_X1 U16348 ( .A1(n13250), .A2(n12914), .B1(n13221), .B2(n12982), .ZN(
        n12918) );
  INV_X1 U16349 ( .A(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12916) );
  INV_X1 U16350 ( .A(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12915) );
  OAI22_X1 U16351 ( .A1(n13053), .A2(n12916), .B1(n12356), .B2(n12915), .ZN(
        n12917) );
  NOR2_X1 U16352 ( .A1(n12918), .A2(n12917), .ZN(n12922) );
  AOI22_X1 U16353 ( .A1(n13275), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13245), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12921) );
  NAND2_X1 U16354 ( .A1(n13056), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n12920) );
  NAND2_X1 U16355 ( .A1(n13874), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n12919) );
  NAND4_X1 U16356 ( .A1(n12922), .A2(n12921), .A3(n12920), .A4(n12919), .ZN(
        n12928) );
  AOI22_X1 U16357 ( .A1(n13255), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n13274), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12926) );
  AOI22_X1 U16358 ( .A1(n13061), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n13254), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12925) );
  AOI22_X1 U16359 ( .A1(n13129), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12392), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12924) );
  AOI22_X1 U16360 ( .A1(n13256), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n13244), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12923) );
  NAND4_X1 U16361 ( .A1(n12926), .A2(n12925), .A3(n12924), .A4(n12923), .ZN(
        n12927) );
  OR2_X1 U16362 ( .A1(n12928), .A2(n12927), .ZN(n12929) );
  NOR2_X1 U16363 ( .A1(n15007), .A2(n15077), .ZN(n12931) );
  INV_X1 U16364 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n12934) );
  XNOR2_X1 U16365 ( .A(n12954), .B(n12934), .ZN(n15473) );
  INV_X1 U16366 ( .A(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13122) );
  NAND2_X1 U16367 ( .A1(n13075), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n12935) );
  OAI21_X1 U16368 ( .B1(n13122), .B2(n13221), .A(n12935), .ZN(n12939) );
  INV_X1 U16369 ( .A(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12937) );
  OAI22_X1 U16370 ( .A1(n13053), .A2(n12937), .B1(n12486), .B2(n12936), .ZN(
        n12938) );
  NOR2_X1 U16371 ( .A1(n12939), .A2(n12938), .ZN(n12943) );
  AOI22_X1 U16372 ( .A1(n13275), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n13274), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12942) );
  NAND2_X1 U16373 ( .A1(n13056), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n12941) );
  NAND2_X1 U16374 ( .A1(n13874), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n12940) );
  NAND4_X1 U16375 ( .A1(n12943), .A2(n12942), .A3(n12941), .A4(n12940), .ZN(
        n12950) );
  AOI22_X1 U16376 ( .A1(n13279), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12944), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12948) );
  AOI22_X1 U16377 ( .A1(n13129), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n13254), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12947) );
  AOI22_X1 U16378 ( .A1(n13255), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n13256), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12946) );
  AOI22_X1 U16379 ( .A1(n13245), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n12392), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12945) );
  NAND4_X1 U16380 ( .A1(n12948), .A2(n12947), .A3(n12946), .A4(n12945), .ZN(
        n12949) );
  NOR2_X1 U16381 ( .A1(n12950), .A2(n12949), .ZN(n12952) );
  AOI22_X1 U16382 ( .A1(n12723), .A2(P1_EAX_REG_17__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n13303), .ZN(n12951) );
  OAI21_X1 U16383 ( .B1(n13299), .B2(n12952), .A(n12951), .ZN(n12953) );
  AOI21_X1 U16384 ( .B1(n15473), .B2(n13526), .A(n12953), .ZN(n14974) );
  INV_X1 U16385 ( .A(n12956), .ZN(n12958) );
  INV_X1 U16386 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n12957) );
  NAND2_X1 U16387 ( .A1(n12958), .A2(n12957), .ZN(n12959) );
  NAND2_X1 U16388 ( .A1(n13001), .A2(n12959), .ZN(n15459) );
  INV_X1 U16389 ( .A(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12961) );
  NAND2_X1 U16390 ( .A1(n13061), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n12960) );
  OAI21_X1 U16391 ( .B1(n12961), .B2(n13221), .A(n12960), .ZN(n12965) );
  INV_X1 U16392 ( .A(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12963) );
  OAI22_X1 U16393 ( .A1(n13053), .A2(n12963), .B1(n12356), .B2(n12962), .ZN(
        n12964) );
  NOR2_X1 U16394 ( .A1(n12965), .A2(n12964), .ZN(n12969) );
  AOI22_X1 U16395 ( .A1(n13275), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n13274), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12968) );
  NAND2_X1 U16396 ( .A1(n13056), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n12967) );
  NAND2_X1 U16397 ( .A1(n13874), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n12966) );
  NAND4_X1 U16398 ( .A1(n12969), .A2(n12968), .A3(n12967), .A4(n12966), .ZN(
        n12975) );
  AOI22_X1 U16399 ( .A1(n13279), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13129), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12973) );
  AOI22_X1 U16400 ( .A1(n13245), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n13254), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12972) );
  AOI22_X1 U16401 ( .A1(n13255), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n13256), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12971) );
  AOI22_X1 U16402 ( .A1(n13075), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12392), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12970) );
  NAND4_X1 U16403 ( .A1(n12973), .A2(n12972), .A3(n12971), .A4(n12970), .ZN(
        n12974) );
  NOR2_X1 U16404 ( .A1(n12975), .A2(n12974), .ZN(n12979) );
  NAND2_X1 U16405 ( .A1(n12682), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12976) );
  NAND2_X1 U16406 ( .A1(n13302), .A2(n12976), .ZN(n12977) );
  AOI21_X1 U16407 ( .B1(n13232), .B2(P1_EAX_REG_18__SCAN_IN), .A(n12977), .ZN(
        n12978) );
  OAI21_X1 U16408 ( .B1(n13299), .B2(n12979), .A(n12978), .ZN(n12980) );
  NAND2_X1 U16409 ( .A1(n12981), .A2(n12980), .ZN(n14963) );
  XNOR2_X1 U16410 ( .A(n13001), .B(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15456) );
  INV_X1 U16411 ( .A(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13176) );
  OAI22_X1 U16412 ( .A1(n13250), .A2(n12982), .B1(n13175), .B2(n13176), .ZN(
        n12986) );
  INV_X1 U16413 ( .A(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12984) );
  OAI22_X1 U16414 ( .A1(n13053), .A2(n12984), .B1(n12486), .B2(n12983), .ZN(
        n12985) );
  NOR2_X1 U16415 ( .A1(n12986), .A2(n12985), .ZN(n12990) );
  AOI22_X1 U16416 ( .A1(n13245), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12392), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12989) );
  NAND2_X1 U16417 ( .A1(n13056), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n12988) );
  NAND2_X1 U16418 ( .A1(n13874), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n12987) );
  NAND4_X1 U16419 ( .A1(n12990), .A2(n12989), .A3(n12988), .A4(n12987), .ZN(
        n12996) );
  AOI22_X1 U16420 ( .A1(n13129), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n13061), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12994) );
  AOI22_X1 U16421 ( .A1(n13275), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n13274), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12993) );
  AOI22_X1 U16422 ( .A1(n13255), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13254), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12992) );
  AOI22_X1 U16423 ( .A1(n13256), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n13244), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12991) );
  NAND4_X1 U16424 ( .A1(n12994), .A2(n12993), .A3(n12992), .A4(n12991), .ZN(
        n12995) );
  OR2_X1 U16425 ( .A1(n12996), .A2(n12995), .ZN(n12999) );
  INV_X1 U16426 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n15265) );
  NAND2_X1 U16427 ( .A1(n12682), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12997) );
  OAI211_X1 U16428 ( .C1(n12884), .C2(n15265), .A(n13302), .B(n12997), .ZN(
        n12998) );
  AOI21_X1 U16429 ( .B1(n13264), .B2(n12999), .A(n12998), .ZN(n13000) );
  AOI21_X1 U16430 ( .B1(n15456), .B2(n13267), .A(n13000), .ZN(n14943) );
  INV_X1 U16431 ( .A(n13002), .ZN(n13004) );
  INV_X1 U16432 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n13003) );
  NAND2_X1 U16433 ( .A1(n13004), .A2(n13003), .ZN(n13005) );
  NAND2_X1 U16434 ( .A1(n13047), .A2(n13005), .ZN(n15447) );
  NAND2_X1 U16435 ( .A1(n13129), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n13009) );
  NAND2_X1 U16436 ( .A1(n13061), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n13008) );
  NAND2_X1 U16437 ( .A1(n13240), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n13007) );
  NAND2_X1 U16438 ( .A1(n13155), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n13006) );
  AND4_X1 U16439 ( .A1(n13009), .A2(n13008), .A3(n13007), .A4(n13006), .ZN(
        n13013) );
  AOI22_X1 U16440 ( .A1(n13274), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n13256), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13012) );
  NAND2_X1 U16441 ( .A1(n13056), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n13011) );
  NAND2_X1 U16442 ( .A1(n13874), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n13010) );
  NAND4_X1 U16443 ( .A1(n13013), .A2(n13012), .A3(n13011), .A4(n13010), .ZN(
        n13022) );
  INV_X1 U16444 ( .A(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n13015) );
  INV_X1 U16445 ( .A(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13014) );
  OAI22_X1 U16446 ( .A1(n13250), .A2(n13015), .B1(n13221), .B2(n13014), .ZN(
        n13016) );
  INV_X1 U16447 ( .A(n13016), .ZN(n13020) );
  AOI22_X1 U16448 ( .A1(n13275), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12391), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13019) );
  AOI22_X1 U16449 ( .A1(n13255), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n13075), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13018) );
  AOI22_X1 U16450 ( .A1(n13254), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n13089), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13017) );
  NAND4_X1 U16451 ( .A1(n13020), .A2(n13019), .A3(n13018), .A4(n13017), .ZN(
        n13021) );
  NOR2_X1 U16452 ( .A1(n13022), .A2(n13021), .ZN(n13025) );
  OAI21_X1 U16453 ( .B1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n21905), .A(
        n12682), .ZN(n13024) );
  NAND2_X1 U16454 ( .A1(n12723), .A2(P1_EAX_REG_20__SCAN_IN), .ZN(n13023) );
  OAI211_X1 U16455 ( .C1(n13299), .C2(n13025), .A(n13024), .B(n13023), .ZN(
        n13026) );
  XNOR2_X1 U16456 ( .A(n13047), .B(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15434) );
  INV_X1 U16457 ( .A(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13028) );
  OAI22_X1 U16458 ( .A1(n13250), .A2(n13028), .B1(n13175), .B2(n21979), .ZN(
        n13032) );
  INV_X1 U16459 ( .A(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13030) );
  INV_X1 U16460 ( .A(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13029) );
  OAI22_X1 U16461 ( .A1(n13053), .A2(n13030), .B1(n12486), .B2(n13029), .ZN(
        n13031) );
  NOR2_X1 U16462 ( .A1(n13032), .A2(n13031), .ZN(n13036) );
  AOI22_X1 U16463 ( .A1(n13254), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n13089), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13035) );
  NAND2_X1 U16464 ( .A1(n13056), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n13034) );
  NAND2_X1 U16465 ( .A1(n13874), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n13033) );
  NAND4_X1 U16466 ( .A1(n13036), .A2(n13035), .A3(n13034), .A4(n13033), .ZN(
        n13042) );
  AOI22_X1 U16467 ( .A1(n13275), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13274), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13040) );
  AOI22_X1 U16468 ( .A1(n13061), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12391), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13039) );
  AOI22_X1 U16469 ( .A1(n13255), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13256), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13038) );
  AOI22_X1 U16470 ( .A1(n13129), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13244), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13037) );
  NAND4_X1 U16471 ( .A1(n13040), .A2(n13039), .A3(n13038), .A4(n13037), .ZN(
        n13041) );
  OR2_X1 U16472 ( .A1(n13042), .A2(n13041), .ZN(n13045) );
  INV_X1 U16473 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n15253) );
  NAND2_X1 U16474 ( .A1(n12682), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n13043) );
  OAI211_X1 U16475 ( .C1(n12884), .C2(n15253), .A(n13302), .B(n13043), .ZN(
        n13044) );
  AOI21_X1 U16476 ( .B1(n13264), .B2(n13045), .A(n13044), .ZN(n13046) );
  AOI21_X1 U16477 ( .B1(n15434), .B2(n13267), .A(n13046), .ZN(n14921) );
  NAND2_X1 U16478 ( .A1(n14919), .A2(n14921), .ZN(n14905) );
  NAND2_X1 U16479 ( .A1(n13048), .A2(n21959), .ZN(n13049) );
  NAND2_X1 U16480 ( .A1(n13113), .A2(n13049), .ZN(n15426) );
  INV_X1 U16481 ( .A(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n13050) );
  INV_X1 U16482 ( .A(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13249) );
  OAI22_X1 U16483 ( .A1(n13250), .A2(n13050), .B1(n13175), .B2(n13249), .ZN(
        n13055) );
  INV_X1 U16484 ( .A(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13052) );
  INV_X1 U16485 ( .A(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n13051) );
  OAI22_X1 U16486 ( .A1(n13053), .A2(n13052), .B1(n12356), .B2(n13051), .ZN(
        n13054) );
  NOR2_X1 U16487 ( .A1(n13055), .A2(n13054), .ZN(n13060) );
  AOI22_X1 U16488 ( .A1(n13255), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n13256), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13059) );
  NAND2_X1 U16489 ( .A1(n13056), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n13058) );
  NAND2_X1 U16490 ( .A1(n13874), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n13057) );
  NAND4_X1 U16491 ( .A1(n13060), .A2(n13059), .A3(n13058), .A4(n13057), .ZN(
        n13067) );
  AOI22_X1 U16492 ( .A1(n13275), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n13245), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13065) );
  AOI22_X1 U16493 ( .A1(n13061), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n13254), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13064) );
  AOI22_X1 U16494 ( .A1(n13274), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12392), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13063) );
  AOI22_X1 U16495 ( .A1(n13129), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13244), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13062) );
  NAND4_X1 U16496 ( .A1(n13065), .A2(n13064), .A3(n13063), .A4(n13062), .ZN(
        n13066) );
  NOR2_X1 U16497 ( .A1(n13067), .A2(n13066), .ZN(n13068) );
  NOR2_X1 U16498 ( .A1(n13299), .A2(n13068), .ZN(n13071) );
  INV_X1 U16499 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n15246) );
  NAND2_X1 U16500 ( .A1(n12682), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n13069) );
  OAI211_X1 U16501 ( .C1(n12884), .C2(n15246), .A(n13302), .B(n13069), .ZN(
        n13070) );
  OAI22_X1 U16502 ( .A1(n15426), .A2(n13302), .B1(n13071), .B2(n13070), .ZN(
        n14907) );
  XNOR2_X1 U16503 ( .A(n13113), .B(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15420) );
  INV_X1 U16504 ( .A(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13072) );
  OAI22_X1 U16505 ( .A1(n13053), .A2(n13072), .B1(n12486), .B2(n12142), .ZN(
        n13074) );
  INV_X1 U16506 ( .A(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13269) );
  NOR2_X1 U16507 ( .A1(n12342), .A2(n13269), .ZN(n13073) );
  AOI211_X1 U16508 ( .C1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .C2(n13129), .A(
        n13074), .B(n13073), .ZN(n13078) );
  AOI22_X1 U16509 ( .A1(n13279), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12365), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n13077) );
  AOI22_X1 U16510 ( .A1(n13061), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n13075), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13076) );
  NAND3_X1 U16511 ( .A1(n13078), .A2(n13077), .A3(n13076), .ZN(n13088) );
  AOI22_X1 U16512 ( .A1(n13255), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n13254), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13080) );
  OAI21_X1 U16513 ( .B1(n13082), .B2(n13081), .A(n13080), .ZN(n13083) );
  AOI21_X1 U16514 ( .B1(n13056), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A(
        n13083), .ZN(n13086) );
  AOI22_X1 U16515 ( .A1(n13274), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n13256), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13085) );
  AOI22_X1 U16516 ( .A1(n13275), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12392), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13084) );
  NAND3_X1 U16517 ( .A1(n13086), .A2(n13085), .A3(n13084), .ZN(n13087) );
  NOR2_X1 U16518 ( .A1(n13088), .A2(n13087), .ZN(n13118) );
  INV_X1 U16519 ( .A(n13089), .ZN(n13093) );
  AOI22_X1 U16520 ( .A1(n13061), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n13240), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13091) );
  NAND2_X1 U16521 ( .A1(n13874), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n13090) );
  OAI211_X1 U16522 ( .C1(n13093), .C2(n13092), .A(n13091), .B(n13090), .ZN(
        n13099) );
  OAI22_X1 U16523 ( .A1(n12335), .A2(n12272), .B1(n13094), .B2(n13250), .ZN(
        n13098) );
  INV_X1 U16524 ( .A(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13096) );
  INV_X1 U16525 ( .A(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13095) );
  OAI22_X1 U16526 ( .A1(n13096), .A2(n13133), .B1(n13282), .B2(n13095), .ZN(
        n13097) );
  OR3_X1 U16527 ( .A1(n13099), .A2(n13098), .A3(n13097), .ZN(n13108) );
  OAI22_X1 U16528 ( .A1(n13221), .A2(n13100), .B1(n12486), .B2(n12258), .ZN(
        n13103) );
  INV_X1 U16529 ( .A(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13101) );
  NOR2_X1 U16530 ( .A1(n12259), .A2(n13101), .ZN(n13102) );
  AOI211_X1 U16531 ( .C1(n13245), .C2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A(
        n13103), .B(n13102), .ZN(n13106) );
  AOI22_X1 U16532 ( .A1(n13129), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n13254), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13105) );
  AOI22_X1 U16533 ( .A1(n13255), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n13125), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13104) );
  NAND3_X1 U16534 ( .A1(n13106), .A2(n13105), .A3(n13104), .ZN(n13107) );
  NOR2_X1 U16535 ( .A1(n13108), .A2(n13107), .ZN(n13117) );
  XOR2_X1 U16536 ( .A(n13118), .B(n13117), .Z(n13111) );
  INV_X1 U16537 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n15240) );
  NOR2_X1 U16538 ( .A1(n21905), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n13109) );
  OAI22_X1 U16539 ( .A1(n12884), .A2(n15240), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n13109), .ZN(n13110) );
  AOI21_X1 U16540 ( .B1(n13111), .B2(n13264), .A(n13110), .ZN(n13112) );
  AOI21_X1 U16541 ( .B1(n15420), .B2(n13526), .A(n13112), .ZN(n14891) );
  INV_X1 U16542 ( .A(n13114), .ZN(n13115) );
  INV_X1 U16543 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n14882) );
  NAND2_X1 U16544 ( .A1(n13115), .A2(n14882), .ZN(n13116) );
  NAND2_X1 U16545 ( .A1(n13165), .A2(n13116), .ZN(n15410) );
  NOR2_X1 U16546 ( .A1(n13118), .A2(n13117), .ZN(n13146) );
  OAI22_X1 U16547 ( .A1(n13053), .A2(n13120), .B1(n12486), .B2(n13119), .ZN(
        n13124) );
  OAI22_X1 U16548 ( .A1(n13250), .A2(n13122), .B1(n13221), .B2(n13121), .ZN(
        n13123) );
  AOI211_X1 U16549 ( .C1(n13056), .C2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A(
        n13124), .B(n13123), .ZN(n13127) );
  AOI22_X1 U16550 ( .A1(n13125), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n13245), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13126) );
  OAI211_X1 U16551 ( .C1(n12342), .C2(n13128), .A(n13127), .B(n13126), .ZN(
        n13139) );
  AOI22_X1 U16552 ( .A1(n13255), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13129), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13131) );
  AOI22_X1 U16553 ( .A1(n13061), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n13244), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13130) );
  NAND2_X1 U16554 ( .A1(n13131), .A2(n13130), .ZN(n13138) );
  INV_X1 U16555 ( .A(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13132) );
  OAI22_X1 U16556 ( .A1(n13133), .A2(n13132), .B1(n13093), .B2(n12762), .ZN(
        n13137) );
  INV_X1 U16557 ( .A(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13134) );
  OAI22_X1 U16558 ( .A1(n12333), .A2(n13135), .B1(n13282), .B2(n13134), .ZN(
        n13136) );
  XNOR2_X1 U16559 ( .A(n13146), .B(n13145), .ZN(n13142) );
  OAI21_X1 U16560 ( .B1(n21905), .B2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n12682), .ZN(n13141) );
  NAND2_X1 U16561 ( .A1(n12723), .A2(P1_EAX_REG_24__SCAN_IN), .ZN(n13140) );
  OAI211_X1 U16562 ( .C1(n13142), .C2(n13299), .A(n13141), .B(n13140), .ZN(
        n13143) );
  OAI21_X1 U16563 ( .B1(n15410), .B2(n13302), .A(n13143), .ZN(n14880) );
  XNOR2_X1 U16564 ( .A(n13165), .B(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15401) );
  INV_X1 U16565 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n15399) );
  NOR2_X1 U16566 ( .A1(n15399), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13144) );
  AOI211_X1 U16567 ( .C1(n13232), .C2(P1_EAX_REG_25__SCAN_IN), .A(n13526), .B(
        n13144), .ZN(n13164) );
  NAND2_X1 U16568 ( .A1(n13146), .A2(n13145), .ZN(n13170) );
  OAI22_X1 U16569 ( .A1(n12332), .A2(n13148), .B1(n13093), .B2(n13147), .ZN(
        n13153) );
  AOI22_X1 U16570 ( .A1(n13129), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n13240), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13150) );
  AOI22_X1 U16571 ( .A1(n13254), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n13256), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13149) );
  OAI211_X1 U16572 ( .C1(n12342), .C2(n13151), .A(n13150), .B(n13149), .ZN(
        n13152) );
  AOI211_X1 U16573 ( .C1(n13056), .C2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A(
        n13153), .B(n13152), .ZN(n13154) );
  INV_X1 U16574 ( .A(n13154), .ZN(n13161) );
  AOI22_X1 U16575 ( .A1(n13279), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13061), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13159) );
  AOI22_X1 U16576 ( .A1(n13274), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n13245), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13158) );
  AOI22_X1 U16577 ( .A1(n12365), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n13155), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13157) );
  AOI22_X1 U16578 ( .A1(n13255), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13244), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13156) );
  NAND4_X1 U16579 ( .A1(n13159), .A2(n13158), .A3(n13157), .A4(n13156), .ZN(
        n13160) );
  NOR2_X1 U16580 ( .A1(n13161), .A2(n13160), .ZN(n13171) );
  XOR2_X1 U16581 ( .A(n13170), .B(n13171), .Z(n13162) );
  NAND2_X1 U16582 ( .A1(n13162), .A2(n13264), .ZN(n13163) );
  AOI22_X1 U16583 ( .A1(n15401), .A2(n13267), .B1(n13164), .B2(n13163), .ZN(
        n14867) );
  INV_X1 U16584 ( .A(n13165), .ZN(n13166) );
  INV_X1 U16585 ( .A(n13167), .ZN(n13168) );
  INV_X1 U16586 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n14854) );
  NAND2_X1 U16587 ( .A1(n13168), .A2(n14854), .ZN(n13169) );
  NAND2_X1 U16588 ( .A1(n13212), .A2(n13169), .ZN(n15395) );
  NOR2_X1 U16589 ( .A1(n13171), .A2(n13170), .ZN(n13192) );
  INV_X1 U16590 ( .A(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13173) );
  OAI22_X1 U16591 ( .A1(n13053), .A2(n13173), .B1(n12486), .B2(n13172), .ZN(
        n13178) );
  OAI22_X1 U16592 ( .A1(n13250), .A2(n13176), .B1(n13175), .B2(n13174), .ZN(
        n13177) );
  AOI211_X1 U16593 ( .C1(n13056), .C2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A(
        n13178), .B(n13177), .ZN(n13186) );
  AOI22_X1 U16594 ( .A1(n13255), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13129), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13182) );
  AOI22_X1 U16595 ( .A1(n13254), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n13256), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13181) );
  AOI22_X1 U16596 ( .A1(n13061), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n13244), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13180) );
  AOI22_X1 U16597 ( .A1(n13274), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12392), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13179) );
  AND4_X1 U16598 ( .A1(n13182), .A2(n13181), .A3(n13180), .A4(n13179), .ZN(
        n13185) );
  AOI22_X1 U16599 ( .A1(n13275), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12391), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13184) );
  NAND2_X1 U16600 ( .A1(n13874), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n13183) );
  NAND4_X1 U16601 ( .A1(n13186), .A2(n13185), .A3(n13184), .A4(n13183), .ZN(
        n13191) );
  XNOR2_X1 U16602 ( .A(n13192), .B(n13191), .ZN(n13189) );
  OAI21_X1 U16603 ( .B1(n21905), .B2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n12682), .ZN(n13188) );
  NAND2_X1 U16604 ( .A1(n12723), .A2(P1_EAX_REG_26__SCAN_IN), .ZN(n13187) );
  OAI211_X1 U16605 ( .C1(n13189), .C2(n13299), .A(n13188), .B(n13187), .ZN(
        n13190) );
  OAI21_X1 U16606 ( .B1(n15395), .B2(n13302), .A(n13190), .ZN(n14852) );
  NOR2_X2 U16607 ( .A1(n14850), .A2(n14852), .ZN(n14833) );
  XNOR2_X1 U16608 ( .A(n13212), .B(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15380) );
  NAND2_X1 U16609 ( .A1(n13192), .A2(n13191), .ZN(n13217) );
  INV_X1 U16610 ( .A(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13193) );
  OAI22_X1 U16611 ( .A1(n13053), .A2(n13193), .B1(n12486), .B2(n12162), .ZN(
        n13196) );
  NOR2_X1 U16612 ( .A1(n12342), .A2(n13194), .ZN(n13195) );
  AOI211_X1 U16613 ( .C1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .C2(n13245), .A(
        n13196), .B(n13195), .ZN(n13199) );
  AOI22_X1 U16614 ( .A1(n13274), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n13244), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13198) );
  AOI22_X1 U16615 ( .A1(n13275), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n13256), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13197) );
  NAND3_X1 U16616 ( .A1(n13199), .A2(n13198), .A3(n13197), .ZN(n13207) );
  INV_X1 U16617 ( .A(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13201) );
  AOI22_X1 U16618 ( .A1(n13279), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12365), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13200) );
  OAI21_X1 U16619 ( .B1(n12333), .B2(n13201), .A(n13200), .ZN(n13202) );
  AOI21_X1 U16620 ( .B1(n13056), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A(
        n13202), .ZN(n13205) );
  AOI22_X1 U16621 ( .A1(n13129), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n13061), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n13204) );
  AOI22_X1 U16622 ( .A1(n13255), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12392), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13203) );
  NAND3_X1 U16623 ( .A1(n13205), .A2(n13204), .A3(n13203), .ZN(n13206) );
  NOR2_X1 U16624 ( .A1(n13207), .A2(n13206), .ZN(n13218) );
  XOR2_X1 U16625 ( .A(n13217), .B(n13218), .Z(n13210) );
  INV_X1 U16626 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n15217) );
  NOR2_X1 U16627 ( .A1(n21905), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n13208) );
  OAI22_X1 U16628 ( .A1(n12884), .A2(n15217), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n13208), .ZN(n13209) );
  AOI21_X1 U16629 ( .B1(n13210), .B2(n13264), .A(n13209), .ZN(n13211) );
  AOI21_X1 U16630 ( .B1(n15380), .B2(n13267), .A(n13211), .ZN(n14834) );
  NAND2_X1 U16631 ( .A1(n14833), .A2(n14834), .ZN(n14821) );
  INV_X1 U16632 ( .A(n13212), .ZN(n13213) );
  NAND2_X1 U16633 ( .A1(n13213), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n13215) );
  INV_X1 U16634 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n13214) );
  NAND2_X1 U16635 ( .A1(n13215), .A2(n13214), .ZN(n13216) );
  NAND2_X1 U16636 ( .A1(n13237), .A2(n13216), .ZN(n15376) );
  NOR2_X1 U16637 ( .A1(n13218), .A2(n13217), .ZN(n13239) );
  INV_X1 U16638 ( .A(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13219) );
  OAI22_X1 U16639 ( .A1(n13053), .A2(n13219), .B1(n12486), .B2(n12116), .ZN(
        n13223) );
  INV_X1 U16640 ( .A(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13220) );
  OAI22_X1 U16641 ( .A1(n21979), .A2(n13250), .B1(n13221), .B2(n13220), .ZN(
        n13222) );
  AOI211_X1 U16642 ( .C1(n13056), .C2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A(
        n13223), .B(n13222), .ZN(n13231) );
  AOI22_X1 U16643 ( .A1(n13255), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n13129), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13227) );
  AOI22_X1 U16644 ( .A1(n13254), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n13256), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13226) );
  AOI22_X1 U16645 ( .A1(n13061), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13244), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13225) );
  AOI22_X1 U16646 ( .A1(n13274), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12392), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13224) );
  AND4_X1 U16647 ( .A1(n13227), .A2(n13226), .A3(n13225), .A4(n13224), .ZN(
        n13230) );
  AOI22_X1 U16648 ( .A1(n13275), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12391), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13229) );
  NAND2_X1 U16649 ( .A1(n13874), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n13228) );
  NAND4_X1 U16650 ( .A1(n13231), .A2(n13230), .A3(n13229), .A4(n13228), .ZN(
        n13238) );
  XNOR2_X1 U16651 ( .A(n13239), .B(n13238), .ZN(n13235) );
  AOI21_X1 U16652 ( .B1(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n12682), .A(
        n13526), .ZN(n13234) );
  NAND2_X1 U16653 ( .A1(n13232), .A2(P1_EAX_REG_28__SCAN_IN), .ZN(n13233) );
  OAI211_X1 U16654 ( .C1(n13235), .C2(n13299), .A(n13234), .B(n13233), .ZN(
        n13236) );
  OAI21_X1 U16655 ( .B1(n15376), .B2(n13302), .A(n13236), .ZN(n14823) );
  XOR2_X1 U16656 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B(n13268), .Z(
        n15364) );
  NAND2_X1 U16657 ( .A1(n13239), .A2(n13238), .ZN(n13293) );
  INV_X1 U16658 ( .A(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13242) );
  AOI22_X1 U16659 ( .A1(n13061), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13240), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13241) );
  OAI21_X1 U16660 ( .B1(n13133), .B2(n13242), .A(n13241), .ZN(n13243) );
  AOI21_X1 U16661 ( .B1(n13874), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A(
        n13243), .ZN(n13248) );
  AOI22_X1 U16662 ( .A1(n12365), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n13244), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13247) );
  AOI22_X1 U16663 ( .A1(n13129), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n13245), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13246) );
  NAND3_X1 U16664 ( .A1(n13248), .A2(n13247), .A3(n13246), .ZN(n13261) );
  OAI22_X1 U16665 ( .A1(n13250), .A2(n13249), .B1(n12486), .B2(n12192), .ZN(
        n13253) );
  INV_X1 U16666 ( .A(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13251) );
  NOR2_X1 U16667 ( .A1(n12259), .A2(n13251), .ZN(n13252) );
  AOI211_X1 U16668 ( .C1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .C2(n13089), .A(
        n13253), .B(n13252), .ZN(n13259) );
  AOI22_X1 U16669 ( .A1(n13255), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13254), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13258) );
  AOI22_X1 U16670 ( .A1(n13275), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n13256), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13257) );
  NAND3_X1 U16671 ( .A1(n13259), .A2(n13258), .A3(n13257), .ZN(n13260) );
  NOR2_X1 U16672 ( .A1(n13261), .A2(n13260), .ZN(n13294) );
  XOR2_X1 U16673 ( .A(n13293), .B(n13294), .Z(n13265) );
  INV_X1 U16674 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n15205) );
  NOR2_X1 U16675 ( .A1(n21905), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13262) );
  OAI22_X1 U16676 ( .A1(n12884), .A2(n15205), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n13262), .ZN(n13263) );
  AOI21_X1 U16677 ( .B1(n13265), .B2(n13264), .A(n13263), .ZN(n13266) );
  INV_X1 U16678 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n13306) );
  INV_X1 U16679 ( .A(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13270) );
  OAI22_X1 U16680 ( .A1(n13053), .A2(n13270), .B1(n12486), .B2(n13269), .ZN(
        n13273) );
  INV_X1 U16681 ( .A(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n13271) );
  NOR2_X1 U16682 ( .A1(n12342), .A2(n13271), .ZN(n13272) );
  AOI211_X1 U16683 ( .C1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .C2(n12391), .A(
        n13273), .B(n13272), .ZN(n13278) );
  AOI22_X1 U16684 ( .A1(n12365), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n13274), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13277) );
  AOI22_X1 U16685 ( .A1(n13275), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n13089), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13276) );
  NAND3_X1 U16686 ( .A1(n13278), .A2(n13277), .A3(n13276), .ZN(n13292) );
  INV_X1 U16687 ( .A(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13283) );
  AOI22_X1 U16688 ( .A1(n13279), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13061), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13281) );
  NAND2_X1 U16689 ( .A1(n13056), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n13280) );
  OAI211_X1 U16690 ( .C1(n13283), .C2(n13282), .A(n13281), .B(n13280), .ZN(
        n13290) );
  OAI22_X1 U16691 ( .A1(n13285), .A2(n12142), .B1(n12335), .B2(n13284), .ZN(
        n13289) );
  INV_X1 U16692 ( .A(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13286) );
  OAI22_X1 U16693 ( .A1(n12334), .A2(n13287), .B1(n12333), .B2(n13286), .ZN(
        n13288) );
  OR3_X1 U16694 ( .A1(n13290), .A2(n13289), .A3(n13288), .ZN(n13291) );
  NOR2_X1 U16695 ( .A1(n13292), .A2(n13291), .ZN(n13296) );
  NOR2_X1 U16696 ( .A1(n13294), .A2(n13293), .ZN(n13295) );
  XOR2_X1 U16697 ( .A(n13296), .B(n13295), .Z(n13300) );
  AOI21_X1 U16698 ( .B1(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n12682), .A(
        n13526), .ZN(n13298) );
  NAND2_X1 U16699 ( .A1(n12723), .A2(P1_EAX_REG_30__SCAN_IN), .ZN(n13297) );
  OAI211_X1 U16700 ( .C1(n13300), .C2(n13299), .A(n13298), .B(n13297), .ZN(
        n13301) );
  OAI21_X1 U16701 ( .B1(n15361), .B2(n13302), .A(n13301), .ZN(n14789) );
  AOI22_X1 U16702 ( .A1(n12723), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n13303), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n13304) );
  NAND3_X1 U16703 ( .A1(n21908), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n17708) );
  INV_X1 U16704 ( .A(n17708), .ZN(n13305) );
  OR2_X2 U16705 ( .A1(n13307), .A2(n13306), .ZN(n13308) );
  INV_X1 U16706 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n13542) );
  XNOR2_X2 U16707 ( .A(n13308), .B(n13542), .ZN(n14799) );
  NAND2_X1 U16708 ( .A1(n21810), .A2(n13312), .ZN(n21911) );
  NAND2_X1 U16709 ( .A1(n21911), .A2(n21908), .ZN(n13309) );
  NAND2_X1 U16710 ( .A1(n21908), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13311) );
  NAND2_X1 U16711 ( .A1(n21905), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13310) );
  NAND2_X1 U16712 ( .A1(n13311), .A2(n13310), .ZN(n13841) );
  INV_X1 U16713 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n22154) );
  NOR2_X1 U16714 ( .A1(n15837), .A2(n22154), .ZN(n13381) );
  AOI21_X1 U16715 ( .B1(n17661), .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n13381), .ZN(n13313) );
  OAI21_X1 U16716 ( .B1(n14799), .B2(n17670), .A(n13313), .ZN(n13314) );
  AOI21_X1 U16717 ( .B1(n14747), .B2(n21328), .A(n13314), .ZN(n13315) );
  NOR3_X1 U16718 ( .A1(n13318), .A2(n13317), .A3(n13316), .ZN(n13320) );
  OAI21_X1 U16719 ( .B1(n13321), .B2(n13320), .A(n13319), .ZN(n14779) );
  AOI21_X1 U16720 ( .B1(n15303), .B2(n15925), .A(n17713), .ZN(n13323) );
  NAND2_X1 U16721 ( .A1(n14779), .A2(n13323), .ZN(n13329) );
  NAND2_X1 U16722 ( .A1(n12289), .A2(n15925), .ZN(n13531) );
  AND2_X1 U16723 ( .A1(n13531), .A2(n21912), .ZN(n13326) );
  NAND2_X1 U16724 ( .A1(n13860), .A2(n12288), .ZN(n13325) );
  AOI21_X1 U16725 ( .B1(n13324), .B2(n13326), .A(n13325), .ZN(n13327) );
  MUX2_X1 U16726 ( .A(n13329), .B(n13328), .S(n13350), .Z(n13336) );
  INV_X1 U16727 ( .A(n13347), .ZN(n13334) );
  INV_X1 U16728 ( .A(n13338), .ZN(n13333) );
  OAI21_X1 U16729 ( .B1(n12320), .B2(n21334), .A(n15300), .ZN(n13330) );
  NAND2_X1 U16730 ( .A1(n13331), .A2(n13330), .ZN(n13353) );
  AOI21_X1 U16731 ( .B1(n13333), .B2(n13353), .A(n14777), .ZN(n13887) );
  AOI21_X1 U16732 ( .B1(n17629), .B2(n13334), .A(n13887), .ZN(n13335) );
  NAND2_X1 U16733 ( .A1(n13336), .A2(n13335), .ZN(n13337) );
  NAND2_X1 U16734 ( .A1(n13885), .A2(n13339), .ZN(n14774) );
  OAI21_X1 U16735 ( .B1(n13489), .B2(n12296), .A(n13340), .ZN(n13341) );
  NOR2_X1 U16736 ( .A1(n14774), .A2(n13341), .ZN(n13342) );
  OAI21_X1 U16737 ( .B1(n13344), .B2(n15094), .A(n13343), .ZN(n13345) );
  INV_X1 U16738 ( .A(n15851), .ZN(n15771) );
  INV_X1 U16739 ( .A(n15091), .ZN(n13741) );
  NAND2_X1 U16740 ( .A1(n12319), .A2(n13741), .ZN(n13356) );
  INV_X1 U16741 ( .A(n13348), .ZN(n13355) );
  OAI211_X1 U16742 ( .C1(n13350), .C2(n13852), .A(n12313), .B(n12672), .ZN(
        n13351) );
  AOI22_X1 U16743 ( .A1(n13352), .A2(n13740), .B1(n15303), .B2(n13351), .ZN(
        n13354) );
  NAND4_X1 U16744 ( .A1(n13356), .A2(n13355), .A3(n13354), .A4(n13353), .ZN(
        n13869) );
  INV_X1 U16745 ( .A(n13869), .ZN(n13358) );
  OAI211_X1 U16746 ( .C1(n13866), .C2(n12288), .A(n13358), .B(n13357), .ZN(
        n13359) );
  NAND2_X1 U16747 ( .A1(n14777), .A2(n15303), .ZN(n15908) );
  NAND3_X1 U16748 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n15818) );
  NAND2_X1 U16749 ( .A1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n13360) );
  NOR2_X1 U16750 ( .A1(n15818), .A2(n13360), .ZN(n15808) );
  AND2_X1 U16751 ( .A1(n15808), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n15799) );
  AND2_X1 U16752 ( .A1(n15799), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15678) );
  NAND2_X1 U16753 ( .A1(n15678), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15757) );
  NAND2_X1 U16754 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n15854) );
  INV_X1 U16755 ( .A(n15854), .ZN(n13361) );
  NAND3_X1 U16756 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n13361), .ZN(n15843) );
  NOR2_X1 U16757 ( .A1(n15756), .A2(n15843), .ZN(n15788) );
  INV_X1 U16758 ( .A(n15788), .ZN(n13362) );
  NOR2_X1 U16759 ( .A1(n15757), .A2(n13362), .ZN(n13375) );
  INV_X1 U16760 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n15679) );
  OAI21_X1 U16761 ( .B1(n15679), .B2(n15751), .A(n15752), .ZN(n15754) );
  INV_X1 U16762 ( .A(n15754), .ZN(n15850) );
  NOR2_X1 U16763 ( .A1(n15850), .A2(n15854), .ZN(n13363) );
  NAND2_X1 U16764 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n13363), .ZN(
        n15817) );
  NAND2_X1 U16765 ( .A1(n15851), .A2(n15817), .ZN(n13365) );
  NAND2_X1 U16766 ( .A1(n15851), .A2(n15757), .ZN(n13366) );
  OAI211_X1 U16767 ( .C1(n15816), .C2(n13375), .A(n15840), .B(n13366), .ZN(
        n15750) );
  NAND2_X1 U16768 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15731) );
  NAND2_X1 U16769 ( .A1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n13367) );
  NOR2_X1 U16770 ( .A1(n15731), .A2(n13367), .ZN(n15703) );
  NAND2_X1 U16771 ( .A1(n15703), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n13368) );
  AND2_X1 U16772 ( .A1(n17681), .A2(n13368), .ZN(n13369) );
  NOR2_X1 U16773 ( .A1(n15750), .A2(n13369), .ZN(n15694) );
  NAND2_X1 U16774 ( .A1(n17681), .A2(n15647), .ZN(n13370) );
  NAND2_X1 U16775 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15659) );
  NAND2_X1 U16776 ( .A1(n17681), .A2(n15659), .ZN(n13371) );
  NAND2_X1 U16777 ( .A1(n15851), .A2(n15650), .ZN(n13372) );
  NAND2_X1 U16778 ( .A1(n13373), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15618) );
  AND2_X1 U16779 ( .A1(n17681), .A2(n15618), .ZN(n13374) );
  INV_X1 U16780 ( .A(n15670), .ZN(n15658) );
  NOR2_X1 U16781 ( .A1(n15658), .A2(n17681), .ZN(n15608) );
  AOI21_X1 U16782 ( .B1(n15616), .B2(n13379), .A(n15608), .ZN(n15595) );
  NOR3_X1 U16783 ( .A1(n15587), .A2(n15608), .A3(n12611), .ZN(n13382) );
  INV_X1 U16784 ( .A(n15816), .ZN(n15842) );
  NAND2_X1 U16785 ( .A1(n15682), .A2(n15679), .ZN(n13916) );
  NAND2_X1 U16786 ( .A1(n15842), .A2(n13916), .ZN(n15793) );
  INV_X1 U16787 ( .A(n13375), .ZN(n15768) );
  INV_X1 U16788 ( .A(n15817), .ZN(n13376) );
  AND2_X1 U16789 ( .A1(n15678), .A2(n13376), .ZN(n15772) );
  AND2_X1 U16790 ( .A1(n15851), .A2(n15772), .ZN(n15680) );
  NAND2_X1 U16791 ( .A1(n15680), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n13377) );
  NAND2_X1 U16792 ( .A1(n15637), .A2(n13377), .ZN(n15714) );
  NAND2_X1 U16793 ( .A1(n15706), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15695) );
  NOR2_X1 U16794 ( .A1(n15695), .A2(n15647), .ZN(n15673) );
  INV_X1 U16795 ( .A(n15659), .ZN(n13378) );
  NAND2_X1 U16796 ( .A1(n15673), .A2(n13378), .ZN(n15638) );
  NOR2_X1 U16797 ( .A1(n15638), .A2(n15384), .ZN(n15612) );
  NAND2_X1 U16798 ( .A1(n15612), .A2(n13379), .ZN(n15592) );
  NOR4_X1 U16799 ( .A1(n15592), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n15367), .A4(n15357), .ZN(n13380) );
  NOR3_X1 U16800 ( .A1(n13382), .A2(n13381), .A3(n13380), .ZN(n13494) );
  INV_X1 U16801 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n13388) );
  NAND2_X1 U16802 ( .A1(n13937), .A2(n13388), .ZN(n13387) );
  NAND2_X1 U16803 ( .A1(n9713), .A2(n15751), .ZN(n13386) );
  NAND3_X1 U16804 ( .A1(n13387), .A2(n14793), .A3(n13386), .ZN(n13390) );
  NAND2_X1 U16805 ( .A1(n13740), .A2(n13388), .ZN(n13389) );
  NAND2_X1 U16806 ( .A1(n13390), .A2(n13389), .ZN(n13392) );
  NAND2_X1 U16807 ( .A1(n9713), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n13391) );
  OAI21_X1 U16808 ( .B1(n13740), .B2(P1_EBX_REG_0__SCAN_IN), .A(n13391), .ZN(
        n13831) );
  XNOR2_X1 U16809 ( .A(n13392), .B(n13831), .ZN(n13911) );
  NAND2_X1 U16810 ( .A1(n13911), .A2(n13937), .ZN(n13913) );
  INV_X1 U16811 ( .A(n13392), .ZN(n13393) );
  NAND2_X1 U16812 ( .A1(n13393), .A2(n13831), .ZN(n13394) );
  NAND2_X1 U16813 ( .A1(n13913), .A2(n13394), .ZN(n14075) );
  NAND2_X1 U16814 ( .A1(n9713), .A2(n15752), .ZN(n13396) );
  INV_X1 U16815 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n13397) );
  NAND2_X1 U16816 ( .A1(n13937), .A2(n13397), .ZN(n13395) );
  NAND3_X1 U16817 ( .A1(n14793), .A2(n13396), .A3(n13395), .ZN(n13399) );
  NAND2_X1 U16818 ( .A1(n13740), .A2(n13397), .ZN(n13398) );
  AND2_X1 U16819 ( .A1(n13399), .A2(n13398), .ZN(n14074) );
  MUX2_X1 U16820 ( .A(n13471), .B(n14793), .S(P1_EBX_REG_3__SCAN_IN), .Z(
        n13402) );
  OR2_X1 U16821 ( .A1(n13485), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13401) );
  AND2_X1 U16822 ( .A1(n13402), .A2(n13401), .ZN(n15190) );
  NAND2_X1 U16823 ( .A1(n14073), .A2(n15190), .ZN(n15170) );
  INV_X1 U16824 ( .A(n9713), .ZN(n13452) );
  MUX2_X1 U16825 ( .A(n13740), .B(n13452), .S(P1_EBX_REG_4__SCAN_IN), .Z(
        n13405) );
  NAND2_X1 U16826 ( .A1(n13452), .A2(n14786), .ZN(n13415) );
  NAND2_X1 U16827 ( .A1(n14786), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13403) );
  NAND2_X1 U16828 ( .A1(n13415), .A2(n13403), .ZN(n13404) );
  NOR2_X1 U16829 ( .A1(n13405), .A2(n13404), .ZN(n15184) );
  INV_X1 U16830 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n13406) );
  NAND2_X1 U16831 ( .A1(n13937), .A2(n13406), .ZN(n13407) );
  OAI211_X1 U16832 ( .C1(n13740), .C2(n15756), .A(n13407), .B(n9713), .ZN(
        n13408) );
  OAI21_X1 U16833 ( .B1(n13471), .B2(P1_EBX_REG_5__SCAN_IN), .A(n13408), .ZN(
        n15171) );
  INV_X1 U16834 ( .A(n13471), .ZN(n13465) );
  INV_X1 U16835 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n21195) );
  NAND2_X1 U16836 ( .A1(n13465), .A2(n21195), .ZN(n13413) );
  INV_X1 U16837 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n13411) );
  NAND2_X1 U16838 ( .A1(n13937), .A2(n21195), .ZN(n13410) );
  OAI211_X1 U16839 ( .C1(n13740), .C2(n13411), .A(n13410), .B(n9713), .ZN(
        n13412) );
  AND2_X1 U16840 ( .A1(n13413), .A2(n13412), .ZN(n15159) );
  MUX2_X1 U16841 ( .A(n14793), .B(n9713), .S(P1_EBX_REG_6__SCAN_IN), .Z(n13417) );
  NAND2_X1 U16842 ( .A1(n14786), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13414) );
  AND2_X1 U16843 ( .A1(n13415), .A2(n13414), .ZN(n13416) );
  NAND2_X1 U16844 ( .A1(n13417), .A2(n13416), .ZN(n15165) );
  INV_X1 U16845 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n13418) );
  NAND2_X1 U16846 ( .A1(n13465), .A2(n13418), .ZN(n13422) );
  INV_X1 U16847 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n13420) );
  NAND2_X1 U16848 ( .A1(n13937), .A2(n13418), .ZN(n13419) );
  OAI211_X1 U16849 ( .C1(n13740), .C2(n13420), .A(n13419), .B(n9713), .ZN(
        n13421) );
  AND2_X1 U16850 ( .A1(n13422), .A2(n13421), .ZN(n15151) );
  MUX2_X1 U16851 ( .A(n14793), .B(n9713), .S(P1_EBX_REG_8__SCAN_IN), .Z(n13424) );
  NAND2_X1 U16852 ( .A1(n14786), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13423) );
  NAND2_X1 U16853 ( .A1(n13424), .A2(n13423), .ZN(n15154) );
  NAND2_X1 U16854 ( .A1(n9713), .A2(n15534), .ZN(n13426) );
  INV_X1 U16855 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n17645) );
  NAND2_X1 U16856 ( .A1(n13937), .A2(n17645), .ZN(n13425) );
  NAND3_X1 U16857 ( .A1(n14793), .A2(n13426), .A3(n13425), .ZN(n13428) );
  NAND2_X1 U16858 ( .A1(n13740), .A2(n17645), .ZN(n13427) );
  NAND2_X1 U16859 ( .A1(n13428), .A2(n13427), .ZN(n15142) );
  MUX2_X1 U16860 ( .A(n13471), .B(n14793), .S(P1_EBX_REG_11__SCAN_IN), .Z(
        n13429) );
  OAI21_X1 U16861 ( .B1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n13485), .A(
        n13429), .ZN(n15082) );
  MUX2_X1 U16862 ( .A(n13740), .B(n13452), .S(P1_EBX_REG_12__SCAN_IN), .Z(
        n13433) );
  NOR2_X1 U16863 ( .A1(n13937), .A2(n15798), .ZN(n13432) );
  NOR2_X1 U16864 ( .A1(n13433), .A2(n13432), .ZN(n15064) );
  MUX2_X1 U16865 ( .A(n13471), .B(n14793), .S(P1_EBX_REG_13__SCAN_IN), .Z(
        n13435) );
  OR2_X1 U16866 ( .A1(n13485), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n13434) );
  NAND2_X1 U16867 ( .A1(n9713), .A2(n15758), .ZN(n13437) );
  INV_X1 U16868 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n15135) );
  NAND2_X1 U16869 ( .A1(n13937), .A2(n15135), .ZN(n13436) );
  NAND3_X1 U16870 ( .A1(n14793), .A2(n13437), .A3(n13436), .ZN(n13439) );
  NAND2_X1 U16871 ( .A1(n13740), .A2(n15135), .ZN(n13438) );
  NAND2_X1 U16872 ( .A1(n13439), .A2(n13438), .ZN(n15030) );
  MUX2_X1 U16873 ( .A(n13471), .B(n14793), .S(P1_EBX_REG_15__SCAN_IN), .Z(
        n13440) );
  OAI21_X1 U16874 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n13485), .A(
        n13440), .ZN(n15015) );
  INV_X1 U16875 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15466) );
  NAND2_X1 U16876 ( .A1(n9713), .A2(n15466), .ZN(n13442) );
  INV_X1 U16877 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n15133) );
  NAND2_X1 U16878 ( .A1(n13937), .A2(n15133), .ZN(n13441) );
  NAND3_X1 U16879 ( .A1(n14793), .A2(n13442), .A3(n13441), .ZN(n13444) );
  NAND2_X1 U16880 ( .A1(n13740), .A2(n15133), .ZN(n13443) );
  NOR2_X4 U16881 ( .A1(n15017), .A2(n14995), .ZN(n14994) );
  MUX2_X1 U16882 ( .A(n13471), .B(n14793), .S(P1_EBX_REG_17__SCAN_IN), .Z(
        n13446) );
  OR2_X1 U16883 ( .A1(n13485), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n13445) );
  INV_X1 U16884 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15708) );
  NAND2_X1 U16885 ( .A1(n9713), .A2(n15708), .ZN(n13448) );
  INV_X1 U16886 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n15132) );
  NAND2_X1 U16887 ( .A1(n13937), .A2(n15132), .ZN(n13447) );
  NAND3_X1 U16888 ( .A1(n14793), .A2(n13448), .A3(n13447), .ZN(n13450) );
  NAND2_X1 U16889 ( .A1(n13740), .A2(n15132), .ZN(n13449) );
  NAND2_X1 U16890 ( .A1(n13450), .A2(n13449), .ZN(n14960) );
  MUX2_X1 U16891 ( .A(n13471), .B(n14793), .S(P1_EBX_REG_19__SCAN_IN), .Z(
        n13451) );
  OAI21_X1 U16892 ( .B1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n13485), .A(
        n13451), .ZN(n14945) );
  MUX2_X1 U16893 ( .A(n13740), .B(n13452), .S(P1_EBX_REG_20__SCAN_IN), .Z(
        n13454) );
  INV_X1 U16894 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15677) );
  NOR2_X1 U16895 ( .A1(n13937), .A2(n15677), .ZN(n13453) );
  NOR2_X1 U16896 ( .A1(n13454), .A2(n13453), .ZN(n14935) );
  MUX2_X1 U16897 ( .A(n13471), .B(n14793), .S(P1_EBX_REG_21__SCAN_IN), .Z(
        n13455) );
  OAI21_X1 U16898 ( .B1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n13485), .A(
        n13455), .ZN(n14926) );
  INV_X1 U16899 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15424) );
  NAND2_X1 U16900 ( .A1(n9713), .A2(n15424), .ZN(n13457) );
  INV_X1 U16901 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n15126) );
  NAND2_X1 U16902 ( .A1(n13937), .A2(n15126), .ZN(n13456) );
  NAND3_X1 U16903 ( .A1(n14793), .A2(n13457), .A3(n13456), .ZN(n13459) );
  NAND2_X1 U16904 ( .A1(n13740), .A2(n15126), .ZN(n13458) );
  NAND2_X1 U16905 ( .A1(n13459), .A2(n13458), .ZN(n14902) );
  NAND2_X1 U16906 ( .A1(n14928), .A2(n14902), .ZN(n14904) );
  MUX2_X1 U16907 ( .A(n13471), .B(n14793), .S(P1_EBX_REG_23__SCAN_IN), .Z(
        n13460) );
  OAI21_X1 U16908 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n13485), .A(
        n13460), .ZN(n14897) );
  INV_X1 U16909 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15403) );
  NAND2_X1 U16910 ( .A1(n9713), .A2(n15403), .ZN(n13462) );
  INV_X1 U16911 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n14883) );
  NAND2_X1 U16912 ( .A1(n13937), .A2(n14883), .ZN(n13461) );
  NAND3_X1 U16913 ( .A1(n14793), .A2(n13462), .A3(n13461), .ZN(n13464) );
  NAND2_X1 U16914 ( .A1(n13740), .A2(n14883), .ZN(n13463) );
  INV_X1 U16915 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n22121) );
  NAND2_X1 U16916 ( .A1(n13465), .A2(n22121), .ZN(n13468) );
  INV_X1 U16917 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15627) );
  NAND2_X1 U16918 ( .A1(n13937), .A2(n22121), .ZN(n13466) );
  OAI211_X1 U16919 ( .C1(n13740), .C2(n15627), .A(n13466), .B(n9713), .ZN(
        n13467) );
  MUX2_X1 U16920 ( .A(n14793), .B(n9713), .S(P1_EBX_REG_26__SCAN_IN), .Z(
        n13470) );
  NAND2_X1 U16921 ( .A1(n14786), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n13469) );
  NAND2_X1 U16922 ( .A1(n13470), .A2(n13469), .ZN(n14848) );
  NAND2_X1 U16923 ( .A1(n14847), .A2(n14848), .ZN(n14840) );
  MUX2_X1 U16924 ( .A(n13471), .B(n14793), .S(P1_EBX_REG_27__SCAN_IN), .Z(
        n13472) );
  OAI21_X1 U16925 ( .B1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n13485), .A(
        n13472), .ZN(n14841) );
  INV_X1 U16926 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15599) );
  NAND2_X1 U16927 ( .A1(n9713), .A2(n15599), .ZN(n13474) );
  INV_X1 U16928 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n13475) );
  NAND2_X1 U16929 ( .A1(n13937), .A2(n13475), .ZN(n13473) );
  NAND3_X1 U16930 ( .A1(n14793), .A2(n13474), .A3(n13473), .ZN(n13477) );
  NAND2_X1 U16931 ( .A1(n13740), .A2(n13475), .ZN(n13476) );
  OR2_X1 U16932 ( .A1(n13485), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13479) );
  INV_X1 U16933 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n15121) );
  NAND2_X1 U16934 ( .A1(n13937), .A2(n15121), .ZN(n13478) );
  NAND2_X1 U16935 ( .A1(n13479), .A2(n13478), .ZN(n14790) );
  NAND2_X1 U16936 ( .A1(n13740), .A2(n15121), .ZN(n13480) );
  OAI21_X1 U16937 ( .B1(n14790), .B2(n13740), .A(n13480), .ZN(n14815) );
  NAND2_X1 U16938 ( .A1(n13485), .A2(P1_EBX_REG_30__SCAN_IN), .ZN(n13482) );
  NAND2_X1 U16939 ( .A1(n14786), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13481) );
  NAND2_X1 U16940 ( .A1(n13482), .A2(n13481), .ZN(n14794) );
  NAND2_X1 U16941 ( .A1(n13484), .A2(n13483), .ZN(n13488) );
  AOI22_X1 U16942 ( .A1(P1_EBX_REG_31__SCAN_IN), .A2(n13485), .B1(n14786), 
        .B2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n13486) );
  INV_X1 U16943 ( .A(n13486), .ZN(n13487) );
  INV_X1 U16944 ( .A(n13489), .ZN(n13491) );
  AOI22_X1 U16945 ( .A1(n13491), .A2(n12296), .B1(n12289), .B2(n13490), .ZN(
        n13492) );
  NOR2_X1 U16946 ( .A1(n13500), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n13501) );
  MUX2_X1 U16947 ( .A(n13502), .B(n13501), .S(n11288), .Z(n15929) );
  NAND2_X1 U16948 ( .A1(n15929), .A2(n11452), .ZN(n13503) );
  XNOR2_X1 U16949 ( .A(n13503), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n13504) );
  AOI22_X1 U16950 ( .A1(n9737), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        n11689), .B2(P2_EAX_REG_31__SCAN_IN), .ZN(n13506) );
  NAND2_X1 U16951 ( .A1(n9739), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n13505) );
  AND2_X1 U16952 ( .A1(n13506), .A2(n13505), .ZN(n13507) );
  AOI22_X1 U16953 ( .A1(n11699), .A2(P2_REIP_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n13509) );
  OAI21_X1 U16954 ( .B1(n13510), .B2(n15931), .A(n13509), .ZN(n13511) );
  AOI21_X1 U16955 ( .B1(n13512), .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A(
        n13511), .ZN(n13513) );
  OAI21_X1 U16956 ( .B1(n17071), .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n13515), .ZN(n13519) );
  INV_X1 U16957 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n15932) );
  NOR2_X1 U16958 ( .A1(n16730), .A2(n15932), .ZN(n14716) );
  NOR4_X1 U16959 ( .A1(n16764), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n13517), .A4(n13516), .ZN(n13518) );
  AOI211_X1 U16960 ( .C1(n13519), .C2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A(
        n14716), .B(n13518), .ZN(n13520) );
  OAI21_X1 U16961 ( .B1(n15927), .B2(n17745), .A(n13520), .ZN(n13521) );
  AOI21_X1 U16962 ( .B1(n16394), .B2(n17741), .A(n13521), .ZN(n13524) );
  INV_X1 U16963 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n13523) );
  INV_X1 U16964 ( .A(n13490), .ZN(n14785) );
  AND2_X1 U16965 ( .A1(n14779), .A2(n14777), .ZN(n14783) );
  NAND2_X1 U16966 ( .A1(n14783), .A2(n14788), .ZN(n13739) );
  NAND2_X1 U16967 ( .A1(n15302), .A2(n13739), .ZN(n21910) );
  INV_X1 U16968 ( .A(n21907), .ZN(n17714) );
  NAND2_X1 U16969 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n17714), .ZN(n17628) );
  AND2_X1 U16970 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n21908), .ZN(n13525) );
  NAND2_X1 U16971 ( .A1(n13526), .A2(n13525), .ZN(n13527) );
  OAI211_X1 U16972 ( .C1(n17628), .C2(n21908), .A(n15837), .B(n13527), .ZN(
        n13528) );
  NAND2_X1 U16973 ( .A1(n14747), .A2(n21212), .ZN(n13550) );
  NOR2_X1 U16974 ( .A1(n15095), .A2(n21334), .ZN(n13541) );
  NAND2_X1 U16975 ( .A1(n15303), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n13537) );
  NAND2_X1 U16976 ( .A1(n21912), .A2(n21905), .ZN(n17622) );
  INV_X1 U16977 ( .A(n17622), .ZN(n13530) );
  NOR2_X1 U16978 ( .A1(n13537), .A2(n13530), .ZN(n13529) );
  AND2_X1 U16979 ( .A1(n13531), .A2(n13530), .ZN(n13539) );
  INV_X1 U16980 ( .A(n21251), .ZN(n14977) );
  INV_X1 U16981 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n15359) );
  INV_X1 U16982 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n22140) );
  INV_X1 U16983 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n21896) );
  INV_X1 U16984 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n21247) );
  INV_X1 U16985 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n21250) );
  NOR4_X1 U16986 ( .A1(n22140), .A2(n21896), .A3(n21247), .A4(n21250), .ZN(
        n21182) );
  INV_X1 U16987 ( .A(n21182), .ZN(n13532) );
  NAND4_X1 U16988 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(P1_REIP_REG_7__SCAN_IN), 
        .A3(P1_REIP_REG_6__SCAN_IN), .A4(P1_REIP_REG_5__SCAN_IN), .ZN(n21171)
         );
  NOR2_X1 U16989 ( .A1(n13532), .A2(n21171), .ZN(n17643) );
  NAND3_X1 U16990 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(P1_REIP_REG_9__SCAN_IN), 
        .A3(n17643), .ZN(n14978) );
  NAND2_X1 U16991 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(P1_REIP_REG_12__SCAN_IN), 
        .ZN(n15047) );
  NAND2_X1 U16992 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(P1_REIP_REG_14__SCAN_IN), 
        .ZN(n13533) );
  NOR2_X1 U16993 ( .A1(n15047), .A2(n13533), .ZN(n14998) );
  NAND2_X1 U16994 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(P1_REIP_REG_15__SCAN_IN), 
        .ZN(n15000) );
  INV_X1 U16995 ( .A(n15000), .ZN(n13534) );
  NAND3_X1 U16996 ( .A1(n14998), .A2(P1_REIP_REG_17__SCAN_IN), .A3(n13534), 
        .ZN(n13535) );
  NOR2_X1 U16997 ( .A1(n14978), .A2(n13535), .ZN(n14976) );
  NAND2_X1 U16998 ( .A1(n14976), .A2(P1_REIP_REG_18__SCAN_IN), .ZN(n14936) );
  NAND2_X1 U16999 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(P1_REIP_REG_19__SCAN_IN), 
        .ZN(n13536) );
  OR2_X1 U17000 ( .A1(n14936), .A2(n13536), .ZN(n14908) );
  INV_X1 U17001 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n21882) );
  NOR2_X1 U17002 ( .A1(n14908), .A2(n21882), .ZN(n14912) );
  AND2_X1 U17003 ( .A1(P1_REIP_REG_22__SCAN_IN), .A2(n14912), .ZN(n14893) );
  NAND2_X1 U17004 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(n14893), .ZN(n14884) );
  INV_X1 U17005 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n15408) );
  NOR2_X1 U17006 ( .A1(n14884), .A2(n15408), .ZN(n14872) );
  AND2_X1 U17007 ( .A1(n14872), .A2(P1_REIP_REG_25__SCAN_IN), .ZN(n14853) );
  NAND2_X1 U17008 ( .A1(n14853), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n14837) );
  INV_X1 U17009 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n21888) );
  INV_X1 U17010 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n22123) );
  OR3_X1 U17011 ( .A1(n14837), .A2(n21888), .A3(n22123), .ZN(n14810) );
  INV_X1 U17012 ( .A(n14810), .ZN(n14811) );
  NAND2_X1 U17013 ( .A1(P1_REIP_REG_29__SCAN_IN), .A2(n14811), .ZN(n14800) );
  NOR2_X1 U17014 ( .A1(n15359), .A2(n14800), .ZN(n13543) );
  OAI21_X1 U17015 ( .B1(n14977), .B2(n13543), .A(n21170), .ZN(n14801) );
  INV_X1 U17016 ( .A(n13537), .ZN(n13538) );
  NOR2_X1 U17017 ( .A1(n13539), .A2(n13538), .ZN(n13540) );
  INV_X1 U17018 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n14365) );
  OAI22_X1 U17019 ( .A1(n21256), .A2(n14365), .B1(n13542), .B2(n21253), .ZN(
        n13546) );
  INV_X1 U17020 ( .A(n13543), .ZN(n13544) );
  NOR3_X1 U17021 ( .A1(n14977), .A2(P1_REIP_REG_31__SCAN_IN), .A3(n13544), 
        .ZN(n13545) );
  AOI211_X1 U17022 ( .C1(P1_REIP_REG_31__SCAN_IN), .C2(n14801), .A(n13546), 
        .B(n13545), .ZN(n13547) );
  NAND2_X1 U17023 ( .A1(n13550), .A2(n13549), .ZN(P1_U2809) );
  NOR2_X1 U17024 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(n21116), .ZN(n13552) );
  NOR4_X1 U17025 ( .A1(P2_BE_N_REG_1__SCAN_IN), .A2(P2_BE_N_REG_2__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n13551) );
  NAND4_X1 U17026 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(n13552), .A3(n13551), .A4(
        n22104), .ZN(n13575) );
  NOR2_X4 U17027 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n13575), .ZN(n17904)
         );
  NOR4_X1 U17028 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(
        P1_ADDRESS_REG_14__SCAN_IN), .A3(P1_ADDRESS_REG_13__SCAN_IN), .A4(
        P1_ADDRESS_REG_12__SCAN_IN), .ZN(n13556) );
  NOR4_X1 U17029 ( .A1(P1_ADDRESS_REG_20__SCAN_IN), .A2(
        P1_ADDRESS_REG_19__SCAN_IN), .A3(P1_ADDRESS_REG_18__SCAN_IN), .A4(
        P1_ADDRESS_REG_16__SCAN_IN), .ZN(n13555) );
  NOR4_X1 U17030 ( .A1(P1_ADDRESS_REG_7__SCAN_IN), .A2(
        P1_ADDRESS_REG_6__SCAN_IN), .A3(P1_ADDRESS_REG_5__SCAN_IN), .A4(
        P1_ADDRESS_REG_4__SCAN_IN), .ZN(n13554) );
  NOR4_X1 U17031 ( .A1(P1_ADDRESS_REG_11__SCAN_IN), .A2(
        P1_ADDRESS_REG_10__SCAN_IN), .A3(P1_ADDRESS_REG_9__SCAN_IN), .A4(
        P1_ADDRESS_REG_8__SCAN_IN), .ZN(n13553) );
  AND4_X1 U17032 ( .A1(n13556), .A2(n13555), .A3(n13554), .A4(n13553), .ZN(
        n13561) );
  NOR4_X1 U17033 ( .A1(P1_ADDRESS_REG_2__SCAN_IN), .A2(
        P1_ADDRESS_REG_1__SCAN_IN), .A3(P1_ADDRESS_REG_0__SCAN_IN), .A4(
        P1_ADDRESS_REG_17__SCAN_IN), .ZN(n13559) );
  NOR4_X1 U17034 ( .A1(P1_ADDRESS_REG_24__SCAN_IN), .A2(
        P1_ADDRESS_REG_23__SCAN_IN), .A3(P1_ADDRESS_REG_22__SCAN_IN), .A4(
        P1_ADDRESS_REG_21__SCAN_IN), .ZN(n13558) );
  NOR4_X1 U17035 ( .A1(P1_ADDRESS_REG_28__SCAN_IN), .A2(
        P1_ADDRESS_REG_27__SCAN_IN), .A3(P1_ADDRESS_REG_26__SCAN_IN), .A4(
        P1_ADDRESS_REG_25__SCAN_IN), .ZN(n13557) );
  AND4_X1 U17036 ( .A1(n13559), .A2(n13558), .A3(n13557), .A4(n13613), .ZN(
        n13560) );
  NAND2_X1 U17037 ( .A1(n13561), .A2(n13560), .ZN(n13562) );
  NOR3_X1 U17038 ( .A1(P1_ADS_N_REG_SCAN_IN), .A2(P1_BE_N_REG_0__SCAN_IN), 
        .A3(n22167), .ZN(n13564) );
  NOR4_X1 U17039 ( .A1(P1_BE_N_REG_1__SCAN_IN), .A2(P1_BE_N_REG_2__SCAN_IN), 
        .A3(P1_BE_N_REG_3__SCAN_IN), .A4(P1_D_C_N_REG_SCAN_IN), .ZN(n13563) );
  NAND4_X1 U17040 ( .A1(n21327), .A2(P1_W_R_N_REG_SCAN_IN), .A3(n13564), .A4(
        n13563), .ZN(U214) );
  NOR4_X1 U17041 ( .A1(P2_ADDRESS_REG_17__SCAN_IN), .A2(
        P2_ADDRESS_REG_15__SCAN_IN), .A3(P2_ADDRESS_REG_13__SCAN_IN), .A4(
        P2_ADDRESS_REG_12__SCAN_IN), .ZN(n13568) );
  NOR4_X1 U17042 ( .A1(P2_ADDRESS_REG_20__SCAN_IN), .A2(
        P2_ADDRESS_REG_19__SCAN_IN), .A3(P2_ADDRESS_REG_16__SCAN_IN), .A4(
        P2_ADDRESS_REG_18__SCAN_IN), .ZN(n13567) );
  NOR4_X1 U17043 ( .A1(P2_ADDRESS_REG_7__SCAN_IN), .A2(
        P2_ADDRESS_REG_6__SCAN_IN), .A3(P2_ADDRESS_REG_5__SCAN_IN), .A4(
        P2_ADDRESS_REG_4__SCAN_IN), .ZN(n13566) );
  NOR4_X1 U17044 ( .A1(P2_ADDRESS_REG_11__SCAN_IN), .A2(
        P2_ADDRESS_REG_8__SCAN_IN), .A3(P2_ADDRESS_REG_10__SCAN_IN), .A4(
        P2_ADDRESS_REG_9__SCAN_IN), .ZN(n13565) );
  AND4_X1 U17045 ( .A1(n13568), .A2(n13567), .A3(n13566), .A4(n13565), .ZN(
        n13573) );
  NOR4_X1 U17046 ( .A1(P2_ADDRESS_REG_3__SCAN_IN), .A2(
        P2_ADDRESS_REG_1__SCAN_IN), .A3(P2_ADDRESS_REG_28__SCAN_IN), .A4(
        P2_ADDRESS_REG_14__SCAN_IN), .ZN(n13571) );
  NOR4_X1 U17047 ( .A1(P2_ADDRESS_REG_24__SCAN_IN), .A2(
        P2_ADDRESS_REG_23__SCAN_IN), .A3(P2_ADDRESS_REG_22__SCAN_IN), .A4(
        P2_ADDRESS_REG_21__SCAN_IN), .ZN(n13570) );
  NOR4_X1 U17048 ( .A1(P2_ADDRESS_REG_25__SCAN_IN), .A2(
        P2_ADDRESS_REG_2__SCAN_IN), .A3(P2_ADDRESS_REG_27__SCAN_IN), .A4(
        P2_ADDRESS_REG_26__SCAN_IN), .ZN(n13569) );
  INV_X1 U17049 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n13584) );
  NOR2_X1 U17050 ( .A1(n13584), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n21144) );
  INV_X1 U17051 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n13576) );
  OAI21_X1 U17052 ( .B1(n13576), .B2(P1_STATE_REG_2__SCAN_IN), .A(
        P1_STATE_REG_0__SCAN_IN), .ZN(n13577) );
  NOR2_X1 U17053 ( .A1(n13577), .A2(n21020), .ZN(n13580) );
  INV_X1 U17054 ( .A(n13580), .ZN(n13583) );
  AOI21_X1 U17055 ( .B1(NA), .B2(n13584), .A(P1_STATE_REG_0__SCAN_IN), .ZN(
        n13578) );
  NOR2_X1 U17056 ( .A1(n21912), .A2(n13584), .ZN(n15921) );
  OAI21_X1 U17057 ( .B1(n13578), .B2(n15921), .A(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n13582) );
  NOR2_X1 U17058 ( .A1(n21143), .A2(n13576), .ZN(n15922) );
  AND2_X1 U17059 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n15922), .ZN(n13579) );
  INV_X1 U17060 ( .A(NA), .ZN(n21010) );
  OAI211_X1 U17061 ( .C1(n13580), .C2(n13579), .A(n21010), .B(n17713), .ZN(
        n13581) );
  OAI211_X1 U17062 ( .C1(n21144), .C2(n13583), .A(n13582), .B(n13581), .ZN(
        P1_U3196) );
  AOI21_X1 U17063 ( .B1(n13584), .B2(n15923), .A(n21020), .ZN(n13585) );
  AOI211_X1 U17064 ( .C1(n21143), .C2(NA), .A(n13576), .B(n13585), .ZN(n13587)
         );
  OAI21_X1 U17065 ( .B1(n15921), .B2(n21143), .A(n15923), .ZN(n13586) );
  OAI21_X1 U17066 ( .B1(n13587), .B2(n21915), .A(n13586), .ZN(P1_U3194) );
  INV_X2 U17067 ( .A(n21915), .ZN(n21916) );
  INV_X1 U17068 ( .A(n13612), .ZN(n13610) );
  INV_X1 U17069 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n13596) );
  INV_X1 U17070 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n15836) );
  INV_X1 U17071 ( .A(P1_ADDRESS_REG_4__SCAN_IN), .ZN(n13588) );
  OAI222_X1 U17072 ( .A1(n13610), .A2(n13596), .B1(n21876), .B2(n15836), .C1(
        n21915), .C2(n13588), .ZN(P1_U3201) );
  INV_X1 U17073 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n17644) );
  AOI22_X1 U17074 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(n13612), .B1(
        P1_ADDRESS_REG_9__SCAN_IN), .B2(n21916), .ZN(n13589) );
  OAI21_X1 U17075 ( .B1(n17644), .B2(n21876), .A(n13589), .ZN(P1_U3206) );
  INV_X1 U17076 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n21880) );
  AOI22_X1 U17077 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(n13612), .B1(
        P1_ADDRESS_REG_12__SCAN_IN), .B2(n21916), .ZN(n13590) );
  OAI21_X1 U17078 ( .B1(n21880), .B2(n21876), .A(n13590), .ZN(P1_U3209) );
  INV_X1 U17079 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n15501) );
  AOI22_X1 U17080 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(n13612), .B1(
        P1_ADDRESS_REG_13__SCAN_IN), .B2(n21916), .ZN(n13591) );
  OAI21_X1 U17081 ( .B1(n15501), .B2(n21876), .A(n13591), .ZN(P1_U3210) );
  INV_X1 U17082 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n21878) );
  AOI22_X1 U17083 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(n13612), .B1(
        P1_ADDRESS_REG_8__SCAN_IN), .B2(n21916), .ZN(n13592) );
  OAI21_X1 U17084 ( .B1(n21878), .B2(n21876), .A(n13592), .ZN(P1_U3205) );
  AOI22_X1 U17085 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(n13612), .B1(
        P1_ADDRESS_REG_1__SCAN_IN), .B2(n21916), .ZN(n13593) );
  OAI21_X1 U17086 ( .B1(n21250), .B2(n21876), .A(n13593), .ZN(P1_U3198) );
  INV_X1 U17087 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n15491) );
  AOI22_X1 U17088 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(n13612), .B1(
        P1_ADDRESS_REG_14__SCAN_IN), .B2(n21916), .ZN(n13594) );
  OAI21_X1 U17089 ( .B1(n15491), .B2(n21876), .A(n13594), .ZN(P1_U3211) );
  AOI22_X1 U17090 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n13612), .B1(
        P1_ADDRESS_REG_5__SCAN_IN), .B2(n21916), .ZN(n13595) );
  OAI21_X1 U17091 ( .B1(n13596), .B2(n21876), .A(n13595), .ZN(P1_U3202) );
  INV_X1 U17092 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n13598) );
  AOI22_X1 U17093 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(n13612), .B1(
        P1_ADDRESS_REG_15__SCAN_IN), .B2(n21916), .ZN(n13597) );
  OAI21_X1 U17094 ( .B1(n13598), .B2(n21876), .A(n13597), .ZN(P1_U3212) );
  AOI22_X1 U17095 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(n13612), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n21916), .ZN(n13599) );
  OAI21_X1 U17096 ( .B1(n21888), .B2(n21876), .A(n13599), .ZN(P1_U3223) );
  AOI22_X1 U17097 ( .A1(P1_REIP_REG_29__SCAN_IN), .A2(n13612), .B1(
        P1_ADDRESS_REG_27__SCAN_IN), .B2(n21916), .ZN(n13600) );
  OAI21_X1 U17098 ( .B1(n22123), .B2(n21876), .A(n13600), .ZN(P1_U3224) );
  INV_X1 U17099 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n22188) );
  AOI22_X1 U17100 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(n13612), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n21916), .ZN(n13601) );
  OAI21_X1 U17101 ( .B1(n22188), .B2(n21876), .A(n13601), .ZN(P1_U3225) );
  INV_X1 U17102 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n22130) );
  AOI22_X1 U17103 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(n13612), .B1(
        P1_ADDRESS_REG_24__SCAN_IN), .B2(n21916), .ZN(n13602) );
  OAI21_X1 U17104 ( .B1(n22130), .B2(n21876), .A(n13602), .ZN(P1_U3221) );
  INV_X1 U17105 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n21884) );
  AOI22_X1 U17106 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(n13612), .B1(
        P1_ADDRESS_REG_22__SCAN_IN), .B2(n21916), .ZN(n13603) );
  OAI21_X1 U17107 ( .B1(n21884), .B2(n21876), .A(n13603), .ZN(P1_U3219) );
  AOI22_X1 U17108 ( .A1(P1_ADDRESS_REG_20__SCAN_IN), .A2(n21916), .B1(
        P1_REIP_REG_22__SCAN_IN), .B2(n13612), .ZN(n13604) );
  OAI21_X1 U17109 ( .B1(n21882), .B2(n21876), .A(n13604), .ZN(P1_U3217) );
  INV_X1 U17110 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n15472) );
  AOI22_X1 U17111 ( .A1(P1_ADDRESS_REG_16__SCAN_IN), .A2(n21916), .B1(
        P1_REIP_REG_18__SCAN_IN), .B2(n13612), .ZN(n13605) );
  OAI21_X1 U17112 ( .B1(n15472), .B2(n21876), .A(n13605), .ZN(P1_U3213) );
  INV_X1 U17113 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n21204) );
  AOI22_X1 U17114 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(n21916), .B1(
        P1_REIP_REG_8__SCAN_IN), .B2(n13612), .ZN(n13606) );
  OAI21_X1 U17115 ( .B1(n21204), .B2(n21876), .A(n13606), .ZN(P1_U3203) );
  INV_X1 U17116 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n15066) );
  AOI22_X1 U17117 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(n21916), .B1(
        P1_REIP_REG_12__SCAN_IN), .B2(n13612), .ZN(n13607) );
  OAI21_X1 U17118 ( .B1(n15066), .B2(n21876), .A(n13607), .ZN(P1_U3207) );
  INV_X1 U17119 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n14956) );
  AOI22_X1 U17120 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(n21916), .B1(
        P1_REIP_REG_20__SCAN_IN), .B2(n13612), .ZN(n13608) );
  OAI21_X1 U17121 ( .B1(n14956), .B2(n21876), .A(n13608), .ZN(P1_U3215) );
  INV_X1 U17122 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n15458) );
  INV_X1 U17123 ( .A(P1_ADDRESS_REG_17__SCAN_IN), .ZN(n13609) );
  OAI222_X1 U17124 ( .A1(n15458), .A2(n21876), .B1(n13610), .B2(n14956), .C1(
        n21915), .C2(n13609), .ZN(P1_U3214) );
  AOI22_X1 U17125 ( .A1(n21916), .A2(P1_ADDRESS_REG_2__SCAN_IN), .B1(
        P1_REIP_REG_4__SCAN_IN), .B2(n13612), .ZN(n13611) );
  OAI21_X1 U17126 ( .B1(n22140), .B2(n21876), .A(n13611), .ZN(P1_U3199) );
  INV_X1 U17127 ( .A(P1_ADDRESS_REG_0__SCAN_IN), .ZN(n22132) );
  OAI222_X1 U17128 ( .A1(n21876), .A2(n21896), .B1(n21250), .B2(n13610), .C1(
        n21915), .C2(n22132), .ZN(P1_U3197) );
  OAI222_X1 U17129 ( .A1(n21876), .A2(n21247), .B1(n21915), .B2(n13613), .C1(
        n15836), .C2(n13610), .ZN(P1_U3200) );
  INV_X1 U17130 ( .A(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n22151) );
  OAI222_X1 U17131 ( .A1(n21876), .A2(n15359), .B1(n21915), .B2(n22151), .C1(
        n22154), .C2(n13610), .ZN(P1_U3226) );
  INV_X1 U17132 ( .A(n13615), .ZN(n13616) );
  NAND2_X1 U17133 ( .A1(n14134), .A2(n13616), .ZN(n16305) );
  INV_X1 U17134 ( .A(n16305), .ZN(n13620) );
  INV_X1 U17135 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n13619) );
  INV_X1 U17136 ( .A(n13632), .ZN(n13618) );
  NOR2_X1 U17137 ( .A1(n20883), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n13627) );
  INV_X1 U17138 ( .A(n13627), .ZN(n13617) );
  OAI211_X1 U17139 ( .C1(n13620), .C2(n13619), .A(n13618), .B(n13617), .ZN(
        P2_U2814) );
  INV_X1 U17140 ( .A(n13629), .ZN(n21128) );
  INV_X1 U17141 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n13622) );
  NAND3_X1 U17142 ( .A1(n21106), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n21135), 
        .ZN(n13621) );
  OAI21_X1 U17143 ( .B1(n21128), .B2(n13622), .A(n13621), .ZN(P2_U2816) );
  INV_X1 U17144 ( .A(n13623), .ZN(n14133) );
  NAND2_X1 U17145 ( .A1(n11257), .A2(n21133), .ZN(n13812) );
  INV_X1 U17146 ( .A(n13812), .ZN(n13624) );
  NOR3_X1 U17147 ( .A1(n13813), .A2(n14133), .A3(n13624), .ZN(n17773) );
  NOR2_X1 U17148 ( .A1(n17773), .A2(n13625), .ZN(n21117) );
  INV_X1 U17149 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n14143) );
  OAI21_X1 U17150 ( .B1(n21117), .B2(n14143), .A(n13626), .ZN(P2_U2819) );
  OAI21_X1 U17151 ( .B1(n13627), .B2(P2_READREQUEST_REG_SCAN_IN), .A(n13629), 
        .ZN(n13628) );
  OAI21_X1 U17152 ( .B1(n13630), .B2(n13629), .A(n13628), .ZN(P2_U3612) );
  AND2_X1 U17153 ( .A1(n21819), .A2(n21871), .ZN(n14950) );
  NAND2_X1 U17154 ( .A1(n15302), .A2(n21149), .ZN(n13738) );
  AOI21_X1 U17155 ( .B1(P1_MEMORYFETCH_REG_SCAN_IN), .B2(n13739), .A(n13738), 
        .ZN(n13631) );
  INV_X1 U17156 ( .A(n13631), .ZN(P1_U2801) );
  AND2_X2 U17157 ( .A1(n13633), .A2(n13716), .ZN(n20352) );
  AOI22_X1 U17158 ( .A1(n20352), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(
        P2_EAX_REG_11__SCAN_IN), .B2(n20348), .ZN(n13636) );
  INV_X1 U17159 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n15215) );
  OR2_X1 U17160 ( .A1(n14329), .A2(n15215), .ZN(n13635) );
  NAND2_X1 U17161 ( .A1(n14329), .A2(BUF2_REG_11__SCAN_IN), .ZN(n13634) );
  NAND2_X1 U17162 ( .A1(n13635), .A2(n13634), .ZN(n16411) );
  NAND2_X1 U17163 ( .A1(n20350), .A2(n16411), .ZN(n13663) );
  NAND2_X1 U17164 ( .A1(n13636), .A2(n13663), .ZN(P2_U2978) );
  AOI22_X1 U17165 ( .A1(n20352), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(
        P2_EAX_REG_19__SCAN_IN), .B2(n20348), .ZN(n13639) );
  INV_X1 U17166 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n15263) );
  OR2_X1 U17167 ( .A1(n14329), .A2(n15263), .ZN(n13638) );
  NAND2_X1 U17168 ( .A1(n14329), .A2(BUF2_REG_3__SCAN_IN), .ZN(n13637) );
  AND2_X1 U17169 ( .A1(n13638), .A2(n13637), .ZN(n20408) );
  INV_X1 U17170 ( .A(n20408), .ZN(n16466) );
  NAND2_X1 U17171 ( .A1(n20350), .A2(n16466), .ZN(n13661) );
  NAND2_X1 U17172 ( .A1(n13639), .A2(n13661), .ZN(P2_U2955) );
  AOI22_X1 U17173 ( .A1(n20352), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(
        P2_EAX_REG_18__SCAN_IN), .B2(n20348), .ZN(n13643) );
  INV_X1 U17174 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n13640) );
  OR2_X1 U17175 ( .A1(n14329), .A2(n13640), .ZN(n13642) );
  NAND2_X1 U17176 ( .A1(n14329), .A2(BUF2_REG_2__SCAN_IN), .ZN(n13641) );
  NAND2_X1 U17177 ( .A1(n13642), .A2(n13641), .ZN(n16518) );
  NAND2_X1 U17178 ( .A1(n20350), .A2(n16518), .ZN(n13688) );
  NAND2_X1 U17179 ( .A1(n13643), .A2(n13688), .ZN(P2_U2954) );
  AOI22_X1 U17180 ( .A1(n20352), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(
        P2_EAX_REG_8__SCAN_IN), .B2(n20348), .ZN(n13647) );
  INV_X1 U17181 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n13644) );
  OR2_X1 U17182 ( .A1(n14329), .A2(n13644), .ZN(n13646) );
  NAND2_X1 U17183 ( .A1(n14329), .A2(BUF2_REG_8__SCAN_IN), .ZN(n13645) );
  AND2_X1 U17184 ( .A1(n13646), .A2(n13645), .ZN(n20287) );
  INV_X1 U17185 ( .A(n20287), .ZN(n16432) );
  NAND2_X1 U17186 ( .A1(n20350), .A2(n16432), .ZN(n13672) );
  NAND2_X1 U17187 ( .A1(n13647), .A2(n13672), .ZN(P2_U2975) );
  AOI22_X1 U17188 ( .A1(n20352), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(
        P2_EAX_REG_7__SCAN_IN), .B2(n20348), .ZN(n13651) );
  INV_X1 U17189 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n13648) );
  OR2_X1 U17190 ( .A1(n14329), .A2(n13648), .ZN(n13650) );
  NAND2_X1 U17191 ( .A1(n14329), .A2(BUF2_REG_7__SCAN_IN), .ZN(n13649) );
  NAND2_X1 U17192 ( .A1(n13650), .A2(n13649), .ZN(n16439) );
  NAND2_X1 U17193 ( .A1(n20350), .A2(n16439), .ZN(n13670) );
  NAND2_X1 U17194 ( .A1(n13651), .A2(n13670), .ZN(P2_U2974) );
  AOI22_X1 U17195 ( .A1(n20352), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(
        P2_EAX_REG_13__SCAN_IN), .B2(n20348), .ZN(n13654) );
  INV_X1 U17196 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n15203) );
  OR2_X1 U17197 ( .A1(n14329), .A2(n15203), .ZN(n13653) );
  NAND2_X1 U17198 ( .A1(n14329), .A2(BUF2_REG_13__SCAN_IN), .ZN(n13652) );
  NAND2_X1 U17199 ( .A1(n13653), .A2(n13652), .ZN(n16399) );
  NAND2_X1 U17200 ( .A1(n20350), .A2(n16399), .ZN(n13659) );
  NAND2_X1 U17201 ( .A1(n13654), .A2(n13659), .ZN(P2_U2980) );
  AOI22_X1 U17202 ( .A1(n20352), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(
        P2_EAX_REG_21__SCAN_IN), .B2(n20348), .ZN(n13658) );
  INV_X1 U17203 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n13655) );
  OR2_X1 U17204 ( .A1(n14329), .A2(n13655), .ZN(n13657) );
  NAND2_X1 U17205 ( .A1(n14329), .A2(BUF2_REG_5__SCAN_IN), .ZN(n13656) );
  NAND2_X1 U17206 ( .A1(n13657), .A2(n13656), .ZN(n20423) );
  NAND2_X1 U17207 ( .A1(n20350), .A2(n20423), .ZN(n13682) );
  NAND2_X1 U17208 ( .A1(n13658), .A2(n13682), .ZN(P2_U2957) );
  AOI22_X1 U17209 ( .A1(n20352), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(
        P2_EAX_REG_29__SCAN_IN), .B2(n20348), .ZN(n13660) );
  NAND2_X1 U17210 ( .A1(n13660), .A2(n13659), .ZN(P2_U2965) );
  AOI22_X1 U17211 ( .A1(n20352), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(
        P2_EAX_REG_3__SCAN_IN), .B2(n20348), .ZN(n13662) );
  NAND2_X1 U17212 ( .A1(n13662), .A2(n13661), .ZN(P2_U2970) );
  AOI22_X1 U17213 ( .A1(n20352), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(
        P2_EAX_REG_27__SCAN_IN), .B2(n20348), .ZN(n13664) );
  NAND2_X1 U17214 ( .A1(n13664), .A2(n13663), .ZN(P2_U2963) );
  AOI22_X1 U17215 ( .A1(n20352), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(
        P2_EAX_REG_1__SCAN_IN), .B2(n20348), .ZN(n13669) );
  INV_X1 U17216 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n13665) );
  OR2_X1 U17217 ( .A1(n14329), .A2(n13665), .ZN(n13667) );
  NAND2_X1 U17218 ( .A1(n14329), .A2(BUF2_REG_1__SCAN_IN), .ZN(n13666) );
  INV_X1 U17219 ( .A(n20393), .ZN(n13668) );
  NAND2_X1 U17220 ( .A1(n20350), .A2(n13668), .ZN(n13686) );
  NAND2_X1 U17221 ( .A1(n13669), .A2(n13686), .ZN(P2_U2968) );
  AOI22_X1 U17222 ( .A1(n20352), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(
        P2_EAX_REG_23__SCAN_IN), .B2(n20348), .ZN(n13671) );
  NAND2_X1 U17223 ( .A1(n13671), .A2(n13670), .ZN(P2_U2959) );
  AOI22_X1 U17224 ( .A1(n20352), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(
        P2_EAX_REG_24__SCAN_IN), .B2(n20348), .ZN(n13673) );
  NAND2_X1 U17225 ( .A1(n13673), .A2(n13672), .ZN(P2_U2960) );
  AOI22_X1 U17226 ( .A1(n20352), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(
        P2_EAX_REG_0__SCAN_IN), .B2(n20348), .ZN(n13677) );
  INV_X1 U17227 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n13674) );
  OR2_X1 U17228 ( .A1(n14329), .A2(n13674), .ZN(n13676) );
  NAND2_X1 U17229 ( .A1(n14329), .A2(BUF2_REG_0__SCAN_IN), .ZN(n13675) );
  AND2_X1 U17230 ( .A1(n13676), .A2(n13675), .ZN(n20381) );
  INV_X1 U17231 ( .A(n20381), .ZN(n16491) );
  NAND2_X1 U17232 ( .A1(n20350), .A2(n16491), .ZN(n13693) );
  NAND2_X1 U17233 ( .A1(n13677), .A2(n13693), .ZN(P2_U2967) );
  AOI22_X1 U17234 ( .A1(n20352), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(
        P2_EAX_REG_20__SCAN_IN), .B2(n20348), .ZN(n13681) );
  INV_X1 U17235 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n13678) );
  OR2_X1 U17236 ( .A1(n14329), .A2(n13678), .ZN(n13680) );
  NAND2_X1 U17237 ( .A1(n14329), .A2(BUF2_REG_4__SCAN_IN), .ZN(n13679) );
  NAND2_X1 U17238 ( .A1(n13680), .A2(n13679), .ZN(n16510) );
  NAND2_X1 U17239 ( .A1(n20350), .A2(n16510), .ZN(n13684) );
  NAND2_X1 U17240 ( .A1(n13681), .A2(n13684), .ZN(P2_U2956) );
  AOI22_X1 U17241 ( .A1(n20352), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(
        P2_EAX_REG_5__SCAN_IN), .B2(n20348), .ZN(n13683) );
  NAND2_X1 U17242 ( .A1(n13683), .A2(n13682), .ZN(P2_U2972) );
  AOI22_X1 U17243 ( .A1(n20352), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(
        P2_EAX_REG_4__SCAN_IN), .B2(n20348), .ZN(n13685) );
  NAND2_X1 U17244 ( .A1(n13685), .A2(n13684), .ZN(P2_U2971) );
  AOI22_X1 U17245 ( .A1(n20352), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(
        P2_EAX_REG_17__SCAN_IN), .B2(n20348), .ZN(n13687) );
  NAND2_X1 U17246 ( .A1(n13687), .A2(n13686), .ZN(P2_U2953) );
  AOI22_X1 U17247 ( .A1(n20352), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(
        P2_EAX_REG_2__SCAN_IN), .B2(n20348), .ZN(n13689) );
  NAND2_X1 U17248 ( .A1(n13689), .A2(n13688), .ZN(P2_U2969) );
  AOI22_X1 U17249 ( .A1(n20352), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(
        P2_EAX_REG_22__SCAN_IN), .B2(n20348), .ZN(n13692) );
  INV_X1 U17250 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n17871) );
  OR2_X1 U17251 ( .A1(n14329), .A2(n17871), .ZN(n13691) );
  NAND2_X1 U17252 ( .A1(n14329), .A2(BUF2_REG_6__SCAN_IN), .ZN(n13690) );
  NAND2_X1 U17253 ( .A1(n13691), .A2(n13690), .ZN(n16446) );
  NAND2_X1 U17254 ( .A1(n20350), .A2(n16446), .ZN(n13695) );
  NAND2_X1 U17255 ( .A1(n13692), .A2(n13695), .ZN(P2_U2958) );
  AOI22_X1 U17256 ( .A1(n20352), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(
        P2_EAX_REG_16__SCAN_IN), .B2(n20348), .ZN(n13694) );
  NAND2_X1 U17257 ( .A1(n13694), .A2(n13693), .ZN(P2_U2952) );
  AOI22_X1 U17258 ( .A1(n20352), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(
        P2_EAX_REG_6__SCAN_IN), .B2(n20348), .ZN(n13696) );
  NAND2_X1 U17259 ( .A1(n13696), .A2(n13695), .ZN(P2_U2973) );
  AOI22_X1 U17260 ( .A1(n20352), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(
        P2_EAX_REG_25__SCAN_IN), .B2(n20348), .ZN(n13699) );
  INV_X1 U17261 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n17866) );
  OR2_X1 U17262 ( .A1(n14329), .A2(n17866), .ZN(n13698) );
  NAND2_X1 U17263 ( .A1(n14329), .A2(BUF2_REG_9__SCAN_IN), .ZN(n13697) );
  NAND2_X1 U17264 ( .A1(n13698), .A2(n13697), .ZN(n16426) );
  NAND2_X1 U17265 ( .A1(n20350), .A2(n16426), .ZN(n13705) );
  NAND2_X1 U17266 ( .A1(n13699), .A2(n13705), .ZN(P2_U2961) );
  INV_X1 U17267 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n13700) );
  OR2_X1 U17268 ( .A1(n14329), .A2(n13700), .ZN(n13702) );
  NAND2_X1 U17269 ( .A1(n14329), .A2(BUF2_REG_15__SCAN_IN), .ZN(n13701) );
  NAND2_X1 U17270 ( .A1(n13702), .A2(n13701), .ZN(n14362) );
  AOI222_X1 U17271 ( .A1(n14362), .A2(n20350), .B1(P2_LWORD_REG_15__SCAN_IN), 
        .B2(n20352), .C1(P2_EAX_REG_15__SCAN_IN), .C2(n20348), .ZN(n13703) );
  INV_X1 U17272 ( .A(n13703), .ZN(P2_U2982) );
  INV_X1 U17273 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n20326) );
  NAND2_X1 U17274 ( .A1(n20352), .A2(P2_LWORD_REG_9__SCAN_IN), .ZN(n13704) );
  OAI211_X1 U17275 ( .C1(n20326), .C2(n13716), .A(n13705), .B(n13704), .ZN(
        P2_U2976) );
  INV_X1 U17276 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n13724) );
  INV_X1 U17277 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n17865) );
  OR2_X1 U17278 ( .A1(n14329), .A2(n17865), .ZN(n13707) );
  NAND2_X1 U17279 ( .A1(n14329), .A2(BUF2_REG_10__SCAN_IN), .ZN(n13706) );
  NAND2_X1 U17280 ( .A1(n13707), .A2(n13706), .ZN(n16418) );
  NAND2_X1 U17281 ( .A1(n20350), .A2(n16418), .ZN(n13710) );
  NAND2_X1 U17282 ( .A1(n20352), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n13708) );
  OAI211_X1 U17283 ( .C1(n13724), .C2(n13716), .A(n13710), .B(n13708), .ZN(
        P2_U2962) );
  INV_X1 U17284 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n22102) );
  NAND2_X1 U17285 ( .A1(n20352), .A2(P2_LWORD_REG_10__SCAN_IN), .ZN(n13709) );
  OAI211_X1 U17286 ( .C1(n22102), .C2(n13716), .A(n13710), .B(n13709), .ZN(
        P2_U2977) );
  INV_X1 U17287 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n22072) );
  INV_X1 U17288 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n22194) );
  OR2_X1 U17289 ( .A1(n14329), .A2(n22194), .ZN(n13712) );
  NAND2_X1 U17290 ( .A1(n14329), .A2(BUF2_REG_12__SCAN_IN), .ZN(n13711) );
  NAND2_X1 U17291 ( .A1(n13712), .A2(n13711), .ZN(n16405) );
  NAND2_X1 U17292 ( .A1(n20350), .A2(n16405), .ZN(n13715) );
  NAND2_X1 U17293 ( .A1(n20352), .A2(P2_LWORD_REG_12__SCAN_IN), .ZN(n13713) );
  OAI211_X1 U17294 ( .C1(n22072), .C2(n13716), .A(n13715), .B(n13713), .ZN(
        P2_U2979) );
  INV_X1 U17295 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n13727) );
  NAND2_X1 U17296 ( .A1(n20352), .A2(P2_UWORD_REG_12__SCAN_IN), .ZN(n13714) );
  OAI211_X1 U17297 ( .C1(n13727), .C2(n13716), .A(n13715), .B(n13714), .ZN(
        P2_U2964) );
  INV_X1 U17298 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n13720) );
  NAND2_X1 U17299 ( .A1(n14134), .A2(n17793), .ZN(n13717) );
  NAND2_X1 U17300 ( .A1(n21132), .A2(n14142), .ZN(n21125) );
  INV_X1 U17301 ( .A(P2_UWORD_REG_4__SCAN_IN), .ZN(n22215) );
  INV_X1 U17302 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n13719) );
  OAI222_X1 U17303 ( .A1(n13720), .A2(n20347), .B1(n21125), .B2(n22215), .C1(
        n13719), .C2(n13746), .ZN(P2_U2931) );
  INV_X1 U17304 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n13722) );
  INV_X1 U17305 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n16480) );
  INV_X1 U17306 ( .A(P2_UWORD_REG_1__SCAN_IN), .ZN(n13721) );
  OAI222_X1 U17307 ( .A1(n13722), .A2(n20347), .B1(n13746), .B2(n16480), .C1(
        n21125), .C2(n13721), .ZN(P2_U2934) );
  INV_X1 U17308 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n13725) );
  INV_X1 U17309 ( .A(P2_UWORD_REG_10__SCAN_IN), .ZN(n13723) );
  OAI222_X1 U17310 ( .A1(n13725), .A2(n20347), .B1(n13746), .B2(n13724), .C1(
        n21125), .C2(n13723), .ZN(P2_U2925) );
  INV_X1 U17311 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n13728) );
  INV_X1 U17312 ( .A(P2_UWORD_REG_12__SCAN_IN), .ZN(n13726) );
  OAI222_X1 U17313 ( .A1(n13728), .A2(n20347), .B1(n13746), .B2(n13727), .C1(
        n21125), .C2(n13726), .ZN(P2_U2923) );
  INV_X1 U17314 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n13731) );
  INV_X1 U17315 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n13730) );
  INV_X1 U17316 ( .A(P2_UWORD_REG_6__SCAN_IN), .ZN(n13729) );
  OAI222_X1 U17317 ( .A1(n13731), .A2(n20347), .B1(n13746), .B2(n13730), .C1(
        n21125), .C2(n13729), .ZN(P2_U2929) );
  INV_X1 U17318 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n13734) );
  INV_X1 U17319 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n13733) );
  INV_X1 U17320 ( .A(P2_UWORD_REG_2__SCAN_IN), .ZN(n13732) );
  OAI222_X1 U17321 ( .A1(n13734), .A2(n20347), .B1(n13746), .B2(n13733), .C1(
        n21125), .C2(n13732), .ZN(P2_U2933) );
  INV_X1 U17322 ( .A(P2_UWORD_REG_0__SCAN_IN), .ZN(n13737) );
  INV_X1 U17323 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n13736) );
  INV_X1 U17324 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n13735) );
  OAI222_X1 U17325 ( .A1(n13737), .A2(n21125), .B1(n13746), .B2(n13736), .C1(
        n13735), .C2(n20347), .ZN(P2_U2935) );
  OR2_X1 U17326 ( .A1(n13738), .A2(P1_READREQUEST_REG_SCAN_IN), .ZN(n13743) );
  INV_X1 U17327 ( .A(n13743), .ZN(n13745) );
  INV_X1 U17328 ( .A(n13739), .ZN(n13742) );
  OAI22_X1 U17329 ( .A1(n13743), .A2(n13742), .B1(n13741), .B2(n13740), .ZN(
        n13744) );
  OAI21_X1 U17330 ( .B1(n13745), .B2(n21910), .A(n13744), .ZN(P1_U3487) );
  INV_X1 U17331 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n13748) );
  AOI22_X1 U17332 ( .A1(n20313), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n20344), 
        .B2(P2_UWORD_REG_8__SCAN_IN), .ZN(n13747) );
  OAI21_X1 U17333 ( .B1(n20347), .B2(n13748), .A(n13747), .ZN(P2_U2927) );
  INV_X1 U17334 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n13750) );
  AOI22_X1 U17335 ( .A1(n20313), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n20344), 
        .B2(P2_UWORD_REG_9__SCAN_IN), .ZN(n13749) );
  OAI21_X1 U17336 ( .B1(n20347), .B2(n13750), .A(n13749), .ZN(P2_U2926) );
  INV_X1 U17337 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n13752) );
  AOI22_X1 U17338 ( .A1(n20313), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n20344), 
        .B2(P2_UWORD_REG_3__SCAN_IN), .ZN(n13751) );
  OAI21_X1 U17339 ( .B1(n20347), .B2(n13752), .A(n13751), .ZN(P2_U2932) );
  INV_X1 U17340 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n13754) );
  AOI22_X1 U17341 ( .A1(n20313), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n20344), 
        .B2(P2_UWORD_REG_5__SCAN_IN), .ZN(n13753) );
  OAI21_X1 U17342 ( .B1(n20347), .B2(n13754), .A(n13753), .ZN(P2_U2930) );
  INV_X1 U17343 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n13756) );
  AOI22_X1 U17344 ( .A1(n20313), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n20344), 
        .B2(P2_UWORD_REG_13__SCAN_IN), .ZN(n13755) );
  OAI21_X1 U17345 ( .B1(n20347), .B2(n13756), .A(n13755), .ZN(P2_U2922) );
  INV_X1 U17346 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n13758) );
  AOI22_X1 U17347 ( .A1(n20313), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n20344), 
        .B2(P2_UWORD_REG_7__SCAN_IN), .ZN(n13757) );
  OAI21_X1 U17348 ( .B1(n20347), .B2(n13758), .A(n13757), .ZN(P2_U2928) );
  INV_X1 U17349 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n13760) );
  AOI22_X1 U17350 ( .A1(n20313), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n20344), 
        .B2(P2_UWORD_REG_11__SCAN_IN), .ZN(n13759) );
  OAI21_X1 U17351 ( .B1(n20347), .B2(n13760), .A(n13759), .ZN(P2_U2924) );
  INV_X1 U17352 ( .A(n20370), .ZN(n20363) );
  INV_X1 U17353 ( .A(n20368), .ZN(n17725) );
  XNOR2_X1 U17354 ( .A(n13761), .B(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17109) );
  INV_X1 U17355 ( .A(n17109), .ZN(n13764) );
  OR2_X1 U17356 ( .A1(n17736), .A2(n16286), .ZN(n13763) );
  NOR2_X1 U17357 ( .A1(n20217), .A2(n21031), .ZN(n17107) );
  INV_X1 U17358 ( .A(n17107), .ZN(n13762) );
  OAI211_X1 U17359 ( .C1(n16762), .C2(n13764), .A(n13763), .B(n13762), .ZN(
        n13765) );
  AOI21_X1 U17360 ( .B1(n17725), .B2(n16286), .A(n13765), .ZN(n13768) );
  OR2_X1 U17361 ( .A1(n13766), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17112) );
  NAND3_X1 U17362 ( .A1(n17112), .A2(n11457), .A3(n17113), .ZN(n13767) );
  OAI211_X1 U17363 ( .C1(n17104), .C2(n20363), .A(n13768), .B(n13767), .ZN(
        P2_U3013) );
  XNOR2_X1 U17364 ( .A(n13769), .B(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13796) );
  NAND2_X1 U17365 ( .A1(n20355), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n13789) );
  INV_X1 U17366 ( .A(n13789), .ZN(n13772) );
  OAI21_X1 U17367 ( .B1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n16298), .A(
        n13770), .ZN(n13793) );
  NOR2_X1 U17368 ( .A1(n16737), .A2(n13793), .ZN(n13771) );
  AOI211_X1 U17369 ( .C1(n13796), .C2(n20357), .A(n13772), .B(n13771), .ZN(
        n13775) );
  OAI21_X1 U17370 ( .B1(n20356), .B2(n13773), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13774) );
  OAI211_X1 U17371 ( .C1(n13790), .C2(n20363), .A(n13775), .B(n13774), .ZN(
        P2_U3014) );
  NAND2_X1 U17372 ( .A1(n17774), .A2(n17776), .ZN(n14137) );
  NAND2_X1 U17373 ( .A1(n14137), .A2(n13776), .ZN(n13777) );
  NAND2_X1 U17374 ( .A1(n13779), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13780) );
  NOR2_X1 U17375 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13783) );
  OAI21_X1 U17376 ( .B1(n13784), .B2(n13783), .A(n13799), .ZN(n13785) );
  INV_X1 U17377 ( .A(n13785), .ZN(n13786) );
  NOR2_X1 U17378 ( .A1(n13790), .A2(n16386), .ZN(n13787) );
  AOI21_X1 U17379 ( .B1(P2_EBX_REG_0__SCAN_IN), .B2(n16386), .A(n13787), .ZN(
        n13788) );
  OAI21_X1 U17380 ( .B1(n16388), .B2(n20673), .A(n13788), .ZN(P2_U2887) );
  OAI21_X1 U17381 ( .B1(n17745), .B2(n13790), .A(n13789), .ZN(n13795) );
  XNOR2_X1 U17382 ( .A(n13792), .B(n13791), .ZN(n20302) );
  OAI22_X1 U17383 ( .A1(n17105), .A2(n20302), .B1(n17101), .B2(n13793), .ZN(
        n13794) );
  AOI211_X1 U17384 ( .C1(n17738), .C2(n13796), .A(n13795), .B(n13794), .ZN(
        n13798) );
  MUX2_X1 U17385 ( .A(n17071), .B(n17103), .S(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .Z(n13797) );
  NAND2_X1 U17386 ( .A1(n13798), .A2(n13797), .ZN(P2_U3046) );
  NAND2_X1 U17387 ( .A1(n13801), .A2(n14056), .ZN(n13803) );
  NAND2_X1 U17388 ( .A1(n20837), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n20838) );
  NAND2_X1 U17389 ( .A1(n21114), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20874) );
  NAND2_X1 U17390 ( .A1(n20838), .A2(n20874), .ZN(n20882) );
  AND2_X1 U17391 ( .A1(n20882), .A2(n20880), .ZN(n20479) );
  AOI21_X1 U17392 ( .B1(n14059), .B2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n20479), .ZN(n13802) );
  NAND2_X1 U17393 ( .A1(n13803), .A2(n13802), .ZN(n13804) );
  NAND2_X1 U17394 ( .A1(n13805), .A2(n13804), .ZN(n13806) );
  NOR2_X1 U17395 ( .A1(n17104), .A2(n16386), .ZN(n13807) );
  AOI21_X1 U17396 ( .B1(P2_EBX_REG_1__SCAN_IN), .B2(n16386), .A(n13807), .ZN(
        n13808) );
  OAI21_X1 U17397 ( .B1(n21099), .B2(n16388), .A(n13808), .ZN(P2_U2886) );
  OAI21_X1 U17398 ( .B1(n13811), .B2(n13810), .A(n13809), .ZN(n20275) );
  OAI22_X1 U17399 ( .A1(n17774), .A2(n14121), .B1(n13813), .B2(n13812), .ZN(
        n14135) );
  AND2_X1 U17400 ( .A1(n13815), .A2(n13814), .ZN(n13816) );
  NAND2_X1 U17401 ( .A1(n16519), .A2(n13818), .ZN(n20298) );
  INV_X1 U17402 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n20330) );
  AND2_X1 U17403 ( .A1(n16519), .A2(n9831), .ZN(n16492) );
  INV_X1 U17404 ( .A(n16492), .ZN(n16481) );
  NAND2_X1 U17405 ( .A1(n13779), .A2(n13819), .ZN(n13820) );
  INV_X1 U17406 ( .A(n14677), .ZN(n13821) );
  INV_X1 U17407 ( .A(n16439), .ZN(n20443) );
  OAI222_X1 U17408 ( .A1(n20275), .A2(n20283), .B1(n20330), .B2(n16519), .C1(
        n20311), .C2(n20443), .ZN(P2_U2912) );
  XOR2_X1 U17409 ( .A(n13822), .B(n13823), .Z(n17051) );
  INV_X1 U17410 ( .A(n17051), .ZN(n13824) );
  INV_X1 U17411 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n20332) );
  INV_X1 U17412 ( .A(n16446), .ZN(n20431) );
  OAI222_X1 U17413 ( .A1(n13824), .A2(n20283), .B1(n20332), .B2(n16519), .C1(
        n20311), .C2(n20431), .ZN(P2_U2913) );
  OAI211_X1 U17414 ( .C1(n9734), .C2(n13827), .A(n13826), .B(n15679), .ZN(
        n13829) );
  NAND2_X1 U17415 ( .A1(n13829), .A2(n13828), .ZN(n13844) );
  OR2_X1 U17416 ( .A1(n13485), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13830) );
  NAND2_X1 U17417 ( .A1(n13831), .A2(n13830), .ZN(n15115) );
  INV_X1 U17418 ( .A(n15682), .ZN(n15769) );
  OAI21_X1 U17419 ( .B1(n15766), .B2(n15769), .A(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13832) );
  NAND2_X1 U17420 ( .A1(n17697), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n13843) );
  OAI211_X1 U17421 ( .C1(n15115), .C2(n15839), .A(n13832), .B(n13843), .ZN(
        n13834) );
  NAND2_X1 U17422 ( .A1(n15851), .A2(n15679), .ZN(n13914) );
  INV_X1 U17423 ( .A(n13914), .ZN(n13833) );
  NOR3_X1 U17424 ( .A1(n13834), .A2(n15765), .A3(n13833), .ZN(n13835) );
  OAI21_X1 U17425 ( .B1(n15864), .B2(n13844), .A(n13835), .ZN(P1_U3031) );
  INV_X1 U17426 ( .A(n13836), .ZN(n13840) );
  INV_X1 U17427 ( .A(n13837), .ZN(n13839) );
  OAI21_X1 U17428 ( .B1(n13840), .B2(n13839), .A(n13838), .ZN(n15119) );
  OAI21_X1 U17429 ( .B1(n17661), .B2(n13841), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13842) );
  OAI211_X1 U17430 ( .C1(n13844), .C2(n21153), .A(n13843), .B(n13842), .ZN(
        n13845) );
  INV_X1 U17431 ( .A(n13845), .ZN(n13846) );
  OAI21_X1 U17432 ( .B1(n15119), .B2(n17671), .A(n13846), .ZN(P1_U2999) );
  OAI21_X1 U17433 ( .B1(n17713), .B2(n13847), .A(n13885), .ZN(n13848) );
  INV_X1 U17434 ( .A(n13848), .ZN(n13855) );
  NOR2_X1 U17435 ( .A1(n13849), .A2(n17713), .ZN(n13850) );
  NAND2_X1 U17436 ( .A1(n14779), .A2(n13850), .ZN(n13888) );
  AND3_X1 U17437 ( .A1(n12296), .A2(n21373), .A3(n13852), .ZN(n13936) );
  NAND2_X1 U17438 ( .A1(n13865), .A2(n13936), .ZN(n13853) );
  NOR2_X1 U17439 ( .A1(n13857), .A2(n13858), .ZN(n13859) );
  INV_X1 U17440 ( .A(n14748), .ZN(n13861) );
  INV_X1 U17441 ( .A(n21327), .ZN(n21329) );
  NAND2_X1 U17442 ( .A1(n21329), .A2(DATAI_0_), .ZN(n13863) );
  NAND2_X1 U17443 ( .A1(n21327), .A2(BUF1_REG_0__SCAN_IN), .ZN(n13862) );
  AND2_X1 U17444 ( .A1(n13863), .A2(n13862), .ZN(n21341) );
  INV_X1 U17445 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n22214) );
  OAI222_X1 U17446 ( .A1(n15299), .A2(n15119), .B1(n15298), .B2(n21341), .C1(
        n15296), .C2(n22214), .ZN(P1_U2904) );
  INV_X1 U17447 ( .A(n13865), .ZN(n13867) );
  INV_X1 U17448 ( .A(n13324), .ZN(n13881) );
  NAND4_X1 U17449 ( .A1(n13867), .A2(n13849), .A3(n13881), .A4(n13866), .ZN(
        n13868) );
  NOR2_X1 U17450 ( .A1(n13869), .A2(n13868), .ZN(n15904) );
  INV_X1 U17451 ( .A(n13934), .ZN(n14776) );
  NAND2_X1 U17452 ( .A1(n14776), .A2(n13885), .ZN(n13903) );
  NOR2_X1 U17453 ( .A1(n12123), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13897) );
  XNOR2_X1 U17454 ( .A(n13897), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13877) );
  XNOR2_X1 U17455 ( .A(n13870), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13875) );
  NOR2_X1 U17456 ( .A1(n12313), .A2(n15091), .ZN(n13871) );
  NAND2_X1 U17457 ( .A1(n13872), .A2(n13871), .ZN(n13900) );
  INV_X1 U17458 ( .A(n13873), .ZN(n13898) );
  AOI21_X1 U17459 ( .B1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n13898), .A(
        n13874), .ZN(n13879) );
  OAI22_X1 U17460 ( .A1(n15908), .A2(n13875), .B1(n13900), .B2(n13879), .ZN(
        n13876) );
  AOI21_X1 U17461 ( .B1(n13903), .B2(n13877), .A(n13876), .ZN(n13878) );
  OAI21_X1 U17462 ( .B1(n9922), .B2(n15904), .A(n13878), .ZN(n15866) );
  INV_X1 U17463 ( .A(n13879), .ZN(n13880) );
  AOI22_X1 U17464 ( .A1(n15866), .A2(n15911), .B1(n15916), .B2(n13880), .ZN(
        n13895) );
  NAND2_X1 U17465 ( .A1(n13881), .A2(n15908), .ZN(n13883) );
  NAND2_X1 U17466 ( .A1(n13847), .A2(n15925), .ZN(n13882) );
  NAND3_X1 U17467 ( .A1(n13883), .A2(n13882), .A3(n21912), .ZN(n13884) );
  AND2_X1 U17468 ( .A1(n13885), .A2(n13884), .ZN(n13886) );
  MUX2_X1 U17469 ( .A(n13886), .B(n14776), .S(n17629), .Z(n13893) );
  INV_X1 U17470 ( .A(n13887), .ZN(n13889) );
  OAI211_X1 U17471 ( .C1(n15094), .C2(n13890), .A(n13889), .B(n13888), .ZN(
        n13891) );
  INV_X1 U17472 ( .A(n13891), .ZN(n13892) );
  INV_X1 U17473 ( .A(n15878), .ZN(n17710) );
  NAND2_X1 U17474 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n17710), .ZN(n17715) );
  OAI22_X1 U17475 ( .A1(n17600), .A2(n21146), .B1(n17715), .B2(n22052), .ZN(
        n13924) );
  NAND2_X1 U17476 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n13947), .ZN(
        n13894) );
  OAI21_X1 U17477 ( .B1(n13895), .B2(n13947), .A(n13894), .ZN(P1_U3469) );
  INV_X1 U17478 ( .A(n13897), .ZN(n13899) );
  NAND2_X1 U17479 ( .A1(n13899), .A2(n13898), .ZN(n13905) );
  XNOR2_X1 U17480 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13901) );
  OAI22_X1 U17481 ( .A1(n15908), .A2(n13901), .B1(n13900), .B2(n13905), .ZN(
        n13902) );
  AOI21_X1 U17482 ( .B1(n13903), .B2(n13905), .A(n13902), .ZN(n13904) );
  OAI21_X1 U17483 ( .B1(n13896), .B2(n15904), .A(n13904), .ZN(n15867) );
  OAI22_X1 U17484 ( .A1(n12611), .A2(n15751), .B1(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n15913) );
  INV_X1 U17485 ( .A(n15913), .ZN(n13907) );
  NOR2_X1 U17486 ( .A1(n21871), .A2(n15679), .ZN(n15914) );
  INV_X1 U17487 ( .A(n13905), .ZN(n13906) );
  AOI222_X1 U17488 ( .A1(n15867), .A2(n15911), .B1(n13907), .B2(n15914), .C1(
        n15916), .C2(n13906), .ZN(n13909) );
  NAND2_X1 U17489 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n13947), .ZN(
        n13908) );
  OAI21_X1 U17490 ( .B1(n13909), .B2(n13947), .A(n13908), .ZN(P1_U3472) );
  XNOR2_X1 U17491 ( .A(n13910), .B(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n14040) );
  OR2_X1 U17492 ( .A1(n13911), .A2(n13937), .ZN(n13912) );
  NAND2_X1 U17493 ( .A1(n13913), .A2(n13912), .ZN(n15107) );
  NOR2_X1 U17494 ( .A1(n15837), .A2(n21896), .ZN(n14037) );
  AOI21_X1 U17495 ( .B1(n15814), .B2(n13914), .A(n15751), .ZN(n13915) );
  AOI211_X1 U17496 ( .C1(n17698), .C2(n15107), .A(n14037), .B(n13915), .ZN(
        n13918) );
  NAND3_X1 U17497 ( .A1(n17681), .A2(n15751), .A3(n13916), .ZN(n13917) );
  OAI211_X1 U17498 ( .C1(n14040), .C2(n15864), .A(n13918), .B(n13917), .ZN(
        P1_U3030) );
  AOI21_X1 U17499 ( .B1(n13920), .B2(n9771), .A(n11572), .ZN(n17010) );
  INV_X1 U17500 ( .A(n17010), .ZN(n20262) );
  INV_X1 U17501 ( .A(n20311), .ZN(n16505) );
  AOI22_X1 U17502 ( .A1(n16505), .A2(n16426), .B1(P2_EAX_REG_9__SCAN_IN), .B2(
        n20303), .ZN(n13921) );
  OAI21_X1 U17503 ( .B1(n20262), .B2(n20283), .A(n13921), .ZN(P2_U2910) );
  INV_X1 U17504 ( .A(n21470), .ZN(n21701) );
  NOR2_X1 U17505 ( .A1(n12445), .A2(n21701), .ZN(n13922) );
  XOR2_X1 U17506 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B(n13922), .Z(
        n21239) );
  INV_X1 U17507 ( .A(n13849), .ZN(n13923) );
  NAND2_X1 U17508 ( .A1(n21239), .A2(n13923), .ZN(n15873) );
  NAND2_X1 U17509 ( .A1(n13924), .A2(n15911), .ZN(n13925) );
  INV_X1 U17510 ( .A(n13947), .ZN(n15919) );
  OAI22_X1 U17511 ( .A1(n15873), .A2(n13925), .B1(n15872), .B2(n15919), .ZN(
        P1_U3468) );
  INV_X1 U17512 ( .A(n18097), .ZN(n13931) );
  INV_X1 U17513 ( .A(P3_REIP_REG_0__SCAN_IN), .ZN(n13930) );
  NAND3_X1 U17514 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n20140), .A3(
        n18242), .ZN(n13929) );
  NOR2_X1 U17515 ( .A1(n20177), .A2(n18818), .ZN(n20192) );
  INV_X1 U17516 ( .A(n20192), .ZN(n18293) );
  NOR2_X1 U17517 ( .A1(n9707), .A2(n18259), .ZN(n13926) );
  INV_X1 U17518 ( .A(P3_EBX_REG_0__SCAN_IN), .ZN(n18669) );
  OAI22_X1 U17519 ( .A1(n18293), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n13926), .B2(n18669), .ZN(n13927) );
  INV_X1 U17520 ( .A(n13927), .ZN(n13928) );
  OAI211_X1 U17521 ( .C1(n13931), .C2(n13930), .A(n13929), .B(n13928), .ZN(
        P3_U2671) );
  OAI21_X1 U17522 ( .B1(n13933), .B2(n13932), .A(n14115), .ZN(n15113) );
  NAND2_X1 U17523 ( .A1(n17629), .A2(n13934), .ZN(n13940) );
  INV_X1 U17524 ( .A(n13935), .ZN(n13938) );
  NAND3_X1 U17525 ( .A1(n13938), .A2(n13937), .A3(n13936), .ZN(n13939) );
  NAND2_X1 U17526 ( .A1(n13940), .A2(n13939), .ZN(n13941) );
  AOI22_X1 U17527 ( .A1(n15175), .A2(n15107), .B1(n15174), .B2(
        P1_EBX_REG_1__SCAN_IN), .ZN(n13942) );
  OAI21_X1 U17528 ( .B1(n15113), .B2(n15195), .A(n13942), .ZN(P1_U2871) );
  INV_X1 U17529 ( .A(n12709), .ZN(n15881) );
  OAI22_X1 U17530 ( .A1(n15881), .A2(n15904), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n15907), .ZN(n17598) );
  INV_X1 U17531 ( .A(n15916), .ZN(n13943) );
  OAI22_X1 U17532 ( .A1(n13943), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n21871), .ZN(n13944) );
  AOI21_X1 U17533 ( .B1(n15911), .B2(n17598), .A(n13944), .ZN(n13948) );
  NOR2_X1 U17534 ( .A1(n15908), .A2(n13945), .ZN(n17597) );
  AOI22_X1 U17535 ( .A1(n17597), .A2(n15911), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n13947), .ZN(n13946) );
  OAI21_X1 U17536 ( .B1(n13948), .B2(n13947), .A(n13946), .ZN(P1_U3474) );
  OAI21_X1 U17537 ( .B1(n15302), .B2(n15303), .A(n13949), .ZN(n13950) );
  INV_X1 U17538 ( .A(n15925), .ZN(n17621) );
  INV_X2 U17539 ( .A(n21281), .ZN(n21299) );
  AOI22_X1 U17540 ( .A1(P1_UWORD_REG_3__SCAN_IN), .A2(n21299), .B1(n21298), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n13951) );
  OAI21_X1 U17541 ( .B1(n15265), .B2(n21270), .A(n13951), .ZN(P1_U2917) );
  AOI22_X1 U17542 ( .A1(P1_UWORD_REG_11__SCAN_IN), .A2(n21299), .B1(n21298), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n13952) );
  OAI21_X1 U17543 ( .B1(n15217), .B2(n21270), .A(n13952), .ZN(P1_U2909) );
  AOI22_X1 U17544 ( .A1(P1_UWORD_REG_13__SCAN_IN), .A2(n21299), .B1(n21298), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n13953) );
  OAI21_X1 U17545 ( .B1(n15205), .B2(n21270), .A(n13953), .ZN(P1_U2907) );
  INV_X1 U17546 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n13955) );
  AOI22_X1 U17547 ( .A1(P1_UWORD_REG_8__SCAN_IN), .A2(n21299), .B1(n21298), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n13954) );
  OAI21_X1 U17548 ( .B1(n13955), .B2(n21270), .A(n13954), .ZN(P1_U2912) );
  INV_X1 U17549 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n13957) );
  AOI22_X1 U17550 ( .A1(P1_UWORD_REG_14__SCAN_IN), .A2(n21299), .B1(n21298), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n13956) );
  OAI21_X1 U17551 ( .B1(n13957), .B2(n21270), .A(n13956), .ZN(P1_U2906) );
  INV_X1 U17552 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n15222) );
  AOI22_X1 U17553 ( .A1(P1_UWORD_REG_10__SCAN_IN), .A2(n21299), .B1(n21298), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n13958) );
  OAI21_X1 U17554 ( .B1(n15222), .B2(n21270), .A(n13958), .ZN(P1_U2910) );
  AOI22_X1 U17555 ( .A1(P1_UWORD_REG_5__SCAN_IN), .A2(n21299), .B1(n21298), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n13959) );
  OAI21_X1 U17556 ( .B1(n15253), .B2(n21270), .A(n13959), .ZN(P1_U2915) );
  INV_X1 U17557 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n13961) );
  AOI22_X1 U17558 ( .A1(P1_UWORD_REG_2__SCAN_IN), .A2(n21299), .B1(n21298), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n13960) );
  OAI21_X1 U17559 ( .B1(n13961), .B2(n21270), .A(n13960), .ZN(P1_U2918) );
  INV_X1 U17560 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n13963) );
  AOI22_X1 U17561 ( .A1(P1_UWORD_REG_4__SCAN_IN), .A2(n21299), .B1(n21298), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n13962) );
  OAI21_X1 U17562 ( .B1(n13963), .B2(n21270), .A(n13962), .ZN(P1_U2916) );
  AOI22_X1 U17563 ( .A1(P1_UWORD_REG_6__SCAN_IN), .A2(n21299), .B1(n21298), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n13964) );
  OAI21_X1 U17564 ( .B1(n15246), .B2(n21270), .A(n13964), .ZN(P1_U2914) );
  INV_X1 U17565 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n13966) );
  AOI22_X1 U17566 ( .A1(P1_UWORD_REG_12__SCAN_IN), .A2(n21299), .B1(n21298), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n13965) );
  OAI21_X1 U17567 ( .B1(n13966), .B2(n21270), .A(n13965), .ZN(P1_U2908) );
  AOI22_X1 U17568 ( .A1(P1_UWORD_REG_7__SCAN_IN), .A2(n21299), .B1(n21298), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n13967) );
  OAI21_X1 U17569 ( .B1(n15240), .B2(n21270), .A(n13967), .ZN(P1_U2913) );
  NOR3_X1 U17570 ( .A1(n13968), .A2(n14012), .A3(n18765), .ZN(n13979) );
  AND2_X1 U17571 ( .A1(n17459), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n13969) );
  NOR2_X1 U17572 ( .A1(n13970), .A2(n13969), .ZN(n14177) );
  INV_X1 U17573 ( .A(n13971), .ZN(n13972) );
  NAND3_X1 U17574 ( .A1(n13973), .A2(n14177), .A3(n13972), .ZN(n13976) );
  NOR2_X1 U17575 ( .A1(n14178), .A2(n13974), .ZN(n13975) );
  NOR2_X1 U17576 ( .A1(n19547), .A2(n13977), .ZN(n19977) );
  INV_X1 U17577 ( .A(n19977), .ZN(n13978) );
  INV_X1 U17578 ( .A(P3_EBX_REG_2__SCAN_IN), .ZN(n18275) );
  INV_X1 U17579 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n18663) );
  NOR2_X1 U17580 ( .A1(n18669), .A2(n18663), .ZN(n18657) );
  INV_X1 U17581 ( .A(n18657), .ZN(n18292) );
  NOR2_X1 U17582 ( .A1(n18275), .A2(n18292), .ZN(n18648) );
  INV_X1 U17583 ( .A(n18640), .ZN(n18652) );
  NAND3_X1 U17584 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(P3_EBX_REG_5__SCAN_IN), 
        .A3(n18652), .ZN(n18642) );
  INV_X1 U17585 ( .A(n18642), .ZN(n18636) );
  NAND3_X1 U17586 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(P3_EBX_REG_7__SCAN_IN), 
        .A3(n18636), .ZN(n18606) );
  NOR2_X1 U17587 ( .A1(n18191), .A2(n18606), .ZN(n18608) );
  NAND4_X1 U17588 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(P3_EBX_REG_9__SCAN_IN), 
        .A3(P3_EBX_REG_8__SCAN_IN), .A4(P3_EBX_REG_7__SCAN_IN), .ZN(n18581) );
  OAI22_X1 U17589 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n18608), .B1(n18642), 
        .B2(n18581), .ZN(n14001) );
  INV_X2 U17590 ( .A(n10660), .ZN(n18403) );
  AOI22_X1 U17591 ( .A1(n18626), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n18403), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13986) );
  AOI22_X1 U17592 ( .A1(n11911), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n14232), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13985) );
  OR2_X1 U17593 ( .A1(n18599), .A2(n13982), .ZN(n13984) );
  NAND2_X1 U17594 ( .A1(n9726), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n13983) );
  NAND4_X1 U17595 ( .A1(n13986), .A2(n13985), .A3(n13984), .A4(n13983), .ZN(
        n13999) );
  NAND2_X1 U17596 ( .A1(n9724), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n13987) );
  OAI21_X1 U17597 ( .B1(n18454), .B2(n18616), .A(n13987), .ZN(n13989) );
  INV_X1 U17598 ( .A(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n19575) );
  OAI22_X1 U17599 ( .A1(n18613), .A2(n22105), .B1(n9723), .B2(n19575), .ZN(
        n13988) );
  NOR2_X1 U17600 ( .A1(n13989), .A2(n13988), .ZN(n13997) );
  AOI22_X1 U17601 ( .A1(n18586), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n18390), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13996) );
  NAND2_X1 U17602 ( .A1(n18620), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n13991) );
  NAND2_X1 U17603 ( .A1(n18489), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n13990) );
  OAI211_X1 U17604 ( .C1(n17550), .C2(n13992), .A(n13991), .B(n13990), .ZN(
        n13993) );
  INV_X1 U17605 ( .A(n13993), .ZN(n13995) );
  INV_X1 U17606 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n18660) );
  NAND2_X1 U17607 ( .A1(n18591), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n13994) );
  NAND4_X1 U17608 ( .A1(n13997), .A2(n13996), .A3(n13995), .A4(n13994), .ZN(
        n13998) );
  OR2_X1 U17609 ( .A1(n13999), .A2(n13998), .ZN(n18786) );
  NAND2_X1 U17610 ( .A1(n18667), .A2(n18786), .ZN(n14000) );
  OAI21_X1 U17611 ( .B1(n14001), .B2(n18667), .A(n14000), .ZN(P3_U2693) );
  INV_X1 U17612 ( .A(DATAI_1_), .ZN(n14003) );
  NAND2_X1 U17613 ( .A1(n21327), .A2(BUF1_REG_1__SCAN_IN), .ZN(n14002) );
  OAI21_X1 U17614 ( .B1(n21327), .B2(n14003), .A(n14002), .ZN(n15306) );
  INV_X1 U17615 ( .A(n15306), .ZN(n21349) );
  INV_X1 U17616 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n21297) );
  OAI222_X1 U17617 ( .A1(n15299), .A2(n15113), .B1(n15298), .B2(n21349), .C1(
        n15296), .C2(n21297), .ZN(P1_U2903) );
  INV_X1 U17618 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n14004) );
  OAI222_X1 U17619 ( .A1(n15115), .A2(n15192), .B1(n14004), .B2(n15194), .C1(
        n15119), .C2(n15187), .ZN(P1_U2872) );
  INV_X1 U17620 ( .A(n14005), .ZN(n14006) );
  AOI21_X1 U17621 ( .B1(n14007), .B2(n13919), .A(n14006), .ZN(n16995) );
  INV_X1 U17622 ( .A(n16995), .ZN(n14009) );
  INV_X1 U17623 ( .A(n16418), .ZN(n14008) );
  OAI222_X1 U17624 ( .A1(n14009), .A2(n20283), .B1(n14008), .B2(n20311), .C1(
        n22102), .C2(n16519), .ZN(P2_U2909) );
  NAND2_X1 U17625 ( .A1(n17927), .A2(n20181), .ZN(n14010) );
  NOR2_X1 U17626 ( .A1(n14010), .A2(n18816), .ZN(n14021) );
  OAI21_X1 U17627 ( .B1(n14012), .B2(n14011), .A(n14110), .ZN(n14013) );
  INV_X1 U17628 ( .A(n14013), .ZN(n14015) );
  NOR3_X1 U17629 ( .A1(n14015), .A2(n14014), .A3(n14026), .ZN(n14192) );
  AND2_X1 U17630 ( .A1(n14192), .A2(n14016), .ZN(n14017) );
  OR2_X1 U17631 ( .A1(n17918), .A2(n14017), .ZN(n14020) );
  INV_X1 U17632 ( .A(n14018), .ZN(n14019) );
  NAND2_X1 U17633 ( .A1(n14020), .A2(n14019), .ZN(n14185) );
  NOR4_X2 U17634 ( .A1(n14022), .A2(n14091), .A3(n14021), .A4(n14185), .ZN(
        n20025) );
  OR2_X1 U17635 ( .A1(n20025), .A2(n20042), .ZN(n14024) );
  INV_X1 U17636 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n19523) );
  NOR3_X1 U17637 ( .A1(n20044), .A2(n20175), .A3(n20187), .ZN(n17578) );
  INV_X1 U17638 ( .A(n17578), .ZN(n20137) );
  NOR2_X1 U17639 ( .A1(n19523), .A2(n20137), .ZN(n17577) );
  NOR2_X1 U17640 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n20138), .ZN(n19531) );
  NOR2_X1 U17641 ( .A1(n17577), .A2(n19531), .ZN(n14023) );
  NOR2_X2 U17642 ( .A1(n14025), .A2(n10371), .ZN(n19349) );
  NOR2_X1 U17643 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n19978), .ZN(
        n19983) );
  NAND2_X1 U17644 ( .A1(n14026), .A2(n20171), .ZN(n14029) );
  INV_X1 U17645 ( .A(n14027), .ZN(n14028) );
  OAI21_X1 U17646 ( .B1(n14030), .B2(n14029), .A(n14028), .ZN(n19975) );
  AND2_X1 U17647 ( .A1(n14110), .A2(n19424), .ZN(n17458) );
  INV_X1 U17648 ( .A(n14031), .ZN(n14032) );
  INV_X1 U17649 ( .A(n18270), .ZN(n19992) );
  NAND2_X1 U17650 ( .A1(n14032), .A2(n19992), .ZN(n18294) );
  OAI22_X1 U17651 ( .A1(n19983), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B1(
        n17458), .B2(n18294), .ZN(n20006) );
  INV_X1 U17652 ( .A(n20140), .ZN(n20188) );
  INV_X1 U17653 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n22165) );
  NOR2_X1 U17654 ( .A1(n20044), .A2(n22165), .ZN(n20153) );
  INV_X1 U17655 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n17443) );
  INV_X1 U17656 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n17394) );
  OAI22_X1 U17657 ( .A1(n17443), .A2(n17394), .B1(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20149) );
  NAND2_X1 U17658 ( .A1(n18236), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n20039) );
  INV_X1 U17659 ( .A(n18294), .ZN(n14033) );
  AOI222_X1 U17660 ( .A1(n20006), .A2(n20188), .B1(n20153), .B2(n20149), .C1(
        n20151), .C2(n14033), .ZN(n14035) );
  NAND2_X1 U17661 ( .A1(n20158), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n14034) );
  OAI21_X1 U17662 ( .B1(n20158), .B2(n14035), .A(n14034), .ZN(P3_U3289) );
  INV_X1 U17663 ( .A(n15113), .ZN(n14038) );
  MUX2_X1 U17664 ( .A(n15576), .B(n17661), .S(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .Z(n14036) );
  AOI211_X1 U17665 ( .C1(n14038), .C2(n21328), .A(n14037), .B(n14036), .ZN(
        n14039) );
  OAI21_X1 U17666 ( .B1(n14040), .B2(n21153), .A(n14039), .ZN(P1_U2998) );
  NAND2_X1 U17667 ( .A1(n14041), .A2(n14056), .ZN(n14043) );
  NAND2_X1 U17668 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n17754) );
  XNOR2_X1 U17669 ( .A(n17754), .B(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n20807) );
  AND2_X1 U17670 ( .A1(n20807), .A2(n20880), .ZN(n20542) );
  AOI21_X1 U17671 ( .B1(n14059), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n20542), .ZN(n14042) );
  NAND2_X1 U17672 ( .A1(n14043), .A2(n14042), .ZN(n14045) );
  OR2_X1 U17673 ( .A1(n14045), .A2(n14044), .ZN(n14046) );
  NAND2_X1 U17674 ( .A1(n14045), .A2(n14044), .ZN(n14054) );
  OR2_X1 U17675 ( .A1(n13800), .A2(n14047), .ZN(n14048) );
  MUX2_X1 U17676 ( .A(n17146), .B(P2_EBX_REG_2__SCAN_IN), .S(n16386), .Z(
        n14052) );
  AOI21_X1 U17677 ( .B1(n20373), .B2(n10619), .A(n14052), .ZN(n14053) );
  INV_X1 U17678 ( .A(n14053), .ZN(P2_U2885) );
  NAND2_X1 U17679 ( .A1(n17733), .A2(n14056), .ZN(n14061) );
  OAI21_X1 U17680 ( .B1(n17754), .B2(n22183), .A(n21096), .ZN(n14057) );
  INV_X1 U17681 ( .A(n17754), .ZN(n20782) );
  NAND2_X1 U17682 ( .A1(n20782), .A2(n20936), .ZN(n20938) );
  AND3_X1 U17683 ( .A1(n14057), .A2(n20938), .A3(n20880), .ZN(n14058) );
  AOI21_X1 U17684 ( .B1(n14059), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n14058), .ZN(n14060) );
  NOR2_X1 U17685 ( .A1(n17744), .A2(n16386), .ZN(n14066) );
  AOI21_X1 U17686 ( .B1(P2_EBX_REG_3__SCAN_IN), .B2(n16386), .A(n14066), .ZN(
        n14067) );
  OAI21_X1 U17687 ( .B1(n21090), .B2(n16388), .A(n14067), .ZN(P2_U2884) );
  AOI22_X1 U17688 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n21299), .B1(n21298), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n14068) );
  OAI21_X1 U17689 ( .B1(n15277), .B2(n21270), .A(n14068), .ZN(P1_U2920) );
  INV_X1 U17690 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n14070) );
  AOI22_X1 U17691 ( .A1(P1_UWORD_REG_1__SCAN_IN), .A2(n21299), .B1(n21298), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n14069) );
  OAI21_X1 U17692 ( .B1(n14070), .B2(n21270), .A(n14069), .ZN(P1_U2919) );
  XNOR2_X1 U17693 ( .A(n14072), .B(n14071), .ZN(n14206) );
  AND2_X1 U17694 ( .A1(n14075), .A2(n14074), .ZN(n14076) );
  OR2_X1 U17695 ( .A1(n14073), .A2(n14076), .ZN(n15099) );
  INV_X1 U17696 ( .A(n15099), .ZN(n14118) );
  NAND2_X1 U17697 ( .A1(n17697), .A2(P1_REIP_REG_2__SCAN_IN), .ZN(n14203) );
  INV_X1 U17698 ( .A(n14203), .ZN(n14080) );
  NOR2_X1 U17699 ( .A1(n15751), .A2(n15793), .ZN(n14078) );
  OAI21_X1 U17700 ( .B1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n15816), .A(
        n15814), .ZN(n14077) );
  MUX2_X1 U17701 ( .A(n14078), .B(n14077), .S(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .Z(n14079) );
  AOI211_X1 U17702 ( .C1(n17698), .C2(n14118), .A(n14080), .B(n14079), .ZN(
        n14084) );
  NOR2_X1 U17703 ( .A1(n15679), .A2(n15751), .ZN(n14081) );
  AOI21_X1 U17704 ( .B1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n14081), .A(
        n15850), .ZN(n14082) );
  OR2_X1 U17705 ( .A1(n15771), .A2(n14082), .ZN(n14083) );
  OAI211_X1 U17706 ( .C1(n14206), .C2(n15864), .A(n14084), .B(n14083), .ZN(
        P1_U3029) );
  AOI21_X1 U17707 ( .B1(n14086), .B2(n14005), .A(n14085), .ZN(n16975) );
  INV_X1 U17708 ( .A(n16975), .ZN(n14088) );
  INV_X1 U17709 ( .A(n16411), .ZN(n14087) );
  INV_X1 U17710 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n20323) );
  OAI222_X1 U17711 ( .A1(n14088), .A2(n20283), .B1(n14087), .B2(n20311), .C1(
        n20323), .C2(n16519), .ZN(P2_U2908) );
  INV_X1 U17712 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n18895) );
  INV_X1 U17713 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n18889) );
  NOR3_X1 U17714 ( .A1(n14089), .A2(n18818), .A3(n20171), .ZN(n14090) );
  NAND2_X1 U17715 ( .A1(n14246), .A2(n19561), .ZN(n18724) );
  NOR3_X1 U17716 ( .A1(n18889), .A2(n18887), .A3(n18724), .ZN(n14223) );
  NAND2_X1 U17717 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n18809), .ZN(n14093) );
  INV_X1 U17718 ( .A(n14093), .ZN(n18814) );
  AOI21_X1 U17719 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n18810), .A(n18814), .ZN(
        n14113) );
  NAND2_X1 U17720 ( .A1(n18585), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n14097) );
  NAND2_X1 U17721 ( .A1(n9724), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n14096) );
  NAND2_X1 U17722 ( .A1(n17547), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n14095) );
  NAND2_X1 U17723 ( .A1(n11911), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n14094) );
  AOI22_X1 U17724 ( .A1(n18586), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17561), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n14103) );
  INV_X1 U17725 ( .A(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n18420) );
  NAND2_X1 U17726 ( .A1(n18620), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n14099) );
  NAND2_X1 U17727 ( .A1(n18619), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n14098) );
  OAI211_X1 U17728 ( .C1(n17550), .C2(n18420), .A(n14099), .B(n14098), .ZN(
        n14100) );
  INV_X1 U17729 ( .A(n14100), .ZN(n14102) );
  NAND2_X1 U17730 ( .A1(n18413), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n14101) );
  NAND4_X1 U17731 ( .A1(n9814), .A2(n14103), .A3(n14102), .A4(n14101), .ZN(
        n14109) );
  AOI22_X1 U17732 ( .A1(n18390), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n18403), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n14107) );
  AOI22_X1 U17733 ( .A1(n18626), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n14232), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n14106) );
  INV_X1 U17734 ( .A(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n18554) );
  OR2_X1 U17735 ( .A1(n18599), .A2(n18554), .ZN(n14105) );
  NAND2_X1 U17736 ( .A1(n9726), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n14104) );
  NAND4_X1 U17737 ( .A1(n14107), .A2(n14106), .A3(n14105), .A4(n14104), .ZN(
        n14108) );
  NOR2_X2 U17738 ( .A1(n14110), .A2(n10253), .ZN(n18785) );
  NAND2_X1 U17739 ( .A1(n14110), .A2(n18784), .ZN(n18815) );
  INV_X1 U17740 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n19546) );
  OAI22_X1 U17741 ( .A1(n17287), .A2(n18812), .B1(n18815), .B2(n19546), .ZN(
        n14111) );
  INV_X1 U17742 ( .A(n14111), .ZN(n14112) );
  OAI21_X1 U17743 ( .B1(n18805), .B2(n14113), .A(n14112), .ZN(P3_U2731) );
  NAND2_X1 U17744 ( .A1(n14114), .A2(n15178), .ZN(n14116) );
  OR2_X1 U17745 ( .A1(n14116), .A2(n14115), .ZN(n15179) );
  NAND2_X1 U17746 ( .A1(n14116), .A2(n14115), .ZN(n14117) );
  AND2_X1 U17747 ( .A1(n15179), .A2(n14117), .ZN(n15093) );
  INV_X1 U17748 ( .A(n15093), .ZN(n14201) );
  AOI22_X1 U17749 ( .A1(n15175), .A2(n14118), .B1(n15174), .B2(
        P1_EBX_REG_2__SCAN_IN), .ZN(n14119) );
  OAI21_X1 U17750 ( .B1(n14201), .B2(n15195), .A(n14119), .ZN(P1_U2870) );
  INV_X1 U17751 ( .A(n14120), .ZN(n17798) );
  AND2_X1 U17752 ( .A1(n14122), .A2(n14121), .ZN(n17155) );
  NOR2_X1 U17753 ( .A1(n10700), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n17148) );
  INV_X1 U17754 ( .A(n14123), .ZN(n14460) );
  OAI22_X1 U17755 ( .A1(n17148), .A2(n14126), .B1(n14460), .B2(n10700), .ZN(
        n14132) );
  INV_X1 U17756 ( .A(n14124), .ZN(n17145) );
  NAND2_X1 U17757 ( .A1(n17733), .A2(n17145), .ZN(n14131) );
  OAI21_X1 U17758 ( .B1(n17147), .B2(n14126), .A(n14125), .ZN(n14129) );
  XNOR2_X1 U17759 ( .A(n10693), .B(n14126), .ZN(n14128) );
  AOI22_X1 U17760 ( .A1(n17152), .A2(n14129), .B1(n14128), .B2(n17150), .ZN(
        n14130) );
  OAI211_X1 U17761 ( .C1(n17155), .C2(n14132), .A(n14131), .B(n14130), .ZN(
        n17753) );
  AOI22_X1 U17762 ( .A1(n20671), .A2(n17798), .B1(n21086), .B2(n17753), .ZN(
        n14145) );
  NAND2_X1 U17763 ( .A1(n14134), .A2(n14133), .ZN(n14140) );
  INV_X1 U17764 ( .A(n14135), .ZN(n14139) );
  AND2_X1 U17765 ( .A1(n14137), .A2(n14136), .ZN(n14138) );
  OAI211_X1 U17766 ( .C1(n14141), .C2(n14140), .A(n14139), .B(n14138), .ZN(
        n17771) );
  NAND2_X1 U17767 ( .A1(n14142), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n17806) );
  OAI22_X1 U17768 ( .A1(n21106), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n14143), 
        .B2(n17806), .ZN(n14144) );
  MUX2_X1 U17769 ( .A(n14145), .B(n14126), .S(n17168), .Z(n14146) );
  INV_X1 U17770 ( .A(n14146), .ZN(P2_U3596) );
  OAI21_X1 U17771 ( .B1(n14085), .B2(n14148), .A(n14147), .ZN(n16964) );
  INV_X1 U17772 ( .A(n16405), .ZN(n14149) );
  OAI222_X1 U17773 ( .A1(n16964), .A2(n20283), .B1(n14149), .B2(n20311), .C1(
        n22072), .C2(n16519), .ZN(P2_U2907) );
  AOI22_X1 U17774 ( .A1(n9724), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n14232), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n14154) );
  AOI22_X1 U17775 ( .A1(n18620), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n18619), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n14153) );
  INV_X1 U17776 ( .A(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n18623) );
  INV_X1 U17777 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n18497) );
  OAI22_X1 U17778 ( .A1(n18616), .A2(n18623), .B1(n11880), .B2(n18497), .ZN(
        n14150) );
  INV_X1 U17779 ( .A(n14150), .ZN(n14152) );
  NAND2_X1 U17780 ( .A1(n18586), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n14151) );
  AOI22_X1 U17781 ( .A1(n18628), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9726), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n14156) );
  AOI22_X1 U17782 ( .A1(n18585), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n18597), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n14155) );
  INV_X1 U17783 ( .A(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17479) );
  NAND2_X1 U17784 ( .A1(n18413), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n14158) );
  NAND2_X1 U17785 ( .A1(n11911), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n14157) );
  OAI211_X1 U17786 ( .C1(n17550), .C2(n17479), .A(n14158), .B(n14157), .ZN(
        n14159) );
  NOR2_X1 U17787 ( .A1(n17296), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17368) );
  NAND2_X1 U17788 ( .A1(n9724), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n14161) );
  NAND2_X1 U17789 ( .A1(n17561), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n14160) );
  INV_X1 U17790 ( .A(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n17502) );
  NAND2_X1 U17791 ( .A1(n18620), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n14163) );
  NAND2_X1 U17792 ( .A1(n18489), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n14162) );
  OAI211_X1 U17793 ( .C1(n17550), .C2(n17502), .A(n14163), .B(n14162), .ZN(
        n14164) );
  NAND2_X1 U17794 ( .A1(n18597), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n14168) );
  NAND2_X1 U17795 ( .A1(n11911), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n14167) );
  NAND2_X1 U17796 ( .A1(n18627), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n14166) );
  NAND2_X1 U17797 ( .A1(n14232), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n14165) );
  AOI22_X1 U17798 ( .A1(n18628), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n9726), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n14173) );
  NAND2_X1 U17799 ( .A1(n18413), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n14171) );
  NAND2_X1 U17800 ( .A1(n18586), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n14170) );
  NAND2_X1 U17801 ( .A1(n18390), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n14169) );
  AND3_X1 U17802 ( .A1(n14171), .A2(n14170), .A3(n14169), .ZN(n14172) );
  NAND2_X1 U17803 ( .A1(n17295), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17294) );
  XNOR2_X1 U17804 ( .A(n17368), .B(n17228), .ZN(n17367) );
  NAND2_X1 U17805 ( .A1(n14175), .A2(n14174), .ZN(n20189) );
  NAND2_X1 U17806 ( .A1(n14178), .A2(n14177), .ZN(n17170) );
  NAND2_X1 U17807 ( .A1(n19539), .A2(n20171), .ZN(n14180) );
  NOR2_X1 U17808 ( .A1(n19555), .A2(n14180), .ZN(n14193) );
  NAND2_X1 U17809 ( .A1(n17170), .A2(n14193), .ZN(n14183) );
  AOI21_X1 U17810 ( .B1(n19535), .B2(n14179), .A(n20170), .ZN(n14181) );
  INV_X1 U17811 ( .A(n20181), .ZN(n20172) );
  AOI21_X1 U17812 ( .B1(n14181), .B2(n14180), .A(n20172), .ZN(n17928) );
  NAND2_X1 U17813 ( .A1(n17928), .A2(n14189), .ZN(n14182) );
  NAND2_X1 U17814 ( .A1(n14183), .A2(n14182), .ZN(n14184) );
  NAND2_X1 U17815 ( .A1(n14184), .A2(n17927), .ZN(n14187) );
  INV_X1 U17816 ( .A(n14185), .ZN(n14186) );
  OAI211_X1 U17817 ( .C1(n14189), .C2(n14188), .A(n14187), .B(n14186), .ZN(
        n14190) );
  NAND2_X1 U17818 ( .A1(n19355), .A2(n19457), .ZN(n19493) );
  AOI211_X1 U17819 ( .C1(n19349), .C2(n22165), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B(n19493), .ZN(n14197) );
  NOR2_X1 U17820 ( .A1(n19986), .A2(n19444), .ZN(n19381) );
  INV_X1 U17821 ( .A(n19381), .ZN(n19306) );
  NAND3_X1 U17822 ( .A1(n19457), .A2(n22165), .A3(n19306), .ZN(n19519) );
  AOI21_X1 U17823 ( .B1(n19512), .B2(n19519), .A(n17443), .ZN(n14196) );
  NAND2_X1 U17824 ( .A1(n14193), .A2(n14192), .ZN(n17398) );
  XNOR2_X1 U17825 ( .A(n17228), .B(n10672), .ZN(n17363) );
  INV_X2 U17826 ( .A(n14191), .ZN(n19508) );
  NAND2_X1 U17827 ( .A1(n19508), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n14194) );
  OAI21_X1 U17828 ( .B1(n19505), .B2(n17363), .A(n14194), .ZN(n14195) );
  NOR3_X1 U17829 ( .A1(n14197), .A2(n14196), .A3(n14195), .ZN(n14198) );
  OAI21_X1 U17830 ( .B1(n17367), .B2(n10011), .A(n14198), .ZN(P3_U2861) );
  INV_X1 U17831 ( .A(DATAI_2_), .ZN(n14200) );
  NAND2_X1 U17832 ( .A1(n21327), .A2(BUF1_REG_2__SCAN_IN), .ZN(n14199) );
  OAI21_X1 U17833 ( .B1(n21327), .B2(n14200), .A(n14199), .ZN(n15308) );
  INV_X1 U17834 ( .A(n15308), .ZN(n21352) );
  INV_X1 U17835 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n21295) );
  OAI222_X1 U17836 ( .A1(n15299), .A2(n14201), .B1(n15298), .B2(n21352), .C1(
        n15296), .C2(n21295), .ZN(P1_U2902) );
  NAND2_X1 U17837 ( .A1(n17661), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n14202) );
  OAI211_X1 U17838 ( .C1(n17670), .C2(n15104), .A(n14203), .B(n14202), .ZN(
        n14204) );
  AOI21_X1 U17839 ( .B1(n15093), .B2(n21328), .A(n14204), .ZN(n14205) );
  OAI21_X1 U17840 ( .B1(n21153), .B2(n14206), .A(n14205), .ZN(P1_U2997) );
  NAND2_X1 U17841 ( .A1(n13779), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n14207) );
  AND2_X1 U17842 ( .A1(n14599), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n14214) );
  INV_X1 U17843 ( .A(n14214), .ZN(n14209) );
  NAND2_X1 U17844 ( .A1(n14210), .A2(n14209), .ZN(n14215) );
  AND2_X1 U17845 ( .A1(n14211), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n14212) );
  NAND2_X1 U17846 ( .A1(n14271), .A2(n14214), .ZN(n14284) );
  OAI21_X1 U17847 ( .B1(n14213), .B2(n14215), .A(n14284), .ZN(n16508) );
  INV_X1 U17848 ( .A(n14216), .ZN(n14220) );
  NAND2_X1 U17849 ( .A1(n14218), .A2(n14217), .ZN(n14219) );
  NAND2_X1 U17850 ( .A1(n14220), .A2(n14219), .ZN(n20362) );
  MUX2_X1 U17851 ( .A(n20362), .B(n14221), .S(n16386), .Z(n14222) );
  OAI21_X1 U17852 ( .B1(n16508), .B2(n16388), .A(n14222), .ZN(P2_U2883) );
  AOI21_X1 U17853 ( .B1(P3_EAX_REG_2__SCAN_IN), .B2(n18810), .A(n14223), .ZN(
        n14245) );
  NAND2_X1 U17854 ( .A1(n18585), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n14227) );
  NAND2_X1 U17855 ( .A1(n9724), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n14226) );
  NAND2_X1 U17856 ( .A1(n17547), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n14225) );
  NAND2_X1 U17857 ( .A1(n17561), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n14224) );
  NAND4_X1 U17858 ( .A1(n14227), .A2(n14226), .A3(n14225), .A4(n14224), .ZN(
        n14231) );
  INV_X1 U17859 ( .A(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17468) );
  NAND2_X1 U17860 ( .A1(n18620), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n14229) );
  NAND2_X1 U17861 ( .A1(n18489), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n14228) );
  OAI211_X1 U17862 ( .C1(n17550), .C2(n17468), .A(n14229), .B(n14228), .ZN(
        n14230) );
  NOR2_X1 U17863 ( .A1(n14231), .A2(n14230), .ZN(n14243) );
  NAND2_X1 U17864 ( .A1(n18597), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n14236) );
  NAND2_X1 U17865 ( .A1(n11911), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n14235) );
  NAND2_X1 U17866 ( .A1(n18627), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n14234) );
  NAND2_X1 U17867 ( .A1(n14232), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n14233) );
  AND4_X1 U17868 ( .A1(n14236), .A2(n14235), .A3(n14234), .A4(n14233), .ZN(
        n14242) );
  AOI22_X1 U17869 ( .A1(n18628), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9726), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n14241) );
  NAND2_X1 U17870 ( .A1(n18413), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n14239) );
  NAND2_X1 U17871 ( .A1(n18586), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n14238) );
  NAND2_X1 U17872 ( .A1(n18390), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n14237) );
  AND3_X1 U17873 ( .A1(n14239), .A2(n14238), .A3(n14237), .ZN(n14240) );
  NAND4_X1 U17874 ( .A1(n14243), .A2(n14242), .A3(n14241), .A4(n14240), .ZN(
        n17278) );
  AOI22_X1 U17875 ( .A1(n17278), .A2(n18785), .B1(n18796), .B2(
        BUF2_REG_2__SCAN_IN), .ZN(n14244) );
  OAI21_X1 U17876 ( .B1(n14245), .B2(n18809), .A(n14244), .ZN(P3_U2733) );
  NOR2_X1 U17877 ( .A1(n18887), .A2(n18724), .ZN(n14248) );
  NOR2_X1 U17878 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n18724), .ZN(n14247) );
  OAI22_X1 U17879 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(n14248), .B1(n14247), .B2(
        n18672), .ZN(n14250) );
  AOI22_X1 U17880 ( .A1(n17295), .A2(n18785), .B1(BUF2_REG_1__SCAN_IN), .B2(
        n18796), .ZN(n14249) );
  NAND2_X1 U17881 ( .A1(n14250), .A2(n14249), .ZN(P3_U2734) );
  XOR2_X1 U17882 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B(n14284), .Z(n14255)
         );
  OAI21_X1 U17883 ( .B1(n14216), .B2(n14252), .A(n14251), .ZN(n16228) );
  INV_X1 U17884 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n14253) );
  MUX2_X1 U17885 ( .A(n16228), .B(n14253), .S(n16386), .Z(n14254) );
  OAI21_X1 U17886 ( .B1(n14255), .B2(n16388), .A(n14254), .ZN(P2_U2882) );
  AOI22_X1 U17887 ( .A1(n17296), .A2(n18785), .B1(BUF2_REG_0__SCAN_IN), .B2(
        n18796), .ZN(n14257) );
  NAND2_X1 U17888 ( .A1(n10253), .A2(P3_EAX_REG_0__SCAN_IN), .ZN(n14256) );
  OAI211_X1 U17889 ( .C1(n18724), .C2(P3_EAX_REG_0__SCAN_IN), .A(n14257), .B(
        n14256), .ZN(P3_U2735) );
  NAND2_X1 U17890 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n14267) );
  NOR2_X1 U17891 ( .A1(n14284), .A2(n14267), .ZN(n14334) );
  XNOR2_X1 U17892 ( .A(n14334), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n14263) );
  AND2_X1 U17893 ( .A1(n14258), .A2(n14259), .ZN(n14260) );
  NOR2_X1 U17894 ( .A1(n14258), .A2(n14259), .ZN(n16197) );
  OR2_X1 U17895 ( .A1(n14260), .A2(n16197), .ZN(n20278) );
  INV_X1 U17896 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n14261) );
  MUX2_X1 U17897 ( .A(n20278), .B(n14261), .S(n16386), .Z(n14262) );
  OAI21_X1 U17898 ( .B1(n14263), .B2(n16388), .A(n14262), .ZN(P2_U2880) );
  OAI21_X1 U17899 ( .B1(n10567), .B2(n10684), .A(n14264), .ZN(n16957) );
  INV_X1 U17900 ( .A(n16399), .ZN(n14265) );
  INV_X1 U17901 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n20320) );
  OAI222_X1 U17902 ( .A1(n16957), .A2(n20283), .B1(n14265), .B2(n20311), .C1(
        n20320), .C2(n16519), .ZN(P2_U2906) );
  INV_X1 U17903 ( .A(n14599), .ZN(n14578) );
  NAND2_X1 U17904 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n14266) );
  NOR2_X1 U17905 ( .A1(n14267), .A2(n14266), .ZN(n14268) );
  NAND3_X1 U17906 ( .A1(n14335), .A2(n14336), .A3(n14268), .ZN(n14269) );
  NOR2_X1 U17907 ( .A1(n14578), .A2(n14269), .ZN(n14270) );
  INV_X1 U17908 ( .A(n14321), .ZN(n14274) );
  INV_X1 U17909 ( .A(n14319), .ZN(n14272) );
  NOR2_X1 U17910 ( .A1(n14321), .A2(n14272), .ZN(n14312) );
  INV_X1 U17911 ( .A(n14312), .ZN(n14273) );
  OAI211_X1 U17912 ( .C1(n14274), .C2(n14319), .A(n14273), .B(n10619), .ZN(
        n14280) );
  INV_X1 U17913 ( .A(n14276), .ZN(n14277) );
  AOI21_X1 U17914 ( .B1(n14278), .B2(n14275), .A(n14277), .ZN(n16987) );
  NAND2_X1 U17915 ( .A1(n16987), .A2(n16363), .ZN(n14279) );
  OAI211_X1 U17916 ( .C1(n16363), .C2(n11185), .A(n14280), .B(n14279), .ZN(
        P2_U2877) );
  NAND2_X1 U17917 ( .A1(n14251), .A2(n14281), .ZN(n14282) );
  NAND2_X1 U17918 ( .A1(n14258), .A2(n14282), .ZN(n17054) );
  NOR2_X1 U17919 ( .A1(n14284), .A2(n14283), .ZN(n14286) );
  INV_X1 U17920 ( .A(n14334), .ZN(n14285) );
  OAI211_X1 U17921 ( .C1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .C2(n14286), .A(
        n14285), .B(n10619), .ZN(n14288) );
  NAND2_X1 U17922 ( .A1(n16386), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n14287) );
  OAI211_X1 U17923 ( .C1(n17054), .C2(n16368), .A(n14288), .B(n14287), .ZN(
        P2_U2881) );
  INV_X1 U17924 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n18899) );
  NAND2_X1 U17925 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n18805), .ZN(n14289) );
  NOR2_X1 U17926 ( .A1(n18899), .A2(n14289), .ZN(n18801) );
  INV_X1 U17927 ( .A(n14289), .ZN(n18808) );
  AOI21_X1 U17928 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n18810), .A(n18808), .ZN(
        n14308) );
  NAND2_X1 U17929 ( .A1(n18585), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n14293) );
  NAND2_X1 U17930 ( .A1(n9724), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n14292) );
  NAND2_X1 U17931 ( .A1(n17547), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n14291) );
  NAND2_X1 U17932 ( .A1(n11911), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n14290) );
  NAND4_X1 U17933 ( .A1(n14293), .A2(n14292), .A3(n14291), .A4(n14290), .ZN(
        n14297) );
  INV_X1 U17934 ( .A(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n18306) );
  NAND2_X1 U17935 ( .A1(n18620), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n14295) );
  NAND2_X1 U17936 ( .A1(n18619), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n14294) );
  OAI211_X1 U17937 ( .C1(n17550), .C2(n18306), .A(n14295), .B(n14294), .ZN(
        n14296) );
  NOR2_X1 U17938 ( .A1(n14297), .A2(n14296), .ZN(n14306) );
  AOI22_X1 U17939 ( .A1(n18390), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n18403), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n14299) );
  AOI22_X1 U17940 ( .A1(n18597), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n14232), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n14298) );
  AND2_X1 U17941 ( .A1(n14299), .A2(n14298), .ZN(n14305) );
  AOI22_X1 U17942 ( .A1(n18628), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n9726), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n14304) );
  INV_X1 U17943 ( .A(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n22203) );
  NAND2_X1 U17944 ( .A1(n18413), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n14301) );
  NAND2_X1 U17945 ( .A1(n18586), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n14300) );
  OAI211_X1 U17946 ( .C1(n18644), .C2(n9723), .A(n14301), .B(n14300), .ZN(
        n14302) );
  INV_X1 U17947 ( .A(n14302), .ZN(n14303) );
  NAND4_X1 U17948 ( .A1(n14306), .A2(n14305), .A3(n14304), .A4(n14303), .ZN(
        n17281) );
  AOI22_X1 U17949 ( .A1(n17281), .A2(n18785), .B1(BUF2_REG_6__SCAN_IN), .B2(
        n18796), .ZN(n14307) );
  OAI21_X1 U17950 ( .B1(n18801), .B2(n14308), .A(n14307), .ZN(P3_U2729) );
  NAND2_X1 U17951 ( .A1(n14276), .A2(n14310), .ZN(n14311) );
  NAND2_X1 U17952 ( .A1(n14309), .A2(n14311), .ZN(n16982) );
  NAND2_X1 U17953 ( .A1(n14312), .A2(n14320), .ZN(n16379) );
  OAI211_X1 U17954 ( .C1(n14312), .C2(n14320), .A(n16379), .B(n10619), .ZN(
        n14314) );
  NAND2_X1 U17955 ( .A1(n16386), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n14313) );
  OAI211_X1 U17956 ( .C1(n16982), .C2(n16368), .A(n14314), .B(n14313), .ZN(
        P2_U2876) );
  NAND2_X1 U17957 ( .A1(n14316), .A2(n14317), .ZN(n14318) );
  NAND2_X1 U17958 ( .A1(n14315), .A2(n14318), .ZN(n20241) );
  OAI211_X1 U17959 ( .C1(n14322), .C2(n14323), .A(n14354), .B(n10619), .ZN(
        n14325) );
  NAND2_X1 U17960 ( .A1(n16368), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n14324) );
  OAI211_X1 U17961 ( .C1(n20241), .C2(n16368), .A(n14325), .B(n14324), .ZN(
        P2_U2873) );
  AOI21_X1 U17962 ( .B1(n14327), .B2(n14264), .A(n14326), .ZN(n20245) );
  INV_X1 U17963 ( .A(n20245), .ZN(n14333) );
  INV_X1 U17964 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n14328) );
  OR2_X1 U17965 ( .A1(n14329), .A2(n14328), .ZN(n14331) );
  NAND2_X1 U17966 ( .A1(n14329), .A2(BUF2_REG_14__SCAN_IN), .ZN(n14330) );
  NAND2_X1 U17967 ( .A1(n14331), .A2(n14330), .ZN(n20349) );
  AOI22_X1 U17968 ( .A1(n16505), .A2(n20349), .B1(P2_EAX_REG_14__SCAN_IN), 
        .B2(n20303), .ZN(n14332) );
  OAI21_X1 U17969 ( .B1(n14333), .B2(n20283), .A(n14332), .ZN(P2_U2905) );
  NAND2_X1 U17970 ( .A1(n14334), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n16389) );
  INV_X1 U17971 ( .A(n14335), .ZN(n16390) );
  NOR2_X1 U17972 ( .A1(n16389), .A2(n16390), .ZN(n16387) );
  OAI211_X1 U17973 ( .C1(n16387), .C2(n14336), .A(n10619), .B(n14321), .ZN(
        n14342) );
  OR2_X1 U17974 ( .A1(n14337), .A2(n14338), .ZN(n14339) );
  NAND2_X1 U17975 ( .A1(n14275), .A2(n14339), .ZN(n20261) );
  INV_X1 U17976 ( .A(n20261), .ZN(n14340) );
  NAND2_X1 U17977 ( .A1(n14340), .A2(n16363), .ZN(n14341) );
  OAI211_X1 U17978 ( .C1(n16363), .C2(n11301), .A(n14342), .B(n14341), .ZN(
        P2_U2878) );
  INV_X1 U17979 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n14351) );
  INV_X1 U17980 ( .A(n16382), .ZN(n14343) );
  NOR2_X1 U17981 ( .A1(n16379), .A2(n14343), .ZN(n16380) );
  INV_X1 U17982 ( .A(n14322), .ZN(n14344) );
  OAI211_X1 U17983 ( .C1(n16380), .C2(n14345), .A(n10619), .B(n14344), .ZN(
        n14350) );
  OR2_X1 U17984 ( .A1(n14346), .A2(n14347), .ZN(n14348) );
  AND2_X1 U17985 ( .A1(n14348), .A2(n14316), .ZN(n16960) );
  NAND2_X1 U17986 ( .A1(n16960), .A2(n16363), .ZN(n14349) );
  OAI211_X1 U17987 ( .C1(n16363), .C2(n14351), .A(n14350), .B(n14349), .ZN(
        P2_U2874) );
  AOI21_X1 U17988 ( .B1(n14353), .B2(n14315), .A(n14352), .ZN(n16922) );
  NAND2_X1 U17989 ( .A1(n16922), .A2(n16363), .ZN(n14357) );
  INV_X1 U17990 ( .A(n14354), .ZN(n14355) );
  OAI211_X1 U17991 ( .C1(n14355), .C2(n9861), .A(n10619), .B(n14366), .ZN(
        n14356) );
  OAI211_X1 U17992 ( .C1(n16363), .C2(n14358), .A(n14357), .B(n14356), .ZN(
        P2_U2872) );
  NOR2_X1 U17993 ( .A1(n14326), .A2(n14360), .ZN(n14361) );
  OR2_X1 U17994 ( .A1(n14359), .A2(n14361), .ZN(n16921) );
  INV_X1 U17995 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n20316) );
  INV_X1 U17996 ( .A(n14362), .ZN(n14363) );
  OAI222_X1 U17997 ( .A1(n16921), .A2(n20283), .B1(n16519), .B2(n20316), .C1(
        n14363), .C2(n20311), .ZN(P2_U2904) );
  OAI22_X1 U17998 ( .A1(n14364), .A2(n15192), .B1(n15194), .B2(n14365), .ZN(
        P1_U2841) );
  AOI22_X1 U17999 ( .A1(n10758), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n14493), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n14373) );
  AOI22_X1 U18000 ( .A1(n10759), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n14477), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n14372) );
  INV_X1 U18001 ( .A(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n14462) );
  NAND2_X1 U18002 ( .A1(n10732), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n14368) );
  NAND2_X1 U18003 ( .A1(n10733), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n14367) );
  OAI211_X1 U18004 ( .C1(n14497), .C2(n14462), .A(n14368), .B(n14367), .ZN(
        n14369) );
  INV_X1 U18005 ( .A(n14369), .ZN(n14371) );
  AOI22_X1 U18006 ( .A1(n10764), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n14444), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n14370) );
  NAND4_X1 U18007 ( .A1(n14373), .A2(n14372), .A3(n14371), .A4(n14370), .ZN(
        n14379) );
  AOI22_X1 U18008 ( .A1(n10769), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n14416), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n14377) );
  AOI22_X1 U18009 ( .A1(n10877), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n14503), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n14376) );
  AOI22_X1 U18010 ( .A1(n14504), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10781), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n14375) );
  NAND2_X1 U18011 ( .A1(n14486), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n14374) );
  NAND4_X1 U18012 ( .A1(n14377), .A2(n14376), .A3(n14375), .A4(n14374), .ZN(
        n14378) );
  NOR2_X1 U18013 ( .A1(n14379), .A2(n14378), .ZN(n16376) );
  INV_X1 U18014 ( .A(n16376), .ZN(n14380) );
  AOI22_X1 U18015 ( .A1(n10758), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n14493), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n14388) );
  AOI22_X1 U18016 ( .A1(n10759), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n14477), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n14387) );
  NAND2_X1 U18017 ( .A1(n10732), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n14383) );
  NAND2_X1 U18018 ( .A1(n10733), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n14382) );
  OAI211_X1 U18019 ( .C1(n14497), .C2(n14514), .A(n14383), .B(n14382), .ZN(
        n14384) );
  INV_X1 U18020 ( .A(n14384), .ZN(n14386) );
  AOI22_X1 U18021 ( .A1(n10764), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n14444), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n14385) );
  NAND4_X1 U18022 ( .A1(n14388), .A2(n14387), .A3(n14386), .A4(n14385), .ZN(
        n14394) );
  INV_X1 U18023 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n22054) );
  AOI22_X1 U18024 ( .A1(n10769), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n14416), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n14392) );
  AOI22_X1 U18025 ( .A1(n10877), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n14503), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n14391) );
  AOI22_X1 U18026 ( .A1(n14504), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n10781), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n14390) );
  NAND2_X1 U18027 ( .A1(n14486), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n14389) );
  NAND4_X1 U18028 ( .A1(n14392), .A2(n14391), .A3(n14390), .A4(n14389), .ZN(
        n14393) );
  NOR2_X1 U18029 ( .A1(n14394), .A2(n14393), .ZN(n16372) );
  AOI22_X1 U18030 ( .A1(n10758), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n14493), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n14402) );
  AOI22_X1 U18031 ( .A1(n10759), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n14477), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n14401) );
  INV_X1 U18032 ( .A(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n14397) );
  NAND2_X1 U18033 ( .A1(n10732), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n14396) );
  NAND2_X1 U18034 ( .A1(n10733), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n14395) );
  OAI211_X1 U18035 ( .C1(n9712), .C2(n14397), .A(n14396), .B(n14395), .ZN(
        n14398) );
  INV_X1 U18036 ( .A(n14398), .ZN(n14400) );
  AOI22_X1 U18037 ( .A1(n10764), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n14444), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n14399) );
  NAND4_X1 U18038 ( .A1(n14402), .A2(n14401), .A3(n14400), .A4(n14399), .ZN(
        n14408) );
  AOI22_X1 U18039 ( .A1(n10769), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n14416), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n14406) );
  AOI22_X1 U18040 ( .A1(n10877), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n14503), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n14405) );
  AOI22_X1 U18041 ( .A1(n14504), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n10781), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n14404) );
  NAND2_X1 U18042 ( .A1(n14486), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n14403) );
  NAND4_X1 U18043 ( .A1(n14406), .A2(n14405), .A3(n14404), .A4(n14403), .ZN(
        n14407) );
  OR2_X1 U18044 ( .A1(n14408), .A2(n14407), .ZN(n16366) );
  AOI22_X1 U18045 ( .A1(n10758), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n14493), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n14415) );
  AOI22_X1 U18046 ( .A1(n10759), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n14477), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n14414) );
  NAND2_X1 U18047 ( .A1(n10732), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n14410) );
  NAND2_X1 U18048 ( .A1(n10733), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n14409) );
  OAI211_X1 U18049 ( .C1(n14497), .C2(n14559), .A(n14410), .B(n14409), .ZN(
        n14411) );
  INV_X1 U18050 ( .A(n14411), .ZN(n14413) );
  AOI22_X1 U18051 ( .A1(n10764), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n14444), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n14412) );
  NAND4_X1 U18052 ( .A1(n14415), .A2(n14414), .A3(n14413), .A4(n14412), .ZN(
        n14427) );
  INV_X1 U18053 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n14420) );
  INV_X1 U18054 ( .A(n10769), .ZN(n14419) );
  INV_X1 U18055 ( .A(n14416), .ZN(n14418) );
  INV_X1 U18056 ( .A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n14417) );
  OAI22_X1 U18057 ( .A1(n14420), .A2(n14419), .B1(n14418), .B2(n14417), .ZN(
        n14421) );
  INV_X1 U18058 ( .A(n14421), .ZN(n14425) );
  AOI22_X1 U18059 ( .A1(n10877), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n14503), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n14424) );
  AOI22_X1 U18060 ( .A1(n14504), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n10781), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n14423) );
  NAND2_X1 U18061 ( .A1(n14486), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n14422) );
  NAND4_X1 U18062 ( .A1(n14425), .A2(n14424), .A3(n14423), .A4(n14422), .ZN(
        n14426) );
  AOI22_X1 U18063 ( .A1(n10758), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n14493), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n14434) );
  AOI22_X1 U18064 ( .A1(n10759), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n14477), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n14433) );
  INV_X1 U18065 ( .A(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n14584) );
  NAND2_X1 U18066 ( .A1(n10732), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n14429) );
  NAND2_X1 U18067 ( .A1(n10733), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n14428) );
  OAI211_X1 U18068 ( .C1(n14497), .C2(n14584), .A(n14429), .B(n14428), .ZN(
        n14430) );
  INV_X1 U18069 ( .A(n14430), .ZN(n14432) );
  AOI22_X1 U18070 ( .A1(n10764), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n14444), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n14431) );
  NAND4_X1 U18071 ( .A1(n14434), .A2(n14433), .A3(n14432), .A4(n14431), .ZN(
        n14440) );
  AOI22_X1 U18072 ( .A1(n10769), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n14416), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n14438) );
  AOI22_X1 U18073 ( .A1(n10877), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n14503), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n14437) );
  AOI22_X1 U18074 ( .A1(n14504), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n10781), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n14436) );
  NAND2_X1 U18075 ( .A1(n14486), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n14435) );
  NAND4_X1 U18076 ( .A1(n14438), .A2(n14437), .A3(n14436), .A4(n14435), .ZN(
        n14439) );
  OR2_X1 U18077 ( .A1(n14440), .A2(n14439), .ZN(n16358) );
  AOI22_X1 U18078 ( .A1(n10758), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n14493), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n14448) );
  AOI22_X1 U18079 ( .A1(n10759), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n14477), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n14447) );
  NAND2_X1 U18080 ( .A1(n10732), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n14442) );
  NAND2_X1 U18081 ( .A1(n10733), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n14441) );
  OAI211_X1 U18082 ( .C1(n9712), .C2(n14609), .A(n14442), .B(n14441), .ZN(
        n14443) );
  INV_X1 U18083 ( .A(n14443), .ZN(n14446) );
  AOI22_X1 U18084 ( .A1(n10764), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n14444), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n14445) );
  NAND4_X1 U18085 ( .A1(n14448), .A2(n14447), .A3(n14446), .A4(n14445), .ZN(
        n14454) );
  AOI22_X1 U18086 ( .A1(n10769), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n14416), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n14452) );
  AOI22_X1 U18087 ( .A1(n10877), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n14503), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n14451) );
  AOI22_X1 U18088 ( .A1(n14504), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n10781), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n14450) );
  NAND2_X1 U18089 ( .A1(n14486), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n14449) );
  NAND4_X1 U18090 ( .A1(n14452), .A2(n14451), .A3(n14450), .A4(n14449), .ZN(
        n14453) );
  NOR2_X1 U18091 ( .A1(n14454), .A2(n14453), .ZN(n16353) );
  INV_X1 U18092 ( .A(n16353), .ZN(n14455) );
  AOI22_X1 U18093 ( .A1(n14632), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n14631), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n14467) );
  AOI22_X1 U18094 ( .A1(n14646), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n14665), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n14466) );
  INV_X1 U18095 ( .A(n14458), .ZN(n14661) );
  INV_X1 U18096 ( .A(n14661), .ZN(n14649) );
  AOI22_X1 U18097 ( .A1(n14649), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17147), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n14465) );
  INV_X1 U18098 ( .A(n14664), .ZN(n14654) );
  NAND2_X1 U18099 ( .A1(n14650), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n14461) );
  NAND2_X1 U18100 ( .A1(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n14459) );
  NAND2_X1 U18101 ( .A1(n14460), .A2(n14459), .ZN(n14655) );
  OAI211_X1 U18102 ( .C1(n14654), .C2(n14462), .A(n14461), .B(n14655), .ZN(
        n14463) );
  INV_X1 U18103 ( .A(n14463), .ZN(n14464) );
  NAND4_X1 U18104 ( .A1(n14467), .A2(n14466), .A3(n14465), .A4(n14464), .ZN(
        n14476) );
  AOI22_X1 U18105 ( .A1(n14646), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n14631), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n14474) );
  AOI22_X1 U18106 ( .A1(n14666), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n14650), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n14473) );
  AOI22_X1 U18107 ( .A1(n14649), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17147), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n14472) );
  INV_X1 U18108 ( .A(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n14469) );
  NAND2_X1 U18109 ( .A1(n14665), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n14468) );
  OAI211_X1 U18110 ( .C1(n14469), .C2(n14654), .A(n14468), .B(n14633), .ZN(
        n14470) );
  INV_X1 U18111 ( .A(n14470), .ZN(n14471) );
  NAND4_X1 U18112 ( .A1(n14474), .A2(n14473), .A3(n14472), .A4(n14471), .ZN(
        n14475) );
  NAND2_X1 U18113 ( .A1(n9736), .A2(n14535), .ZN(n14530) );
  AOI22_X1 U18114 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n10759), .B1(
        n14477), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14485) );
  AOI22_X1 U18115 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n14493), .B1(
        n10758), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n14484) );
  INV_X1 U18116 ( .A(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n14480) );
  NAND2_X1 U18117 ( .A1(n10732), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n14479) );
  NAND2_X1 U18118 ( .A1(n10733), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n14478) );
  OAI211_X1 U18119 ( .C1(n14497), .C2(n14480), .A(n14479), .B(n14478), .ZN(
        n14481) );
  INV_X1 U18120 ( .A(n14481), .ZN(n14483) );
  AOI22_X1 U18121 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n10764), .B1(
        n14444), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n14482) );
  NAND4_X1 U18122 ( .A1(n14485), .A2(n14484), .A3(n14483), .A4(n14482), .ZN(
        n14492) );
  AOI22_X1 U18123 ( .A1(n10769), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n14416), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n14490) );
  AOI22_X1 U18124 ( .A1(n10877), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n14503), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n14489) );
  AOI22_X1 U18125 ( .A1(n14504), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n10781), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n14488) );
  NAND2_X1 U18126 ( .A1(n14486), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n14487) );
  NAND4_X1 U18127 ( .A1(n14490), .A2(n14489), .A3(n14488), .A4(n14487), .ZN(
        n14491) );
  XNOR2_X1 U18128 ( .A(n14530), .B(n14538), .ZN(n14511) );
  AOI22_X1 U18129 ( .A1(n10758), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n14493), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n14502) );
  AOI22_X1 U18130 ( .A1(n10759), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n14477), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n14501) );
  NAND2_X1 U18131 ( .A1(n10732), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n14495) );
  NAND2_X1 U18132 ( .A1(n10733), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n14494) );
  OAI211_X1 U18133 ( .C1(n14497), .C2(n14496), .A(n14495), .B(n14494), .ZN(
        n14498) );
  INV_X1 U18134 ( .A(n14498), .ZN(n14500) );
  AOI22_X1 U18135 ( .A1(n10764), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n14444), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n14499) );
  NAND4_X1 U18136 ( .A1(n14502), .A2(n14501), .A3(n14500), .A4(n14499), .ZN(
        n14510) );
  AOI22_X1 U18137 ( .A1(n10769), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n14416), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n14508) );
  AOI22_X1 U18138 ( .A1(n10877), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n14503), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n14507) );
  AOI22_X1 U18139 ( .A1(n14504), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n10781), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n14506) );
  NAND2_X1 U18140 ( .A1(n14486), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n14505) );
  NAND4_X1 U18141 ( .A1(n14508), .A2(n14507), .A3(n14506), .A4(n14505), .ZN(
        n14509) );
  NAND2_X1 U18142 ( .A1(n14511), .A2(n16349), .ZN(n14512) );
  INV_X1 U18143 ( .A(n14511), .ZN(n16344) );
  NAND2_X1 U18144 ( .A1(n9735), .A2(n14535), .ZN(n16343) );
  NAND2_X1 U18145 ( .A1(n14538), .A2(n14535), .ZN(n14529) );
  AOI22_X1 U18146 ( .A1(n14646), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n14631), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n14519) );
  AOI22_X1 U18147 ( .A1(n14632), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n14665), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n14518) );
  AOI22_X1 U18148 ( .A1(n14649), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17147), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n14517) );
  NAND2_X1 U18149 ( .A1(n14650), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n14513) );
  OAI211_X1 U18150 ( .C1(n14654), .C2(n14514), .A(n14513), .B(n14655), .ZN(
        n14515) );
  INV_X1 U18151 ( .A(n14515), .ZN(n14516) );
  NAND4_X1 U18152 ( .A1(n14519), .A2(n14518), .A3(n14517), .A4(n14516), .ZN(
        n14528) );
  AOI22_X1 U18153 ( .A1(n14646), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n14631), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n14526) );
  AOI22_X1 U18154 ( .A1(n14632), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n14665), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n14525) );
  AOI22_X1 U18155 ( .A1(n14649), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n17147), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n14524) );
  NAND2_X1 U18156 ( .A1(n14650), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n14520) );
  OAI211_X1 U18157 ( .C1(n14521), .C2(n14654), .A(n14520), .B(n14633), .ZN(
        n14522) );
  INV_X1 U18158 ( .A(n14522), .ZN(n14523) );
  NAND4_X1 U18159 ( .A1(n14526), .A2(n14525), .A3(n14524), .A4(n14523), .ZN(
        n14527) );
  NAND2_X1 U18160 ( .A1(n14528), .A2(n14527), .ZN(n14536) );
  OAI21_X1 U18161 ( .B1(n14578), .B2(n14529), .A(n14536), .ZN(n14534) );
  INV_X1 U18162 ( .A(n14530), .ZN(n14532) );
  INV_X1 U18163 ( .A(n14536), .ZN(n14531) );
  NAND3_X1 U18164 ( .A1(n14532), .A2(n14531), .A3(n14538), .ZN(n14533) );
  AND2_X1 U18165 ( .A1(n14534), .A2(n14533), .ZN(n16338) );
  INV_X1 U18166 ( .A(n14535), .ZN(n14537) );
  NOR2_X1 U18167 ( .A1(n14537), .A2(n14536), .ZN(n14539) );
  AND2_X1 U18168 ( .A1(n14539), .A2(n14538), .ZN(n14556) );
  AOI22_X1 U18169 ( .A1(n14646), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n14565), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n14546) );
  AOI22_X1 U18170 ( .A1(n14632), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n14665), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n14545) );
  AOI22_X1 U18171 ( .A1(n14649), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n9733), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n14544) );
  INV_X1 U18172 ( .A(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n14541) );
  NAND2_X1 U18173 ( .A1(n14650), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n14540) );
  OAI211_X1 U18174 ( .C1(n14659), .C2(n14541), .A(n14540), .B(n14655), .ZN(
        n14542) );
  INV_X1 U18175 ( .A(n14542), .ZN(n14543) );
  NAND4_X1 U18176 ( .A1(n14546), .A2(n14545), .A3(n14544), .A4(n14543), .ZN(
        n14555) );
  AOI22_X1 U18177 ( .A1(n14646), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n14666), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n14553) );
  AOI22_X1 U18178 ( .A1(n14631), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n14665), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n14552) );
  AOI22_X1 U18179 ( .A1(n14649), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17147), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n14551) );
  INV_X1 U18180 ( .A(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n14548) );
  NAND2_X1 U18181 ( .A1(n14650), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n14547) );
  OAI211_X1 U18182 ( .C1(n14548), .C2(n14654), .A(n14547), .B(n14633), .ZN(
        n14549) );
  INV_X1 U18183 ( .A(n14549), .ZN(n14550) );
  NAND4_X1 U18184 ( .A1(n14553), .A2(n14552), .A3(n14551), .A4(n14550), .ZN(
        n14554) );
  AND2_X1 U18185 ( .A1(n14555), .A2(n14554), .ZN(n14557) );
  NAND2_X1 U18186 ( .A1(n14556), .A2(n14557), .ZN(n14582) );
  OAI211_X1 U18187 ( .C1(n14556), .C2(n14557), .A(n14599), .B(n14582), .ZN(
        n14576) );
  NAND2_X1 U18188 ( .A1(n9735), .A2(n14557), .ZN(n16333) );
  AOI22_X1 U18189 ( .A1(n14646), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n14631), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n14564) );
  AOI22_X1 U18190 ( .A1(n14632), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n14665), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n14563) );
  AOI22_X1 U18191 ( .A1(n14649), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17147), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n14562) );
  NAND2_X1 U18192 ( .A1(n14650), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n14558) );
  OAI211_X1 U18193 ( .C1(n14654), .C2(n14559), .A(n14558), .B(n14655), .ZN(
        n14560) );
  INV_X1 U18194 ( .A(n14560), .ZN(n14561) );
  NAND4_X1 U18195 ( .A1(n14564), .A2(n14563), .A3(n14562), .A4(n14561), .ZN(
        n14574) );
  AOI22_X1 U18196 ( .A1(n14646), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n14565), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n14572) );
  AOI22_X1 U18197 ( .A1(n14632), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n14665), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n14571) );
  AOI22_X1 U18198 ( .A1(n14649), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17147), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n14570) );
  NAND2_X1 U18199 ( .A1(n14650), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n14566) );
  OAI211_X1 U18200 ( .C1(n14567), .C2(n14654), .A(n14566), .B(n14633), .ZN(
        n14568) );
  INV_X1 U18201 ( .A(n14568), .ZN(n14569) );
  NAND4_X1 U18202 ( .A1(n14572), .A2(n14571), .A3(n14570), .A4(n14569), .ZN(
        n14573) );
  NAND2_X1 U18203 ( .A1(n14574), .A2(n14573), .ZN(n16325) );
  OR2_X1 U18204 ( .A1(n16333), .A2(n16325), .ZN(n14575) );
  NOR2_X1 U18205 ( .A1(n16322), .A2(n14575), .ZN(n14581) );
  INV_X1 U18206 ( .A(n14582), .ZN(n14577) );
  XOR2_X1 U18207 ( .A(n16325), .B(n14577), .Z(n14579) );
  NOR2_X1 U18208 ( .A1(n14579), .A2(n14578), .ZN(n16327) );
  NOR2_X1 U18209 ( .A1(n14581), .A2(n14580), .ZN(n14602) );
  NOR2_X1 U18210 ( .A1(n14582), .A2(n16325), .ZN(n14600) );
  AOI22_X1 U18211 ( .A1(n14646), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n14631), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n14589) );
  AOI22_X1 U18212 ( .A1(n14632), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n14665), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n14588) );
  AOI22_X1 U18213 ( .A1(n14649), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17147), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n14587) );
  NAND2_X1 U18214 ( .A1(n14650), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n14583) );
  OAI211_X1 U18215 ( .C1(n14654), .C2(n14584), .A(n14583), .B(n14655), .ZN(
        n14585) );
  INV_X1 U18216 ( .A(n14585), .ZN(n14586) );
  NAND4_X1 U18217 ( .A1(n14589), .A2(n14588), .A3(n14587), .A4(n14586), .ZN(
        n14598) );
  AOI22_X1 U18218 ( .A1(n14646), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n14631), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n14596) );
  AOI22_X1 U18219 ( .A1(n14632), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n14665), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n14595) );
  AOI22_X1 U18220 ( .A1(n14649), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17147), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n14594) );
  INV_X1 U18221 ( .A(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n14591) );
  NAND2_X1 U18222 ( .A1(n14650), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n14590) );
  OAI211_X1 U18223 ( .C1(n14591), .C2(n14654), .A(n14590), .B(n14633), .ZN(
        n14592) );
  INV_X1 U18224 ( .A(n14592), .ZN(n14593) );
  NAND4_X1 U18225 ( .A1(n14596), .A2(n14595), .A3(n14594), .A4(n14593), .ZN(
        n14597) );
  AND2_X1 U18226 ( .A1(n14598), .A2(n14597), .ZN(n14604) );
  NAND2_X1 U18227 ( .A1(n14600), .A2(n14604), .ZN(n16311) );
  OAI211_X1 U18228 ( .C1(n14600), .C2(n14604), .A(n16311), .B(n14599), .ZN(
        n14601) );
  NAND2_X1 U18229 ( .A1(n14602), .A2(n14601), .ZN(n14603) );
  INV_X1 U18230 ( .A(n14604), .ZN(n14605) );
  NOR2_X1 U18231 ( .A1(n9736), .A2(n14605), .ZN(n16319) );
  AOI22_X1 U18232 ( .A1(n14646), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n14631), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n14614) );
  AOI22_X1 U18233 ( .A1(n14632), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n14665), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n14613) );
  AOI22_X1 U18234 ( .A1(n14649), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17147), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n14612) );
  NAND2_X1 U18235 ( .A1(n14650), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n14608) );
  OAI211_X1 U18236 ( .C1(n14654), .C2(n14609), .A(n14608), .B(n14655), .ZN(
        n14610) );
  INV_X1 U18237 ( .A(n14610), .ZN(n14611) );
  NAND4_X1 U18238 ( .A1(n14614), .A2(n14613), .A3(n14612), .A4(n14611), .ZN(
        n14623) );
  AOI22_X1 U18239 ( .A1(n14646), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n14631), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n14621) );
  AOI22_X1 U18240 ( .A1(n14632), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n14665), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n14620) );
  AOI22_X1 U18241 ( .A1(n14649), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17147), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n14619) );
  NAND2_X1 U18242 ( .A1(n14650), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n14615) );
  OAI211_X1 U18243 ( .C1(n14616), .C2(n14654), .A(n14615), .B(n14633), .ZN(
        n14617) );
  INV_X1 U18244 ( .A(n14617), .ZN(n14618) );
  NAND4_X1 U18245 ( .A1(n14621), .A2(n14620), .A3(n14619), .A4(n14618), .ZN(
        n14622) );
  NAND2_X1 U18246 ( .A1(n14623), .A2(n14622), .ZN(n16314) );
  AOI22_X1 U18247 ( .A1(n14632), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n14631), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n14630) );
  AOI22_X1 U18248 ( .A1(n9730), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n14665), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n14629) );
  AOI22_X1 U18249 ( .A1(n9733), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17147), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n14628) );
  NAND2_X1 U18250 ( .A1(n14650), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n14624) );
  OAI211_X1 U18251 ( .C1(n14661), .C2(n14625), .A(n14624), .B(n14655), .ZN(
        n14626) );
  INV_X1 U18252 ( .A(n14626), .ZN(n14627) );
  NAND4_X1 U18253 ( .A1(n14630), .A2(n14629), .A3(n14628), .A4(n14627), .ZN(
        n14642) );
  AOI22_X1 U18254 ( .A1(n14646), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n14631), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n14640) );
  AOI22_X1 U18255 ( .A1(n14632), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n14665), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n14639) );
  AOI22_X1 U18256 ( .A1(n14649), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17147), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n14638) );
  NAND2_X1 U18257 ( .A1(n14650), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n14634) );
  OAI211_X1 U18258 ( .C1(n14635), .C2(n14654), .A(n14634), .B(n14633), .ZN(
        n14636) );
  INV_X1 U18259 ( .A(n14636), .ZN(n14637) );
  NAND4_X1 U18260 ( .A1(n14640), .A2(n14639), .A3(n14638), .A4(n14637), .ZN(
        n14641) );
  NAND2_X1 U18261 ( .A1(n14642), .A2(n14641), .ZN(n14644) );
  OR3_X1 U18262 ( .A1(n16311), .A2(n9735), .A3(n16314), .ZN(n14643) );
  NOR2_X1 U18263 ( .A1(n14643), .A2(n14644), .ZN(n14645) );
  AOI21_X1 U18264 ( .B1(n14644), .B2(n14643), .A(n14645), .ZN(n16307) );
  NOR2_X1 U18265 ( .A1(n16398), .A2(n14645), .ZN(n14674) );
  AOI22_X1 U18266 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n14631), .B1(
        n14666), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n14648) );
  AOI22_X1 U18267 ( .A1(n14646), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n14665), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n14647) );
  NAND2_X1 U18268 ( .A1(n14648), .A2(n14647), .ZN(n14672) );
  INV_X1 U18269 ( .A(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n14653) );
  AOI22_X1 U18270 ( .A1(n14649), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17147), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n14652) );
  AOI21_X1 U18271 ( .B1(n14650), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A(
        n14655), .ZN(n14651) );
  OAI211_X1 U18272 ( .C1(n14654), .C2(n14653), .A(n14652), .B(n14651), .ZN(
        n14671) );
  OAI21_X1 U18273 ( .B1(n14657), .B2(n14656), .A(n14655), .ZN(n14663) );
  INV_X1 U18274 ( .A(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n14660) );
  INV_X1 U18275 ( .A(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n14658) );
  OAI22_X1 U18276 ( .A1(n14661), .A2(n14660), .B1(n14659), .B2(n14658), .ZN(
        n14662) );
  AOI211_X1 U18277 ( .C1(n9733), .C2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A(
        n14663), .B(n14662), .ZN(n14669) );
  AOI22_X1 U18278 ( .A1(n14631), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n14665), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n14668) );
  AOI22_X1 U18279 ( .A1(n9730), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n14666), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n14667) );
  NAND3_X1 U18280 ( .A1(n14669), .A2(n14668), .A3(n14667), .ZN(n14670) );
  OAI21_X1 U18281 ( .B1(n14672), .B2(n14671), .A(n14670), .ZN(n14673) );
  XNOR2_X1 U18282 ( .A(n14674), .B(n14673), .ZN(n14683) );
  NOR2_X1 U18283 ( .A1(n14741), .A2(n16386), .ZN(n14675) );
  AOI21_X1 U18284 ( .B1(P2_EBX_REG_30__SCAN_IN), .B2(n16386), .A(n14675), .ZN(
        n14676) );
  OAI21_X1 U18285 ( .B1(n14683), .B2(n16388), .A(n14676), .ZN(P2_U2857) );
  INV_X1 U18286 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n15199) );
  NAND2_X1 U18287 ( .A1(n16490), .A2(BUF2_REG_30__SCAN_IN), .ZN(n14679) );
  AOI22_X1 U18288 ( .A1(n16492), .A2(n20349), .B1(P2_EAX_REG_30__SCAN_IN), 
        .B2(n20303), .ZN(n14678) );
  OAI211_X1 U18289 ( .C1(n16495), .C2(n15199), .A(n14679), .B(n14678), .ZN(
        n14680) );
  AOI21_X1 U18290 ( .B1(n14681), .B2(n20304), .A(n14680), .ZN(n14682) );
  OAI21_X1 U18291 ( .B1(n14683), .B2(n20298), .A(n14682), .ZN(P2_U2889) );
  INV_X1 U18292 ( .A(n14684), .ZN(n16272) );
  OR2_X1 U18293 ( .A1(n14686), .A2(n14685), .ZN(n14687) );
  NAND2_X1 U18294 ( .A1(n14688), .A2(n14687), .ZN(n14706) );
  INV_X1 U18295 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n14689) );
  OR2_X1 U18296 ( .A1(n17736), .A2(n14689), .ZN(n14691) );
  INV_X1 U18297 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n21034) );
  NOR2_X1 U18298 ( .A1(n20217), .A2(n21034), .ZN(n14702) );
  INV_X1 U18299 ( .A(n14702), .ZN(n14690) );
  OAI211_X1 U18300 ( .C1(n16762), .C2(n14706), .A(n14691), .B(n14690), .ZN(
        n14692) );
  AOI21_X1 U18301 ( .B1(n17725), .B2(n16272), .A(n14692), .ZN(n14695) );
  OR2_X1 U18302 ( .A1(n14693), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n14710) );
  NAND3_X1 U18303 ( .A1(n14710), .A2(n11457), .A3(n14711), .ZN(n14694) );
  OAI211_X1 U18304 ( .C1(n14714), .C2(n20363), .A(n14695), .B(n14694), .ZN(
        P2_U3012) );
  AND2_X1 U18305 ( .A1(n14697), .A2(n14696), .ZN(n14708) );
  OR2_X1 U18306 ( .A1(n14699), .A2(n14698), .ZN(n14700) );
  NAND2_X1 U18307 ( .A1(n14701), .A2(n14700), .ZN(n21104) );
  AOI21_X1 U18308 ( .B1(n17741), .B2(n21104), .A(n14702), .ZN(n14705) );
  OAI21_X1 U18309 ( .B1(n14703), .B2(n17069), .A(n17070), .ZN(n14704) );
  OAI211_X1 U18310 ( .C1(n14706), .C2(n17082), .A(n14705), .B(n14704), .ZN(
        n14707) );
  AOI211_X1 U18311 ( .C1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .C2(n14709), .A(
        n14708), .B(n14707), .ZN(n14713) );
  NAND3_X1 U18312 ( .A1(n17748), .A2(n14711), .A3(n14710), .ZN(n14712) );
  OAI211_X1 U18313 ( .C1(n17745), .C2(n14714), .A(n14713), .B(n14712), .ZN(
        P2_U3044) );
  INV_X1 U18314 ( .A(n14715), .ZN(n14722) );
  INV_X1 U18315 ( .A(n16103), .ZN(n14718) );
  AOI21_X1 U18316 ( .B1(n20356), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n14716), .ZN(n14717) );
  INV_X1 U18317 ( .A(n14719), .ZN(n14720) );
  OAI21_X1 U18318 ( .B1(n14724), .B2(n16737), .A(n14723), .ZN(P2_U2983) );
  AOI21_X1 U18319 ( .B1(n15955), .B2(n14726), .A(n14725), .ZN(n16397) );
  INV_X1 U18320 ( .A(n14727), .ZN(n16778) );
  INV_X1 U18321 ( .A(n16764), .ZN(n14728) );
  NAND2_X1 U18322 ( .A1(n14728), .A2(n16777), .ZN(n16776) );
  NAND2_X1 U18323 ( .A1(n16778), .A2(n16776), .ZN(n16767) );
  AOI21_X1 U18324 ( .B1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n14730), .A(
        n22042), .ZN(n14729) );
  AOI211_X1 U18325 ( .C1(n14730), .C2(n22042), .A(n14729), .B(n16764), .ZN(
        n14731) );
  AOI211_X1 U18326 ( .C1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n16767), .A(
        n14732), .B(n14731), .ZN(n14733) );
  INV_X1 U18327 ( .A(n14736), .ZN(n14743) );
  AOI21_X1 U18328 ( .B1(n20356), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n14737), .ZN(n14738) );
  OAI21_X1 U18329 ( .B1(n15928), .B2(n20368), .A(n14738), .ZN(n14739) );
  INV_X1 U18330 ( .A(n14739), .ZN(n14740) );
  AOI21_X1 U18331 ( .B1(n20357), .B2(n14743), .A(n14742), .ZN(n14744) );
  OAI21_X1 U18332 ( .B1(n14745), .B2(n16737), .A(n14744), .ZN(P2_U2984) );
  INV_X1 U18333 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n17837) );
  NAND2_X1 U18334 ( .A1(n14747), .A2(n14746), .ZN(n14750) );
  AOI22_X1 U18335 ( .A1(n15281), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n15291), .ZN(n14749) );
  OAI211_X1 U18336 ( .C1(n15274), .C2(n17837), .A(n14750), .B(n14749), .ZN(
        P1_U2873) );
  NOR2_X1 U18337 ( .A1(n17070), .A2(n17738), .ZN(n14752) );
  OR2_X1 U18338 ( .A1(n16911), .A2(n14752), .ZN(n14759) );
  NAND2_X1 U18339 ( .A1(n16989), .A2(n14753), .ZN(n14754) );
  NAND2_X1 U18340 ( .A1(n16993), .A2(n14754), .ZN(n16978) );
  AND2_X1 U18341 ( .A1(n17111), .A2(n14761), .ZN(n14755) );
  INV_X1 U18342 ( .A(n14756), .ZN(n17019) );
  AND2_X1 U18343 ( .A1(n17019), .A2(n16924), .ZN(n14757) );
  NOR2_X1 U18344 ( .A1(n16926), .A2(n14757), .ZN(n14758) );
  NAND2_X1 U18345 ( .A1(n16989), .A2(n14760), .ZN(n16938) );
  OAI22_X1 U18346 ( .A1(n16643), .A2(n17082), .B1(n16924), .B2(n16892), .ZN(
        n14771) );
  OAI21_X1 U18347 ( .B1(n9766), .B2(n14763), .A(n14762), .ZN(n16642) );
  OR2_X1 U18348 ( .A1(n14352), .A2(n14764), .ZN(n14765) );
  AND2_X1 U18349 ( .A1(n9792), .A2(n14765), .ZN(n16639) );
  NOR2_X1 U18350 ( .A1(n16730), .A2(n21056), .ZN(n16636) );
  OAI21_X1 U18351 ( .B1(n14359), .B2(n14767), .A(n14766), .ZN(n20224) );
  NOR2_X1 U18352 ( .A1(n20224), .A2(n17105), .ZN(n14768) );
  AOI211_X1 U18353 ( .C1(n17076), .C2(n16639), .A(n16636), .B(n14768), .ZN(
        n14769) );
  OAI21_X1 U18354 ( .B1(n16642), .B2(n17101), .A(n14769), .ZN(n14770) );
  AOI21_X1 U18355 ( .B1(n14771), .B2(n14773), .A(n14770), .ZN(n14772) );
  OAI21_X1 U18356 ( .B1(n16907), .B2(n14773), .A(n14772), .ZN(P2_U3030) );
  INV_X1 U18357 ( .A(n14774), .ZN(n14775) );
  MUX2_X1 U18358 ( .A(n14776), .B(n14775), .S(n17629), .Z(n14782) );
  INV_X1 U18359 ( .A(n14777), .ZN(n14778) );
  NOR2_X1 U18360 ( .A1(n14779), .A2(n14778), .ZN(n14780) );
  AOI21_X1 U18361 ( .B1(n17629), .B2(n13490), .A(n14780), .ZN(n14781) );
  NAND2_X1 U18362 ( .A1(n14782), .A2(n14781), .ZN(n17612) );
  INV_X1 U18363 ( .A(n14783), .ZN(n14784) );
  AOI22_X1 U18364 ( .A1(n17629), .A2(n15091), .B1(n14785), .B2(n14784), .ZN(
        n21145) );
  NAND3_X1 U18365 ( .A1(n14786), .A2(n15091), .A3(n15925), .ZN(n14787) );
  NAND2_X1 U18366 ( .A1(n14787), .A2(n21912), .ZN(n21904) );
  NAND2_X1 U18367 ( .A1(n21145), .A2(n21904), .ZN(n17610) );
  AND2_X1 U18368 ( .A1(n17610), .A2(n14788), .ZN(n21154) );
  MUX2_X1 U18369 ( .A(P1_MORE_REG_SCAN_IN), .B(n17612), .S(n21154), .Z(
        P1_U3484) );
  INV_X1 U18370 ( .A(n14790), .ZN(n14791) );
  NAND2_X1 U18371 ( .A1(n14824), .A2(n14791), .ZN(n14792) );
  OAI21_X1 U18372 ( .B1(n14814), .B2(n14793), .A(n14792), .ZN(n14796) );
  INV_X1 U18373 ( .A(n14794), .ZN(n14795) );
  XNOR2_X1 U18374 ( .A(n14796), .B(n14795), .ZN(n15589) );
  INV_X1 U18375 ( .A(n14797), .ZN(n14798) );
  AOI22_X1 U18376 ( .A1(n21223), .A2(P1_EBX_REG_30__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n21233), .ZN(n14804) );
  NOR2_X1 U18377 ( .A1(n14977), .A2(n14800), .ZN(n14802) );
  OAI21_X1 U18378 ( .B1(n14802), .B2(P1_REIP_REG_30__SCAN_IN), .A(n14801), 
        .ZN(n14803) );
  OAI211_X1 U18379 ( .C1(n21263), .C2(n15361), .A(n14804), .B(n14803), .ZN(
        n14805) );
  AOI21_X1 U18380 ( .B1(n15589), .B2(n21259), .A(n14805), .ZN(n14806) );
  OAI21_X1 U18381 ( .B1(n15202), .B2(n17648), .A(n14806), .ZN(P1_U2810) );
  INV_X1 U18382 ( .A(n21170), .ZN(n21249) );
  AOI21_X1 U18383 ( .B1(n21251), .B2(n14810), .A(n21249), .ZN(n14826) );
  AOI22_X1 U18384 ( .A1(n21223), .A2(P1_EBX_REG_29__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n21233), .ZN(n14813) );
  NAND3_X1 U18385 ( .A1(n21251), .A2(n14811), .A3(n22188), .ZN(n14812) );
  OAI211_X1 U18386 ( .C1(n14826), .C2(n22188), .A(n14813), .B(n14812), .ZN(
        n14819) );
  OR2_X1 U18387 ( .A1(n14824), .A2(n14815), .ZN(n14816) );
  AOI211_X1 U18388 ( .C1(n21174), .C2(n15364), .A(n14819), .B(n14818), .ZN(
        n14820) );
  OAI21_X1 U18389 ( .B1(n15372), .B2(n17648), .A(n14820), .ZN(P1_U2811) );
  AOI21_X1 U18390 ( .B1(n14823), .B2(n14822), .A(n14807), .ZN(n15378) );
  INV_X1 U18391 ( .A(n15378), .ZN(n15214) );
  AOI21_X1 U18392 ( .B1(n14825), .B2(n14843), .A(n14824), .ZN(n15603) );
  AOI22_X1 U18393 ( .A1(n21223), .A2(P1_EBX_REG_28__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n21233), .ZN(n14830) );
  NOR3_X1 U18394 ( .A1(n14977), .A2(n21888), .A3(n14837), .ZN(n14828) );
  INV_X1 U18395 ( .A(n14826), .ZN(n14827) );
  OAI21_X1 U18396 ( .B1(n14828), .B2(P1_REIP_REG_28__SCAN_IN), .A(n14827), 
        .ZN(n14829) );
  OAI211_X1 U18397 ( .C1(n21263), .C2(n15376), .A(n14830), .B(n14829), .ZN(
        n14831) );
  AOI21_X1 U18398 ( .B1(n15603), .B2(n21259), .A(n14831), .ZN(n14832) );
  OAI21_X1 U18399 ( .B1(n15214), .B2(n17648), .A(n14832), .ZN(P1_U2812) );
  OAI21_X1 U18400 ( .B1(n14833), .B2(n14834), .A(n14822), .ZN(n15389) );
  INV_X1 U18401 ( .A(n14837), .ZN(n14835) );
  NAND2_X1 U18402 ( .A1(n21170), .A2(n14835), .ZN(n14836) );
  NAND2_X1 U18403 ( .A1(n21217), .A2(n14836), .ZN(n14858) );
  AOI22_X1 U18404 ( .A1(n21223), .A2(P1_EBX_REG_27__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n21233), .ZN(n14839) );
  OR3_X1 U18405 ( .A1(n14977), .A2(P1_REIP_REG_27__SCAN_IN), .A3(n14837), .ZN(
        n14838) );
  OAI211_X1 U18406 ( .C1(n14858), .C2(n21888), .A(n14839), .B(n14838), .ZN(
        n14845) );
  NAND2_X1 U18407 ( .A1(n14840), .A2(n14841), .ZN(n14842) );
  NAND2_X1 U18408 ( .A1(n14843), .A2(n14842), .ZN(n15615) );
  NOR2_X1 U18409 ( .A1(n15615), .A2(n17647), .ZN(n14844) );
  AOI211_X1 U18410 ( .C1(n21174), .C2(n15380), .A(n14845), .B(n14844), .ZN(
        n14846) );
  OAI21_X1 U18411 ( .B1(n15389), .B2(n17648), .A(n14846), .ZN(P1_U2813) );
  OR2_X1 U18412 ( .A1(n14847), .A2(n14848), .ZN(n14849) );
  NAND2_X1 U18413 ( .A1(n14840), .A2(n14849), .ZN(n15619) );
  AOI21_X1 U18414 ( .B1(n14852), .B2(n14851), .A(n14833), .ZN(n15397) );
  NAND2_X1 U18415 ( .A1(n15397), .A2(n21212), .ZN(n14862) );
  INV_X1 U18416 ( .A(n15395), .ZN(n14860) );
  AOI21_X1 U18417 ( .B1(n21251), .B2(n14853), .A(P1_REIP_REG_26__SCAN_IN), 
        .ZN(n14857) );
  INV_X1 U18418 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n22185) );
  OAI22_X1 U18419 ( .A1(n21256), .A2(n22185), .B1(n14854), .B2(n21253), .ZN(
        n14855) );
  INV_X1 U18420 ( .A(n14855), .ZN(n14856) );
  OAI21_X1 U18421 ( .B1(n14858), .B2(n14857), .A(n14856), .ZN(n14859) );
  AOI21_X1 U18422 ( .B1(n21174), .B2(n14860), .A(n14859), .ZN(n14861) );
  OAI211_X1 U18423 ( .C1(n15619), .C2(n17647), .A(n14862), .B(n14861), .ZN(
        P1_U2814) );
  NOR2_X1 U18424 ( .A1(n14863), .A2(n14864), .ZN(n14865) );
  OR2_X1 U18425 ( .A1(n14847), .A2(n14865), .ZN(n15634) );
  OAI21_X1 U18426 ( .B1(n14866), .B2(n14867), .A(n14851), .ZN(n15406) );
  INV_X1 U18427 ( .A(n15406), .ZN(n14868) );
  NAND2_X1 U18428 ( .A1(n14868), .A2(n21212), .ZN(n14878) );
  NAND2_X1 U18429 ( .A1(n21251), .A2(n14884), .ZN(n14869) );
  NAND2_X1 U18430 ( .A1(n14869), .A2(n21170), .ZN(n14892) );
  NAND2_X1 U18431 ( .A1(n14892), .A2(P1_REIP_REG_25__SCAN_IN), .ZN(n14875) );
  OAI22_X1 U18432 ( .A1(n21256), .A2(n22121), .B1(n15399), .B2(n21253), .ZN(
        n14870) );
  INV_X1 U18433 ( .A(n14870), .ZN(n14874) );
  NAND2_X1 U18434 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(P1_REIP_REG_25__SCAN_IN), 
        .ZN(n14871) );
  OAI211_X1 U18435 ( .C1(P1_REIP_REG_25__SCAN_IN), .C2(n14872), .A(n21251), 
        .B(n14871), .ZN(n14873) );
  NAND3_X1 U18436 ( .A1(n14875), .A2(n14874), .A3(n14873), .ZN(n14876) );
  AOI21_X1 U18437 ( .B1(n21174), .B2(n15401), .A(n14876), .ZN(n14877) );
  OAI211_X1 U18438 ( .C1(n17647), .C2(n15634), .A(n14878), .B(n14877), .ZN(
        P1_U2815) );
  AOI21_X1 U18439 ( .B1(n14880), .B2(n14879), .A(n14866), .ZN(n15412) );
  INV_X1 U18440 ( .A(n15412), .ZN(n15237) );
  AOI21_X1 U18441 ( .B1(n14881), .B2(n9788), .A(n14863), .ZN(n15642) );
  OAI22_X1 U18442 ( .A1(n21256), .A2(n14883), .B1(n14882), .B2(n21253), .ZN(
        n14886) );
  NOR3_X1 U18443 ( .A1(n14977), .A2(P1_REIP_REG_24__SCAN_IN), .A3(n14884), 
        .ZN(n14885) );
  AOI211_X1 U18444 ( .C1(P1_REIP_REG_24__SCAN_IN), .C2(n14892), .A(n14886), 
        .B(n14885), .ZN(n14887) );
  OAI21_X1 U18445 ( .B1(n21263), .B2(n15410), .A(n14887), .ZN(n14888) );
  AOI21_X1 U18446 ( .B1(n15642), .B2(n21259), .A(n14888), .ZN(n14889) );
  OAI21_X1 U18447 ( .B1(n15237), .B2(n17648), .A(n14889), .ZN(P1_U2816) );
  OAI21_X1 U18448 ( .B1(n14890), .B2(n14891), .A(n14879), .ZN(n15417) );
  INV_X1 U18449 ( .A(n14892), .ZN(n14896) );
  AOI21_X1 U18450 ( .B1(n21251), .B2(n14893), .A(P1_REIP_REG_23__SCAN_IN), 
        .ZN(n14895) );
  AOI22_X1 U18451 ( .A1(n21223), .A2(P1_EBX_REG_23__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n21233), .ZN(n14894) );
  OAI21_X1 U18452 ( .B1(n14896), .B2(n14895), .A(n14894), .ZN(n14900) );
  NAND2_X1 U18453 ( .A1(n14904), .A2(n14897), .ZN(n14898) );
  NAND2_X1 U18454 ( .A1(n9788), .A2(n14898), .ZN(n15646) );
  NOR2_X1 U18455 ( .A1(n15646), .A2(n17647), .ZN(n14899) );
  AOI211_X1 U18456 ( .C1(n21174), .C2(n15420), .A(n14900), .B(n14899), .ZN(
        n14901) );
  OAI21_X1 U18457 ( .B1(n15417), .B2(n17648), .A(n14901), .ZN(P1_U2817) );
  OR2_X1 U18458 ( .A1(n14928), .A2(n14902), .ZN(n14903) );
  NAND2_X1 U18459 ( .A1(n14904), .A2(n14903), .ZN(n15662) );
  AOI21_X1 U18460 ( .B1(n14907), .B2(n14906), .A(n14890), .ZN(n15430) );
  NAND2_X1 U18461 ( .A1(n15430), .A2(n21212), .ZN(n14918) );
  INV_X1 U18462 ( .A(n15426), .ZN(n14916) );
  INV_X1 U18463 ( .A(n14908), .ZN(n14922) );
  NAND2_X1 U18464 ( .A1(n21170), .A2(n14922), .ZN(n14909) );
  NAND2_X1 U18465 ( .A1(n21217), .A2(n14909), .ZN(n14938) );
  INV_X1 U18466 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n15427) );
  OAI22_X1 U18467 ( .A1(n21256), .A2(n15126), .B1(n21959), .B2(n21253), .ZN(
        n14910) );
  INV_X1 U18468 ( .A(n14910), .ZN(n14914) );
  NAND2_X1 U18469 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(P1_REIP_REG_22__SCAN_IN), 
        .ZN(n14911) );
  OAI211_X1 U18470 ( .C1(P1_REIP_REG_22__SCAN_IN), .C2(n14912), .A(n21251), 
        .B(n14911), .ZN(n14913) );
  OAI211_X1 U18471 ( .C1(n14938), .C2(n15427), .A(n14914), .B(n14913), .ZN(
        n14915) );
  AOI21_X1 U18472 ( .B1(n21174), .B2(n14916), .A(n14915), .ZN(n14917) );
  OAI211_X1 U18473 ( .C1(n15662), .C2(n17647), .A(n14918), .B(n14917), .ZN(
        P1_U2818) );
  OAI21_X1 U18474 ( .B1(n14920), .B2(n14921), .A(n14906), .ZN(n15440) );
  AOI22_X1 U18475 ( .A1(n21223), .A2(P1_EBX_REG_21__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n21233), .ZN(n14924) );
  NAND3_X1 U18476 ( .A1(n21251), .A2(n14922), .A3(n21882), .ZN(n14923) );
  OAI211_X1 U18477 ( .C1(n14938), .C2(n21882), .A(n14924), .B(n14923), .ZN(
        n14925) );
  AOI21_X1 U18478 ( .B1(n21174), .B2(n15434), .A(n14925), .ZN(n14930) );
  AND2_X1 U18479 ( .A1(n14933), .A2(n14926), .ZN(n14927) );
  NOR2_X1 U18480 ( .A1(n14928), .A2(n14927), .ZN(n15666) );
  NAND2_X1 U18481 ( .A1(n15666), .A2(n21259), .ZN(n14929) );
  OAI211_X1 U18482 ( .C1(n15440), .C2(n17648), .A(n14930), .B(n14929), .ZN(
        P1_U2819) );
  AOI21_X1 U18483 ( .B1(n9883), .B2(n14932), .A(n14920), .ZN(n15449) );
  INV_X1 U18484 ( .A(n15449), .ZN(n15262) );
  INV_X1 U18485 ( .A(n14933), .ZN(n14934) );
  AOI21_X1 U18486 ( .B1(n14935), .B2(n14947), .A(n14934), .ZN(n15689) );
  INV_X1 U18487 ( .A(n14936), .ZN(n14948) );
  AND2_X1 U18488 ( .A1(n21251), .A2(n14948), .ZN(n14953) );
  AOI21_X1 U18489 ( .B1(n14953), .B2(P1_REIP_REG_19__SCAN_IN), .A(
        P1_REIP_REG_20__SCAN_IN), .ZN(n14939) );
  AOI22_X1 U18490 ( .A1(n21223), .A2(P1_EBX_REG_20__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n21233), .ZN(n14937) );
  OAI21_X1 U18491 ( .B1(n14939), .B2(n14938), .A(n14937), .ZN(n14941) );
  NOR2_X1 U18492 ( .A1(n21263), .A2(n15447), .ZN(n14940) );
  AOI211_X1 U18493 ( .C1(n15689), .C2(n21259), .A(n14941), .B(n14940), .ZN(
        n14942) );
  OAI21_X1 U18494 ( .B1(n15262), .B2(n17648), .A(n14942), .ZN(P1_U2820) );
  OAI21_X1 U18495 ( .B1(n14943), .B2(n9850), .A(n14932), .ZN(n15453) );
  NAND2_X1 U18496 ( .A1(n14944), .A2(n14945), .ZN(n14946) );
  AND2_X1 U18497 ( .A1(n14947), .A2(n14946), .ZN(n15698) );
  NAND2_X1 U18498 ( .A1(n21170), .A2(n14948), .ZN(n14949) );
  NAND2_X1 U18499 ( .A1(n21217), .A2(n14949), .ZN(n14968) );
  NAND2_X1 U18500 ( .A1(n21174), .A2(n15456), .ZN(n14955) );
  INV_X1 U18501 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n15130) );
  NAND2_X1 U18502 ( .A1(n21170), .A2(n14950), .ZN(n21235) );
  NAND2_X1 U18503 ( .A1(n21233), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14951) );
  OAI211_X1 U18504 ( .C1(n21256), .C2(n15130), .A(n21235), .B(n14951), .ZN(
        n14952) );
  AOI21_X1 U18505 ( .B1(n14953), .B2(n14956), .A(n14952), .ZN(n14954) );
  OAI211_X1 U18506 ( .C1(n14956), .C2(n14968), .A(n14955), .B(n14954), .ZN(
        n14957) );
  AOI21_X1 U18507 ( .B1(n21259), .B2(n15698), .A(n14957), .ZN(n14958) );
  OAI21_X1 U18508 ( .B1(n15453), .B2(n17648), .A(n14958), .ZN(P1_U2821) );
  OR2_X1 U18509 ( .A1(n14959), .A2(n14960), .ZN(n14961) );
  NAND2_X1 U18510 ( .A1(n14944), .A2(n14961), .ZN(n15702) );
  AOI21_X1 U18511 ( .B1(n14963), .B2(n14962), .A(n9850), .ZN(n15131) );
  NAND2_X1 U18512 ( .A1(n15131), .A2(n21212), .ZN(n14972) );
  INV_X1 U18513 ( .A(n15459), .ZN(n14970) );
  AOI21_X1 U18514 ( .B1(n21251), .B2(n14976), .A(P1_REIP_REG_18__SCAN_IN), 
        .ZN(n14967) );
  NAND2_X1 U18515 ( .A1(n21233), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14964) );
  OAI211_X1 U18516 ( .C1(n21256), .C2(n15132), .A(n21235), .B(n14964), .ZN(
        n14965) );
  INV_X1 U18517 ( .A(n14965), .ZN(n14966) );
  OAI21_X1 U18518 ( .B1(n14968), .B2(n14967), .A(n14966), .ZN(n14969) );
  AOI21_X1 U18519 ( .B1(n21174), .B2(n14970), .A(n14969), .ZN(n14971) );
  OAI211_X1 U18520 ( .C1(n15702), .C2(n17647), .A(n14972), .B(n14971), .ZN(
        P1_U2822) );
  NAND2_X1 U18521 ( .A1(n14973), .A2(n14974), .ZN(n14975) );
  NAND2_X1 U18522 ( .A1(n14962), .A2(n14975), .ZN(n15477) );
  OAI21_X1 U18523 ( .B1(n14977), .B2(n14976), .A(n21170), .ZN(n14987) );
  INV_X1 U18524 ( .A(n14978), .ZN(n14997) );
  NAND2_X1 U18525 ( .A1(n21251), .A2(n14997), .ZN(n15080) );
  INV_X1 U18526 ( .A(n14998), .ZN(n14979) );
  NOR2_X1 U18527 ( .A1(n15080), .A2(n14979), .ZN(n15020) );
  INV_X1 U18528 ( .A(n15020), .ZN(n14980) );
  OAI21_X1 U18529 ( .B1(n14980), .B2(n15000), .A(n15472), .ZN(n14986) );
  INV_X1 U18530 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n22213) );
  INV_X1 U18531 ( .A(n21235), .ZN(n21221) );
  AOI21_X1 U18532 ( .B1(n21233), .B2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n21221), .ZN(n14981) );
  OAI21_X1 U18533 ( .B1(n21256), .B2(n22213), .A(n14981), .ZN(n14985) );
  NOR2_X1 U18534 ( .A1(n14994), .A2(n14982), .ZN(n14983) );
  OR2_X1 U18535 ( .A1(n14959), .A2(n14983), .ZN(n15717) );
  OAI22_X1 U18536 ( .A1(n21263), .A2(n15473), .B1(n17647), .B2(n15717), .ZN(
        n14984) );
  AOI211_X1 U18537 ( .C1(n14987), .C2(n14986), .A(n14985), .B(n14984), .ZN(
        n14988) );
  OAI21_X1 U18538 ( .B1(n15477), .B2(n17648), .A(n14988), .ZN(P1_U2823) );
  INV_X1 U18539 ( .A(n14989), .ZN(n15008) );
  INV_X1 U18540 ( .A(n14990), .ZN(n14991) );
  NAND4_X1 U18541 ( .A1(n15008), .A2(n14991), .A3(n15013), .A4(n15028), .ZN(
        n15012) );
  INV_X1 U18542 ( .A(n15012), .ZN(n14993) );
  OAI21_X1 U18543 ( .B1(n14993), .B2(n14992), .A(n14973), .ZN(n15486) );
  AOI21_X1 U18544 ( .B1(n14995), .B2(n15017), .A(n14994), .ZN(n14996) );
  INV_X1 U18545 ( .A(n14996), .ZN(n15727) );
  AND2_X1 U18546 ( .A1(n21170), .A2(n14997), .ZN(n15078) );
  NAND2_X1 U18547 ( .A1(n15078), .A2(n14998), .ZN(n14999) );
  AND2_X1 U18548 ( .A1(n21217), .A2(n14999), .ZN(n15035) );
  OAI211_X1 U18549 ( .C1(P1_REIP_REG_15__SCAN_IN), .C2(P1_REIP_REG_16__SCAN_IN), .A(n15020), .B(n15000), .ZN(n15002) );
  AOI21_X1 U18550 ( .B1(n21233), .B2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n21221), .ZN(n15001) );
  OAI211_X1 U18551 ( .C1(n15133), .C2(n21256), .A(n15002), .B(n15001), .ZN(
        n15003) );
  AOI21_X1 U18552 ( .B1(P1_REIP_REG_16__SCAN_IN), .B2(n15035), .A(n15003), 
        .ZN(n15004) );
  OAI21_X1 U18553 ( .B1(n15727), .B2(n17647), .A(n15004), .ZN(n15005) );
  AOI21_X1 U18554 ( .B1(n15489), .B2(n21174), .A(n15005), .ZN(n15006) );
  OAI21_X1 U18555 ( .B1(n15486), .B2(n17648), .A(n15006), .ZN(P1_U2824) );
  AOI21_X1 U18556 ( .B1(n15077), .B2(n15008), .A(n15043), .ZN(n15010) );
  INV_X1 U18557 ( .A(n15028), .ZN(n15011) );
  NOR2_X1 U18558 ( .A1(n15045), .A2(n15011), .ZN(n15026) );
  OAI21_X1 U18559 ( .B1(n15026), .B2(n15013), .A(n15012), .ZN(n15500) );
  INV_X1 U18560 ( .A(n15492), .ZN(n15024) );
  NAND2_X1 U18561 ( .A1(n15014), .A2(n15015), .ZN(n15016) );
  NAND2_X1 U18562 ( .A1(n15017), .A2(n15016), .ZN(n15736) );
  INV_X1 U18563 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n15134) );
  NAND2_X1 U18564 ( .A1(n21233), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15018) );
  OAI211_X1 U18565 ( .C1(n21256), .C2(n15134), .A(n21235), .B(n15018), .ZN(
        n15019) );
  AOI21_X1 U18566 ( .B1(n15020), .B2(n15491), .A(n15019), .ZN(n15022) );
  NAND2_X1 U18567 ( .A1(n15035), .A2(P1_REIP_REG_15__SCAN_IN), .ZN(n15021) );
  OAI211_X1 U18568 ( .C1(n15736), .C2(n17647), .A(n15022), .B(n15021), .ZN(
        n15023) );
  AOI21_X1 U18569 ( .B1(n21174), .B2(n15024), .A(n15023), .ZN(n15025) );
  OAI21_X1 U18570 ( .B1(n15500), .B2(n17648), .A(n15025), .ZN(P1_U2825) );
  INV_X1 U18571 ( .A(n15045), .ZN(n15029) );
  INV_X1 U18572 ( .A(n15026), .ZN(n15027) );
  INV_X1 U18573 ( .A(n15502), .ZN(n15040) );
  OR2_X1 U18574 ( .A1(n15052), .A2(n15030), .ZN(n15031) );
  NAND2_X1 U18575 ( .A1(n15014), .A2(n15031), .ZN(n15747) );
  INV_X1 U18576 ( .A(n15747), .ZN(n15034) );
  NAND2_X1 U18577 ( .A1(n21233), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15032) );
  OAI211_X1 U18578 ( .C1(n21256), .C2(n15135), .A(n21235), .B(n15032), .ZN(
        n15033) );
  AOI21_X1 U18579 ( .B1(n15034), .B2(n21259), .A(n15033), .ZN(n15038) );
  OR2_X1 U18580 ( .A1(n15080), .A2(n15047), .ZN(n15056) );
  OAI21_X1 U18581 ( .B1(n15056), .B2(n21880), .A(n15501), .ZN(n15036) );
  NAND2_X1 U18582 ( .A1(n15036), .A2(n15035), .ZN(n15037) );
  NAND2_X1 U18583 ( .A1(n15038), .A2(n15037), .ZN(n15039) );
  AOI21_X1 U18584 ( .B1(n21174), .B2(n15040), .A(n15039), .ZN(n15041) );
  OAI21_X1 U18585 ( .B1(n15511), .B2(n17648), .A(n15041), .ZN(P1_U2826) );
  AOI21_X1 U18586 ( .B1(n15042), .B2(n14989), .A(n15043), .ZN(n15076) );
  AOI21_X1 U18587 ( .B1(n15076), .B2(n15077), .A(n15043), .ZN(n15062) );
  INV_X1 U18588 ( .A(n15044), .ZN(n15061) );
  NOR2_X1 U18589 ( .A1(n15062), .A2(n15061), .ZN(n15060) );
  OAI21_X1 U18590 ( .B1(n15060), .B2(n15046), .A(n15045), .ZN(n15522) );
  INV_X1 U18591 ( .A(n15047), .ZN(n15048) );
  INV_X1 U18592 ( .A(n21217), .ZN(n15079) );
  AOI21_X1 U18593 ( .B1(n15048), .B2(n15078), .A(n15079), .ZN(n15067) );
  OAI21_X1 U18594 ( .B1(n21253), .B2(n15049), .A(n21235), .ZN(n15054) );
  NOR2_X1 U18595 ( .A1(n9856), .A2(n15050), .ZN(n15051) );
  OR2_X1 U18596 ( .A1(n15052), .A2(n15051), .ZN(n15773) );
  NOR2_X1 U18597 ( .A1(n15773), .A2(n17647), .ZN(n15053) );
  AOI211_X1 U18598 ( .C1(P1_EBX_REG_13__SCAN_IN), .C2(n21223), .A(n15054), .B(
        n15053), .ZN(n15055) );
  OAI21_X1 U18599 ( .B1(P1_REIP_REG_13__SCAN_IN), .B2(n15056), .A(n15055), 
        .ZN(n15058) );
  NOR2_X1 U18600 ( .A1(n21263), .A2(n15512), .ZN(n15057) );
  AOI211_X1 U18601 ( .C1(P1_REIP_REG_13__SCAN_IN), .C2(n15067), .A(n15058), 
        .B(n15057), .ZN(n15059) );
  OAI21_X1 U18602 ( .B1(n15522), .B2(n17648), .A(n15059), .ZN(P1_U2827) );
  AOI21_X1 U18603 ( .B1(n15062), .B2(n15061), .A(n15060), .ZN(n15063) );
  INV_X1 U18604 ( .A(n15063), .ZN(n15531) );
  INV_X1 U18605 ( .A(n15524), .ZN(n15074) );
  AND2_X1 U18606 ( .A1(n15084), .A2(n15064), .ZN(n15065) );
  OR2_X1 U18607 ( .A1(n15065), .A2(n9856), .ZN(n15794) );
  NOR2_X1 U18608 ( .A1(n15080), .A2(n15066), .ZN(n15068) );
  OAI21_X1 U18609 ( .B1(P1_REIP_REG_12__SCAN_IN), .B2(n15068), .A(n15067), 
        .ZN(n15072) );
  OAI21_X1 U18610 ( .B1(n21253), .B2(n15069), .A(n21235), .ZN(n15070) );
  AOI21_X1 U18611 ( .B1(n21223), .B2(P1_EBX_REG_12__SCAN_IN), .A(n15070), .ZN(
        n15071) );
  OAI211_X1 U18612 ( .C1(n15794), .C2(n17647), .A(n15072), .B(n15071), .ZN(
        n15073) );
  AOI21_X1 U18613 ( .B1(n21174), .B2(n15074), .A(n15073), .ZN(n15075) );
  OAI21_X1 U18614 ( .B1(n15531), .B2(n17648), .A(n15075), .ZN(P1_U2828) );
  XOR2_X1 U18615 ( .A(n15077), .B(n15076), .Z(n15540) );
  NAND2_X1 U18616 ( .A1(n15540), .A2(n21212), .ZN(n15090) );
  NOR2_X1 U18617 ( .A1(n15079), .A2(n15078), .ZN(n17653) );
  NOR2_X1 U18618 ( .A1(n15080), .A2(P1_REIP_REG_11__SCAN_IN), .ZN(n15088) );
  NAND2_X1 U18619 ( .A1(n15081), .A2(n15082), .ZN(n15083) );
  NAND2_X1 U18620 ( .A1(n15084), .A2(n15083), .ZN(n15804) );
  INV_X1 U18621 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n15138) );
  NOR2_X1 U18622 ( .A1(n21256), .A2(n15138), .ZN(n15085) );
  AOI211_X1 U18623 ( .C1(n21233), .C2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n21221), .B(n15085), .ZN(n15086) );
  OAI21_X1 U18624 ( .B1(n17647), .B2(n15804), .A(n15086), .ZN(n15087) );
  AOI211_X1 U18625 ( .C1(n17653), .C2(P1_REIP_REG_11__SCAN_IN), .A(n15088), 
        .B(n15087), .ZN(n15089) );
  OAI211_X1 U18626 ( .C1(n21263), .C2(n15538), .A(n15090), .B(n15089), .ZN(
        P1_U2829) );
  NOR2_X1 U18627 ( .A1(n15095), .A2(n15091), .ZN(n15092) );
  NAND2_X1 U18628 ( .A1(n21265), .A2(n15093), .ZN(n15103) );
  NOR2_X1 U18629 ( .A1(n15095), .A2(n15094), .ZN(n21240) );
  INV_X1 U18630 ( .A(n21240), .ZN(n21252) );
  AOI22_X1 U18631 ( .A1(n21233), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n21249), .B2(P1_REIP_REG_2__SCAN_IN), .ZN(n15096) );
  OAI21_X1 U18632 ( .B1(n21252), .B2(n13896), .A(n15096), .ZN(n15101) );
  NAND2_X1 U18633 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_2__SCAN_IN), 
        .ZN(n15097) );
  OAI211_X1 U18634 ( .C1(P1_REIP_REG_2__SCAN_IN), .C2(P1_REIP_REG_1__SCAN_IN), 
        .A(n21251), .B(n15097), .ZN(n15098) );
  OAI21_X1 U18635 ( .B1(n17647), .B2(n15099), .A(n15098), .ZN(n15100) );
  AOI211_X1 U18636 ( .C1(n21223), .C2(P1_EBX_REG_2__SCAN_IN), .A(n15101), .B(
        n15100), .ZN(n15102) );
  OAI211_X1 U18637 ( .C1(n21263), .C2(n15104), .A(n15103), .B(n15102), .ZN(
        P1_U2838) );
  MUX2_X1 U18638 ( .A(n21263), .B(n21253), .S(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .Z(n15111) );
  NOR2_X1 U18639 ( .A1(n21170), .A2(n21896), .ZN(n15106) );
  AOI21_X1 U18640 ( .B1(n21240), .B2(n21778), .A(n15106), .ZN(n15110) );
  AOI22_X1 U18641 ( .A1(n21259), .A2(n15107), .B1(n21251), .B2(n21896), .ZN(
        n15109) );
  OR2_X1 U18642 ( .A1(n21256), .A2(n13388), .ZN(n15108) );
  OAI21_X1 U18643 ( .B1(n21225), .B2(n15113), .A(n15112), .ZN(P1_U2839) );
  AOI22_X1 U18644 ( .A1(n21223), .A2(P1_EBX_REG_0__SCAN_IN), .B1(n12709), .B2(
        n21240), .ZN(n15114) );
  OAI21_X1 U18645 ( .B1(n17647), .B2(n15115), .A(n15114), .ZN(n15116) );
  AOI21_X1 U18646 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(n21217), .A(n15116), .ZN(
        n15118) );
  OAI21_X1 U18647 ( .B1(n21174), .B2(n21233), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n15117) );
  OAI211_X1 U18648 ( .C1(n21225), .C2(n15119), .A(n15118), .B(n15117), .ZN(
        P1_U2840) );
  AOI22_X1 U18649 ( .A1(n15589), .A2(n15175), .B1(P1_EBX_REG_30__SCAN_IN), 
        .B2(n15174), .ZN(n15120) );
  OAI21_X1 U18650 ( .B1(n15202), .B2(n15195), .A(n15120), .ZN(P1_U2842) );
  OAI222_X1 U18651 ( .A1(n15187), .A2(n15372), .B1(n15121), .B2(n15194), .C1(
        n15598), .C2(n15192), .ZN(P1_U2843) );
  AOI22_X1 U18652 ( .A1(n15603), .A2(n15175), .B1(P1_EBX_REG_28__SCAN_IN), 
        .B2(n15174), .ZN(n15122) );
  OAI21_X1 U18653 ( .B1(n15214), .B2(n15195), .A(n15122), .ZN(P1_U2844) );
  INV_X1 U18654 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n15123) );
  OAI222_X1 U18655 ( .A1(n15187), .A2(n15389), .B1(n15123), .B2(n15194), .C1(
        n15615), .C2(n15192), .ZN(P1_U2845) );
  INV_X1 U18656 ( .A(n15397), .ZN(n15226) );
  OAI222_X1 U18657 ( .A1(n15187), .A2(n15226), .B1(n22185), .B2(n15194), .C1(
        n15619), .C2(n15192), .ZN(P1_U2846) );
  OAI222_X1 U18658 ( .A1(n15187), .A2(n15406), .B1(n22121), .B2(n15194), .C1(
        n15634), .C2(n15192), .ZN(P1_U2847) );
  AOI22_X1 U18659 ( .A1(n15642), .A2(n15175), .B1(P1_EBX_REG_24__SCAN_IN), 
        .B2(n15174), .ZN(n15124) );
  OAI21_X1 U18660 ( .B1(n15237), .B2(n15195), .A(n15124), .ZN(P1_U2848) );
  INV_X1 U18661 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n15125) );
  OAI222_X1 U18662 ( .A1(n15417), .A2(n15195), .B1(n15125), .B2(n15194), .C1(
        n15646), .C2(n15192), .ZN(P1_U2849) );
  INV_X1 U18663 ( .A(n15430), .ZN(n15250) );
  OAI222_X1 U18664 ( .A1(n15250), .A2(n15195), .B1(n15126), .B2(n15194), .C1(
        n15662), .C2(n15192), .ZN(P1_U2850) );
  AOI22_X1 U18665 ( .A1(n15666), .A2(n15175), .B1(P1_EBX_REG_21__SCAN_IN), 
        .B2(n15174), .ZN(n15127) );
  OAI21_X1 U18666 ( .B1(n15440), .B2(n15195), .A(n15127), .ZN(P1_U2851) );
  AOI22_X1 U18667 ( .A1(n15689), .A2(n15175), .B1(P1_EBX_REG_20__SCAN_IN), 
        .B2(n15174), .ZN(n15128) );
  OAI21_X1 U18668 ( .B1(n15262), .B2(n15195), .A(n15128), .ZN(P1_U2852) );
  INV_X1 U18669 ( .A(n15698), .ZN(n15129) );
  OAI222_X1 U18670 ( .A1(n15453), .A2(n15195), .B1(n15130), .B2(n15194), .C1(
        n15129), .C2(n15192), .ZN(P1_U2853) );
  INV_X1 U18671 ( .A(n15131), .ZN(n15465) );
  OAI222_X1 U18672 ( .A1(n15465), .A2(n15195), .B1(n15132), .B2(n15194), .C1(
        n15702), .C2(n15192), .ZN(P1_U2854) );
  OAI222_X1 U18673 ( .A1(n15477), .A2(n15187), .B1(n22213), .B2(n15194), .C1(
        n15717), .C2(n15192), .ZN(P1_U2855) );
  OAI222_X1 U18674 ( .A1(n15486), .A2(n15187), .B1(n15133), .B2(n15194), .C1(
        n15727), .C2(n15192), .ZN(P1_U2856) );
  OAI222_X1 U18675 ( .A1(n15500), .A2(n15187), .B1(n15134), .B2(n15194), .C1(
        n15736), .C2(n15192), .ZN(P1_U2857) );
  OAI222_X1 U18676 ( .A1(n15511), .A2(n15187), .B1(n15135), .B2(n15194), .C1(
        n15747), .C2(n15192), .ZN(P1_U2858) );
  INV_X1 U18677 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n15136) );
  OAI222_X1 U18678 ( .A1(n15522), .A2(n15187), .B1(n15136), .B2(n15194), .C1(
        n15773), .C2(n15192), .ZN(P1_U2859) );
  INV_X1 U18679 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n15137) );
  OAI222_X1 U18680 ( .A1(n15794), .A2(n15192), .B1(n15137), .B2(n15194), .C1(
        n15531), .C2(n15187), .ZN(P1_U2860) );
  INV_X1 U18681 ( .A(n15540), .ZN(n15288) );
  OAI222_X1 U18682 ( .A1(n15288), .A2(n15187), .B1(n15138), .B2(n15194), .C1(
        n15804), .C2(n15192), .ZN(P1_U2861) );
  OR2_X1 U18683 ( .A1(n15139), .A2(n15140), .ZN(n15141) );
  NAND2_X1 U18684 ( .A1(n14989), .A2(n15141), .ZN(n17649) );
  INV_X1 U18685 ( .A(n17649), .ZN(n15146) );
  OR2_X1 U18686 ( .A1(n9873), .A2(n15142), .ZN(n15143) );
  NAND2_X1 U18687 ( .A1(n15081), .A2(n15143), .ZN(n17646) );
  OAI22_X1 U18688 ( .A1(n15192), .A2(n17646), .B1(n17645), .B2(n15194), .ZN(
        n15144) );
  AOI21_X1 U18689 ( .B1(n15146), .B2(n15145), .A(n15144), .ZN(n15147) );
  INV_X1 U18690 ( .A(n15147), .ZN(P1_U2862) );
  AND2_X1 U18691 ( .A1(n15148), .A2(n15149), .ZN(n15150) );
  OR2_X1 U18692 ( .A1(n15139), .A2(n15150), .ZN(n21173) );
  AOI21_X1 U18693 ( .B1(n9881), .B2(n15154), .A(n15151), .ZN(n15152) );
  OR2_X1 U18694 ( .A1(n15152), .A2(n9873), .ZN(n15827) );
  INV_X1 U18695 ( .A(n15827), .ZN(n21172) );
  AOI22_X1 U18696 ( .A1(n21172), .A2(n15175), .B1(P1_EBX_REG_9__SCAN_IN), .B2(
        n15174), .ZN(n15153) );
  OAI21_X1 U18697 ( .B1(n21173), .B2(n15187), .A(n15153), .ZN(P1_U2863) );
  OAI21_X1 U18698 ( .B1(n12755), .B2(n9884), .A(n15148), .ZN(n21184) );
  INV_X1 U18699 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n15155) );
  XNOR2_X1 U18700 ( .A(n9881), .B(n15154), .ZN(n17679) );
  OAI222_X1 U18701 ( .A1(n15187), .A2(n21184), .B1(n15155), .B2(n15194), .C1(
        n15192), .C2(n17679), .ZN(P1_U2864) );
  OR2_X1 U18702 ( .A1(n15156), .A2(n15157), .ZN(n15158) );
  INV_X1 U18703 ( .A(n21200), .ZN(n15295) );
  INV_X1 U18704 ( .A(n15172), .ZN(n15166) );
  AOI21_X1 U18705 ( .B1(n15166), .B2(n15165), .A(n15159), .ZN(n15160) );
  NOR2_X1 U18706 ( .A1(n15160), .A2(n9881), .ZN(n21199) );
  AOI22_X1 U18707 ( .A1(n15175), .A2(n21199), .B1(n15174), .B2(
        P1_EBX_REG_7__SCAN_IN), .ZN(n15161) );
  OAI21_X1 U18708 ( .B1(n15295), .B2(n15195), .A(n15161), .ZN(P1_U2865) );
  AND2_X1 U18709 ( .A1(n15162), .A2(n15163), .ZN(n15164) );
  OR2_X1 U18710 ( .A1(n15156), .A2(n15164), .ZN(n17667) );
  INV_X1 U18711 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n15167) );
  XNOR2_X1 U18712 ( .A(n15166), .B(n15165), .ZN(n17696) );
  OAI222_X1 U18713 ( .A1(n15187), .A2(n17667), .B1(n15167), .B2(n15194), .C1(
        n15192), .C2(n17696), .ZN(P1_U2866) );
  OR2_X1 U18714 ( .A1(n15177), .A2(n15168), .ZN(n15169) );
  NAND2_X1 U18715 ( .A1(n15162), .A2(n15169), .ZN(n21226) );
  OAI21_X1 U18716 ( .B1(n15170), .B2(n15184), .A(n15171), .ZN(n15173) );
  NAND2_X1 U18717 ( .A1(n15173), .A2(n15172), .ZN(n15838) );
  INV_X1 U18718 ( .A(n15838), .ZN(n21222) );
  AOI22_X1 U18719 ( .A1(n15175), .A2(n21222), .B1(n15174), .B2(
        P1_EBX_REG_5__SCAN_IN), .ZN(n15176) );
  OAI21_X1 U18720 ( .B1(n21226), .B2(n15195), .A(n15176), .ZN(P1_U2867) );
  NAND2_X1 U18721 ( .A1(n15179), .A2(n15178), .ZN(n15189) );
  NAND2_X1 U18722 ( .A1(n15189), .A2(n15180), .ZN(n15188) );
  INV_X1 U18723 ( .A(n15181), .ZN(n15182) );
  NAND2_X1 U18724 ( .A1(n15188), .A2(n15182), .ZN(n15183) );
  NAND2_X1 U18725 ( .A1(n10273), .A2(n15183), .ZN(n21230) );
  INV_X1 U18726 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n21236) );
  INV_X1 U18727 ( .A(n15184), .ZN(n15185) );
  XNOR2_X1 U18728 ( .A(n15170), .B(n15185), .ZN(n21232) );
  INV_X1 U18729 ( .A(n21232), .ZN(n15186) );
  OAI222_X1 U18730 ( .A1(n15187), .A2(n21230), .B1(n15194), .B2(n21236), .C1(
        n15192), .C2(n15186), .ZN(P1_U2868) );
  OAI21_X1 U18731 ( .B1(n15189), .B2(n15180), .A(n15188), .ZN(n15581) );
  INV_X1 U18732 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n21255) );
  OR2_X1 U18733 ( .A1(n14073), .A2(n15190), .ZN(n15191) );
  AND2_X1 U18734 ( .A1(n15170), .A2(n15191), .ZN(n21260) );
  INV_X1 U18735 ( .A(n21260), .ZN(n15193) );
  OAI222_X1 U18736 ( .A1(n15581), .A2(n15195), .B1(n15194), .B2(n21255), .C1(
        n15193), .C2(n15192), .ZN(P1_U2869) );
  INV_X1 U18737 ( .A(DATAI_14_), .ZN(n15197) );
  NAND2_X1 U18738 ( .A1(n21327), .A2(BUF1_REG_14__SCAN_IN), .ZN(n15196) );
  OAI21_X1 U18739 ( .B1(n21327), .B2(n15197), .A(n15196), .ZN(n21310) );
  AOI22_X1 U18740 ( .A1(n15272), .A2(n21310), .B1(n15291), .B2(
        P1_EAX_REG_30__SCAN_IN), .ZN(n15198) );
  OAI21_X1 U18741 ( .B1(n15199), .B2(n15274), .A(n15198), .ZN(n15200) );
  AOI21_X1 U18742 ( .B1(n15281), .B2(DATAI_30_), .A(n15200), .ZN(n15201) );
  OAI21_X1 U18743 ( .B1(n15202), .B2(n15299), .A(n15201), .ZN(P1_U2874) );
  INV_X1 U18744 ( .A(DATAI_13_), .ZN(n15204) );
  MUX2_X1 U18745 ( .A(n15204), .B(n15203), .S(n21327), .Z(n15325) );
  OAI22_X1 U18746 ( .A1(n15278), .A2(n15325), .B1(n15296), .B2(n15205), .ZN(
        n15206) );
  AOI21_X1 U18747 ( .B1(n15280), .B2(BUF1_REG_29__SCAN_IN), .A(n15206), .ZN(
        n15208) );
  NAND2_X1 U18748 ( .A1(n15281), .A2(DATAI_29_), .ZN(n15207) );
  OAI211_X1 U18749 ( .C1(n15372), .C2(n15299), .A(n15208), .B(n15207), .ZN(
        P1_U2875) );
  INV_X1 U18750 ( .A(DATAI_12_), .ZN(n15210) );
  NAND2_X1 U18751 ( .A1(n21327), .A2(BUF1_REG_12__SCAN_IN), .ZN(n15209) );
  OAI21_X1 U18752 ( .B1(n21327), .B2(n15210), .A(n15209), .ZN(n21308) );
  AOI22_X1 U18753 ( .A1(n15272), .A2(n21308), .B1(n15291), .B2(
        P1_EAX_REG_28__SCAN_IN), .ZN(n15211) );
  OAI21_X1 U18754 ( .B1(n15274), .B2(n17841), .A(n15211), .ZN(n15212) );
  AOI21_X1 U18755 ( .B1(n15281), .B2(DATAI_28_), .A(n15212), .ZN(n15213) );
  OAI21_X1 U18756 ( .B1(n15214), .B2(n15299), .A(n15213), .ZN(P1_U2876) );
  INV_X1 U18757 ( .A(DATAI_11_), .ZN(n15216) );
  MUX2_X1 U18758 ( .A(n15216), .B(n15215), .S(n21327), .Z(n21305) );
  OAI22_X1 U18759 ( .A1(n15278), .A2(n21305), .B1(n15296), .B2(n15217), .ZN(
        n15218) );
  AOI21_X1 U18760 ( .B1(n15280), .B2(BUF1_REG_27__SCAN_IN), .A(n15218), .ZN(
        n15220) );
  NAND2_X1 U18761 ( .A1(n15281), .A2(DATAI_27_), .ZN(n15219) );
  OAI211_X1 U18762 ( .C1(n15389), .C2(n15299), .A(n15220), .B(n15219), .ZN(
        P1_U2877) );
  INV_X1 U18763 ( .A(DATAI_10_), .ZN(n15221) );
  MUX2_X1 U18764 ( .A(n15221), .B(n17865), .S(n21327), .Z(n15322) );
  OAI22_X1 U18765 ( .A1(n15278), .A2(n15322), .B1(n15296), .B2(n15222), .ZN(
        n15223) );
  AOI21_X1 U18766 ( .B1(n15280), .B2(BUF1_REG_26__SCAN_IN), .A(n15223), .ZN(
        n15225) );
  NAND2_X1 U18767 ( .A1(n15281), .A2(DATAI_26_), .ZN(n15224) );
  OAI211_X1 U18768 ( .C1(n15226), .C2(n15299), .A(n15225), .B(n15224), .ZN(
        P1_U2878) );
  INV_X1 U18769 ( .A(DATAI_9_), .ZN(n15227) );
  MUX2_X1 U18770 ( .A(n15227), .B(n17866), .S(n21327), .Z(n21302) );
  INV_X1 U18771 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n15228) );
  OAI22_X1 U18772 ( .A1(n15278), .A2(n21302), .B1(n15296), .B2(n15228), .ZN(
        n15229) );
  AOI21_X1 U18773 ( .B1(n15280), .B2(BUF1_REG_25__SCAN_IN), .A(n15229), .ZN(
        n15231) );
  NAND2_X1 U18774 ( .A1(n15281), .A2(DATAI_25_), .ZN(n15230) );
  OAI211_X1 U18775 ( .C1(n15406), .C2(n15299), .A(n15231), .B(n15230), .ZN(
        P1_U2879) );
  INV_X1 U18776 ( .A(DATAI_8_), .ZN(n15233) );
  NAND2_X1 U18777 ( .A1(n21327), .A2(BUF1_REG_8__SCAN_IN), .ZN(n15232) );
  OAI21_X1 U18778 ( .B1(n21327), .B2(n15233), .A(n15232), .ZN(n15320) );
  AOI22_X1 U18779 ( .A1(n15272), .A2(n15320), .B1(n15291), .B2(
        P1_EAX_REG_24__SCAN_IN), .ZN(n15234) );
  OAI21_X1 U18780 ( .B1(n15274), .B2(n17846), .A(n15234), .ZN(n15235) );
  AOI21_X1 U18781 ( .B1(n15281), .B2(DATAI_24_), .A(n15235), .ZN(n15236) );
  OAI21_X1 U18782 ( .B1(n15237), .B2(n15299), .A(n15236), .ZN(P1_U2880) );
  NAND2_X1 U18783 ( .A1(n21329), .A2(DATAI_7_), .ZN(n15239) );
  NAND2_X1 U18784 ( .A1(n21327), .A2(BUF1_REG_7__SCAN_IN), .ZN(n15238) );
  AND2_X1 U18785 ( .A1(n15239), .A2(n15238), .ZN(n21376) );
  OAI22_X1 U18786 ( .A1(n15278), .A2(n21376), .B1(n15296), .B2(n15240), .ZN(
        n15241) );
  AOI21_X1 U18787 ( .B1(n15280), .B2(BUF1_REG_23__SCAN_IN), .A(n15241), .ZN(
        n15243) );
  NAND2_X1 U18788 ( .A1(n15281), .A2(DATAI_23_), .ZN(n15242) );
  OAI211_X1 U18789 ( .C1(n15417), .C2(n15299), .A(n15243), .B(n15242), .ZN(
        P1_U2881) );
  NAND2_X1 U18790 ( .A1(n21329), .A2(DATAI_6_), .ZN(n15245) );
  NAND2_X1 U18791 ( .A1(n21327), .A2(BUF1_REG_6__SCAN_IN), .ZN(n15244) );
  AND2_X1 U18792 ( .A1(n15245), .A2(n15244), .ZN(n21366) );
  OAI22_X1 U18793 ( .A1(n15278), .A2(n21366), .B1(n15296), .B2(n15246), .ZN(
        n15247) );
  AOI21_X1 U18794 ( .B1(n15280), .B2(BUF1_REG_22__SCAN_IN), .A(n15247), .ZN(
        n15249) );
  NAND2_X1 U18795 ( .A1(n15281), .A2(DATAI_22_), .ZN(n15248) );
  OAI211_X1 U18796 ( .C1(n15250), .C2(n15299), .A(n15249), .B(n15248), .ZN(
        P1_U2882) );
  NAND2_X1 U18797 ( .A1(n21329), .A2(DATAI_5_), .ZN(n15252) );
  NAND2_X1 U18798 ( .A1(n21327), .A2(BUF1_REG_5__SCAN_IN), .ZN(n15251) );
  AND2_X1 U18799 ( .A1(n15252), .A2(n15251), .ZN(n21362) );
  OAI22_X1 U18800 ( .A1(n15278), .A2(n21362), .B1(n15296), .B2(n15253), .ZN(
        n15254) );
  AOI21_X1 U18801 ( .B1(n15280), .B2(BUF1_REG_21__SCAN_IN), .A(n15254), .ZN(
        n15256) );
  NAND2_X1 U18802 ( .A1(n15281), .A2(DATAI_21_), .ZN(n15255) );
  OAI211_X1 U18803 ( .C1(n15440), .C2(n15299), .A(n15256), .B(n15255), .ZN(
        P1_U2883) );
  INV_X1 U18804 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n17851) );
  INV_X1 U18805 ( .A(DATAI_4_), .ZN(n15258) );
  NAND2_X1 U18806 ( .A1(n21327), .A2(BUF1_REG_4__SCAN_IN), .ZN(n15257) );
  OAI21_X1 U18807 ( .B1(n21327), .B2(n15258), .A(n15257), .ZN(n15312) );
  AOI22_X1 U18808 ( .A1(n15272), .A2(n15312), .B1(n15291), .B2(
        P1_EAX_REG_20__SCAN_IN), .ZN(n15259) );
  OAI21_X1 U18809 ( .B1(n15274), .B2(n17851), .A(n15259), .ZN(n15260) );
  AOI21_X1 U18810 ( .B1(n15281), .B2(DATAI_20_), .A(n15260), .ZN(n15261) );
  OAI21_X1 U18811 ( .B1(n15262), .B2(n15299), .A(n15261), .ZN(P1_U2884) );
  INV_X1 U18812 ( .A(DATAI_3_), .ZN(n15264) );
  MUX2_X1 U18813 ( .A(n15264), .B(n15263), .S(n21327), .Z(n21355) );
  OAI22_X1 U18814 ( .A1(n15278), .A2(n21355), .B1(n15296), .B2(n15265), .ZN(
        n15266) );
  AOI21_X1 U18815 ( .B1(n15280), .B2(BUF1_REG_19__SCAN_IN), .A(n15266), .ZN(
        n15268) );
  NAND2_X1 U18816 ( .A1(n15281), .A2(DATAI_19_), .ZN(n15267) );
  OAI211_X1 U18817 ( .C1(n15453), .C2(n15299), .A(n15268), .B(n15267), .ZN(
        P1_U2885) );
  AOI22_X1 U18818 ( .A1(n15272), .A2(n15308), .B1(n15291), .B2(
        P1_EAX_REG_18__SCAN_IN), .ZN(n15269) );
  OAI21_X1 U18819 ( .B1(n15274), .B2(n17854), .A(n15269), .ZN(n15270) );
  AOI21_X1 U18820 ( .B1(n15281), .B2(DATAI_18_), .A(n15270), .ZN(n15271) );
  OAI21_X1 U18821 ( .B1(n15465), .B2(n15299), .A(n15271), .ZN(P1_U2886) );
  INV_X1 U18822 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n16479) );
  AOI22_X1 U18823 ( .A1(n15272), .A2(n15306), .B1(n15291), .B2(
        P1_EAX_REG_17__SCAN_IN), .ZN(n15273) );
  OAI21_X1 U18824 ( .B1(n15274), .B2(n16479), .A(n15273), .ZN(n15275) );
  AOI21_X1 U18825 ( .B1(n15281), .B2(DATAI_17_), .A(n15275), .ZN(n15276) );
  OAI21_X1 U18826 ( .B1(n15477), .B2(n15299), .A(n15276), .ZN(P1_U2887) );
  OAI22_X1 U18827 ( .A1(n15278), .A2(n21341), .B1(n15296), .B2(n15277), .ZN(
        n15279) );
  AOI21_X1 U18828 ( .B1(n15280), .B2(BUF1_REG_16__SCAN_IN), .A(n15279), .ZN(
        n15283) );
  NAND2_X1 U18829 ( .A1(n15281), .A2(DATAI_16_), .ZN(n15282) );
  OAI211_X1 U18830 ( .C1(n15486), .C2(n15299), .A(n15283), .B(n15282), .ZN(
        P1_U2888) );
  MUX2_X1 U18831 ( .A(DATAI_15_), .B(BUF1_REG_15__SCAN_IN), .S(n21327), .Z(
        n15349) );
  AOI22_X1 U18832 ( .A1(n15292), .A2(n15349), .B1(P1_EAX_REG_15__SCAN_IN), 
        .B2(n15291), .ZN(n15284) );
  OAI21_X1 U18833 ( .B1(n15500), .B2(n15299), .A(n15284), .ZN(P1_U2889) );
  AOI22_X1 U18834 ( .A1(n15292), .A2(n21310), .B1(P1_EAX_REG_14__SCAN_IN), 
        .B2(n15291), .ZN(n15285) );
  OAI21_X1 U18835 ( .B1(n15511), .B2(n15299), .A(n15285), .ZN(P1_U2890) );
  OAI222_X1 U18836 ( .A1(n15522), .A2(n15299), .B1(n15325), .B2(n15298), .C1(
        n22101), .C2(n15296), .ZN(P1_U2891) );
  AOI22_X1 U18837 ( .A1(n15292), .A2(n21308), .B1(P1_EAX_REG_12__SCAN_IN), 
        .B2(n15291), .ZN(n15286) );
  OAI21_X1 U18838 ( .B1(n15531), .B2(n15299), .A(n15286), .ZN(P1_U2892) );
  INV_X1 U18839 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n15287) );
  OAI222_X1 U18840 ( .A1(n15288), .A2(n15299), .B1(n21305), .B2(n15298), .C1(
        n15287), .C2(n15296), .ZN(P1_U2893) );
  INV_X1 U18841 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n15289) );
  OAI222_X1 U18842 ( .A1(n17649), .A2(n15299), .B1(n15322), .B2(n15298), .C1(
        n15289), .C2(n15296), .ZN(P1_U2894) );
  INV_X1 U18843 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n15290) );
  OAI222_X1 U18844 ( .A1(n21173), .A2(n15299), .B1(n21302), .B2(n15298), .C1(
        n15290), .C2(n15296), .ZN(P1_U2895) );
  AOI22_X1 U18845 ( .A1(n15292), .A2(n15320), .B1(P1_EAX_REG_8__SCAN_IN), .B2(
        n15291), .ZN(n15293) );
  OAI21_X1 U18846 ( .B1(n21184), .B2(n15299), .A(n15293), .ZN(P1_U2896) );
  INV_X1 U18847 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n15294) );
  OAI222_X1 U18848 ( .A1(n15295), .A2(n15299), .B1(n21376), .B2(n15298), .C1(
        n15294), .C2(n15296), .ZN(P1_U2897) );
  OAI222_X1 U18849 ( .A1(n15299), .A2(n17667), .B1(n21366), .B2(n15298), .C1(
        n15296), .C2(n12726), .ZN(P1_U2898) );
  INV_X1 U18850 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n22197) );
  OAI222_X1 U18851 ( .A1(n15299), .A2(n21226), .B1(n21362), .B2(n15298), .C1(
        n15296), .C2(n22197), .ZN(P1_U2899) );
  INV_X1 U18852 ( .A(n15312), .ZN(n21358) );
  INV_X1 U18853 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n21292) );
  OAI222_X1 U18854 ( .A1(n21230), .A2(n15299), .B1(n15298), .B2(n21358), .C1(
        n21292), .C2(n15296), .ZN(P1_U2900) );
  INV_X1 U18855 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n15297) );
  OAI222_X1 U18856 ( .A1(n15581), .A2(n15299), .B1(n15298), .B2(n21355), .C1(
        n15297), .C2(n15296), .ZN(P1_U2901) );
  AOI22_X1 U18857 ( .A1(n21322), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_UWORD_REG_0__SCAN_IN), .B2(n15346), .ZN(n15305) );
  INV_X1 U18858 ( .A(n21341), .ZN(n15304) );
  NAND2_X1 U18859 ( .A1(n21311), .A2(n15304), .ZN(n15328) );
  NAND2_X1 U18860 ( .A1(n15305), .A2(n15328), .ZN(P1_U2937) );
  AOI22_X1 U18861 ( .A1(n21322), .A2(P1_EAX_REG_17__SCAN_IN), .B1(
        P1_UWORD_REG_1__SCAN_IN), .B2(n15346), .ZN(n15307) );
  NAND2_X1 U18862 ( .A1(n21311), .A2(n15306), .ZN(n15330) );
  NAND2_X1 U18863 ( .A1(n15307), .A2(n15330), .ZN(P1_U2938) );
  AOI22_X1 U18864 ( .A1(n21322), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_UWORD_REG_2__SCAN_IN), .B2(n15346), .ZN(n15309) );
  NAND2_X1 U18865 ( .A1(n21311), .A2(n15308), .ZN(n15332) );
  NAND2_X1 U18866 ( .A1(n15309), .A2(n15332), .ZN(P1_U2939) );
  AOI22_X1 U18867 ( .A1(n21322), .A2(P1_EAX_REG_19__SCAN_IN), .B1(
        P1_UWORD_REG_3__SCAN_IN), .B2(n15346), .ZN(n15311) );
  INV_X1 U18868 ( .A(n21355), .ZN(n15310) );
  NAND2_X1 U18869 ( .A1(n21311), .A2(n15310), .ZN(n15334) );
  NAND2_X1 U18870 ( .A1(n15311), .A2(n15334), .ZN(P1_U2940) );
  AOI22_X1 U18871 ( .A1(n21322), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_UWORD_REG_4__SCAN_IN), .B2(n15346), .ZN(n15313) );
  NAND2_X1 U18872 ( .A1(n21311), .A2(n15312), .ZN(n15336) );
  NAND2_X1 U18873 ( .A1(n15313), .A2(n15336), .ZN(P1_U2941) );
  AOI22_X1 U18874 ( .A1(n21322), .A2(P1_EAX_REG_21__SCAN_IN), .B1(
        P1_UWORD_REG_5__SCAN_IN), .B2(n15346), .ZN(n15315) );
  INV_X1 U18875 ( .A(n21362), .ZN(n15314) );
  NAND2_X1 U18876 ( .A1(n21311), .A2(n15314), .ZN(n15338) );
  NAND2_X1 U18877 ( .A1(n15315), .A2(n15338), .ZN(P1_U2942) );
  AOI22_X1 U18878 ( .A1(n21322), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_UWORD_REG_6__SCAN_IN), .B2(n15346), .ZN(n15317) );
  INV_X1 U18879 ( .A(n21366), .ZN(n15316) );
  NAND2_X1 U18880 ( .A1(n21311), .A2(n15316), .ZN(n15340) );
  NAND2_X1 U18881 ( .A1(n15317), .A2(n15340), .ZN(P1_U2943) );
  AOI22_X1 U18882 ( .A1(n21322), .A2(P1_EAX_REG_23__SCAN_IN), .B1(
        P1_UWORD_REG_7__SCAN_IN), .B2(n15346), .ZN(n15319) );
  INV_X1 U18883 ( .A(n21376), .ZN(n15318) );
  NAND2_X1 U18884 ( .A1(n21311), .A2(n15318), .ZN(n15342) );
  NAND2_X1 U18885 ( .A1(n15319), .A2(n15342), .ZN(P1_U2944) );
  INV_X1 U18886 ( .A(P1_UWORD_REG_8__SCAN_IN), .ZN(n21994) );
  NAND2_X1 U18887 ( .A1(n21311), .A2(n15320), .ZN(n15344) );
  NAND2_X1 U18888 ( .A1(n21322), .A2(P1_EAX_REG_24__SCAN_IN), .ZN(n15321) );
  OAI211_X1 U18889 ( .C1(n15352), .C2(n21994), .A(n15344), .B(n15321), .ZN(
        P1_U2945) );
  AOI22_X1 U18890 ( .A1(n21322), .A2(P1_EAX_REG_26__SCAN_IN), .B1(
        P1_UWORD_REG_10__SCAN_IN), .B2(n15346), .ZN(n15324) );
  INV_X1 U18891 ( .A(n15322), .ZN(n15323) );
  NAND2_X1 U18892 ( .A1(n21311), .A2(n15323), .ZN(n21315) );
  NAND2_X1 U18893 ( .A1(n15324), .A2(n21315), .ZN(P1_U2947) );
  AOI22_X1 U18894 ( .A1(n21322), .A2(P1_EAX_REG_29__SCAN_IN), .B1(
        P1_UWORD_REG_13__SCAN_IN), .B2(n15346), .ZN(n15327) );
  INV_X1 U18895 ( .A(n15325), .ZN(n15326) );
  NAND2_X1 U18896 ( .A1(n21311), .A2(n15326), .ZN(n15347) );
  NAND2_X1 U18897 ( .A1(n15327), .A2(n15347), .ZN(P1_U2950) );
  AOI22_X1 U18898 ( .A1(n21322), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_LWORD_REG_0__SCAN_IN), .B2(n15346), .ZN(n15329) );
  NAND2_X1 U18899 ( .A1(n15329), .A2(n15328), .ZN(P1_U2952) );
  AOI22_X1 U18900 ( .A1(n21322), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_LWORD_REG_1__SCAN_IN), .B2(n15346), .ZN(n15331) );
  NAND2_X1 U18901 ( .A1(n15331), .A2(n15330), .ZN(P1_U2953) );
  AOI22_X1 U18902 ( .A1(n21322), .A2(P1_EAX_REG_2__SCAN_IN), .B1(
        P1_LWORD_REG_2__SCAN_IN), .B2(n15346), .ZN(n15333) );
  NAND2_X1 U18903 ( .A1(n15333), .A2(n15332), .ZN(P1_U2954) );
  AOI22_X1 U18904 ( .A1(n21322), .A2(P1_EAX_REG_3__SCAN_IN), .B1(
        P1_LWORD_REG_3__SCAN_IN), .B2(n15346), .ZN(n15335) );
  NAND2_X1 U18905 ( .A1(n15335), .A2(n15334), .ZN(P1_U2955) );
  AOI22_X1 U18906 ( .A1(n21322), .A2(P1_EAX_REG_4__SCAN_IN), .B1(
        P1_LWORD_REG_4__SCAN_IN), .B2(n21321), .ZN(n15337) );
  NAND2_X1 U18907 ( .A1(n15337), .A2(n15336), .ZN(P1_U2956) );
  AOI22_X1 U18908 ( .A1(n21322), .A2(P1_EAX_REG_5__SCAN_IN), .B1(
        P1_LWORD_REG_5__SCAN_IN), .B2(n15346), .ZN(n15339) );
  NAND2_X1 U18909 ( .A1(n15339), .A2(n15338), .ZN(P1_U2957) );
  AOI22_X1 U18910 ( .A1(n21322), .A2(P1_EAX_REG_6__SCAN_IN), .B1(
        P1_LWORD_REG_6__SCAN_IN), .B2(n21321), .ZN(n15341) );
  NAND2_X1 U18911 ( .A1(n15341), .A2(n15340), .ZN(P1_U2958) );
  AOI22_X1 U18912 ( .A1(n21322), .A2(P1_EAX_REG_7__SCAN_IN), .B1(
        P1_LWORD_REG_7__SCAN_IN), .B2(n15346), .ZN(n15343) );
  NAND2_X1 U18913 ( .A1(n15343), .A2(n15342), .ZN(P1_U2959) );
  INV_X1 U18914 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n21287) );
  NAND2_X1 U18915 ( .A1(n21321), .A2(P1_LWORD_REG_8__SCAN_IN), .ZN(n15345) );
  OAI211_X1 U18916 ( .C1(n15354), .C2(n21287), .A(n15345), .B(n15344), .ZN(
        P1_U2960) );
  AOI22_X1 U18917 ( .A1(n21322), .A2(P1_EAX_REG_13__SCAN_IN), .B1(
        P1_LWORD_REG_13__SCAN_IN), .B2(n15346), .ZN(n15348) );
  NAND2_X1 U18918 ( .A1(n15348), .A2(n15347), .ZN(P1_U2965) );
  INV_X1 U18919 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n15353) );
  INV_X1 U18920 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n21274) );
  INV_X1 U18921 ( .A(n21311), .ZN(n15351) );
  INV_X1 U18922 ( .A(n15349), .ZN(n15350) );
  OAI222_X1 U18923 ( .A1(n15354), .A2(n15353), .B1(n15352), .B2(n21274), .C1(
        n15351), .C2(n15350), .ZN(P1_U2967) );
  NAND2_X1 U18924 ( .A1(n15355), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15356) );
  XNOR2_X1 U18925 ( .A(n15358), .B(n15357), .ZN(n15590) );
  NOR2_X1 U18926 ( .A1(n15837), .A2(n15359), .ZN(n15588) );
  AOI21_X1 U18927 ( .B1(n17661), .B2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n15588), .ZN(n15360) );
  OAI21_X1 U18928 ( .B1(n15361), .B2(n17670), .A(n15360), .ZN(n15362) );
  OAI21_X1 U18929 ( .B1(n21153), .B2(n15590), .A(n15363), .ZN(P1_U2969) );
  NOR2_X1 U18930 ( .A1(n15837), .A2(n22188), .ZN(n15594) );
  INV_X1 U18931 ( .A(n15364), .ZN(n15365) );
  NOR2_X1 U18932 ( .A1(n15365), .A2(n17670), .ZN(n15366) );
  AOI211_X1 U18933 ( .C1(n17661), .C2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n15594), .B(n15366), .ZN(n15371) );
  XNOR2_X1 U18934 ( .A(n15554), .B(n15367), .ZN(n15368) );
  XNOR2_X1 U18935 ( .A(n15369), .B(n15368), .ZN(n15591) );
  NAND2_X1 U18936 ( .A1(n15591), .A2(n12669), .ZN(n15370) );
  OAI211_X1 U18937 ( .C1(n15372), .C2(n17671), .A(n15371), .B(n15370), .ZN(
        P1_U2970) );
  NAND2_X1 U18938 ( .A1(n15554), .A2(n15618), .ZN(n15392) );
  INV_X1 U18939 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15611) );
  MUX2_X1 U18940 ( .A(n15611), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .S(
        n15554), .Z(n15373) );
  XNOR2_X1 U18941 ( .A(n15374), .B(n15599), .ZN(n15606) );
  NOR2_X1 U18942 ( .A1(n15837), .A2(n22123), .ZN(n15601) );
  AOI21_X1 U18943 ( .B1(n17661), .B2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n15601), .ZN(n15375) );
  OAI21_X1 U18944 ( .B1(n15376), .B2(n17670), .A(n15375), .ZN(n15377) );
  AOI21_X1 U18945 ( .B1(n15378), .B2(n21328), .A(n15377), .ZN(n15379) );
  NOR2_X1 U18946 ( .A1(n15837), .A2(n21888), .ZN(n15610) );
  INV_X1 U18947 ( .A(n15380), .ZN(n15381) );
  NOR2_X1 U18948 ( .A1(n15381), .A2(n17670), .ZN(n15382) );
  AOI211_X1 U18949 ( .C1(n17661), .C2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n15610), .B(n15382), .ZN(n15388) );
  INV_X1 U18950 ( .A(n15384), .ZN(n15385) );
  NAND2_X1 U18951 ( .A1(n15402), .A2(n15385), .ZN(n15387) );
  NAND2_X1 U18952 ( .A1(n15390), .A2(n15650), .ZN(n15391) );
  INV_X1 U18953 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n15393) );
  NOR2_X1 U18954 ( .A1(n15837), .A2(n15393), .ZN(n15621) );
  AOI21_X1 U18955 ( .B1(n17661), .B2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n15621), .ZN(n15394) );
  OAI21_X1 U18956 ( .B1(n15395), .B2(n17670), .A(n15394), .ZN(n15396) );
  AOI21_X1 U18957 ( .B1(n15397), .B2(n21328), .A(n15396), .ZN(n15398) );
  NOR2_X1 U18958 ( .A1(n15837), .A2(n22130), .ZN(n15629) );
  NOR2_X1 U18959 ( .A1(n17676), .A2(n15399), .ZN(n15400) );
  AOI211_X1 U18960 ( .C1(n15401), .C2(n15576), .A(n15629), .B(n15400), .ZN(
        n15405) );
  NAND2_X1 U18961 ( .A1(n15626), .A2(n12669), .ZN(n15404) );
  OAI211_X1 U18962 ( .C1(n15406), .C2(n17671), .A(n15405), .B(n15404), .ZN(
        P1_U2974) );
  XNOR2_X1 U18963 ( .A(n15407), .B(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15645) );
  NOR2_X1 U18964 ( .A1(n15837), .A2(n15408), .ZN(n15640) );
  AOI21_X1 U18965 ( .B1(n17661), .B2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n15640), .ZN(n15409) );
  OAI21_X1 U18966 ( .B1(n15410), .B2(n17670), .A(n15409), .ZN(n15411) );
  AOI21_X1 U18967 ( .B1(n15412), .B2(n21328), .A(n15411), .ZN(n15413) );
  OAI21_X1 U18968 ( .B1(n21153), .B2(n15645), .A(n15413), .ZN(P1_U2975) );
  XNOR2_X1 U18969 ( .A(n15554), .B(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15414) );
  XNOR2_X1 U18970 ( .A(n15415), .B(n15414), .ZN(n15655) );
  NAND2_X1 U18971 ( .A1(n17697), .A2(P1_REIP_REG_23__SCAN_IN), .ZN(n15649) );
  OAI21_X1 U18972 ( .B1(n17676), .B2(n15416), .A(n15649), .ZN(n15419) );
  NOR2_X1 U18973 ( .A1(n15417), .A2(n17671), .ZN(n15418) );
  AOI211_X1 U18974 ( .C1(n15576), .C2(n15420), .A(n15419), .B(n15418), .ZN(
        n15421) );
  OAI21_X1 U18975 ( .B1(n15655), .B2(n21153), .A(n15421), .ZN(P1_U2976) );
  NAND2_X1 U18976 ( .A1(n15423), .A2(n15422), .ZN(n15425) );
  XNOR2_X1 U18977 ( .A(n15425), .B(n15424), .ZN(n15665) );
  NOR2_X1 U18978 ( .A1(n17670), .A2(n15426), .ZN(n15429) );
  OR2_X1 U18979 ( .A1(n15837), .A2(n15427), .ZN(n15656) );
  OAI21_X1 U18980 ( .B1(n17676), .B2(n21959), .A(n15656), .ZN(n15428) );
  AOI211_X1 U18981 ( .C1(n15430), .C2(n21328), .A(n15429), .B(n15428), .ZN(
        n15431) );
  OAI21_X1 U18982 ( .B1(n21153), .B2(n15665), .A(n15431), .ZN(P1_U2977) );
  NOR2_X1 U18983 ( .A1(n15837), .A2(n21882), .ZN(n15668) );
  NOR2_X1 U18984 ( .A1(n17676), .A2(n15432), .ZN(n15433) );
  AOI211_X1 U18985 ( .C1(n15576), .C2(n15434), .A(n15668), .B(n15433), .ZN(
        n15439) );
  MUX2_X1 U18986 ( .A(n15436), .B(n15435), .S(n15545), .Z(n15437) );
  XNOR2_X1 U18987 ( .A(n15437), .B(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15667) );
  NAND2_X1 U18988 ( .A1(n15667), .A2(n12669), .ZN(n15438) );
  OAI211_X1 U18989 ( .C1(n15440), .C2(n17671), .A(n15439), .B(n15438), .ZN(
        P1_U2978) );
  INV_X1 U18990 ( .A(n15441), .ZN(n15442) );
  NAND2_X1 U18991 ( .A1(n15442), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15443) );
  MUX2_X1 U18992 ( .A(n15444), .B(n15443), .S(n15554), .Z(n15445) );
  XOR2_X1 U18993 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .B(n15445), .Z(
        n15691) );
  NAND2_X1 U18994 ( .A1(n17697), .A2(P1_REIP_REG_20__SCAN_IN), .ZN(n15686) );
  NAND2_X1 U18995 ( .A1(n17661), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15446) );
  OAI211_X1 U18996 ( .C1(n17670), .C2(n15447), .A(n15686), .B(n15446), .ZN(
        n15448) );
  AOI21_X1 U18997 ( .B1(n15449), .B2(n21328), .A(n15448), .ZN(n15450) );
  OAI21_X1 U18998 ( .B1(n21153), .B2(n15691), .A(n15450), .ZN(P1_U2979) );
  NOR2_X1 U18999 ( .A1(n15554), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15451) );
  MUX2_X1 U19000 ( .A(n15554), .B(n15451), .S(n15441), .Z(n15452) );
  XNOR2_X1 U19001 ( .A(n15452), .B(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15700) );
  NAND2_X1 U19002 ( .A1(n17697), .A2(P1_REIP_REG_19__SCAN_IN), .ZN(n15692) );
  OAI21_X1 U19003 ( .B1(n17676), .B2(n10055), .A(n15692), .ZN(n15455) );
  NOR2_X1 U19004 ( .A1(n15453), .A2(n17671), .ZN(n15454) );
  AOI211_X1 U19005 ( .C1(n15576), .C2(n15456), .A(n15455), .B(n15454), .ZN(
        n15457) );
  OAI21_X1 U19006 ( .B1(n21153), .B2(n15700), .A(n15457), .ZN(P1_U2980) );
  NOR2_X1 U19007 ( .A1(n15837), .A2(n15458), .ZN(n15710) );
  NOR2_X1 U19008 ( .A1(n17670), .A2(n15459), .ZN(n15460) );
  AOI211_X1 U19009 ( .C1(n17661), .C2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n15710), .B(n15460), .ZN(n15464) );
  OR2_X1 U19010 ( .A1(n15462), .A2(n15461), .ZN(n15701) );
  NAND3_X1 U19011 ( .A1(n15701), .A2(n12669), .A3(n15441), .ZN(n15463) );
  OAI211_X1 U19012 ( .C1(n15465), .C2(n17671), .A(n15464), .B(n15463), .ZN(
        P1_U2981) );
  NAND2_X1 U19013 ( .A1(n15545), .A2(n15466), .ZN(n15470) );
  INV_X1 U19014 ( .A(n15468), .ZN(n15480) );
  MUX2_X1 U19015 ( .A(n15545), .B(n15470), .S(n15469), .Z(n15471) );
  XNOR2_X1 U19016 ( .A(n15471), .B(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15716) );
  NAND2_X1 U19017 ( .A1(n15716), .A2(n12669), .ZN(n15476) );
  NOR2_X1 U19018 ( .A1(n15837), .A2(n15472), .ZN(n15718) );
  NOR2_X1 U19019 ( .A1(n17670), .A2(n15473), .ZN(n15474) );
  AOI211_X1 U19020 ( .C1(n17661), .C2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n15718), .B(n15474), .ZN(n15475) );
  OAI211_X1 U19021 ( .C1(n17671), .C2(n15477), .A(n15476), .B(n15475), .ZN(
        P1_U2982) );
  INV_X1 U19022 ( .A(n15478), .ZN(n15506) );
  NOR2_X1 U19023 ( .A1(n15506), .A2(n15479), .ZN(n15494) );
  NOR2_X1 U19024 ( .A1(n15494), .A2(n15480), .ZN(n15482) );
  NOR2_X1 U19025 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15729) );
  NOR2_X1 U19026 ( .A1(n15482), .A2(n15729), .ZN(n15484) );
  OAI22_X1 U19027 ( .A1(n15484), .A2(n15483), .B1(n15482), .B2(n15481), .ZN(
        n15734) );
  NAND2_X1 U19028 ( .A1(n17697), .A2(P1_REIP_REG_16__SCAN_IN), .ZN(n15726) );
  OAI21_X1 U19029 ( .B1(n17676), .B2(n15485), .A(n15726), .ZN(n15488) );
  NOR2_X1 U19030 ( .A1(n15486), .A2(n17671), .ZN(n15487) );
  AOI211_X1 U19031 ( .C1(n15576), .C2(n15489), .A(n15488), .B(n15487), .ZN(
        n15490) );
  OAI21_X1 U19032 ( .B1(n21153), .B2(n15734), .A(n15490), .ZN(P1_U2983) );
  NOR2_X1 U19033 ( .A1(n15837), .A2(n15491), .ZN(n15737) );
  NOR2_X1 U19034 ( .A1(n17670), .A2(n15492), .ZN(n15493) );
  AOI211_X1 U19035 ( .C1(n17661), .C2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n15737), .B(n15493), .ZN(n15499) );
  AOI21_X1 U19036 ( .B1(n15545), .B2(n15495), .A(n15494), .ZN(n15497) );
  XNOR2_X1 U19037 ( .A(n15554), .B(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15496) );
  XNOR2_X1 U19038 ( .A(n15497), .B(n15496), .ZN(n15735) );
  NAND2_X1 U19039 ( .A1(n15735), .A2(n12669), .ZN(n15498) );
  OAI211_X1 U19040 ( .C1(n15500), .C2(n17671), .A(n15499), .B(n15498), .ZN(
        P1_U2984) );
  NOR2_X1 U19041 ( .A1(n15837), .A2(n15501), .ZN(n15749) );
  NOR2_X1 U19042 ( .A1(n17670), .A2(n15502), .ZN(n15503) );
  AOI211_X1 U19043 ( .C1(n17661), .C2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n15749), .B(n15503), .ZN(n15510) );
  OAI22_X1 U19044 ( .A1(n15506), .A2(n15505), .B1(n15554), .B2(n15504), .ZN(
        n15508) );
  XNOR2_X1 U19045 ( .A(n15554), .B(n15758), .ZN(n15507) );
  XNOR2_X1 U19046 ( .A(n15508), .B(n15507), .ZN(n15746) );
  NAND2_X1 U19047 ( .A1(n15746), .A2(n12669), .ZN(n15509) );
  OAI211_X1 U19048 ( .C1(n15511), .C2(n17671), .A(n15510), .B(n15509), .ZN(
        P1_U2985) );
  NOR2_X1 U19049 ( .A1(n15837), .A2(n21880), .ZN(n15774) );
  NOR2_X1 U19050 ( .A1(n17670), .A2(n15512), .ZN(n15513) );
  AOI211_X1 U19051 ( .C1(n17661), .C2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n15774), .B(n15513), .ZN(n15521) );
  AOI22_X1 U19052 ( .A1(n15542), .A2(n15516), .B1(n15545), .B2(n15515), .ZN(
        n15528) );
  AOI21_X1 U19053 ( .B1(n15545), .B2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n12596), .ZN(n15527) );
  NAND2_X1 U19054 ( .A1(n15528), .A2(n15527), .ZN(n15526) );
  NAND2_X1 U19055 ( .A1(n15526), .A2(n15517), .ZN(n15519) );
  XNOR2_X1 U19056 ( .A(n15519), .B(n15518), .ZN(n15763) );
  NAND2_X1 U19057 ( .A1(n15763), .A2(n12669), .ZN(n15520) );
  OAI211_X1 U19058 ( .C1(n15522), .C2(n17671), .A(n15521), .B(n15520), .ZN(
        P1_U2986) );
  INV_X1 U19059 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n15523) );
  NOR2_X1 U19060 ( .A1(n15837), .A2(n15523), .ZN(n15796) );
  NOR2_X1 U19061 ( .A1(n17670), .A2(n15524), .ZN(n15525) );
  AOI211_X1 U19062 ( .C1(n17661), .C2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n15796), .B(n15525), .ZN(n15530) );
  OAI21_X1 U19063 ( .B1(n15528), .B2(n15527), .A(n15526), .ZN(n15787) );
  NAND2_X1 U19064 ( .A1(n15787), .A2(n12669), .ZN(n15529) );
  OAI211_X1 U19065 ( .C1(n15531), .C2(n17671), .A(n15530), .B(n15529), .ZN(
        P1_U2987) );
  XNOR2_X1 U19066 ( .A(n15532), .B(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17658) );
  NOR2_X1 U19067 ( .A1(n17657), .A2(n17658), .ZN(n17656) );
  AOI21_X1 U19068 ( .B1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n15532), .A(
        n17656), .ZN(n15564) );
  NAND2_X1 U19069 ( .A1(n15554), .A2(n15533), .ZN(n15562) );
  NAND3_X1 U19070 ( .A1(n15543), .A2(n15545), .A3(n15534), .ZN(n15548) );
  NAND3_X1 U19071 ( .A1(n15542), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        n15554), .ZN(n15535) );
  NAND2_X1 U19072 ( .A1(n15548), .A2(n15535), .ZN(n15536) );
  XNOR2_X1 U19073 ( .A(n15536), .B(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n15811) );
  NAND2_X1 U19074 ( .A1(n17697), .A2(P1_REIP_REG_11__SCAN_IN), .ZN(n15803) );
  NAND2_X1 U19075 ( .A1(n17661), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n15537) );
  OAI211_X1 U19076 ( .C1(n17670), .C2(n15538), .A(n15803), .B(n15537), .ZN(
        n15539) );
  AOI21_X1 U19077 ( .B1(n15540), .B2(n21328), .A(n15539), .ZN(n15541) );
  OAI21_X1 U19078 ( .B1(n15811), .B2(n21153), .A(n15541), .ZN(P1_U2988) );
  XNOR2_X1 U19079 ( .A(n15542), .B(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15547) );
  INV_X1 U19080 ( .A(n15543), .ZN(n15544) );
  NAND2_X1 U19081 ( .A1(n15544), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15546) );
  MUX2_X1 U19082 ( .A(n15547), .B(n15546), .S(n15545), .Z(n15549) );
  NAND2_X1 U19083 ( .A1(n15549), .A2(n15548), .ZN(n15813) );
  NAND2_X1 U19084 ( .A1(n15813), .A2(n12669), .ZN(n15553) );
  NAND2_X1 U19085 ( .A1(n17697), .A2(P1_REIP_REG_10__SCAN_IN), .ZN(n15821) );
  OAI21_X1 U19086 ( .B1(n17676), .B2(n15550), .A(n15821), .ZN(n15551) );
  AOI21_X1 U19087 ( .B1(n15576), .B2(n17642), .A(n15551), .ZN(n15552) );
  OAI211_X1 U19088 ( .C1(n17671), .C2(n17649), .A(n15553), .B(n15552), .ZN(
        P1_U2989) );
  XNOR2_X1 U19089 ( .A(n15554), .B(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15555) );
  XNOR2_X1 U19090 ( .A(n15556), .B(n15555), .ZN(n15833) );
  NAND2_X1 U19091 ( .A1(n17697), .A2(P1_REIP_REG_9__SCAN_IN), .ZN(n15826) );
  OAI21_X1 U19092 ( .B1(n17676), .B2(n15557), .A(n15826), .ZN(n15559) );
  NOR2_X1 U19093 ( .A1(n21173), .A2(n17671), .ZN(n15558) );
  AOI211_X1 U19094 ( .C1(n15576), .C2(n21175), .A(n15559), .B(n15558), .ZN(
        n15560) );
  OAI21_X1 U19095 ( .B1(n15833), .B2(n21153), .A(n15560), .ZN(P1_U2990) );
  XNOR2_X1 U19096 ( .A(n15562), .B(n15561), .ZN(n15563) );
  XNOR2_X1 U19097 ( .A(n15564), .B(n15563), .ZN(n17687) );
  NAND2_X1 U19098 ( .A1(n17687), .A2(n12669), .ZN(n15568) );
  INV_X1 U19099 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n15565) );
  NOR2_X1 U19100 ( .A1(n15837), .A2(n15565), .ZN(n17680) );
  NOR2_X1 U19101 ( .A1(n17670), .A2(n21186), .ZN(n15566) );
  AOI211_X1 U19102 ( .C1(n17661), .C2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n17680), .B(n15566), .ZN(n15567) );
  OAI211_X1 U19103 ( .C1(n17671), .C2(n21184), .A(n15568), .B(n15567), .ZN(
        P1_U2991) );
  XNOR2_X1 U19104 ( .A(n15570), .B(n15569), .ZN(n15580) );
  AOI22_X1 U19105 ( .A1(n15580), .A2(n15579), .B1(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n15570), .ZN(n15573) );
  XNOR2_X1 U19106 ( .A(n15571), .B(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n15572) );
  XNOR2_X1 U19107 ( .A(n15573), .B(n15572), .ZN(n15848) );
  NAND2_X1 U19108 ( .A1(n15848), .A2(n12669), .ZN(n15578) );
  NOR2_X1 U19109 ( .A1(n15837), .A2(n21247), .ZN(n15853) );
  INV_X1 U19110 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n15574) );
  NOR2_X1 U19111 ( .A1(n17676), .A2(n15574), .ZN(n15575) );
  AOI211_X1 U19112 ( .C1(n15576), .C2(n21231), .A(n15853), .B(n15575), .ZN(
        n15577) );
  OAI211_X1 U19113 ( .C1(n17671), .C2(n21230), .A(n15578), .B(n15577), .ZN(
        P1_U2995) );
  XNOR2_X1 U19114 ( .A(n15580), .B(n15579), .ZN(n15865) );
  INV_X1 U19115 ( .A(n15581), .ZN(n21266) );
  NOR2_X1 U19116 ( .A1(n15837), .A2(n22140), .ZN(n15859) );
  AOI21_X1 U19117 ( .B1(n17661), .B2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n15859), .ZN(n15582) );
  OAI21_X1 U19118 ( .B1(n21262), .B2(n17670), .A(n15582), .ZN(n15583) );
  AOI21_X1 U19119 ( .B1(n21266), .B2(n21328), .A(n15583), .ZN(n15584) );
  OAI21_X1 U19120 ( .B1(n21153), .B2(n15865), .A(n15584), .ZN(P1_U2996) );
  INV_X1 U19121 ( .A(n15592), .ZN(n15585) );
  AOI21_X1 U19122 ( .B1(n15585), .B2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15586) );
  NAND2_X1 U19123 ( .A1(n15591), .A2(n17700), .ZN(n15597) );
  NOR2_X1 U19124 ( .A1(n15592), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15593) );
  AOI211_X1 U19125 ( .C1(n15595), .C2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n15594), .B(n15593), .ZN(n15596) );
  OAI211_X1 U19126 ( .C1(n15839), .C2(n15598), .A(n15597), .B(n15596), .ZN(
        P1_U3002) );
  XNOR2_X1 U19127 ( .A(n15599), .B(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15602) );
  NOR3_X1 U19128 ( .A1(n15616), .A2(n15608), .A3(n15599), .ZN(n15600) );
  AOI211_X1 U19129 ( .C1(n15612), .C2(n15602), .A(n15601), .B(n15600), .ZN(
        n15605) );
  NAND2_X1 U19130 ( .A1(n15603), .A2(n17698), .ZN(n15604) );
  OAI211_X1 U19131 ( .C1(n15606), .C2(n15864), .A(n15605), .B(n15604), .ZN(
        P1_U3003) );
  NAND2_X1 U19132 ( .A1(n15607), .A2(n17700), .ZN(n15614) );
  NOR3_X1 U19133 ( .A1(n15616), .A2(n15608), .A3(n15611), .ZN(n15609) );
  AOI211_X1 U19134 ( .C1(n15612), .C2(n15611), .A(n15610), .B(n15609), .ZN(
        n15613) );
  OAI211_X1 U19135 ( .C1(n15839), .C2(n15615), .A(n15614), .B(n15613), .ZN(
        P1_U3004) );
  INV_X1 U19136 ( .A(n15616), .ZN(n15623) );
  OAI21_X1 U19137 ( .B1(n15638), .B2(n15618), .A(n15617), .ZN(n15622) );
  NOR2_X1 U19138 ( .A1(n15619), .A2(n15839), .ZN(n15620) );
  AOI211_X1 U19139 ( .C1(n15623), .C2(n15622), .A(n15621), .B(n15620), .ZN(
        n15624) );
  OAI21_X1 U19140 ( .B1(n15625), .B2(n15864), .A(n15624), .ZN(P1_U3005) );
  NAND2_X1 U19141 ( .A1(n15626), .A2(n17700), .ZN(n15633) );
  NAND2_X1 U19142 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15628) );
  OAI21_X1 U19143 ( .B1(n15638), .B2(n15628), .A(n15627), .ZN(n15631) );
  AOI21_X1 U19144 ( .B1(n15631), .B2(n15630), .A(n15629), .ZN(n15632) );
  OAI211_X1 U19145 ( .C1(n15839), .C2(n15634), .A(n15633), .B(n15632), .ZN(
        P1_U3006) );
  INV_X1 U19146 ( .A(n15635), .ZN(n15636) );
  OAI21_X1 U19147 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n15637), .A(
        n15636), .ZN(n15641) );
  NOR3_X1 U19148 ( .A1(n15638), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        n15650), .ZN(n15639) );
  AOI211_X1 U19149 ( .C1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .C2(n15641), .A(
        n15640), .B(n15639), .ZN(n15644) );
  NAND2_X1 U19150 ( .A1(n15642), .A2(n17698), .ZN(n15643) );
  OAI211_X1 U19151 ( .C1(n15645), .C2(n15864), .A(n15644), .B(n15643), .ZN(
        P1_U3007) );
  INV_X1 U19152 ( .A(n15646), .ZN(n15653) );
  OR4_X1 U19153 ( .A1(n15695), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n15647), .A4(n15659), .ZN(n15648) );
  OAI211_X1 U19154 ( .C1(n15651), .C2(n15650), .A(n15649), .B(n15648), .ZN(
        n15652) );
  AOI21_X1 U19155 ( .B1(n15653), .B2(n17698), .A(n15652), .ZN(n15654) );
  OAI21_X1 U19156 ( .B1(n15655), .B2(n15864), .A(n15654), .ZN(P1_U3008) );
  INV_X1 U19157 ( .A(n15656), .ZN(n15657) );
  AOI21_X1 U19158 ( .B1(n15658), .B2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n15657), .ZN(n15661) );
  OAI211_X1 U19159 ( .C1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n15673), .B(n15659), .ZN(
        n15660) );
  OAI211_X1 U19160 ( .C1(n15662), .C2(n15839), .A(n15661), .B(n15660), .ZN(
        n15663) );
  INV_X1 U19161 ( .A(n15663), .ZN(n15664) );
  OAI21_X1 U19162 ( .B1(n15665), .B2(n15864), .A(n15664), .ZN(P1_U3009) );
  INV_X1 U19163 ( .A(n15666), .ZN(n15676) );
  NAND2_X1 U19164 ( .A1(n15667), .A2(n17700), .ZN(n15675) );
  INV_X1 U19165 ( .A(n15668), .ZN(n15669) );
  OAI21_X1 U19166 ( .B1(n15670), .B2(n15672), .A(n15669), .ZN(n15671) );
  AOI21_X1 U19167 ( .B1(n15673), .B2(n15672), .A(n15671), .ZN(n15674) );
  OAI211_X1 U19168 ( .C1(n15839), .C2(n15676), .A(n15675), .B(n15674), .ZN(
        P1_U3010) );
  NAND2_X1 U19169 ( .A1(n15677), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15687) );
  INV_X1 U19170 ( .A(n15694), .ZN(n15684) );
  NAND2_X1 U19171 ( .A1(n15788), .A2(n15678), .ZN(n15777) );
  NOR3_X1 U19172 ( .A1(n15764), .A2(n15777), .A3(n15679), .ZN(n15681) );
  NOR2_X1 U19173 ( .A1(n15681), .A2(n15680), .ZN(n15782) );
  AOI21_X1 U19174 ( .B1(n15782), .B2(n15682), .A(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15683) );
  OAI21_X1 U19175 ( .B1(n15684), .B2(n15683), .A(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15685) );
  OAI211_X1 U19176 ( .C1(n15695), .C2(n15687), .A(n15686), .B(n15685), .ZN(
        n15688) );
  AOI21_X1 U19177 ( .B1(n15689), .B2(n17698), .A(n15688), .ZN(n15690) );
  OAI21_X1 U19178 ( .B1(n15691), .B2(n15864), .A(n15690), .ZN(P1_U3011) );
  INV_X1 U19179 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15693) );
  OAI21_X1 U19180 ( .B1(n15694), .B2(n15693), .A(n15692), .ZN(n15697) );
  NOR2_X1 U19181 ( .A1(n15695), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15696) );
  AOI211_X1 U19182 ( .C1(n15698), .C2(n17698), .A(n15697), .B(n15696), .ZN(
        n15699) );
  OAI21_X1 U19183 ( .B1(n15700), .B2(n15864), .A(n15699), .ZN(P1_U3012) );
  NAND3_X1 U19184 ( .A1(n15701), .A2(n17700), .A3(n15441), .ZN(n15713) );
  INV_X1 U19185 ( .A(n15702), .ZN(n15711) );
  INV_X1 U19186 ( .A(n15703), .ZN(n15704) );
  AND2_X1 U19187 ( .A1(n17681), .A2(n15704), .ZN(n15705) );
  NOR2_X1 U19188 ( .A1(n15750), .A2(n15705), .ZN(n15723) );
  NAND2_X1 U19189 ( .A1(n15706), .A2(n15708), .ZN(n15707) );
  OAI21_X1 U19190 ( .B1(n15723), .B2(n15708), .A(n15707), .ZN(n15709) );
  AOI211_X1 U19191 ( .C1(n15711), .C2(n17698), .A(n15710), .B(n15709), .ZN(
        n15712) );
  NAND2_X1 U19192 ( .A1(n15713), .A2(n15712), .ZN(P1_U3013) );
  INV_X1 U19193 ( .A(n15731), .ZN(n15715) );
  AOI21_X1 U19194 ( .B1(n15740), .B2(n15715), .A(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15722) );
  NAND2_X1 U19195 ( .A1(n15716), .A2(n17700), .ZN(n15721) );
  INV_X1 U19196 ( .A(n15717), .ZN(n15719) );
  AOI21_X1 U19197 ( .B1(n15719), .B2(n17698), .A(n15718), .ZN(n15720) );
  OAI211_X1 U19198 ( .C1(n15723), .C2(n15722), .A(n15721), .B(n15720), .ZN(
        P1_U3014) );
  INV_X1 U19199 ( .A(n15750), .ZN(n15725) );
  NAND2_X1 U19200 ( .A1(n17681), .A2(n15758), .ZN(n15724) );
  NAND2_X1 U19201 ( .A1(n15725), .A2(n15724), .ZN(n15741) );
  OAI21_X1 U19202 ( .B1(n15727), .B2(n15839), .A(n15726), .ZN(n15728) );
  AOI21_X1 U19203 ( .B1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n15741), .A(
        n15728), .ZN(n15733) );
  INV_X1 U19204 ( .A(n15729), .ZN(n15730) );
  NAND3_X1 U19205 ( .A1(n15740), .A2(n15731), .A3(n15730), .ZN(n15732) );
  OAI211_X1 U19206 ( .C1(n15734), .C2(n15864), .A(n15733), .B(n15732), .ZN(
        P1_U3015) );
  NAND2_X1 U19207 ( .A1(n15735), .A2(n17700), .ZN(n15745) );
  INV_X1 U19208 ( .A(n15736), .ZN(n15738) );
  AOI21_X1 U19209 ( .B1(n15738), .B2(n17698), .A(n15737), .ZN(n15744) );
  NAND2_X1 U19210 ( .A1(n15740), .A2(n15739), .ZN(n15743) );
  NAND2_X1 U19211 ( .A1(n15741), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15742) );
  NAND4_X1 U19212 ( .A1(n15745), .A2(n15744), .A3(n15743), .A4(n15742), .ZN(
        P1_U3016) );
  INV_X1 U19213 ( .A(n15746), .ZN(n15762) );
  NOR2_X1 U19214 ( .A1(n15747), .A2(n15839), .ZN(n15748) );
  AOI211_X1 U19215 ( .C1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n15750), .A(
        n15749), .B(n15748), .ZN(n15761) );
  NOR2_X1 U19216 ( .A1(n15752), .A2(n15751), .ZN(n15815) );
  INV_X1 U19217 ( .A(n15815), .ZN(n15753) );
  NOR2_X1 U19218 ( .A1(n15793), .A2(n15753), .ZN(n17685) );
  AND2_X1 U19219 ( .A1(n15851), .A2(n15754), .ZN(n15755) );
  INV_X1 U19220 ( .A(n15855), .ZN(n15861) );
  INV_X1 U19221 ( .A(n15757), .ZN(n15759) );
  NAND3_X1 U19222 ( .A1(n17699), .A2(n15759), .A3(n15758), .ZN(n15760) );
  OAI211_X1 U19223 ( .C1(n15762), .C2(n15864), .A(n15761), .B(n15760), .ZN(
        P1_U3017) );
  INV_X1 U19224 ( .A(n15763), .ZN(n15786) );
  INV_X1 U19225 ( .A(n15764), .ZN(n15767) );
  AOI211_X1 U19226 ( .C1(n15777), .C2(n15767), .A(n15766), .B(n15765), .ZN(
        n15770) );
  NAND2_X1 U19227 ( .A1(n15769), .A2(n15768), .ZN(n15776) );
  OAI211_X1 U19228 ( .C1(n15772), .C2(n15771), .A(n15770), .B(n15776), .ZN(
        n15784) );
  INV_X1 U19229 ( .A(n15773), .ZN(n15775) );
  AOI21_X1 U19230 ( .B1(n15775), .B2(n17698), .A(n15774), .ZN(n15781) );
  INV_X1 U19231 ( .A(n15776), .ZN(n15779) );
  INV_X1 U19232 ( .A(n15777), .ZN(n15778) );
  NAND2_X1 U19233 ( .A1(n15779), .A2(n15778), .ZN(n15780) );
  OAI211_X1 U19234 ( .C1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .C2(n15782), .A(
        n15781), .B(n15780), .ZN(n15783) );
  AOI21_X1 U19235 ( .B1(n15784), .B2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n15783), .ZN(n15785) );
  OAI21_X1 U19236 ( .B1(n15786), .B2(n15864), .A(n15785), .ZN(P1_U3018) );
  INV_X1 U19237 ( .A(n15787), .ZN(n15802) );
  AND2_X1 U19238 ( .A1(n15808), .A2(n15788), .ZN(n15791) );
  INV_X1 U19239 ( .A(n15799), .ZN(n15789) );
  NAND2_X1 U19240 ( .A1(n15851), .A2(n15789), .ZN(n15790) );
  OAI211_X1 U19241 ( .C1(n15816), .C2(n15791), .A(n15840), .B(n15790), .ZN(
        n15806) );
  INV_X1 U19242 ( .A(n15806), .ZN(n15792) );
  OAI21_X1 U19243 ( .B1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n15793), .A(
        n15792), .ZN(n15797) );
  NOR2_X1 U19244 ( .A1(n15794), .A2(n15839), .ZN(n15795) );
  AOI211_X1 U19245 ( .C1(n15797), .C2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n15796), .B(n15795), .ZN(n15801) );
  NAND3_X1 U19246 ( .A1(n17699), .A2(n15799), .A3(n15798), .ZN(n15800) );
  OAI211_X1 U19247 ( .C1(n15802), .C2(n15864), .A(n15801), .B(n15800), .ZN(
        P1_U3019) );
  OAI21_X1 U19248 ( .B1(n15804), .B2(n15839), .A(n15803), .ZN(n15805) );
  AOI21_X1 U19249 ( .B1(n15806), .B2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n15805), .ZN(n15810) );
  NAND3_X1 U19250 ( .A1(n17699), .A2(n15808), .A3(n15807), .ZN(n15809) );
  OAI211_X1 U19251 ( .C1(n15811), .C2(n15864), .A(n15810), .B(n15809), .ZN(
        P1_U3020) );
  XNOR2_X1 U19252 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .B(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15825) );
  INV_X1 U19253 ( .A(n15818), .ZN(n15812) );
  NAND2_X1 U19254 ( .A1(n17699), .A2(n15812), .ZN(n15828) );
  NAND2_X1 U19255 ( .A1(n15813), .A2(n17700), .ZN(n15824) );
  OAI21_X1 U19256 ( .B1(n15816), .B2(n15815), .A(n15814), .ZN(n15849) );
  INV_X1 U19257 ( .A(n15849), .ZN(n15820) );
  OAI21_X1 U19258 ( .B1(n15818), .B2(n15817), .A(n17681), .ZN(n15819) );
  NAND2_X1 U19259 ( .A1(n15820), .A2(n15819), .ZN(n15831) );
  OAI21_X1 U19260 ( .B1(n15839), .B2(n17646), .A(n15821), .ZN(n15822) );
  AOI21_X1 U19261 ( .B1(n15831), .B2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n15822), .ZN(n15823) );
  OAI211_X1 U19262 ( .C1(n15825), .C2(n15828), .A(n15824), .B(n15823), .ZN(
        P1_U3021) );
  OAI21_X1 U19263 ( .B1(n15839), .B2(n15827), .A(n15826), .ZN(n15830) );
  NOR2_X1 U19264 ( .A1(n15828), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15829) );
  AOI211_X1 U19265 ( .C1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n15831), .A(
        n15830), .B(n15829), .ZN(n15832) );
  OAI21_X1 U19266 ( .B1(n15833), .B2(n15864), .A(n15832), .ZN(P1_U3022) );
  XOR2_X1 U19267 ( .A(n15834), .B(n15835), .Z(n17673) );
  INV_X1 U19268 ( .A(n17673), .ZN(n15847) );
  NOR2_X1 U19269 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n15854), .ZN(
        n17684) );
  OR2_X1 U19270 ( .A1(n15837), .A2(n15836), .ZN(n17674) );
  OAI21_X1 U19271 ( .B1(n15839), .B2(n15838), .A(n17674), .ZN(n15845) );
  INV_X1 U19272 ( .A(n15840), .ZN(n15841) );
  AOI21_X1 U19273 ( .B1(n15843), .B2(n15842), .A(n15841), .ZN(n17682) );
  NOR2_X1 U19274 ( .A1(n17682), .A2(n15756), .ZN(n15844) );
  AOI211_X1 U19275 ( .C1(n17684), .C2(n15855), .A(n15845), .B(n15844), .ZN(
        n15846) );
  OAI21_X1 U19276 ( .B1(n15847), .B2(n15864), .A(n15846), .ZN(P1_U3026) );
  INV_X1 U19277 ( .A(n15848), .ZN(n15858) );
  AOI21_X1 U19278 ( .B1(n15851), .B2(n15850), .A(n15849), .ZN(n15860) );
  NOR2_X1 U19279 ( .A1(n10095), .A2(n15860), .ZN(n15852) );
  AOI211_X1 U19280 ( .C1(n17698), .C2(n21232), .A(n15853), .B(n15852), .ZN(
        n15857) );
  OAI211_X1 U19281 ( .C1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(n15855), .B(n15854), .ZN(n15856) );
  OAI211_X1 U19282 ( .C1(n15858), .C2(n15864), .A(n15857), .B(n15856), .ZN(
        P1_U3027) );
  AOI21_X1 U19283 ( .B1(n17698), .B2(n21260), .A(n15859), .ZN(n15863) );
  MUX2_X1 U19284 ( .A(n15861), .B(n15860), .S(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .Z(n15862) );
  OAI211_X1 U19285 ( .C1(n15865), .C2(n15864), .A(n15863), .B(n15862), .ZN(
        P1_U3028) );
  NOR2_X1 U19286 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n21871), .ZN(n15868) );
  MUX2_X1 U19287 ( .A(n15866), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n17600), .Z(n17607) );
  AOI22_X1 U19288 ( .A1(n15868), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n21871), .B2(n17607), .ZN(n15870) );
  MUX2_X1 U19289 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n15867), .S(
        n15877), .Z(n17604) );
  AOI22_X1 U19290 ( .A1(n15868), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n17604), .B2(n21871), .ZN(n15869) );
  NOR2_X1 U19291 ( .A1(n15870), .A2(n15869), .ZN(n17615) );
  INV_X1 U19292 ( .A(n15871), .ZN(n15906) );
  NAND2_X1 U19293 ( .A1(n17615), .A2(n15906), .ZN(n15880) );
  NOR2_X1 U19294 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n15872), .ZN(n15875) );
  NAND2_X1 U19295 ( .A1(n15873), .A2(n15877), .ZN(n15874) );
  MUX2_X1 U19296 ( .A(n15875), .B(n15874), .S(n21871), .Z(n15876) );
  OAI21_X1 U19297 ( .B1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n15877), .A(
        n15876), .ZN(n17616) );
  AND3_X1 U19298 ( .A1(n15880), .A2(n22052), .A3(n17616), .ZN(n15879) );
  AND3_X1 U19299 ( .A1(n15880), .A2(n17710), .A3(n17616), .ZN(n17619) );
  NAND2_X1 U19300 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n21704), .ZN(n15898) );
  INV_X1 U19301 ( .A(n15898), .ZN(n15887) );
  OAI22_X1 U19302 ( .A1(n9734), .A2(n21810), .B1(n15881), .B2(n15887), .ZN(
        n15882) );
  OAI21_X1 U19303 ( .B1(n17619), .B2(n15882), .A(n21325), .ZN(n15883) );
  OAI21_X1 U19304 ( .B1(n21325), .B2(n21729), .A(n15883), .ZN(P1_U3478) );
  NAND2_X1 U19305 ( .A1(n15884), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n15895) );
  OAI21_X1 U19306 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n15884), .A(n21815), 
        .ZN(n15885) );
  OAI21_X1 U19307 ( .B1(n21702), .B2(n15887), .A(n15885), .ZN(n15886) );
  MUX2_X1 U19308 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n15886), .S(
        n21325), .Z(P1_U3477) );
  NOR2_X1 U19309 ( .A1(n13896), .A2(n15887), .ZN(n15891) );
  NOR2_X1 U19310 ( .A1(n15895), .A2(n21810), .ZN(n15889) );
  MUX2_X1 U19311 ( .A(n15889), .B(n21815), .S(n21330), .Z(n15890) );
  OAI21_X1 U19312 ( .B1(n15891), .B2(n15890), .A(n21325), .ZN(n15892) );
  OAI21_X1 U19313 ( .B1(n21325), .B2(n21586), .A(n15892), .ZN(P1_U3476) );
  INV_X1 U19314 ( .A(n21325), .ZN(n15903) );
  INV_X1 U19315 ( .A(n15893), .ZN(n15894) );
  OAI22_X1 U19316 ( .A1(n21776), .A2(n15884), .B1(n21561), .B2(n15895), .ZN(
        n15897) );
  NAND2_X1 U19317 ( .A1(n15897), .A2(n21584), .ZN(n15900) );
  AOI21_X1 U19318 ( .B1(n15896), .B2(n21905), .A(n21810), .ZN(n15899) );
  AOI22_X1 U19319 ( .A1(n15900), .A2(n15899), .B1(n15898), .B2(n21585), .ZN(
        n15902) );
  NAND2_X1 U19320 ( .A1(n15903), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n15901) );
  OAI21_X1 U19321 ( .B1(n15903), .B2(n15902), .A(n15901), .ZN(P1_U3475) );
  INV_X1 U19322 ( .A(n15904), .ZN(n15910) );
  INV_X1 U19323 ( .A(n12123), .ZN(n15905) );
  NAND2_X1 U19324 ( .A1(n15906), .A2(n15905), .ZN(n15912) );
  OAI22_X1 U19325 ( .A1(n15908), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B1(
        n15912), .B2(n15907), .ZN(n15909) );
  AOI21_X1 U19326 ( .B1(n21778), .B2(n15910), .A(n15909), .ZN(n17599) );
  INV_X1 U19327 ( .A(n15911), .ZN(n15918) );
  INV_X1 U19328 ( .A(n15912), .ZN(n15915) );
  AOI22_X1 U19329 ( .A1(n15916), .A2(n15915), .B1(n15914), .B2(n15913), .ZN(
        n15917) );
  OAI21_X1 U19330 ( .B1(n17599), .B2(n15918), .A(n15917), .ZN(n15920) );
  MUX2_X1 U19331 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n15920), .S(
        n15919), .Z(P1_U3473) );
  AOI21_X1 U19332 ( .B1(n21144), .B2(HOLD), .A(n15921), .ZN(n15926) );
  OAI21_X1 U19333 ( .B1(n21020), .B2(n15923), .A(n15922), .ZN(n15924) );
  NAND3_X1 U19334 ( .A1(n15926), .A2(n15925), .A3(n15924), .ZN(P1_U3195) );
  INV_X1 U19335 ( .A(n16394), .ZN(n15940) );
  INV_X1 U19336 ( .A(n15927), .ZN(n16306) );
  NAND2_X1 U19337 ( .A1(n16174), .A2(n15928), .ZN(n15936) );
  NAND2_X1 U19338 ( .A1(n15929), .A2(n9708), .ZN(n15935) );
  OAI22_X1 U19339 ( .A1(n20269), .A2(n15932), .B1(n15931), .B2(n15930), .ZN(
        n15933) );
  AOI21_X1 U19340 ( .B1(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n20240), .A(
        n15933), .ZN(n15934) );
  OAI211_X1 U19341 ( .C1(n15937), .C2(n15936), .A(n15935), .B(n15934), .ZN(
        n15938) );
  AOI21_X1 U19342 ( .B1(n16306), .B2(n20242), .A(n15938), .ZN(n15939) );
  OAI21_X1 U19343 ( .B1(n15940), .B2(n20276), .A(n15939), .ZN(P2_U2824) );
  NAND2_X1 U19344 ( .A1(n16397), .A2(n20244), .ZN(n15951) );
  AOI21_X1 U19345 ( .B1(n15941), .B2(n20227), .A(n16299), .ZN(n15942) );
  NOR2_X1 U19346 ( .A1(n15942), .A2(n15943), .ZN(n15948) );
  NAND3_X1 U19347 ( .A1(n15944), .A2(n16174), .A3(n15943), .ZN(n15946) );
  AOI22_X1 U19348 ( .A1(n20256), .A2(P2_REIP_REG_29__SCAN_IN), .B1(
        P2_EBX_REG_29__SCAN_IN), .B2(n20271), .ZN(n15945) );
  OAI211_X1 U19349 ( .C1(n20260), .C2(n10416), .A(n15946), .B(n15945), .ZN(
        n15947) );
  OAI211_X1 U19350 ( .C1(n20277), .C2(n16310), .A(n15951), .B(n15950), .ZN(
        P2_U2826) );
  OR2_X1 U19351 ( .A1(n15952), .A2(n15953), .ZN(n15954) );
  INV_X1 U19352 ( .A(n15956), .ZN(n15971) );
  AOI21_X1 U19353 ( .B1(n15958), .B2(n15971), .A(n15957), .ZN(n16763) );
  XNOR2_X1 U19354 ( .A(n15959), .B(n16531), .ZN(n15965) );
  NAND2_X1 U19355 ( .A1(n15960), .A2(n9708), .ZN(n15964) );
  OAI22_X1 U19356 ( .A1(n16528), .A2(n20269), .B1(n20231), .B2(n15961), .ZN(
        n15962) );
  AOI21_X1 U19357 ( .B1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n20240), .A(
        n15962), .ZN(n15963) );
  OAI211_X1 U19358 ( .C1(n21006), .C2(n15965), .A(n15964), .B(n15963), .ZN(
        n15966) );
  AOI21_X1 U19359 ( .B1(n16763), .B2(n20242), .A(n15966), .ZN(n15967) );
  OAI21_X1 U19360 ( .B1(n16770), .B2(n20276), .A(n15967), .ZN(P2_U2827) );
  INV_X1 U19361 ( .A(n15952), .ZN(n15969) );
  OAI21_X1 U19362 ( .B1(n15968), .B2(n15970), .A(n15969), .ZN(n16779) );
  AOI21_X1 U19363 ( .B1(n15972), .B2(n10533), .A(n15956), .ZN(n16782) );
  OAI21_X1 U19364 ( .B1(n15973), .B2(n21006), .A(n16261), .ZN(n15977) );
  INV_X1 U19365 ( .A(n15978), .ZN(n16535) );
  NAND3_X1 U19366 ( .A1(n15973), .A2(n16174), .A3(n16535), .ZN(n15975) );
  AOI22_X1 U19367 ( .A1(n20256), .A2(P2_REIP_REG_27__SCAN_IN), .B1(
        P2_EBX_REG_27__SCAN_IN), .B2(n20271), .ZN(n15974) );
  OAI211_X1 U19368 ( .C1(n20260), .C2(n16536), .A(n15975), .B(n15974), .ZN(
        n15976) );
  AOI21_X1 U19369 ( .B1(n15978), .B2(n15977), .A(n15976), .ZN(n15979) );
  OAI21_X1 U19370 ( .B1(n15980), .B2(n20273), .A(n15979), .ZN(n15981) );
  AOI21_X1 U19371 ( .B1(n16782), .B2(n20242), .A(n15981), .ZN(n15982) );
  OAI21_X1 U19372 ( .B1(n16779), .B2(n20276), .A(n15982), .ZN(P2_U2828) );
  OR2_X1 U19373 ( .A1(n15983), .A2(n15984), .ZN(n15985) );
  NAND2_X1 U19374 ( .A1(n10533), .A2(n15985), .ZN(n16794) );
  AND2_X1 U19375 ( .A1(n9781), .A2(n15986), .ZN(n15987) );
  NOR2_X1 U19376 ( .A1(n15968), .A2(n15987), .ZN(n16797) );
  NAND2_X1 U19377 ( .A1(n16797), .A2(n20244), .ZN(n15995) );
  XNOR2_X1 U19378 ( .A(n15988), .B(n16548), .ZN(n15991) );
  AOI22_X1 U19379 ( .A1(n20256), .A2(P2_REIP_REG_26__SCAN_IN), .B1(
        P2_EBX_REG_26__SCAN_IN), .B2(n20271), .ZN(n15990) );
  NAND2_X1 U19380 ( .A1(n20240), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15989) );
  OAI211_X1 U19381 ( .C1(n15991), .C2(n21006), .A(n15990), .B(n15989), .ZN(
        n15992) );
  AOI21_X1 U19382 ( .B1(n15993), .B2(n9708), .A(n15992), .ZN(n15994) );
  OAI211_X1 U19383 ( .C1(n20277), .C2(n16794), .A(n15995), .B(n15994), .ZN(
        P2_U2829) );
  XNOR2_X1 U19384 ( .A(n15996), .B(n15997), .ZN(n16806) );
  AOI21_X1 U19385 ( .B1(n15999), .B2(n15998), .A(n15983), .ZN(n16799) );
  XNOR2_X1 U19386 ( .A(n11438), .B(P2_EBX_REG_25__SCAN_IN), .ZN(n16007) );
  OAI21_X1 U19387 ( .B1(n16000), .B2(n21006), .A(n16261), .ZN(n16004) );
  NAND3_X1 U19388 ( .A1(n16000), .A2(n16174), .A3(n11778), .ZN(n16002) );
  AOI22_X1 U19389 ( .A1(n20256), .A2(P2_REIP_REG_25__SCAN_IN), .B1(
        P2_EBX_REG_25__SCAN_IN), .B2(n20271), .ZN(n16001) );
  OAI211_X1 U19390 ( .C1(n20260), .C2(n22107), .A(n16002), .B(n16001), .ZN(
        n16003) );
  AOI21_X1 U19391 ( .B1(n16005), .B2(n16004), .A(n16003), .ZN(n16006) );
  OAI21_X1 U19392 ( .B1(n16007), .B2(n20273), .A(n16006), .ZN(n16008) );
  AOI21_X1 U19393 ( .B1(n16799), .B2(n20242), .A(n16008), .ZN(n16009) );
  OAI21_X1 U19394 ( .B1(n16806), .B2(n20276), .A(n16009), .ZN(P2_U2830) );
  OR2_X1 U19395 ( .A1(n16027), .A2(n16010), .ZN(n16011) );
  NAND2_X1 U19396 ( .A1(n15996), .A2(n16011), .ZN(n16818) );
  INV_X1 U19397 ( .A(n15998), .ZN(n16013) );
  AOI21_X1 U19398 ( .B1(n16014), .B2(n16012), .A(n16013), .ZN(n16816) );
  XNOR2_X1 U19399 ( .A(n11431), .B(P2_EBX_REG_24__SCAN_IN), .ZN(n16021) );
  XOR2_X1 U19400 ( .A(n16565), .B(n16015), .Z(n16019) );
  AOI22_X1 U19401 ( .A1(n20256), .A2(P2_REIP_REG_24__SCAN_IN), .B1(
        P2_EBX_REG_24__SCAN_IN), .B2(n20271), .ZN(n16016) );
  OAI21_X1 U19402 ( .B1(n20260), .B2(n16017), .A(n16016), .ZN(n16018) );
  AOI21_X1 U19403 ( .B1(n16019), .B2(n20227), .A(n16018), .ZN(n16020) );
  OAI21_X1 U19404 ( .B1(n16021), .B2(n20273), .A(n16020), .ZN(n16022) );
  AOI21_X1 U19405 ( .B1(n16816), .B2(n20242), .A(n16022), .ZN(n16023) );
  OAI21_X1 U19406 ( .B1(n16818), .B2(n20276), .A(n16023), .ZN(P2_U2831) );
  OAI21_X1 U19407 ( .B1(n9741), .B2(n16024), .A(n16012), .ZN(n16827) );
  AND2_X1 U19408 ( .A1(n16048), .A2(n16025), .ZN(n16026) );
  NOR2_X1 U19409 ( .A1(n16027), .A2(n16026), .ZN(n16830) );
  NAND2_X1 U19410 ( .A1(n16830), .A2(n20244), .ZN(n16038) );
  AOI21_X1 U19411 ( .B1(n16028), .B2(n20227), .A(n16299), .ZN(n16029) );
  NOR2_X1 U19412 ( .A1(n16029), .A2(n16572), .ZN(n16035) );
  INV_X1 U19413 ( .A(n16028), .ZN(n16030) );
  NAND3_X1 U19414 ( .A1(n16030), .A2(n16174), .A3(n16572), .ZN(n16032) );
  AOI22_X1 U19415 ( .A1(n20256), .A2(P2_REIP_REG_23__SCAN_IN), .B1(
        P2_EBX_REG_23__SCAN_IN), .B2(n20271), .ZN(n16031) );
  OAI211_X1 U19416 ( .C1(n20260), .C2(n16033), .A(n16032), .B(n16031), .ZN(
        n16034) );
  AOI211_X1 U19417 ( .C1(n16036), .C2(n9708), .A(n16035), .B(n16034), .ZN(
        n16037) );
  OAI211_X1 U19418 ( .C1(n16827), .C2(n20277), .A(n16038), .B(n16037), .ZN(
        P2_U2832) );
  AOI21_X1 U19419 ( .B1(n16039), .B2(n16055), .A(n9741), .ZN(n16836) );
  INV_X1 U19420 ( .A(n16836), .ZN(n16053) );
  XNOR2_X1 U19421 ( .A(n16040), .B(n16583), .ZN(n16044) );
  INV_X1 U19422 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n16581) );
  OAI22_X1 U19423 ( .A1(n16581), .A2(n20269), .B1(n20231), .B2(n16041), .ZN(
        n16042) );
  AOI21_X1 U19424 ( .B1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n20240), .A(
        n16042), .ZN(n16043) );
  OAI21_X1 U19425 ( .B1(n16044), .B2(n21006), .A(n16043), .ZN(n16045) );
  AOI21_X1 U19426 ( .B1(n16046), .B2(n9708), .A(n16045), .ZN(n16052) );
  INV_X1 U19427 ( .A(n16048), .ZN(n16049) );
  AOI21_X1 U19428 ( .B1(n16050), .B2(n16047), .A(n16049), .ZN(n16844) );
  NAND2_X1 U19429 ( .A1(n16844), .A2(n20244), .ZN(n16051) );
  OAI211_X1 U19430 ( .C1(n16053), .C2(n20277), .A(n16052), .B(n16051), .ZN(
        P2_U2833) );
  OAI21_X1 U19431 ( .B1(n16054), .B2(n9868), .A(n16055), .ZN(n16854) );
  INV_X1 U19432 ( .A(n16047), .ZN(n16058) );
  AOI21_X1 U19433 ( .B1(n16059), .B2(n16057), .A(n16058), .ZN(n16857) );
  NAND2_X1 U19434 ( .A1(n16857), .A2(n20244), .ZN(n16070) );
  INV_X1 U19435 ( .A(n16060), .ZN(n16061) );
  AOI21_X1 U19436 ( .B1(n16061), .B2(n20227), .A(n16299), .ZN(n16062) );
  NOR2_X1 U19437 ( .A1(n16062), .A2(n16595), .ZN(n16067) );
  INV_X1 U19438 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n16065) );
  AOI22_X1 U19439 ( .A1(n20256), .A2(P2_REIP_REG_21__SCAN_IN), .B1(
        P2_EBX_REG_21__SCAN_IN), .B2(n20271), .ZN(n16064) );
  NAND3_X1 U19440 ( .A1(n16174), .A2(n16060), .A3(n16595), .ZN(n16063) );
  OAI211_X1 U19441 ( .C1(n20260), .C2(n16065), .A(n16064), .B(n16063), .ZN(
        n16066) );
  AOI211_X1 U19442 ( .C1(n16068), .C2(n9708), .A(n16067), .B(n16066), .ZN(
        n16069) );
  OAI211_X1 U19443 ( .C1(n20277), .C2(n16854), .A(n16070), .B(n16069), .ZN(
        P2_U2834) );
  OAI21_X1 U19444 ( .B1(n16071), .B2(n16072), .A(n16057), .ZN(n16874) );
  AOI21_X1 U19445 ( .B1(n16073), .B2(n12104), .A(n16054), .ZN(n16872) );
  NAND2_X1 U19446 ( .A1(n16872), .A2(n20242), .ZN(n16081) );
  XNOR2_X1 U19447 ( .A(n16074), .B(n16609), .ZN(n16077) );
  AOI22_X1 U19448 ( .A1(n20256), .A2(P2_REIP_REG_20__SCAN_IN), .B1(
        P2_EBX_REG_20__SCAN_IN), .B2(n20271), .ZN(n16076) );
  NAND2_X1 U19449 ( .A1(n20240), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n16075) );
  OAI211_X1 U19450 ( .C1(n16077), .C2(n21006), .A(n16076), .B(n16075), .ZN(
        n16078) );
  AOI21_X1 U19451 ( .B1(n16079), .B2(n9708), .A(n16078), .ZN(n16080) );
  OAI211_X1 U19452 ( .C1(n20276), .C2(n16874), .A(n16081), .B(n16080), .ZN(
        P2_U2835) );
  NOR2_X1 U19453 ( .A1(n16082), .A2(n16083), .ZN(n16084) );
  OR2_X1 U19454 ( .A1(n16071), .A2(n16084), .ZN(n16887) );
  AOI21_X1 U19455 ( .B1(n20227), .B2(n16087), .A(n16299), .ZN(n16094) );
  NAND2_X1 U19456 ( .A1(n16085), .A2(n9708), .ZN(n16092) );
  AOI21_X1 U19457 ( .B1(n20271), .B2(P2_EBX_REG_19__SCAN_IN), .A(n20355), .ZN(
        n16086) );
  OAI21_X1 U19458 ( .B1(n20269), .B2(n21061), .A(n16086), .ZN(n16090) );
  INV_X1 U19459 ( .A(n16093), .ZN(n16088) );
  NOR3_X1 U19460 ( .A1(n16302), .A2(n16088), .A3(n16087), .ZN(n16089) );
  AOI211_X1 U19461 ( .C1(n20240), .C2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n16090), .B(n16089), .ZN(n16091) );
  OAI211_X1 U19462 ( .C1(n16094), .C2(n16093), .A(n16092), .B(n16091), .ZN(
        n16095) );
  AOI21_X1 U19463 ( .B1(n16880), .B2(n20242), .A(n16095), .ZN(n16096) );
  OAI21_X1 U19464 ( .B1(n16887), .B2(n20276), .A(n16096), .ZN(P2_U2836) );
  AND2_X1 U19465 ( .A1(n9794), .A2(n16097), .ZN(n16098) );
  OR2_X1 U19466 ( .A1(n16098), .A2(n12105), .ZN(n16902) );
  AND2_X1 U19467 ( .A1(n16099), .A2(n16100), .ZN(n16101) );
  NOR2_X1 U19468 ( .A1(n16082), .A2(n16101), .ZN(n16899) );
  NAND2_X1 U19469 ( .A1(n16899), .A2(n20244), .ZN(n16115) );
  INV_X1 U19470 ( .A(n16619), .ZN(n16111) );
  INV_X1 U19471 ( .A(n16102), .ZN(n16104) );
  NAND2_X1 U19472 ( .A1(n16174), .A2(n16104), .ZN(n16120) );
  INV_X1 U19473 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n16618) );
  NAND2_X1 U19474 ( .A1(n16104), .A2(n16103), .ZN(n16105) );
  NAND3_X1 U19475 ( .A1(n16105), .A2(n20227), .A3(n16111), .ZN(n16106) );
  NAND2_X1 U19476 ( .A1(n16106), .A2(n20217), .ZN(n16107) );
  AOI21_X1 U19477 ( .B1(n20271), .B2(P2_EBX_REG_18__SCAN_IN), .A(n16107), .ZN(
        n16108) );
  OAI21_X1 U19478 ( .B1(n20269), .B2(n16618), .A(n16108), .ZN(n16109) );
  AOI21_X1 U19479 ( .B1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n20240), .A(
        n16109), .ZN(n16110) );
  OAI21_X1 U19480 ( .B1(n16111), .B2(n16120), .A(n16110), .ZN(n16112) );
  AOI21_X1 U19481 ( .B1(n16113), .B2(n9708), .A(n16112), .ZN(n16114) );
  OAI211_X1 U19482 ( .C1(n16902), .C2(n20277), .A(n16115), .B(n16114), .ZN(
        P2_U2837) );
  NAND2_X1 U19483 ( .A1(n9792), .A2(n16116), .ZN(n16117) );
  NAND2_X1 U19484 ( .A1(n9794), .A2(n16117), .ZN(n16910) );
  INV_X1 U19485 ( .A(n16099), .ZN(n16118) );
  AOI21_X1 U19486 ( .B1(n16119), .B2(n14766), .A(n16118), .ZN(n16917) );
  NAND2_X1 U19487 ( .A1(n16917), .A2(n20244), .ZN(n16130) );
  INV_X1 U19488 ( .A(n16629), .ZN(n16122) );
  AOI21_X1 U19489 ( .B1(n16122), .B2(n16121), .A(n16120), .ZN(n16127) );
  INV_X1 U19490 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n21058) );
  AOI21_X1 U19491 ( .B1(n20271), .B2(P2_EBX_REG_17__SCAN_IN), .A(n20355), .ZN(
        n16123) );
  OAI21_X1 U19492 ( .B1(n20269), .B2(n21058), .A(n16123), .ZN(n16124) );
  AOI21_X1 U19493 ( .B1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n20240), .A(
        n16124), .ZN(n16125) );
  OAI21_X1 U19494 ( .B1(n16629), .B2(n16261), .A(n16125), .ZN(n16126) );
  AOI211_X1 U19495 ( .C1(n16128), .C2(n9708), .A(n16127), .B(n16126), .ZN(
        n16129) );
  OAI211_X1 U19496 ( .C1(n20277), .C2(n16910), .A(n16130), .B(n16129), .ZN(
        P2_U2838) );
  INV_X1 U19497 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n21055) );
  AOI21_X1 U19498 ( .B1(n20271), .B2(P2_EBX_REG_15__SCAN_IN), .A(n20355), .ZN(
        n16131) );
  OAI21_X1 U19499 ( .B1(n20269), .B2(n21055), .A(n16131), .ZN(n16132) );
  AOI21_X1 U19500 ( .B1(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n20240), .A(
        n16132), .ZN(n16138) );
  NAND2_X1 U19501 ( .A1(n20250), .A2(n16133), .ZN(n16135) );
  XNOR2_X1 U19502 ( .A(n16135), .B(n16134), .ZN(n16136) );
  NAND2_X1 U19503 ( .A1(n16136), .A2(n20227), .ZN(n16137) );
  OAI211_X1 U19504 ( .C1(n16139), .C2(n20273), .A(n16138), .B(n16137), .ZN(
        n16140) );
  AOI21_X1 U19505 ( .B1(n16922), .B2(n20242), .A(n16140), .ZN(n16141) );
  OAI21_X1 U19506 ( .B1(n16921), .B2(n20276), .A(n16141), .ZN(P2_U2840) );
  AOI21_X1 U19507 ( .B1(n20227), .B2(n16145), .A(n16299), .ZN(n16151) );
  NAND2_X1 U19508 ( .A1(n16142), .A2(n9708), .ZN(n16150) );
  INV_X1 U19509 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n16144) );
  AOI21_X1 U19510 ( .B1(n20271), .B2(P2_EBX_REG_13__SCAN_IN), .A(n20355), .ZN(
        n16143) );
  OAI21_X1 U19511 ( .B1(n20269), .B2(n16144), .A(n16143), .ZN(n16148) );
  INV_X1 U19512 ( .A(n16669), .ZN(n16146) );
  NOR3_X1 U19513 ( .A1(n16302), .A2(n16146), .A3(n16145), .ZN(n16147) );
  AOI211_X1 U19514 ( .C1(n20240), .C2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n16148), .B(n16147), .ZN(n16149) );
  OAI211_X1 U19515 ( .C1(n16151), .C2(n16669), .A(n16150), .B(n16149), .ZN(
        n16152) );
  AOI21_X1 U19516 ( .B1(n16960), .B2(n20242), .A(n16152), .ZN(n16153) );
  OAI21_X1 U19517 ( .B1(n20276), .B2(n16957), .A(n16153), .ZN(P2_U2842) );
  INV_X1 U19518 ( .A(n14346), .ZN(n16156) );
  NAND2_X1 U19519 ( .A1(n14309), .A2(n16154), .ZN(n16155) );
  NAND2_X1 U19520 ( .A1(n16156), .A2(n16155), .ZN(n16969) );
  INV_X1 U19521 ( .A(n16969), .ZN(n16167) );
  OAI21_X1 U19522 ( .B1(n21006), .B2(n16172), .A(n16261), .ZN(n16162) );
  INV_X1 U19523 ( .A(n16172), .ZN(n16157) );
  NOR3_X1 U19524 ( .A1(n16302), .A2(n16163), .A3(n16157), .ZN(n16161) );
  INV_X1 U19525 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n21050) );
  NAND2_X1 U19526 ( .A1(n20240), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n16159) );
  AOI21_X1 U19527 ( .B1(n20271), .B2(P2_EBX_REG_12__SCAN_IN), .A(n20355), .ZN(
        n16158) );
  OAI211_X1 U19528 ( .C1(n21050), .C2(n20269), .A(n16159), .B(n16158), .ZN(
        n16160) );
  AOI211_X1 U19529 ( .C1(n16163), .C2(n16162), .A(n16161), .B(n16160), .ZN(
        n16164) );
  OAI21_X1 U19530 ( .B1(n16165), .B2(n20273), .A(n16164), .ZN(n16166) );
  AOI21_X1 U19531 ( .B1(n16167), .B2(n20242), .A(n16166), .ZN(n16168) );
  OAI21_X1 U19532 ( .B1(n20276), .B2(n16964), .A(n16168), .ZN(P2_U2843) );
  NAND2_X1 U19533 ( .A1(n16975), .A2(n20244), .ZN(n16181) );
  INV_X1 U19534 ( .A(n16697), .ZN(n16177) );
  INV_X1 U19535 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n16694) );
  AOI21_X1 U19536 ( .B1(n20271), .B2(P2_EBX_REG_11__SCAN_IN), .A(n20355), .ZN(
        n16169) );
  OAI21_X1 U19537 ( .B1(n20269), .B2(n16694), .A(n16169), .ZN(n16170) );
  AOI21_X1 U19538 ( .B1(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n20240), .A(
        n16170), .ZN(n16176) );
  NAND2_X1 U19539 ( .A1(n16697), .A2(n16171), .ZN(n16173) );
  NAND3_X1 U19540 ( .A1(n16174), .A2(n16173), .A3(n16172), .ZN(n16175) );
  OAI211_X1 U19541 ( .C1(n16261), .C2(n16177), .A(n16176), .B(n16175), .ZN(
        n16178) );
  AOI21_X1 U19542 ( .B1(n16179), .B2(n9708), .A(n16178), .ZN(n16180) );
  OAI211_X1 U19543 ( .C1(n16982), .C2(n20277), .A(n16181), .B(n16180), .ZN(
        P2_U2844) );
  INV_X1 U19544 ( .A(n16987), .ZN(n16193) );
  AOI21_X1 U19545 ( .B1(n20227), .B2(n16183), .A(n16299), .ZN(n16188) );
  INV_X1 U19546 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n22182) );
  AOI21_X1 U19547 ( .B1(n20271), .B2(P2_EBX_REG_10__SCAN_IN), .A(n20355), .ZN(
        n16182) );
  OAI21_X1 U19548 ( .B1(n20269), .B2(n22182), .A(n16182), .ZN(n16186) );
  INV_X1 U19549 ( .A(n16707), .ZN(n16184) );
  NOR3_X1 U19550 ( .A1(n16302), .A2(n16184), .A3(n16183), .ZN(n16185) );
  AOI211_X1 U19551 ( .C1(n20240), .C2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n16186), .B(n16185), .ZN(n16187) );
  OAI21_X1 U19552 ( .B1(n16188), .B2(n16707), .A(n16187), .ZN(n16189) );
  AOI21_X1 U19553 ( .B1(n16190), .B2(n9708), .A(n16189), .ZN(n16192) );
  NAND2_X1 U19554 ( .A1(n16995), .A2(n20244), .ZN(n16191) );
  OAI211_X1 U19555 ( .C1(n16193), .C2(n20277), .A(n16192), .B(n16191), .ZN(
        P2_U2845) );
  NAND2_X1 U19556 ( .A1(n13809), .A2(n16194), .ZN(n16195) );
  AND2_X1 U19557 ( .A1(n9771), .A2(n16195), .ZN(n20285) );
  INV_X1 U19558 ( .A(n20285), .ZN(n16211) );
  NOR2_X1 U19559 ( .A1(n16197), .A2(n16196), .ZN(n16198) );
  OR2_X1 U19560 ( .A1(n14337), .A2(n16198), .ZN(n17031) );
  INV_X1 U19561 ( .A(n17031), .ZN(n16734) );
  NAND2_X1 U19562 ( .A1(n20250), .A2(n16199), .ZN(n20268) );
  OAI22_X1 U19563 ( .A1(n16302), .A2(n16200), .B1(n21006), .B2(n20268), .ZN(
        n16206) );
  AND2_X1 U19564 ( .A1(n20227), .A2(n16214), .ZN(n16212) );
  NAND3_X1 U19565 ( .A1(n16757), .A2(n16212), .A3(n16200), .ZN(n16201) );
  AOI21_X1 U19566 ( .B1(n16261), .B2(n16201), .A(n16732), .ZN(n16205) );
  INV_X1 U19567 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n21044) );
  NAND2_X1 U19568 ( .A1(n20240), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16203) );
  AOI21_X1 U19569 ( .B1(n20271), .B2(P2_EBX_REG_8__SCAN_IN), .A(n20355), .ZN(
        n16202) );
  OAI211_X1 U19570 ( .C1(n20269), .C2(n21044), .A(n16203), .B(n16202), .ZN(
        n16204) );
  AOI211_X1 U19571 ( .C1(n16732), .C2(n16206), .A(n16205), .B(n16204), .ZN(
        n16207) );
  OAI21_X1 U19572 ( .B1(n16208), .B2(n20273), .A(n16207), .ZN(n16209) );
  AOI21_X1 U19573 ( .B1(n16734), .B2(n20242), .A(n16209), .ZN(n16210) );
  OAI21_X1 U19574 ( .B1(n20276), .B2(n16211), .A(n16210), .ZN(P2_U2847) );
  NAND2_X1 U19575 ( .A1(n17051), .A2(n20244), .ZN(n16223) );
  NOR2_X1 U19576 ( .A1(n16299), .A2(n16212), .ZN(n16219) );
  AOI21_X1 U19577 ( .B1(n20271), .B2(P2_EBX_REG_6__SCAN_IN), .A(n20355), .ZN(
        n16213) );
  OAI21_X1 U19578 ( .B1(n20269), .B2(n21040), .A(n16213), .ZN(n16217) );
  INV_X1 U19579 ( .A(n16757), .ZN(n16215) );
  NOR3_X1 U19580 ( .A1(n16302), .A2(n16215), .A3(n16214), .ZN(n16216) );
  AOI211_X1 U19581 ( .C1(n20240), .C2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n16217), .B(n16216), .ZN(n16218) );
  OAI21_X1 U19582 ( .B1(n16219), .B2(n16757), .A(n16218), .ZN(n16220) );
  AOI21_X1 U19583 ( .B1(n9708), .B2(n16221), .A(n16220), .ZN(n16222) );
  OAI211_X1 U19584 ( .C1(n17054), .C2(n20277), .A(n16223), .B(n16222), .ZN(
        P2_U2849) );
  OR2_X1 U19585 ( .A1(n16225), .A2(n16224), .ZN(n16226) );
  NAND2_X1 U19586 ( .A1(n16227), .A2(n16226), .ZN(n17079) );
  INV_X1 U19587 ( .A(n16228), .ZN(n17718) );
  OAI21_X1 U19588 ( .B1(n16229), .B2(n21006), .A(n16261), .ZN(n16235) );
  INV_X1 U19589 ( .A(n16229), .ZN(n16230) );
  NOR3_X1 U19590 ( .A1(n16302), .A2(n17717), .A3(n16230), .ZN(n16234) );
  INV_X1 U19591 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n21038) );
  NAND2_X1 U19592 ( .A1(n20240), .A2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n16232) );
  AOI21_X1 U19593 ( .B1(n20271), .B2(P2_EBX_REG_5__SCAN_IN), .A(n20355), .ZN(
        n16231) );
  OAI211_X1 U19594 ( .C1(n21038), .C2(n20269), .A(n16232), .B(n16231), .ZN(
        n16233) );
  AOI211_X1 U19595 ( .C1(n17717), .C2(n16235), .A(n16234), .B(n16233), .ZN(
        n16236) );
  OAI21_X1 U19596 ( .B1(n16237), .B2(n20273), .A(n16236), .ZN(n16238) );
  AOI21_X1 U19597 ( .B1(n17718), .B2(n20242), .A(n16238), .ZN(n16239) );
  OAI21_X1 U19598 ( .B1(n20276), .B2(n17079), .A(n16239), .ZN(P2_U2850) );
  XNOR2_X1 U19599 ( .A(n16240), .B(n9882), .ZN(n17096) );
  INV_X1 U19600 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n21036) );
  AOI21_X1 U19601 ( .B1(n20271), .B2(P2_EBX_REG_4__SCAN_IN), .A(n20355), .ZN(
        n16241) );
  OAI21_X1 U19602 ( .B1(n20269), .B2(n21036), .A(n16241), .ZN(n16242) );
  INV_X1 U19603 ( .A(n16242), .ZN(n16248) );
  NOR2_X1 U19604 ( .A1(n20233), .A2(n16243), .ZN(n16246) );
  INV_X1 U19605 ( .A(n20367), .ZN(n16245) );
  AOI21_X1 U19606 ( .B1(n16245), .B2(n16246), .A(n21006), .ZN(n16244) );
  OAI21_X1 U19607 ( .B1(n16246), .B2(n16245), .A(n16244), .ZN(n16247) );
  OAI211_X1 U19608 ( .C1(n20260), .C2(n10423), .A(n16248), .B(n16247), .ZN(
        n16249) );
  AOI21_X1 U19609 ( .B1(n9708), .B2(n16250), .A(n16249), .ZN(n16251) );
  OAI21_X1 U19610 ( .B1(n20362), .B2(n20277), .A(n16251), .ZN(n16252) );
  AOI21_X1 U19611 ( .B1(n20244), .B2(n17096), .A(n16252), .ZN(n16253) );
  OAI21_X1 U19612 ( .B1(n16508), .B2(n16305), .A(n16253), .ZN(P2_U2851) );
  NAND2_X1 U19613 ( .A1(n16255), .A2(n16254), .ZN(n16256) );
  INV_X1 U19614 ( .A(n20288), .ZN(n21089) );
  INV_X1 U19615 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n21035) );
  NAND2_X1 U19616 ( .A1(n20271), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n16257) );
  OAI21_X1 U19617 ( .B1(n20269), .B2(n21035), .A(n16257), .ZN(n16260) );
  INV_X1 U19618 ( .A(n16262), .ZN(n16258) );
  NOR3_X1 U19619 ( .A1(n16302), .A2(n16258), .A3(n17724), .ZN(n16259) );
  AOI211_X1 U19620 ( .C1(n20240), .C2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n16260), .B(n16259), .ZN(n16266) );
  OAI21_X1 U19621 ( .B1(n21006), .B2(n16262), .A(n16261), .ZN(n16264) );
  AOI22_X1 U19622 ( .A1(n16264), .A2(n17724), .B1(n9708), .B2(n10190), .ZN(
        n16265) );
  OAI211_X1 U19623 ( .C1(n21089), .C2(n20276), .A(n16266), .B(n16265), .ZN(
        n16267) );
  AOI21_X1 U19624 ( .B1(n17733), .B2(n20242), .A(n16267), .ZN(n16268) );
  OAI21_X1 U19625 ( .B1(n21090), .B2(n16305), .A(n16268), .ZN(P2_U2852) );
  INV_X1 U19626 ( .A(n16269), .ZN(n16270) );
  OAI21_X1 U19627 ( .B1(n10662), .B2(n16272), .A(n20227), .ZN(n16271) );
  AOI21_X1 U19628 ( .B1(n10662), .B2(n16272), .A(n16271), .ZN(n16277) );
  AOI22_X1 U19629 ( .A1(n20256), .A2(P2_REIP_REG_2__SCAN_IN), .B1(
        P2_EBX_REG_2__SCAN_IN), .B2(n20271), .ZN(n16274) );
  NAND2_X1 U19630 ( .A1(n20240), .A2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n16273) );
  OAI211_X1 U19631 ( .C1(n20273), .C2(n16275), .A(n16274), .B(n16273), .ZN(
        n16276) );
  AOI211_X1 U19632 ( .C1(n20244), .C2(n21104), .A(n16277), .B(n16276), .ZN(
        n16279) );
  NAND2_X1 U19633 ( .A1(n17146), .A2(n20242), .ZN(n16278) );
  OAI211_X1 U19634 ( .C1(n21100), .C2(n16305), .A(n16279), .B(n16278), .ZN(
        P2_U2853) );
  OR2_X1 U19635 ( .A1(n16281), .A2(n16280), .ZN(n16283) );
  NAND2_X1 U19636 ( .A1(n16283), .A2(n16282), .ZN(n20295) );
  NAND2_X1 U19637 ( .A1(n16294), .A2(n16284), .ZN(n16285) );
  NAND2_X1 U19638 ( .A1(n10662), .A2(n16285), .ZN(n17137) );
  NOR2_X1 U19639 ( .A1(n17137), .A2(n21006), .ZN(n16291) );
  AOI22_X1 U19640 ( .A1(n20240), .A2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B1(
        n16299), .B2(n16286), .ZN(n16288) );
  AOI22_X1 U19641 ( .A1(n20256), .A2(P2_REIP_REG_1__SCAN_IN), .B1(
        P2_EBX_REG_1__SCAN_IN), .B2(n20271), .ZN(n16287) );
  OAI211_X1 U19642 ( .C1(n16289), .C2(n20273), .A(n16288), .B(n16287), .ZN(
        n16290) );
  AOI211_X1 U19643 ( .C1(n20244), .C2(n20295), .A(n16291), .B(n16290), .ZN(
        n16293) );
  NAND2_X1 U19644 ( .A1(n13801), .A2(n20242), .ZN(n16292) );
  OAI211_X1 U19645 ( .C1(n21099), .C2(n16305), .A(n16293), .B(n16292), .ZN(
        P2_U2854) );
  INV_X1 U19646 ( .A(n16294), .ZN(n17129) );
  INV_X1 U19647 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n16295) );
  NOR2_X1 U19648 ( .A1(n20231), .A2(n16295), .ZN(n16297) );
  INV_X1 U19649 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n20211) );
  OAI22_X1 U19650 ( .A1(n20269), .A2(n20211), .B1(n20276), .B2(n20302), .ZN(
        n16296) );
  AOI211_X1 U19651 ( .C1(n9708), .C2(n16298), .A(n16297), .B(n16296), .ZN(
        n16301) );
  OAI21_X1 U19652 ( .B1(n20240), .B2(n16299), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n16300) );
  OAI211_X1 U19653 ( .C1(n17129), .C2(n16302), .A(n16301), .B(n16300), .ZN(
        n16303) );
  AOI21_X1 U19654 ( .B1(n13778), .B2(n20242), .A(n16303), .ZN(n16304) );
  OAI21_X1 U19655 ( .B1(n20673), .B2(n16305), .A(n16304), .ZN(P2_U2855) );
  MUX2_X1 U19656 ( .A(n16306), .B(P2_EBX_REG_31__SCAN_IN), .S(n16368), .Z(
        P2_U2856) );
  NAND2_X1 U19657 ( .A1(n16386), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n16308) );
  OAI211_X1 U19658 ( .C1(n16368), .C2(n16310), .A(n16309), .B(n16308), .ZN(
        P2_U2858) );
  NAND2_X1 U19659 ( .A1(n16312), .A2(n16311), .ZN(n16313) );
  XOR2_X1 U19660 ( .A(n16314), .B(n16313), .Z(n16410) );
  NAND2_X1 U19661 ( .A1(n16368), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n16316) );
  NAND2_X1 U19662 ( .A1(n16763), .A2(n16363), .ZN(n16315) );
  OAI211_X1 U19663 ( .C1(n16410), .C2(n16388), .A(n16316), .B(n16315), .ZN(
        P2_U2859) );
  OAI21_X1 U19664 ( .B1(n16317), .B2(n16319), .A(n16318), .ZN(n16417) );
  NAND2_X1 U19665 ( .A1(n16368), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n16321) );
  NAND2_X1 U19666 ( .A1(n16782), .A2(n16363), .ZN(n16320) );
  OAI211_X1 U19667 ( .C1(n16417), .C2(n16388), .A(n16321), .B(n16320), .ZN(
        P2_U2860) );
  NOR2_X1 U19668 ( .A1(n16323), .A2(n16333), .ZN(n16332) );
  NOR2_X1 U19669 ( .A1(n16332), .A2(n16324), .ZN(n16329) );
  NOR2_X1 U19670 ( .A1(n9736), .A2(n16325), .ZN(n16326) );
  XNOR2_X1 U19671 ( .A(n16327), .B(n16326), .ZN(n16328) );
  XNOR2_X1 U19672 ( .A(n16329), .B(n16328), .ZN(n16424) );
  NOR2_X1 U19673 ( .A1(n16794), .A2(n16386), .ZN(n16330) );
  AOI21_X1 U19674 ( .B1(P2_EBX_REG_26__SCAN_IN), .B2(n16386), .A(n16330), .ZN(
        n16331) );
  OAI21_X1 U19675 ( .B1(n16424), .B2(n16388), .A(n16331), .ZN(P2_U2861) );
  INV_X1 U19676 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n16336) );
  AOI21_X1 U19677 ( .B1(n16323), .B2(n16333), .A(n16332), .ZN(n16425) );
  NAND2_X1 U19678 ( .A1(n16425), .A2(n10619), .ZN(n16335) );
  NAND2_X1 U19679 ( .A1(n16799), .A2(n16363), .ZN(n16334) );
  OAI211_X1 U19680 ( .C1(n16363), .C2(n16336), .A(n16335), .B(n16334), .ZN(
        P2_U2862) );
  NAND2_X1 U19681 ( .A1(n16816), .A2(n16363), .ZN(n16341) );
  OR2_X1 U19682 ( .A1(n16339), .A2(n16338), .ZN(n16436) );
  NAND3_X1 U19683 ( .A1(n16337), .A2(n10619), .A3(n16436), .ZN(n16340) );
  OAI211_X1 U19684 ( .C1(n16363), .C2(n16342), .A(n16341), .B(n16340), .ZN(
        P2_U2863) );
  NAND2_X1 U19685 ( .A1(n9751), .A2(n16349), .ZN(n16348) );
  XNOR2_X1 U19686 ( .A(n16344), .B(n16343), .ZN(n16345) );
  XNOR2_X1 U19687 ( .A(n16348), .B(n16345), .ZN(n16445) );
  NOR2_X1 U19688 ( .A1(n16827), .A2(n16386), .ZN(n16346) );
  AOI21_X1 U19689 ( .B1(P2_EBX_REG_23__SCAN_IN), .B2(n16386), .A(n16346), .ZN(
        n16347) );
  OAI21_X1 U19690 ( .B1(n16445), .B2(n16388), .A(n16347), .ZN(P2_U2864) );
  OAI21_X1 U19691 ( .B1(n9751), .B2(n16349), .A(n16348), .ZN(n16452) );
  NAND2_X1 U19692 ( .A1(n16836), .A2(n16363), .ZN(n16351) );
  NAND2_X1 U19693 ( .A1(n16368), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n16350) );
  OAI211_X1 U19694 ( .C1(n16452), .C2(n16388), .A(n16351), .B(n16350), .ZN(
        P2_U2865) );
  AOI21_X1 U19695 ( .B1(n16353), .B2(n16352), .A(n9751), .ZN(n16453) );
  NAND2_X1 U19696 ( .A1(n16453), .A2(n10619), .ZN(n16355) );
  NAND2_X1 U19697 ( .A1(n16386), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n16354) );
  OAI211_X1 U19698 ( .C1(n16368), .C2(n16854), .A(n16355), .B(n16354), .ZN(
        P2_U2866) );
  OAI21_X1 U19699 ( .B1(n16357), .B2(n16358), .A(n16352), .ZN(n16465) );
  NAND2_X1 U19700 ( .A1(n16872), .A2(n16363), .ZN(n16360) );
  NAND2_X1 U19701 ( .A1(n16386), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n16359) );
  OAI211_X1 U19702 ( .C1(n16465), .C2(n16388), .A(n16360), .B(n16359), .ZN(
        P2_U2867) );
  INV_X1 U19703 ( .A(n16357), .ZN(n16361) );
  OAI21_X1 U19704 ( .B1(n9857), .B2(n16362), .A(n16361), .ZN(n16473) );
  NAND2_X1 U19705 ( .A1(n16368), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n16365) );
  NAND2_X1 U19706 ( .A1(n16880), .A2(n16363), .ZN(n16364) );
  OAI211_X1 U19707 ( .C1(n16473), .C2(n16388), .A(n16365), .B(n16364), .ZN(
        P2_U2868) );
  NOR2_X1 U19708 ( .A1(n9787), .A2(n16366), .ZN(n16367) );
  OR2_X1 U19709 ( .A1(n9857), .A2(n16367), .ZN(n16478) );
  MUX2_X1 U19710 ( .A(n16902), .B(n16369), .S(n16368), .Z(n16370) );
  OAI21_X1 U19711 ( .B1(n16388), .B2(n16478), .A(n16370), .ZN(P2_U2869) );
  AOI21_X1 U19712 ( .B1(n16372), .B2(n16371), .A(n9787), .ZN(n16484) );
  NAND2_X1 U19713 ( .A1(n16484), .A2(n10619), .ZN(n16374) );
  NAND2_X1 U19714 ( .A1(n16368), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n16373) );
  OAI211_X1 U19715 ( .C1(n16910), .C2(n16368), .A(n16374), .B(n16373), .ZN(
        P2_U2870) );
  INV_X1 U19716 ( .A(n16639), .ZN(n20225) );
  INV_X1 U19717 ( .A(n16371), .ZN(n16375) );
  AOI21_X1 U19718 ( .B1(n16376), .B2(n14366), .A(n16375), .ZN(n16489) );
  NAND2_X1 U19719 ( .A1(n16489), .A2(n10619), .ZN(n16378) );
  NAND2_X1 U19720 ( .A1(n16368), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n16377) );
  OAI211_X1 U19721 ( .C1(n20225), .C2(n16368), .A(n16378), .B(n16377), .ZN(
        P2_U2871) );
  INV_X1 U19722 ( .A(n16379), .ZN(n16383) );
  INV_X1 U19723 ( .A(n16380), .ZN(n16381) );
  OAI211_X1 U19724 ( .C1(n16383), .C2(n16382), .A(n16381), .B(n10619), .ZN(
        n16385) );
  NAND2_X1 U19725 ( .A1(n16368), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n16384) );
  OAI211_X1 U19726 ( .C1(n16969), .C2(n16386), .A(n16385), .B(n16384), .ZN(
        P2_U2875) );
  NOR2_X1 U19727 ( .A1(n17031), .A2(n16386), .ZN(n16392) );
  AOI211_X1 U19728 ( .C1(n16390), .C2(n16389), .A(n16388), .B(n16387), .ZN(
        n16391) );
  AOI211_X1 U19729 ( .C1(P2_EBX_REG_8__SCAN_IN), .C2(n16386), .A(n16392), .B(
        n16391), .ZN(n16393) );
  INV_X1 U19730 ( .A(n16393), .ZN(P2_U2879) );
  NAND2_X1 U19731 ( .A1(n16394), .A2(n20304), .ZN(n16396) );
  AOI22_X1 U19732 ( .A1(n16490), .A2(BUF2_REG_31__SCAN_IN), .B1(
        P2_EAX_REG_31__SCAN_IN), .B2(n20303), .ZN(n16395) );
  OAI211_X1 U19733 ( .C1(n17837), .C2(n16495), .A(n16396), .B(n16395), .ZN(
        P2_U2888) );
  INV_X1 U19734 ( .A(n16397), .ZN(n16404) );
  INV_X1 U19735 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n16401) );
  AOI22_X1 U19736 ( .A1(n16492), .A2(n16399), .B1(P2_EAX_REG_29__SCAN_IN), 
        .B2(n20303), .ZN(n16400) );
  OAI21_X1 U19737 ( .B1(n16495), .B2(n16401), .A(n16400), .ZN(n16402) );
  AOI21_X1 U19738 ( .B1(n16490), .B2(BUF2_REG_29__SCAN_IN), .A(n16402), .ZN(
        n16403) );
  AOI22_X1 U19739 ( .A1(n16492), .A2(n16405), .B1(P2_EAX_REG_28__SCAN_IN), 
        .B2(n20303), .ZN(n16406) );
  OAI21_X1 U19740 ( .B1(n16495), .B2(n17841), .A(n16406), .ZN(n16408) );
  NOR2_X1 U19741 ( .A1(n16770), .A2(n16487), .ZN(n16407) );
  OAI21_X1 U19742 ( .B1(n16410), .B2(n20298), .A(n16409), .ZN(P2_U2891) );
  INV_X1 U19743 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n16413) );
  AOI22_X1 U19744 ( .A1(n16492), .A2(n16411), .B1(P2_EAX_REG_27__SCAN_IN), 
        .B2(n20303), .ZN(n16412) );
  OAI21_X1 U19745 ( .B1(n16495), .B2(n16413), .A(n16412), .ZN(n16415) );
  NOR2_X1 U19746 ( .A1(n16779), .A2(n16487), .ZN(n16414) );
  AOI211_X1 U19747 ( .C1(n16490), .C2(BUF2_REG_27__SCAN_IN), .A(n16415), .B(
        n16414), .ZN(n16416) );
  OAI21_X1 U19748 ( .B1(n16417), .B2(n20298), .A(n16416), .ZN(P2_U2892) );
  INV_X1 U19749 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n16421) );
  NAND2_X1 U19750 ( .A1(n16490), .A2(BUF2_REG_26__SCAN_IN), .ZN(n16420) );
  AOI22_X1 U19751 ( .A1(n16492), .A2(n16418), .B1(P2_EAX_REG_26__SCAN_IN), 
        .B2(n20303), .ZN(n16419) );
  OAI211_X1 U19752 ( .C1(n16495), .C2(n16421), .A(n16420), .B(n16419), .ZN(
        n16422) );
  AOI21_X1 U19753 ( .B1(n16797), .B2(n20304), .A(n16422), .ZN(n16423) );
  OAI21_X1 U19754 ( .B1(n16424), .B2(n20298), .A(n16423), .ZN(P2_U2893) );
  INV_X1 U19755 ( .A(n20298), .ZN(n20306) );
  NAND2_X1 U19756 ( .A1(n16425), .A2(n20306), .ZN(n16431) );
  INV_X1 U19757 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n16428) );
  AOI22_X1 U19758 ( .A1(n16492), .A2(n16426), .B1(P2_EAX_REG_25__SCAN_IN), 
        .B2(n20303), .ZN(n16427) );
  OAI21_X1 U19759 ( .B1(n16495), .B2(n16428), .A(n16427), .ZN(n16429) );
  AOI21_X1 U19760 ( .B1(n16490), .B2(BUF2_REG_25__SCAN_IN), .A(n16429), .ZN(
        n16430) );
  OAI211_X1 U19761 ( .C1(n16806), .C2(n16487), .A(n16431), .B(n16430), .ZN(
        P2_U2894) );
  AOI22_X1 U19762 ( .A1(n16492), .A2(n16432), .B1(P2_EAX_REG_24__SCAN_IN), 
        .B2(n20303), .ZN(n16433) );
  OAI21_X1 U19763 ( .B1(n16495), .B2(n17846), .A(n16433), .ZN(n16435) );
  NOR2_X1 U19764 ( .A1(n16818), .A2(n16487), .ZN(n16434) );
  AOI211_X1 U19765 ( .C1(n16490), .C2(BUF2_REG_24__SCAN_IN), .A(n16435), .B(
        n16434), .ZN(n16438) );
  NAND3_X1 U19766 ( .A1(n16337), .A2(n20306), .A3(n16436), .ZN(n16437) );
  NAND2_X1 U19767 ( .A1(n16438), .A2(n16437), .ZN(P2_U2895) );
  INV_X1 U19768 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n16442) );
  NAND2_X1 U19769 ( .A1(n16490), .A2(BUF2_REG_23__SCAN_IN), .ZN(n16441) );
  AOI22_X1 U19770 ( .A1(n16492), .A2(n16439), .B1(P2_EAX_REG_23__SCAN_IN), 
        .B2(n20303), .ZN(n16440) );
  OAI211_X1 U19771 ( .C1(n16442), .C2(n16495), .A(n16441), .B(n16440), .ZN(
        n16443) );
  AOI21_X1 U19772 ( .B1(n16830), .B2(n20304), .A(n16443), .ZN(n16444) );
  OAI21_X1 U19773 ( .B1(n16445), .B2(n20298), .A(n16444), .ZN(P2_U2896) );
  INV_X1 U19774 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n16449) );
  NAND2_X1 U19775 ( .A1(n16490), .A2(BUF2_REG_22__SCAN_IN), .ZN(n16448) );
  AOI22_X1 U19776 ( .A1(n16492), .A2(n16446), .B1(P2_EAX_REG_22__SCAN_IN), 
        .B2(n20303), .ZN(n16447) );
  OAI211_X1 U19777 ( .C1(n16449), .C2(n16495), .A(n16448), .B(n16447), .ZN(
        n16450) );
  AOI21_X1 U19778 ( .B1(n16844), .B2(n20304), .A(n16450), .ZN(n16451) );
  OAI21_X1 U19779 ( .B1(n20298), .B2(n16452), .A(n16451), .ZN(P2_U2897) );
  INV_X1 U19780 ( .A(n16453), .ZN(n16459) );
  INV_X1 U19781 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n16456) );
  NAND2_X1 U19782 ( .A1(n16490), .A2(BUF2_REG_21__SCAN_IN), .ZN(n16455) );
  AOI22_X1 U19783 ( .A1(n16492), .A2(n20423), .B1(P2_EAX_REG_21__SCAN_IN), 
        .B2(n20303), .ZN(n16454) );
  OAI211_X1 U19784 ( .C1(n16456), .C2(n16495), .A(n16455), .B(n16454), .ZN(
        n16457) );
  AOI21_X1 U19785 ( .B1(n16857), .B2(n20304), .A(n16457), .ZN(n16458) );
  OAI21_X1 U19786 ( .B1(n16459), .B2(n20298), .A(n16458), .ZN(P2_U2898) );
  INV_X1 U19787 ( .A(n16874), .ZN(n16463) );
  NAND2_X1 U19788 ( .A1(n16490), .A2(BUF2_REG_20__SCAN_IN), .ZN(n16461) );
  AOI22_X1 U19789 ( .A1(n16492), .A2(n16510), .B1(P2_EAX_REG_20__SCAN_IN), 
        .B2(n20303), .ZN(n16460) );
  OAI211_X1 U19790 ( .C1(n17851), .C2(n16495), .A(n16461), .B(n16460), .ZN(
        n16462) );
  AOI21_X1 U19791 ( .B1(n16463), .B2(n20304), .A(n16462), .ZN(n16464) );
  OAI21_X1 U19792 ( .B1(n20298), .B2(n16465), .A(n16464), .ZN(P2_U2899) );
  INV_X1 U19793 ( .A(n16887), .ZN(n16471) );
  INV_X1 U19794 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n16469) );
  NAND2_X1 U19795 ( .A1(n16490), .A2(BUF2_REG_19__SCAN_IN), .ZN(n16468) );
  AOI22_X1 U19796 ( .A1(n16492), .A2(n16466), .B1(P2_EAX_REG_19__SCAN_IN), 
        .B2(n20303), .ZN(n16467) );
  OAI211_X1 U19797 ( .C1(n16469), .C2(n16495), .A(n16468), .B(n16467), .ZN(
        n16470) );
  AOI21_X1 U19798 ( .B1(n16471), .B2(n20304), .A(n16470), .ZN(n16472) );
  OAI21_X1 U19799 ( .B1(n20298), .B2(n16473), .A(n16472), .ZN(P2_U2900) );
  NAND2_X1 U19800 ( .A1(n16490), .A2(BUF2_REG_18__SCAN_IN), .ZN(n16475) );
  AOI22_X1 U19801 ( .A1(n16492), .A2(n16518), .B1(P2_EAX_REG_18__SCAN_IN), 
        .B2(n20303), .ZN(n16474) );
  OAI211_X1 U19802 ( .C1(n17854), .C2(n16495), .A(n16475), .B(n16474), .ZN(
        n16476) );
  AOI21_X1 U19803 ( .B1(n16899), .B2(n20304), .A(n16476), .ZN(n16477) );
  OAI21_X1 U19804 ( .B1(n20298), .B2(n16478), .A(n16477), .ZN(P2_U2901) );
  INV_X1 U19805 ( .A(n16917), .ZN(n16488) );
  NOR2_X1 U19806 ( .A1(n16495), .A2(n16479), .ZN(n16483) );
  OAI22_X1 U19807 ( .A1(n16481), .A2(n20393), .B1(n16519), .B2(n16480), .ZN(
        n16482) );
  AOI211_X1 U19808 ( .C1(n16490), .C2(BUF2_REG_17__SCAN_IN), .A(n16483), .B(
        n16482), .ZN(n16486) );
  NAND2_X1 U19809 ( .A1(n16484), .A2(n20306), .ZN(n16485) );
  OAI211_X1 U19810 ( .C1(n16488), .C2(n16487), .A(n16486), .B(n16485), .ZN(
        P2_U2902) );
  INV_X1 U19811 ( .A(n16489), .ZN(n16499) );
  INV_X1 U19812 ( .A(n20224), .ZN(n16497) );
  NAND2_X1 U19813 ( .A1(n16490), .A2(BUF2_REG_16__SCAN_IN), .ZN(n16494) );
  AOI22_X1 U19814 ( .A1(n16492), .A2(n16491), .B1(n20303), .B2(
        P2_EAX_REG_16__SCAN_IN), .ZN(n16493) );
  OAI211_X1 U19815 ( .C1(n17857), .C2(n16495), .A(n16494), .B(n16493), .ZN(
        n16496) );
  AOI21_X1 U19816 ( .B1(n16497), .B2(n20304), .A(n16496), .ZN(n16498) );
  OAI21_X1 U19817 ( .B1(n16499), .B2(n20298), .A(n16498), .ZN(P2_U2903) );
  INV_X1 U19818 ( .A(n21104), .ZN(n16503) );
  XNOR2_X1 U19819 ( .A(n20373), .B(n21104), .ZN(n16517) );
  OR2_X1 U19820 ( .A1(n20672), .A2(n20295), .ZN(n16501) );
  NAND2_X1 U19821 ( .A1(n20672), .A2(n20295), .ZN(n16500) );
  NAND2_X1 U19822 ( .A1(n16501), .A2(n16500), .ZN(n20297) );
  NOR2_X1 U19823 ( .A1(n20673), .A2(n20302), .ZN(n20305) );
  NOR2_X1 U19824 ( .A1(n20297), .A2(n20305), .ZN(n20296) );
  INV_X1 U19825 ( .A(n16501), .ZN(n16502) );
  NOR2_X1 U19826 ( .A1(n20296), .A2(n16502), .ZN(n16516) );
  NOR2_X1 U19827 ( .A1(n16517), .A2(n16516), .ZN(n16515) );
  AOI21_X1 U19828 ( .B1(n16503), .B2(n21100), .A(n16515), .ZN(n20291) );
  XNOR2_X1 U19829 ( .A(n20671), .B(n20288), .ZN(n20290) );
  NOR2_X1 U19830 ( .A1(n20291), .A2(n20290), .ZN(n20289) );
  AOI21_X1 U19831 ( .B1(n21090), .B2(n21089), .A(n20289), .ZN(n16504) );
  NOR2_X1 U19832 ( .A1(n16504), .A2(n17096), .ZN(n16509) );
  OR3_X1 U19833 ( .A1(n16509), .A2(n16508), .A3(n20298), .ZN(n16507) );
  AOI22_X1 U19834 ( .A1(n16505), .A2(n20423), .B1(n20303), .B2(
        P2_EAX_REG_5__SCAN_IN), .ZN(n16506) );
  OAI211_X1 U19835 ( .C1(n20283), .C2(n17079), .A(n16507), .B(n16506), .ZN(
        P2_U2914) );
  XNOR2_X1 U19836 ( .A(n16509), .B(n16508), .ZN(n16514) );
  INV_X1 U19837 ( .A(n16510), .ZN(n20416) );
  INV_X1 U19838 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n16511) );
  OAI22_X1 U19839 ( .A1(n20311), .A2(n20416), .B1(n16519), .B2(n16511), .ZN(
        n16512) );
  AOI21_X1 U19840 ( .B1(n20304), .B2(n17096), .A(n16512), .ZN(n16513) );
  OAI21_X1 U19841 ( .B1(n16514), .B2(n20298), .A(n16513), .ZN(P2_U2915) );
  AOI21_X1 U19842 ( .B1(n16517), .B2(n16516), .A(n16515), .ZN(n16522) );
  INV_X1 U19843 ( .A(n16518), .ZN(n20401) );
  INV_X1 U19844 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n20339) );
  OAI22_X1 U19845 ( .A1(n20311), .A2(n20401), .B1(n16519), .B2(n20339), .ZN(
        n16520) );
  AOI21_X1 U19846 ( .B1(n20304), .B2(n21104), .A(n16520), .ZN(n16521) );
  OAI21_X1 U19847 ( .B1(n16522), .B2(n20298), .A(n16521), .ZN(P2_U2917) );
  XNOR2_X1 U19848 ( .A(n16525), .B(n22042), .ZN(n16526) );
  XNOR2_X1 U19849 ( .A(n16527), .B(n16526), .ZN(n16774) );
  NAND2_X1 U19850 ( .A1(n16763), .A2(n20370), .ZN(n16530) );
  NOR2_X1 U19851 ( .A1(n16730), .A2(n16528), .ZN(n16766) );
  AOI21_X1 U19852 ( .B1(n20356), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n16766), .ZN(n16529) );
  OAI211_X1 U19853 ( .C1(n20368), .C2(n16531), .A(n16530), .B(n16529), .ZN(
        n16532) );
  AOI21_X1 U19854 ( .B1(n20357), .B2(n16772), .A(n16532), .ZN(n16533) );
  OAI21_X1 U19855 ( .B1(n16774), .B2(n16737), .A(n16533), .ZN(P2_U2986) );
  XNOR2_X1 U19856 ( .A(n16534), .B(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16787) );
  NOR2_X1 U19857 ( .A1(n20368), .A2(n16535), .ZN(n16538) );
  OR2_X1 U19858 ( .A1(n16730), .A2(n21074), .ZN(n16775) );
  OAI21_X1 U19859 ( .B1(n17736), .B2(n16536), .A(n16775), .ZN(n16537) );
  AOI211_X1 U19860 ( .C1(n16782), .C2(n20370), .A(n16538), .B(n16537), .ZN(
        n16540) );
  NAND2_X1 U19861 ( .A1(n10066), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n16544) );
  NAND2_X1 U19862 ( .A1(n16544), .A2(n16777), .ZN(n16783) );
  NAND3_X1 U19863 ( .A1(n16784), .A2(n20357), .A3(n16783), .ZN(n16539) );
  OAI211_X1 U19864 ( .C1(n16787), .C2(n16737), .A(n16540), .B(n16539), .ZN(
        P2_U2987) );
  INV_X1 U19865 ( .A(n16794), .ZN(n16545) );
  NAND2_X1 U19866 ( .A1(n16545), .A2(n20370), .ZN(n16547) );
  INV_X1 U19867 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n21072) );
  NOR2_X1 U19868 ( .A1(n20217), .A2(n21072), .ZN(n16792) );
  AOI21_X1 U19869 ( .B1(n20356), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n16792), .ZN(n16546) );
  OAI211_X1 U19870 ( .C1(n20368), .C2(n16548), .A(n16547), .B(n16546), .ZN(
        n16549) );
  NOR2_X1 U19871 ( .A1(n16551), .A2(n11442), .ZN(n16552) );
  XNOR2_X1 U19872 ( .A(n16541), .B(n16552), .ZN(n16810) );
  OAI21_X1 U19873 ( .B1(n16553), .B2(n16813), .A(n16554), .ZN(n16555) );
  AND2_X1 U19874 ( .A1(n16556), .A2(n16555), .ZN(n16808) );
  NAND2_X1 U19875 ( .A1(n16799), .A2(n20370), .ZN(n16558) );
  INV_X1 U19876 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n21070) );
  NOR2_X1 U19877 ( .A1(n16730), .A2(n21070), .ZN(n16802) );
  AOI21_X1 U19878 ( .B1(n20356), .B2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n16802), .ZN(n16557) );
  OAI211_X1 U19879 ( .C1(n11778), .C2(n20368), .A(n16558), .B(n16557), .ZN(
        n16559) );
  AOI21_X1 U19880 ( .B1(n20357), .B2(n16808), .A(n16559), .ZN(n16560) );
  OAI21_X1 U19881 ( .B1(n16810), .B2(n16737), .A(n16560), .ZN(P2_U2989) );
  XNOR2_X1 U19882 ( .A(n16553), .B(n16813), .ZN(n16822) );
  XNOR2_X1 U19883 ( .A(n16561), .B(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n16562) );
  XNOR2_X1 U19884 ( .A(n16563), .B(n16562), .ZN(n16820) );
  NAND2_X1 U19885 ( .A1(n16820), .A2(n11457), .ZN(n16568) );
  NAND2_X1 U19886 ( .A1(n20355), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n16811) );
  NAND2_X1 U19887 ( .A1(n20356), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n16564) );
  OAI211_X1 U19888 ( .C1(n20368), .C2(n16565), .A(n16811), .B(n16564), .ZN(
        n16566) );
  AOI21_X1 U19889 ( .B1(n16816), .B2(n20370), .A(n16566), .ZN(n16567) );
  OAI211_X1 U19890 ( .C1(n16822), .C2(n16762), .A(n16568), .B(n16567), .ZN(
        P2_U2990) );
  OAI21_X1 U19891 ( .B1(n16580), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n16553), .ZN(n16834) );
  XOR2_X1 U19892 ( .A(n16570), .B(n16569), .Z(n16831) );
  NOR2_X1 U19893 ( .A1(n16827), .A2(n20363), .ZN(n16574) );
  NAND2_X1 U19894 ( .A1(n20355), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n16826) );
  NAND2_X1 U19895 ( .A1(n20356), .A2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n16571) );
  OAI211_X1 U19896 ( .C1(n20368), .C2(n16572), .A(n16826), .B(n16571), .ZN(
        n16573) );
  AOI211_X1 U19897 ( .C1(n16831), .C2(n11457), .A(n16574), .B(n16573), .ZN(
        n16575) );
  OAI21_X1 U19898 ( .B1(n16834), .B2(n16762), .A(n16575), .ZN(P2_U2991) );
  INV_X1 U19899 ( .A(n16576), .ZN(n16578) );
  NAND2_X1 U19900 ( .A1(n16578), .A2(n16577), .ZN(n16579) );
  XNOR2_X1 U19901 ( .A(n9801), .B(n16579), .ZN(n16847) );
  NOR2_X1 U19902 ( .A1(n16730), .A2(n16581), .ZN(n16837) );
  AOI21_X1 U19903 ( .B1(n20356), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n16837), .ZN(n16582) );
  OAI21_X1 U19904 ( .B1(n20368), .B2(n16583), .A(n16582), .ZN(n16584) );
  AOI21_X1 U19905 ( .B1(n16836), .B2(n20370), .A(n16584), .ZN(n16585) );
  OAI211_X1 U19906 ( .C1(n16847), .C2(n16737), .A(n16586), .B(n16585), .ZN(
        P2_U2992) );
  INV_X1 U19907 ( .A(n16600), .ZN(n16589) );
  AOI21_X1 U19908 ( .B1(n16603), .B2(n16589), .A(n16601), .ZN(n16593) );
  NAND2_X1 U19909 ( .A1(n16591), .A2(n16590), .ZN(n16592) );
  XNOR2_X1 U19910 ( .A(n16593), .B(n16592), .ZN(n16859) );
  INV_X1 U19911 ( .A(n16854), .ZN(n16598) );
  INV_X1 U19912 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n21064) );
  NOR2_X1 U19913 ( .A1(n16730), .A2(n21064), .ZN(n16850) );
  AOI21_X1 U19914 ( .B1(n20356), .B2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n16850), .ZN(n16594) );
  OAI21_X1 U19915 ( .B1(n20368), .B2(n16595), .A(n16594), .ZN(n16597) );
  OAI21_X1 U19916 ( .B1(n16859), .B2(n16737), .A(n16599), .ZN(P2_U2993) );
  NOR2_X1 U19917 ( .A1(n16601), .A2(n16600), .ZN(n16602) );
  NAND2_X1 U19918 ( .A1(n16872), .A2(n20370), .ZN(n16608) );
  NOR2_X1 U19919 ( .A1(n16730), .A2(n16606), .ZN(n16867) );
  AOI21_X1 U19920 ( .B1(n20356), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n16867), .ZN(n16607) );
  OAI211_X1 U19921 ( .C1(n16609), .C2(n20368), .A(n16608), .B(n16607), .ZN(
        n16610) );
  AOI21_X1 U19922 ( .B1(n16876), .B2(n20357), .A(n16610), .ZN(n16611) );
  NAND2_X1 U19923 ( .A1(n16612), .A2(n16615), .ZN(n16613) );
  AOI22_X1 U19924 ( .A1(n16616), .A2(n16615), .B1(n16614), .B2(n16613), .ZN(
        n16906) );
  NOR2_X1 U19925 ( .A1(n16730), .A2(n16618), .ZN(n16894) );
  NOR2_X1 U19926 ( .A1(n20368), .A2(n16619), .ZN(n16620) );
  AOI211_X1 U19927 ( .C1(n20356), .C2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n16894), .B(n16620), .ZN(n16621) );
  OAI21_X1 U19928 ( .B1(n16902), .B2(n20363), .A(n16621), .ZN(n16622) );
  OAI21_X1 U19929 ( .B1(n16906), .B2(n16737), .A(n16623), .ZN(P2_U2996) );
  NAND2_X1 U19930 ( .A1(n16625), .A2(n16624), .ZN(n16626) );
  XNOR2_X1 U19931 ( .A(n9838), .B(n16626), .ZN(n16920) );
  OAI211_X1 U19932 ( .C1(n16911), .C2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n20357), .B(n16627), .ZN(n16633) );
  INV_X1 U19933 ( .A(n16910), .ZN(n16631) );
  NAND2_X1 U19934 ( .A1(n20355), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n16909) );
  NAND2_X1 U19935 ( .A1(n20356), .A2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n16628) );
  OAI211_X1 U19936 ( .C1(n20368), .C2(n16629), .A(n16909), .B(n16628), .ZN(
        n16630) );
  AOI21_X1 U19937 ( .B1(n16631), .B2(n20370), .A(n16630), .ZN(n16632) );
  OAI211_X1 U19938 ( .C1(n16920), .C2(n16737), .A(n16633), .B(n16632), .ZN(
        P2_U2997) );
  INV_X1 U19939 ( .A(n16643), .ZN(n16635) );
  INV_X1 U19940 ( .A(n16911), .ZN(n16634) );
  OAI211_X1 U19941 ( .C1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n16635), .A(
        n16634), .B(n20357), .ZN(n16641) );
  AOI21_X1 U19942 ( .B1(n20356), .B2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n16636), .ZN(n16637) );
  OAI21_X1 U19943 ( .B1(n20368), .B2(n20223), .A(n16637), .ZN(n16638) );
  AOI21_X1 U19944 ( .B1(n16639), .B2(n20370), .A(n16638), .ZN(n16640) );
  OAI211_X1 U19945 ( .C1(n16642), .C2(n16737), .A(n16641), .B(n16640), .ZN(
        P2_U2998) );
  OAI21_X1 U19946 ( .B1(n16653), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n16643), .ZN(n16935) );
  NOR2_X1 U19947 ( .A1(n16730), .A2(n21055), .ZN(n16923) );
  AOI21_X1 U19948 ( .B1(n20356), .B2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n16923), .ZN(n16644) );
  OAI21_X1 U19949 ( .B1(n20368), .B2(n16645), .A(n16644), .ZN(n16651) );
  NAND2_X1 U19950 ( .A1(n16647), .A2(n16646), .ZN(n16648) );
  XNOR2_X1 U19951 ( .A(n16649), .B(n16648), .ZN(n16930) );
  NOR2_X1 U19952 ( .A1(n16930), .A2(n16737), .ZN(n16650) );
  AOI211_X1 U19953 ( .C1(n20370), .C2(n16922), .A(n16651), .B(n16650), .ZN(
        n16652) );
  OAI21_X1 U19954 ( .B1(n16762), .B2(n16935), .A(n16652), .ZN(P2_U2999) );
  OAI21_X1 U19955 ( .B1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n16666), .A(
        n10004), .ZN(n16949) );
  NAND2_X1 U19956 ( .A1(n16655), .A2(n16654), .ZN(n16656) );
  XNOR2_X1 U19957 ( .A(n16657), .B(n16656), .ZN(n16946) );
  INV_X1 U19958 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n21053) );
  NOR2_X1 U19959 ( .A1(n16730), .A2(n21053), .ZN(n16939) );
  NOR2_X1 U19960 ( .A1(n20368), .A2(n20234), .ZN(n16658) );
  AOI211_X1 U19961 ( .C1(n20356), .C2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n16939), .B(n16658), .ZN(n16659) );
  OAI21_X1 U19962 ( .B1(n20241), .B2(n20363), .A(n16659), .ZN(n16660) );
  AOI21_X1 U19963 ( .B1(n16946), .B2(n11457), .A(n16660), .ZN(n16661) );
  OAI21_X1 U19964 ( .B1(n16949), .B2(n16762), .A(n16661), .ZN(P2_U3000) );
  NAND2_X1 U19965 ( .A1(n16663), .A2(n16662), .ZN(n16664) );
  XNOR2_X1 U19966 ( .A(n16665), .B(n16664), .ZN(n16963) );
  AOI21_X1 U19967 ( .B1(n16667), .B2(n16674), .A(n16666), .ZN(n16950) );
  NAND2_X1 U19968 ( .A1(n16950), .A2(n20357), .ZN(n16672) );
  NAND2_X1 U19969 ( .A1(n20355), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n16953) );
  NAND2_X1 U19970 ( .A1(n20356), .A2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n16668) );
  OAI211_X1 U19971 ( .C1(n20368), .C2(n16669), .A(n16953), .B(n16668), .ZN(
        n16670) );
  AOI21_X1 U19972 ( .B1(n16960), .B2(n20370), .A(n16670), .ZN(n16671) );
  OAI21_X1 U19973 ( .B1(n16673), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n16674), .ZN(n16974) );
  NAND2_X1 U19974 ( .A1(n16676), .A2(n16675), .ZN(n16677) );
  XNOR2_X1 U19975 ( .A(n16678), .B(n16677), .ZN(n16972) );
  NOR2_X1 U19976 ( .A1(n16730), .A2(n21050), .ZN(n16965) );
  NOR2_X1 U19977 ( .A1(n20368), .A2(n16679), .ZN(n16680) );
  AOI211_X1 U19978 ( .C1(n20356), .C2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n16965), .B(n16680), .ZN(n16681) );
  OAI21_X1 U19979 ( .B1(n16969), .B2(n20363), .A(n16681), .ZN(n16682) );
  AOI21_X1 U19980 ( .B1(n16972), .B2(n11457), .A(n16682), .ZN(n16683) );
  OAI21_X1 U19981 ( .B1(n16974), .B2(n16762), .A(n16683), .ZN(P2_U3002) );
  NOR2_X1 U19982 ( .A1(n16712), .A2(n16992), .ZN(n16709) );
  INV_X1 U19983 ( .A(n16673), .ZN(n16684) );
  OAI21_X1 U19984 ( .B1(n16709), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n16684), .ZN(n16986) );
  INV_X1 U19985 ( .A(n16756), .ZN(n16686) );
  INV_X1 U19986 ( .A(n16742), .ZN(n16687) );
  OAI21_X1 U19987 ( .B1(n16744), .B2(n16687), .A(n16741), .ZN(n16725) );
  INV_X1 U19988 ( .A(n16722), .ZN(n16688) );
  INV_X1 U19989 ( .A(n16701), .ZN(n16690) );
  NAND2_X1 U19990 ( .A1(n16692), .A2(n16691), .ZN(n16693) );
  NOR2_X1 U19991 ( .A1(n20217), .A2(n16694), .ZN(n16977) );
  NOR2_X1 U19992 ( .A1(n17736), .A2(n16695), .ZN(n16696) );
  AOI211_X1 U19993 ( .C1(n16697), .C2(n17725), .A(n16977), .B(n16696), .ZN(
        n16698) );
  OAI21_X1 U19994 ( .B1(n16982), .B2(n20363), .A(n16698), .ZN(n16699) );
  AOI21_X1 U19995 ( .B1(n16984), .B2(n11457), .A(n16699), .ZN(n16700) );
  OAI21_X1 U19996 ( .B1(n16986), .B2(n16762), .A(n16700), .ZN(P2_U3003) );
  NAND2_X1 U19997 ( .A1(n16702), .A2(n16701), .ZN(n16705) );
  NAND2_X1 U19998 ( .A1(n16703), .A2(n16715), .ZN(n16704) );
  XOR2_X1 U19999 ( .A(n16705), .B(n16704), .Z(n17000) );
  NOR2_X1 U20000 ( .A1(n20217), .A2(n22182), .ZN(n16988) );
  AOI21_X1 U20001 ( .B1(n20356), .B2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n16988), .ZN(n16706) );
  OAI21_X1 U20002 ( .B1(n20368), .B2(n16707), .A(n16706), .ZN(n16708) );
  AOI21_X1 U20003 ( .B1(n16987), .B2(n20370), .A(n16708), .ZN(n16711) );
  INV_X1 U20004 ( .A(n16709), .ZN(n16997) );
  NAND2_X1 U20005 ( .A1(n16712), .A2(n16992), .ZN(n16996) );
  NAND3_X1 U20006 ( .A1(n16997), .A2(n20357), .A3(n16996), .ZN(n16710) );
  OAI211_X1 U20007 ( .C1(n17000), .C2(n16737), .A(n16711), .B(n16710), .ZN(
        P2_U3004) );
  OAI21_X1 U20008 ( .B1(n16713), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n16712), .ZN(n17014) );
  NAND2_X1 U20009 ( .A1(n16715), .A2(n16714), .ZN(n16716) );
  XNOR2_X1 U20010 ( .A(n16717), .B(n16716), .ZN(n17011) );
  INV_X1 U20011 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n21046) );
  NOR2_X1 U20012 ( .A1(n20217), .A2(n21046), .ZN(n17002) );
  NOR2_X1 U20013 ( .A1(n17736), .A2(n20259), .ZN(n16718) );
  AOI211_X1 U20014 ( .C1(n20251), .C2(n17725), .A(n17002), .B(n16718), .ZN(
        n16719) );
  OAI21_X1 U20015 ( .B1(n20261), .B2(n20363), .A(n16719), .ZN(n16720) );
  AOI21_X1 U20016 ( .B1(n17011), .B2(n11457), .A(n16720), .ZN(n16721) );
  OAI21_X1 U20017 ( .B1(n17014), .B2(n16762), .A(n16721), .ZN(P2_U3005) );
  NAND2_X1 U20018 ( .A1(n16723), .A2(n16722), .ZN(n16724) );
  XNOR2_X1 U20019 ( .A(n16725), .B(n16724), .ZN(n17035) );
  NAND2_X1 U20020 ( .A1(n16728), .A2(n16729), .ZN(n17015) );
  NAND3_X1 U20021 ( .A1(n16727), .A2(n17015), .A3(n20357), .ZN(n16736) );
  NOR2_X1 U20022 ( .A1(n16730), .A2(n21044), .ZN(n17028) );
  AOI21_X1 U20023 ( .B1(n20356), .B2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n17028), .ZN(n16731) );
  OAI21_X1 U20024 ( .B1(n20368), .B2(n16732), .A(n16731), .ZN(n16733) );
  AOI21_X1 U20025 ( .B1(n16734), .B2(n20370), .A(n16733), .ZN(n16735) );
  OAI211_X1 U20026 ( .C1(n17035), .C2(n16737), .A(n16736), .B(n16735), .ZN(
        P2_U3006) );
  XNOR2_X1 U20027 ( .A(n16739), .B(n22145), .ZN(n16740) );
  XNOR2_X1 U20028 ( .A(n16738), .B(n16740), .ZN(n17046) );
  NAND2_X1 U20029 ( .A1(n16742), .A2(n16741), .ZN(n16743) );
  XNOR2_X1 U20030 ( .A(n16744), .B(n16743), .ZN(n17044) );
  NOR2_X1 U20031 ( .A1(n20217), .A2(n21042), .ZN(n17036) );
  AOI21_X1 U20032 ( .B1(n20356), .B2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n17036), .ZN(n16746) );
  NAND2_X1 U20033 ( .A1(n17725), .A2(n20267), .ZN(n16745) );
  OAI211_X1 U20034 ( .C1(n20278), .C2(n20363), .A(n16746), .B(n16745), .ZN(
        n16747) );
  AOI21_X1 U20035 ( .B1(n17044), .B2(n11457), .A(n16747), .ZN(n16748) );
  OAI21_X1 U20036 ( .B1(n17046), .B2(n16762), .A(n16748), .ZN(P2_U3007) );
  MUX2_X1 U20037 ( .A(n16753), .B(n16751), .S(n16752), .Z(n16754) );
  XNOR2_X1 U20038 ( .A(n16755), .B(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17058) );
  NOR2_X1 U20039 ( .A1(n20217), .A2(n21040), .ZN(n17049) );
  NOR2_X1 U20040 ( .A1(n20368), .A2(n16757), .ZN(n16758) );
  AOI211_X1 U20041 ( .C1(n20356), .C2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n17049), .B(n16758), .ZN(n16759) );
  OAI21_X1 U20042 ( .B1(n17054), .B2(n20363), .A(n16759), .ZN(n16760) );
  AOI21_X1 U20043 ( .B1(n17056), .B2(n11457), .A(n16760), .ZN(n16761) );
  OAI21_X1 U20044 ( .B1(n17058), .B2(n16762), .A(n16761), .ZN(P2_U3008) );
  NAND2_X1 U20045 ( .A1(n16763), .A2(n17076), .ZN(n16769) );
  NOR3_X1 U20046 ( .A1(n16764), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        n16777), .ZN(n16765) );
  AOI211_X1 U20047 ( .C1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n16767), .A(
        n16766), .B(n16765), .ZN(n16768) );
  OAI211_X1 U20048 ( .C1(n16770), .C2(n17105), .A(n16769), .B(n16768), .ZN(
        n16771) );
  AOI21_X1 U20049 ( .B1(n17738), .B2(n16772), .A(n16771), .ZN(n16773) );
  OAI21_X1 U20050 ( .B1(n16774), .B2(n17101), .A(n16773), .ZN(P2_U3018) );
  OAI211_X1 U20051 ( .C1(n16778), .C2(n16777), .A(n16776), .B(n16775), .ZN(
        n16781) );
  NOR2_X1 U20052 ( .A1(n16779), .A2(n17105), .ZN(n16780) );
  AOI211_X1 U20053 ( .C1(n16782), .C2(n17076), .A(n16781), .B(n16780), .ZN(
        n16786) );
  NAND3_X1 U20054 ( .A1(n16784), .A2(n17738), .A3(n16783), .ZN(n16785) );
  OAI211_X1 U20055 ( .C1(n16787), .C2(n17101), .A(n16786), .B(n16785), .ZN(
        P2_U3019) );
  NAND2_X1 U20056 ( .A1(n16789), .A2(n16813), .ZN(n16812) );
  NAND2_X1 U20057 ( .A1(n16814), .A2(n16812), .ZN(n16803) );
  NOR2_X1 U20058 ( .A1(n11149), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n16790) );
  INV_X1 U20059 ( .A(n16789), .ZN(n16800) );
  AOI211_X1 U20060 ( .C1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(n16790), .B(n16800), .ZN(
        n16791) );
  AOI211_X1 U20061 ( .C1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .C2(n16803), .A(
        n16792), .B(n16791), .ZN(n16793) );
  OAI21_X1 U20062 ( .B1(n16794), .B2(n17745), .A(n16793), .ZN(n16796) );
  NAND2_X1 U20063 ( .A1(n16799), .A2(n17076), .ZN(n16805) );
  NOR3_X1 U20064 ( .A1(n16800), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        n16813), .ZN(n16801) );
  AOI211_X1 U20065 ( .C1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .C2(n16803), .A(
        n16802), .B(n16801), .ZN(n16804) );
  OAI211_X1 U20066 ( .C1(n16806), .C2(n17105), .A(n16805), .B(n16804), .ZN(
        n16807) );
  AOI21_X1 U20067 ( .B1(n17738), .B2(n16808), .A(n16807), .ZN(n16809) );
  OAI21_X1 U20068 ( .B1(n16810), .B2(n17101), .A(n16809), .ZN(P2_U3021) );
  OAI211_X1 U20069 ( .C1(n16814), .C2(n16813), .A(n16812), .B(n16811), .ZN(
        n16815) );
  AOI21_X1 U20070 ( .B1(n16816), .B2(n17076), .A(n16815), .ZN(n16817) );
  OAI21_X1 U20071 ( .B1(n17105), .B2(n16818), .A(n16817), .ZN(n16819) );
  AOI21_X1 U20072 ( .B1(n17748), .B2(n16820), .A(n16819), .ZN(n16821) );
  OAI21_X1 U20073 ( .B1(n17082), .B2(n16822), .A(n16821), .ZN(P2_U3022) );
  INV_X1 U20074 ( .A(n16823), .ZN(n16838) );
  OAI211_X1 U20075 ( .C1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n16838), .B(n16824), .ZN(
        n16825) );
  OAI211_X1 U20076 ( .C1(n16842), .C2(n22170), .A(n16826), .B(n16825), .ZN(
        n16829) );
  NOR2_X1 U20077 ( .A1(n16827), .A2(n17745), .ZN(n16828) );
  AOI211_X1 U20078 ( .C1(n16830), .C2(n17741), .A(n16829), .B(n16828), .ZN(
        n16833) );
  NAND2_X1 U20079 ( .A1(n16831), .A2(n17748), .ZN(n16832) );
  OAI211_X1 U20080 ( .C1(n16834), .C2(n17082), .A(n16833), .B(n16832), .ZN(
        P2_U3023) );
  NAND2_X1 U20081 ( .A1(n16835), .A2(n17738), .ZN(n16846) );
  NAND2_X1 U20082 ( .A1(n16836), .A2(n17076), .ZN(n16840) );
  AOI21_X1 U20083 ( .B1(n16838), .B2(n16841), .A(n16837), .ZN(n16839) );
  OAI211_X1 U20084 ( .C1(n16842), .C2(n16841), .A(n16840), .B(n16839), .ZN(
        n16843) );
  AOI21_X1 U20085 ( .B1(n17741), .B2(n16844), .A(n16843), .ZN(n16845) );
  OAI211_X1 U20086 ( .C1(n16847), .C2(n17101), .A(n16846), .B(n16845), .ZN(
        P2_U3024) );
  INV_X1 U20087 ( .A(n16989), .ZN(n16976) );
  OAI21_X1 U20088 ( .B1(n16976), .B2(n16849), .A(n16848), .ZN(n16852) );
  AOI21_X1 U20089 ( .B1(n16852), .B2(n16851), .A(n16850), .ZN(n16853) );
  OAI21_X1 U20090 ( .B1(n16854), .B2(n17745), .A(n16853), .ZN(n16856) );
  OAI21_X1 U20091 ( .B1(n16859), .B2(n17101), .A(n16858), .ZN(P2_U3025) );
  NAND2_X1 U20092 ( .A1(n16861), .A2(n16860), .ZN(n16870) );
  AND2_X1 U20093 ( .A1(n17111), .A2(n16893), .ZN(n16862) );
  NOR2_X1 U20094 ( .A1(n16926), .A2(n16862), .ZN(n16897) );
  NAND2_X1 U20095 ( .A1(n17111), .A2(n22065), .ZN(n16863) );
  NAND2_X1 U20096 ( .A1(n16897), .A2(n16863), .ZN(n16884) );
  NAND3_X1 U20097 ( .A1(n16865), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n16864), .ZN(n16866) );
  NOR2_X1 U20098 ( .A1(n16892), .A2(n16866), .ZN(n16882) );
  OAI21_X1 U20099 ( .B1(n16884), .B2(n16882), .A(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n16869) );
  INV_X1 U20100 ( .A(n16867), .ZN(n16868) );
  OAI211_X1 U20101 ( .C1(n16892), .C2(n16870), .A(n16869), .B(n16868), .ZN(
        n16871) );
  AOI21_X1 U20102 ( .B1(n16872), .B2(n17076), .A(n16871), .ZN(n16873) );
  OAI21_X1 U20103 ( .B1(n17105), .B2(n16874), .A(n16873), .ZN(n16875) );
  AOI21_X1 U20104 ( .B1(n16876), .B2(n17738), .A(n16875), .ZN(n16877) );
  OAI21_X1 U20105 ( .B1(n16878), .B2(n17101), .A(n16877), .ZN(P2_U3026) );
  NAND2_X1 U20106 ( .A1(n16880), .A2(n17076), .ZN(n16886) );
  OR2_X1 U20107 ( .A1(n16882), .A2(n16881), .ZN(n16883) );
  AOI21_X1 U20108 ( .B1(n16884), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n16883), .ZN(n16885) );
  OAI211_X1 U20109 ( .C1(n16887), .C2(n17105), .A(n16886), .B(n16885), .ZN(
        n16888) );
  AOI21_X1 U20110 ( .B1(n16889), .B2(n17738), .A(n16888), .ZN(n16890) );
  OAI21_X1 U20111 ( .B1(n16891), .B2(n17101), .A(n16890), .ZN(P2_U3027) );
  INV_X1 U20112 ( .A(n16892), .ZN(n16925) );
  NOR2_X1 U20113 ( .A1(n16893), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n16895) );
  AOI21_X1 U20114 ( .B1(n16925), .B2(n16895), .A(n16894), .ZN(n16896) );
  OAI21_X1 U20115 ( .B1(n16897), .B2(n22065), .A(n16896), .ZN(n16898) );
  INV_X1 U20116 ( .A(n16898), .ZN(n16901) );
  NAND2_X1 U20117 ( .A1(n16899), .A2(n17741), .ZN(n16900) );
  OAI211_X1 U20118 ( .C1(n16902), .C2(n17745), .A(n16901), .B(n16900), .ZN(
        n16903) );
  AOI21_X1 U20119 ( .B1(n16904), .B2(n17738), .A(n16903), .ZN(n16905) );
  OAI21_X1 U20120 ( .B1(n16906), .B2(n17101), .A(n16905), .ZN(P2_U3028) );
  OAI21_X1 U20121 ( .B1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17071), .A(
        n16907), .ZN(n16908) );
  NAND2_X1 U20122 ( .A1(n16908), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n16919) );
  OAI21_X1 U20123 ( .B1(n16910), .B2(n17745), .A(n16909), .ZN(n16916) );
  NAND2_X1 U20124 ( .A1(n16925), .A2(n16912), .ZN(n16913) );
  OAI211_X1 U20125 ( .C1(n16920), .C2(n17101), .A(n16919), .B(n16918), .ZN(
        P2_U3029) );
  INV_X1 U20126 ( .A(n16921), .ZN(n16933) );
  INV_X1 U20127 ( .A(n16922), .ZN(n16929) );
  AOI21_X1 U20128 ( .B1(n16925), .B2(n16924), .A(n16923), .ZN(n16928) );
  NAND2_X1 U20129 ( .A1(n16926), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16927) );
  OAI211_X1 U20130 ( .C1(n16929), .C2(n17745), .A(n16928), .B(n16927), .ZN(
        n16932) );
  NOR2_X1 U20131 ( .A1(n16930), .A2(n17101), .ZN(n16931) );
  AOI211_X1 U20132 ( .C1(n17741), .C2(n16933), .A(n16932), .B(n16931), .ZN(
        n16934) );
  OAI21_X1 U20133 ( .B1(n17082), .B2(n16935), .A(n16934), .ZN(P2_U3031) );
  NOR2_X1 U20134 ( .A1(n16938), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n16951) );
  NOR2_X1 U20135 ( .A1(n16938), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n16966) );
  OR2_X1 U20136 ( .A1(n16966), .A2(n16978), .ZN(n16952) );
  NOR2_X1 U20137 ( .A1(n16951), .A2(n16952), .ZN(n16943) );
  INV_X1 U20138 ( .A(n16936), .ZN(n16937) );
  OR3_X1 U20139 ( .A1(n16938), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        n16937), .ZN(n16941) );
  INV_X1 U20140 ( .A(n16939), .ZN(n16940) );
  OAI211_X1 U20141 ( .C1(n16943), .C2(n16942), .A(n16941), .B(n16940), .ZN(
        n16945) );
  NOR2_X1 U20142 ( .A1(n20241), .A2(n17745), .ZN(n16944) );
  AOI211_X1 U20143 ( .C1(n20245), .C2(n17741), .A(n16945), .B(n16944), .ZN(
        n16948) );
  NAND2_X1 U20144 ( .A1(n16946), .A2(n17748), .ZN(n16947) );
  OAI211_X1 U20145 ( .C1(n16949), .C2(n17082), .A(n16948), .B(n16947), .ZN(
        P2_U3032) );
  NAND2_X1 U20146 ( .A1(n16950), .A2(n17738), .ZN(n16962) );
  INV_X1 U20147 ( .A(n16951), .ZN(n16956) );
  NAND2_X1 U20148 ( .A1(n16952), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n16954) );
  OAI211_X1 U20149 ( .C1(n16956), .C2(n16955), .A(n16954), .B(n16953), .ZN(
        n16959) );
  NOR2_X1 U20150 ( .A1(n16957), .A2(n17105), .ZN(n16958) );
  AOI211_X1 U20151 ( .C1(n16960), .C2(n17076), .A(n16959), .B(n16958), .ZN(
        n16961) );
  OAI211_X1 U20152 ( .C1(n16963), .C2(n17101), .A(n16962), .B(n16961), .ZN(
        P2_U3033) );
  NOR2_X1 U20153 ( .A1(n16964), .A2(n17105), .ZN(n16971) );
  NOR2_X1 U20154 ( .A1(n16966), .A2(n16965), .ZN(n16968) );
  NAND2_X1 U20155 ( .A1(n16978), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n16967) );
  OAI211_X1 U20156 ( .C1(n16969), .C2(n17745), .A(n16968), .B(n16967), .ZN(
        n16970) );
  AOI211_X1 U20157 ( .C1(n16972), .C2(n17748), .A(n16971), .B(n16970), .ZN(
        n16973) );
  OAI21_X1 U20158 ( .B1(n16974), .B2(n17082), .A(n16973), .ZN(P2_U3034) );
  NAND2_X1 U20159 ( .A1(n16975), .A2(n17741), .ZN(n16981) );
  OAI21_X1 U20160 ( .B1(n16976), .B2(n16992), .A(n22118), .ZN(n16979) );
  AOI21_X1 U20161 ( .B1(n16979), .B2(n16978), .A(n16977), .ZN(n16980) );
  OAI211_X1 U20162 ( .C1(n16982), .C2(n17745), .A(n16981), .B(n16980), .ZN(
        n16983) );
  AOI21_X1 U20163 ( .B1(n16984), .B2(n17748), .A(n16983), .ZN(n16985) );
  OAI21_X1 U20164 ( .B1(n16986), .B2(n17082), .A(n16985), .ZN(P2_U3035) );
  NAND2_X1 U20165 ( .A1(n16987), .A2(n17076), .ZN(n16991) );
  AOI21_X1 U20166 ( .B1(n16989), .B2(n16992), .A(n16988), .ZN(n16990) );
  OAI211_X1 U20167 ( .C1(n16993), .C2(n16992), .A(n16991), .B(n16990), .ZN(
        n16994) );
  AOI21_X1 U20168 ( .B1(n17741), .B2(n16995), .A(n16994), .ZN(n16999) );
  NAND3_X1 U20169 ( .A1(n16997), .A2(n17738), .A3(n16996), .ZN(n16998) );
  OAI211_X1 U20170 ( .C1(n17000), .C2(n17101), .A(n16999), .B(n16998), .ZN(
        P2_U3036) );
  INV_X1 U20171 ( .A(n17023), .ZN(n17004) );
  NOR2_X1 U20172 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n17001), .ZN(
        n17003) );
  AOI21_X1 U20173 ( .B1(n17004), .B2(n17003), .A(n17002), .ZN(n17005) );
  OAI21_X1 U20174 ( .B1(n17007), .B2(n17006), .A(n17005), .ZN(n17009) );
  NOR2_X1 U20175 ( .A1(n20261), .A2(n17745), .ZN(n17008) );
  AOI211_X1 U20176 ( .C1(n17010), .C2(n17741), .A(n17009), .B(n17008), .ZN(
        n17013) );
  NAND2_X1 U20177 ( .A1(n17011), .A2(n17748), .ZN(n17012) );
  OAI211_X1 U20178 ( .C1(n17014), .C2(n17082), .A(n17013), .B(n17012), .ZN(
        P2_U3037) );
  NAND3_X1 U20179 ( .A1(n16727), .A2(n17015), .A3(n17738), .ZN(n17034) );
  INV_X1 U20180 ( .A(n17026), .ZN(n17024) );
  NAND2_X1 U20181 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n17024), .ZN(
        n17018) );
  INV_X1 U20182 ( .A(n17016), .ZN(n17017) );
  AOI22_X1 U20183 ( .A1(n17019), .A2(n17018), .B1(n17070), .B2(n17017), .ZN(
        n17020) );
  NAND2_X1 U20184 ( .A1(n17021), .A2(n17020), .ZN(n17050) );
  AND2_X1 U20185 ( .A1(n17070), .A2(n22168), .ZN(n17022) );
  NOR2_X1 U20186 ( .A1(n17050), .A2(n17022), .ZN(n17039) );
  NOR2_X1 U20187 ( .A1(n17069), .A2(n17023), .ZN(n17072) );
  NAND4_X1 U20188 ( .A1(n22145), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A3(
        n17072), .A4(n17024), .ZN(n17038) );
  AOI21_X1 U20189 ( .B1(n17039), .B2(n17038), .A(n17025), .ZN(n17029) );
  INV_X1 U20190 ( .A(n17072), .ZN(n17752) );
  OR2_X1 U20191 ( .A1(n17026), .A2(n17752), .ZN(n17047) );
  NAND2_X1 U20192 ( .A1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n21952) );
  NOR3_X1 U20193 ( .A1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n17047), .A3(
        n21952), .ZN(n17027) );
  NOR3_X1 U20194 ( .A1(n17029), .A2(n17028), .A3(n17027), .ZN(n17030) );
  OAI21_X1 U20195 ( .B1(n17745), .B2(n17031), .A(n17030), .ZN(n17032) );
  AOI21_X1 U20196 ( .B1(n17741), .B2(n20285), .A(n17032), .ZN(n17033) );
  OAI211_X1 U20197 ( .C1(n17035), .C2(n17101), .A(n17034), .B(n17033), .ZN(
        P2_U3038) );
  INV_X1 U20198 ( .A(n20278), .ZN(n17041) );
  INV_X1 U20199 ( .A(n17036), .ZN(n17037) );
  OAI211_X1 U20200 ( .C1(n17039), .C2(n22145), .A(n17038), .B(n17037), .ZN(
        n17040) );
  AOI21_X1 U20201 ( .B1(n17076), .B2(n17041), .A(n17040), .ZN(n17042) );
  OAI21_X1 U20202 ( .B1(n17105), .B2(n20275), .A(n17042), .ZN(n17043) );
  AOI21_X1 U20203 ( .B1(n17044), .B2(n17748), .A(n17043), .ZN(n17045) );
  OAI21_X1 U20204 ( .B1(n17046), .B2(n17082), .A(n17045), .ZN(P2_U3039) );
  NOR2_X1 U20205 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n17047), .ZN(
        n17048) );
  AOI211_X1 U20206 ( .C1(n17050), .C2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n17049), .B(n17048), .ZN(n17053) );
  NAND2_X1 U20207 ( .A1(n17051), .A2(n17741), .ZN(n17052) );
  OAI211_X1 U20208 ( .C1(n17054), .C2(n17745), .A(n17053), .B(n17052), .ZN(
        n17055) );
  AOI21_X1 U20209 ( .B1(n17056), .B2(n17748), .A(n17055), .ZN(n17057) );
  OAI21_X1 U20210 ( .B1(n17058), .B2(n17082), .A(n17057), .ZN(P2_U3040) );
  OR2_X1 U20211 ( .A1(n16751), .A2(n17059), .ZN(n17064) );
  OR2_X1 U20212 ( .A1(n17062), .A2(n17061), .ZN(n17063) );
  INV_X1 U20213 ( .A(n17720), .ZN(n17083) );
  INV_X1 U20214 ( .A(n17065), .ZN(n17066) );
  XNOR2_X1 U20215 ( .A(n17067), .B(n17066), .ZN(n17719) );
  AOI21_X1 U20216 ( .B1(n17070), .B2(n17069), .A(n17068), .ZN(n17750) );
  OAI21_X1 U20217 ( .B1(n17071), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n17750), .ZN(n17092) );
  NAND2_X1 U20218 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n17072), .ZN(
        n17091) );
  AOI221_X1 U20219 ( .B1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .C1(n17073), .C2(n17097), .A(
        n17091), .ZN(n17075) );
  NOR2_X1 U20220 ( .A1(n20217), .A2(n21038), .ZN(n17074) );
  AOI211_X1 U20221 ( .C1(n17092), .C2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n17075), .B(n17074), .ZN(n17078) );
  NAND2_X1 U20222 ( .A1(n17718), .A2(n17076), .ZN(n17077) );
  OAI211_X1 U20223 ( .C1(n17079), .C2(n17105), .A(n17078), .B(n17077), .ZN(
        n17080) );
  AOI21_X1 U20224 ( .B1(n17719), .B2(n17748), .A(n17080), .ZN(n17081) );
  OAI21_X1 U20225 ( .B1(n17083), .B2(n17082), .A(n17081), .ZN(P2_U3041) );
  INV_X1 U20226 ( .A(n17084), .ZN(n17085) );
  NAND2_X1 U20227 ( .A1(n17085), .A2(n17751), .ZN(n17727) );
  NAND2_X1 U20228 ( .A1(n17084), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n17726) );
  NAND2_X1 U20229 ( .A1(n17726), .A2(n17086), .ZN(n17087) );
  NAND2_X1 U20230 ( .A1(n17727), .A2(n17087), .ZN(n17090) );
  XNOR2_X1 U20231 ( .A(n17088), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n17089) );
  XNOR2_X1 U20232 ( .A(n17090), .B(n17089), .ZN(n20359) );
  INV_X1 U20233 ( .A(n20359), .ZN(n17102) );
  OAI22_X1 U20234 ( .A1(n20362), .A2(n17745), .B1(n21036), .B2(n20217), .ZN(
        n17095) );
  INV_X1 U20235 ( .A(n17091), .ZN(n17093) );
  MUX2_X1 U20236 ( .A(n17093), .B(n17092), .S(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .Z(n17094) );
  AOI211_X1 U20237 ( .C1(n17741), .C2(n17096), .A(n17095), .B(n17094), .ZN(
        n17100) );
  XNOR2_X1 U20238 ( .A(n17098), .B(n17097), .ZN(n20358) );
  NAND2_X1 U20239 ( .A1(n20358), .A2(n17738), .ZN(n17099) );
  OAI211_X1 U20240 ( .C1(n17102), .C2(n17101), .A(n17100), .B(n17099), .ZN(
        P2_U3042) );
  INV_X1 U20241 ( .A(n17103), .ZN(n17108) );
  INV_X1 U20242 ( .A(n20295), .ZN(n17122) );
  OAI22_X1 U20243 ( .A1(n17105), .A2(n17122), .B1(n17104), .B2(n17745), .ZN(
        n17106) );
  AOI211_X1 U20244 ( .C1(n17108), .C2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n17107), .B(n17106), .ZN(n17117) );
  NAND2_X1 U20245 ( .A1(n17738), .A2(n17109), .ZN(n17116) );
  OAI211_X1 U20246 ( .C1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(n17111), .B(n17110), .ZN(n17115) );
  NAND3_X1 U20247 ( .A1(n17748), .A2(n17113), .A3(n17112), .ZN(n17114) );
  NAND4_X1 U20248 ( .A1(n17117), .A2(n17116), .A3(n17115), .A4(n17114), .ZN(
        P2_U3045) );
  INV_X1 U20249 ( .A(n21110), .ZN(n17119) );
  AND2_X1 U20250 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n17118) );
  OR2_X1 U20251 ( .A1(n17119), .A2(n17118), .ZN(n17120) );
  MUX2_X1 U20252 ( .A(n21098), .B(n17120), .S(n20672), .Z(n17121) );
  OAI21_X1 U20253 ( .B1(n17122), .B2(n21106), .A(n17121), .ZN(n17125) );
  INV_X1 U20254 ( .A(n17806), .ZN(n17640) );
  OAI21_X1 U20255 ( .B1(n21119), .B2(P2_FLUSH_REG_SCAN_IN), .A(n17640), .ZN(
        n17123) );
  INV_X1 U20256 ( .A(n17123), .ZN(n17124) );
  OR2_X1 U20257 ( .A1(n20941), .A2(n17124), .ZN(n21112) );
  INV_X1 U20258 ( .A(n21112), .ZN(n21115) );
  MUX2_X1 U20259 ( .A(n17125), .B(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        n21115), .Z(P2_U3604) );
  NAND2_X1 U20260 ( .A1(n17127), .A2(n17126), .ZN(n17139) );
  MUX2_X1 U20261 ( .A(n17139), .B(n17150), .S(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n17128) );
  AOI21_X1 U20262 ( .B1(n13778), .B2(n17145), .A(n17128), .ZN(n17758) );
  OAI21_X1 U20263 ( .B1(n17758), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n11279), 
        .ZN(n17133) );
  MUX2_X1 U20264 ( .A(n17130), .B(n17129), .S(n20250), .Z(n17131) );
  NOR2_X1 U20265 ( .A1(n17131), .A2(n11279), .ZN(n17159) );
  INV_X1 U20266 ( .A(n17159), .ZN(n17132) );
  AOI22_X1 U20267 ( .A1(n17798), .A2(n21111), .B1(n17133), .B2(n17132), .ZN(
        n17135) );
  NAND2_X1 U20268 ( .A1(n17168), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n17134) );
  OAI21_X1 U20269 ( .B1(n17135), .B2(n17168), .A(n17134), .ZN(P2_U3601) );
  NAND2_X1 U20270 ( .A1(n20233), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17136) );
  NAND2_X1 U20271 ( .A1(n17137), .A2(n17136), .ZN(n17160) );
  INV_X1 U20272 ( .A(n17160), .ZN(n17142) );
  NAND2_X1 U20273 ( .A1(n13801), .A2(n17145), .ZN(n17141) );
  AOI22_X1 U20274 ( .A1(n17150), .A2(n10702), .B1(n17139), .B2(n17138), .ZN(
        n17140) );
  NAND2_X1 U20275 ( .A1(n17141), .A2(n17140), .ZN(n17755) );
  AOI222_X1 U20276 ( .A1(n20672), .A2(n17798), .B1(n17159), .B2(n17142), .C1(
        n17755), .C2(n21086), .ZN(n17144) );
  NAND2_X1 U20277 ( .A1(n17168), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n17143) );
  OAI21_X1 U20278 ( .B1(n17144), .B2(n17168), .A(n17143), .ZN(P2_U3600) );
  NAND2_X1 U20279 ( .A1(n17146), .A2(n17145), .ZN(n17158) );
  NOR2_X1 U20280 ( .A1(n17148), .A2(n17147), .ZN(n17154) );
  NOR2_X1 U20281 ( .A1(n17149), .A2(n10693), .ZN(n17151) );
  AOI22_X1 U20282 ( .A1(n17152), .A2(n17154), .B1(n17151), .B2(n17150), .ZN(
        n17153) );
  OAI21_X1 U20283 ( .B1(n17155), .B2(n17154), .A(n17153), .ZN(n17156) );
  INV_X1 U20284 ( .A(n17156), .ZN(n17157) );
  NAND2_X1 U20285 ( .A1(n17158), .A2(n17157), .ZN(n17761) );
  AOI222_X1 U20286 ( .A1(n17160), .A2(n17159), .B1(n20373), .B2(n17798), .C1(
        n17761), .C2(n21086), .ZN(n17162) );
  NAND2_X1 U20287 ( .A1(n17168), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n17161) );
  OAI21_X1 U20288 ( .B1(n17162), .B2(n17168), .A(n17161), .ZN(P2_U3599) );
  INV_X1 U20289 ( .A(n17163), .ZN(n17164) );
  NAND2_X1 U20290 ( .A1(n17165), .A2(n17164), .ZN(n17166) );
  NOR2_X1 U20291 ( .A1(n17167), .A2(n17166), .ZN(n17767) );
  AND2_X1 U20292 ( .A1(n17767), .A2(n21086), .ZN(n17169) );
  MUX2_X1 U20293 ( .A(n17169), .B(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n17168), .Z(P2_U3595) );
  NAND2_X1 U20294 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n19521) );
  NAND2_X1 U20295 ( .A1(n20138), .A2(n19521), .ZN(n20178) );
  NAND2_X1 U20296 ( .A1(n17927), .A2(n17170), .ZN(n20014) );
  INV_X1 U20297 ( .A(n20014), .ZN(n17171) );
  NAND2_X1 U20298 ( .A1(n20015), .A2(n17171), .ZN(n17172) );
  NOR2_X1 U20299 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n18996), .ZN(
        n17829) );
  INV_X1 U20300 ( .A(n19068), .ZN(n19113) );
  NAND2_X1 U20301 ( .A1(n20044), .A2(n20187), .ZN(n20174) );
  NAND3_X1 U20302 ( .A1(n20187), .A2(n20138), .A3(P3_STATEBS16_REG_SCAN_IN), 
        .ZN(n19830) );
  NOR2_X1 U20303 ( .A1(n19882), .A2(n9880), .ZN(n17819) );
  AOI211_X1 U20304 ( .C1(n17174), .C2(n19113), .A(n19231), .B(n17819), .ZN(
        n17175) );
  INV_X1 U20305 ( .A(n17175), .ZN(n17818) );
  NOR2_X1 U20306 ( .A1(n17829), .A2(n17818), .ZN(n17813) );
  INV_X1 U20307 ( .A(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n18574) );
  OAI22_X1 U20308 ( .A1(n18613), .A2(n17176), .B1(n18615), .B2(n18574), .ZN(
        n17178) );
  INV_X1 U20309 ( .A(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n18565) );
  INV_X1 U20310 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n18654) );
  OAI22_X1 U20311 ( .A1(n18616), .A2(n18565), .B1(n11880), .B2(n18654), .ZN(
        n17177) );
  NOR2_X1 U20312 ( .A1(n17178), .A2(n17177), .ZN(n17185) );
  INV_X1 U20313 ( .A(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17515) );
  NAND2_X1 U20314 ( .A1(n18620), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n17180) );
  INV_X1 U20315 ( .A(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n18430) );
  NAND2_X1 U20316 ( .A1(n18619), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n17179) );
  OAI211_X1 U20317 ( .C1(n17550), .C2(n17515), .A(n17180), .B(n17179), .ZN(
        n17181) );
  INV_X1 U20318 ( .A(n17181), .ZN(n17184) );
  AOI22_X1 U20319 ( .A1(n18586), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11911), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17183) );
  NAND2_X1 U20320 ( .A1(n18413), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n17182) );
  NAND4_X1 U20321 ( .A1(n17185), .A2(n17184), .A3(n17183), .A4(n17182), .ZN(
        n17191) );
  AOI22_X1 U20322 ( .A1(n18626), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n18390), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17189) );
  AOI22_X1 U20323 ( .A1(n9724), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n18403), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17188) );
  INV_X1 U20324 ( .A(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n18576) );
  OR2_X1 U20325 ( .A1(n18599), .A2(n18576), .ZN(n17187) );
  NAND2_X1 U20326 ( .A1(n9726), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n17186) );
  NAND4_X1 U20327 ( .A1(n17189), .A2(n17188), .A3(n17187), .A4(n17186), .ZN(
        n17190) );
  NAND2_X1 U20328 ( .A1(n17547), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n17195) );
  NAND2_X1 U20329 ( .A1(n9724), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n17194) );
  NAND2_X1 U20330 ( .A1(n18597), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n17193) );
  INV_X1 U20331 ( .A(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n18391) );
  NAND2_X1 U20332 ( .A1(n14232), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n17192) );
  AND4_X1 U20333 ( .A1(n17195), .A2(n17194), .A3(n17193), .A4(n17192), .ZN(
        n17202) );
  NAND2_X1 U20334 ( .A1(n18620), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n17197) );
  NAND2_X1 U20335 ( .A1(n18489), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n17196) );
  OAI211_X1 U20336 ( .C1(n17550), .C2(n17542), .A(n17197), .B(n17196), .ZN(
        n17198) );
  INV_X1 U20337 ( .A(n17198), .ZN(n17201) );
  AOI22_X1 U20338 ( .A1(n18586), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17561), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17200) );
  NAND2_X1 U20339 ( .A1(n18413), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n17199) );
  NAND4_X1 U20340 ( .A1(n17202), .A2(n17201), .A3(n17200), .A4(n17199), .ZN(
        n17208) );
  AOI22_X1 U20341 ( .A1(n18585), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11911), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n17206) );
  AOI22_X1 U20342 ( .A1(n18390), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n18403), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n17205) );
  INV_X1 U20343 ( .A(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n18396) );
  OR2_X1 U20344 ( .A1(n18599), .A2(n18396), .ZN(n17204) );
  NAND2_X1 U20345 ( .A1(n9726), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n17203) );
  NAND4_X1 U20346 ( .A1(n17206), .A2(n17205), .A3(n17204), .A4(n17203), .ZN(
        n17207) );
  OR2_X1 U20347 ( .A1(n18806), .A2(n17287), .ZN(n17209) );
  INV_X1 U20348 ( .A(n17281), .ZN(n17283) );
  AOI22_X1 U20349 ( .A1(n17547), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n9724), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n17214) );
  AOI22_X1 U20350 ( .A1(n18620), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n18619), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n17213) );
  INV_X1 U20351 ( .A(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n18506) );
  INV_X1 U20352 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n18637) );
  OAI22_X1 U20353 ( .A1(n18613), .A2(n18506), .B1(n9723), .B2(n18637), .ZN(
        n17210) );
  INV_X1 U20354 ( .A(n17210), .ZN(n17212) );
  NAND2_X1 U20355 ( .A1(n18586), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n17211) );
  AOI22_X1 U20356 ( .A1(n18390), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n18403), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n17218) );
  INV_X1 U20357 ( .A(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n21957) );
  AOI22_X1 U20358 ( .A1(n18626), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11911), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n17217) );
  INV_X1 U20359 ( .A(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n18318) );
  OR2_X1 U20360 ( .A1(n18599), .A2(n18318), .ZN(n17216) );
  NAND2_X1 U20361 ( .A1(n9726), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n17215) );
  INV_X1 U20362 ( .A(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17221) );
  NAND2_X1 U20363 ( .A1(n18591), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n17220) );
  NAND2_X1 U20364 ( .A1(n14232), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n17219) );
  OAI211_X1 U20365 ( .C1(n17550), .C2(n17221), .A(n17220), .B(n17219), .ZN(
        n17222) );
  INV_X1 U20366 ( .A(n17222), .ZN(n17223) );
  INV_X1 U20367 ( .A(n17226), .ZN(n17235) );
  OR2_X1 U20368 ( .A1(n17295), .A2(n17278), .ZN(n17227) );
  NAND2_X1 U20369 ( .A1(n17235), .A2(n17227), .ZN(n17231) );
  XNOR2_X1 U20370 ( .A(n17231), .B(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n17355) );
  NAND2_X1 U20371 ( .A1(n17228), .A2(n10672), .ZN(n17230) );
  OR2_X1 U20372 ( .A1(n17295), .A2(n17443), .ZN(n17229) );
  NAND2_X1 U20373 ( .A1(n17230), .A2(n17229), .ZN(n17354) );
  NAND2_X1 U20374 ( .A1(n17355), .A2(n17354), .ZN(n17234) );
  INV_X1 U20375 ( .A(n17231), .ZN(n17232) );
  NAND2_X1 U20376 ( .A1(n17232), .A2(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n17233) );
  NAND2_X1 U20377 ( .A1(n17234), .A2(n17233), .ZN(n19238) );
  XNOR2_X1 U20378 ( .A(n18811), .B(n17235), .ZN(n19236) );
  INV_X1 U20379 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n19511) );
  NAND2_X1 U20380 ( .A1(n19236), .A2(n19511), .ZN(n17236) );
  INV_X1 U20381 ( .A(n19236), .ZN(n17237) );
  NAND2_X1 U20382 ( .A1(n17237), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n17238) );
  XNOR2_X1 U20383 ( .A(n17239), .B(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n19224) );
  INV_X1 U20384 ( .A(n17239), .ZN(n17240) );
  NAND2_X1 U20385 ( .A1(n17240), .A2(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n17241) );
  OR2_X1 U20386 ( .A1(n17242), .A2(n17287), .ZN(n17243) );
  XNOR2_X1 U20387 ( .A(n17243), .B(n18806), .ZN(n19209) );
  INV_X1 U20388 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n19482) );
  NAND2_X1 U20389 ( .A1(n19209), .A2(n19482), .ZN(n17244) );
  INV_X1 U20390 ( .A(n19209), .ZN(n17245) );
  NAND2_X1 U20391 ( .A1(n17245), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n17246) );
  XNOR2_X1 U20392 ( .A(n17247), .B(n17281), .ZN(n17249) );
  INV_X1 U20393 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n17248) );
  XNOR2_X1 U20394 ( .A(n17249), .B(n17248), .ZN(n19195) );
  NAND2_X1 U20395 ( .A1(n17407), .A2(n18802), .ZN(n17250) );
  NAND2_X1 U20396 ( .A1(n19185), .A2(n17250), .ZN(n17251) );
  XNOR2_X1 U20397 ( .A(n17253), .B(n17251), .ZN(n17350) );
  INV_X1 U20398 ( .A(n17251), .ZN(n17252) );
  NAND2_X1 U20399 ( .A1(n17253), .A2(n17252), .ZN(n17254) );
  NAND2_X1 U20400 ( .A1(n17257), .A2(n19185), .ZN(n19161) );
  NAND2_X1 U20401 ( .A1(n19377), .A2(n19101), .ZN(n19364) );
  OR2_X1 U20402 ( .A1(n19364), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n17258) );
  NAND2_X1 U20403 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n19146) );
  NOR2_X1 U20404 ( .A1(n19146), .A2(n19138), .ZN(n19423) );
  NAND2_X1 U20405 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n19423), .ZN(
        n19122) );
  NAND2_X1 U20406 ( .A1(n19379), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n19362) );
  INV_X1 U20407 ( .A(n19327), .ZN(n19062) );
  MUX2_X1 U20408 ( .A(n19185), .B(n17260), .S(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .Z(n17259) );
  NAND2_X1 U20409 ( .A1(n17262), .A2(n17259), .ZN(n19052) );
  OAI21_X2 U20410 ( .B1(n19052), .B2(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n19185), .ZN(n19020) );
  INV_X1 U20411 ( .A(n17260), .ZN(n17261) );
  NAND2_X1 U20412 ( .A1(n19064), .A2(n19331), .ZN(n17263) );
  NAND2_X1 U20413 ( .A1(n19020), .A2(n17263), .ZN(n19045) );
  AND2_X1 U20414 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17337) );
  NOR2_X1 U20415 ( .A1(n22088), .A2(n19319), .ZN(n19297) );
  AND2_X1 U20416 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n19297), .ZN(
        n17264) );
  AND2_X1 U20417 ( .A1(n18978), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n17265) );
  AND2_X1 U20418 ( .A1(n19045), .A2(n17265), .ZN(n17268) );
  NAND2_X1 U20419 ( .A1(n18978), .A2(n19331), .ZN(n17406) );
  NOR2_X1 U20420 ( .A1(n17406), .A2(n18988), .ZN(n17320) );
  INV_X1 U20421 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17266) );
  NAND2_X1 U20422 ( .A1(n19043), .A2(n19319), .ZN(n17267) );
  NOR2_X1 U20423 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17267), .ZN(
        n19010) );
  INV_X1 U20424 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n19286) );
  INV_X1 U20425 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n19288) );
  INV_X1 U20426 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17269) );
  INV_X1 U20427 ( .A(n17372), .ZN(n17416) );
  OAI21_X1 U20428 ( .B1(n18958), .B2(n17416), .A(n19063), .ZN(n17270) );
  INV_X1 U20429 ( .A(n17408), .ZN(n18939) );
  NAND3_X1 U20430 ( .A1(n18939), .A2(n19063), .A3(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17593) );
  INV_X1 U20431 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n17825) );
  INV_X1 U20432 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n19259) );
  INV_X1 U20433 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n21976) );
  INV_X1 U20434 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n17817) );
  OAI22_X1 U20435 ( .A1(n17272), .A2(n17632), .B1(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n17817), .ZN(n17276) );
  XNOR2_X1 U20436 ( .A(n19185), .B(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n17274) );
  AND2_X1 U20437 ( .A1(n17817), .A2(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n17317) );
  NOR2_X1 U20438 ( .A1(n17274), .A2(n17317), .ZN(n17275) );
  NOR2_X1 U20439 ( .A1(n17632), .A2(n19063), .ZN(n17273) );
  NAND2_X1 U20440 ( .A1(n17396), .A2(n19172), .ZN(n17331) );
  NOR2_X1 U20441 ( .A1(n20044), .A2(n17926), .ZN(n19067) );
  INV_X1 U20442 ( .A(n19067), .ZN(n19218) );
  INV_X1 U20443 ( .A(n17278), .ZN(n17291) );
  NAND2_X1 U20444 ( .A1(n17292), .A2(n17291), .ZN(n17289) );
  AND2_X1 U20445 ( .A1(n17289), .A2(n17279), .ZN(n17288) );
  INV_X1 U20446 ( .A(n17287), .ZN(n17280) );
  NAND2_X1 U20447 ( .A1(n17288), .A2(n17280), .ZN(n17285) );
  NOR2_X1 U20448 ( .A1(n17285), .A2(n18806), .ZN(n17284) );
  NAND2_X1 U20449 ( .A1(n17284), .A2(n17281), .ZN(n17282) );
  NOR2_X1 U20450 ( .A1(n18802), .A2(n17282), .ZN(n17314) );
  XOR2_X1 U20451 ( .A(n18802), .B(n17282), .Z(n17348) );
  XNOR2_X1 U20452 ( .A(n17284), .B(n17283), .ZN(n17307) );
  XOR2_X1 U20453 ( .A(n18806), .B(n17285), .Z(n17286) );
  NAND2_X1 U20454 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n17286), .ZN(
        n17306) );
  XOR2_X1 U20455 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B(n17286), .Z(
        n19206) );
  XNOR2_X1 U20456 ( .A(n17288), .B(n17287), .ZN(n17304) );
  NAND2_X1 U20457 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n17290), .ZN(
        n17302) );
  XNOR2_X1 U20458 ( .A(n17292), .B(n17291), .ZN(n17293) );
  NAND2_X1 U20459 ( .A1(n17293), .A2(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n17301) );
  XNOR2_X1 U20460 ( .A(n17293), .B(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n17357) );
  NAND2_X1 U20461 ( .A1(n17294), .A2(n22165), .ZN(n17298) );
  INV_X1 U20462 ( .A(n17295), .ZN(n17297) );
  MUX2_X1 U20463 ( .A(n17298), .B(n17297), .S(n17296), .Z(n17300) );
  NAND2_X1 U20464 ( .A1(n17300), .A2(n17299), .ZN(n17356) );
  NAND2_X1 U20465 ( .A1(n17304), .A2(n17303), .ZN(n17305) );
  NAND2_X1 U20466 ( .A1(n17307), .A2(n17308), .ZN(n17309) );
  INV_X1 U20467 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n19470) );
  NAND2_X1 U20468 ( .A1(n17314), .A2(n17310), .ZN(n17315) );
  NAND2_X1 U20469 ( .A1(n17348), .A2(n17347), .ZN(n17312) );
  NAND2_X1 U20470 ( .A1(n17314), .A2(n17313), .ZN(n17311) );
  OAI211_X1 U20471 ( .C1(n17314), .C2(n17313), .A(n17312), .B(n17311), .ZN(
        n19177) );
  NAND2_X1 U20472 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n19177), .ZN(
        n19176) );
  INV_X1 U20473 ( .A(n18956), .ZN(n17316) );
  AND2_X2 U20474 ( .A1(n17372), .A2(n17316), .ZN(n17425) );
  AND2_X1 U20475 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17318) );
  NAND2_X1 U20476 ( .A1(n17425), .A2(n17318), .ZN(n17824) );
  AND3_X1 U20477 ( .A1(n17394), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n17322) );
  INV_X1 U20478 ( .A(n17322), .ZN(n17391) );
  INV_X1 U20479 ( .A(n17317), .ZN(n17386) );
  NAND2_X1 U20480 ( .A1(n17318), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n17810) );
  INV_X1 U20481 ( .A(n17810), .ZN(n17379) );
  NAND2_X1 U20482 ( .A1(n17379), .A2(n17425), .ZN(n17809) );
  NAND2_X1 U20483 ( .A1(n17809), .A2(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n17319) );
  INV_X1 U20484 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n22186) );
  NOR2_X2 U20485 ( .A1(n19187), .A2(n17256), .ZN(n19418) );
  NAND2_X1 U20486 ( .A1(n19418), .A2(n19354), .ZN(n19104) );
  NAND2_X1 U20487 ( .A1(n19366), .A2(n17320), .ZN(n18969) );
  NOR2_X1 U20488 ( .A1(n22186), .A2(n18969), .ZN(n18950) );
  NAND2_X1 U20489 ( .A1(n17372), .A2(n18950), .ZN(n17422) );
  NOR2_X1 U20490 ( .A1(n17422), .A2(n17810), .ZN(n17808) );
  NAND2_X1 U20491 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17321) );
  NOR2_X1 U20492 ( .A1(n17422), .A2(n17321), .ZN(n17820) );
  NAND2_X1 U20493 ( .A1(n17820), .A2(n17322), .ZN(n17323) );
  OAI211_X1 U20494 ( .C1(n17808), .C2(n17394), .A(n17323), .B(n17386), .ZN(
        n17383) );
  NAND2_X1 U20495 ( .A1(n19145), .A2(n17383), .ZN(n17324) );
  NAND2_X1 U20496 ( .A1(n19508), .A2(P3_REIP_REG_31__SCAN_IN), .ZN(n17385) );
  OAI211_X1 U20497 ( .C1(n17325), .C2(n19235), .A(n17324), .B(n17385), .ZN(
        n17329) );
  AOI21_X1 U20498 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n17326), .A(
        n19921), .ZN(n19026) );
  INV_X1 U20499 ( .A(n19026), .ZN(n19070) );
  NAND2_X1 U20500 ( .A1(n9880), .A2(n19070), .ZN(n17814) );
  XNOR2_X1 U20501 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(
        P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n17327) );
  NOR2_X1 U20502 ( .A1(n17814), .A2(n17327), .ZN(n17328) );
  AOI211_X1 U20503 ( .C1(n19128), .C2(n17277), .A(n17329), .B(n17328), .ZN(
        n17330) );
  OAI211_X1 U20504 ( .C1(n17813), .C2(n17332), .A(n17331), .B(n17330), .ZN(
        P3_U2799) );
  INV_X1 U20505 ( .A(n17333), .ZN(n17336) );
  INV_X1 U20506 ( .A(n17334), .ZN(n17335) );
  AOI21_X1 U20507 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17336), .A(
        n17335), .ZN(n17432) );
  INV_X1 U20508 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n19263) );
  NAND2_X1 U20509 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17418) );
  AND3_X1 U20510 ( .A1(n19331), .A2(n17337), .A3(n19297), .ZN(n19283) );
  INV_X1 U20511 ( .A(n19283), .ZN(n19287) );
  INV_X1 U20512 ( .A(n19418), .ZN(n19144) );
  NOR3_X1 U20513 ( .A1(n19288), .A2(n19287), .A3(n19079), .ZN(n18975) );
  INV_X1 U20514 ( .A(n17422), .ZN(n17338) );
  OAI22_X1 U20515 ( .A1(n17338), .A2(n19105), .B1(n17425), .B2(n19235), .ZN(
        n18946) );
  INV_X1 U20516 ( .A(n17339), .ZN(n17340) );
  OAI21_X1 U20517 ( .B1(n17340), .B2(n19068), .A(n19207), .ZN(n17341) );
  AOI21_X1 U20518 ( .B1(n19067), .B2(n18924), .A(n17341), .ZN(n18922) );
  AOI21_X1 U20519 ( .B1(n11795), .B2(n19921), .A(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17343) );
  OAI21_X1 U20520 ( .B1(n19128), .B2(n17326), .A(n17984), .ZN(n17342) );
  NAND2_X1 U20521 ( .A1(n19508), .A2(P3_REIP_REG_26__SCAN_IN), .ZN(n17428) );
  OAI211_X1 U20522 ( .C1(n18922), .C2(n17343), .A(n17342), .B(n17428), .ZN(
        n17344) );
  NAND2_X1 U20523 ( .A1(n19118), .A2(n18996), .ZN(n19215) );
  NAND2_X1 U20524 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18206), .ZN(
        n18217) );
  NAND2_X1 U20525 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n9894), .ZN(
        n18197) );
  INV_X1 U20526 ( .A(n18197), .ZN(n17345) );
  AOI21_X1 U20527 ( .B1(n19165), .B2(n18217), .A(n17345), .ZN(n18208) );
  INV_X1 U20528 ( .A(n18208), .ZN(n17353) );
  NOR2_X1 U20529 ( .A1(n10079), .A2(n19882), .ZN(n19166) );
  OAI21_X1 U20530 ( .B1(n19218), .B2(n18206), .A(n19207), .ZN(n19178) );
  INV_X1 U20531 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n20084) );
  NOR2_X1 U20532 ( .A1(n14191), .A2(n20084), .ZN(n19467) );
  AOI221_X1 U20533 ( .B1(n19166), .B2(n19165), .C1(n19178), .C2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A(n19467), .ZN(n17352) );
  AOI21_X1 U20534 ( .B1(n17348), .B2(n17347), .A(n17346), .ZN(n17349) );
  XOR2_X1 U20535 ( .A(n17349), .B(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .Z(
        n19462) );
  INV_X1 U20536 ( .A(n19239), .ZN(n19190) );
  XOR2_X1 U20537 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B(n17350), .Z(
        n19463) );
  AOI22_X1 U20538 ( .A1(n10167), .A2(n19462), .B1(n19190), .B2(n19463), .ZN(
        n17351) );
  OAI211_X1 U20539 ( .C1(n19248), .C2(n17353), .A(n17352), .B(n17351), .ZN(
        P3_U2823) );
  XNOR2_X1 U20540 ( .A(n17355), .B(n17354), .ZN(n17450) );
  INV_X1 U20541 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n19230) );
  NAND2_X1 U20542 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n18254) );
  OAI21_X1 U20543 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n18254), .ZN(n18284) );
  NAND2_X1 U20544 ( .A1(n17357), .A2(n17356), .ZN(n17358) );
  NAND2_X1 U20545 ( .A1(n17359), .A2(n17358), .ZN(n17451) );
  OAI22_X1 U20546 ( .A1(n19248), .A2(n18284), .B1(n19235), .B2(n17451), .ZN(
        n17360) );
  AOI221_X1 U20547 ( .B1(n19231), .B2(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .C1(
        n19921), .C2(n19230), .A(n17360), .ZN(n17361) );
  NAND2_X1 U20548 ( .A1(n19508), .A2(P3_REIP_REG_2__SCAN_IN), .ZN(n17456) );
  OAI211_X1 U20549 ( .C1(n17450), .C2(n19239), .A(n17361), .B(n17456), .ZN(
        P3_U2828) );
  AOI22_X1 U20550 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n19194), .B1(
        n19215), .B2(n18301), .ZN(n17366) );
  INV_X1 U20551 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n17362) );
  OAI22_X1 U20552 ( .A1(n19239), .A2(n17363), .B1(n14191), .B2(n17362), .ZN(
        n17364) );
  INV_X1 U20553 ( .A(n17364), .ZN(n17365) );
  OAI211_X1 U20554 ( .C1(n17367), .C2(n19235), .A(n17366), .B(n17365), .ZN(
        P3_U2829) );
  NOR2_X1 U20555 ( .A1(n17368), .A2(n10672), .ZN(n19516) );
  NAND3_X1 U20556 ( .A1(n20044), .A2(n19207), .A3(n19068), .ZN(n17369) );
  AOI22_X1 U20557 ( .A1(n19508), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17369), .ZN(n17371) );
  NAND2_X1 U20558 ( .A1(n19190), .A2(n19516), .ZN(n17370) );
  OAI211_X1 U20559 ( .C1(n19516), .C2(n19235), .A(n17371), .B(n17370), .ZN(
        P3_U2830) );
  INV_X1 U20560 ( .A(n17418), .ZN(n19264) );
  NAND2_X1 U20561 ( .A1(n17372), .A2(n19264), .ZN(n19250) );
  NOR2_X1 U20562 ( .A1(n19259), .A2(n19250), .ZN(n18921) );
  NAND3_X1 U20563 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n19325) );
  NAND3_X1 U20564 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n19323) );
  INV_X1 U20565 ( .A(n19323), .ZN(n17374) );
  INV_X1 U20566 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n17452) );
  NOR2_X1 U20567 ( .A1(n17452), .A2(n17443), .ZN(n19490) );
  NAND2_X1 U20568 ( .A1(n17374), .A2(n19490), .ZN(n19441) );
  NOR2_X1 U20569 ( .A1(n19325), .A2(n19441), .ZN(n19348) );
  INV_X1 U20570 ( .A(n19348), .ZN(n17373) );
  NOR2_X1 U20571 ( .A1(n22165), .A2(n17373), .ZN(n19413) );
  NAND2_X1 U20572 ( .A1(n19327), .A2(n19413), .ZN(n19352) );
  NOR2_X1 U20573 ( .A1(n17406), .A2(n19352), .ZN(n17419) );
  AOI21_X1 U20574 ( .B1(n18921), .B2(n17419), .A(n19424), .ZN(n17378) );
  NOR2_X1 U20575 ( .A1(n19062), .A2(n17373), .ZN(n19328) );
  INV_X1 U20576 ( .A(n19328), .ZN(n17388) );
  NOR3_X1 U20577 ( .A1(n17406), .A2(n17388), .A3(n19250), .ZN(n17376) );
  INV_X1 U20578 ( .A(n19331), .ZN(n17375) );
  OAI21_X1 U20579 ( .B1(n17443), .B2(n22165), .A(n17452), .ZN(n19322) );
  NAND2_X1 U20580 ( .A1(n17374), .A2(n19322), .ZN(n19443) );
  NOR2_X1 U20581 ( .A1(n19443), .A2(n19325), .ZN(n19350) );
  NAND2_X1 U20582 ( .A1(n19327), .A2(n19350), .ZN(n19280) );
  NOR2_X1 U20583 ( .A1(n17375), .A2(n19280), .ZN(n19330) );
  NAND2_X1 U20584 ( .A1(n18978), .A2(n19330), .ZN(n17417) );
  NAND2_X1 U20585 ( .A1(n19444), .A2(n17417), .ZN(n17437) );
  OAI21_X1 U20586 ( .B1(n19349), .B2(n17376), .A(n17437), .ZN(n17377) );
  AOI211_X1 U20587 ( .C1(n19444), .C2(n19250), .A(n17378), .B(n17377), .ZN(
        n17399) );
  OR2_X1 U20588 ( .A1(n17399), .A2(n19517), .ZN(n17382) );
  OAI21_X1 U20589 ( .B1(n19493), .B2(n17379), .A(n19512), .ZN(n17380) );
  INV_X1 U20590 ( .A(n17380), .ZN(n17381) );
  AND2_X1 U20591 ( .A1(n17382), .A2(n17381), .ZN(n17639) );
  INV_X1 U20592 ( .A(n19505), .ZN(n19515) );
  NAND3_X1 U20593 ( .A1(n19515), .A2(n18802), .A3(n17383), .ZN(n17384) );
  OAI211_X1 U20594 ( .C1(n19493), .C2(n17386), .A(n17385), .B(n17384), .ZN(
        n17387) );
  AOI21_X1 U20595 ( .B1(n19986), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n19978), .ZN(n19320) );
  OAI22_X1 U20596 ( .A1(n20019), .A2(n19280), .B1(n19320), .B2(n17388), .ZN(
        n17405) );
  INV_X1 U20597 ( .A(n17405), .ZN(n17389) );
  NOR2_X1 U20598 ( .A1(n17389), .A2(n17406), .ZN(n19265) );
  AND2_X1 U20599 ( .A1(n18921), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n17390) );
  NAND2_X1 U20600 ( .A1(n19265), .A2(n17390), .ZN(n17587) );
  OR3_X1 U20601 ( .A1(n17587), .A2(n19517), .A3(n17391), .ZN(n17392) );
  OAI211_X1 U20602 ( .C1(n17639), .C2(n17394), .A(n17393), .B(n17392), .ZN(
        n17395) );
  AOI21_X1 U20603 ( .B1(n17396), .B2(n19455), .A(n17395), .ZN(n17397) );
  INV_X1 U20604 ( .A(n17397), .ZN(P3_U2831) );
  OR2_X1 U20605 ( .A1(n19188), .A2(n17398), .ZN(n19452) );
  NAND2_X1 U20606 ( .A1(n20019), .A2(n19349), .ZN(n19430) );
  OAI21_X1 U20607 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n19422), .A(
        n17399), .ZN(n17589) );
  AOI211_X1 U20608 ( .C1(n19416), .C2(n17824), .A(n19473), .B(n17589), .ZN(
        n17403) );
  XNOR2_X1 U20609 ( .A(n19185), .B(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n18932) );
  NAND2_X1 U20610 ( .A1(n17408), .A2(n19063), .ZN(n18941) );
  NAND2_X1 U20611 ( .A1(n18941), .A2(n17409), .ZN(n18931) );
  OAI211_X1 U20612 ( .C1(n17408), .C2(n17407), .A(n20015), .B(n19188), .ZN(
        n17400) );
  AOI21_X1 U20613 ( .B1(n18932), .B2(n18931), .A(n17400), .ZN(n17401) );
  INV_X1 U20614 ( .A(n17401), .ZN(n17402) );
  OAI211_X1 U20615 ( .C1(n17820), .C2(n19452), .A(n17403), .B(n17402), .ZN(
        n17404) );
  NAND3_X1 U20616 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n14191), .A3(
        n17404), .ZN(n17414) );
  OAI22_X1 U20617 ( .A1(n10378), .A2(n19415), .B1(n19144), .B2(n19452), .ZN(
        n19326) );
  AOI21_X1 U20618 ( .B1(n19326), .B2(n19327), .A(n17405), .ZN(n19293) );
  NOR2_X1 U20619 ( .A1(n17406), .A2(n19293), .ZN(n19273) );
  INV_X1 U20620 ( .A(n19273), .ZN(n19249) );
  NOR2_X1 U20621 ( .A1(n19517), .A2(n19249), .ZN(n17441) );
  NAND3_X1 U20622 ( .A1(n18921), .A2(n17441), .A3(n21976), .ZN(n17413) );
  NAND2_X1 U20623 ( .A1(n19508), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n18926) );
  NOR3_X1 U20624 ( .A1(n17408), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        n17407), .ZN(n17411) );
  NOR2_X1 U20625 ( .A1(n17409), .A2(n18932), .ZN(n17410) );
  OAI21_X1 U20626 ( .B1(n17411), .B2(n17410), .A(n19455), .ZN(n17412) );
  NAND4_X1 U20627 ( .A1(n17414), .A2(n17413), .A3(n18926), .A4(n17412), .ZN(
        P3_U2834) );
  INV_X1 U20628 ( .A(n19455), .ZN(n19428) );
  NAND2_X1 U20629 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n19264), .ZN(
        n17415) );
  NOR2_X1 U20630 ( .A1(n19249), .A2(n17415), .ZN(n17426) );
  AOI22_X1 U20631 ( .A1(n19978), .A2(n19263), .B1(n17416), .B2(n19306), .ZN(
        n17424) );
  INV_X1 U20632 ( .A(n19452), .ZN(n19282) );
  OAI21_X1 U20633 ( .B1(n17418), .B2(n17417), .A(n19444), .ZN(n17421) );
  AOI21_X1 U20634 ( .B1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n19424), .A(
        n17419), .ZN(n19285) );
  NAND2_X1 U20635 ( .A1(n19328), .A2(n19283), .ZN(n17420) );
  INV_X1 U20636 ( .A(n19488), .ZN(n19442) );
  OAI21_X1 U20637 ( .B1(n19285), .B2(n17420), .A(n19442), .ZN(n17435) );
  OAI211_X1 U20638 ( .C1(n19488), .C2(n19264), .A(n17421), .B(n17435), .ZN(
        n19261) );
  AOI21_X1 U20639 ( .B1(n19282), .B2(n17422), .A(n19261), .ZN(n17423) );
  OAI211_X1 U20640 ( .C1(n17425), .C2(n10378), .A(n17424), .B(n17423), .ZN(
        n19251) );
  MUX2_X1 U20641 ( .A(n17426), .B(n19251), .S(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .Z(n17427) );
  NAND2_X1 U20642 ( .A1(n17427), .A2(n19457), .ZN(n17431) );
  INV_X1 U20643 ( .A(n17428), .ZN(n17429) );
  AOI21_X1 U20644 ( .B1(n19473), .B2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n17429), .ZN(n17430) );
  OAI211_X1 U20645 ( .C1(n17432), .C2(n19428), .A(n17431), .B(n17430), .ZN(
        P3_U2836) );
  INV_X1 U20646 ( .A(n18957), .ZN(n17433) );
  AOI21_X1 U20647 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n17434), .A(
        n17433), .ZN(n18972) );
  NOR2_X1 U20648 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n18988), .ZN(
        n18974) );
  NOR2_X1 U20649 ( .A1(n14191), .A2(n20114), .ZN(n18964) );
  INV_X1 U20650 ( .A(n19355), .ZN(n19447) );
  OAI211_X1 U20651 ( .C1(n18968), .C2(n10378), .A(n19512), .B(n17435), .ZN(
        n17436) );
  AOI21_X1 U20652 ( .B1(n19282), .B2(n18969), .A(n17436), .ZN(n17439) );
  NAND3_X1 U20653 ( .A1(n17437), .A2(n17439), .A3(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17438) );
  NAND2_X1 U20654 ( .A1(n17438), .A2(n14191), .ZN(n19277) );
  AOI211_X1 U20655 ( .C1(n19447), .C2(n17439), .A(n22186), .B(n19277), .ZN(
        n17440) );
  AOI211_X1 U20656 ( .C1(n18974), .C2(n17441), .A(n18964), .B(n17440), .ZN(
        n17442) );
  OAI21_X1 U20657 ( .B1(n18972), .B2(n19428), .A(n17442), .ZN(P3_U2838) );
  NOR2_X1 U20658 ( .A1(n17443), .A2(n19320), .ZN(n17448) );
  NOR2_X1 U20659 ( .A1(n17443), .A2(n22165), .ZN(n17445) );
  NAND2_X1 U20660 ( .A1(n19986), .A2(n22165), .ZN(n19489) );
  AOI21_X1 U20661 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n19489), .A(
        n19488), .ZN(n17444) );
  AOI21_X1 U20662 ( .B1(n17445), .B2(n19444), .A(n17444), .ZN(n17446) );
  INV_X1 U20663 ( .A(n17446), .ZN(n17447) );
  MUX2_X1 U20664 ( .A(n17448), .B(n17447), .S(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .Z(n17449) );
  NOR2_X1 U20665 ( .A1(n20019), .A2(n19322), .ZN(n19492) );
  OAI21_X1 U20666 ( .B1(n17449), .B2(n19492), .A(n19457), .ZN(n17457) );
  OR2_X1 U20667 ( .A1(n19505), .A2(n17450), .ZN(n17455) );
  OAI22_X1 U20668 ( .A1(n17452), .A2(n19512), .B1(n10011), .B2(n17451), .ZN(
        n17453) );
  INV_X1 U20669 ( .A(n17453), .ZN(n17454) );
  NAND4_X1 U20670 ( .A1(n17457), .A2(n17456), .A3(n17455), .A4(n17454), .ZN(
        P3_U2860) );
  MUX2_X1 U20671 ( .A(n17458), .B(n19349), .S(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n20003) );
  AOI22_X1 U20672 ( .A1(n20151), .A2(n17459), .B1(P3_STATE2_REG_1__SCAN_IN), 
        .B2(n22165), .ZN(n17460) );
  OAI21_X1 U20673 ( .B1(n20003), .B2(n20140), .A(n17460), .ZN(n17461) );
  MUX2_X1 U20674 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(n17461), .S(
        n20155), .Z(P3_U3290) );
  NAND3_X1 U20675 ( .A1(n17462), .A2(P3_EBX_REG_6__SCAN_IN), .A3(
        P3_EBX_REG_5__SCAN_IN), .ZN(n18582) );
  INV_X1 U20676 ( .A(P3_EBX_REG_12__SCAN_IN), .ZN(n18561) );
  NAND3_X1 U20678 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(P3_EBX_REG_13__SCAN_IN), 
        .A3(n17574), .ZN(n18521) );
  NAND2_X1 U20679 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n18520), .ZN(n18504) );
  INV_X1 U20680 ( .A(n18461), .ZN(n18481) );
  AND2_X1 U20681 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .ZN(n18339) );
  NOR3_X1 U20682 ( .A1(n18338), .A2(n18002), .A3(n18389), .ZN(n17463) );
  NAND4_X1 U20683 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n17558), .A3(n18339), 
        .A4(n17463), .ZN(n18303) );
  NOR2_X1 U20684 ( .A1(n18304), .A2(n18303), .ZN(n18333) );
  NAND2_X1 U20685 ( .A1(n18661), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n17465) );
  NAND2_X1 U20686 ( .A1(n18333), .A2(n19561), .ZN(n17464) );
  OAI22_X1 U20687 ( .A1(n18333), .A2(n17465), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n17464), .ZN(P3_U2672) );
  OAI22_X1 U20688 ( .A1(n18466), .A2(n18454), .B1(n9786), .B2(n22105), .ZN(
        n17470) );
  AOI22_X1 U20689 ( .A1(n9724), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n14232), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17467) );
  NAND2_X1 U20690 ( .A1(n17547), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n17466) );
  OAI211_X1 U20691 ( .C1(n17468), .C2(n9723), .A(n17467), .B(n17466), .ZN(
        n17469) );
  AOI211_X1 U20692 ( .C1(n11937), .C2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A(
        n17470), .B(n17469), .ZN(n17472) );
  AOI22_X1 U20693 ( .A1(n18586), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n18403), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17471) );
  OAI211_X1 U20694 ( .C1(n9718), .C2(n18447), .A(n17472), .B(n17471), .ZN(
        n17477) );
  AOI22_X1 U20695 ( .A1(n18628), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n9726), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17475) );
  AOI22_X1 U20696 ( .A1(n18585), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11911), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17474) );
  AOI22_X1 U20697 ( .A1(n18626), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n18390), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17473) );
  NAND3_X1 U20698 ( .A1(n17475), .A2(n17474), .A3(n17473), .ZN(n17476) );
  NOR2_X1 U20699 ( .A1(n17477), .A2(n17476), .ZN(n18354) );
  INV_X1 U20700 ( .A(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n18486) );
  OAI22_X1 U20701 ( .A1(n18611), .A2(n18486), .B1(n17478), .B2(n18613), .ZN(
        n17486) );
  INV_X1 U20702 ( .A(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n18485) );
  INV_X1 U20703 ( .A(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17480) );
  OAI22_X1 U20704 ( .A1(n18616), .A2(n17480), .B1(n9723), .B2(n17479), .ZN(
        n17482) );
  NOR2_X1 U20705 ( .A1(n11861), .A2(n18623), .ZN(n17481) );
  AOI211_X1 U20706 ( .C1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .C2(n14232), .A(
        n17482), .B(n17481), .ZN(n17484) );
  AOI22_X1 U20707 ( .A1(n18620), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n18619), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17483) );
  OAI211_X1 U20708 ( .C1(n17550), .C2(n18485), .A(n17484), .B(n17483), .ZN(
        n17485) );
  AOI211_X1 U20709 ( .C1(n18591), .C2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A(
        n17486), .B(n17485), .ZN(n17490) );
  AOI22_X1 U20710 ( .A1(n18626), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n18403), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17489) );
  AOI22_X1 U20711 ( .A1(n18390), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n9724), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17488) );
  AOI22_X1 U20712 ( .A1(n18628), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n9726), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17487) );
  AND4_X1 U20713 ( .A1(n17490), .A2(n17489), .A3(n17488), .A4(n17487), .ZN(
        n18365) );
  OAI22_X1 U20714 ( .A1(n18611), .A2(n11841), .B1(n19777), .B2(n18615), .ZN(
        n17497) );
  AOI22_X1 U20715 ( .A1(n17547), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n18597), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n17495) );
  AOI22_X1 U20716 ( .A1(n18620), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n18619), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n17494) );
  AOI22_X1 U20717 ( .A1(n9724), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17561), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n17493) );
  INV_X1 U20718 ( .A(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n17491) );
  OR2_X1 U20719 ( .A1(n17550), .A2(n17491), .ZN(n17492) );
  NAND4_X1 U20720 ( .A1(n17495), .A2(n17494), .A3(n17493), .A4(n17492), .ZN(
        n17496) );
  AOI211_X1 U20721 ( .C1(n18591), .C2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A(
        n17497), .B(n17496), .ZN(n17501) );
  AOI22_X1 U20722 ( .A1(n18390), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11911), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17500) );
  AOI22_X1 U20723 ( .A1(n18585), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n18403), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n17499) );
  AOI22_X1 U20724 ( .A1(n18628), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n9726), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n17498) );
  AND4_X1 U20725 ( .A1(n17501), .A2(n17500), .A3(n17499), .A4(n17498), .ZN(
        n18364) );
  NOR2_X1 U20726 ( .A1(n18365), .A2(n18364), .ZN(n18361) );
  INV_X1 U20727 ( .A(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n18474) );
  NOR2_X1 U20728 ( .A1(n18616), .A2(n18474), .ZN(n17504) );
  INV_X1 U20729 ( .A(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n18598) );
  OAI22_X1 U20730 ( .A1(n18613), .A2(n18598), .B1(n9723), .B2(n17502), .ZN(
        n17503) );
  AOI211_X1 U20731 ( .C1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .C2(n9724), .A(
        n17504), .B(n17503), .ZN(n17506) );
  AOI22_X1 U20732 ( .A1(n18620), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n18619), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n17505) );
  OAI211_X1 U20733 ( .C1(n17550), .C2(n17507), .A(n17506), .B(n17505), .ZN(
        n17510) );
  AOI22_X1 U20734 ( .A1(n18586), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n18390), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n17508) );
  OAI21_X1 U20735 ( .B1(n9718), .B2(n11951), .A(n17508), .ZN(n17509) );
  NOR2_X1 U20736 ( .A1(n17510), .A2(n17509), .ZN(n17514) );
  AOI22_X1 U20737 ( .A1(n11911), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n14232), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n17513) );
  AOI22_X1 U20738 ( .A1(n18626), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n18403), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17512) );
  AOI22_X1 U20739 ( .A1(n18628), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n9726), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n17511) );
  NAND4_X1 U20740 ( .A1(n17514), .A2(n17513), .A3(n17512), .A4(n17511), .ZN(
        n18360) );
  NAND2_X1 U20741 ( .A1(n18361), .A2(n18360), .ZN(n18359) );
  NOR2_X1 U20742 ( .A1(n18354), .A2(n18359), .ZN(n18353) );
  INV_X1 U20743 ( .A(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n18572) );
  NOR2_X1 U20744 ( .A1(n18616), .A2(n18574), .ZN(n17517) );
  INV_X1 U20745 ( .A(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n18573) );
  OAI22_X1 U20746 ( .A1(n18613), .A2(n18573), .B1(n9723), .B2(n17515), .ZN(
        n17516) );
  AOI211_X1 U20747 ( .C1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .C2(n9724), .A(
        n17517), .B(n17516), .ZN(n17519) );
  AOI22_X1 U20748 ( .A1(n18620), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n18619), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17518) );
  OAI211_X1 U20749 ( .C1(n17550), .C2(n18572), .A(n17519), .B(n17518), .ZN(
        n17522) );
  AOI22_X1 U20750 ( .A1(n18586), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n18390), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17520) );
  OAI21_X1 U20751 ( .B1(n9718), .B2(n18431), .A(n17520), .ZN(n17521) );
  NOR2_X1 U20752 ( .A1(n17522), .A2(n17521), .ZN(n17526) );
  AOI22_X1 U20753 ( .A1(n11911), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n14232), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17525) );
  AOI22_X1 U20754 ( .A1(n18626), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n18403), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17524) );
  AOI22_X1 U20755 ( .A1(n18628), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n9726), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17523) );
  NAND4_X1 U20756 ( .A1(n17526), .A2(n17525), .A3(n17524), .A4(n17523), .ZN(
        n18349) );
  NAND2_X1 U20757 ( .A1(n18353), .A2(n18349), .ZN(n18348) );
  INV_X1 U20758 ( .A(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n18553) );
  NAND2_X1 U20759 ( .A1(n9724), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n17527) );
  OAI21_X1 U20760 ( .B1(n18553), .B2(n18616), .A(n17527), .ZN(n17529) );
  INV_X1 U20761 ( .A(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n18552) );
  OAI22_X1 U20762 ( .A1(n18613), .A2(n18552), .B1(n9723), .B2(n18420), .ZN(
        n17528) );
  NOR2_X1 U20763 ( .A1(n17529), .A2(n17528), .ZN(n17536) );
  AOI22_X1 U20764 ( .A1(n18586), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n18403), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17535) );
  INV_X1 U20765 ( .A(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n18550) );
  INV_X1 U20766 ( .A(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n19667) );
  NAND2_X1 U20767 ( .A1(n18620), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n17531) );
  NAND2_X1 U20768 ( .A1(n18489), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n17530) );
  OAI211_X1 U20769 ( .C1(n17550), .C2(n18550), .A(n17531), .B(n17530), .ZN(
        n17532) );
  INV_X1 U20770 ( .A(n17532), .ZN(n17534) );
  NAND2_X1 U20771 ( .A1(n18591), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n17533) );
  NAND4_X1 U20772 ( .A1(n17536), .A2(n17535), .A3(n17534), .A4(n17533), .ZN(
        n17541) );
  AOI22_X1 U20773 ( .A1(n18628), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n9726), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17539) );
  AOI22_X1 U20774 ( .A1(n11911), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n14232), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17538) );
  AOI22_X1 U20775 ( .A1(n18626), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n18390), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n17537) );
  NAND3_X1 U20776 ( .A1(n17539), .A2(n17538), .A3(n17537), .ZN(n17540) );
  NOR2_X1 U20777 ( .A1(n17541), .A2(n17540), .ZN(n18343) );
  NOR2_X1 U20778 ( .A1(n18348), .A2(n18343), .ZN(n18342) );
  INV_X1 U20779 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n18645) );
  OAI22_X1 U20780 ( .A1(n18611), .A2(n18396), .B1(n10660), .B2(n18645), .ZN(
        n17552) );
  INV_X1 U20781 ( .A(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n17543) );
  OAI22_X1 U20782 ( .A1(n18613), .A2(n17543), .B1(n9723), .B2(n17542), .ZN(
        n17546) );
  INV_X1 U20783 ( .A(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n17544) );
  NOR2_X1 U20784 ( .A1(n18556), .A2(n17544), .ZN(n17545) );
  AOI211_X1 U20785 ( .C1(n17547), .C2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A(
        n17546), .B(n17545), .ZN(n17549) );
  AOI22_X1 U20786 ( .A1(n18620), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n18489), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n17548) );
  OAI211_X1 U20787 ( .C1(n17550), .C2(n18393), .A(n17549), .B(n17548), .ZN(
        n17551) );
  AOI211_X1 U20788 ( .C1(n18591), .C2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A(
        n17552), .B(n17551), .ZN(n17556) );
  AOI22_X1 U20789 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n11911), .B1(
        n14232), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n17555) );
  AOI22_X1 U20790 ( .A1(n18626), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n18390), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n17554) );
  AOI22_X1 U20791 ( .A1(n18628), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n9726), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n17553) );
  NAND4_X1 U20792 ( .A1(n17556), .A2(n17555), .A3(n17554), .A4(n17553), .ZN(
        n17557) );
  NAND2_X1 U20793 ( .A1(n18342), .A2(n17557), .ZN(n18335) );
  OAI21_X1 U20794 ( .B1(n18342), .B2(n17557), .A(n18335), .ZN(n18694) );
  NAND2_X1 U20795 ( .A1(n19561), .A2(n18670), .ZN(n18664) );
  NAND3_X1 U20796 ( .A1(n19561), .A2(P3_EBX_REG_21__SCAN_IN), .A3(n17558), 
        .ZN(n18352) );
  NAND2_X1 U20797 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n18357), .ZN(n18347) );
  NAND2_X1 U20798 ( .A1(n18661), .A2(n18347), .ZN(n18345) );
  OAI21_X1 U20799 ( .B1(n18339), .B2(n18664), .A(n18345), .ZN(n18337) );
  NOR3_X1 U20800 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n18346), .A3(n18347), .ZN(
        n17559) );
  AOI21_X1 U20801 ( .B1(P3_EBX_REG_28__SCAN_IN), .B2(n18337), .A(n17559), .ZN(
        n17560) );
  OAI21_X1 U20802 ( .B1(n18694), .B2(n18661), .A(n17560), .ZN(P3_U2675) );
  AOI22_X1 U20803 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n17547), .B1(
        n9724), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n17566) );
  AOI22_X1 U20804 ( .A1(n18585), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17561), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n17565) );
  AOI22_X1 U20805 ( .A1(n18620), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n18619), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n17564) );
  INV_X1 U20806 ( .A(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n17562) );
  OR2_X1 U20807 ( .A1(n17550), .A2(n17562), .ZN(n17563) );
  AND4_X1 U20808 ( .A1(n17566), .A2(n17565), .A3(n17564), .A4(n17563), .ZN(
        n17568) );
  AOI22_X1 U20809 ( .A1(n18586), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n18597), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n17567) );
  OAI211_X1 U20810 ( .C1(n18645), .C2(n9718), .A(n17568), .B(n17567), .ZN(
        n17573) );
  INV_X1 U20811 ( .A(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n17569) );
  OAI22_X1 U20812 ( .A1(n18525), .A2(n18393), .B1(n17569), .B2(n18615), .ZN(
        n17572) );
  OAI22_X1 U20813 ( .A1(n9783), .A2(n18391), .B1(n17543), .B2(n18599), .ZN(
        n17571) );
  OAI22_X1 U20814 ( .A1(n10660), .A2(n18396), .B1(n11861), .B2(n18395), .ZN(
        n17570) );
  NOR4_X1 U20815 ( .A1(n17573), .A2(n17572), .A3(n17571), .A4(n17570), .ZN(
        n18770) );
  OAI22_X1 U20816 ( .A1(n18667), .A2(n17574), .B1(P3_EBX_REG_13__SCAN_IN), 
        .B2(n18664), .ZN(n18540) );
  OAI21_X1 U20817 ( .B1(P3_EBX_REG_13__SCAN_IN), .B2(n17574), .A(n18540), .ZN(
        n17575) );
  OAI21_X1 U20818 ( .B1(n18770), .B2(n18661), .A(n17575), .ZN(P3_U2690) );
  NOR2_X1 U20819 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20138), .ZN(
        n19566) );
  NOR2_X1 U20820 ( .A1(n17576), .A2(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n17585) );
  NAND2_X1 U20821 ( .A1(n18599), .A2(n17585), .ZN(n19522) );
  INV_X1 U20822 ( .A(n19565), .ZN(n19833) );
  AOI211_X1 U20823 ( .C1(n17578), .C2(n19522), .A(n19833), .B(n17577), .ZN(
        n17579) );
  NOR2_X1 U20824 ( .A1(n19566), .A2(n17579), .ZN(n17581) );
  INV_X1 U20825 ( .A(n17579), .ZN(n19528) );
  OAI22_X1 U20826 ( .A1(n19067), .A2(n20178), .B1(n11982), .B2(n20138), .ZN(
        n17584) );
  NAND3_X1 U20827 ( .A1(n20002), .A2(n19528), .A3(n17584), .ZN(n17580) );
  OAI221_X1 U20828 ( .B1(n20002), .B2(n17581), .C1(n20002), .C2(n19830), .A(
        n17580), .ZN(P3_U2864) );
  OR2_X1 U20829 ( .A1(n19067), .A2(n20178), .ZN(n17582) );
  OAI221_X1 U20830 ( .B1(n20138), .B2(n19681), .C1(n17582), .C2(n19681), .A(
        n17581), .ZN(n17583) );
  INV_X1 U20831 ( .A(n17583), .ZN(n19527) );
  INV_X1 U20832 ( .A(n19830), .ZN(n19707) );
  OAI221_X1 U20833 ( .B1(n19707), .B2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .C1(n19707), .C2(n17584), .A(n19528), .ZN(n19525) );
  AOI22_X1 U20834 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n19527), .B1(
        n19525), .B2(n20011), .ZN(P3_U2865) );
  NOR2_X1 U20835 ( .A1(n17585), .A2(n20013), .ZN(n20024) );
  NAND3_X1 U20836 ( .A1(n20155), .A2(n20188), .A3(n20024), .ZN(n17586) );
  OAI21_X1 U20837 ( .B1(n20155), .B2(n18236), .A(n17586), .ZN(P3_U3284) );
  OAI21_X1 U20838 ( .B1(n17824), .B2(n10378), .A(n17587), .ZN(n17588) );
  OAI221_X1 U20839 ( .B1(n17588), .B2(n17820), .C1(n17588), .C2(n19282), .A(
        n19457), .ZN(n17635) );
  AOI211_X1 U20840 ( .C1(n19355), .C2(n21976), .A(n19517), .B(n17589), .ZN(
        n17591) );
  NOR3_X1 U20841 ( .A1(n17808), .A2(n19188), .A3(n19505), .ZN(n17590) );
  AOI21_X1 U20842 ( .B1(n19388), .B2(n17809), .A(n17590), .ZN(n17638) );
  OAI21_X1 U20843 ( .B1(n19508), .B2(n17591), .A(n17638), .ZN(n17595) );
  NAND2_X1 U20844 ( .A1(n17593), .A2(n17592), .ZN(n17594) );
  XOR2_X1 U20845 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B(n17594), .Z(
        n17828) );
  AOI22_X1 U20846 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n17595), .B1(
        n19455), .B2(n17828), .ZN(n17596) );
  NAND2_X1 U20847 ( .A1(n19508), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n17831) );
  OAI211_X1 U20848 ( .C1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n17635), .A(
        n17596), .B(n17831), .ZN(P3_U2833) );
  NOR3_X1 U20849 ( .A1(n17598), .A2(n17597), .A3(n21729), .ZN(n17601) );
  NAND2_X1 U20850 ( .A1(n17601), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n17603) );
  OAI22_X1 U20851 ( .A1(n17601), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(
        n17600), .B2(n17599), .ZN(n17602) );
  NAND2_X1 U20852 ( .A1(n17603), .A2(n17602), .ZN(n17606) );
  INV_X1 U20853 ( .A(n17604), .ZN(n17605) );
  AOI222_X1 U20854 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n17606), 
        .B1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n17605), .C1(n17606), 
        .C2(n17605), .ZN(n17608) );
  AOI222_X1 U20855 ( .A1(n17608), .A2(n21636), .B1(n17608), .B2(n17607), .C1(
        n21636), .C2(n17607), .ZN(n17618) );
  INV_X1 U20856 ( .A(n17609), .ZN(n17614) );
  INV_X1 U20857 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n17611) );
  AOI21_X1 U20858 ( .B1(n22052), .B2(n17611), .A(n17610), .ZN(n17613) );
  NOR4_X1 U20859 ( .A1(n17615), .A2(n17614), .A3(n17613), .A4(n17612), .ZN(
        n17617) );
  OAI211_X1 U20860 ( .C1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .C2(n17618), .A(
        n17617), .B(n17616), .ZN(n17626) );
  AOI21_X1 U20861 ( .B1(n17625), .B2(n17626), .A(n17619), .ZN(n17620) );
  OAI211_X1 U20862 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n21912), .A(n17620), 
        .B(n17628), .ZN(n17627) );
  NOR3_X1 U20863 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n12682), .A3(n21912), 
        .ZN(n17624) );
  NAND3_X1 U20864 ( .A1(n13490), .A2(n12289), .A3(n17621), .ZN(n17623) );
  OAI22_X1 U20865 ( .A1(n17625), .A2(n17624), .B1(n17623), .B2(n17622), .ZN(
        n17709) );
  AOI221_X1 U20866 ( .B1(n21908), .B2(n21871), .C1(n17626), .C2(n21871), .A(
        n17709), .ZN(n17706) );
  NOR2_X1 U20867 ( .A1(n17627), .A2(n17706), .ZN(n17631) );
  OAI21_X1 U20868 ( .B1(n17629), .B2(n17628), .A(n21908), .ZN(n17630) );
  OAI22_X1 U20869 ( .A1(n21908), .A2(n17631), .B1(n17706), .B2(n17630), .ZN(
        P1_U3161) );
  NOR2_X1 U20870 ( .A1(n17633), .A2(n17632), .ZN(n17634) );
  XNOR2_X1 U20871 ( .A(n17634), .B(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n17816) );
  NOR2_X1 U20872 ( .A1(n14191), .A2(n20129), .ZN(n17811) );
  NOR3_X1 U20873 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n17825), .A3(
        n17635), .ZN(n17636) );
  AOI211_X1 U20874 ( .C1(n19455), .C2(n17816), .A(n17811), .B(n17636), .ZN(
        n17637) );
  OAI221_X1 U20875 ( .B1(n17817), .B2(n17639), .C1(n17817), .C2(n17638), .A(
        n17637), .ZN(P3_U2832) );
  INV_X1 U20876 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n17912) );
  NOR2_X1 U20877 ( .A1(n21285), .A2(n17912), .ZN(P1_U2905) );
  NOR2_X1 U20878 ( .A1(n21133), .A2(n21003), .ZN(n17791) );
  NOR4_X1 U20879 ( .A1(n17641), .A2(n21135), .A3(n17640), .A4(n17791), .ZN(
        P2_U3178) );
  INV_X1 U20880 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n17765) );
  NOR2_X1 U20881 ( .A1(n17765), .A2(n21112), .ZN(P2_U3047) );
  AOI22_X1 U20882 ( .A1(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n21233), .B1(
        n17642), .B2(n21174), .ZN(n17655) );
  NAND2_X1 U20883 ( .A1(n21251), .A2(n17643), .ZN(n21177) );
  OAI21_X1 U20884 ( .B1(n21177), .B2(n21878), .A(n17644), .ZN(n17652) );
  OAI22_X1 U20885 ( .A1(n17647), .A2(n17646), .B1(n17645), .B2(n21256), .ZN(
        n17651) );
  NOR2_X1 U20886 ( .A1(n17649), .A2(n17648), .ZN(n17650) );
  AOI211_X1 U20887 ( .C1(n17653), .C2(n17652), .A(n17651), .B(n17650), .ZN(
        n17654) );
  NAND3_X1 U20888 ( .A1(n17655), .A2(n17654), .A3(n21235), .ZN(P1_U2830) );
  AOI22_X1 U20889 ( .A1(n17661), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n17697), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n17660) );
  AOI21_X1 U20890 ( .B1(n17658), .B2(n17657), .A(n17656), .ZN(n17692) );
  AOI22_X1 U20891 ( .A1(n17692), .A2(n12669), .B1(n21328), .B2(n21200), .ZN(
        n17659) );
  OAI211_X1 U20892 ( .C1(n17670), .C2(n21196), .A(n17660), .B(n17659), .ZN(
        P1_U2992) );
  AOI22_X1 U20893 ( .A1(n17661), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n17697), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n17669) );
  INV_X1 U20894 ( .A(n17663), .ZN(n17665) );
  NAND2_X1 U20895 ( .A1(n17665), .A2(n17664), .ZN(n17666) );
  XNOR2_X1 U20896 ( .A(n17662), .B(n17666), .ZN(n17701) );
  INV_X1 U20897 ( .A(n17667), .ZN(n21211) );
  AOI22_X1 U20898 ( .A1(n17701), .A2(n12669), .B1(n21211), .B2(n21328), .ZN(
        n17668) );
  OAI211_X1 U20899 ( .C1(n17670), .C2(n21206), .A(n17669), .B(n17668), .ZN(
        P1_U2993) );
  OAI22_X1 U20900 ( .A1(n21226), .A2(n17671), .B1(n21218), .B2(n17670), .ZN(
        n17672) );
  AOI21_X1 U20901 ( .B1(n17673), .B2(n12669), .A(n17672), .ZN(n17675) );
  OAI211_X1 U20902 ( .C1(n17677), .C2(n17676), .A(n17675), .B(n17674), .ZN(
        P1_U2994) );
  NAND2_X1 U20903 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n17699), .ZN(
        n17695) );
  NAND2_X1 U20904 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n17678) );
  OAI21_X1 U20905 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n17678), .ZN(n17690) );
  INV_X1 U20906 ( .A(n17679), .ZN(n21183) );
  AOI21_X1 U20907 ( .B1(n17698), .B2(n21183), .A(n17680), .ZN(n17689) );
  INV_X1 U20908 ( .A(n17681), .ZN(n17686) );
  INV_X1 U20909 ( .A(n17682), .ZN(n17683) );
  AOI21_X1 U20910 ( .B1(n17685), .B2(n17684), .A(n17683), .ZN(n17705) );
  OAI21_X1 U20911 ( .B1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n17686), .A(
        n17705), .ZN(n17691) );
  AOI22_X1 U20912 ( .A1(n17687), .A2(n17700), .B1(
        P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n17691), .ZN(n17688) );
  OAI211_X1 U20913 ( .C1(n17695), .C2(n17690), .A(n17689), .B(n17688), .ZN(
        P1_U3023) );
  AOI22_X1 U20914 ( .A1(n17698), .A2(n21199), .B1(n17697), .B2(
        P1_REIP_REG_7__SCAN_IN), .ZN(n17694) );
  AOI22_X1 U20915 ( .A1(n17692), .A2(n17700), .B1(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n17691), .ZN(n17693) );
  OAI211_X1 U20916 ( .C1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n17695), .A(
        n17694), .B(n17693), .ZN(P1_U3024) );
  INV_X1 U20917 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n17704) );
  INV_X1 U20918 ( .A(n17696), .ZN(n21205) );
  AOI22_X1 U20919 ( .A1(n17698), .A2(n21205), .B1(n17697), .B2(
        P1_REIP_REG_6__SCAN_IN), .ZN(n17703) );
  AOI22_X1 U20920 ( .A1(n17701), .A2(n17700), .B1(n17699), .B2(n17704), .ZN(
        n17702) );
  OAI211_X1 U20921 ( .C1(n17705), .C2(n17704), .A(n17703), .B(n17702), .ZN(
        P1_U3025) );
  NOR2_X1 U20922 ( .A1(n17706), .A2(n21908), .ZN(n17716) );
  NAND4_X1 U20923 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .A3(n12682), .A4(n21912), .ZN(n17707) );
  NAND2_X1 U20924 ( .A1(n17708), .A2(n17707), .ZN(n21872) );
  OAI21_X1 U20925 ( .B1(n17710), .B2(n21872), .A(n17709), .ZN(n17711) );
  OAI21_X1 U20926 ( .B1(P1_STATE2_REG_1__SCAN_IN), .B2(n17716), .A(n17711), 
        .ZN(n17712) );
  AOI221_X1 U20927 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n17714), .C1(n17713), 
        .C2(n17714), .A(n17712), .ZN(P1_U3162) );
  OAI21_X1 U20928 ( .B1(n17716), .B2(n21704), .A(n17715), .ZN(P1_U3466) );
  AOI22_X1 U20929 ( .A1(n17725), .A2(n17717), .B1(P2_REIP_REG_5__SCAN_IN), 
        .B2(n20355), .ZN(n17722) );
  AOI222_X1 U20930 ( .A1(n17720), .A2(n20357), .B1(n11457), .B2(n17719), .C1(
        n20370), .C2(n17718), .ZN(n17721) );
  OAI211_X1 U20931 ( .C1(n17736), .C2(n17723), .A(n17722), .B(n17721), .ZN(
        P2_U3009) );
  NOR2_X1 U20932 ( .A1(n20217), .A2(n21035), .ZN(n17740) );
  AOI21_X1 U20933 ( .B1(n17725), .B2(n17724), .A(n17740), .ZN(n17735) );
  NAND2_X1 U20934 ( .A1(n17727), .A2(n17726), .ZN(n17729) );
  XNOR2_X1 U20935 ( .A(n17729), .B(n17728), .ZN(n17747) );
  INV_X1 U20936 ( .A(n17730), .ZN(n17731) );
  AOI21_X1 U20937 ( .B1(n17732), .B2(n11315), .A(n17731), .ZN(n17739) );
  AOI222_X1 U20938 ( .A1(n17747), .A2(n11457), .B1(n20357), .B2(n17739), .C1(
        n17733), .C2(n20370), .ZN(n17734) );
  OAI211_X1 U20939 ( .C1(n17737), .C2(n17736), .A(n17735), .B(n17734), .ZN(
        P2_U3011) );
  NAND2_X1 U20940 ( .A1(n17739), .A2(n17738), .ZN(n17743) );
  AOI21_X1 U20941 ( .B1(n17741), .B2(n20288), .A(n17740), .ZN(n17742) );
  OAI211_X1 U20942 ( .C1(n17745), .C2(n17744), .A(n17743), .B(n17742), .ZN(
        n17746) );
  AOI21_X1 U20943 ( .B1(n17748), .B2(n17747), .A(n17746), .ZN(n17749) );
  OAI221_X1 U20944 ( .B1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n17752), .C1(
        n17751), .C2(n17750), .A(n17749), .ZN(P2_U3043) );
  MUX2_X1 U20945 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n17753), .S(
        n17771), .Z(n17787) );
  OAI21_X1 U20946 ( .B1(n17755), .B2(n21114), .A(n17754), .ZN(n17757) );
  OAI21_X1 U20947 ( .B1(n17755), .B2(n20837), .A(n17771), .ZN(n17756) );
  AOI21_X1 U20948 ( .B1(n17758), .B2(n17757), .A(n17756), .ZN(n17760) );
  OR2_X1 U20949 ( .A1(n17761), .A2(n22183), .ZN(n17759) );
  OAI211_X1 U20950 ( .C1(n17787), .C2(n21096), .A(n17760), .B(n17759), .ZN(
        n17764) );
  MUX2_X1 U20951 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n17761), .S(
        n17771), .Z(n17788) );
  NAND2_X1 U20952 ( .A1(n21096), .A2(n22183), .ZN(n20483) );
  INV_X1 U20953 ( .A(n20483), .ZN(n20508) );
  NAND2_X1 U20954 ( .A1(n17788), .A2(n20508), .ZN(n17763) );
  NAND2_X1 U20955 ( .A1(n17787), .A2(n21096), .ZN(n17762) );
  NAND3_X1 U20956 ( .A1(n17764), .A2(n17763), .A3(n17762), .ZN(n17766) );
  NAND2_X1 U20957 ( .A1(n17766), .A2(n17765), .ZN(n17790) );
  NOR2_X1 U20958 ( .A1(n21118), .A2(n17767), .ZN(n17769) );
  OAI211_X1 U20959 ( .C1(n17771), .C2(n17770), .A(n17769), .B(n17768), .ZN(
        n17772) );
  INV_X1 U20960 ( .A(n17772), .ZN(n17785) );
  OAI21_X1 U20961 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(P2_MORE_REG_SCAN_IN), .A(
        n17773), .ZN(n17784) );
  MUX2_X1 U20962 ( .A(n17776), .B(n17775), .S(n17774), .Z(n17783) );
  INV_X1 U20963 ( .A(n17777), .ZN(n17780) );
  OAI22_X1 U20964 ( .A1(n17781), .A2(n17780), .B1(n17779), .B2(n17778), .ZN(
        n17782) );
  NOR2_X1 U20965 ( .A1(n17783), .A2(n17782), .ZN(n21121) );
  NAND3_X1 U20966 ( .A1(n17785), .A2(n17784), .A3(n21121), .ZN(n17786) );
  AOI21_X1 U20967 ( .B1(n17788), .B2(n17787), .A(n17786), .ZN(n17789) );
  NAND2_X1 U20968 ( .A1(n17790), .A2(n17789), .ZN(n17799) );
  AOI211_X1 U20969 ( .C1(n17793), .C2(n17799), .A(n17792), .B(n17791), .ZN(
        n17805) );
  INV_X1 U20970 ( .A(n21133), .ZN(n21126) );
  OR2_X1 U20971 ( .A1(n17795), .A2(n17794), .ZN(n17797) );
  AND2_X1 U20972 ( .A1(n17797), .A2(n10671), .ZN(n17800) );
  AOI22_X1 U20973 ( .A1(n17798), .A2(n21135), .B1(n21126), .B2(n17800), .ZN(
        n17803) );
  OAI21_X1 U20974 ( .B1(n17799), .B2(P2_STATE2_REG_1__SCAN_IN), .A(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n17801) );
  NAND2_X1 U20975 ( .A1(n17801), .A2(n17800), .ZN(n21002) );
  AND2_X1 U20976 ( .A1(n21002), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n17807) );
  INV_X1 U20977 ( .A(n17807), .ZN(n17802) );
  OAI21_X1 U20978 ( .B1(P2_STATE2_REG_0__SCAN_IN), .B2(n17803), .A(n17802), 
        .ZN(n17804) );
  OAI211_X1 U20979 ( .C1(n21119), .C2(n17806), .A(n17805), .B(n17804), .ZN(
        P2_U3176) );
  OAI21_X1 U20980 ( .B1(n17807), .B2(n21106), .A(n17806), .ZN(P2_U3593) );
  OR2_X1 U20981 ( .A1(n19105), .A2(n17808), .ZN(n17821) );
  NAND2_X1 U20982 ( .A1(n10167), .A2(n17809), .ZN(n17823) );
  AOI21_X1 U20983 ( .B1(n19128), .B2(n17947), .A(n17811), .ZN(n17812) );
  OAI221_X1 U20984 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n17814), .C1(
        n17948), .C2(n17813), .A(n17812), .ZN(n17815) );
  AOI22_X1 U20985 ( .A1(n9895), .A2(n17819), .B1(
        P3_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n17818), .ZN(n17833) );
  INV_X1 U20986 ( .A(n17820), .ZN(n17822) );
  AOI21_X1 U20987 ( .B1(n17822), .B2(n17825), .A(n17821), .ZN(n17827) );
  AOI21_X1 U20988 ( .B1(n17825), .B2(n17824), .A(n17823), .ZN(n17826) );
  AOI211_X1 U20989 ( .C1(n19172), .C2(n17828), .A(n17827), .B(n17826), .ZN(
        n17832) );
  OAI21_X1 U20990 ( .B1(n17829), .B2(n19128), .A(n17955), .ZN(n17830) );
  NAND4_X1 U20991 ( .A1(n17833), .A2(n17832), .A3(n17831), .A4(n17830), .ZN(
        P3_U2801) );
  NOR3_X1 U20992 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(P3_BE_N_REG_0__SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .ZN(n17835) );
  NOR4_X1 U20993 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n17834) );
  NAND4_X1 U20994 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n17835), .A3(n17834), .A4(
        U215), .ZN(U213) );
  INV_X1 U20995 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n20312) );
  INV_X2 U20996 ( .A(U214), .ZN(n17879) );
  OAI222_X1 U20997 ( .A1(U212), .A2(n20312), .B1(n17878), .B2(n17837), .C1(
        U214), .C2(n17912), .ZN(U216) );
  AOI222_X1 U20998 ( .A1(n17879), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n17880), 
        .B2(BUF1_REG_30__SCAN_IN), .C1(n17876), .C2(P2_DATAO_REG_30__SCAN_IN), 
        .ZN(n17838) );
  INV_X1 U20999 ( .A(n17838), .ZN(U217) );
  AOI22_X1 U21000 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n17879), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n17876), .ZN(n17839) );
  OAI21_X1 U21001 ( .B1(n16401), .B2(n17878), .A(n17839), .ZN(U218) );
  INV_X1 U21002 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n17841) );
  AOI22_X1 U21003 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n17879), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n17876), .ZN(n17840) );
  OAI21_X1 U21004 ( .B1(n17841), .B2(n17878), .A(n17840), .ZN(U219) );
  AOI22_X1 U21005 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n17879), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n17876), .ZN(n17842) );
  OAI21_X1 U21006 ( .B1(n16413), .B2(n17878), .A(n17842), .ZN(U220) );
  AOI22_X1 U21007 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n17879), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n17876), .ZN(n17843) );
  OAI21_X1 U21008 ( .B1(n16421), .B2(n17878), .A(n17843), .ZN(U221) );
  AOI222_X1 U21009 ( .A1(n17876), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(n17880), 
        .B2(BUF1_REG_25__SCAN_IN), .C1(n17879), .C2(P1_DATAO_REG_25__SCAN_IN), 
        .ZN(n17844) );
  INV_X1 U21010 ( .A(n17844), .ZN(U222) );
  INV_X1 U21011 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n17846) );
  AOI22_X1 U21012 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n17879), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n17876), .ZN(n17845) );
  OAI21_X1 U21013 ( .B1(n17846), .B2(n17878), .A(n17845), .ZN(U223) );
  AOI22_X1 U21014 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n17879), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n17876), .ZN(n17847) );
  OAI21_X1 U21015 ( .B1(n16442), .B2(n17878), .A(n17847), .ZN(U224) );
  AOI22_X1 U21016 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n17879), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n17876), .ZN(n17848) );
  OAI21_X1 U21017 ( .B1(n16449), .B2(n17878), .A(n17848), .ZN(U225) );
  AOI22_X1 U21018 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n17880), .B1(
        P1_DATAO_REG_21__SCAN_IN), .B2(n17879), .ZN(n17849) );
  OAI21_X1 U21019 ( .B1(n13754), .B2(U212), .A(n17849), .ZN(U226) );
  AOI22_X1 U21020 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n17879), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n17876), .ZN(n17850) );
  OAI21_X1 U21021 ( .B1(n17851), .B2(n17878), .A(n17850), .ZN(U227) );
  AOI22_X1 U21022 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n17879), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n17876), .ZN(n17852) );
  OAI21_X1 U21023 ( .B1(n16469), .B2(n17878), .A(n17852), .ZN(U228) );
  INV_X1 U21024 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n17854) );
  AOI22_X1 U21025 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n17879), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n17876), .ZN(n17853) );
  OAI21_X1 U21026 ( .B1(n17854), .B2(n17878), .A(n17853), .ZN(U229) );
  AOI22_X1 U21027 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n17879), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n17876), .ZN(n17855) );
  OAI21_X1 U21028 ( .B1(n16479), .B2(n17878), .A(n17855), .ZN(U230) );
  INV_X1 U21029 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n17857) );
  AOI22_X1 U21030 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n17879), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n17876), .ZN(n17856) );
  OAI21_X1 U21031 ( .B1(n17857), .B2(n17878), .A(n17856), .ZN(U231) );
  INV_X1 U21032 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n17896) );
  AOI22_X1 U21033 ( .A1(BUF1_REG_15__SCAN_IN), .A2(n17880), .B1(
        P1_DATAO_REG_15__SCAN_IN), .B2(n17879), .ZN(n17858) );
  OAI21_X1 U21034 ( .B1(n17896), .B2(U212), .A(n17858), .ZN(U232) );
  INV_X1 U21035 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n17860) );
  AOI22_X1 U21036 ( .A1(BUF1_REG_14__SCAN_IN), .A2(n17880), .B1(
        P1_DATAO_REG_14__SCAN_IN), .B2(n17879), .ZN(n17859) );
  OAI21_X1 U21037 ( .B1(n17860), .B2(U212), .A(n17859), .ZN(U233) );
  INV_X1 U21038 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n17894) );
  AOI22_X1 U21039 ( .A1(BUF1_REG_13__SCAN_IN), .A2(n17880), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(n17879), .ZN(n17861) );
  OAI21_X1 U21040 ( .B1(n17894), .B2(U212), .A(n17861), .ZN(U234) );
  AOI22_X1 U21041 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n17879), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n17876), .ZN(n17862) );
  OAI21_X1 U21042 ( .B1(n22194), .B2(n17878), .A(n17862), .ZN(U235) );
  INV_X1 U21043 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n17892) );
  AOI22_X1 U21044 ( .A1(BUF1_REG_11__SCAN_IN), .A2(n17880), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n17879), .ZN(n17863) );
  OAI21_X1 U21045 ( .B1(n17892), .B2(U212), .A(n17863), .ZN(U236) );
  AOI22_X1 U21046 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n17879), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n17876), .ZN(n17864) );
  OAI21_X1 U21047 ( .B1(n17865), .B2(n17878), .A(n17864), .ZN(U237) );
  INV_X1 U21048 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n17890) );
  INV_X1 U21049 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n22210) );
  OAI222_X1 U21050 ( .A1(U212), .A2(n17890), .B1(n17878), .B2(n17866), .C1(
        U214), .C2(n22210), .ZN(U238) );
  INV_X1 U21051 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n17868) );
  AOI22_X1 U21052 ( .A1(BUF1_REG_8__SCAN_IN), .A2(n17880), .B1(
        P1_DATAO_REG_8__SCAN_IN), .B2(n17879), .ZN(n17867) );
  OAI21_X1 U21053 ( .B1(n17868), .B2(U212), .A(n17867), .ZN(U239) );
  INV_X1 U21054 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n17888) );
  AOI22_X1 U21055 ( .A1(BUF1_REG_7__SCAN_IN), .A2(n17880), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n17879), .ZN(n17869) );
  OAI21_X1 U21056 ( .B1(n17888), .B2(U212), .A(n17869), .ZN(U240) );
  AOI22_X1 U21057 ( .A1(P1_DATAO_REG_6__SCAN_IN), .A2(n17879), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n17876), .ZN(n17870) );
  OAI21_X1 U21058 ( .B1(n17871), .B2(n17878), .A(n17870), .ZN(U241) );
  INV_X1 U21059 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n17886) );
  AOI22_X1 U21060 ( .A1(BUF1_REG_5__SCAN_IN), .A2(n17880), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(n17879), .ZN(n17872) );
  OAI21_X1 U21061 ( .B1(n17886), .B2(U212), .A(n17872), .ZN(U242) );
  AOI22_X1 U21062 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n17879), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n17876), .ZN(n17873) );
  OAI21_X1 U21063 ( .B1(n13678), .B2(n17878), .A(n17873), .ZN(U243) );
  AOI22_X1 U21064 ( .A1(P1_DATAO_REG_3__SCAN_IN), .A2(n17879), .B1(
        P2_DATAO_REG_3__SCAN_IN), .B2(n17876), .ZN(n17874) );
  OAI21_X1 U21065 ( .B1(n15263), .B2(n17878), .A(n17874), .ZN(U244) );
  AOI22_X1 U21066 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n17879), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n17876), .ZN(n17875) );
  OAI21_X1 U21067 ( .B1(n13640), .B2(n17878), .A(n17875), .ZN(U245) );
  AOI22_X1 U21068 ( .A1(P1_DATAO_REG_1__SCAN_IN), .A2(n17879), .B1(
        P2_DATAO_REG_1__SCAN_IN), .B2(n17876), .ZN(n17877) );
  OAI21_X1 U21069 ( .B1(n13665), .B2(n17878), .A(n17877), .ZN(U246) );
  INV_X1 U21070 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n22173) );
  AOI22_X1 U21071 ( .A1(BUF1_REG_0__SCAN_IN), .A2(n17880), .B1(
        P1_DATAO_REG_0__SCAN_IN), .B2(n17879), .ZN(n17881) );
  OAI21_X1 U21072 ( .B1(n22173), .B2(U212), .A(n17881), .ZN(U247) );
  AOI22_X1 U21073 ( .A1(n17904), .A2(n22173), .B1(n22011), .B2(U215), .ZN(U251) );
  OAI22_X1 U21074 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n17904), .ZN(n17882) );
  INV_X1 U21075 ( .A(n17882), .ZN(U252) );
  OAI22_X1 U21076 ( .A1(U215), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n17904), .ZN(n17883) );
  INV_X1 U21077 ( .A(n17883), .ZN(U253) );
  OAI22_X1 U21078 ( .A1(U215), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n17904), .ZN(n17884) );
  INV_X1 U21079 ( .A(n17884), .ZN(U254) );
  OAI22_X1 U21080 ( .A1(U215), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n17904), .ZN(n17885) );
  INV_X1 U21081 ( .A(n17885), .ZN(U255) );
  INV_X1 U21082 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n19550) );
  AOI22_X1 U21083 ( .A1(n17904), .A2(n17886), .B1(n19550), .B2(U215), .ZN(U256) );
  OAI22_X1 U21084 ( .A1(U215), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n17904), .ZN(n17887) );
  INV_X1 U21085 ( .A(n17887), .ZN(U257) );
  INV_X1 U21086 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n19558) );
  AOI22_X1 U21087 ( .A1(n17904), .A2(n17888), .B1(n19558), .B2(U215), .ZN(U258) );
  OAI22_X1 U21088 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n17904), .ZN(n17889) );
  INV_X1 U21089 ( .A(n17889), .ZN(U259) );
  INV_X1 U21090 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n18795) );
  AOI22_X1 U21091 ( .A1(n17904), .A2(n17890), .B1(n18795), .B2(U215), .ZN(U260) );
  OAI22_X1 U21092 ( .A1(U215), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n17904), .ZN(n17891) );
  INV_X1 U21093 ( .A(n17891), .ZN(U261) );
  INV_X1 U21094 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n18782) );
  AOI22_X1 U21095 ( .A1(n17904), .A2(n17892), .B1(n18782), .B2(U215), .ZN(U262) );
  OAI22_X1 U21096 ( .A1(U215), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n17904), .ZN(n17893) );
  INV_X1 U21097 ( .A(n17893), .ZN(U263) );
  INV_X1 U21098 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n18773) );
  AOI22_X1 U21099 ( .A1(n17904), .A2(n17894), .B1(n18773), .B2(U215), .ZN(U264) );
  OAI22_X1 U21100 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n17904), .ZN(n17895) );
  INV_X1 U21101 ( .A(n17895), .ZN(U265) );
  INV_X1 U21102 ( .A(BUF2_REG_15__SCAN_IN), .ZN(n22198) );
  AOI22_X1 U21103 ( .A1(n17904), .A2(n17896), .B1(n22198), .B2(U215), .ZN(U266) );
  OAI22_X1 U21104 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n17904), .ZN(n17897) );
  INV_X1 U21105 ( .A(n17897), .ZN(U267) );
  OAI22_X1 U21106 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17904), .ZN(n17898) );
  INV_X1 U21107 ( .A(n17898), .ZN(U268) );
  OAI22_X1 U21108 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n17904), .ZN(n17899) );
  INV_X1 U21109 ( .A(n17899), .ZN(U269) );
  OAI22_X1 U21110 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n17904), .ZN(n17900) );
  INV_X1 U21111 ( .A(n17900), .ZN(U270) );
  OAI22_X1 U21112 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n17904), .ZN(n17901) );
  INV_X1 U21113 ( .A(n17901), .ZN(U271) );
  INV_X1 U21114 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n17902) );
  AOI22_X1 U21115 ( .A1(n17904), .A2(n13754), .B1(n17902), .B2(U215), .ZN(U272) );
  OAI22_X1 U21116 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n17904), .ZN(n17903) );
  INV_X1 U21117 ( .A(n17903), .ZN(U273) );
  OAI22_X1 U21118 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n17904), .ZN(n17905) );
  INV_X1 U21119 ( .A(n17905), .ZN(U274) );
  OAI22_X1 U21120 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n17904), .ZN(n17906) );
  INV_X1 U21121 ( .A(n17906), .ZN(U275) );
  OAI22_X1 U21122 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n17904), .ZN(n17907) );
  INV_X1 U21123 ( .A(n17907), .ZN(U276) );
  OAI22_X1 U21124 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n17904), .ZN(n17908) );
  INV_X1 U21125 ( .A(n17908), .ZN(U277) );
  OAI22_X1 U21126 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n17904), .ZN(n17909) );
  INV_X1 U21127 ( .A(n17909), .ZN(U278) );
  OAI22_X1 U21128 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n17904), .ZN(n17910) );
  INV_X1 U21129 ( .A(n17910), .ZN(U279) );
  OAI22_X1 U21130 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n17904), .ZN(n17911) );
  INV_X1 U21131 ( .A(n17911), .ZN(U280) );
  INV_X1 U21132 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n22204) );
  INV_X1 U21133 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n18681) );
  AOI22_X1 U21134 ( .A1(n17904), .A2(n22204), .B1(n18681), .B2(U215), .ZN(U281) );
  INV_X1 U21135 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n18679) );
  AOI22_X1 U21136 ( .A1(n17904), .A2(n20312), .B1(n18679), .B2(U215), .ZN(U282) );
  AOI222_X1 U21137 ( .A1(n20312), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(n17912), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .C1(n18817), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n17913) );
  INV_X2 U21138 ( .A(n17915), .ZN(n17914) );
  INV_X1 U21139 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n20090) );
  INV_X1 U21140 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n21048) );
  AOI22_X1 U21141 ( .A1(n17914), .A2(n20090), .B1(n21048), .B2(n17915), .ZN(
        U347) );
  INV_X1 U21142 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n20088) );
  INV_X1 U21143 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n21047) );
  AOI22_X1 U21144 ( .A1(n17914), .A2(n20088), .B1(n21047), .B2(n17915), .ZN(
        U348) );
  INV_X1 U21145 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n20087) );
  INV_X1 U21146 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n21045) );
  AOI22_X1 U21147 ( .A1(n17914), .A2(n20087), .B1(n21045), .B2(n17915), .ZN(
        U349) );
  INV_X1 U21148 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n20085) );
  INV_X1 U21149 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n21043) );
  AOI22_X1 U21150 ( .A1(n17914), .A2(n20085), .B1(n21043), .B2(n17915), .ZN(
        U350) );
  INV_X1 U21151 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n22006) );
  INV_X1 U21152 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n21041) );
  AOI22_X1 U21153 ( .A1(n17914), .A2(n22006), .B1(n21041), .B2(n17915), .ZN(
        U351) );
  INV_X1 U21154 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n20081) );
  INV_X1 U21155 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n21039) );
  AOI22_X1 U21156 ( .A1(n17914), .A2(n20081), .B1(n21039), .B2(n17915), .ZN(
        U352) );
  INV_X1 U21157 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n20080) );
  INV_X1 U21158 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n21037) );
  AOI22_X1 U21159 ( .A1(n17914), .A2(n20080), .B1(n21037), .B2(n17915), .ZN(
        U353) );
  INV_X1 U21160 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n20078) );
  INV_X1 U21161 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n22020) );
  AOI22_X1 U21162 ( .A1(n17914), .A2(n20078), .B1(n22020), .B2(n17915), .ZN(
        U354) );
  INV_X1 U21163 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n20128) );
  INV_X1 U21164 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n21079) );
  AOI22_X1 U21165 ( .A1(n17914), .A2(n20128), .B1(n21079), .B2(n17915), .ZN(
        U355) );
  INV_X1 U21166 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n20126) );
  INV_X1 U21167 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n22233) );
  AOI22_X1 U21168 ( .A1(n17914), .A2(n20126), .B1(n22233), .B2(n17915), .ZN(
        U356) );
  INV_X1 U21169 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n20122) );
  INV_X1 U21170 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n21075) );
  AOI22_X1 U21171 ( .A1(n17914), .A2(n20122), .B1(n21075), .B2(n17915), .ZN(
        U357) );
  INV_X1 U21172 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n20121) );
  INV_X1 U21173 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n21073) );
  AOI22_X1 U21174 ( .A1(n17914), .A2(n20121), .B1(n21073), .B2(n17915), .ZN(
        U358) );
  INV_X1 U21175 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n20119) );
  INV_X1 U21176 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n22117) );
  AOI22_X1 U21177 ( .A1(n17914), .A2(n20119), .B1(n22117), .B2(n17915), .ZN(
        U359) );
  INV_X1 U21178 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n22195) );
  INV_X1 U21179 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n21071) );
  AOI22_X1 U21180 ( .A1(n17914), .A2(n22195), .B1(n21071), .B2(n17915), .ZN(
        U360) );
  INV_X1 U21181 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n20115) );
  INV_X1 U21182 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n21069) );
  AOI22_X1 U21183 ( .A1(n17914), .A2(n20115), .B1(n21069), .B2(n17915), .ZN(
        U361) );
  INV_X1 U21184 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n20112) );
  INV_X1 U21185 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n21068) );
  AOI22_X1 U21186 ( .A1(n17914), .A2(n20112), .B1(n21068), .B2(n17915), .ZN(
        U362) );
  INV_X1 U21187 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n20111) );
  INV_X1 U21188 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n21066) );
  AOI22_X1 U21189 ( .A1(n17914), .A2(n20111), .B1(n21066), .B2(n17915), .ZN(
        U363) );
  INV_X1 U21190 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n20109) );
  INV_X1 U21191 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n21065) );
  AOI22_X1 U21192 ( .A1(n17914), .A2(n20109), .B1(n21065), .B2(n17915), .ZN(
        U364) );
  INV_X1 U21193 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n20076) );
  INV_X1 U21194 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n21033) );
  AOI22_X1 U21195 ( .A1(n17914), .A2(n20076), .B1(n21033), .B2(n17915), .ZN(
        U365) );
  INV_X1 U21196 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n22155) );
  INV_X1 U21197 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n21063) );
  AOI22_X1 U21198 ( .A1(n17914), .A2(n22155), .B1(n21063), .B2(n17915), .ZN(
        U366) );
  INV_X1 U21199 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n20106) );
  INV_X1 U21200 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n21062) );
  AOI22_X1 U21201 ( .A1(n17914), .A2(n20106), .B1(n21062), .B2(n17915), .ZN(
        U367) );
  INV_X1 U21202 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n22048) );
  INV_X1 U21203 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n21060) );
  AOI22_X1 U21204 ( .A1(n17914), .A2(n22048), .B1(n21060), .B2(n17915), .ZN(
        U368) );
  INV_X1 U21205 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n20103) );
  INV_X1 U21206 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n21059) );
  AOI22_X1 U21207 ( .A1(n17914), .A2(n20103), .B1(n21059), .B2(n17915), .ZN(
        U369) );
  INV_X1 U21208 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n20101) );
  INV_X1 U21209 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n21057) );
  AOI22_X1 U21210 ( .A1(n17914), .A2(n20101), .B1(n21057), .B2(n17915), .ZN(
        U370) );
  INV_X1 U21211 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n20099) );
  INV_X1 U21212 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n22066) );
  AOI22_X1 U21213 ( .A1(n17913), .A2(n20099), .B1(n22066), .B2(n17915), .ZN(
        U371) );
  INV_X1 U21214 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n20097) );
  INV_X1 U21215 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n21054) );
  AOI22_X1 U21216 ( .A1(n17914), .A2(n20097), .B1(n21054), .B2(n17915), .ZN(
        U372) );
  INV_X1 U21217 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n20096) );
  INV_X1 U21218 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n21052) );
  AOI22_X1 U21219 ( .A1(n17913), .A2(n20096), .B1(n21052), .B2(n17915), .ZN(
        U373) );
  INV_X1 U21220 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n20094) );
  INV_X1 U21221 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n21051) );
  AOI22_X1 U21222 ( .A1(n17913), .A2(n20094), .B1(n21051), .B2(n17915), .ZN(
        U374) );
  INV_X1 U21223 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n20092) );
  INV_X1 U21224 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n21049) );
  AOI22_X1 U21225 ( .A1(n17913), .A2(n20092), .B1(n21049), .B2(n17915), .ZN(
        U375) );
  INV_X1 U21226 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n20074) );
  AOI22_X1 U21227 ( .A1(n17914), .A2(n20074), .B1(n21032), .B2(n17915), .ZN(
        U376) );
  NOR2_X1 U21228 ( .A1(n20073), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n17916) );
  NOR2_X1 U21229 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(P3_STATE_REG_1__SCAN_IN), 
        .ZN(n20058) );
  AOI21_X1 U21230 ( .B1(P3_STATE_REG_1__SCAN_IN), .B2(n17916), .A(n20058), 
        .ZN(n20055) );
  INV_X1 U21231 ( .A(n20055), .ZN(n20136) );
  AOI21_X1 U21232 ( .B1(P3_STATE_REG_0__SCAN_IN), .B2(P3_ADS_N_REG_SCAN_IN), 
        .A(n20136), .ZN(n17917) );
  INV_X1 U21233 ( .A(n17917), .ZN(P3_U2633) );
  NAND2_X1 U21234 ( .A1(n20187), .A2(n20138), .ZN(n17923) );
  INV_X1 U21235 ( .A(n20048), .ZN(n17922) );
  NOR2_X1 U21236 ( .A1(n17919), .A2(n17918), .ZN(n17920) );
  OAI21_X1 U21237 ( .B1(n17920), .B2(n18857), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n17921) );
  OAI21_X1 U21238 ( .B1(n17923), .B2(n17922), .A(n17921), .ZN(P3_U2634) );
  NOR2_X1 U21239 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n17925) );
  AOI22_X1 U21240 ( .A1(P3_D_C_N_REG_SCAN_IN), .A2(n20185), .B1(n17925), .B2(
        n20073), .ZN(n17924) );
  OAI21_X1 U21241 ( .B1(P3_CODEFETCH_REG_SCAN_IN), .B2(n20185), .A(n17924), 
        .ZN(P3_U2635) );
  OAI21_X1 U21242 ( .B1(BS16), .B2(n17925), .A(n20136), .ZN(n20135) );
  OAI21_X1 U21243 ( .B1(n20136), .B2(n17926), .A(n20135), .ZN(P3_U2636) );
  INV_X1 U21244 ( .A(n17927), .ZN(n20017) );
  AOI211_X1 U21245 ( .C1(n18858), .C2(n17929), .A(n17928), .B(n20017), .ZN(
        n20026) );
  NOR2_X1 U21246 ( .A1(n20026), .A2(n20042), .ZN(n20168) );
  OAI21_X1 U21247 ( .B1(n20168), .B2(n19523), .A(n17930), .ZN(P3_U2637) );
  NOR4_X1 U21248 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_12__SCAN_IN), .A3(P3_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_14__SCAN_IN), .ZN(n17940) );
  NOR4_X1 U21249 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_6__SCAN_IN), .A3(P3_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_9__SCAN_IN), .ZN(n17939) );
  NOR4_X1 U21250 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_2__SCAN_IN), .A3(P3_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_4__SCAN_IN), .ZN(n17931) );
  INV_X1 U21251 ( .A(P3_DATAWIDTH_REG_8__SCAN_IN), .ZN(n22108) );
  INV_X1 U21252 ( .A(P3_DATAWIDTH_REG_11__SCAN_IN), .ZN(n22026) );
  NAND3_X1 U21253 ( .A1(n17931), .A2(n22108), .A3(n22026), .ZN(n17937) );
  NOR4_X1 U21254 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_20__SCAN_IN), .A3(P3_DATAWIDTH_REG_21__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_22__SCAN_IN), .ZN(n17935) );
  NOR4_X1 U21255 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_15__SCAN_IN), .A3(P3_DATAWIDTH_REG_16__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_18__SCAN_IN), .ZN(n17934) );
  NOR4_X1 U21256 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_28__SCAN_IN), .A3(P3_DATAWIDTH_REG_29__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_30__SCAN_IN), .ZN(n17933) );
  NOR4_X1 U21257 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_24__SCAN_IN), .A3(P3_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n17932) );
  NAND4_X1 U21258 ( .A1(n17935), .A2(n17934), .A3(n17933), .A4(n17932), .ZN(
        n17936) );
  AOI211_X1 U21259 ( .C1(P3_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(n17937), .B(n17936), .ZN(n17938) );
  NAND3_X1 U21260 ( .A1(n17940), .A2(n17939), .A3(n17938), .ZN(n20166) );
  INV_X1 U21261 ( .A(n20166), .ZN(n20160) );
  INV_X1 U21262 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n17941) );
  NOR2_X1 U21263 ( .A1(P3_DATAWIDTH_REG_1__SCAN_IN), .A2(n20166), .ZN(n17942)
         );
  INV_X1 U21264 ( .A(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n20162) );
  NAND3_X1 U21265 ( .A1(n17942), .A2(n13930), .A3(n20162), .ZN(n17943) );
  OAI221_X1 U21266 ( .B1(n20160), .B2(n17941), .C1(n20166), .C2(n17362), .A(
        n17943), .ZN(P3_U2638) );
  INV_X1 U21267 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n17944) );
  NAND2_X1 U21268 ( .A1(n17942), .A2(n17362), .ZN(n20163) );
  OAI211_X1 U21269 ( .C1(n20160), .C2(n17944), .A(n17943), .B(n20163), .ZN(
        P3_U2639) );
  NAND2_X1 U21270 ( .A1(n18259), .A2(n17945), .ZN(n17956) );
  OAI22_X1 U21271 ( .A1(n17961), .A2(n20129), .B1(n17948), .B2(n18252), .ZN(
        n17950) );
  OAI21_X1 U21272 ( .B1(n9707), .B2(n17951), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n17952) );
  AOI22_X1 U21273 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n18288), .B1(
        n9707), .B2(P3_EBX_REG_29__SCAN_IN), .ZN(n17960) );
  INV_X1 U21274 ( .A(n17963), .ZN(n17957) );
  AOI21_X1 U21275 ( .B1(P3_EBX_REG_29__SCAN_IN), .B2(n17957), .A(n17956), .ZN(
        n17958) );
  INV_X1 U21276 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n20123) );
  NAND2_X1 U21277 ( .A1(P3_REIP_REG_27__SCAN_IN), .A2(n20123), .ZN(n17972) );
  AOI22_X1 U21278 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n18288), .B1(
        n9707), .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n17971) );
  INV_X1 U21279 ( .A(n17981), .ZN(n17962) );
  OAI21_X1 U21280 ( .B1(P3_REIP_REG_27__SCAN_IN), .B2(n17980), .A(n17962), 
        .ZN(n17969) );
  AOI211_X1 U21281 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n17977), .A(n17963), .B(
        n18295), .ZN(n17968) );
  AOI211_X1 U21282 ( .C1(n17966), .C2(n17965), .A(n17964), .B(n20051), .ZN(
        n17967) );
  AOI211_X1 U21283 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n17969), .A(n17968), 
        .B(n17967), .ZN(n17970) );
  OAI211_X1 U21284 ( .C1(n17980), .C2(n17972), .A(n17971), .B(n17970), .ZN(
        P3_U2643) );
  AOI211_X1 U21285 ( .C1(n18937), .C2(n17974), .A(n17973), .B(n20051), .ZN(
        n17976) );
  OAI22_X1 U21286 ( .A1(n18943), .A2(n18252), .B1(n18290), .B2(n18346), .ZN(
        n17975) );
  AOI211_X1 U21287 ( .C1(P3_REIP_REG_27__SCAN_IN), .C2(n17981), .A(n17976), 
        .B(n17975), .ZN(n17979) );
  OAI211_X1 U21288 ( .C1(n17985), .C2(n18346), .A(n18259), .B(n17977), .ZN(
        n17978) );
  OAI211_X1 U21289 ( .C1(P3_REIP_REG_27__SCAN_IN), .C2(n17980), .A(n17979), 
        .B(n17978), .ZN(P3_U2644) );
  AOI22_X1 U21290 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(n17981), .B1(n9707), 
        .B2(P3_EBX_REG_26__SCAN_IN), .ZN(n17990) );
  INV_X1 U21291 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n20118) );
  AOI211_X1 U21292 ( .C1(n17984), .C2(n17983), .A(n17982), .B(n20051), .ZN(
        n17987) );
  AOI211_X1 U21293 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n17998), .A(n17985), .B(
        n18295), .ZN(n17986) );
  AOI211_X1 U21294 ( .C1(n17988), .C2(n20118), .A(n17987), .B(n17986), .ZN(
        n17989) );
  OAI211_X1 U21295 ( .C1(n10470), .C2(n18252), .A(n17990), .B(n17989), .ZN(
        P3_U2645) );
  OAI21_X1 U21296 ( .B1(P3_REIP_REG_24__SCAN_IN), .B2(n18291), .A(n18015), 
        .ZN(n17991) );
  AOI22_X1 U21297 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n18288), .B1(
        P3_REIP_REG_25__SCAN_IN), .B2(n17991), .ZN(n18001) );
  OAI21_X1 U21298 ( .B1(n18002), .B2(n18003), .A(n18259), .ZN(n17992) );
  INV_X1 U21299 ( .A(n17992), .ZN(n17999) );
  AOI211_X1 U21300 ( .C1(n17995), .C2(n17994), .A(n17993), .B(n20051), .ZN(
        n17997) );
  AND3_X1 U21301 ( .A1(n20117), .A2(n18009), .A3(P3_REIP_REG_24__SCAN_IN), 
        .ZN(n17996) );
  AOI211_X1 U21302 ( .C1(n17999), .C2(n17998), .A(n17997), .B(n17996), .ZN(
        n18000) );
  OAI211_X1 U21303 ( .C1(n18290), .C2(n18002), .A(n18001), .B(n18000), .ZN(
        P3_U2646) );
  AOI22_X1 U21304 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n18288), .B1(
        n9707), .B2(P3_EBX_REG_24__SCAN_IN), .ZN(n18011) );
  AOI211_X1 U21305 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n18018), .A(n18003), .B(
        n18295), .ZN(n18008) );
  INV_X1 U21306 ( .A(n18004), .ZN(n18005) );
  AOI211_X1 U21307 ( .C1(n18963), .C2(n18006), .A(n18005), .B(n20051), .ZN(
        n18007) );
  AOI211_X1 U21308 ( .C1(n18009), .C2(n20114), .A(n18008), .B(n18007), .ZN(
        n18010) );
  OAI211_X1 U21309 ( .C1(n20114), .C2(n18015), .A(n18011), .B(n18010), .ZN(
        P3_U2647) );
  NOR2_X1 U21310 ( .A1(n18099), .A2(n18022), .ZN(n18038) );
  NAND2_X1 U21311 ( .A1(n18038), .A2(n20113), .ZN(n18021) );
  AOI211_X1 U21312 ( .C1(n18014), .C2(n18013), .A(n18012), .B(n20051), .ZN(
        n18017) );
  OAI22_X1 U21313 ( .A1(n20113), .A2(n18015), .B1(n18290), .B2(n22099), .ZN(
        n18016) );
  AOI211_X1 U21314 ( .C1(n18288), .C2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n18017), .B(n18016), .ZN(n18020) );
  OAI211_X1 U21315 ( .C1(n18025), .C2(n22099), .A(n18259), .B(n18018), .ZN(
        n18019) );
  OAI211_X1 U21316 ( .C1(n18030), .C2(n18021), .A(n18020), .B(n18019), .ZN(
        P3_U2648) );
  OAI21_X1 U21317 ( .B1(n18022), .B2(n18096), .A(n18097), .ZN(n18052) );
  INV_X1 U21318 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n20110) );
  AOI211_X1 U21319 ( .C1(n18997), .C2(n18024), .A(n18023), .B(n20051), .ZN(
        n18029) );
  AOI211_X1 U21320 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n18039), .A(n18025), .B(
        n18295), .ZN(n18028) );
  OAI22_X1 U21321 ( .A1(n18026), .A2(n18252), .B1(n18290), .B2(n18358), .ZN(
        n18027) );
  NOR3_X1 U21322 ( .A1(n18029), .A2(n18028), .A3(n18027), .ZN(n18032) );
  OAI211_X1 U21323 ( .C1(P3_REIP_REG_22__SCAN_IN), .C2(P3_REIP_REG_21__SCAN_IN), .A(n18038), .B(n18030), .ZN(n18031) );
  OAI211_X1 U21324 ( .C1(n18052), .C2(n20110), .A(n18032), .B(n18031), .ZN(
        P3_U2649) );
  AOI22_X1 U21325 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n18288), .B1(
        n9707), .B2(P3_EBX_REG_21__SCAN_IN), .ZN(n18042) );
  INV_X1 U21326 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n20108) );
  INV_X1 U21327 ( .A(n18052), .ZN(n18037) );
  INV_X1 U21328 ( .A(n18033), .ZN(n18034) );
  AOI211_X1 U21329 ( .C1(n19004), .C2(n18035), .A(n18034), .B(n20051), .ZN(
        n18036) );
  AOI221_X1 U21330 ( .B1(n18038), .B2(n20108), .C1(n18037), .C2(
        P3_REIP_REG_21__SCAN_IN), .A(n18036), .ZN(n18041) );
  OAI211_X1 U21331 ( .C1(n18046), .C2(n18389), .A(n18259), .B(n18039), .ZN(
        n18040) );
  NAND3_X1 U21332 ( .A1(n18042), .A2(n18041), .A3(n18040), .ZN(P3_U2650) );
  NAND2_X1 U21333 ( .A1(n18098), .A2(n18043), .ZN(n18053) );
  INV_X1 U21334 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n20107) );
  AOI211_X1 U21335 ( .C1(n19018), .C2(n18045), .A(n18044), .B(n20051), .ZN(
        n18050) );
  AOI211_X1 U21336 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n18063), .A(n18046), .B(
        n18295), .ZN(n18049) );
  AOI22_X1 U21337 ( .A1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n18288), .B1(
        n9707), .B2(P3_EBX_REG_20__SCAN_IN), .ZN(n18047) );
  INV_X1 U21338 ( .A(n18047), .ZN(n18048) );
  NOR3_X1 U21339 ( .A1(n18050), .A2(n18049), .A3(n18048), .ZN(n18051) );
  OAI221_X1 U21340 ( .B1(P3_REIP_REG_20__SCAN_IN), .B2(n18053), .C1(n20107), 
        .C2(n18052), .A(n18051), .ZN(P3_U2651) );
  AOI22_X1 U21341 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n18288), .B1(
        n9707), .B2(P3_EBX_REG_19__SCAN_IN), .ZN(n18067) );
  OR2_X1 U21342 ( .A1(n18054), .A2(n18227), .ZN(n18071) );
  INV_X1 U21343 ( .A(n19025), .ZN(n18078) );
  NOR2_X1 U21344 ( .A1(n19041), .A2(n18078), .ZN(n18056) );
  OAI21_X1 U21345 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n18056), .A(
        n18055), .ZN(n19029) );
  XOR2_X1 U21346 ( .A(n18071), .B(n19029), .Z(n18062) );
  INV_X1 U21347 ( .A(n18058), .ZN(n18057) );
  OAI21_X1 U21348 ( .B1(n18057), .B2(n18096), .A(n18097), .ZN(n18085) );
  INV_X1 U21349 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n20104) );
  NAND3_X1 U21350 ( .A1(n18098), .A2(n18058), .A3(n20104), .ZN(n18076) );
  AOI21_X1 U21351 ( .B1(n18085), .B2(n18076), .A(n20105), .ZN(n18061) );
  NOR3_X1 U21352 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(n18099), .A3(n18059), 
        .ZN(n18060) );
  AOI211_X1 U21353 ( .C1(n18062), .C2(n18280), .A(n18061), .B(n18060), .ZN(
        n18066) );
  OAI211_X1 U21354 ( .C1(n18072), .C2(n18064), .A(n18259), .B(n18063), .ZN(
        n18065) );
  NAND4_X1 U21355 ( .A1(n18067), .A2(n18066), .A3(n14191), .A4(n18065), .ZN(
        P3_U2652) );
  AOI22_X1 U21356 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n18078), .B1(
        n19025), .B2(n19041), .ZN(n19038) );
  NAND2_X1 U21357 ( .A1(n18227), .A2(n18280), .ZN(n18285) );
  INV_X1 U21358 ( .A(n18068), .ZN(n18069) );
  OAI21_X1 U21359 ( .B1(n18069), .B2(n19038), .A(n18280), .ZN(n18070) );
  AOI22_X1 U21360 ( .A1(n19038), .A2(n18071), .B1(n18285), .B2(n18070), .ZN(
        n18075) );
  AOI211_X1 U21361 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n18081), .A(n18072), .B(
        n18295), .ZN(n18074) );
  OAI22_X1 U21362 ( .A1(n19041), .A2(n18252), .B1(n18290), .B2(n18462), .ZN(
        n18073) );
  NOR4_X1 U21363 ( .A1(n19508), .A2(n18075), .A3(n18074), .A4(n18073), .ZN(
        n18077) );
  OAI211_X1 U21364 ( .C1(n18085), .C2(n20104), .A(n18077), .B(n18076), .ZN(
        P3_U2653) );
  INV_X1 U21365 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n18105) );
  NOR2_X1 U21366 ( .A1(n18105), .A2(n18108), .ZN(n18079) );
  OAI21_X1 U21367 ( .B1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n18079), .A(
        n18078), .ZN(n19054) );
  NOR2_X1 U21368 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18301), .ZN(
        n18281) );
  AOI21_X1 U21369 ( .B1(n19053), .B2(n18281), .A(n18227), .ZN(n18080) );
  XOR2_X1 U21370 ( .A(n19054), .B(n18080), .Z(n18091) );
  OAI211_X1 U21371 ( .C1(n18092), .C2(n18083), .A(n18259), .B(n18081), .ZN(
        n18082) );
  OAI211_X1 U21372 ( .C1(n18290), .C2(n18083), .A(n14191), .B(n18082), .ZN(
        n18089) );
  NOR2_X1 U21373 ( .A1(n18099), .A2(n18084), .ZN(n18087) );
  INV_X1 U21374 ( .A(n18085), .ZN(n18086) );
  MUX2_X1 U21375 ( .A(n18087), .B(n18086), .S(P3_REIP_REG_17__SCAN_IN), .Z(
        n18088) );
  AOI211_X1 U21376 ( .C1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .C2(n18288), .A(
        n18089), .B(n18088), .ZN(n18090) );
  OAI21_X1 U21377 ( .B1(n20051), .B2(n18091), .A(n18090), .ZN(P3_U2654) );
  AOI211_X1 U21378 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n18106), .A(n18092), .B(
        n18295), .ZN(n18093) );
  AOI211_X1 U21379 ( .C1(n9707), .C2(P3_EBX_REG_16__SCAN_IN), .A(n19508), .B(
        n18093), .ZN(n18104) );
  NOR2_X1 U21380 ( .A1(n18094), .A2(n18227), .ZN(n18109) );
  INV_X1 U21381 ( .A(n18108), .ZN(n18095) );
  AOI22_X1 U21382 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n18108), .B1(
        n18095), .B2(n18105), .ZN(n19075) );
  XNOR2_X1 U21383 ( .A(n18109), .B(n19075), .ZN(n18102) );
  NAND2_X1 U21384 ( .A1(n18097), .A2(n18096), .ZN(n18117) );
  INV_X1 U21385 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n20098) );
  NAND2_X1 U21386 ( .A1(n18098), .A2(n20098), .ZN(n18114) );
  INV_X1 U21387 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n20100) );
  AOI21_X1 U21388 ( .B1(n18117), .B2(n18114), .A(n20100), .ZN(n18101) );
  NOR3_X1 U21389 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(n18099), .A3(n20098), 
        .ZN(n18100) );
  AOI211_X1 U21390 ( .C1(n18102), .C2(n18280), .A(n18101), .B(n18100), .ZN(
        n18103) );
  OAI211_X1 U21391 ( .C1(n18105), .C2(n18252), .A(n18104), .B(n18103), .ZN(
        P3_U2655) );
  OAI211_X1 U21392 ( .C1(n18119), .C2(n18522), .A(n18259), .B(n18106), .ZN(
        n18107) );
  OAI211_X1 U21393 ( .C1(n18290), .C2(n18522), .A(n14191), .B(n18107), .ZN(
        n18113) );
  NOR2_X1 U21394 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n20051), .ZN(
        n18286) );
  INV_X1 U21395 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n19084) );
  INV_X1 U21396 ( .A(n18285), .ZN(n18287) );
  AOI21_X1 U21397 ( .B1(n18286), .B2(n19084), .A(n18287), .ZN(n18111) );
  OAI21_X1 U21398 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n19069), .A(
        n18108), .ZN(n19081) );
  NAND3_X1 U21399 ( .A1(n18280), .A2(n18109), .A3(n19081), .ZN(n18110) );
  OAI21_X1 U21400 ( .B1(n18111), .B2(n19081), .A(n18110), .ZN(n18112) );
  AOI211_X1 U21401 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(n18288), .A(
        n18113), .B(n18112), .ZN(n18115) );
  OAI211_X1 U21402 ( .C1(n18117), .C2(n20098), .A(n18115), .B(n18114), .ZN(
        P3_U2656) );
  INV_X1 U21403 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n18120) );
  NAND2_X1 U21404 ( .A1(n19098), .A2(n18116), .ZN(n18127) );
  AOI21_X1 U21405 ( .B1(n18120), .B2(n18127), .A(n19069), .ZN(n19099) );
  INV_X1 U21406 ( .A(n19098), .ZN(n19115) );
  NAND2_X1 U21407 ( .A1(n9890), .A2(n18281), .ZN(n18146) );
  OAI21_X1 U21408 ( .B1(n19115), .B2(n18146), .A(n18289), .ZN(n18138) );
  INV_X1 U21409 ( .A(n19099), .ZN(n18126) );
  AOI21_X1 U21410 ( .B1(n18286), .B2(n18120), .A(n18287), .ZN(n18125) );
  AOI21_X1 U21411 ( .B1(n22146), .B2(n18118), .A(n18117), .ZN(n18123) );
  AOI211_X1 U21412 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n18130), .A(n18119), .B(
        n18295), .ZN(n18122) );
  INV_X1 U21413 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n18541) );
  OAI22_X1 U21414 ( .A1(n18120), .A2(n18252), .B1(n18290), .B2(n18541), .ZN(
        n18121) );
  NOR4_X1 U21415 ( .A1(n19508), .A2(n18123), .A3(n18122), .A4(n18121), .ZN(
        n18124) );
  OAI221_X1 U21416 ( .B1(n19099), .B2(n18138), .C1(n18126), .C2(n18125), .A(
        n18124), .ZN(P3_U2657) );
  NOR2_X1 U21417 ( .A1(n18145), .A2(n19112), .ZN(n18144) );
  OAI21_X1 U21418 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n18144), .A(
        n18127), .ZN(n19117) );
  INV_X1 U21419 ( .A(n19117), .ZN(n18139) );
  AOI21_X1 U21420 ( .B1(n18144), .B2(n18286), .A(n18287), .ZN(n18137) );
  OAI21_X1 U21421 ( .B1(n18143), .B2(n18291), .A(n18242), .ZN(n18162) );
  NOR2_X1 U21422 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n18291), .ZN(n18142) );
  NOR3_X1 U21423 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(n18291), .A3(n18128), 
        .ZN(n18129) );
  AOI211_X1 U21424 ( .C1(n9707), .C2(P3_EBX_REG_13__SCAN_IN), .A(n19508), .B(
        n18129), .ZN(n18133) );
  OAI211_X1 U21425 ( .C1(n18140), .C2(n18131), .A(n18259), .B(n18130), .ZN(
        n18132) );
  OAI211_X1 U21426 ( .C1(n18252), .C2(n18134), .A(n18133), .B(n18132), .ZN(
        n18135) );
  AOI221_X1 U21427 ( .B1(n18162), .B2(P3_REIP_REG_13__SCAN_IN), .C1(n18142), 
        .C2(P3_REIP_REG_13__SCAN_IN), .A(n18135), .ZN(n18136) );
  OAI221_X1 U21428 ( .B1(n18139), .B2(n18138), .C1(n19117), .C2(n18137), .A(
        n18136), .ZN(P3_U2658) );
  AOI211_X1 U21429 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n18156), .A(n18140), .B(
        n18295), .ZN(n18141) );
  AOI21_X1 U21430 ( .B1(P3_EBX_REG_12__SCAN_IN), .B2(n9707), .A(n18141), .ZN(
        n18151) );
  AOI22_X1 U21431 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n18288), .B1(
        n18143), .B2(n18142), .ZN(n18150) );
  AOI21_X1 U21432 ( .B1(n18145), .B2(n19112), .A(n18144), .ZN(n19127) );
  NAND2_X1 U21433 ( .A1(n17277), .A2(n18146), .ZN(n18147) );
  XNOR2_X1 U21434 ( .A(n19127), .B(n18147), .ZN(n18148) );
  AOI22_X1 U21435 ( .A1(n18280), .A2(n18148), .B1(P3_REIP_REG_12__SCAN_IN), 
        .B2(n18162), .ZN(n18149) );
  NAND4_X1 U21436 ( .A1(n18151), .A2(n18150), .A3(n18149), .A4(n14191), .ZN(
        P3_U2659) );
  NOR2_X1 U21437 ( .A1(n18291), .A2(n18174), .ZN(n18222) );
  OAI21_X1 U21438 ( .B1(n18152), .B2(n18205), .A(n20091), .ZN(n18161) );
  INV_X1 U21439 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n18159) );
  INV_X1 U21440 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n19152) );
  NOR2_X1 U21441 ( .A1(n19152), .A2(n18184), .ZN(n18170) );
  OAI21_X1 U21442 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n18170), .A(
        n19112), .ZN(n19140) );
  NAND2_X1 U21443 ( .A1(n18171), .A2(n18281), .ZN(n18153) );
  OAI21_X1 U21444 ( .B1(n19152), .B2(n18153), .A(n17277), .ZN(n18155) );
  AOI21_X1 U21445 ( .B1(n19140), .B2(n18155), .A(n20051), .ZN(n18154) );
  OAI21_X1 U21446 ( .B1(n19140), .B2(n18155), .A(n18154), .ZN(n18158) );
  OAI211_X1 U21447 ( .C1(n18165), .C2(n18164), .A(n18259), .B(n18156), .ZN(
        n18157) );
  OAI211_X1 U21448 ( .C1(n18252), .C2(n18159), .A(n18158), .B(n18157), .ZN(
        n18160) );
  AOI21_X1 U21449 ( .B1(n18162), .B2(n18161), .A(n18160), .ZN(n18163) );
  OAI211_X1 U21450 ( .C1(n18290), .C2(n18164), .A(n18163), .B(n14191), .ZN(
        P3_U2660) );
  AOI22_X1 U21451 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n18288), .B1(
        n9707), .B2(P3_EBX_REG_10__SCAN_IN), .ZN(n18179) );
  NOR2_X1 U21452 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(n18205), .ZN(n18168) );
  AOI211_X1 U21453 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n18166), .A(n18165), .B(
        n18295), .ZN(n18167) );
  AOI211_X1 U21454 ( .C1(n18169), .C2(n18168), .A(n19508), .B(n18167), .ZN(
        n18178) );
  AOI21_X1 U21455 ( .B1(n19152), .B2(n18184), .A(n18170), .ZN(n19153) );
  AOI21_X1 U21456 ( .B1(n18171), .B2(n18281), .A(n18227), .ZN(n18185) );
  AOI21_X1 U21457 ( .B1(n19153), .B2(n18185), .A(n20051), .ZN(n18172) );
  OAI21_X1 U21458 ( .B1(n19153), .B2(n18185), .A(n18172), .ZN(n18177) );
  NOR3_X1 U21459 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n18173), .A3(n18205), .ZN(
        n18189) );
  INV_X1 U21460 ( .A(n18173), .ZN(n18175) );
  AOI21_X1 U21461 ( .B1(n18272), .B2(n18174), .A(n18298), .ZN(n18230) );
  OAI21_X1 U21462 ( .B1(n18175), .B2(n18291), .A(n18230), .ZN(n18180) );
  OAI21_X1 U21463 ( .B1(n18189), .B2(n18180), .A(P3_REIP_REG_10__SCAN_IN), 
        .ZN(n18176) );
  NAND4_X1 U21464 ( .A1(n18179), .A2(n18178), .A3(n18177), .A4(n18176), .ZN(
        P3_U2661) );
  INV_X1 U21465 ( .A(n18180), .ZN(n18204) );
  INV_X1 U21466 ( .A(n18181), .ZN(n18182) );
  AOI211_X1 U21467 ( .C1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .C2(n18288), .A(
        n19508), .B(n18182), .ZN(n18193) );
  NOR2_X1 U21468 ( .A1(n18183), .A2(n18295), .ZN(n18195) );
  INV_X1 U21469 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n19179) );
  NOR2_X1 U21470 ( .A1(n19179), .A2(n18197), .ZN(n18196) );
  OAI21_X1 U21471 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n18196), .A(
        n18184), .ZN(n19167) );
  INV_X1 U21472 ( .A(n18185), .ZN(n18188) );
  INV_X1 U21473 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n18186) );
  AOI211_X1 U21474 ( .C1(n18196), .C2(n18186), .A(n18227), .B(n19167), .ZN(
        n18187) );
  AOI211_X1 U21475 ( .C1(n19167), .C2(n18188), .A(n18187), .B(n20051), .ZN(
        n18190) );
  AOI211_X1 U21476 ( .C1(n18195), .C2(n18191), .A(n18190), .B(n18189), .ZN(
        n18192) );
  OAI211_X1 U21477 ( .C1(n18204), .C2(n22085), .A(n18193), .B(n18192), .ZN(
        P3_U2662) );
  INV_X1 U21478 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n20086) );
  NAND2_X1 U21479 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n18212), .ZN(n18194) );
  AOI22_X1 U21480 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n9707), .B1(n18195), .B2(
        n18194), .ZN(n18203) );
  AOI21_X1 U21481 ( .B1(n19179), .B2(n18197), .A(n18196), .ZN(n19184) );
  OAI21_X1 U21482 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n18197), .A(
        n17277), .ZN(n18198) );
  XNOR2_X1 U21483 ( .A(n19184), .B(n18198), .ZN(n18201) );
  NAND3_X1 U21484 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(P3_REIP_REG_6__SCAN_IN), 
        .A3(n20086), .ZN(n18199) );
  OAI22_X1 U21485 ( .A1(n19179), .A2(n18252), .B1(n18205), .B2(n18199), .ZN(
        n18200) );
  AOI211_X1 U21486 ( .C1(n18280), .C2(n18201), .A(n19508), .B(n18200), .ZN(
        n18202) );
  OAI211_X1 U21487 ( .C1(n18204), .C2(n20086), .A(n18203), .B(n18202), .ZN(
        P3_U2663) );
  OAI21_X1 U21488 ( .B1(P3_REIP_REG_6__SCAN_IN), .B2(n18205), .A(n18230), .ZN(
        n18223) );
  AOI21_X1 U21489 ( .B1(n18206), .B2(n18281), .A(n18227), .ZN(n18218) );
  OAI21_X1 U21490 ( .B1(n18208), .B2(n18218), .A(n18280), .ZN(n18207) );
  AOI21_X1 U21491 ( .B1(n18208), .B2(n18218), .A(n18207), .ZN(n18211) );
  NAND3_X1 U21492 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n18222), .A3(n20084), 
        .ZN(n18209) );
  OAI211_X1 U21493 ( .C1(n19165), .C2(n18252), .A(n14191), .B(n18209), .ZN(
        n18210) );
  AOI211_X1 U21494 ( .C1(P3_REIP_REG_7__SCAN_IN), .C2(n18223), .A(n18211), .B(
        n18210), .ZN(n18214) );
  OAI211_X1 U21495 ( .C1(n18215), .C2(n18633), .A(n18259), .B(n18212), .ZN(
        n18213) );
  OAI211_X1 U21496 ( .C1(n18633), .C2(n18290), .A(n18214), .B(n18213), .ZN(
        P3_U2664) );
  AOI211_X1 U21497 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n18232), .A(n18215), .B(
        n18295), .ZN(n18216) );
  AOI211_X1 U21498 ( .C1(n9707), .C2(P3_EBX_REG_6__SCAN_IN), .A(n19508), .B(
        n18216), .ZN(n18225) );
  AOI21_X1 U21499 ( .B1(n18286), .B2(n22084), .A(n18287), .ZN(n18220) );
  NOR2_X1 U21500 ( .A1(n18301), .A2(n19193), .ZN(n18226) );
  OAI21_X1 U21501 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n18226), .A(
        n18217), .ZN(n19200) );
  NAND3_X1 U21502 ( .A1(n18280), .A2(n18218), .A3(n19200), .ZN(n18219) );
  OAI21_X1 U21503 ( .B1(n18220), .B2(n19200), .A(n18219), .ZN(n18221) );
  AOI221_X1 U21504 ( .B1(P3_REIP_REG_6__SCAN_IN), .B2(n18223), .C1(n18222), 
        .C2(n18223), .A(n18221), .ZN(n18224) );
  OAI211_X1 U21505 ( .C1(n22084), .C2(n18252), .A(n18225), .B(n18224), .ZN(
        P3_U2665) );
  NOR3_X1 U21506 ( .A1(n18291), .A2(n20077), .A3(n18271), .ZN(n18249) );
  AOI21_X1 U21507 ( .B1(P3_REIP_REG_4__SCAN_IN), .B2(n18249), .A(
        P3_REIP_REG_5__SCAN_IN), .ZN(n18229) );
  NAND3_X1 U21508 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A3(n10078), .ZN(n18245) );
  AOI21_X1 U21509 ( .B1(n10077), .B2(n18245), .A(n18226), .ZN(n19216) );
  AOI21_X1 U21510 ( .B1(n19208), .B2(n18281), .A(n18227), .ZN(n18246) );
  XNOR2_X1 U21511 ( .A(n19216), .B(n18246), .ZN(n18228) );
  OAI22_X1 U21512 ( .A1(n18230), .A2(n18229), .B1(n20051), .B2(n18228), .ZN(
        n18231) );
  AOI211_X1 U21513 ( .C1(n9707), .C2(P3_EBX_REG_5__SCAN_IN), .A(n19508), .B(
        n18231), .ZN(n18234) );
  OAI211_X1 U21514 ( .C1(n18235), .C2(n18641), .A(n18259), .B(n18232), .ZN(
        n18233) );
  OAI211_X1 U21515 ( .C1(n18252), .C2(n10077), .A(n18234), .B(n18233), .ZN(
        P3_U2666) );
  AOI211_X1 U21516 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n18258), .A(n18235), .B(
        n18295), .ZN(n18241) );
  NAND2_X1 U21517 ( .A1(n9723), .A2(n18236), .ZN(n18237) );
  NAND2_X1 U21518 ( .A1(n20192), .A2(n18237), .ZN(n18239) );
  NAND2_X1 U21519 ( .A1(n9707), .A2(P3_EBX_REG_4__SCAN_IN), .ZN(n18238) );
  NAND3_X1 U21520 ( .A1(n18239), .A2(n18238), .A3(n14191), .ZN(n18240) );
  NOR2_X1 U21521 ( .A1(n18241), .A2(n18240), .ZN(n18251) );
  OAI21_X1 U21522 ( .B1(n18243), .B2(n18291), .A(n18242), .ZN(n18263) );
  INV_X1 U21523 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n20079) );
  NOR2_X1 U21524 ( .A1(n18244), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n19221) );
  NOR2_X1 U21525 ( .A1(n18301), .A2(n18244), .ZN(n18253) );
  OAI21_X1 U21526 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n18253), .A(
        n18245), .ZN(n19225) );
  AOI22_X1 U21527 ( .A1(n18281), .A2(n19221), .B1(n18246), .B2(n19225), .ZN(
        n18247) );
  OAI22_X1 U21528 ( .A1(n18247), .A2(n20051), .B1(n19225), .B2(n18285), .ZN(
        n18248) );
  AOI221_X1 U21529 ( .B1(n18263), .B2(P3_REIP_REG_4__SCAN_IN), .C1(n18249), 
        .C2(n20079), .A(n18248), .ZN(n18250) );
  OAI211_X1 U21530 ( .C1(n22149), .C2(n18252), .A(n18251), .B(n18250), .ZN(
        P3_U2667) );
  INV_X1 U21531 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n19240) );
  AOI21_X1 U21532 ( .B1(n19240), .B2(n18254), .A(n18253), .ZN(n19229) );
  OAI21_X1 U21533 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n18254), .A(
        n17277), .ZN(n18278) );
  XOR2_X1 U21534 ( .A(n19229), .B(n18278), .Z(n18266) );
  AOI22_X1 U21535 ( .A1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n18288), .B1(
        n9707), .B2(P3_EBX_REG_3__SCAN_IN), .ZN(n18265) );
  NOR2_X1 U21536 ( .A1(n18291), .A2(n18271), .ZN(n18262) );
  NAND2_X1 U21537 ( .A1(n18256), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n18269) );
  NAND2_X1 U21538 ( .A1(n18269), .A2(n20146), .ZN(n18257) );
  NAND2_X1 U21539 ( .A1(n18257), .A2(n9723), .ZN(n20141) );
  OAI211_X1 U21540 ( .C1(n18267), .C2(n18649), .A(n18259), .B(n18258), .ZN(
        n18260) );
  OAI21_X1 U21541 ( .B1(n18293), .B2(n20141), .A(n18260), .ZN(n18261) );
  AOI221_X1 U21542 ( .B1(n18263), .B2(P3_REIP_REG_3__SCAN_IN), .C1(n18262), 
        .C2(n20077), .A(n18261), .ZN(n18264) );
  OAI211_X1 U21543 ( .C1(n20051), .C2(n18266), .A(n18265), .B(n18264), .ZN(
        P3_U2668) );
  NAND2_X1 U21544 ( .A1(n18669), .A2(n18663), .ZN(n18268) );
  AOI211_X1 U21545 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n18268), .A(n18267), .B(
        n18295), .ZN(n18277) );
  INV_X1 U21546 ( .A(n18269), .ZN(n19981) );
  NOR2_X1 U21547 ( .A1(n18270), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n19982) );
  NOR2_X1 U21548 ( .A1(n19981), .A2(n19982), .ZN(n20150) );
  AOI22_X1 U21549 ( .A1(P3_REIP_REG_2__SCAN_IN), .A2(n18298), .B1(n20150), 
        .B2(n20192), .ZN(n18274) );
  OAI211_X1 U21550 ( .C1(P3_REIP_REG_1__SCAN_IN), .C2(P3_REIP_REG_2__SCAN_IN), 
        .A(n18272), .B(n18271), .ZN(n18273) );
  OAI211_X1 U21551 ( .C1(n18275), .C2(n18290), .A(n18274), .B(n18273), .ZN(
        n18276) );
  AOI211_X1 U21552 ( .C1(n18288), .C2(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n18277), .B(n18276), .ZN(n18283) );
  INV_X1 U21553 ( .A(n18278), .ZN(n18279) );
  OAI211_X1 U21554 ( .C1(n18281), .C2(n18284), .A(n18280), .B(n18279), .ZN(
        n18282) );
  OAI211_X1 U21555 ( .C1(n18285), .C2(n18284), .A(n18283), .B(n18282), .ZN(
        P3_U2669) );
  NOR2_X1 U21556 ( .A1(n18287), .A2(n18286), .ZN(n18302) );
  AOI21_X1 U21557 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n18289), .A(
        n18288), .ZN(n18300) );
  OAI22_X1 U21558 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n18291), .B1(n18290), 
        .B2(n18663), .ZN(n18297) );
  OAI21_X1 U21559 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(P3_EBX_REG_1__SCAN_IN), 
        .A(n18292), .ZN(n18665) );
  OAI22_X1 U21560 ( .A1(n18295), .A2(n18665), .B1(n18294), .B2(n18293), .ZN(
        n18296) );
  AOI211_X1 U21561 ( .C1(P3_REIP_REG_1__SCAN_IN), .C2(n18298), .A(n18297), .B(
        n18296), .ZN(n18299) );
  OAI221_X1 U21562 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n18302), .C1(
        n18301), .C2(n18300), .A(n18299), .ZN(P3_U2670) );
  NAND2_X1 U21563 ( .A1(n18304), .A2(n18303), .ZN(n18305) );
  NAND2_X1 U21564 ( .A1(n18305), .A2(n18661), .ZN(n18332) );
  INV_X1 U21565 ( .A(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n22036) );
  INV_X1 U21566 ( .A(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n18528) );
  INV_X1 U21567 ( .A(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n19675) );
  OAI22_X1 U21568 ( .A1(n22203), .A2(n18613), .B1(n19675), .B2(n18466), .ZN(
        n18311) );
  OAI22_X1 U21569 ( .A1(n9786), .A2(n18527), .B1(n9723), .B2(n18306), .ZN(
        n18307) );
  AOI21_X1 U21570 ( .B1(n18626), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A(
        n18307), .ZN(n18309) );
  AOI22_X1 U21571 ( .A1(n18390), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11911), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n18308) );
  OAI211_X1 U21572 ( .C1(n9718), .C2(n18369), .A(n18309), .B(n18308), .ZN(
        n18310) );
  AOI211_X1 U21573 ( .C1(n9726), .C2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A(
        n18311), .B(n18310), .ZN(n18312) );
  OAI21_X1 U21574 ( .B1(n18615), .B2(n18528), .A(n18312), .ZN(n18314) );
  INV_X1 U21575 ( .A(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n18524) );
  OAI22_X1 U21576 ( .A1(n10660), .A2(n18644), .B1(n17550), .B2(n18524), .ZN(
        n18313) );
  AOI211_X1 U21577 ( .C1(n18586), .C2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A(
        n18314), .B(n18313), .ZN(n18316) );
  AOI22_X1 U21578 ( .A1(n17547), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n9724), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n18315) );
  OAI211_X1 U21579 ( .C1(n22036), .C2(n18599), .A(n18316), .B(n18315), .ZN(
        n18317) );
  INV_X1 U21580 ( .A(n18317), .ZN(n18336) );
  NOR2_X1 U21581 ( .A1(n18336), .A2(n18335), .ZN(n18334) );
  OAI22_X1 U21582 ( .A1(n18611), .A2(n18318), .B1(n18525), .B2(n21957), .ZN(
        n18326) );
  AOI22_X1 U21583 ( .A1(n17547), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n9724), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n18324) );
  AOI22_X1 U21584 ( .A1(n18620), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n18619), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n18323) );
  INV_X1 U21585 ( .A(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n18319) );
  OAI22_X1 U21586 ( .A1(n18613), .A2(n18319), .B1(n9723), .B2(n17221), .ZN(
        n18320) );
  INV_X1 U21587 ( .A(n18320), .ZN(n18322) );
  OR2_X1 U21588 ( .A1(n17550), .A2(n22079), .ZN(n18321) );
  NAND4_X1 U21589 ( .A1(n18324), .A2(n18323), .A3(n18322), .A4(n18321), .ZN(
        n18325) );
  AOI211_X1 U21590 ( .C1(n18413), .C2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A(
        n18326), .B(n18325), .ZN(n18330) );
  AOI22_X1 U21591 ( .A1(n11911), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n14232), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n18329) );
  AOI22_X1 U21592 ( .A1(n18597), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n18403), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n18328) );
  AOI22_X1 U21593 ( .A1(n18628), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n9726), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n18327) );
  NAND4_X1 U21594 ( .A1(n18330), .A2(n18329), .A3(n18328), .A4(n18327), .ZN(
        n18331) );
  XNOR2_X1 U21595 ( .A(n18334), .B(n18331), .ZN(n18682) );
  OAI22_X1 U21596 ( .A1(n18333), .A2(n18332), .B1(n18682), .B2(n18661), .ZN(
        P3_U2673) );
  AOI21_X1 U21597 ( .B1(n18336), .B2(n18335), .A(n18334), .ZN(n18686) );
  AOI22_X1 U21598 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n18337), .B1(n18686), 
        .B2(n18667), .ZN(n18341) );
  NAND4_X1 U21599 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n18357), .A3(n18339), 
        .A4(n18338), .ZN(n18340) );
  NAND2_X1 U21600 ( .A1(n18341), .A2(n18340), .ZN(P3_U2674) );
  AOI21_X1 U21601 ( .B1(n18343), .B2(n18348), .A(n18342), .ZN(n18695) );
  NAND2_X1 U21602 ( .A1(n18667), .A2(n18695), .ZN(n18344) );
  OAI221_X1 U21603 ( .B1(P3_EBX_REG_27__SCAN_IN), .B2(n18347), .C1(n18346), 
        .C2(n18345), .A(n18344), .ZN(P3_U2676) );
  INV_X1 U21604 ( .A(n18347), .ZN(n18351) );
  AOI21_X1 U21605 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n18661), .A(n18357), .ZN(
        n18350) );
  OAI21_X1 U21606 ( .B1(n18353), .B2(n18349), .A(n18348), .ZN(n18704) );
  OAI22_X1 U21607 ( .A1(n18351), .A2(n18350), .B1(n18661), .B2(n18704), .ZN(
        P3_U2677) );
  INV_X1 U21608 ( .A(n18352), .ZN(n18363) );
  AOI21_X1 U21609 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n18661), .A(n18363), .ZN(
        n18356) );
  AOI21_X1 U21610 ( .B1(n18354), .B2(n18359), .A(n18353), .ZN(n18705) );
  INV_X1 U21611 ( .A(n18705), .ZN(n18355) );
  OAI22_X1 U21612 ( .A1(n18357), .A2(n18356), .B1(n18661), .B2(n18355), .ZN(
        P3_U2678) );
  NOR3_X1 U21613 ( .A1(n18765), .A2(n18389), .A3(n9795), .ZN(n18386) );
  INV_X1 U21614 ( .A(n18386), .ZN(n18409) );
  AOI21_X1 U21615 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n18661), .A(n18367), .ZN(
        n18362) );
  OAI21_X1 U21616 ( .B1(n18361), .B2(n18360), .A(n18359), .ZN(n18714) );
  OAI22_X1 U21617 ( .A1(n18363), .A2(n18362), .B1(n18661), .B2(n18714), .ZN(
        P3_U2679) );
  AOI21_X1 U21618 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n18661), .A(n18388), .ZN(
        n18366) );
  XNOR2_X1 U21619 ( .A(n18365), .B(n18364), .ZN(n18717) );
  OAI22_X1 U21620 ( .A1(n18367), .A2(n18366), .B1(n18661), .B2(n18717), .ZN(
        P3_U2680) );
  NAND2_X1 U21621 ( .A1(n9724), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n18368) );
  OAI21_X1 U21622 ( .B1(n18524), .B2(n18616), .A(n18368), .ZN(n18372) );
  INV_X1 U21623 ( .A(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n18370) );
  OAI22_X1 U21624 ( .A1(n18613), .A2(n18370), .B1(n9723), .B2(n18369), .ZN(
        n18371) );
  NOR2_X1 U21625 ( .A1(n18372), .A2(n18371), .ZN(n18379) );
  AOI22_X1 U21626 ( .A1(n18586), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n18390), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n18378) );
  NAND2_X1 U21627 ( .A1(n18620), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n18374) );
  NAND2_X1 U21628 ( .A1(n18619), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n18373) );
  OAI211_X1 U21629 ( .C1(n17550), .C2(n19675), .A(n18374), .B(n18373), .ZN(
        n18375) );
  INV_X1 U21630 ( .A(n18375), .ZN(n18377) );
  NAND2_X1 U21631 ( .A1(n18413), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n18376) );
  NAND4_X1 U21632 ( .A1(n18379), .A2(n18378), .A3(n18377), .A4(n18376), .ZN(
        n18385) );
  AOI22_X1 U21633 ( .A1(n18626), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n18403), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n18383) );
  AOI22_X1 U21634 ( .A1(n11911), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n14232), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n18382) );
  OR2_X1 U21635 ( .A1(n18599), .A2(n18644), .ZN(n18381) );
  NAND2_X1 U21636 ( .A1(n9726), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n18380) );
  NAND4_X1 U21637 ( .A1(n18383), .A2(n18382), .A3(n18381), .A4(n18380), .ZN(
        n18384) );
  NOR2_X1 U21638 ( .A1(n18385), .A2(n18384), .ZN(n18721) );
  AOI21_X1 U21639 ( .B1(P3_EBX_REG_22__SCAN_IN), .B2(n18661), .A(n18386), .ZN(
        n18387) );
  OAI22_X1 U21640 ( .A1(n18721), .A2(n18661), .B1(n18388), .B2(n18387), .ZN(
        P3_U2681) );
  AOI21_X1 U21641 ( .B1(n18389), .B2(n9795), .A(n18667), .ZN(n18408) );
  INV_X1 U21642 ( .A(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n18392) );
  OAI22_X1 U21643 ( .A1(n18611), .A2(n18392), .B1(n18525), .B2(n18391), .ZN(
        n18402) );
  INV_X1 U21644 ( .A(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n19670) );
  OAI22_X1 U21645 ( .A1(n18556), .A2(n18394), .B1(n18616), .B2(n18393), .ZN(
        n18398) );
  OAI22_X1 U21646 ( .A1(n18613), .A2(n18396), .B1(n9723), .B2(n18395), .ZN(
        n18397) );
  NOR2_X1 U21647 ( .A1(n18398), .A2(n18397), .ZN(n18400) );
  AOI22_X1 U21648 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18620), .B1(
        n18489), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n18399) );
  OAI211_X1 U21649 ( .C1(n19670), .C2(n17550), .A(n18400), .B(n18399), .ZN(
        n18401) );
  AOI211_X1 U21650 ( .C1(n18413), .C2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A(
        n18402), .B(n18401), .ZN(n18407) );
  AOI22_X1 U21651 ( .A1(n11911), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n14232), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n18406) );
  AOI22_X1 U21652 ( .A1(n18597), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n18403), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n18405) );
  AOI22_X1 U21653 ( .A1(n18628), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n9726), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n18404) );
  NAND4_X1 U21654 ( .A1(n18407), .A2(n18406), .A3(n18405), .A4(n18404), .ZN(
        n18730) );
  AOI22_X1 U21655 ( .A1(n18409), .A2(n18408), .B1(n18730), .B2(n18667), .ZN(
        n18410) );
  INV_X1 U21656 ( .A(n18410), .ZN(P3_U2682) );
  AOI22_X1 U21657 ( .A1(n18597), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n18390), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n18426) );
  INV_X1 U21658 ( .A(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n18416) );
  OAI22_X1 U21659 ( .A1(n18611), .A2(n18411), .B1(n10660), .B2(n18552), .ZN(
        n18412) );
  AOI21_X1 U21660 ( .B1(n18413), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A(
        n18412), .ZN(n18415) );
  AOI22_X1 U21661 ( .A1(n18585), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n9724), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n18414) );
  OAI211_X1 U21662 ( .C1(n9783), .C2(n18416), .A(n18415), .B(n18414), .ZN(
        n18424) );
  AOI22_X1 U21663 ( .A1(n18620), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n18489), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n18417) );
  OAI21_X1 U21664 ( .B1(n17550), .B2(n19667), .A(n18417), .ZN(n18423) );
  OAI22_X1 U21665 ( .A1(n18616), .A2(n18550), .B1(n9723), .B2(n18418), .ZN(
        n18422) );
  INV_X1 U21666 ( .A(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n18419) );
  OAI22_X1 U21667 ( .A1(n11861), .A2(n18420), .B1(n18615), .B2(n18419), .ZN(
        n18421) );
  NOR4_X1 U21668 ( .A1(n18424), .A2(n18423), .A3(n18422), .A4(n18421), .ZN(
        n18425) );
  OAI211_X1 U21669 ( .C1(n18599), .C2(n18650), .A(n18426), .B(n18425), .ZN(
        n18735) );
  INV_X1 U21670 ( .A(n18735), .ZN(n18428) );
  OAI21_X1 U21671 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n18445), .A(n9795), .ZN(
        n18427) );
  AOI22_X1 U21672 ( .A1(n18667), .A2(n18428), .B1(n18427), .B2(n18661), .ZN(
        P3_U2683) );
  OAI21_X1 U21673 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n18429), .A(n18661), .ZN(
        n18444) );
  OAI22_X1 U21674 ( .A1(n18611), .A2(n18575), .B1(n18551), .B2(n18430), .ZN(
        n18439) );
  AOI22_X1 U21675 ( .A1(n18390), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n9724), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n18437) );
  AOI22_X1 U21676 ( .A1(n18620), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n18619), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n18436) );
  OAI22_X1 U21677 ( .A1(n18616), .A2(n18572), .B1(n9723), .B2(n18431), .ZN(
        n18432) );
  INV_X1 U21678 ( .A(n18432), .ZN(n18435) );
  INV_X1 U21679 ( .A(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n18433) );
  OR2_X1 U21680 ( .A1(n17550), .A2(n18433), .ZN(n18434) );
  NAND4_X1 U21681 ( .A1(n18437), .A2(n18436), .A3(n18435), .A4(n18434), .ZN(
        n18438) );
  AOI211_X1 U21682 ( .C1(n18591), .C2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A(
        n18439), .B(n18438), .ZN(n18443) );
  AOI22_X1 U21683 ( .A1(n18585), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11911), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n18442) );
  AOI22_X1 U21684 ( .A1(n18627), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n14232), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n18441) );
  AOI22_X1 U21685 ( .A1(n18628), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n9726), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n18440) );
  AND4_X1 U21686 ( .A1(n18443), .A2(n18442), .A3(n18441), .A4(n18440), .ZN(
        n18742) );
  OAI22_X1 U21687 ( .A1(n18445), .A2(n18444), .B1(n18742), .B2(n18661), .ZN(
        P3_U2684) );
  INV_X1 U21688 ( .A(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n18446) );
  OAI22_X1 U21689 ( .A1(n18611), .A2(n22105), .B1(n18525), .B2(n18446), .ZN(
        n18456) );
  NOR2_X1 U21690 ( .A1(n9723), .A2(n18447), .ZN(n18451) );
  OAI22_X1 U21691 ( .A1(n18556), .A2(n18449), .B1(n18616), .B2(n18448), .ZN(
        n18450) );
  AOI211_X1 U21692 ( .C1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .C2(n18585), .A(
        n18451), .B(n18450), .ZN(n18453) );
  AOI22_X1 U21693 ( .A1(n18620), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n18619), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n18452) );
  OAI211_X1 U21694 ( .C1(n17550), .C2(n18454), .A(n18453), .B(n18452), .ZN(
        n18455) );
  AOI211_X1 U21695 ( .C1(n18591), .C2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A(
        n18456), .B(n18455), .ZN(n18460) );
  AOI22_X1 U21696 ( .A1(n11911), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n14232), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n18459) );
  AOI22_X1 U21697 ( .A1(n18626), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n18627), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n18458) );
  AOI22_X1 U21698 ( .A1(n18628), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n9726), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n18457) );
  NAND4_X1 U21699 ( .A1(n18460), .A2(n18459), .A3(n18458), .A4(n18457), .ZN(
        n18743) );
  OAI33_X1 U21700 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n18481), .A3(n18765), 
        .B1(n18462), .B2(n18667), .B3(n18461), .ZN(n18463) );
  AOI21_X1 U21701 ( .B1(n18667), .B2(n18743), .A(n18463), .ZN(n18464) );
  INV_X1 U21702 ( .A(n18464), .ZN(P3_U2685) );
  INV_X1 U21703 ( .A(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n18473) );
  INV_X1 U21704 ( .A(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n18594) );
  INV_X1 U21705 ( .A(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n18465) );
  OAI22_X1 U21706 ( .A1(n18466), .A2(n18594), .B1(n9786), .B2(n18465), .ZN(
        n18470) );
  AOI22_X1 U21707 ( .A1(n17547), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11911), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n18468) );
  AOI22_X1 U21708 ( .A1(n9724), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n14232), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n18467) );
  NAND2_X1 U21709 ( .A1(n18468), .A2(n18467), .ZN(n18469) );
  AOI211_X1 U21710 ( .C1(n18586), .C2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A(
        n18470), .B(n18469), .ZN(n18472) );
  AOI22_X1 U21711 ( .A1(n11937), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n18585), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n18471) );
  OAI211_X1 U21712 ( .C1(n9718), .C2(n18473), .A(n18472), .B(n18471), .ZN(
        n18480) );
  INV_X1 U21713 ( .A(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n18475) );
  OAI22_X1 U21714 ( .A1(n18551), .A2(n18475), .B1(n18525), .B2(n18474), .ZN(
        n18479) );
  OAI22_X1 U21715 ( .A1(n10660), .A2(n18598), .B1(n11951), .B2(n9723), .ZN(
        n18478) );
  INV_X1 U21716 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n18662) );
  OAI22_X1 U21717 ( .A1(n9783), .A2(n18476), .B1(n18599), .B2(n18662), .ZN(
        n18477) );
  NOR4_X1 U21718 ( .A1(n18480), .A2(n18479), .A3(n18478), .A4(n18477), .ZN(
        n18753) );
  INV_X1 U21719 ( .A(n18504), .ZN(n18482) );
  OAI211_X1 U21720 ( .C1(P3_EBX_REG_17__SCAN_IN), .C2(n18482), .A(n18481), .B(
        n18661), .ZN(n18483) );
  OAI21_X1 U21721 ( .B1(n18753), .B2(n18661), .A(n18483), .ZN(P3_U2686) );
  NAND2_X1 U21722 ( .A1(n9724), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n18484) );
  OAI21_X1 U21723 ( .B1(n18485), .B2(n18616), .A(n18484), .ZN(n18488) );
  OAI22_X1 U21724 ( .A1(n18613), .A2(n18486), .B1(n9723), .B2(n18609), .ZN(
        n18487) );
  NOR2_X1 U21725 ( .A1(n18488), .A2(n18487), .ZN(n18496) );
  AOI22_X1 U21726 ( .A1(n18586), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n18390), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n18495) );
  INV_X1 U21727 ( .A(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n22148) );
  NAND2_X1 U21728 ( .A1(n18620), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n18491) );
  NAND2_X1 U21729 ( .A1(n18489), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n18490) );
  OAI211_X1 U21730 ( .C1(n17550), .C2(n22148), .A(n18491), .B(n18490), .ZN(
        n18492) );
  INV_X1 U21731 ( .A(n18492), .ZN(n18494) );
  NAND2_X1 U21732 ( .A1(n18591), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n18493) );
  NAND4_X1 U21733 ( .A1(n18496), .A2(n18495), .A3(n18494), .A4(n18493), .ZN(
        n18503) );
  AOI22_X1 U21734 ( .A1(n18597), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n18627), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n18501) );
  AOI22_X1 U21735 ( .A1(n11911), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n14232), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n18500) );
  OR2_X1 U21736 ( .A1(n18599), .A2(n18497), .ZN(n18499) );
  NAND2_X1 U21737 ( .A1(n9726), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n18498) );
  NAND4_X1 U21738 ( .A1(n18501), .A2(n18500), .A3(n18499), .A4(n18498), .ZN(
        n18502) );
  NOR2_X1 U21739 ( .A1(n18503), .A2(n18502), .ZN(n18754) );
  OAI21_X1 U21740 ( .B1(P3_EBX_REG_16__SCAN_IN), .B2(n18520), .A(n18504), .ZN(
        n18505) );
  AOI22_X1 U21741 ( .A1(n18667), .A2(n18754), .B1(n18505), .B2(n18661), .ZN(
        P3_U2687) );
  OAI22_X1 U21742 ( .A1(n18611), .A2(n18506), .B1(n18525), .B2(n22079), .ZN(
        n18515) );
  AOI22_X1 U21743 ( .A1(n17547), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n9724), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n18513) );
  AOI22_X1 U21744 ( .A1(n18620), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n18619), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n18512) );
  INV_X1 U21745 ( .A(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n18507) );
  OAI22_X1 U21746 ( .A1(n18613), .A2(n11841), .B1(n9723), .B2(n18507), .ZN(
        n18508) );
  INV_X1 U21747 ( .A(n18508), .ZN(n18511) );
  INV_X1 U21748 ( .A(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n18509) );
  OR2_X1 U21749 ( .A1(n17550), .A2(n18509), .ZN(n18510) );
  NAND4_X1 U21750 ( .A1(n18513), .A2(n18512), .A3(n18511), .A4(n18510), .ZN(
        n18514) );
  AOI211_X1 U21751 ( .C1(n18591), .C2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A(
        n18515), .B(n18514), .ZN(n18519) );
  AOI22_X1 U21752 ( .A1(n11911), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n14232), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n18518) );
  AOI22_X1 U21753 ( .A1(n18626), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n18627), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n18517) );
  AOI22_X1 U21754 ( .A1(n18628), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n9726), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n18516) );
  NAND4_X1 U21755 ( .A1(n18519), .A2(n18518), .A3(n18517), .A4(n18516), .ZN(
        n18762) );
  AOI21_X1 U21756 ( .B1(n18522), .B2(n18521), .A(n18520), .ZN(n18523) );
  MUX2_X1 U21757 ( .A(n18762), .B(n18523), .S(n18661), .Z(P3_U2688) );
  INV_X1 U21758 ( .A(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n18526) );
  OAI22_X1 U21759 ( .A1(n18611), .A2(n18526), .B1(n18525), .B2(n18524), .ZN(
        n18535) );
  INV_X1 U21760 ( .A(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n18533) );
  OAI22_X1 U21761 ( .A1(n18613), .A2(n18527), .B1(n9723), .B2(n22036), .ZN(
        n18530) );
  NOR2_X1 U21762 ( .A1(n18556), .A2(n18528), .ZN(n18529) );
  AOI211_X1 U21763 ( .C1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .C2(n17547), .A(
        n18530), .B(n18529), .ZN(n18532) );
  AOI22_X1 U21764 ( .A1(n18620), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n18619), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n18531) );
  OAI211_X1 U21765 ( .C1(n17550), .C2(n18533), .A(n18532), .B(n18531), .ZN(
        n18534) );
  AOI211_X1 U21766 ( .C1(n18591), .C2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A(
        n18535), .B(n18534), .ZN(n18539) );
  AOI22_X1 U21767 ( .A1(n11911), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n14232), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n18538) );
  AOI22_X1 U21768 ( .A1(n18626), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n18627), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n18537) );
  AOI22_X1 U21769 ( .A1(n18628), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n9726), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n18536) );
  NAND4_X1 U21770 ( .A1(n18539), .A2(n18538), .A3(n18537), .A4(n18536), .ZN(
        n18766) );
  AOI22_X1 U21771 ( .A1(n18540), .A2(P3_EBX_REG_14__SCAN_IN), .B1(n18667), 
        .B2(n18766), .ZN(n18543) );
  NOR2_X1 U21772 ( .A1(n18765), .A2(n18582), .ZN(n18562) );
  NAND4_X1 U21773 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(P3_EBX_REG_12__SCAN_IN), 
        .A3(n18562), .A4(n18541), .ZN(n18542) );
  NAND2_X1 U21774 ( .A1(n18543), .A2(n18542), .ZN(P3_U2689) );
  AOI22_X1 U21775 ( .A1(n18585), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17547), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n18547) );
  AOI22_X1 U21776 ( .A1(n18620), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n18619), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n18546) );
  AOI22_X1 U21777 ( .A1(n14232), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17561), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n18545) );
  OR2_X1 U21778 ( .A1(n17550), .A2(n21977), .ZN(n18544) );
  AND4_X1 U21779 ( .A1(n18547), .A2(n18546), .A3(n18545), .A4(n18544), .ZN(
        n18549) );
  AOI22_X1 U21780 ( .A1(n18586), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11911), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n18548) );
  OAI211_X1 U21781 ( .C1(n18650), .C2(n9718), .A(n18549), .B(n18548), .ZN(
        n18560) );
  OAI22_X1 U21782 ( .A1(n18419), .A2(n18551), .B1(n18525), .B2(n18550), .ZN(
        n18559) );
  OAI22_X1 U21783 ( .A1(n9783), .A2(n18553), .B1(n18599), .B2(n18552), .ZN(
        n18558) );
  INV_X1 U21784 ( .A(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n18555) );
  OAI22_X1 U21785 ( .A1(n18556), .A2(n18555), .B1(n10660), .B2(n18554), .ZN(
        n18557) );
  NOR4_X1 U21786 ( .A1(n18560), .A2(n18559), .A3(n18558), .A4(n18557), .ZN(
        n18775) );
  AND2_X1 U21787 ( .A1(n18661), .A2(n18582), .ZN(n18563) );
  AOI22_X1 U21788 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n18563), .B1(n18562), 
        .B2(n18561), .ZN(n18564) );
  OAI21_X1 U21789 ( .B1(n18775), .B2(n18661), .A(n18564), .ZN(P3_U2691) );
  AOI22_X1 U21790 ( .A1(n17547), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n9724), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n18569) );
  AOI22_X1 U21791 ( .A1(n18620), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n18619), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n18568) );
  AOI22_X1 U21792 ( .A1(n11911), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17561), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n18567) );
  OR2_X1 U21793 ( .A1(n17550), .A2(n18565), .ZN(n18566) );
  AND4_X1 U21794 ( .A1(n18569), .A2(n18568), .A3(n18567), .A4(n18566), .ZN(
        n18571) );
  AOI22_X1 U21795 ( .A1(n18586), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n18597), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n18570) );
  OAI211_X1 U21796 ( .C1(n18654), .C2(n9718), .A(n18571), .B(n18570), .ZN(
        n18580) );
  OAI22_X1 U21797 ( .A1(n18525), .A2(n18572), .B1(n21980), .B2(n18615), .ZN(
        n18579) );
  OAI22_X1 U21798 ( .A1(n9783), .A2(n18574), .B1(n18599), .B2(n18573), .ZN(
        n18578) );
  OAI22_X1 U21799 ( .A1(n10660), .A2(n18576), .B1(n18613), .B2(n18575), .ZN(
        n18577) );
  NOR4_X1 U21800 ( .A1(n18580), .A2(n18579), .A3(n18578), .A4(n18577), .ZN(
        n18779) );
  NOR2_X1 U21801 ( .A1(n18581), .A2(n18642), .ZN(n18583) );
  OAI211_X1 U21802 ( .C1(P3_EBX_REG_11__SCAN_IN), .C2(n18583), .A(n18582), .B(
        n18661), .ZN(n18584) );
  OAI21_X1 U21803 ( .B1(n18779), .B2(n18661), .A(n18584), .ZN(P3_U2692) );
  AOI22_X1 U21804 ( .A1(n17547), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n9724), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n18590) );
  AOI22_X1 U21805 ( .A1(n18585), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11911), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n18589) );
  AOI22_X1 U21806 ( .A1(n18620), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n18619), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n18588) );
  NAND2_X1 U21807 ( .A1(n18586), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n18587) );
  NAND4_X1 U21808 ( .A1(n18590), .A2(n18589), .A3(n18588), .A4(n18587), .ZN(
        n18596) );
  NAND2_X1 U21809 ( .A1(n18591), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n18593) );
  NAND2_X1 U21810 ( .A1(n14232), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n18592) );
  OAI211_X1 U21811 ( .C1(n18594), .C2(n17550), .A(n18593), .B(n18592), .ZN(
        n18595) );
  OR2_X1 U21812 ( .A1(n18596), .A2(n18595), .ZN(n18605) );
  AOI22_X1 U21813 ( .A1(n18597), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n18390), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n18603) );
  AOI22_X1 U21814 ( .A1(n18627), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17561), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n18602) );
  OR2_X1 U21815 ( .A1(n18599), .A2(n18598), .ZN(n18601) );
  NAND2_X1 U21816 ( .A1(n9726), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n18600) );
  NAND4_X1 U21817 ( .A1(n18603), .A2(n18602), .A3(n18601), .A4(n18600), .ZN(
        n18604) );
  NOR2_X1 U21818 ( .A1(n18605), .A2(n18604), .ZN(n18792) );
  INV_X1 U21819 ( .A(n18606), .ZN(n18635) );
  OAI21_X1 U21820 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n18635), .A(n18661), .ZN(
        n18607) );
  OAI22_X1 U21821 ( .A1(n18792), .A2(n18661), .B1(n18608), .B2(n18607), .ZN(
        P3_U2694) );
  OAI22_X1 U21822 ( .A1(n18611), .A2(n18610), .B1(n11861), .B2(n18609), .ZN(
        n18625) );
  NOR2_X1 U21823 ( .A1(n18613), .A2(n18612), .ZN(n18618) );
  INV_X1 U21824 ( .A(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n18614) );
  OAI22_X1 U21825 ( .A1(n18616), .A2(n22148), .B1(n18615), .B2(n18614), .ZN(
        n18617) );
  AOI211_X1 U21826 ( .C1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .C2(n9724), .A(
        n18618), .B(n18617), .ZN(n18622) );
  AOI22_X1 U21827 ( .A1(n18620), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n18619), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n18621) );
  OAI211_X1 U21828 ( .C1(n17550), .C2(n18623), .A(n18622), .B(n18621), .ZN(
        n18624) );
  AOI211_X1 U21829 ( .C1(n18591), .C2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A(
        n18625), .B(n18624), .ZN(n18632) );
  AOI22_X1 U21830 ( .A1(n18626), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n18390), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n18631) );
  AOI22_X1 U21831 ( .A1(n18627), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17561), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n18630) );
  AOI22_X1 U21832 ( .A1(n18628), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n9726), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n18629) );
  AND4_X1 U21833 ( .A1(n18632), .A2(n18631), .A3(n18630), .A4(n18629), .ZN(
        n18800) );
  NOR2_X1 U21834 ( .A1(n18633), .A2(n18642), .ZN(n18639) );
  AOI22_X1 U21835 ( .A1(n19561), .A2(n18639), .B1(P3_EBX_REG_8__SCAN_IN), .B2(
        n18661), .ZN(n18634) );
  OAI22_X1 U21836 ( .A1(n18800), .A2(n18661), .B1(n18635), .B2(n18634), .ZN(
        P3_U2695) );
  OAI21_X1 U21837 ( .B1(P3_EBX_REG_7__SCAN_IN), .B2(n18636), .A(n18661), .ZN(
        n18638) );
  OAI22_X1 U21838 ( .A1(n18639), .A2(n18638), .B1(n18637), .B2(n18661), .ZN(
        P3_U2696) );
  NOR2_X1 U21839 ( .A1(n18641), .A2(n18640), .ZN(n18647) );
  OAI21_X1 U21840 ( .B1(P3_EBX_REG_6__SCAN_IN), .B2(n18647), .A(n18642), .ZN(
        n18643) );
  AOI22_X1 U21841 ( .A1(n18667), .A2(n18644), .B1(n18643), .B2(n18661), .ZN(
        P3_U2697) );
  OAI21_X1 U21842 ( .B1(P3_EBX_REG_5__SCAN_IN), .B2(n18652), .A(n18661), .ZN(
        n18646) );
  OAI22_X1 U21843 ( .A1(n18647), .A2(n18646), .B1(n18645), .B2(n18661), .ZN(
        P3_U2698) );
  INV_X1 U21844 ( .A(n18664), .ZN(n18666) );
  NAND2_X1 U21845 ( .A1(n18648), .A2(n18666), .ZN(n18653) );
  NOR2_X1 U21846 ( .A1(n18649), .A2(n18653), .ZN(n18656) );
  AOI21_X1 U21847 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n18661), .A(n18656), .ZN(
        n18651) );
  OAI22_X1 U21848 ( .A1(n18652), .A2(n18651), .B1(n18650), .B2(n18661), .ZN(
        P3_U2699) );
  INV_X1 U21849 ( .A(n18653), .ZN(n18658) );
  AOI21_X1 U21850 ( .B1(P3_EBX_REG_3__SCAN_IN), .B2(n18661), .A(n18658), .ZN(
        n18655) );
  OAI22_X1 U21851 ( .A1(n18656), .A2(n18655), .B1(n18654), .B2(n18661), .ZN(
        P3_U2700) );
  AOI211_X1 U21852 ( .C1(n18667), .C2(n18660), .A(n18659), .B(n18658), .ZN(
        P3_U2701) );
  OAI222_X1 U21853 ( .A1(n18665), .A2(n18664), .B1(n18663), .B2(n18670), .C1(
        n18662), .C2(n18661), .ZN(P3_U2702) );
  AOI22_X1 U21854 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18667), .B1(
        n18666), .B2(n18669), .ZN(n18668) );
  OAI21_X1 U21855 ( .B1(n18670), .B2(n18669), .A(n18668), .ZN(P3_U2703) );
  NOR2_X2 U21856 ( .A1(n18810), .A2(n19555), .ZN(n18756) );
  INV_X1 U21857 ( .A(n18756), .ZN(n18700) );
  NAND4_X1 U21858 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(P3_EAX_REG_4__SCAN_IN), 
        .A3(P3_EAX_REG_3__SCAN_IN), .A4(P3_EAX_REG_2__SCAN_IN), .ZN(n18671) );
  INV_X1 U21859 ( .A(n18797), .ZN(n18676) );
  NAND4_X1 U21860 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(P3_EAX_REG_11__SCAN_IN), 
        .A3(P3_EAX_REG_10__SCAN_IN), .A4(P3_EAX_REG_9__SCAN_IN), .ZN(n18674)
         );
  NAND3_X1 U21861 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(P3_EAX_REG_8__SCAN_IN), 
        .A3(P3_EAX_REG_14__SCAN_IN), .ZN(n18673) );
  NAND2_X1 U21862 ( .A1(P3_EAX_REG_17__SCAN_IN), .A2(P3_EAX_REG_18__SCAN_IN), 
        .ZN(n18723) );
  NAND2_X1 U21863 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(P3_EAX_REG_20__SCAN_IN), 
        .ZN(n18725) );
  NAND3_X1 U21864 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(P3_EAX_REG_19__SCAN_IN), 
        .A3(n18677), .ZN(n18716) );
  NAND2_X1 U21865 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n18696), .ZN(n18691) );
  INV_X1 U21866 ( .A(n18691), .ZN(n18688) );
  NAND2_X1 U21867 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n18688), .ZN(n18687) );
  NOR2_X1 U21868 ( .A1(P3_EAX_REG_31__SCAN_IN), .A2(n18687), .ZN(n18678) );
  INV_X1 U21869 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n18885) );
  INV_X1 U21870 ( .A(n18680), .ZN(n19551) );
  OAI22_X1 U21871 ( .A1(n18682), .A2(n18812), .B1(n18681), .B2(n18700), .ZN(
        n18683) );
  AOI21_X1 U21872 ( .B1(BUF2_REG_14__SCAN_IN), .B2(n18748), .A(n18683), .ZN(
        n18684) );
  OAI221_X1 U21873 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n18687), .C1(n18885), 
        .C2(n18685), .A(n18684), .ZN(P3_U2705) );
  INV_X1 U21874 ( .A(BUF2_REG_29__SCAN_IN), .ZN(n22049) );
  AOI22_X1 U21875 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n18748), .B1(n18785), .B2(
        n18686), .ZN(n18690) );
  OAI211_X1 U21876 ( .C1(n18688), .C2(P3_EAX_REG_29__SCAN_IN), .A(n18810), .B(
        n18687), .ZN(n18689) );
  OAI211_X1 U21877 ( .C1(n18700), .C2(n22049), .A(n18690), .B(n18689), .ZN(
        P3_U2706) );
  AOI22_X1 U21878 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n18748), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n18756), .ZN(n18693) );
  OAI211_X1 U21879 ( .C1(n18696), .C2(P3_EAX_REG_28__SCAN_IN), .A(n18810), .B(
        n18691), .ZN(n18692) );
  OAI211_X1 U21880 ( .C1(n18694), .C2(n18812), .A(n18693), .B(n18692), .ZN(
        P3_U2707) );
  AOI22_X1 U21881 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n18748), .B1(n18785), .B2(
        n18695), .ZN(n18699) );
  AOI211_X1 U21882 ( .C1(n22041), .C2(n18701), .A(n18696), .B(n18784), .ZN(
        n18697) );
  INV_X1 U21883 ( .A(n18697), .ZN(n18698) );
  OAI211_X1 U21884 ( .C1(n18700), .C2(n22056), .A(n18699), .B(n18698), .ZN(
        P3_U2708) );
  AOI22_X1 U21885 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n18748), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n18756), .ZN(n18703) );
  OAI211_X1 U21886 ( .C1(n9852), .C2(P3_EAX_REG_26__SCAN_IN), .A(n18810), .B(
        n18701), .ZN(n18702) );
  OAI211_X1 U21887 ( .C1(n18704), .C2(n18812), .A(n18703), .B(n18702), .ZN(
        P3_U2709) );
  AOI22_X1 U21888 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n18756), .B1(n18785), .B2(
        n18705), .ZN(n18708) );
  AOI211_X1 U21889 ( .C1(n18877), .C2(n18710), .A(n9852), .B(n18784), .ZN(
        n18706) );
  INV_X1 U21890 ( .A(n18706), .ZN(n18707) );
  OAI211_X1 U21891 ( .C1(n18760), .C2(n18795), .A(n18708), .B(n18707), .ZN(
        P3_U2710) );
  AOI22_X1 U21892 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n18748), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n18756), .ZN(n18713) );
  OAI21_X1 U21893 ( .B1(n18875), .B2(n18784), .A(n18709), .ZN(n18711) );
  NAND2_X1 U21894 ( .A1(n18711), .A2(n18710), .ZN(n18712) );
  OAI211_X1 U21895 ( .C1(n18714), .C2(n18812), .A(n18713), .B(n18712), .ZN(
        P3_U2711) );
  AOI211_X1 U21896 ( .C1(n18873), .C2(n18716), .A(n18784), .B(n18715), .ZN(
        n18719) );
  OAI22_X1 U21897 ( .A1(n19558), .A2(n18760), .B1(n18812), .B2(n18717), .ZN(
        n18718) );
  AOI211_X1 U21898 ( .C1(n18756), .C2(BUF2_REG_23__SCAN_IN), .A(n18719), .B(
        n18718), .ZN(n18720) );
  INV_X1 U21899 ( .A(n18720), .ZN(P3_U2712) );
  INV_X1 U21900 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n19554) );
  INV_X1 U21901 ( .A(n18721), .ZN(n18722) );
  AOI22_X1 U21902 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n18756), .B1(n18785), .B2(
        n18722), .ZN(n18729) );
  INV_X1 U21903 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n18867) );
  NAND2_X1 U21904 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n18744), .ZN(n18739) );
  OR2_X1 U21905 ( .A1(n18867), .A2(n18739), .ZN(n18734) );
  NAND2_X1 U21906 ( .A1(n18810), .A2(n18734), .ZN(n18731) );
  OAI21_X1 U21907 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n18724), .A(n18731), .ZN(
        n18727) );
  NOR3_X1 U21908 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n18725), .A3(n18739), .ZN(
        n18726) );
  AOI21_X1 U21909 ( .B1(P3_EAX_REG_22__SCAN_IN), .B2(n18727), .A(n18726), .ZN(
        n18728) );
  OAI211_X1 U21910 ( .C1(n19554), .C2(n18760), .A(n18729), .B(n18728), .ZN(
        P3_U2713) );
  AOI22_X1 U21911 ( .A1(BUF2_REG_21__SCAN_IN), .A2(n18756), .B1(n18785), .B2(
        n18730), .ZN(n18733) );
  INV_X1 U21912 ( .A(n18731), .ZN(n18736) );
  AOI22_X1 U21913 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n18748), .B1(
        P3_EAX_REG_21__SCAN_IN), .B2(n18736), .ZN(n18732) );
  OAI211_X1 U21914 ( .C1(P3_EAX_REG_21__SCAN_IN), .C2(n18734), .A(n18733), .B(
        n18732), .ZN(P3_U2714) );
  AOI22_X1 U21915 ( .A1(BUF2_REG_20__SCAN_IN), .A2(n18756), .B1(n18785), .B2(
        n18735), .ZN(n18738) );
  AOI22_X1 U21916 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n18748), .B1(
        P3_EAX_REG_20__SCAN_IN), .B2(n18736), .ZN(n18737) );
  OAI211_X1 U21917 ( .C1(P3_EAX_REG_20__SCAN_IN), .C2(n18739), .A(n18738), .B(
        n18737), .ZN(P3_U2715) );
  AOI22_X1 U21918 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n18748), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n18756), .ZN(n18741) );
  OAI211_X1 U21919 ( .C1(n18744), .C2(P3_EAX_REG_19__SCAN_IN), .A(n18810), .B(
        n18739), .ZN(n18740) );
  OAI211_X1 U21920 ( .C1(n18742), .C2(n18812), .A(n18741), .B(n18740), .ZN(
        P3_U2716) );
  INV_X1 U21921 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n19538) );
  AOI22_X1 U21922 ( .A1(BUF2_REG_18__SCAN_IN), .A2(n18756), .B1(n18785), .B2(
        n18743), .ZN(n18747) );
  INV_X1 U21923 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n18863) );
  INV_X1 U21924 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n22200) );
  OR2_X1 U21925 ( .A1(n18757), .A2(n22200), .ZN(n18749) );
  AOI211_X1 U21926 ( .C1(n18863), .C2(n18749), .A(n18744), .B(n18784), .ZN(
        n18745) );
  INV_X1 U21927 ( .A(n18745), .ZN(n18746) );
  OAI211_X1 U21928 ( .C1(n18760), .C2(n19538), .A(n18747), .B(n18746), .ZN(
        P3_U2717) );
  AOI22_X1 U21929 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n18748), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n18756), .ZN(n18752) );
  INV_X1 U21930 ( .A(n18757), .ZN(n18750) );
  OAI211_X1 U21931 ( .C1(n18750), .C2(P3_EAX_REG_17__SCAN_IN), .A(n18810), .B(
        n18749), .ZN(n18751) );
  OAI211_X1 U21932 ( .C1(n18753), .C2(n18812), .A(n18752), .B(n18751), .ZN(
        P3_U2718) );
  INV_X1 U21933 ( .A(n18754), .ZN(n18755) );
  AOI22_X1 U21934 ( .A1(BUF2_REG_16__SCAN_IN), .A2(n18756), .B1(n18785), .B2(
        n18755), .ZN(n18759) );
  OAI211_X1 U21935 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n9875), .A(n18810), .B(
        n18757), .ZN(n18758) );
  OAI211_X1 U21936 ( .C1(n18760), .C2(n22011), .A(n18759), .B(n18758), .ZN(
        P3_U2719) );
  OR2_X1 U21937 ( .A1(n18765), .A2(n18761), .ZN(n18764) );
  NAND2_X1 U21938 ( .A1(n18810), .A2(n18761), .ZN(n18768) );
  AOI22_X1 U21939 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n18796), .B1(n18785), .B2(
        n18762), .ZN(n18763) );
  OAI221_X1 U21940 ( .B1(P3_EAX_REG_15__SCAN_IN), .B2(n18764), .C1(n18920), 
        .C2(n18768), .A(n18763), .ZN(P3_U2720) );
  INV_X1 U21941 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n22098) );
  INV_X1 U21942 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n18908) );
  NOR2_X1 U21943 ( .A1(n18765), .A2(n18797), .ZN(n18804) );
  NAND3_X1 U21944 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(P3_EAX_REG_8__SCAN_IN), 
        .A3(n18804), .ZN(n18791) );
  NAND2_X1 U21945 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(n18783), .ZN(n18774) );
  NAND2_X1 U21946 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n18777), .ZN(n18769) );
  INV_X1 U21947 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n18916) );
  AOI22_X1 U21948 ( .A1(n18766), .A2(n18785), .B1(BUF2_REG_14__SCAN_IN), .B2(
        n18796), .ZN(n18767) );
  OAI221_X1 U21949 ( .B1(P3_EAX_REG_14__SCAN_IN), .B2(n18769), .C1(n18916), 
        .C2(n18768), .A(n18767), .ZN(P3_U2721) );
  INV_X1 U21950 ( .A(n18769), .ZN(n18772) );
  AOI21_X1 U21951 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n18810), .A(n18777), .ZN(
        n18771) );
  OAI222_X1 U21952 ( .A1(n18815), .A2(n18773), .B1(n18772), .B2(n18771), .C1(
        n18812), .C2(n18770), .ZN(P3_U2722) );
  INV_X1 U21953 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n18778) );
  INV_X1 U21954 ( .A(n18774), .ZN(n18781) );
  AOI21_X1 U21955 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n18810), .A(n18781), .ZN(
        n18776) );
  OAI222_X1 U21956 ( .A1(n18815), .A2(n18778), .B1(n18777), .B2(n18776), .C1(
        n18812), .C2(n18775), .ZN(P3_U2723) );
  AOI21_X1 U21957 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n18810), .A(n18783), .ZN(
        n18780) );
  OAI222_X1 U21958 ( .A1(n18815), .A2(n18782), .B1(n18781), .B2(n18780), .C1(
        n18812), .C2(n18779), .ZN(P3_U2724) );
  INV_X1 U21959 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n18790) );
  AOI211_X1 U21960 ( .C1(n18908), .C2(n18791), .A(n18784), .B(n18783), .ZN(
        n18788) );
  AND2_X1 U21961 ( .A1(n18786), .A2(n18785), .ZN(n18787) );
  NOR2_X1 U21962 ( .A1(n18788), .A2(n18787), .ZN(n18789) );
  OAI21_X1 U21963 ( .B1(n18790), .B2(n18815), .A(n18789), .ZN(P3_U2725) );
  INV_X1 U21964 ( .A(n18791), .ZN(n18794) );
  AOI22_X1 U21965 ( .A1(n18804), .A2(P3_EAX_REG_8__SCAN_IN), .B1(
        P3_EAX_REG_9__SCAN_IN), .B2(n18810), .ZN(n18793) );
  OAI222_X1 U21966 ( .A1(n18815), .A2(n18795), .B1(n18794), .B2(n18793), .C1(
        n18812), .C2(n18792), .ZN(P3_U2726) );
  INV_X1 U21967 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n18904) );
  AOI22_X1 U21968 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n18796), .B1(n18804), .B2(
        n18904), .ZN(n18799) );
  NAND3_X1 U21969 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n18810), .A3(n18797), .ZN(
        n18798) );
  OAI211_X1 U21970 ( .C1(n18800), .C2(n18812), .A(n18799), .B(n18798), .ZN(
        P3_U2727) );
  AOI21_X1 U21971 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n18810), .A(n18801), .ZN(
        n18803) );
  OAI222_X1 U21972 ( .A1(n19558), .A2(n18815), .B1(n18804), .B2(n18803), .C1(
        n18812), .C2(n18802), .ZN(P3_U2728) );
  AOI21_X1 U21973 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n18810), .A(n18805), .ZN(
        n18807) );
  OAI222_X1 U21974 ( .A1(n19550), .A2(n18815), .B1(n18808), .B2(n18807), .C1(
        n18812), .C2(n18806), .ZN(P3_U2730) );
  INV_X1 U21975 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n19542) );
  AOI21_X1 U21976 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n18810), .A(n18809), .ZN(
        n18813) );
  OAI222_X1 U21977 ( .A1(n19542), .A2(n18815), .B1(n18814), .B2(n18813), .C1(
        n18812), .C2(n18811), .ZN(P3_U2732) );
  NAND2_X1 U21978 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n19113), .ZN(n18854) );
  NOR2_X1 U21979 ( .A1(n18853), .A2(n18817), .ZN(P3_U2736) );
  INV_X2 U21980 ( .A(n18854), .ZN(n18851) );
  AOI22_X1 U21981 ( .A1(n18851), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n18850), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n18819) );
  OAI21_X1 U21982 ( .B1(n18885), .B2(n18834), .A(n18819), .ZN(P3_U2737) );
  INV_X1 U21983 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n18883) );
  AOI22_X1 U21984 ( .A1(n18851), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n18850), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n18820) );
  OAI21_X1 U21985 ( .B1(n18883), .B2(n18834), .A(n18820), .ZN(P3_U2738) );
  INV_X1 U21986 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n18881) );
  AOI22_X1 U21987 ( .A1(n18851), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n18850), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n18821) );
  OAI21_X1 U21988 ( .B1(n18881), .B2(n18834), .A(n18821), .ZN(P3_U2739) );
  AOI22_X1 U21989 ( .A1(n18851), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n18850), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n18822) );
  OAI21_X1 U21990 ( .B1(n22041), .B2(n18834), .A(n18822), .ZN(P3_U2740) );
  AOI22_X1 U21991 ( .A1(n18851), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n18850), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n18823) );
  OAI21_X1 U21992 ( .B1(n10256), .B2(n18834), .A(n18823), .ZN(P3_U2741) );
  AOI22_X1 U21993 ( .A1(n18851), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n18850), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n18824) );
  OAI21_X1 U21994 ( .B1(n18877), .B2(n18834), .A(n18824), .ZN(P3_U2742) );
  AOI22_X1 U21995 ( .A1(n18851), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n18850), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n18825) );
  OAI21_X1 U21996 ( .B1(n18875), .B2(n18834), .A(n18825), .ZN(P3_U2743) );
  AOI22_X1 U21997 ( .A1(n18851), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n18850), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n18826) );
  OAI21_X1 U21998 ( .B1(n18873), .B2(n18834), .A(n18826), .ZN(P3_U2744) );
  INV_X1 U21999 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n18871) );
  AOI22_X1 U22000 ( .A1(n18851), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n18850), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n18827) );
  OAI21_X1 U22001 ( .B1(n18871), .B2(n18834), .A(n18827), .ZN(P3_U2745) );
  INV_X1 U22002 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n18869) );
  AOI22_X1 U22003 ( .A1(n18851), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n18850), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n18828) );
  OAI21_X1 U22004 ( .B1(n18869), .B2(n18834), .A(n18828), .ZN(P3_U2746) );
  AOI22_X1 U22005 ( .A1(n18851), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n18850), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n18829) );
  OAI21_X1 U22006 ( .B1(n18867), .B2(n18834), .A(n18829), .ZN(P3_U2747) );
  INV_X1 U22007 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n18865) );
  AOI22_X1 U22008 ( .A1(n18851), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n18850), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n18830) );
  OAI21_X1 U22009 ( .B1(n18865), .B2(n18834), .A(n18830), .ZN(P3_U2748) );
  AOI22_X1 U22010 ( .A1(n18851), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n18850), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n18831) );
  OAI21_X1 U22011 ( .B1(n18863), .B2(n18834), .A(n18831), .ZN(P3_U2749) );
  AOI22_X1 U22012 ( .A1(n18851), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n18850), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n18832) );
  OAI21_X1 U22013 ( .B1(n22200), .B2(n18834), .A(n18832), .ZN(P3_U2750) );
  INV_X1 U22014 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n18860) );
  AOI22_X1 U22015 ( .A1(n18851), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n18850), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n18833) );
  OAI21_X1 U22016 ( .B1(n18860), .B2(n18834), .A(n18833), .ZN(P3_U2751) );
  AOI22_X1 U22017 ( .A1(n18851), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n18850), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n18835) );
  OAI21_X1 U22018 ( .B1(n18920), .B2(n18855), .A(n18835), .ZN(P3_U2752) );
  AOI22_X1 U22019 ( .A1(n18851), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n18850), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n18836) );
  OAI21_X1 U22020 ( .B1(n18916), .B2(n18855), .A(n18836), .ZN(P3_U2753) );
  INV_X1 U22021 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n18914) );
  AOI22_X1 U22022 ( .A1(n18851), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n18850), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n18837) );
  OAI21_X1 U22023 ( .B1(n18914), .B2(n18855), .A(n18837), .ZN(P3_U2754) );
  AOI22_X1 U22024 ( .A1(n18851), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n18850), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n18838) );
  OAI21_X1 U22025 ( .B1(n22098), .B2(n18855), .A(n18838), .ZN(P3_U2755) );
  INV_X1 U22026 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n18910) );
  AOI22_X1 U22027 ( .A1(n18851), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n18850), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n18839) );
  OAI21_X1 U22028 ( .B1(n18910), .B2(n18855), .A(n18839), .ZN(P3_U2756) );
  AOI22_X1 U22029 ( .A1(P3_DATAO_REG_10__SCAN_IN), .A2(n18850), .B1(n18851), 
        .B2(P3_LWORD_REG_10__SCAN_IN), .ZN(n18840) );
  OAI21_X1 U22030 ( .B1(n18908), .B2(n18855), .A(n18840), .ZN(P3_U2757) );
  INV_X1 U22031 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n18906) );
  AOI22_X1 U22032 ( .A1(n18851), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n18850), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n18841) );
  OAI21_X1 U22033 ( .B1(n18906), .B2(n18855), .A(n18841), .ZN(P3_U2758) );
  AOI22_X1 U22034 ( .A1(n18851), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n18850), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n18842) );
  OAI21_X1 U22035 ( .B1(n18904), .B2(n18855), .A(n18842), .ZN(P3_U2759) );
  INV_X1 U22036 ( .A(P3_LWORD_REG_7__SCAN_IN), .ZN(n22082) );
  AOI22_X1 U22037 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(n18843), .B1(n18850), .B2(
        P3_DATAO_REG_7__SCAN_IN), .ZN(n18844) );
  OAI21_X1 U22038 ( .B1(n22082), .B2(n18854), .A(n18844), .ZN(P3_U2760) );
  AOI22_X1 U22039 ( .A1(n18851), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n18850), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n18845) );
  OAI21_X1 U22040 ( .B1(n18899), .B2(n18855), .A(n18845), .ZN(P3_U2761) );
  INV_X1 U22041 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n18897) );
  AOI22_X1 U22042 ( .A1(n18851), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n18850), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n18846) );
  OAI21_X1 U22043 ( .B1(n18897), .B2(n18855), .A(n18846), .ZN(P3_U2762) );
  AOI22_X1 U22044 ( .A1(n18851), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n18850), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n18847) );
  OAI21_X1 U22045 ( .B1(n18895), .B2(n18855), .A(n18847), .ZN(P3_U2763) );
  INV_X1 U22046 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n18893) );
  AOI22_X1 U22047 ( .A1(n18851), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n18850), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n18848) );
  OAI21_X1 U22048 ( .B1(n18893), .B2(n18855), .A(n18848), .ZN(P3_U2764) );
  INV_X1 U22049 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n18891) );
  AOI22_X1 U22050 ( .A1(n18851), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n18850), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n18849) );
  OAI21_X1 U22051 ( .B1(n18891), .B2(n18855), .A(n18849), .ZN(P3_U2765) );
  AOI22_X1 U22052 ( .A1(n18851), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n18850), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n18852) );
  OAI21_X1 U22053 ( .B1(n18889), .B2(n18855), .A(n18852), .ZN(P3_U2766) );
  INV_X1 U22054 ( .A(P3_LWORD_REG_0__SCAN_IN), .ZN(n22201) );
  INV_X1 U22055 ( .A(P3_DATAO_REG_0__SCAN_IN), .ZN(n22120) );
  OAI222_X1 U22056 ( .A1(n18855), .A2(n18887), .B1(n18854), .B2(n22201), .C1(
        n22120), .C2(n18853), .ZN(P3_U2767) );
  INV_X1 U22057 ( .A(n18856), .ZN(n20035) );
  NOR2_X4 U22058 ( .A1(n19535), .A2(n18917), .ZN(n18911) );
  AOI22_X1 U22059 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n18911), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n18917), .ZN(n18859) );
  OAI21_X1 U22060 ( .B1(n18860), .B2(n18919), .A(n18859), .ZN(P3_U2768) );
  AOI22_X1 U22061 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n18911), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n18917), .ZN(n18861) );
  OAI21_X1 U22062 ( .B1(n22200), .B2(n18919), .A(n18861), .ZN(P3_U2769) );
  AOI22_X1 U22063 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n18911), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n18917), .ZN(n18862) );
  OAI21_X1 U22064 ( .B1(n18863), .B2(n18919), .A(n18862), .ZN(P3_U2770) );
  AOI22_X1 U22065 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n18911), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n18917), .ZN(n18864) );
  OAI21_X1 U22066 ( .B1(n18865), .B2(n18919), .A(n18864), .ZN(P3_U2771) );
  AOI22_X1 U22067 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n18911), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n18917), .ZN(n18866) );
  OAI21_X1 U22068 ( .B1(n18867), .B2(n18919), .A(n18866), .ZN(P3_U2772) );
  AOI22_X1 U22069 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n18911), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n18917), .ZN(n18868) );
  OAI21_X1 U22070 ( .B1(n18869), .B2(n18919), .A(n18868), .ZN(P3_U2773) );
  AOI22_X1 U22071 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n18911), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n18917), .ZN(n18870) );
  OAI21_X1 U22072 ( .B1(n18871), .B2(n18919), .A(n18870), .ZN(P3_U2774) );
  AOI22_X1 U22073 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n18911), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n18917), .ZN(n18872) );
  OAI21_X1 U22074 ( .B1(n18873), .B2(n18919), .A(n18872), .ZN(P3_U2775) );
  AOI22_X1 U22075 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n18911), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n18917), .ZN(n18874) );
  OAI21_X1 U22076 ( .B1(n18875), .B2(n18919), .A(n18874), .ZN(P3_U2776) );
  AOI22_X1 U22077 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n18911), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n18917), .ZN(n18876) );
  OAI21_X1 U22078 ( .B1(n18877), .B2(n18919), .A(n18876), .ZN(P3_U2777) );
  AOI22_X1 U22079 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n18911), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n18917), .ZN(n18878) );
  OAI21_X1 U22080 ( .B1(n10256), .B2(n18919), .A(n18878), .ZN(P3_U2778) );
  AOI22_X1 U22081 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n18911), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n18917), .ZN(n18879) );
  OAI21_X1 U22082 ( .B1(n22041), .B2(n18919), .A(n18879), .ZN(P3_U2779) );
  AOI22_X1 U22083 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n18911), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n18917), .ZN(n18880) );
  OAI21_X1 U22084 ( .B1(n18881), .B2(n18919), .A(n18880), .ZN(P3_U2780) );
  AOI22_X1 U22085 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n18911), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n18917), .ZN(n18882) );
  OAI21_X1 U22086 ( .B1(n18883), .B2(n18919), .A(n18882), .ZN(P3_U2781) );
  AOI22_X1 U22087 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n18911), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n18917), .ZN(n18884) );
  OAI21_X1 U22088 ( .B1(n18885), .B2(n18919), .A(n18884), .ZN(P3_U2782) );
  AOI22_X1 U22089 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n18911), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n18917), .ZN(n18886) );
  OAI21_X1 U22090 ( .B1(n18887), .B2(n18919), .A(n18886), .ZN(P3_U2783) );
  AOI22_X1 U22091 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n18911), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n18917), .ZN(n18888) );
  OAI21_X1 U22092 ( .B1(n18889), .B2(n18919), .A(n18888), .ZN(P3_U2784) );
  AOI22_X1 U22093 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n18911), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n18917), .ZN(n18890) );
  OAI21_X1 U22094 ( .B1(n18891), .B2(n18919), .A(n18890), .ZN(P3_U2785) );
  AOI22_X1 U22095 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n18911), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n18917), .ZN(n18892) );
  OAI21_X1 U22096 ( .B1(n18893), .B2(n18919), .A(n18892), .ZN(P3_U2786) );
  AOI22_X1 U22097 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n18911), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n18917), .ZN(n18894) );
  OAI21_X1 U22098 ( .B1(n18895), .B2(n18919), .A(n18894), .ZN(P3_U2787) );
  AOI22_X1 U22099 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n18911), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n18917), .ZN(n18896) );
  OAI21_X1 U22100 ( .B1(n18897), .B2(n18919), .A(n18896), .ZN(P3_U2788) );
  AOI22_X1 U22101 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n18911), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n18917), .ZN(n18898) );
  OAI21_X1 U22102 ( .B1(n18899), .B2(n18919), .A(n18898), .ZN(P3_U2789) );
  AOI22_X1 U22103 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n18911), .B1(
        P3_EAX_REG_7__SCAN_IN), .B2(n18900), .ZN(n18901) );
  OAI21_X1 U22104 ( .B1(n18902), .B2(n22082), .A(n18901), .ZN(P3_U2790) );
  AOI22_X1 U22105 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n18911), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n18917), .ZN(n18903) );
  OAI21_X1 U22106 ( .B1(n18904), .B2(n18919), .A(n18903), .ZN(P3_U2791) );
  AOI22_X1 U22107 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n18911), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n18917), .ZN(n18905) );
  OAI21_X1 U22108 ( .B1(n18906), .B2(n18919), .A(n18905), .ZN(P3_U2792) );
  AOI22_X1 U22109 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n18911), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n18917), .ZN(n18907) );
  OAI21_X1 U22110 ( .B1(n18908), .B2(n18919), .A(n18907), .ZN(P3_U2793) );
  AOI22_X1 U22111 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n18911), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n18917), .ZN(n18909) );
  OAI21_X1 U22112 ( .B1(n18910), .B2(n18919), .A(n18909), .ZN(P3_U2794) );
  AOI22_X1 U22113 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n18911), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n18917), .ZN(n18912) );
  OAI21_X1 U22114 ( .B1(n22098), .B2(n18919), .A(n18912), .ZN(P3_U2795) );
  AOI22_X1 U22115 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n18911), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n18917), .ZN(n18913) );
  OAI21_X1 U22116 ( .B1(n18914), .B2(n18919), .A(n18913), .ZN(P3_U2796) );
  AOI22_X1 U22117 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n18911), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n18917), .ZN(n18915) );
  OAI21_X1 U22118 ( .B1(n18916), .B2(n18919), .A(n18915), .ZN(P3_U2797) );
  AOI22_X1 U22119 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n18911), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n18917), .ZN(n18918) );
  OAI21_X1 U22120 ( .B1(n18920), .B2(n18919), .A(n18918), .ZN(P3_U2798) );
  NAND2_X1 U22121 ( .A1(n18921), .A2(n21976), .ZN(n18936) );
  OAI21_X1 U22122 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n18996), .A(
        n18922), .ZN(n18938) );
  NOR2_X1 U22123 ( .A1(n19145), .A2(n10167), .ZN(n19019) );
  NOR2_X1 U22124 ( .A1(n19259), .A2(n18946), .ZN(n18923) );
  NOR3_X1 U22125 ( .A1(n19019), .A2(n18923), .A3(n21976), .ZN(n18930) );
  NOR2_X1 U22126 ( .A1(n19026), .A2(n18924), .ZN(n18944) );
  OAI211_X1 U22127 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(n18944), .B(n18925), .ZN(n18927) );
  OAI211_X1 U22128 ( .C1(n19118), .C2(n18928), .A(n18927), .B(n18926), .ZN(
        n18929) );
  AOI211_X1 U22129 ( .C1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .C2(n18938), .A(
        n18930), .B(n18929), .ZN(n18935) );
  XOR2_X1 U22130 ( .A(n18932), .B(n18931), .Z(n18933) );
  NAND2_X1 U22131 ( .A1(n18933), .A2(n19172), .ZN(n18934) );
  OAI211_X1 U22132 ( .C1(n18989), .C2(n18936), .A(n18935), .B(n18934), .ZN(
        P3_U2802) );
  AOI22_X1 U22133 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n18938), .B1(
        n19128), .B2(n18937), .ZN(n18949) );
  OAI21_X1 U22134 ( .B1(n18939), .B2(n18942), .A(n19185), .ZN(n18940) );
  OAI21_X1 U22135 ( .B1(n18942), .B2(n18941), .A(n18940), .ZN(n19255) );
  AOI22_X1 U22136 ( .A1(n19172), .A2(n19255), .B1(n18944), .B2(n18943), .ZN(
        n18948) );
  NOR2_X1 U22137 ( .A1(n19250), .A2(n18989), .ZN(n18945) );
  AOI22_X1 U22138 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18946), .B1(
        n18945), .B2(n19259), .ZN(n18947) );
  NAND2_X1 U22139 ( .A1(n19508), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n19257) );
  NAND4_X1 U22140 ( .A1(n18949), .A2(n18948), .A3(n18947), .A4(n19257), .ZN(
        P3_U2803) );
  XOR2_X1 U22141 ( .A(n18950), .B(n19263), .Z(n19268) );
  OAI21_X1 U22142 ( .B1(n18951), .B2(n19068), .A(n19207), .ZN(n18952) );
  AOI21_X1 U22143 ( .B1(n19921), .B2(n11799), .A(n18952), .ZN(n18983) );
  OAI21_X1 U22144 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n18996), .A(
        n18983), .ZN(n18965) );
  NOR2_X1 U22145 ( .A1(n19026), .A2(n11799), .ZN(n18967) );
  OAI211_X1 U22146 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n18967), .B(n18953), .ZN(n18954) );
  NAND2_X1 U22147 ( .A1(n19508), .A2(P3_REIP_REG_25__SCAN_IN), .ZN(n19270) );
  OAI211_X1 U22148 ( .C1(n19118), .C2(n18955), .A(n18954), .B(n19270), .ZN(
        n18961) );
  XOR2_X1 U22149 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B(n18956), .Z(
        n19260) );
  MUX2_X1 U22150 ( .A(n18958), .B(n18957), .S(n19185), .Z(n18959) );
  XOR2_X1 U22151 ( .A(n18959), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n19272) );
  OAI22_X1 U22152 ( .A1(n19235), .A2(n19260), .B1(n19150), .B2(n19272), .ZN(
        n18960) );
  AOI211_X1 U22153 ( .C1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .C2(n18965), .A(
        n18961), .B(n18960), .ZN(n18962) );
  OAI21_X1 U22154 ( .B1(n19105), .B2(n19268), .A(n18962), .ZN(P3_U2805) );
  AOI221_X1 U22155 ( .B1(n18967), .B2(n18966), .C1(n18965), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n18964), .ZN(n18977) );
  OR2_X1 U22156 ( .A1(n18968), .A2(n19235), .ZN(n18971) );
  NAND2_X1 U22157 ( .A1(n19145), .A2(n18969), .ZN(n18970) );
  AND2_X1 U22158 ( .A1(n18971), .A2(n18970), .ZN(n18987) );
  OAI22_X1 U22159 ( .A1(n18987), .A2(n22186), .B1(n18972), .B2(n19150), .ZN(
        n18973) );
  AOI21_X1 U22160 ( .B1(n18975), .B2(n18974), .A(n18973), .ZN(n18976) );
  OAI211_X1 U22161 ( .C1(n19118), .C2(n11809), .A(n18977), .B(n18976), .ZN(
        P3_U2806) );
  INV_X1 U22162 ( .A(n19020), .ZN(n18992) );
  AOI21_X1 U22163 ( .B1(n19045), .B2(n18978), .A(n18990), .ZN(n18979) );
  AOI211_X1 U22164 ( .C1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n19185), .A(
        n18992), .B(n18979), .ZN(n18980) );
  XNOR2_X1 U22165 ( .A(n18980), .B(n18988), .ZN(n19275) );
  NOR2_X1 U22166 ( .A1(n14191), .A2(n20113), .ZN(n19274) );
  AOI21_X1 U22167 ( .B1(n18981), .B2(n19921), .A(
        P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n18982) );
  OAI22_X1 U22168 ( .A1(n19248), .A2(n18984), .B1(n18983), .B2(n18982), .ZN(
        n18985) );
  AOI211_X1 U22169 ( .C1(n19275), .C2(n19172), .A(n19274), .B(n18985), .ZN(
        n18986) );
  OAI221_X1 U22170 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n18989), 
        .C1(n18988), .C2(n18987), .A(n18986), .ZN(P3_U2807) );
  AOI21_X1 U22171 ( .B1(n19064), .B2(n19283), .A(n18990), .ZN(n18991) );
  NOR2_X1 U22172 ( .A1(n18992), .A2(n18991), .ZN(n18993) );
  XNOR2_X1 U22173 ( .A(n18993), .B(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n19292) );
  NOR2_X1 U22174 ( .A1(n19287), .A2(n19079), .ZN(n19002) );
  NOR2_X1 U22175 ( .A1(n19366), .A2(n19105), .ZN(n19092) );
  AOI21_X1 U22176 ( .B1(n10167), .B2(n19279), .A(n19092), .ZN(n19078) );
  OAI21_X1 U22177 ( .B1(n19283), .B2(n19019), .A(n19078), .ZN(n19012) );
  OAI21_X1 U22178 ( .B1(n18994), .B2(n19068), .A(n19207), .ZN(n18995) );
  AOI21_X1 U22179 ( .B1(n19067), .B2(n9888), .A(n18995), .ZN(n19015) );
  OAI21_X1 U22180 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n18996), .A(
        n19015), .ZN(n19006) );
  AOI22_X1 U22181 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n19006), .B1(
        n19128), .B2(n18997), .ZN(n19000) );
  NOR2_X1 U22182 ( .A1(n19026), .A2(n9888), .ZN(n19008) );
  OAI211_X1 U22183 ( .C1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A(n19008), .B(n18998), .ZN(n18999) );
  OAI211_X1 U22184 ( .C1(n20110), .C2(n14191), .A(n19000), .B(n18999), .ZN(
        n19001) );
  AOI221_X1 U22185 ( .B1(n19002), .B2(n19288), .C1(n19012), .C2(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n19001), .ZN(n19003) );
  OAI21_X1 U22186 ( .B1(n19150), .B2(n19292), .A(n19003), .ZN(P3_U2808) );
  NAND2_X1 U22187 ( .A1(n19297), .A2(n19286), .ZN(n19301) );
  NAND2_X1 U22188 ( .A1(n19331), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n19295) );
  OAI22_X1 U22189 ( .A1(n14191), .A2(n20108), .B1(n19118), .B2(n11806), .ZN(
        n19005) );
  AOI221_X1 U22190 ( .B1(n19008), .B2(n19007), .C1(n19006), .C2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(n19005), .ZN(n19014) );
  INV_X1 U22191 ( .A(n19045), .ZN(n19031) );
  NAND4_X1 U22192 ( .A1(n19064), .A2(n19331), .A3(n19063), .A4(
        P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n19032) );
  INV_X1 U22193 ( .A(n19032), .ZN(n19009) );
  AOI22_X1 U22194 ( .A1(n19031), .A2(n19010), .B1(n19297), .B2(n19009), .ZN(
        n19011) );
  XNOR2_X1 U22195 ( .A(n19011), .B(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n19294) );
  AOI22_X1 U22196 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n19012), .B1(
        n19172), .B2(n19294), .ZN(n19013) );
  OAI211_X1 U22197 ( .C1(n19301), .C2(n19037), .A(n19014), .B(n19013), .ZN(
        P3_U2809) );
  NAND2_X1 U22198 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n22088), .ZN(
        n19313) );
  AOI221_X1 U22199 ( .B1(n9789), .B2(n19016), .C1(n19882), .C2(n19016), .A(
        n19015), .ZN(n19017) );
  NOR2_X1 U22200 ( .A1(n14191), .A2(n20107), .ZN(n19309) );
  AOI211_X1 U22201 ( .C1(n19018), .C2(n19215), .A(n19017), .B(n19309), .ZN(
        n19024) );
  NOR2_X1 U22202 ( .A1(n19319), .A2(n19295), .ZN(n19303) );
  OAI21_X1 U22203 ( .B1(n19019), .B2(n19303), .A(n19078), .ZN(n19034) );
  OAI21_X1 U22204 ( .B1(n19043), .B2(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n19020), .ZN(n19021) );
  AOI21_X1 U22205 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n19032), .A(
        n19021), .ZN(n19022) );
  XNOR2_X1 U22206 ( .A(n19022), .B(n22088), .ZN(n19310) );
  AOI22_X1 U22207 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n19034), .B1(
        n19172), .B2(n19310), .ZN(n19023) );
  OAI211_X1 U22208 ( .C1(n19037), .C2(n19313), .A(n19024), .B(n19023), .ZN(
        P3_U2810) );
  AOI21_X1 U22209 ( .B1(n19067), .B2(n11801), .A(n19231), .ZN(n19055) );
  OAI21_X1 U22210 ( .B1(n19025), .B2(n19068), .A(n19055), .ZN(n19040) );
  NOR2_X1 U22211 ( .A1(n19026), .A2(n11801), .ZN(n19042) );
  OAI211_X1 U22212 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n19042), .B(n19027), .ZN(n19028) );
  NAND2_X1 U22213 ( .A1(n19508), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n19316) );
  OAI211_X1 U22214 ( .C1(n19118), .C2(n19029), .A(n19028), .B(n19316), .ZN(
        n19030) );
  AOI21_X1 U22215 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n19040), .A(
        n19030), .ZN(n19036) );
  NAND2_X1 U22216 ( .A1(n19031), .A2(n19043), .ZN(n19048) );
  NAND2_X1 U22217 ( .A1(n19048), .A2(n19032), .ZN(n19033) );
  XNOR2_X1 U22218 ( .A(n19033), .B(n19319), .ZN(n19315) );
  AOI22_X1 U22219 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n19034), .B1(
        n19172), .B2(n19315), .ZN(n19035) );
  OAI211_X1 U22220 ( .C1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n19037), .A(
        n19036), .B(n19035), .ZN(P3_U2811) );
  NAND2_X1 U22221 ( .A1(n19331), .A2(n17266), .ZN(n19338) );
  OAI22_X1 U22222 ( .A1(n14191), .A2(n20104), .B1(n19118), .B2(n19038), .ZN(
        n19039) );
  AOI221_X1 U22223 ( .B1(n19042), .B2(n19041), .C1(n19040), .C2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n19039), .ZN(n19051) );
  OAI21_X1 U22224 ( .B1(n19331), .B2(n19079), .A(n19078), .ZN(n19059) );
  NAND2_X1 U22225 ( .A1(n19063), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n19047) );
  INV_X1 U22226 ( .A(n19043), .ZN(n19044) );
  NAND2_X1 U22227 ( .A1(n19044), .A2(n19047), .ZN(n19046) );
  MUX2_X1 U22228 ( .A(n19047), .B(n19046), .S(n19045), .Z(n19049) );
  NAND2_X1 U22229 ( .A1(n19049), .A2(n19048), .ZN(n19334) );
  AOI22_X1 U22230 ( .A1(n19059), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .B1(
        n19172), .B2(n19334), .ZN(n19050) );
  OAI211_X1 U22231 ( .C1(n19079), .C2(n19338), .A(n19051), .B(n19050), .ZN(
        P3_U2812) );
  INV_X1 U22232 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n19339) );
  NAND2_X1 U22233 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n19339), .ZN(
        n19347) );
  XNOR2_X1 U22234 ( .A(n19052), .B(n19339), .ZN(n19343) );
  INV_X1 U22235 ( .A(n19343), .ZN(n19058) );
  NOR2_X1 U22236 ( .A1(n14191), .A2(n20102), .ZN(n19341) );
  AOI21_X1 U22237 ( .B1(n19053), .B2(n19921), .A(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n19056) );
  OAI22_X1 U22238 ( .A1(n19056), .A2(n19055), .B1(n19248), .B2(n19054), .ZN(
        n19057) );
  AOI211_X1 U22239 ( .C1(n19172), .C2(n19058), .A(n19341), .B(n19057), .ZN(
        n19061) );
  NAND2_X1 U22240 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n19059), .ZN(
        n19060) );
  OAI211_X1 U22241 ( .C1(n19347), .C2(n19079), .A(n19061), .B(n19060), .ZN(
        P3_U2813) );
  INV_X1 U22242 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n19360) );
  NAND2_X1 U22243 ( .A1(n10281), .A2(n19063), .ZN(n19164) );
  OAI22_X1 U22244 ( .A1(n19064), .A2(n19063), .B1(n19164), .B2(n19062), .ZN(
        n19065) );
  XOR2_X1 U22245 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B(n19065), .Z(
        n19357) );
  AOI21_X1 U22246 ( .B1(n19067), .B2(n19066), .A(n19231), .ZN(n19110) );
  OAI21_X1 U22247 ( .B1(n19069), .B2(n19068), .A(n19110), .ZN(n19083) );
  AOI22_X1 U22248 ( .A1(n19508), .A2(P3_REIP_REG_16__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n19083), .ZN(n19074) );
  NAND2_X1 U22249 ( .A1(n9890), .A2(n19070), .ZN(n19131) );
  NOR2_X1 U22250 ( .A1(n19071), .A2(n19131), .ZN(n19085) );
  OAI211_X1 U22251 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n19085), .B(n19072), .ZN(n19073) );
  OAI211_X1 U22252 ( .C1(n19118), .C2(n19075), .A(n19074), .B(n19073), .ZN(
        n19076) );
  AOI21_X1 U22253 ( .B1(n19172), .B2(n19357), .A(n19076), .ZN(n19077) );
  OAI221_X1 U22254 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n19079), 
        .C1(n19360), .C2(n19078), .A(n19077), .ZN(P3_U2814) );
  NAND2_X1 U22255 ( .A1(n19379), .A2(n19080), .ZN(n19396) );
  NOR3_X1 U22256 ( .A1(n10460), .A2(n19101), .A3(n19396), .ZN(n19100) );
  NOR2_X1 U22257 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n19100), .ZN(
        n19372) );
  NAND2_X1 U22258 ( .A1(n10167), .A2(n19279), .ZN(n19095) );
  NAND2_X1 U22259 ( .A1(n19508), .A2(P3_REIP_REG_15__SCAN_IN), .ZN(n19375) );
  OAI21_X1 U22260 ( .B1(n19118), .B2(n19081), .A(n19375), .ZN(n19082) );
  AOI221_X1 U22261 ( .B1(n19085), .B2(n19084), .C1(n19083), .C2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(n19082), .ZN(n19094) );
  NOR2_X1 U22262 ( .A1(n19101), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n19090) );
  INV_X1 U22263 ( .A(n19102), .ZN(n19088) );
  INV_X1 U22264 ( .A(n19423), .ZN(n19402) );
  NOR4_X1 U22265 ( .A1(n19086), .A2(n10460), .A3(n19402), .A4(n19101), .ZN(
        n19087) );
  NOR2_X1 U22266 ( .A1(n19088), .A2(n19087), .ZN(n19089) );
  AOI211_X1 U22267 ( .C1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n19185), .A(
        n19090), .B(n19089), .ZN(n19091) );
  XOR2_X1 U22268 ( .A(n19091), .B(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .Z(
        n19373) );
  NAND2_X1 U22269 ( .A1(n19104), .A2(n19377), .ZN(n19367) );
  AOI22_X1 U22270 ( .A1(n19172), .A2(n19373), .B1(n19092), .B2(n19367), .ZN(
        n19093) );
  OAI211_X1 U22271 ( .C1(n19372), .C2(n19095), .A(n19094), .B(n19093), .ZN(
        P3_U2815) );
  NOR2_X1 U22272 ( .A1(n19096), .A2(n19882), .ZN(n19169) );
  INV_X1 U22273 ( .A(n19169), .ZN(n19151) );
  NOR2_X1 U22274 ( .A1(n19097), .A2(n19151), .ZN(n19142) );
  AOI21_X1 U22275 ( .B1(n19098), .B2(n19142), .A(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n19109) );
  AOI22_X1 U22276 ( .A1(n19508), .A2(P3_REIP_REG_14__SCAN_IN), .B1(n19099), 
        .B2(n19215), .ZN(n19108) );
  AOI221_X1 U22277 ( .B1(n19415), .B2(n19101), .C1(n19362), .C2(n19101), .A(
        n19100), .ZN(n19387) );
  OAI22_X1 U22278 ( .A1(n19102), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B1(
        n19362), .B2(n19164), .ZN(n19103) );
  XNOR2_X1 U22279 ( .A(n19103), .B(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n19392) );
  NAND2_X1 U22280 ( .A1(n19418), .A2(n19379), .ZN(n19111) );
  INV_X1 U22281 ( .A(n19111), .ZN(n19393) );
  OAI221_X1 U22282 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .C1(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n19393), .A(n19104), .ZN(
        n19386) );
  OAI22_X1 U22283 ( .A1(n19392), .A2(n19150), .B1(n19105), .B2(n19386), .ZN(
        n19106) );
  AOI21_X1 U22284 ( .B1(n10167), .B2(n19387), .A(n19106), .ZN(n19107) );
  OAI211_X1 U22285 ( .C1(n19110), .C2(n19109), .A(n19108), .B(n19107), .ZN(
        P3_U2816) );
  AOI22_X1 U22286 ( .A1(n19145), .A2(n19111), .B1(n10167), .B2(n19396), .ZN(
        n19135) );
  AOI21_X1 U22287 ( .B1(n19113), .B2(n19112), .A(n19231), .ZN(n19114) );
  OAI21_X1 U22288 ( .B1(n9890), .B2(n19218), .A(n19114), .ZN(n19129) );
  NOR2_X1 U22289 ( .A1(n14191), .A2(n20095), .ZN(n19120) );
  OAI21_X1 U22290 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(n19115), .ZN(n19116) );
  OAI22_X1 U22291 ( .A1(n19118), .A2(n19117), .B1(n19131), .B2(n19116), .ZN(
        n19119) );
  AOI211_X1 U22292 ( .C1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n19129), .A(
        n19120), .B(n19119), .ZN(n19124) );
  OAI22_X1 U22293 ( .A1(n19125), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B1(
        n19164), .B2(n19122), .ZN(n19121) );
  XOR2_X1 U22294 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n19121), .Z(
        n19399) );
  NOR2_X1 U22295 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n19122), .ZN(
        n19398) );
  AOI22_X1 U22296 ( .A1(n19172), .A2(n19399), .B1(n19398), .B2(n19147), .ZN(
        n19123) );
  OAI211_X1 U22297 ( .C1(n19135), .C2(n10460), .A(n19124), .B(n19123), .ZN(
        P3_U2817) );
  INV_X1 U22298 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n22114) );
  OAI21_X1 U22299 ( .B1(n19402), .B2(n19164), .A(n19125), .ZN(n19126) );
  XOR2_X1 U22300 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B(n19126), .Z(
        n19407) );
  INV_X1 U22301 ( .A(n19147), .ZN(n19175) );
  NOR3_X1 U22302 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n19175), .A3(
        n19402), .ZN(n19133) );
  AOI22_X1 U22303 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n19129), .B1(
        n19128), .B2(n19127), .ZN(n19130) );
  NAND2_X1 U22304 ( .A1(n19508), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n19409) );
  OAI211_X1 U22305 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(n19131), .A(
        n19130), .B(n19409), .ZN(n19132) );
  AOI211_X1 U22306 ( .C1(n19172), .C2(n19407), .A(n19133), .B(n19132), .ZN(
        n19134) );
  OAI21_X1 U22307 ( .B1(n19135), .B2(n22114), .A(n19134), .ZN(P3_U2818) );
  INV_X1 U22308 ( .A(n19164), .ZN(n19137) );
  INV_X1 U22309 ( .A(n19146), .ZN(n19421) );
  AOI21_X1 U22310 ( .B1(n19137), .B2(n19421), .A(n19136), .ZN(n19139) );
  XNOR2_X1 U22311 ( .A(n19139), .B(n19138), .ZN(n19429) );
  AOI22_X1 U22312 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n19169), .B1(
        P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n19194), .ZN(n19141) );
  OAI22_X1 U22313 ( .A1(n19142), .A2(n19141), .B1(n19248), .B2(n19140), .ZN(
        n19143) );
  AOI21_X1 U22314 ( .B1(n19508), .B2(P3_REIP_REG_11__SCAN_IN), .A(n19143), 
        .ZN(n19149) );
  AOI22_X1 U22315 ( .A1(n19145), .A2(n19144), .B1(n10167), .B2(n19415), .ZN(
        n19174) );
  OAI21_X1 U22316 ( .B1(n19421), .B2(n19175), .A(n19174), .ZN(n19156) );
  NOR2_X1 U22317 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n19146), .ZN(
        n19411) );
  AOI22_X1 U22318 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n19156), .B1(
        n19411), .B2(n19147), .ZN(n19148) );
  OAI211_X1 U22319 ( .C1(n19429), .C2(n19150), .A(n19149), .B(n19148), .ZN(
        P3_U2819) );
  NOR2_X1 U22320 ( .A1(n19152), .A2(n19151), .ZN(n19160) );
  AOI21_X1 U22321 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n19194), .A(
        n19169), .ZN(n19159) );
  AOI22_X1 U22322 ( .A1(n19508), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n19153), 
        .B2(n19215), .ZN(n19158) );
  OAI21_X1 U22323 ( .B1(n19164), .B2(n10290), .A(n19162), .ZN(n19154) );
  XOR2_X1 U22324 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B(n19154), .Z(
        n19432) );
  OAI21_X1 U22325 ( .B1(n19175), .B2(n10290), .A(n10463), .ZN(n19155) );
  AOI22_X1 U22326 ( .A1(n19172), .A2(n19432), .B1(n19156), .B2(n19155), .ZN(
        n19157) );
  OAI211_X1 U22327 ( .C1(n19160), .C2(n19159), .A(n19158), .B(n19157), .ZN(
        P3_U2820) );
  NAND3_X1 U22328 ( .A1(n19164), .A2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(
        n19161), .ZN(n19163) );
  OAI211_X1 U22329 ( .C1(n19164), .C2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n19163), .B(n19162), .ZN(n19438) );
  NOR2_X1 U22330 ( .A1(n14191), .A2(n22085), .ZN(n19171) );
  NOR2_X1 U22331 ( .A1(n19165), .A2(n19179), .ZN(n19182) );
  AOI22_X1 U22332 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n19194), .B1(
        n19166), .B2(n19182), .ZN(n19168) );
  OAI22_X1 U22333 ( .A1(n19169), .A2(n19168), .B1(n19248), .B2(n19167), .ZN(
        n19170) );
  AOI211_X1 U22334 ( .C1(n19172), .C2(n19438), .A(n19171), .B(n19170), .ZN(
        n19173) );
  OAI221_X1 U22335 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n19175), .C1(
        n10290), .C2(n19174), .A(n19173), .ZN(P3_U2821) );
  OAI21_X1 U22336 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n19177), .A(
        n19176), .ZN(n19460) );
  NOR2_X1 U22337 ( .A1(n14191), .A2(n20086), .ZN(n19448) );
  OAI21_X1 U22338 ( .B1(n9894), .B2(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n19921), .ZN(n19181) );
  INV_X1 U22339 ( .A(n19178), .ZN(n19180) );
  OAI22_X1 U22340 ( .A1(n19182), .A2(n19181), .B1(n19180), .B2(n19179), .ZN(
        n19183) );
  AOI211_X1 U22341 ( .C1(n19184), .C2(n19215), .A(n19448), .B(n19183), .ZN(
        n19192) );
  NOR2_X1 U22342 ( .A1(n19450), .A2(n19185), .ZN(n19186) );
  NOR2_X1 U22343 ( .A1(n19187), .A2(n19186), .ZN(n19454) );
  MUX2_X1 U22344 ( .A(n19450), .B(n19454), .S(n19188), .Z(n19189) );
  NAND2_X1 U22345 ( .A1(n19190), .A2(n19189), .ZN(n19191) );
  OAI211_X1 U22346 ( .C1(n19235), .C2(n19460), .A(n19192), .B(n19191), .ZN(
        P3_U2822) );
  OR2_X1 U22347 ( .A1(n19193), .A2(n19882), .ZN(n19197) );
  NAND2_X1 U22348 ( .A1(n19194), .A2(n19197), .ZN(n19212) );
  XNOR2_X1 U22349 ( .A(n19196), .B(n19195), .ZN(n19474) );
  OAI22_X1 U22350 ( .A1(n19239), .A2(n19474), .B1(
        P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n19197), .ZN(n19202) );
  OAI21_X1 U22351 ( .B1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n19199), .A(
        n19198), .ZN(n19475) );
  OAI22_X1 U22352 ( .A1(n19248), .A2(n19200), .B1(n19235), .B2(n19475), .ZN(
        n19201) );
  AOI211_X1 U22353 ( .C1(n19508), .C2(P3_REIP_REG_6__SCAN_IN), .A(n19202), .B(
        n19201), .ZN(n19203) );
  OAI21_X1 U22354 ( .B1(n22084), .B2(n19212), .A(n19203), .ZN(P3_U2824) );
  OAI21_X1 U22355 ( .B1(n19206), .B2(n19205), .A(n19204), .ZN(n19484) );
  AOI21_X1 U22356 ( .B1(n19208), .B2(n19207), .A(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n19213) );
  XNOR2_X1 U22357 ( .A(n19209), .B(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n19210) );
  XNOR2_X1 U22358 ( .A(n19211), .B(n19210), .ZN(n19485) );
  OAI22_X1 U22359 ( .A1(n19213), .A2(n19212), .B1(n19239), .B2(n19485), .ZN(
        n19214) );
  AOI21_X1 U22360 ( .B1(n19216), .B2(n19215), .A(n19214), .ZN(n19217) );
  NAND2_X1 U22361 ( .A1(n19508), .A2(P3_REIP_REG_5__SCAN_IN), .ZN(n19480) );
  OAI211_X1 U22362 ( .C1(n19235), .C2(n19484), .A(n19217), .B(n19480), .ZN(
        P3_U2825) );
  NOR2_X1 U22363 ( .A1(n10078), .A2(n19218), .ZN(n19245) );
  NOR2_X1 U22364 ( .A1(n19231), .A2(n19245), .ZN(n19241) );
  OAI21_X1 U22365 ( .B1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n19220), .A(
        n19219), .ZN(n19500) );
  INV_X1 U22366 ( .A(n19221), .ZN(n19222) );
  OAI22_X1 U22367 ( .A1(n19235), .A2(n19500), .B1(n19882), .B2(n19222), .ZN(
        n19227) );
  XNOR2_X1 U22368 ( .A(n19224), .B(n19223), .ZN(n19494) );
  OAI22_X1 U22369 ( .A1(n19248), .A2(n19225), .B1(n19239), .B2(n19494), .ZN(
        n19226) );
  AOI211_X1 U22370 ( .C1(n19508), .C2(P3_REIP_REG_4__SCAN_IN), .A(n19227), .B(
        n19226), .ZN(n19228) );
  OAI21_X1 U22371 ( .B1(n19241), .B2(n22149), .A(n19228), .ZN(P3_U2826) );
  INV_X1 U22372 ( .A(n19229), .ZN(n19247) );
  NOR2_X1 U22373 ( .A1(n19231), .A2(n19230), .ZN(n19244) );
  OAI21_X1 U22374 ( .B1(n19234), .B2(n19233), .A(n19232), .ZN(n19503) );
  OAI22_X1 U22375 ( .A1(n19235), .A2(n19503), .B1(n14191), .B2(n20077), .ZN(
        n19243) );
  XNOR2_X1 U22376 ( .A(n19236), .B(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n19237) );
  XNOR2_X1 U22377 ( .A(n19238), .B(n19237), .ZN(n19504) );
  OAI22_X1 U22378 ( .A1(n19241), .A2(n19240), .B1(n19239), .B2(n19504), .ZN(
        n19242) );
  AOI211_X1 U22379 ( .C1(n19245), .C2(n19244), .A(n19243), .B(n19242), .ZN(
        n19246) );
  OAI21_X1 U22380 ( .B1(n19248), .B2(n19247), .A(n19246), .ZN(P3_U2827) );
  NOR2_X1 U22381 ( .A1(n19250), .A2(n19249), .ZN(n19254) );
  AOI21_X1 U22382 ( .B1(n19978), .B2(n17269), .A(n19251), .ZN(n19252) );
  INV_X1 U22383 ( .A(n19252), .ZN(n19253) );
  MUX2_X1 U22384 ( .A(n19254), .B(n19253), .S(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .Z(n19256) );
  AOI22_X1 U22385 ( .A1(n19457), .A2(n19256), .B1(n19455), .B2(n19255), .ZN(
        n19258) );
  OAI211_X1 U22386 ( .C1(n19512), .C2(n19259), .A(n19258), .B(n19257), .ZN(
        P3_U2835) );
  INV_X1 U22387 ( .A(n19260), .ZN(n19262) );
  AOI22_X1 U22388 ( .A1(n19416), .A2(n19262), .B1(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n19261), .ZN(n19267) );
  NAND3_X1 U22389 ( .A1(n19265), .A2(n19264), .A3(n19263), .ZN(n19266) );
  OAI211_X1 U22390 ( .C1(n19268), .C2(n19452), .A(n19267), .B(n19266), .ZN(
        n19269) );
  AOI22_X1 U22391 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n19473), .B1(
        n19457), .B2(n19269), .ZN(n19271) );
  OAI211_X1 U22392 ( .C1(n19272), .C2(n19428), .A(n19271), .B(n19270), .ZN(
        P3_U2837) );
  AOI21_X1 U22393 ( .B1(n19273), .B2(n19512), .A(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n19278) );
  AOI21_X1 U22394 ( .B1(n19275), .B2(n19455), .A(n19274), .ZN(n19276) );
  OAI21_X1 U22395 ( .B1(n19278), .B2(n19277), .A(n19276), .ZN(P3_U2839) );
  OAI221_X1 U22396 ( .B1(n19349), .B2(n19328), .C1(n19349), .C2(n19303), .A(
        n19281), .ZN(n19305) );
  NOR2_X1 U22397 ( .A1(n19416), .A2(n19282), .ZN(n19420) );
  OAI22_X1 U22398 ( .A1(n19349), .A2(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n19283), .B2(n19420), .ZN(n19284) );
  AOI22_X1 U22399 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n19473), .B1(
        n19457), .B2(n19289), .ZN(n19291) );
  NAND2_X1 U22400 ( .A1(n19508), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n19290) );
  OAI211_X1 U22401 ( .C1(n19292), .C2(n19428), .A(n19291), .B(n19290), .ZN(
        P3_U2840) );
  NOR3_X1 U22402 ( .A1(n19517), .A2(n19295), .A3(n19293), .ZN(n19314) );
  INV_X1 U22403 ( .A(n19314), .ZN(n19312) );
  AOI22_X1 U22404 ( .A1(n19508), .A2(P3_REIP_REG_21__SCAN_IN), .B1(n19455), 
        .B2(n19294), .ZN(n19300) );
  OAI21_X1 U22405 ( .B1(n19352), .B2(n19295), .A(n19986), .ZN(n19302) );
  OAI211_X1 U22406 ( .C1(n19297), .C2(n19381), .A(n19296), .B(n19302), .ZN(
        n19298) );
  OAI211_X1 U22407 ( .C1(n19517), .C2(n19298), .A(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n14191), .ZN(n19299) );
  OAI211_X1 U22408 ( .C1(n19312), .C2(n19301), .A(n19300), .B(n19299), .ZN(
        P3_U2841) );
  OAI211_X1 U22409 ( .C1(n19303), .C2(n19420), .A(n19512), .B(n19302), .ZN(
        n19304) );
  OAI21_X1 U22410 ( .B1(n19305), .B2(n19304), .A(n14191), .ZN(n19318) );
  NAND3_X1 U22411 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n19319), .A3(n19306), 
        .ZN(n19307) );
  AOI21_X1 U22412 ( .B1(n19318), .B2(n19307), .A(n22088), .ZN(n19308) );
  AOI211_X1 U22413 ( .C1(n19310), .C2(n19455), .A(n19309), .B(n19308), .ZN(
        n19311) );
  OAI21_X1 U22414 ( .B1(n19313), .B2(n19312), .A(n19311), .ZN(P3_U2842) );
  AOI22_X1 U22415 ( .A1(n19455), .A2(n19315), .B1(n19314), .B2(n19319), .ZN(
        n19317) );
  OAI211_X1 U22416 ( .C1(n19319), .C2(n19318), .A(n19317), .B(n19316), .ZN(
        P3_U2843) );
  INV_X1 U22417 ( .A(n19320), .ZN(n19321) );
  AOI22_X1 U22418 ( .A1(n19444), .A2(n19322), .B1(n19321), .B2(n19490), .ZN(
        n19502) );
  NOR2_X1 U22419 ( .A1(n19502), .A2(n19323), .ZN(n19461) );
  INV_X1 U22420 ( .A(n19461), .ZN(n19324) );
  NOR2_X1 U22421 ( .A1(n19325), .A2(n19324), .ZN(n19363) );
  NOR2_X1 U22422 ( .A1(n19326), .A2(n19363), .ZN(n19403) );
  NAND2_X1 U22423 ( .A1(n19327), .A2(n19437), .ZN(n19361) );
  NAND3_X1 U22424 ( .A1(n19328), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n19489), .ZN(n19333) );
  OR2_X1 U22425 ( .A1(n19517), .A2(n19329), .ZN(n19356) );
  OAI22_X1 U22426 ( .A1(n19331), .A2(n19420), .B1(n19330), .B2(n20019), .ZN(
        n19332) );
  AOI211_X1 U22427 ( .C1(n19442), .C2(n19333), .A(n19356), .B(n19332), .ZN(
        n19340) );
  AOI221_X1 U22428 ( .B1(n19488), .B2(n19340), .C1(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n19340), .A(n19508), .ZN(
        n19335) );
  AOI22_X1 U22429 ( .A1(n19335), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .B1(
        n19455), .B2(n19334), .ZN(n19337) );
  NAND2_X1 U22430 ( .A1(n19508), .A2(P3_REIP_REG_18__SCAN_IN), .ZN(n19336) );
  OAI211_X1 U22431 ( .C1(n19338), .C2(n19361), .A(n19337), .B(n19336), .ZN(
        P3_U2844) );
  NOR3_X1 U22432 ( .A1(n19508), .A2(n19340), .A3(n19339), .ZN(n19345) );
  INV_X1 U22433 ( .A(n19341), .ZN(n19342) );
  OAI21_X1 U22434 ( .B1(n19343), .B2(n19428), .A(n19342), .ZN(n19344) );
  NOR2_X1 U22435 ( .A1(n19345), .A2(n19344), .ZN(n19346) );
  OAI21_X1 U22436 ( .B1(n19361), .B2(n19347), .A(n19346), .ZN(P3_U2845) );
  OAI22_X1 U22437 ( .A1(n20019), .A2(n19350), .B1(n19349), .B2(n19348), .ZN(
        n19351) );
  INV_X1 U22438 ( .A(n19351), .ZN(n19412) );
  OAI21_X1 U22439 ( .B1(n19377), .B2(n19986), .A(n19352), .ZN(n19353) );
  OAI211_X1 U22440 ( .C1(n19354), .C2(n19422), .A(n19412), .B(n19353), .ZN(
        n19365) );
  OAI221_X1 U22441 ( .B1(n19356), .B2(n19355), .C1(n19356), .C2(n19365), .A(
        n14191), .ZN(n19359) );
  AOI22_X1 U22442 ( .A1(n19508), .A2(P3_REIP_REG_16__SCAN_IN), .B1(n19455), 
        .B2(n19357), .ZN(n19358) );
  OAI221_X1 U22443 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n19361), 
        .C1(n19360), .C2(n19359), .A(n19358), .ZN(P3_U2846) );
  INV_X1 U22444 ( .A(n19362), .ZN(n19380) );
  AND2_X1 U22445 ( .A1(n19380), .A2(n19363), .ZN(n19378) );
  OAI211_X1 U22446 ( .C1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n19378), .A(
        n19365), .B(n19364), .ZN(n19370) );
  NOR2_X1 U22447 ( .A1(n19366), .A2(n19452), .ZN(n19368) );
  NAND2_X1 U22448 ( .A1(n19368), .A2(n19367), .ZN(n19369) );
  OAI211_X1 U22449 ( .C1(n19372), .C2(n19371), .A(n19370), .B(n19369), .ZN(
        n19374) );
  AOI22_X1 U22450 ( .A1(n19457), .A2(n19374), .B1(n19455), .B2(n19373), .ZN(
        n19376) );
  OAI211_X1 U22451 ( .C1(n19512), .C2(n19377), .A(n19376), .B(n19375), .ZN(
        P3_U2847) );
  AOI22_X1 U22452 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n19473), .B1(
        n19508), .B2(P3_REIP_REG_14__SCAN_IN), .ZN(n19391) );
  INV_X1 U22453 ( .A(n19378), .ZN(n19384) );
  OAI221_X1 U22454 ( .B1(n19424), .B2(n19379), .C1(n19424), .C2(n19413), .A(
        n19412), .ZN(n19395) );
  OAI22_X1 U22455 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n19381), .B1(
        n19380), .B2(n19422), .ZN(n19382) );
  NOR2_X1 U22456 ( .A1(n19395), .A2(n19382), .ZN(n19383) );
  MUX2_X1 U22457 ( .A(n19384), .B(n19383), .S(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .Z(n19385) );
  OAI21_X1 U22458 ( .B1(n19452), .B2(n19386), .A(n19385), .ZN(n19389) );
  AOI22_X1 U22459 ( .A1(n19457), .A2(n19389), .B1(n19388), .B2(n19387), .ZN(
        n19390) );
  OAI211_X1 U22460 ( .C1(n19392), .C2(n19428), .A(n19391), .B(n19390), .ZN(
        P3_U2848) );
  OAI22_X1 U22461 ( .A1(n19423), .A2(n19422), .B1(n19393), .B2(n19452), .ZN(
        n19394) );
  AOI211_X1 U22462 ( .C1(n19416), .C2(n19396), .A(n19395), .B(n19394), .ZN(
        n19404) );
  OAI211_X1 U22463 ( .C1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n19422), .A(
        n19457), .B(n19404), .ZN(n19397) );
  NAND2_X1 U22464 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n19397), .ZN(
        n19401) );
  AOI22_X1 U22465 ( .A1(n19455), .A2(n19399), .B1(n19437), .B2(n19398), .ZN(
        n19400) );
  OAI221_X1 U22466 ( .B1(n19508), .B2(n19401), .C1(n14191), .C2(n20095), .A(
        n19400), .ZN(P3_U2849) );
  NOR2_X1 U22467 ( .A1(n19403), .A2(n19402), .ZN(n19406) );
  INV_X1 U22468 ( .A(n19404), .ZN(n19405) );
  MUX2_X1 U22469 ( .A(n19406), .B(n19405), .S(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .Z(n19408) );
  AOI22_X1 U22470 ( .A1(n19457), .A2(n19408), .B1(n19455), .B2(n19407), .ZN(
        n19410) );
  OAI211_X1 U22471 ( .C1(n19512), .C2(n22114), .A(n19410), .B(n19409), .ZN(
        P3_U2850) );
  AOI22_X1 U22472 ( .A1(n19508), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n19437), 
        .B2(n19411), .ZN(n19427) );
  OAI211_X1 U22473 ( .C1(n19424), .C2(n19413), .A(n19457), .B(n19412), .ZN(
        n19414) );
  AOI21_X1 U22474 ( .B1(n19416), .B2(n19415), .A(n19414), .ZN(n19417) );
  OAI21_X1 U22475 ( .B1(n19418), .B2(n19452), .A(n19417), .ZN(n19436) );
  AOI21_X1 U22476 ( .B1(n19986), .B2(n10290), .A(n19436), .ZN(n19419) );
  OAI21_X1 U22477 ( .B1(n19421), .B2(n19420), .A(n19419), .ZN(n19431) );
  OAI22_X1 U22478 ( .A1(n19424), .A2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B1(
        n19423), .B2(n19422), .ZN(n19425) );
  OAI211_X1 U22479 ( .C1(n19431), .C2(n19425), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n14191), .ZN(n19426) );
  OAI211_X1 U22480 ( .C1(n19429), .C2(n19428), .A(n19427), .B(n19426), .ZN(
        P3_U2851) );
  NAND2_X1 U22481 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n19437), .ZN(
        n19435) );
  OAI221_X1 U22482 ( .B1(n19431), .B2(n10290), .C1(n19431), .C2(n19430), .A(
        n14191), .ZN(n19434) );
  AOI22_X1 U22483 ( .A1(n19508), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n19455), 
        .B2(n19432), .ZN(n19433) );
  OAI221_X1 U22484 ( .B1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n19435), 
        .C1(n10463), .C2(n19434), .A(n19433), .ZN(P3_U2852) );
  NAND2_X1 U22485 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n19436), .ZN(
        n19440) );
  AOI22_X1 U22486 ( .A1(n19455), .A2(n19438), .B1(n19437), .B2(n10290), .ZN(
        n19439) );
  OAI221_X1 U22487 ( .B1(n19508), .B2(n19440), .C1(n14191), .C2(n22085), .A(
        n19439), .ZN(P3_U2853) );
  OAI21_X1 U22488 ( .B1(n19447), .B2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n19446) );
  AOI22_X1 U22489 ( .A1(n19444), .A2(n19443), .B1(n19442), .B2(n19441), .ZN(
        n19445) );
  AOI21_X1 U22490 ( .B1(n19445), .B2(n19489), .A(n19517), .ZN(n19472) );
  AOI21_X1 U22491 ( .B1(n19457), .B2(n19446), .A(n19472), .ZN(n19471) );
  OAI21_X1 U22492 ( .B1(n19447), .B2(n19471), .A(n19512), .ZN(n19449) );
  AOI21_X1 U22493 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n19449), .A(
        n19448), .ZN(n19459) );
  INV_X1 U22494 ( .A(n19450), .ZN(n19453) );
  NAND4_X1 U22495 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(n19461), .A4(n17256), .ZN(
        n19451) );
  OAI21_X1 U22496 ( .B1(n19453), .B2(n19452), .A(n19451), .ZN(n19456) );
  AOI22_X1 U22497 ( .A1(n19457), .A2(n19456), .B1(n19455), .B2(n19454), .ZN(
        n19458) );
  OAI211_X1 U22498 ( .C1(n10011), .C2(n19460), .A(n19459), .B(n19458), .ZN(
        P3_U2854) );
  NAND2_X1 U22499 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n19461), .ZN(
        n19469) );
  INV_X1 U22500 ( .A(n19462), .ZN(n19465) );
  INV_X1 U22501 ( .A(n19463), .ZN(n19464) );
  OAI22_X1 U22502 ( .A1(n10011), .A2(n19465), .B1(n19464), .B2(n19505), .ZN(
        n19466) );
  AOI211_X1 U22503 ( .C1(n19473), .C2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n19467), .B(n19466), .ZN(n19468) );
  OAI221_X1 U22504 ( .B1(n19471), .B2(n19470), .C1(n19471), .C2(n19469), .A(
        n19468), .ZN(P3_U2855) );
  NOR2_X1 U22505 ( .A1(n19473), .A2(n19472), .ZN(n19481) );
  NOR3_X1 U22506 ( .A1(n19502), .A2(n19517), .A3(n19511), .ZN(n19498) );
  NAND2_X1 U22507 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n19498), .ZN(
        n19483) );
  NOR2_X1 U22508 ( .A1(n19483), .A2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n19477) );
  OAI22_X1 U22509 ( .A1(n10011), .A2(n19475), .B1(n19505), .B2(n19474), .ZN(
        n19476) );
  AOI21_X1 U22510 ( .B1(n19477), .B2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n19476), .ZN(n19479) );
  NAND2_X1 U22511 ( .A1(n19508), .A2(P3_REIP_REG_6__SCAN_IN), .ZN(n19478) );
  OAI211_X1 U22512 ( .C1(n19481), .C2(n17248), .A(n19479), .B(n19478), .ZN(
        P3_U2856) );
  OAI221_X1 U22513 ( .B1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n19483), .C1(
        n19482), .C2(n19481), .A(n19480), .ZN(n19487) );
  OAI22_X1 U22514 ( .A1(n19505), .A2(n19485), .B1(n10011), .B2(n19484), .ZN(
        n19486) );
  OR2_X1 U22515 ( .A1(n19487), .A2(n19486), .ZN(P3_U2857) );
  INV_X1 U22516 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n19497) );
  AOI21_X1 U22517 ( .B1(n19490), .B2(n19489), .A(n19488), .ZN(n19491) );
  NOR3_X1 U22518 ( .A1(n19492), .A2(n19491), .A3(n19511), .ZN(n19501) );
  OAI21_X1 U22519 ( .B1(n19501), .B2(n19493), .A(n19512), .ZN(n19496) );
  OAI22_X1 U22520 ( .A1(n19505), .A2(n19494), .B1(n20079), .B2(n14191), .ZN(
        n19495) );
  AOI221_X1 U22521 ( .B1(n19498), .B2(n19497), .C1(n19496), .C2(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A(n19495), .ZN(n19499) );
  OAI21_X1 U22522 ( .B1(n10011), .B2(n19500), .A(n19499), .ZN(P3_U2858) );
  AOI211_X1 U22523 ( .C1(n19502), .C2(n19511), .A(n19501), .B(n19517), .ZN(
        n19507) );
  OAI22_X1 U22524 ( .A1(n19505), .A2(n19504), .B1(n10011), .B2(n19503), .ZN(
        n19506) );
  NOR2_X1 U22525 ( .A1(n19507), .A2(n19506), .ZN(n19510) );
  NAND2_X1 U22526 ( .A1(n19508), .A2(P3_REIP_REG_3__SCAN_IN), .ZN(n19509) );
  OAI211_X1 U22527 ( .C1(n19512), .C2(n19511), .A(n19510), .B(n19509), .ZN(
        P3_U2859) );
  NOR2_X1 U22528 ( .A1(n14191), .A2(n13930), .ZN(n19514) );
  NOR2_X1 U22529 ( .A1(n10011), .A2(n19516), .ZN(n19513) );
  AOI211_X1 U22530 ( .C1(n19516), .C2(n19515), .A(n19514), .B(n19513), .ZN(
        n19520) );
  OAI211_X1 U22531 ( .C1(n19978), .C2(n19517), .A(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B(n14191), .ZN(n19518) );
  NAND3_X1 U22532 ( .A1(n19520), .A2(n19519), .A3(n19518), .ZN(P3_U2862) );
  AOI21_X1 U22533 ( .B1(n19523), .B2(n19522), .A(n19521), .ZN(n20036) );
  OAI21_X1 U22534 ( .B1(n20036), .B2(n19566), .A(n19528), .ZN(n19524) );
  OAI221_X1 U22535 ( .B1(n11982), .B2(n20178), .C1(n11982), .C2(n19528), .A(
        n19524), .ZN(P3_U2863) );
  INV_X1 U22536 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20021) );
  NAND2_X1 U22537 ( .A1(n20011), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19778) );
  INV_X1 U22538 ( .A(n19778), .ZN(n19802) );
  INV_X1 U22539 ( .A(n19656), .ZN(n19706) );
  NOR2_X1 U22540 ( .A1(n19802), .A2(n19706), .ZN(n19526) );
  OAI22_X1 U22541 ( .A1(n19527), .A2(n20021), .B1(n19526), .B2(n19525), .ZN(
        P3_U2866) );
  NOR2_X1 U22542 ( .A1(n20022), .A2(n19528), .ZN(P3_U2867) );
  NAND2_X1 U22543 ( .A1(n19921), .A2(BUF2_REG_16__SCAN_IN), .ZN(n19888) );
  NAND2_X1 U22544 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19681), .ZN(
        n19914) );
  NOR2_X2 U22545 ( .A1(n19914), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19910) );
  NAND2_X1 U22546 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19856) );
  NOR2_X2 U22547 ( .A1(n19856), .A2(n19752), .ZN(n19958) );
  NAND2_X1 U22548 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n19921), .ZN(n19925) );
  INV_X1 U22549 ( .A(n19925), .ZN(n19881) );
  NOR2_X2 U22550 ( .A1(n19565), .A2(n22011), .ZN(n19916) );
  INV_X1 U22551 ( .A(n19914), .ZN(n19919) );
  NAND2_X1 U22552 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19919), .ZN(
        n19602) );
  NOR2_X1 U22553 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19611) );
  NOR2_X2 U22554 ( .A1(n20007), .A2(n19567), .ZN(n19618) );
  NAND2_X1 U22555 ( .A1(n19602), .A2(n19631), .ZN(n19529) );
  INV_X1 U22556 ( .A(n19529), .ZN(n19590) );
  NOR2_X1 U22557 ( .A1(n19915), .A2(n19590), .ZN(n19559) );
  AOI22_X1 U22558 ( .A1(n19958), .A2(n19881), .B1(n19916), .B2(n19559), .ZN(
        n19534) );
  INV_X1 U22559 ( .A(n19958), .ZN(n19974) );
  AOI21_X1 U22560 ( .B1(n19880), .B2(n19974), .A(n19565), .ZN(n19885) );
  AOI21_X1 U22561 ( .B1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        P3_STATE2_REG_3__SCAN_IN), .A(n19565), .ZN(n19682) );
  AOI22_X1 U22562 ( .A1(n19707), .A2(n19885), .B1(n19682), .B2(n19529), .ZN(
        n19562) );
  NAND2_X1 U22563 ( .A1(n19531), .A2(n19530), .ZN(n19560) );
  NOR2_X2 U22564 ( .A1(n19532), .A2(n19560), .ZN(n19922) );
  AOI22_X1 U22565 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19562), .B1(
        n19618), .B2(n19922), .ZN(n19533) );
  OAI211_X1 U22566 ( .C1(n19888), .C2(n19880), .A(n19534), .B(n19533), .ZN(
        P3_U2868) );
  NAND2_X1 U22567 ( .A1(n19921), .A2(BUF2_REG_17__SCAN_IN), .ZN(n19931) );
  NAND2_X1 U22568 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n19921), .ZN(n19892) );
  INV_X1 U22569 ( .A(n19892), .ZN(n19927) );
  AND2_X1 U22570 ( .A1(n19833), .A2(BUF2_REG_1__SCAN_IN), .ZN(n19926) );
  AOI22_X1 U22571 ( .A1(n19958), .A2(n19927), .B1(n19559), .B2(n19926), .ZN(
        n19537) );
  NOR2_X2 U22572 ( .A1(n19535), .A2(n19560), .ZN(n19928) );
  AOI22_X1 U22573 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19562), .B1(
        n19618), .B2(n19928), .ZN(n19536) );
  OAI211_X1 U22574 ( .C1(n19880), .C2(n19931), .A(n19537), .B(n19536), .ZN(
        P3_U2869) );
  NAND2_X1 U22575 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n19921), .ZN(n19811) );
  INV_X1 U22576 ( .A(n19811), .ZN(n19933) );
  NOR2_X2 U22577 ( .A1(n19565), .A2(n19538), .ZN(n19932) );
  AOI22_X1 U22578 ( .A1(n19958), .A2(n19933), .B1(n19559), .B2(n19932), .ZN(
        n19541) );
  NOR2_X2 U22579 ( .A1(n19539), .A2(n19560), .ZN(n19934) );
  AOI22_X1 U22580 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19562), .B1(
        n19618), .B2(n19934), .ZN(n19540) );
  OAI211_X1 U22581 ( .C1(n19880), .C2(n19937), .A(n19541), .B(n19540), .ZN(
        P3_U2870) );
  INV_X1 U22582 ( .A(n19895), .ZN(n19943) );
  INV_X1 U22583 ( .A(n19898), .ZN(n19939) );
  NOR2_X2 U22584 ( .A1(n19565), .A2(n19542), .ZN(n19938) );
  AOI22_X1 U22585 ( .A1(n19910), .A2(n19939), .B1(n19559), .B2(n19938), .ZN(
        n19545) );
  NOR2_X2 U22586 ( .A1(n19543), .A2(n19560), .ZN(n19940) );
  AOI22_X1 U22587 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19562), .B1(
        n19618), .B2(n19940), .ZN(n19544) );
  OAI211_X1 U22588 ( .C1(n19974), .C2(n19943), .A(n19545), .B(n19544), .ZN(
        P3_U2871) );
  NAND2_X1 U22589 ( .A1(n19921), .A2(BUF2_REG_20__SCAN_IN), .ZN(n19902) );
  INV_X1 U22590 ( .A(n19902), .ZN(n19945) );
  NOR2_X2 U22591 ( .A1(n19565), .A2(n19546), .ZN(n19944) );
  AOI22_X1 U22592 ( .A1(n19910), .A2(n19945), .B1(n19559), .B2(n19944), .ZN(
        n19549) );
  NOR2_X2 U22593 ( .A1(n19547), .A2(n19560), .ZN(n19946) );
  AOI22_X1 U22594 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19562), .B1(
        n19618), .B2(n19946), .ZN(n19548) );
  OAI211_X1 U22595 ( .C1(n19974), .C2(n19949), .A(n19549), .B(n19548), .ZN(
        P3_U2872) );
  NAND2_X1 U22596 ( .A1(n19921), .A2(BUF2_REG_21__SCAN_IN), .ZN(n19819) );
  NAND2_X1 U22597 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n19921), .ZN(n19955) );
  INV_X1 U22598 ( .A(n19955), .ZN(n19816) );
  NOR2_X2 U22599 ( .A1(n19565), .A2(n19550), .ZN(n19950) );
  AOI22_X1 U22600 ( .A1(n19958), .A2(n19816), .B1(n19559), .B2(n19950), .ZN(
        n19553) );
  NOR2_X2 U22601 ( .A1(n19551), .A2(n19560), .ZN(n19952) );
  AOI22_X1 U22602 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19562), .B1(
        n19618), .B2(n19952), .ZN(n19552) );
  OAI211_X1 U22603 ( .C1(n19880), .C2(n19819), .A(n19553), .B(n19552), .ZN(
        P3_U2873) );
  NAND2_X1 U22604 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n19921), .ZN(n19963) );
  NOR2_X2 U22605 ( .A1(n19565), .A2(n19554), .ZN(n19956) );
  AOI22_X1 U22606 ( .A1(n19958), .A2(n19872), .B1(n19559), .B2(n19956), .ZN(
        n19557) );
  NOR2_X2 U22607 ( .A1(n19555), .A2(n19560), .ZN(n19959) );
  AOI22_X1 U22608 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19562), .B1(
        n19618), .B2(n19959), .ZN(n19556) );
  OAI211_X1 U22609 ( .C1(n19880), .C2(n19875), .A(n19557), .B(n19556), .ZN(
        P3_U2874) );
  NAND2_X1 U22610 ( .A1(n19921), .A2(BUF2_REG_23__SCAN_IN), .ZN(n19973) );
  NAND2_X1 U22611 ( .A1(n19921), .A2(BUF2_REG_31__SCAN_IN), .ZN(n19829) );
  INV_X1 U22612 ( .A(n19829), .ZN(n19965) );
  NOR2_X2 U22613 ( .A1(n19565), .A2(n19558), .ZN(n19967) );
  AOI22_X1 U22614 ( .A1(n19958), .A2(n19965), .B1(n19559), .B2(n19967), .ZN(
        n19564) );
  NOR2_X2 U22615 ( .A1(n19561), .A2(n19560), .ZN(n19968) );
  AOI22_X1 U22616 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19562), .B1(
        n19618), .B2(n19968), .ZN(n19563) );
  OAI211_X1 U22617 ( .C1(n19880), .C2(n19973), .A(n19564), .B(n19563), .ZN(
        P3_U2875) );
  INV_X1 U22618 ( .A(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n19570) );
  NOR2_X1 U22619 ( .A1(n19566), .A2(n19565), .ZN(n19918) );
  NAND2_X1 U22620 ( .A1(n19918), .A2(n20002), .ZN(n19855) );
  OAI22_X1 U22621 ( .A1(n19882), .A2(n19914), .B1(n19567), .B2(n19855), .ZN(
        n19579) );
  NAND2_X1 U22622 ( .A1(n20002), .A2(n20046), .ZN(n19854) );
  NOR2_X1 U22623 ( .A1(n19567), .A2(n19854), .ZN(n19586) );
  AOI22_X1 U22624 ( .A1(n19910), .A2(n19881), .B1(n19916), .B2(n19586), .ZN(
        n19569) );
  INV_X1 U22625 ( .A(n19888), .ZN(n19917) );
  INV_X1 U22626 ( .A(n19602), .ZN(n19969) );
  NOR2_X2 U22627 ( .A1(n19567), .A2(n19752), .ZN(n19645) );
  AOI22_X1 U22628 ( .A1(n19917), .A2(n19969), .B1(n19922), .B2(n19645), .ZN(
        n19568) );
  OAI211_X1 U22629 ( .C1(n19570), .C2(n19579), .A(n19569), .B(n19568), .ZN(
        P3_U2876) );
  INV_X1 U22630 ( .A(n19931), .ZN(n19889) );
  AOI22_X1 U22631 ( .A1(n19969), .A2(n19889), .B1(n19926), .B2(n19586), .ZN(
        n19572) );
  AOI22_X1 U22632 ( .A1(n19910), .A2(n19927), .B1(n19928), .B2(n19645), .ZN(
        n19571) );
  OAI211_X1 U22633 ( .C1(n18473), .C2(n19579), .A(n19572), .B(n19571), .ZN(
        P3_U2877) );
  AOI22_X1 U22634 ( .A1(n19969), .A2(n19808), .B1(n19932), .B2(n19586), .ZN(
        n19574) );
  AOI22_X1 U22635 ( .A1(n19910), .A2(n19933), .B1(n19934), .B2(n19645), .ZN(
        n19573) );
  OAI211_X1 U22636 ( .C1(n19575), .C2(n19579), .A(n19574), .B(n19573), .ZN(
        P3_U2878) );
  INV_X1 U22637 ( .A(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n19578) );
  AOI22_X1 U22638 ( .A1(n19969), .A2(n19939), .B1(n19938), .B2(n19586), .ZN(
        n19577) );
  AOI22_X1 U22639 ( .A1(n19910), .A2(n19895), .B1(n19940), .B2(n19645), .ZN(
        n19576) );
  OAI211_X1 U22640 ( .C1(n19578), .C2(n19579), .A(n19577), .B(n19576), .ZN(
        P3_U2879) );
  AOI22_X1 U22641 ( .A1(n19969), .A2(n19945), .B1(n19944), .B2(n19586), .ZN(
        n19581) );
  INV_X1 U22642 ( .A(n19579), .ZN(n19587) );
  AOI22_X1 U22643 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19587), .B1(
        n19946), .B2(n19645), .ZN(n19580) );
  OAI211_X1 U22644 ( .C1(n19880), .C2(n19949), .A(n19581), .B(n19580), .ZN(
        P3_U2880) );
  INV_X1 U22645 ( .A(n19819), .ZN(n19951) );
  AOI22_X1 U22646 ( .A1(n19969), .A2(n19951), .B1(n19950), .B2(n19586), .ZN(
        n19583) );
  AOI22_X1 U22647 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19587), .B1(
        n19952), .B2(n19645), .ZN(n19582) );
  OAI211_X1 U22648 ( .C1(n19880), .C2(n19955), .A(n19583), .B(n19582), .ZN(
        P3_U2881) );
  AOI22_X1 U22649 ( .A1(n19910), .A2(n19872), .B1(n19956), .B2(n19586), .ZN(
        n19585) );
  AOI22_X1 U22650 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19587), .B1(
        n19959), .B2(n19645), .ZN(n19584) );
  OAI211_X1 U22651 ( .C1(n19602), .C2(n19875), .A(n19585), .B(n19584), .ZN(
        P3_U2882) );
  AOI22_X1 U22652 ( .A1(n19910), .A2(n19965), .B1(n19967), .B2(n19586), .ZN(
        n19589) );
  AOI22_X1 U22653 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19587), .B1(
        n19968), .B2(n19645), .ZN(n19588) );
  OAI211_X1 U22654 ( .C1(n19602), .C2(n19973), .A(n19589), .B(n19588), .ZN(
        P3_U2883) );
  NOR2_X2 U22655 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19655), .ZN(
        n19671) );
  NOR2_X1 U22656 ( .A1(n19645), .A2(n19671), .ZN(n19633) );
  NOR2_X1 U22657 ( .A1(n19915), .A2(n19633), .ZN(n19607) );
  AOI22_X1 U22658 ( .A1(n19969), .A2(n19881), .B1(n19916), .B2(n19607), .ZN(
        n19593) );
  OAI21_X1 U22659 ( .B1(n19590), .B2(n19830), .A(n19633), .ZN(n19591) );
  OAI211_X1 U22660 ( .C1(n19671), .C2(n20138), .A(n19833), .B(n19591), .ZN(
        n19608) );
  AOI22_X1 U22661 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19608), .B1(
        n19922), .B2(n19671), .ZN(n19592) );
  OAI211_X1 U22662 ( .C1(n19888), .C2(n19631), .A(n19593), .B(n19592), .ZN(
        P3_U2884) );
  AOI22_X1 U22663 ( .A1(n19969), .A2(n19927), .B1(n19926), .B2(n19607), .ZN(
        n19595) );
  AOI22_X1 U22664 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19608), .B1(
        n19928), .B2(n19671), .ZN(n19594) );
  OAI211_X1 U22665 ( .C1(n19631), .C2(n19931), .A(n19595), .B(n19594), .ZN(
        P3_U2885) );
  AOI22_X1 U22666 ( .A1(n19618), .A2(n19808), .B1(n19932), .B2(n19607), .ZN(
        n19597) );
  AOI22_X1 U22667 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19608), .B1(
        n19934), .B2(n19671), .ZN(n19596) );
  OAI211_X1 U22668 ( .C1(n19602), .C2(n19811), .A(n19597), .B(n19596), .ZN(
        P3_U2886) );
  AOI22_X1 U22669 ( .A1(n19969), .A2(n19895), .B1(n19938), .B2(n19607), .ZN(
        n19599) );
  AOI22_X1 U22670 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19608), .B1(
        n19940), .B2(n19671), .ZN(n19598) );
  OAI211_X1 U22671 ( .C1(n19631), .C2(n19898), .A(n19599), .B(n19598), .ZN(
        P3_U2887) );
  AOI22_X1 U22672 ( .A1(n19618), .A2(n19945), .B1(n19944), .B2(n19607), .ZN(
        n19601) );
  AOI22_X1 U22673 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19608), .B1(
        n19946), .B2(n19671), .ZN(n19600) );
  OAI211_X1 U22674 ( .C1(n19602), .C2(n19949), .A(n19601), .B(n19600), .ZN(
        P3_U2888) );
  AOI22_X1 U22675 ( .A1(n19969), .A2(n19816), .B1(n19950), .B2(n19607), .ZN(
        n19604) );
  AOI22_X1 U22676 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19608), .B1(
        n19952), .B2(n19671), .ZN(n19603) );
  OAI211_X1 U22677 ( .C1(n19631), .C2(n19819), .A(n19604), .B(n19603), .ZN(
        P3_U2889) );
  AOI22_X1 U22678 ( .A1(n19969), .A2(n19872), .B1(n19956), .B2(n19607), .ZN(
        n19606) );
  AOI22_X1 U22679 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19608), .B1(
        n19959), .B2(n19671), .ZN(n19605) );
  OAI211_X1 U22680 ( .C1(n19631), .C2(n19875), .A(n19606), .B(n19605), .ZN(
        P3_U2890) );
  AOI22_X1 U22681 ( .A1(n19969), .A2(n19965), .B1(n19967), .B2(n19607), .ZN(
        n19610) );
  AOI22_X1 U22682 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19608), .B1(
        n19968), .B2(n19671), .ZN(n19609) );
  OAI211_X1 U22683 ( .C1(n19631), .C2(n19973), .A(n19610), .B(n19609), .ZN(
        P3_U2891) );
  NOR2_X1 U22684 ( .A1(n19915), .A2(n19655), .ZN(n19627) );
  AOI22_X1 U22685 ( .A1(n19917), .A2(n19645), .B1(n19916), .B2(n19627), .ZN(
        n19613) );
  OAI211_X1 U22686 ( .C1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n19707), .A(
        n19611), .B(n19918), .ZN(n19628) );
  NOR2_X2 U22687 ( .A1(n11982), .A2(n19655), .ZN(n19692) );
  AOI22_X1 U22688 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19628), .B1(
        n19922), .B2(n19692), .ZN(n19612) );
  OAI211_X1 U22689 ( .C1(n19631), .C2(n19925), .A(n19613), .B(n19612), .ZN(
        P3_U2892) );
  AOI22_X1 U22690 ( .A1(n19618), .A2(n19927), .B1(n19926), .B2(n19627), .ZN(
        n19615) );
  AOI22_X1 U22691 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19628), .B1(
        n19928), .B2(n19692), .ZN(n19614) );
  OAI211_X1 U22692 ( .C1(n19931), .C2(n19654), .A(n19615), .B(n19614), .ZN(
        P3_U2893) );
  AOI22_X1 U22693 ( .A1(n19618), .A2(n19933), .B1(n19932), .B2(n19627), .ZN(
        n19617) );
  AOI22_X1 U22694 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19628), .B1(
        n19934), .B2(n19692), .ZN(n19616) );
  OAI211_X1 U22695 ( .C1(n19937), .C2(n19654), .A(n19617), .B(n19616), .ZN(
        P3_U2894) );
  AOI22_X1 U22696 ( .A1(n19618), .A2(n19895), .B1(n19938), .B2(n19627), .ZN(
        n19620) );
  AOI22_X1 U22697 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19628), .B1(
        n19940), .B2(n19692), .ZN(n19619) );
  OAI211_X1 U22698 ( .C1(n19898), .C2(n19654), .A(n19620), .B(n19619), .ZN(
        P3_U2895) );
  AOI22_X1 U22699 ( .A1(n19945), .A2(n19645), .B1(n19944), .B2(n19627), .ZN(
        n19622) );
  AOI22_X1 U22700 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19628), .B1(
        n19946), .B2(n19692), .ZN(n19621) );
  OAI211_X1 U22701 ( .C1(n19631), .C2(n19949), .A(n19622), .B(n19621), .ZN(
        P3_U2896) );
  AOI22_X1 U22702 ( .A1(n19951), .A2(n19645), .B1(n19950), .B2(n19627), .ZN(
        n19624) );
  AOI22_X1 U22703 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19628), .B1(
        n19952), .B2(n19692), .ZN(n19623) );
  OAI211_X1 U22704 ( .C1(n19631), .C2(n19955), .A(n19624), .B(n19623), .ZN(
        P3_U2897) );
  INV_X1 U22705 ( .A(n19875), .ZN(n19957) );
  AOI22_X1 U22706 ( .A1(n19957), .A2(n19645), .B1(n19956), .B2(n19627), .ZN(
        n19626) );
  AOI22_X1 U22707 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19628), .B1(
        n19959), .B2(n19692), .ZN(n19625) );
  OAI211_X1 U22708 ( .C1(n19631), .C2(n19963), .A(n19626), .B(n19625), .ZN(
        P3_U2898) );
  INV_X1 U22709 ( .A(n19973), .ZN(n19824) );
  AOI22_X1 U22710 ( .A1(n19824), .A2(n19645), .B1(n19967), .B2(n19627), .ZN(
        n19630) );
  AOI22_X1 U22711 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19628), .B1(
        n19968), .B2(n19692), .ZN(n19629) );
  OAI211_X1 U22712 ( .C1(n19631), .C2(n19829), .A(n19630), .B(n19629), .ZN(
        P3_U2899) );
  NOR2_X2 U22713 ( .A1(n20007), .A2(n19656), .ZN(n19720) );
  NAND2_X1 U22714 ( .A1(n19705), .A2(n19727), .ZN(n19683) );
  INV_X1 U22715 ( .A(n19683), .ZN(n19632) );
  NOR2_X1 U22716 ( .A1(n19915), .A2(n19632), .ZN(n19650) );
  AOI22_X1 U22717 ( .A1(n19917), .A2(n19671), .B1(n19916), .B2(n19650), .ZN(
        n19636) );
  OAI21_X1 U22718 ( .B1(n19633), .B2(n19830), .A(n19632), .ZN(n19634) );
  OAI211_X1 U22719 ( .C1(n19720), .C2(n20138), .A(n19833), .B(n19634), .ZN(
        n19651) );
  AOI22_X1 U22720 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19651), .B1(
        n19922), .B2(n19720), .ZN(n19635) );
  OAI211_X1 U22721 ( .C1(n19925), .C2(n19654), .A(n19636), .B(n19635), .ZN(
        P3_U2900) );
  AOI22_X1 U22722 ( .A1(n19889), .A2(n19671), .B1(n19926), .B2(n19650), .ZN(
        n19638) );
  AOI22_X1 U22723 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19651), .B1(
        n19928), .B2(n19720), .ZN(n19637) );
  OAI211_X1 U22724 ( .C1(n19892), .C2(n19654), .A(n19638), .B(n19637), .ZN(
        P3_U2901) );
  AOI22_X1 U22725 ( .A1(n19933), .A2(n19645), .B1(n19932), .B2(n19650), .ZN(
        n19640) );
  AOI22_X1 U22726 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19651), .B1(
        n19934), .B2(n19720), .ZN(n19639) );
  OAI211_X1 U22727 ( .C1(n19937), .C2(n19680), .A(n19640), .B(n19639), .ZN(
        P3_U2902) );
  AOI22_X1 U22728 ( .A1(n19895), .A2(n19645), .B1(n19938), .B2(n19650), .ZN(
        n19642) );
  AOI22_X1 U22729 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19651), .B1(
        n19940), .B2(n19720), .ZN(n19641) );
  OAI211_X1 U22730 ( .C1(n19898), .C2(n19680), .A(n19642), .B(n19641), .ZN(
        P3_U2903) );
  AOI22_X1 U22731 ( .A1(n19945), .A2(n19671), .B1(n19944), .B2(n19650), .ZN(
        n19644) );
  AOI22_X1 U22732 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19651), .B1(
        n19946), .B2(n19720), .ZN(n19643) );
  OAI211_X1 U22733 ( .C1(n19949), .C2(n19654), .A(n19644), .B(n19643), .ZN(
        P3_U2904) );
  AOI22_X1 U22734 ( .A1(n19816), .A2(n19645), .B1(n19950), .B2(n19650), .ZN(
        n19647) );
  AOI22_X1 U22735 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19651), .B1(
        n19952), .B2(n19720), .ZN(n19646) );
  OAI211_X1 U22736 ( .C1(n19819), .C2(n19680), .A(n19647), .B(n19646), .ZN(
        P3_U2905) );
  AOI22_X1 U22737 ( .A1(n19957), .A2(n19671), .B1(n19956), .B2(n19650), .ZN(
        n19649) );
  AOI22_X1 U22738 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19651), .B1(
        n19959), .B2(n19720), .ZN(n19648) );
  OAI211_X1 U22739 ( .C1(n19963), .C2(n19654), .A(n19649), .B(n19648), .ZN(
        P3_U2906) );
  AOI22_X1 U22740 ( .A1(n19824), .A2(n19671), .B1(n19967), .B2(n19650), .ZN(
        n19653) );
  AOI22_X1 U22741 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19651), .B1(
        n19968), .B2(n19720), .ZN(n19652) );
  OAI211_X1 U22742 ( .C1(n19829), .C2(n19654), .A(n19653), .B(n19652), .ZN(
        P3_U2907) );
  OAI22_X1 U22743 ( .A1(n19882), .A2(n19655), .B1(n19656), .B2(n19855), .ZN(
        n19674) );
  NOR2_X1 U22744 ( .A1(n19656), .A2(n19854), .ZN(n19676) );
  AOI22_X1 U22745 ( .A1(n19917), .A2(n19692), .B1(n19916), .B2(n19676), .ZN(
        n19658) );
  NOR2_X2 U22746 ( .A1(n19656), .A2(n19752), .ZN(n19740) );
  AOI22_X1 U22747 ( .A1(n19922), .A2(n19740), .B1(n19881), .B2(n19671), .ZN(
        n19657) );
  OAI211_X1 U22748 ( .C1(n22148), .C2(n19674), .A(n19658), .B(n19657), .ZN(
        P3_U2908) );
  AOI22_X1 U22749 ( .A1(n19889), .A2(n19692), .B1(n19926), .B2(n19676), .ZN(
        n19660) );
  INV_X1 U22750 ( .A(n19674), .ZN(n19677) );
  AOI22_X1 U22751 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19677), .B1(
        n19928), .B2(n19740), .ZN(n19659) );
  OAI211_X1 U22752 ( .C1(n19892), .C2(n19680), .A(n19660), .B(n19659), .ZN(
        P3_U2909) );
  AOI22_X1 U22753 ( .A1(n19808), .A2(n19692), .B1(n19932), .B2(n19676), .ZN(
        n19662) );
  AOI22_X1 U22754 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19677), .B1(
        n19934), .B2(n19740), .ZN(n19661) );
  OAI211_X1 U22755 ( .C1(n19811), .C2(n19680), .A(n19662), .B(n19661), .ZN(
        P3_U2910) );
  AOI22_X1 U22756 ( .A1(n19938), .A2(n19676), .B1(n19939), .B2(n19692), .ZN(
        n19664) );
  AOI22_X1 U22757 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19677), .B1(
        n19940), .B2(n19740), .ZN(n19663) );
  OAI211_X1 U22758 ( .C1(n19943), .C2(n19680), .A(n19664), .B(n19663), .ZN(
        P3_U2911) );
  INV_X1 U22759 ( .A(n19949), .ZN(n19899) );
  AOI22_X1 U22760 ( .A1(n19899), .A2(n19671), .B1(n19944), .B2(n19676), .ZN(
        n19666) );
  AOI22_X1 U22761 ( .A1(n19946), .A2(n19740), .B1(n19945), .B2(n19692), .ZN(
        n19665) );
  OAI211_X1 U22762 ( .C1(n19667), .C2(n19674), .A(n19666), .B(n19665), .ZN(
        P3_U2912) );
  AOI22_X1 U22763 ( .A1(n19816), .A2(n19671), .B1(n19950), .B2(n19676), .ZN(
        n19669) );
  AOI22_X1 U22764 ( .A1(n19951), .A2(n19692), .B1(n19952), .B2(n19740), .ZN(
        n19668) );
  OAI211_X1 U22765 ( .C1(n19670), .C2(n19674), .A(n19669), .B(n19668), .ZN(
        P3_U2913) );
  AOI22_X1 U22766 ( .A1(n19872), .A2(n19671), .B1(n19956), .B2(n19676), .ZN(
        n19673) );
  AOI22_X1 U22767 ( .A1(n19957), .A2(n19692), .B1(n19959), .B2(n19740), .ZN(
        n19672) );
  OAI211_X1 U22768 ( .C1(n19675), .C2(n19674), .A(n19673), .B(n19672), .ZN(
        P3_U2914) );
  AOI22_X1 U22769 ( .A1(n19824), .A2(n19692), .B1(n19967), .B2(n19676), .ZN(
        n19679) );
  AOI22_X1 U22770 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19677), .B1(
        n19968), .B2(n19740), .ZN(n19678) );
  OAI211_X1 U22771 ( .C1(n19829), .C2(n19680), .A(n19679), .B(n19678), .ZN(
        P3_U2915) );
  NAND2_X1 U22772 ( .A1(n19681), .A2(n20021), .ZN(n19751) );
  NOR2_X1 U22773 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19751), .ZN(
        n19685) );
  INV_X1 U22774 ( .A(n19685), .ZN(n19743) );
  NAND2_X1 U22775 ( .A1(n19750), .A2(n19743), .ZN(n19684) );
  INV_X1 U22776 ( .A(n19684), .ZN(n19728) );
  NOR2_X1 U22777 ( .A1(n19915), .A2(n19728), .ZN(n19701) );
  AOI22_X1 U22778 ( .A1(n19917), .A2(n19720), .B1(n19916), .B2(n19701), .ZN(
        n19687) );
  OAI221_X1 U22779 ( .B1(n19684), .B2(n19707), .C1(n19684), .C2(n19683), .A(
        n19682), .ZN(n19702) );
  CLKBUF_X1 U22780 ( .A(n19685), .Z(n19773) );
  AOI22_X1 U22781 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19702), .B1(
        n19922), .B2(n19773), .ZN(n19686) );
  OAI211_X1 U22782 ( .C1(n19925), .C2(n19705), .A(n19687), .B(n19686), .ZN(
        P3_U2916) );
  AOI22_X1 U22783 ( .A1(n19889), .A2(n19720), .B1(n19926), .B2(n19701), .ZN(
        n19689) );
  AOI22_X1 U22784 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19702), .B1(
        n19928), .B2(n19773), .ZN(n19688) );
  OAI211_X1 U22785 ( .C1(n19892), .C2(n19705), .A(n19689), .B(n19688), .ZN(
        P3_U2917) );
  AOI22_X1 U22786 ( .A1(n19808), .A2(n19720), .B1(n19932), .B2(n19701), .ZN(
        n19691) );
  AOI22_X1 U22787 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19702), .B1(
        n19934), .B2(n19773), .ZN(n19690) );
  OAI211_X1 U22788 ( .C1(n19811), .C2(n19705), .A(n19691), .B(n19690), .ZN(
        P3_U2918) );
  AOI22_X1 U22789 ( .A1(n19895), .A2(n19692), .B1(n19938), .B2(n19701), .ZN(
        n19694) );
  AOI22_X1 U22790 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19702), .B1(
        n19940), .B2(n19773), .ZN(n19693) );
  OAI211_X1 U22791 ( .C1(n19898), .C2(n19727), .A(n19694), .B(n19693), .ZN(
        P3_U2919) );
  AOI22_X1 U22792 ( .A1(n19945), .A2(n19720), .B1(n19944), .B2(n19701), .ZN(
        n19696) );
  AOI22_X1 U22793 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19702), .B1(
        n19946), .B2(n19773), .ZN(n19695) );
  OAI211_X1 U22794 ( .C1(n19949), .C2(n19705), .A(n19696), .B(n19695), .ZN(
        P3_U2920) );
  AOI22_X1 U22795 ( .A1(n19951), .A2(n19720), .B1(n19950), .B2(n19701), .ZN(
        n19698) );
  AOI22_X1 U22796 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19702), .B1(
        n19952), .B2(n19773), .ZN(n19697) );
  OAI211_X1 U22797 ( .C1(n19955), .C2(n19705), .A(n19698), .B(n19697), .ZN(
        P3_U2921) );
  AOI22_X1 U22798 ( .A1(n19957), .A2(n19720), .B1(n19956), .B2(n19701), .ZN(
        n19700) );
  AOI22_X1 U22799 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19702), .B1(
        n19959), .B2(n19773), .ZN(n19699) );
  OAI211_X1 U22800 ( .C1(n19963), .C2(n19705), .A(n19700), .B(n19699), .ZN(
        P3_U2922) );
  AOI22_X1 U22801 ( .A1(n19824), .A2(n19720), .B1(n19967), .B2(n19701), .ZN(
        n19704) );
  AOI22_X1 U22802 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19702), .B1(
        n19968), .B2(n19773), .ZN(n19703) );
  OAI211_X1 U22803 ( .C1(n19829), .C2(n19705), .A(n19704), .B(n19703), .ZN(
        P3_U2923) );
  NOR2_X1 U22804 ( .A1(n19915), .A2(n19751), .ZN(n19723) );
  AOI22_X1 U22805 ( .A1(n19917), .A2(n19740), .B1(n19916), .B2(n19723), .ZN(
        n19709) );
  OAI211_X1 U22806 ( .C1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n19707), .A(
        n19706), .B(n19918), .ZN(n19724) );
  NOR2_X1 U22807 ( .A1(n11982), .A2(n19751), .ZN(n19792) );
  AOI22_X1 U22808 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19724), .B1(
        n19922), .B2(n19792), .ZN(n19708) );
  OAI211_X1 U22809 ( .C1(n19925), .C2(n19727), .A(n19709), .B(n19708), .ZN(
        P3_U2924) );
  AOI22_X1 U22810 ( .A1(n19889), .A2(n19740), .B1(n19926), .B2(n19723), .ZN(
        n19711) );
  AOI22_X1 U22811 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19724), .B1(
        n19928), .B2(n19785), .ZN(n19710) );
  OAI211_X1 U22812 ( .C1(n19892), .C2(n19727), .A(n19711), .B(n19710), .ZN(
        P3_U2925) );
  AOI22_X1 U22813 ( .A1(n19933), .A2(n19720), .B1(n19932), .B2(n19723), .ZN(
        n19713) );
  AOI22_X1 U22814 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19724), .B1(
        n19934), .B2(n19785), .ZN(n19712) );
  OAI211_X1 U22815 ( .C1(n19937), .C2(n19750), .A(n19713), .B(n19712), .ZN(
        P3_U2926) );
  AOI22_X1 U22816 ( .A1(n19938), .A2(n19723), .B1(n19939), .B2(n19740), .ZN(
        n19715) );
  AOI22_X1 U22817 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19724), .B1(
        n19940), .B2(n19785), .ZN(n19714) );
  OAI211_X1 U22818 ( .C1(n19943), .C2(n19727), .A(n19715), .B(n19714), .ZN(
        P3_U2927) );
  AOI22_X1 U22819 ( .A1(n19899), .A2(n19720), .B1(n19944), .B2(n19723), .ZN(
        n19717) );
  AOI22_X1 U22820 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19724), .B1(
        n19946), .B2(n19792), .ZN(n19716) );
  OAI211_X1 U22821 ( .C1(n19902), .C2(n19750), .A(n19717), .B(n19716), .ZN(
        P3_U2928) );
  AOI22_X1 U22822 ( .A1(n19951), .A2(n19740), .B1(n19950), .B2(n19723), .ZN(
        n19719) );
  AOI22_X1 U22823 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19724), .B1(
        n19952), .B2(n19785), .ZN(n19718) );
  OAI211_X1 U22824 ( .C1(n19955), .C2(n19727), .A(n19719), .B(n19718), .ZN(
        P3_U2929) );
  AOI22_X1 U22825 ( .A1(n19872), .A2(n19720), .B1(n19956), .B2(n19723), .ZN(
        n19722) );
  AOI22_X1 U22826 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19724), .B1(
        n19959), .B2(n19785), .ZN(n19721) );
  OAI211_X1 U22827 ( .C1(n19875), .C2(n19750), .A(n19722), .B(n19721), .ZN(
        P3_U2930) );
  AOI22_X1 U22828 ( .A1(n19824), .A2(n19740), .B1(n19967), .B2(n19723), .ZN(
        n19726) );
  AOI22_X1 U22829 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19724), .B1(
        n19968), .B2(n19785), .ZN(n19725) );
  OAI211_X1 U22830 ( .C1(n19829), .C2(n19727), .A(n19726), .B(n19725), .ZN(
        P3_U2931) );
  NOR2_X2 U22831 ( .A1(n20007), .A2(n19778), .ZN(n19820) );
  NOR2_X1 U22832 ( .A1(n19785), .A2(n19820), .ZN(n19779) );
  NOR2_X1 U22833 ( .A1(n19915), .A2(n19779), .ZN(n19746) );
  AOI22_X1 U22834 ( .A1(n19917), .A2(n19773), .B1(n19916), .B2(n19746), .ZN(
        n19731) );
  OAI21_X1 U22835 ( .B1(n19728), .B2(n19830), .A(n19779), .ZN(n19729) );
  OAI211_X1 U22836 ( .C1(n19820), .C2(n20138), .A(n19833), .B(n19729), .ZN(
        n19747) );
  AOI22_X1 U22837 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19747), .B1(
        n19922), .B2(n19820), .ZN(n19730) );
  OAI211_X1 U22838 ( .C1(n19925), .C2(n19750), .A(n19731), .B(n19730), .ZN(
        P3_U2932) );
  AOI22_X1 U22839 ( .A1(n19889), .A2(n19773), .B1(n19926), .B2(n19746), .ZN(
        n19733) );
  AOI22_X1 U22840 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19747), .B1(
        n19928), .B2(n19820), .ZN(n19732) );
  OAI211_X1 U22841 ( .C1(n19892), .C2(n19750), .A(n19733), .B(n19732), .ZN(
        P3_U2933) );
  AOI22_X1 U22842 ( .A1(n19933), .A2(n19740), .B1(n19932), .B2(n19746), .ZN(
        n19735) );
  AOI22_X1 U22843 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19747), .B1(
        n19934), .B2(n19820), .ZN(n19734) );
  OAI211_X1 U22844 ( .C1(n19937), .C2(n19743), .A(n19735), .B(n19734), .ZN(
        P3_U2934) );
  AOI22_X1 U22845 ( .A1(n19895), .A2(n19740), .B1(n19938), .B2(n19746), .ZN(
        n19737) );
  AOI22_X1 U22846 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19747), .B1(
        n19940), .B2(n19820), .ZN(n19736) );
  OAI211_X1 U22847 ( .C1(n19898), .C2(n19743), .A(n19737), .B(n19736), .ZN(
        P3_U2935) );
  AOI22_X1 U22848 ( .A1(n19899), .A2(n19740), .B1(n19944), .B2(n19746), .ZN(
        n19739) );
  AOI22_X1 U22849 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19747), .B1(
        n19946), .B2(n19820), .ZN(n19738) );
  OAI211_X1 U22850 ( .C1(n19902), .C2(n19743), .A(n19739), .B(n19738), .ZN(
        P3_U2936) );
  AOI22_X1 U22851 ( .A1(n19816), .A2(n19740), .B1(n19950), .B2(n19746), .ZN(
        n19742) );
  AOI22_X1 U22852 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19747), .B1(
        n19952), .B2(n19820), .ZN(n19741) );
  OAI211_X1 U22853 ( .C1(n19819), .C2(n19743), .A(n19742), .B(n19741), .ZN(
        P3_U2937) );
  AOI22_X1 U22854 ( .A1(n19957), .A2(n19773), .B1(n19956), .B2(n19746), .ZN(
        n19745) );
  AOI22_X1 U22855 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19747), .B1(
        n19959), .B2(n19820), .ZN(n19744) );
  OAI211_X1 U22856 ( .C1(n19963), .C2(n19750), .A(n19745), .B(n19744), .ZN(
        P3_U2938) );
  AOI22_X1 U22857 ( .A1(n19824), .A2(n19773), .B1(n19967), .B2(n19746), .ZN(
        n19749) );
  AOI22_X1 U22858 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19747), .B1(
        n19968), .B2(n19820), .ZN(n19748) );
  OAI211_X1 U22859 ( .C1(n19829), .C2(n19750), .A(n19749), .B(n19748), .ZN(
        P3_U2939) );
  OAI22_X1 U22860 ( .A1(n19882), .A2(n19751), .B1(n19778), .B2(n19855), .ZN(
        n19776) );
  NOR2_X1 U22861 ( .A1(n19778), .A2(n19854), .ZN(n19772) );
  AOI22_X1 U22862 ( .A1(n19917), .A2(n19792), .B1(n19916), .B2(n19772), .ZN(
        n19754) );
  NOR2_X2 U22863 ( .A1(n19778), .A2(n19752), .ZN(n19849) );
  AOI22_X1 U22864 ( .A1(n19922), .A2(n19849), .B1(n19881), .B2(n19773), .ZN(
        n19753) );
  OAI211_X1 U22865 ( .C1(n19755), .C2(n19776), .A(n19754), .B(n19753), .ZN(
        P3_U2940) );
  AOI22_X1 U22866 ( .A1(n19927), .A2(n19773), .B1(n19926), .B2(n19772), .ZN(
        n19757) );
  AOI22_X1 U22867 ( .A1(n19889), .A2(n19792), .B1(n19928), .B2(n19849), .ZN(
        n19756) );
  OAI211_X1 U22868 ( .C1(n19758), .C2(n19776), .A(n19757), .B(n19756), .ZN(
        P3_U2941) );
  INV_X1 U22869 ( .A(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n22139) );
  AOI22_X1 U22870 ( .A1(n19808), .A2(n19785), .B1(n19932), .B2(n19772), .ZN(
        n19760) );
  AOI22_X1 U22871 ( .A1(n19934), .A2(n19849), .B1(n19933), .B2(n19773), .ZN(
        n19759) );
  OAI211_X1 U22872 ( .C1(n22139), .C2(n19776), .A(n19760), .B(n19759), .ZN(
        P3_U2942) );
  INV_X1 U22873 ( .A(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n19763) );
  AOI22_X1 U22874 ( .A1(n19895), .A2(n19773), .B1(n19938), .B2(n19772), .ZN(
        n19762) );
  AOI22_X1 U22875 ( .A1(n19940), .A2(n19849), .B1(n19939), .B2(n19792), .ZN(
        n19761) );
  OAI211_X1 U22876 ( .C1(n19763), .C2(n19776), .A(n19762), .B(n19761), .ZN(
        P3_U2943) );
  AOI22_X1 U22877 ( .A1(n19945), .A2(n19785), .B1(n19944), .B2(n19772), .ZN(
        n19765) );
  AOI22_X1 U22878 ( .A1(n19899), .A2(n19773), .B1(n19946), .B2(n19849), .ZN(
        n19764) );
  OAI211_X1 U22879 ( .C1(n18419), .C2(n19776), .A(n19765), .B(n19764), .ZN(
        P3_U2944) );
  INV_X1 U22880 ( .A(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n19768) );
  AOI22_X1 U22881 ( .A1(n19951), .A2(n19792), .B1(n19950), .B2(n19772), .ZN(
        n19767) );
  AOI22_X1 U22882 ( .A1(n19952), .A2(n19849), .B1(n19816), .B2(n19773), .ZN(
        n19766) );
  OAI211_X1 U22883 ( .C1(n19768), .C2(n19776), .A(n19767), .B(n19766), .ZN(
        P3_U2945) );
  INV_X1 U22884 ( .A(n19792), .ZN(n19801) );
  AOI22_X1 U22885 ( .A1(n19872), .A2(n19773), .B1(n19956), .B2(n19772), .ZN(
        n19771) );
  INV_X1 U22886 ( .A(n19776), .ZN(n19769) );
  AOI22_X1 U22887 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19769), .B1(
        n19959), .B2(n19849), .ZN(n19770) );
  OAI211_X1 U22888 ( .C1(n19875), .C2(n19801), .A(n19771), .B(n19770), .ZN(
        P3_U2946) );
  AOI22_X1 U22889 ( .A1(n19824), .A2(n19792), .B1(n19967), .B2(n19772), .ZN(
        n19775) );
  AOI22_X1 U22890 ( .A1(n19968), .A2(n19849), .B1(n19965), .B2(n19773), .ZN(
        n19774) );
  OAI211_X1 U22891 ( .C1(n19777), .C2(n19776), .A(n19775), .B(n19774), .ZN(
        P3_U2947) );
  NAND2_X1 U22892 ( .A1(n11982), .A2(n19803), .ZN(n19871) );
  INV_X1 U22893 ( .A(n19871), .ZN(n19876) );
  NOR2_X1 U22894 ( .A1(n19849), .A2(n19876), .ZN(n19831) );
  NOR2_X1 U22895 ( .A1(n19915), .A2(n19831), .ZN(n19797) );
  AOI22_X1 U22896 ( .A1(n19916), .A2(n19797), .B1(n19881), .B2(n19785), .ZN(
        n19782) );
  OAI21_X1 U22897 ( .B1(n19779), .B2(n19830), .A(n19831), .ZN(n19780) );
  OAI211_X1 U22898 ( .C1(n19876), .C2(n20138), .A(n19833), .B(n19780), .ZN(
        n19798) );
  AOI22_X1 U22899 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19798), .B1(
        n19922), .B2(n19876), .ZN(n19781) );
  OAI211_X1 U22900 ( .C1(n19888), .C2(n19828), .A(n19782), .B(n19781), .ZN(
        P3_U2948) );
  AOI22_X1 U22901 ( .A1(n19927), .A2(n19785), .B1(n19926), .B2(n19797), .ZN(
        n19784) );
  AOI22_X1 U22902 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19798), .B1(
        n19928), .B2(n19876), .ZN(n19783) );
  OAI211_X1 U22903 ( .C1(n19931), .C2(n19828), .A(n19784), .B(n19783), .ZN(
        P3_U2949) );
  AOI22_X1 U22904 ( .A1(n19933), .A2(n19785), .B1(n19932), .B2(n19797), .ZN(
        n19787) );
  AOI22_X1 U22905 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19798), .B1(
        n19934), .B2(n19876), .ZN(n19786) );
  OAI211_X1 U22906 ( .C1(n19937), .C2(n19828), .A(n19787), .B(n19786), .ZN(
        P3_U2950) );
  AOI22_X1 U22907 ( .A1(n19895), .A2(n19792), .B1(n19938), .B2(n19797), .ZN(
        n19789) );
  AOI22_X1 U22908 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19798), .B1(
        n19940), .B2(n19876), .ZN(n19788) );
  OAI211_X1 U22909 ( .C1(n19898), .C2(n19828), .A(n19789), .B(n19788), .ZN(
        P3_U2951) );
  AOI22_X1 U22910 ( .A1(n19945), .A2(n19820), .B1(n19944), .B2(n19797), .ZN(
        n19791) );
  AOI22_X1 U22911 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19798), .B1(
        n19946), .B2(n19876), .ZN(n19790) );
  OAI211_X1 U22912 ( .C1(n19949), .C2(n19801), .A(n19791), .B(n19790), .ZN(
        P3_U2952) );
  AOI22_X1 U22913 ( .A1(n19816), .A2(n19792), .B1(n19950), .B2(n19797), .ZN(
        n19794) );
  AOI22_X1 U22914 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19798), .B1(
        n19952), .B2(n19876), .ZN(n19793) );
  OAI211_X1 U22915 ( .C1(n19819), .C2(n19828), .A(n19794), .B(n19793), .ZN(
        P3_U2953) );
  AOI22_X1 U22916 ( .A1(n19957), .A2(n19820), .B1(n19956), .B2(n19797), .ZN(
        n19796) );
  AOI22_X1 U22917 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19798), .B1(
        n19959), .B2(n19876), .ZN(n19795) );
  OAI211_X1 U22918 ( .C1(n19963), .C2(n19801), .A(n19796), .B(n19795), .ZN(
        P3_U2954) );
  AOI22_X1 U22919 ( .A1(n19824), .A2(n19820), .B1(n19967), .B2(n19797), .ZN(
        n19800) );
  AOI22_X1 U22920 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19798), .B1(
        n19968), .B2(n19876), .ZN(n19799) );
  OAI211_X1 U22921 ( .C1(n19829), .C2(n19801), .A(n19800), .B(n19799), .ZN(
        P3_U2955) );
  INV_X1 U22922 ( .A(n19803), .ZN(n19857) );
  NOR2_X1 U22923 ( .A1(n19915), .A2(n19857), .ZN(n19823) );
  AOI22_X1 U22924 ( .A1(n19917), .A2(n19849), .B1(n19916), .B2(n19823), .ZN(
        n19805) );
  AOI22_X1 U22925 ( .A1(n19921), .A2(n19802), .B1(n19918), .B2(n19803), .ZN(
        n19825) );
  NAND2_X1 U22926 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19803), .ZN(
        n19907) );
  INV_X1 U22927 ( .A(n19907), .ZN(n19908) );
  AOI22_X1 U22928 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19825), .B1(
        n19922), .B2(n19908), .ZN(n19804) );
  OAI211_X1 U22929 ( .C1(n19925), .C2(n19828), .A(n19805), .B(n19804), .ZN(
        P3_U2956) );
  INV_X1 U22930 ( .A(n19849), .ZN(n19846) );
  AOI22_X1 U22931 ( .A1(n19927), .A2(n19820), .B1(n19926), .B2(n19823), .ZN(
        n19807) );
  AOI22_X1 U22932 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19825), .B1(
        n19928), .B2(n19908), .ZN(n19806) );
  OAI211_X1 U22933 ( .C1(n19931), .C2(n19846), .A(n19807), .B(n19806), .ZN(
        P3_U2957) );
  AOI22_X1 U22934 ( .A1(n19808), .A2(n19849), .B1(n19932), .B2(n19823), .ZN(
        n19810) );
  AOI22_X1 U22935 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19825), .B1(
        n19934), .B2(n19908), .ZN(n19809) );
  OAI211_X1 U22936 ( .C1(n19811), .C2(n19828), .A(n19810), .B(n19809), .ZN(
        P3_U2958) );
  AOI22_X1 U22937 ( .A1(n19938), .A2(n19823), .B1(n19939), .B2(n19849), .ZN(
        n19813) );
  AOI22_X1 U22938 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19825), .B1(
        n19940), .B2(n19908), .ZN(n19812) );
  OAI211_X1 U22939 ( .C1(n19943), .C2(n19828), .A(n19813), .B(n19812), .ZN(
        P3_U2959) );
  AOI22_X1 U22940 ( .A1(n19945), .A2(n19849), .B1(n19944), .B2(n19823), .ZN(
        n19815) );
  AOI22_X1 U22941 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19825), .B1(
        n19946), .B2(n19908), .ZN(n19814) );
  OAI211_X1 U22942 ( .C1(n19949), .C2(n19828), .A(n19815), .B(n19814), .ZN(
        P3_U2960) );
  AOI22_X1 U22943 ( .A1(n19816), .A2(n19820), .B1(n19950), .B2(n19823), .ZN(
        n19818) );
  AOI22_X1 U22944 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19825), .B1(
        n19952), .B2(n19908), .ZN(n19817) );
  OAI211_X1 U22945 ( .C1(n19819), .C2(n19846), .A(n19818), .B(n19817), .ZN(
        P3_U2961) );
  AOI22_X1 U22946 ( .A1(n19872), .A2(n19820), .B1(n19956), .B2(n19823), .ZN(
        n19822) );
  AOI22_X1 U22947 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19825), .B1(
        n19959), .B2(n19908), .ZN(n19821) );
  OAI211_X1 U22948 ( .C1(n19875), .C2(n19846), .A(n19822), .B(n19821), .ZN(
        P3_U2962) );
  AOI22_X1 U22949 ( .A1(n19824), .A2(n19849), .B1(n19967), .B2(n19823), .ZN(
        n19827) );
  AOI22_X1 U22950 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19825), .B1(
        n19968), .B2(n19908), .ZN(n19826) );
  OAI211_X1 U22951 ( .C1(n19829), .C2(n19828), .A(n19827), .B(n19826), .ZN(
        P3_U2963) );
  NOR2_X2 U22952 ( .A1(n20007), .A2(n19856), .ZN(n19964) );
  NOR2_X1 U22953 ( .A1(n19908), .A2(n19964), .ZN(n19883) );
  NOR2_X1 U22954 ( .A1(n19915), .A2(n19883), .ZN(n19850) );
  AOI22_X1 U22955 ( .A1(n19916), .A2(n19850), .B1(n19881), .B2(n19849), .ZN(
        n19835) );
  OAI21_X1 U22956 ( .B1(n19831), .B2(n19830), .A(n19883), .ZN(n19832) );
  OAI211_X1 U22957 ( .C1(n19964), .C2(n20138), .A(n19833), .B(n19832), .ZN(
        n19851) );
  AOI22_X1 U22958 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19851), .B1(
        n19922), .B2(n19964), .ZN(n19834) );
  OAI211_X1 U22959 ( .C1(n19888), .C2(n19871), .A(n19835), .B(n19834), .ZN(
        P3_U2964) );
  AOI22_X1 U22960 ( .A1(n19889), .A2(n19876), .B1(n19926), .B2(n19850), .ZN(
        n19837) );
  AOI22_X1 U22961 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19851), .B1(
        n19928), .B2(n19964), .ZN(n19836) );
  OAI211_X1 U22962 ( .C1(n19892), .C2(n19846), .A(n19837), .B(n19836), .ZN(
        P3_U2965) );
  AOI22_X1 U22963 ( .A1(n19933), .A2(n19849), .B1(n19932), .B2(n19850), .ZN(
        n19839) );
  AOI22_X1 U22964 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19851), .B1(
        n19934), .B2(n19964), .ZN(n19838) );
  OAI211_X1 U22965 ( .C1(n19937), .C2(n19871), .A(n19839), .B(n19838), .ZN(
        P3_U2966) );
  AOI22_X1 U22966 ( .A1(n19895), .A2(n19849), .B1(n19938), .B2(n19850), .ZN(
        n19841) );
  AOI22_X1 U22967 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19851), .B1(
        n19940), .B2(n19964), .ZN(n19840) );
  OAI211_X1 U22968 ( .C1(n19898), .C2(n19871), .A(n19841), .B(n19840), .ZN(
        P3_U2967) );
  AOI22_X1 U22969 ( .A1(n19945), .A2(n19876), .B1(n19944), .B2(n19850), .ZN(
        n19843) );
  AOI22_X1 U22970 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19851), .B1(
        n19946), .B2(n19964), .ZN(n19842) );
  OAI211_X1 U22971 ( .C1(n19949), .C2(n19846), .A(n19843), .B(n19842), .ZN(
        P3_U2968) );
  AOI22_X1 U22972 ( .A1(n19951), .A2(n19876), .B1(n19950), .B2(n19850), .ZN(
        n19845) );
  AOI22_X1 U22973 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19851), .B1(
        n19952), .B2(n19964), .ZN(n19844) );
  OAI211_X1 U22974 ( .C1(n19955), .C2(n19846), .A(n19845), .B(n19844), .ZN(
        P3_U2969) );
  AOI22_X1 U22975 ( .A1(n19872), .A2(n19849), .B1(n19956), .B2(n19850), .ZN(
        n19848) );
  AOI22_X1 U22976 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19851), .B1(
        n19959), .B2(n19964), .ZN(n19847) );
  OAI211_X1 U22977 ( .C1(n19875), .C2(n19871), .A(n19848), .B(n19847), .ZN(
        P3_U2970) );
  AOI22_X1 U22978 ( .A1(n19967), .A2(n19850), .B1(n19965), .B2(n19849), .ZN(
        n19853) );
  AOI22_X1 U22979 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19851), .B1(
        n19968), .B2(n19964), .ZN(n19852) );
  OAI211_X1 U22980 ( .C1(n19973), .C2(n19871), .A(n19853), .B(n19852), .ZN(
        P3_U2971) );
  NOR2_X1 U22981 ( .A1(n19856), .A2(n19854), .ZN(n19920) );
  AOI22_X1 U22982 ( .A1(n19916), .A2(n19920), .B1(n19881), .B2(n19876), .ZN(
        n19860) );
  OAI22_X1 U22983 ( .A1(n19882), .A2(n19857), .B1(n19856), .B2(n19855), .ZN(
        n19858) );
  INV_X1 U22984 ( .A(n19858), .ZN(n19877) );
  AOI22_X1 U22985 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19877), .B1(
        n19958), .B2(n19922), .ZN(n19859) );
  OAI211_X1 U22986 ( .C1(n19888), .C2(n19907), .A(n19860), .B(n19859), .ZN(
        P3_U2972) );
  AOI22_X1 U22987 ( .A1(n19889), .A2(n19908), .B1(n19926), .B2(n19920), .ZN(
        n19862) );
  AOI22_X1 U22988 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19877), .B1(
        n19958), .B2(n19928), .ZN(n19861) );
  OAI211_X1 U22989 ( .C1(n19892), .C2(n19871), .A(n19862), .B(n19861), .ZN(
        P3_U2973) );
  AOI22_X1 U22990 ( .A1(n19933), .A2(n19876), .B1(n19932), .B2(n19920), .ZN(
        n19864) );
  AOI22_X1 U22991 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19877), .B1(
        n19958), .B2(n19934), .ZN(n19863) );
  OAI211_X1 U22992 ( .C1(n19937), .C2(n19907), .A(n19864), .B(n19863), .ZN(
        P3_U2974) );
  AOI22_X1 U22993 ( .A1(n19895), .A2(n19876), .B1(n19938), .B2(n19920), .ZN(
        n19866) );
  AOI22_X1 U22994 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19877), .B1(
        n19958), .B2(n19940), .ZN(n19865) );
  OAI211_X1 U22995 ( .C1(n19898), .C2(n19907), .A(n19866), .B(n19865), .ZN(
        P3_U2975) );
  AOI22_X1 U22996 ( .A1(n19899), .A2(n19876), .B1(n19944), .B2(n19920), .ZN(
        n19868) );
  AOI22_X1 U22997 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19877), .B1(
        n19958), .B2(n19946), .ZN(n19867) );
  OAI211_X1 U22998 ( .C1(n19902), .C2(n19907), .A(n19868), .B(n19867), .ZN(
        P3_U2976) );
  AOI22_X1 U22999 ( .A1(n19951), .A2(n19908), .B1(n19950), .B2(n19920), .ZN(
        n19870) );
  AOI22_X1 U23000 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19877), .B1(
        n19958), .B2(n19952), .ZN(n19869) );
  OAI211_X1 U23001 ( .C1(n19955), .C2(n19871), .A(n19870), .B(n19869), .ZN(
        P3_U2977) );
  AOI22_X1 U23002 ( .A1(n19872), .A2(n19876), .B1(n19956), .B2(n19920), .ZN(
        n19874) );
  AOI22_X1 U23003 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19877), .B1(
        n19958), .B2(n19959), .ZN(n19873) );
  OAI211_X1 U23004 ( .C1(n19875), .C2(n19907), .A(n19874), .B(n19873), .ZN(
        P3_U2978) );
  AOI22_X1 U23005 ( .A1(n19967), .A2(n19920), .B1(n19965), .B2(n19876), .ZN(
        n19879) );
  AOI22_X1 U23006 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19877), .B1(
        n19958), .B2(n19968), .ZN(n19878) );
  OAI211_X1 U23007 ( .C1(n19973), .C2(n19907), .A(n19879), .B(n19878), .ZN(
        P3_U2979) );
  INV_X1 U23008 ( .A(n19964), .ZN(n19962) );
  AOI21_X1 U23009 ( .B1(n19880), .B2(n19974), .A(n19915), .ZN(n19909) );
  AOI22_X1 U23010 ( .A1(n19916), .A2(n19909), .B1(n19881), .B2(n19908), .ZN(
        n19887) );
  NOR2_X1 U23011 ( .A1(n19883), .A2(n19882), .ZN(n19884) );
  OAI22_X1 U23012 ( .A1(n19910), .A2(n20138), .B1(n19885), .B2(n19884), .ZN(
        n19911) );
  AOI22_X1 U23013 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19911), .B1(
        n19910), .B2(n19922), .ZN(n19886) );
  OAI211_X1 U23014 ( .C1(n19888), .C2(n19962), .A(n19887), .B(n19886), .ZN(
        P3_U2980) );
  AOI22_X1 U23015 ( .A1(n19889), .A2(n19964), .B1(n19926), .B2(n19909), .ZN(
        n19891) );
  AOI22_X1 U23016 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19911), .B1(
        n19910), .B2(n19928), .ZN(n19890) );
  OAI211_X1 U23017 ( .C1(n19892), .C2(n19907), .A(n19891), .B(n19890), .ZN(
        P3_U2981) );
  AOI22_X1 U23018 ( .A1(n19933), .A2(n19908), .B1(n19932), .B2(n19909), .ZN(
        n19894) );
  AOI22_X1 U23019 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19911), .B1(
        n19910), .B2(n19934), .ZN(n19893) );
  OAI211_X1 U23020 ( .C1(n19937), .C2(n19962), .A(n19894), .B(n19893), .ZN(
        P3_U2982) );
  AOI22_X1 U23021 ( .A1(n19895), .A2(n19908), .B1(n19938), .B2(n19909), .ZN(
        n19897) );
  AOI22_X1 U23022 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19911), .B1(
        n19910), .B2(n19940), .ZN(n19896) );
  OAI211_X1 U23023 ( .C1(n19898), .C2(n19962), .A(n19897), .B(n19896), .ZN(
        P3_U2983) );
  AOI22_X1 U23024 ( .A1(n19899), .A2(n19908), .B1(n19944), .B2(n19909), .ZN(
        n19901) );
  AOI22_X1 U23025 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19911), .B1(
        n19910), .B2(n19946), .ZN(n19900) );
  OAI211_X1 U23026 ( .C1(n19902), .C2(n19962), .A(n19901), .B(n19900), .ZN(
        P3_U2984) );
  AOI22_X1 U23027 ( .A1(n19951), .A2(n19964), .B1(n19950), .B2(n19909), .ZN(
        n19904) );
  AOI22_X1 U23028 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19911), .B1(
        n19910), .B2(n19952), .ZN(n19903) );
  OAI211_X1 U23029 ( .C1(n19955), .C2(n19907), .A(n19904), .B(n19903), .ZN(
        P3_U2985) );
  AOI22_X1 U23030 ( .A1(n19957), .A2(n19964), .B1(n19956), .B2(n19909), .ZN(
        n19906) );
  AOI22_X1 U23031 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19911), .B1(
        n19910), .B2(n19959), .ZN(n19905) );
  OAI211_X1 U23032 ( .C1(n19963), .C2(n19907), .A(n19906), .B(n19905), .ZN(
        P3_U2986) );
  AOI22_X1 U23033 ( .A1(n19967), .A2(n19909), .B1(n19965), .B2(n19908), .ZN(
        n19913) );
  AOI22_X1 U23034 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19911), .B1(
        n19910), .B2(n19968), .ZN(n19912) );
  OAI211_X1 U23035 ( .C1(n19973), .C2(n19962), .A(n19913), .B(n19912), .ZN(
        P3_U2987) );
  NOR2_X1 U23036 ( .A1(n19915), .A2(n19914), .ZN(n19966) );
  AOI22_X1 U23037 ( .A1(n19917), .A2(n19958), .B1(n19916), .B2(n19966), .ZN(
        n19924) );
  AOI22_X1 U23038 ( .A1(n19921), .A2(n19920), .B1(n19919), .B2(n19918), .ZN(
        n19970) );
  AOI22_X1 U23039 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19970), .B1(
        n19969), .B2(n19922), .ZN(n19923) );
  OAI211_X1 U23040 ( .C1(n19925), .C2(n19962), .A(n19924), .B(n19923), .ZN(
        P3_U2988) );
  AOI22_X1 U23041 ( .A1(n19927), .A2(n19964), .B1(n19926), .B2(n19966), .ZN(
        n19930) );
  AOI22_X1 U23042 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19970), .B1(
        n19969), .B2(n19928), .ZN(n19929) );
  OAI211_X1 U23043 ( .C1(n19974), .C2(n19931), .A(n19930), .B(n19929), .ZN(
        P3_U2989) );
  AOI22_X1 U23044 ( .A1(n19933), .A2(n19964), .B1(n19932), .B2(n19966), .ZN(
        n19936) );
  AOI22_X1 U23045 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19970), .B1(
        n19969), .B2(n19934), .ZN(n19935) );
  OAI211_X1 U23046 ( .C1(n19974), .C2(n19937), .A(n19936), .B(n19935), .ZN(
        P3_U2990) );
  AOI22_X1 U23047 ( .A1(n19958), .A2(n19939), .B1(n19938), .B2(n19966), .ZN(
        n19942) );
  AOI22_X1 U23048 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19970), .B1(
        n19969), .B2(n19940), .ZN(n19941) );
  OAI211_X1 U23049 ( .C1(n19943), .C2(n19962), .A(n19942), .B(n19941), .ZN(
        P3_U2991) );
  AOI22_X1 U23050 ( .A1(n19958), .A2(n19945), .B1(n19944), .B2(n19966), .ZN(
        n19948) );
  AOI22_X1 U23051 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19970), .B1(
        n19969), .B2(n19946), .ZN(n19947) );
  OAI211_X1 U23052 ( .C1(n19949), .C2(n19962), .A(n19948), .B(n19947), .ZN(
        P3_U2992) );
  AOI22_X1 U23053 ( .A1(n19958), .A2(n19951), .B1(n19950), .B2(n19966), .ZN(
        n19954) );
  AOI22_X1 U23054 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19970), .B1(
        n19969), .B2(n19952), .ZN(n19953) );
  OAI211_X1 U23055 ( .C1(n19955), .C2(n19962), .A(n19954), .B(n19953), .ZN(
        P3_U2993) );
  AOI22_X1 U23056 ( .A1(n19958), .A2(n19957), .B1(n19956), .B2(n19966), .ZN(
        n19961) );
  AOI22_X1 U23057 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19970), .B1(
        n19969), .B2(n19959), .ZN(n19960) );
  OAI211_X1 U23058 ( .C1(n19963), .C2(n19962), .A(n19961), .B(n19960), .ZN(
        P3_U2994) );
  AOI22_X1 U23059 ( .A1(n19967), .A2(n19966), .B1(n19965), .B2(n19964), .ZN(
        n19972) );
  AOI22_X1 U23060 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19970), .B1(
        n19969), .B2(n19968), .ZN(n19971) );
  OAI211_X1 U23061 ( .C1(n19974), .C2(n19973), .A(n19972), .B(n19971), .ZN(
        P3_U2995) );
  AOI21_X1 U23062 ( .B1(n19977), .B2(n19976), .A(n19975), .ZN(n19989) );
  NAND2_X1 U23063 ( .A1(n19978), .A2(n19997), .ZN(n19980) );
  INV_X1 U23064 ( .A(n19982), .ZN(n19979) );
  OAI211_X1 U23065 ( .C1(n19981), .C2(n19989), .A(n19980), .B(n19979), .ZN(
        n20145) );
  NOR2_X1 U23066 ( .A1(n20025), .A2(n20145), .ZN(n19985) );
  OAI22_X1 U23067 ( .A1(n19983), .A2(n19997), .B1(n20019), .B2(n19982), .ZN(
        n20144) );
  NAND2_X1 U23068 ( .A1(n20146), .A2(n20144), .ZN(n19984) );
  OAI22_X1 U23069 ( .A1(n19985), .A2(n20146), .B1(n20025), .B2(n19984), .ZN(
        n20033) );
  INV_X1 U23070 ( .A(n20025), .ZN(n20001) );
  NAND2_X1 U23071 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n19986), .ZN(
        n19987) );
  NAND2_X1 U23072 ( .A1(n19987), .A2(n19990), .ZN(n19988) );
  NAND2_X1 U23073 ( .A1(n19988), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n19994) );
  OAI21_X1 U23074 ( .B1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n19990), .A(
        n19989), .ZN(n19991) );
  NAND2_X1 U23075 ( .A1(n19992), .A2(n19991), .ZN(n19993) );
  MUX2_X1 U23076 ( .A(n19994), .B(n19993), .S(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n20000) );
  INV_X1 U23077 ( .A(n20013), .ZN(n19998) );
  INV_X1 U23078 ( .A(n19995), .ZN(n19996) );
  NAND3_X1 U23079 ( .A1(n19998), .A2(n19997), .A3(n19996), .ZN(n19999) );
  OAI211_X1 U23080 ( .C1(n20019), .C2(n20150), .A(n20000), .B(n19999), .ZN(
        n20154) );
  OAI22_X1 U23081 ( .A1(n20001), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n20154), .B2(n20025), .ZN(n20012) );
  INV_X1 U23082 ( .A(n20012), .ZN(n20010) );
  NOR2_X1 U23083 ( .A1(n20003), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20005) );
  NAND3_X1 U23084 ( .A1(n20003), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20004) );
  OAI21_X1 U23085 ( .B1(n20006), .B2(n20005), .A(n20004), .ZN(n20008) );
  OAI21_X1 U23086 ( .B1(n20025), .B2(n20008), .A(n20007), .ZN(n20009) );
  AOI222_X1 U23087 ( .A1(n20011), .A2(n20010), .B1(n20011), .B2(n20009), .C1(
        n20010), .C2(n20009), .ZN(n20030) );
  OAI221_X1 U23088 ( .B1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C1(
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .C2(n20030), .A(n20012), .ZN(
        n20032) );
  NAND2_X1 U23089 ( .A1(n9798), .A2(n20013), .ZN(n20016) );
  AOI22_X1 U23090 ( .A1(n20017), .A2(n20016), .B1(n20015), .B2(n20014), .ZN(
        n20018) );
  OAI221_X1 U23091 ( .B1(n20020), .B2(n20019), .C1(n20020), .C2(n10378), .A(
        n20018), .ZN(n20169) );
  NAND2_X1 U23092 ( .A1(n20022), .A2(n20021), .ZN(n20029) );
  AOI211_X1 U23093 ( .C1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .C2(n20025), .A(
        n20024), .B(n20023), .ZN(n20028) );
  OAI21_X1 U23094 ( .B1(P3_MORE_REG_SCAN_IN), .B2(P3_FLUSH_REG_SCAN_IN), .A(
        n20026), .ZN(n20027) );
  OAI211_X1 U23095 ( .C1(n20030), .C2(n20029), .A(n20028), .B(n20027), .ZN(
        n20031) );
  AOI211_X1 U23096 ( .C1(n20033), .C2(n20032), .A(n20169), .B(n20031), .ZN(
        n20043) );
  NAND2_X1 U23097 ( .A1(n20172), .A2(n18851), .ZN(n20050) );
  OAI211_X1 U23098 ( .C1(n20035), .C2(n20034), .A(n20179), .B(n20043), .ZN(
        n20047) );
  AND2_X1 U23099 ( .A1(n20047), .A2(P3_STATE2_REG_0__SCAN_IN), .ZN(n20139) );
  NAND2_X1 U23100 ( .A1(n20172), .A2(n20187), .ZN(n20045) );
  INV_X1 U23101 ( .A(n20036), .ZN(n20037) );
  NAND3_X1 U23102 ( .A1(n20139), .A2(n20045), .A3(n20037), .ZN(n20038) );
  OAI211_X1 U23103 ( .C1(n20174), .C2(n20039), .A(n20050), .B(n20038), .ZN(
        n20040) );
  OAI211_X1 U23104 ( .C1(n20043), .C2(n20042), .A(n20041), .B(n20040), .ZN(
        P3_U2996) );
  OR3_X1 U23105 ( .A1(n20044), .A2(n20175), .A3(n20045), .ZN(n20052) );
  NAND4_X1 U23106 ( .A1(n20048), .A2(n20047), .A3(n20046), .A4(n20045), .ZN(
        n20049) );
  NAND4_X1 U23107 ( .A1(n20051), .A2(n20050), .A3(n20052), .A4(n20049), .ZN(
        P3_U2997) );
  AND4_X1 U23108 ( .A1(n20174), .A2(n20053), .A3(n20137), .A4(n20052), .ZN(
        P3_U2998) );
  AND2_X1 U23109 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n20055), .ZN(
        P3_U2999) );
  AND2_X1 U23110 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n20055), .ZN(
        P3_U3000) );
  AND2_X1 U23111 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n20055), .ZN(
        P3_U3001) );
  AND2_X1 U23112 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n20055), .ZN(
        P3_U3002) );
  AND2_X1 U23113 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n20055), .ZN(
        P3_U3003) );
  AND2_X1 U23114 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n20055), .ZN(
        P3_U3004) );
  INV_X1 U23115 ( .A(P3_DATAWIDTH_REG_25__SCAN_IN), .ZN(n22212) );
  NOR2_X1 U23116 ( .A1(n22212), .A2(n20136), .ZN(P3_U3005) );
  AND2_X1 U23117 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n20055), .ZN(
        P3_U3006) );
  AND2_X1 U23118 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n20055), .ZN(
        P3_U3007) );
  AND2_X1 U23119 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n20055), .ZN(
        P3_U3008) );
  AND2_X1 U23120 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n20055), .ZN(
        P3_U3009) );
  AND2_X1 U23121 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n20054), .ZN(
        P3_U3010) );
  AND2_X1 U23122 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n20054), .ZN(
        P3_U3011) );
  AND2_X1 U23123 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n20054), .ZN(
        P3_U3012) );
  AND2_X1 U23124 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n20054), .ZN(
        P3_U3013) );
  AND2_X1 U23125 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n20054), .ZN(
        P3_U3014) );
  AND2_X1 U23126 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n20054), .ZN(
        P3_U3015) );
  AND2_X1 U23127 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n20054), .ZN(
        P3_U3016) );
  AND2_X1 U23128 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n20054), .ZN(
        P3_U3017) );
  AND2_X1 U23129 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n20054), .ZN(
        P3_U3018) );
  NOR2_X1 U23130 ( .A1(n22026), .A2(n20136), .ZN(P3_U3019) );
  AND2_X1 U23131 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n20054), .ZN(
        P3_U3020) );
  AND2_X1 U23132 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n20054), .ZN(P3_U3021) );
  NOR2_X1 U23133 ( .A1(n22108), .A2(n20136), .ZN(P3_U3022) );
  AND2_X1 U23134 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n20054), .ZN(P3_U3023) );
  AND2_X1 U23135 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n20055), .ZN(P3_U3024) );
  AND2_X1 U23136 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n20055), .ZN(P3_U3025) );
  AND2_X1 U23137 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n20055), .ZN(P3_U3026) );
  AND2_X1 U23138 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n20054), .ZN(P3_U3027) );
  AND2_X1 U23139 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n20055), .ZN(P3_U3028) );
  INV_X1 U23140 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n20064) );
  AOI221_X1 U23141 ( .B1(P3_STATE_REG_1__SCAN_IN), .B2(HOLD), .C1(
        P3_STATE_REG_2__SCAN_IN), .C2(HOLD), .A(n20064), .ZN(n20057) );
  NAND2_X1 U23142 ( .A1(n20172), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n20067) );
  INV_X1 U23143 ( .A(n20067), .ZN(n20061) );
  NOR2_X1 U23144 ( .A1(n20061), .A2(n20073), .ZN(n20056) );
  AOI211_X1 U23145 ( .C1(NA), .C2(n20058), .A(n20056), .B(n20066), .ZN(n20070)
         );
  OAI22_X1 U23146 ( .A1(n20184), .A2(n20057), .B1(n20056), .B2(n20070), .ZN(
        P3_U3029) );
  NOR2_X1 U23147 ( .A1(HOLD), .A2(n20058), .ZN(n20060) );
  AOI22_X1 U23148 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n20066), .B1(n20060), 
        .B2(n20059), .ZN(n20065) );
  AND2_X1 U23149 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n20062) );
  AOI211_X1 U23150 ( .C1(n20062), .C2(n20066), .A(n20061), .B(n20170), .ZN(
        n20063) );
  OAI21_X1 U23151 ( .B1(n20065), .B2(n20064), .A(n20063), .ZN(P3_U3030) );
  NOR2_X1 U23152 ( .A1(n20066), .A2(n21020), .ZN(n20069) );
  OAI22_X1 U23153 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(NA), .B2(n20067), .ZN(n20068) );
  OAI22_X1 U23154 ( .A1(n20069), .A2(n20068), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n20072) );
  INV_X1 U23155 ( .A(n20070), .ZN(n20071) );
  OAI21_X1 U23156 ( .B1(n20073), .B2(n20072), .A(n20071), .ZN(P3_U3031) );
  INV_X1 U23157 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n20075) );
  OAI222_X1 U23158 ( .A1(n20130), .A2(n17362), .B1(n20074), .B2(n20184), .C1(
        n20075), .C2(n20116), .ZN(P3_U3032) );
  CLKBUF_X1 U23159 ( .A(n20130), .Z(n20124) );
  OAI222_X1 U23160 ( .A1(n20077), .A2(n20116), .B1(n20076), .B2(n20184), .C1(
        n20075), .C2(n20124), .ZN(P3_U3033) );
  OAI222_X1 U23161 ( .A1(n20079), .A2(n20116), .B1(n20078), .B2(n20184), .C1(
        n20077), .C2(n20124), .ZN(P3_U3034) );
  INV_X1 U23162 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n20082) );
  OAI222_X1 U23163 ( .A1(n20082), .A2(n20116), .B1(n20080), .B2(n20184), .C1(
        n20079), .C2(n20124), .ZN(P3_U3035) );
  INV_X1 U23164 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n20083) );
  OAI222_X1 U23165 ( .A1(n20124), .A2(n20082), .B1(n20081), .B2(n20184), .C1(
        n20083), .C2(n20116), .ZN(P3_U3036) );
  OAI222_X1 U23166 ( .A1(n20084), .A2(n20116), .B1(n22006), .B2(n20184), .C1(
        n20083), .C2(n20124), .ZN(P3_U3037) );
  OAI222_X1 U23167 ( .A1(n20086), .A2(n20116), .B1(n20085), .B2(n20184), .C1(
        n20084), .C2(n20130), .ZN(P3_U3038) );
  OAI222_X1 U23168 ( .A1(n22085), .A2(n20116), .B1(n20087), .B2(n20184), .C1(
        n20086), .C2(n20130), .ZN(P3_U3039) );
  INV_X1 U23169 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n20089) );
  OAI222_X1 U23170 ( .A1(n20089), .A2(n20116), .B1(n20088), .B2(n20184), .C1(
        n22085), .C2(n20130), .ZN(P3_U3040) );
  OAI222_X1 U23171 ( .A1(n20091), .A2(n20116), .B1(n20090), .B2(n20184), .C1(
        n20089), .C2(n20130), .ZN(P3_U3041) );
  INV_X1 U23172 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n20093) );
  OAI222_X1 U23173 ( .A1(n20093), .A2(n20116), .B1(n20092), .B2(n20184), .C1(
        n20091), .C2(n20130), .ZN(P3_U3042) );
  OAI222_X1 U23174 ( .A1(n20095), .A2(n20116), .B1(n20094), .B2(n20184), .C1(
        n20093), .C2(n20130), .ZN(P3_U3043) );
  OAI222_X1 U23175 ( .A1(n22146), .A2(n20116), .B1(n20096), .B2(n20184), .C1(
        n20095), .C2(n20124), .ZN(P3_U3044) );
  OAI222_X1 U23176 ( .A1(n20130), .A2(n22146), .B1(n20097), .B2(n20184), .C1(
        n20098), .C2(n20116), .ZN(P3_U3045) );
  OAI222_X1 U23177 ( .A1(n20100), .A2(n20116), .B1(n20099), .B2(n20184), .C1(
        n20098), .C2(n20124), .ZN(P3_U3046) );
  OAI222_X1 U23178 ( .A1(n20102), .A2(n20116), .B1(n20101), .B2(n20184), .C1(
        n20100), .C2(n20124), .ZN(P3_U3047) );
  OAI222_X1 U23179 ( .A1(n20104), .A2(n20116), .B1(n20103), .B2(n20184), .C1(
        n20102), .C2(n20124), .ZN(P3_U3048) );
  OAI222_X1 U23180 ( .A1(n20105), .A2(n20116), .B1(n22048), .B2(n20184), .C1(
        n20104), .C2(n20124), .ZN(P3_U3049) );
  OAI222_X1 U23181 ( .A1(n20107), .A2(n20116), .B1(n20106), .B2(n20184), .C1(
        n20105), .C2(n20124), .ZN(P3_U3050) );
  OAI222_X1 U23182 ( .A1(n20124), .A2(n20107), .B1(n22155), .B2(n20184), .C1(
        n20108), .C2(n20116), .ZN(P3_U3051) );
  OAI222_X1 U23183 ( .A1(n20110), .A2(n20116), .B1(n20109), .B2(n20184), .C1(
        n20108), .C2(n20124), .ZN(P3_U3052) );
  OAI222_X1 U23184 ( .A1(n20113), .A2(n20116), .B1(n20111), .B2(n20184), .C1(
        n20110), .C2(n20124), .ZN(P3_U3053) );
  OAI222_X1 U23185 ( .A1(n20130), .A2(n20113), .B1(n20112), .B2(n20184), .C1(
        n20114), .C2(n20116), .ZN(P3_U3054) );
  OAI222_X1 U23186 ( .A1(n20117), .A2(n20116), .B1(n20115), .B2(n20184), .C1(
        n20114), .C2(n20130), .ZN(P3_U3055) );
  OAI222_X1 U23187 ( .A1(n20118), .A2(n20116), .B1(n22195), .B2(n20184), .C1(
        n20117), .C2(n20124), .ZN(P3_U3056) );
  INV_X1 U23188 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n20120) );
  OAI222_X1 U23189 ( .A1(n20120), .A2(n20116), .B1(n20119), .B2(n20184), .C1(
        n20118), .C2(n20124), .ZN(P3_U3057) );
  OAI222_X1 U23190 ( .A1(n20123), .A2(n20116), .B1(n20121), .B2(n20184), .C1(
        n20120), .C2(n20124), .ZN(P3_U3058) );
  OAI222_X1 U23191 ( .A1(n20124), .A2(n20123), .B1(n20122), .B2(n20184), .C1(
        n20125), .C2(n20116), .ZN(P3_U3059) );
  OAI222_X1 U23192 ( .A1(n20129), .A2(n20116), .B1(n20126), .B2(n20184), .C1(
        n20125), .C2(n20124), .ZN(P3_U3060) );
  OAI222_X1 U23193 ( .A1(n20130), .A2(n20129), .B1(n20128), .B2(n20184), .C1(
        n20127), .C2(n20116), .ZN(P3_U3061) );
  OAI22_X1 U23194 ( .A1(n20185), .A2(P3_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P3_BE_N_REG_3__SCAN_IN), .B2(n20184), .ZN(n20131) );
  INV_X1 U23195 ( .A(n20131), .ZN(P3_U3274) );
  MUX2_X1 U23196 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .B(P3_BE_N_REG_2__SCAN_IN), .S(n20185), .Z(P3_U3275) );
  OAI22_X1 U23197 ( .A1(n20185), .A2(P3_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P3_BE_N_REG_1__SCAN_IN), .B2(n20184), .ZN(n20132) );
  INV_X1 U23198 ( .A(n20132), .ZN(P3_U3276) );
  OAI22_X1 U23199 ( .A1(n20185), .A2(P3_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P3_BE_N_REG_0__SCAN_IN), .B2(n20184), .ZN(n20133) );
  INV_X1 U23200 ( .A(n20133), .ZN(P3_U3277) );
  OAI21_X1 U23201 ( .B1(n20136), .B2(P3_DATAWIDTH_REG_0__SCAN_IN), .A(n20135), 
        .ZN(n20134) );
  INV_X1 U23202 ( .A(n20134), .ZN(P3_U3280) );
  INV_X1 U23203 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n22180) );
  OAI21_X1 U23204 ( .B1(n20136), .B2(n22180), .A(n20135), .ZN(P3_U3281) );
  OAI21_X1 U23205 ( .B1(n20139), .B2(n20138), .A(n20137), .ZN(P3_U3282) );
  NOR2_X1 U23206 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n20140), .ZN(
        n20143) );
  INV_X1 U23207 ( .A(n20141), .ZN(n20142) );
  AOI22_X1 U23208 ( .A1(n20144), .A2(n20143), .B1(n20151), .B2(n20142), .ZN(
        n20148) );
  AOI21_X1 U23209 ( .B1(n20188), .B2(n20145), .A(n20158), .ZN(n20147) );
  OAI22_X1 U23210 ( .A1(n20158), .A2(n20148), .B1(n20147), .B2(n20146), .ZN(
        P3_U3285) );
  INV_X1 U23211 ( .A(n20149), .ZN(n20152) );
  AOI222_X1 U23212 ( .A1(n20154), .A2(n20188), .B1(n20153), .B2(n20152), .C1(
        n20151), .C2(n20150), .ZN(n20156) );
  AOI22_X1 U23213 ( .A1(n20158), .A2(n20157), .B1(n20156), .B2(n20155), .ZN(
        P3_U3288) );
  NAND3_X1 U23214 ( .A1(n20160), .A2(n17362), .A3(n13930), .ZN(n20164) );
  OAI21_X1 U23215 ( .B1(n13930), .B2(n17362), .A(n20160), .ZN(n20159) );
  OAI21_X1 U23216 ( .B1(P3_BYTEENABLE_REG_2__SCAN_IN), .B2(n20160), .A(n20159), 
        .ZN(n20161) );
  OAI221_X1 U23217 ( .B1(P3_DATAWIDTH_REG_0__SCAN_IN), .B2(n20163), .C1(n20162), .C2(n20164), .A(n20161), .ZN(P3_U3292) );
  INV_X1 U23218 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n22017) );
  INV_X1 U23219 ( .A(n20164), .ZN(n20165) );
  AOI21_X1 U23220 ( .B1(n22017), .B2(n20166), .A(n20165), .ZN(P3_U3293) );
  INV_X1 U23221 ( .A(P3_READREQUEST_REG_SCAN_IN), .ZN(n20191) );
  OAI22_X1 U23222 ( .A1(n20185), .A2(n20191), .B1(P3_W_R_N_REG_SCAN_IN), .B2(
        n20184), .ZN(n20167) );
  INV_X1 U23223 ( .A(n20167), .ZN(P3_U3294) );
  MUX2_X1 U23224 ( .A(P3_MORE_REG_SCAN_IN), .B(n20169), .S(n20168), .Z(
        P3_U3295) );
  OAI21_X1 U23225 ( .B1(P3_STATEBS16_REG_SCAN_IN), .B2(n20171), .A(n20170), 
        .ZN(n20173) );
  AOI211_X1 U23226 ( .C1(n20189), .C2(n20173), .A(n20172), .B(n20187), .ZN(
        n20176) );
  OAI21_X1 U23227 ( .B1(n20176), .B2(n20175), .A(n20174), .ZN(n20183) );
  OAI21_X1 U23228 ( .B1(n20179), .B2(n20178), .A(n20177), .ZN(n20180) );
  AOI21_X1 U23229 ( .B1(n18851), .B2(n20181), .A(n20180), .ZN(n20182) );
  MUX2_X1 U23230 ( .A(n20183), .B(P3_REQUESTPENDING_REG_SCAN_IN), .S(n20182), 
        .Z(P3_U3296) );
  OAI22_X1 U23231 ( .A1(n20185), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .B1(
        P3_M_IO_N_REG_SCAN_IN), .B2(n20184), .ZN(n20186) );
  INV_X1 U23232 ( .A(n20186), .ZN(P3_U3297) );
  AOI21_X1 U23233 ( .B1(n20188), .B2(n20187), .A(n20190), .ZN(n20194) );
  AOI22_X1 U23234 ( .A1(n20194), .A2(n20191), .B1(n20190), .B2(n20189), .ZN(
        P3_U3298) );
  INV_X1 U23235 ( .A(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n20193) );
  AOI21_X1 U23236 ( .B1(n20194), .B2(n20193), .A(n20192), .ZN(P3_U3299) );
  NAND2_X1 U23237 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n21030), .ZN(n21019) );
  AOI22_X1 U23238 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n21019), .B1(
        P2_STATE_REG_1__SCAN_IN), .B2(n21011), .ZN(n21085) );
  AOI21_X1 U23239 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(P2_ADS_N_REG_SCAN_IN), 
        .A(n21085), .ZN(n20195) );
  INV_X1 U23240 ( .A(n20195), .ZN(P2_U2815) );
  NAND2_X1 U23241 ( .A1(n21011), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n21141) );
  AOI21_X1 U23242 ( .B1(n21011), .B2(n21030), .A(P2_D_C_N_REG_SCAN_IN), .ZN(
        n20196) );
  AOI22_X1 U23243 ( .A1(n21140), .A2(P2_CODEFETCH_REG_SCAN_IN), .B1(n20196), 
        .B2(n21141), .ZN(P2_U2817) );
  OAI21_X1 U23244 ( .B1(n21013), .B2(BS16), .A(n21085), .ZN(n21083) );
  OAI21_X1 U23245 ( .B1(n21085), .B2(n20842), .A(n21083), .ZN(P2_U2818) );
  NOR4_X1 U23246 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_11__SCAN_IN), .A3(P2_DATAWIDTH_REG_12__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_13__SCAN_IN), .ZN(n20206) );
  NOR4_X1 U23247 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_7__SCAN_IN), .A3(P2_DATAWIDTH_REG_8__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_9__SCAN_IN), .ZN(n20205) );
  AOI211_X1 U23248 ( .C1(P2_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_1__SCAN_IN), .A(P2_DATAWIDTH_REG_3__SCAN_IN), .B(
        P2_DATAWIDTH_REG_4__SCAN_IN), .ZN(n20197) );
  INV_X1 U23249 ( .A(P2_DATAWIDTH_REG_5__SCAN_IN), .ZN(n22137) );
  INV_X1 U23250 ( .A(P2_DATAWIDTH_REG_19__SCAN_IN), .ZN(n22071) );
  NAND3_X1 U23251 ( .A1(n20197), .A2(n22137), .A3(n22071), .ZN(n20203) );
  NOR4_X1 U23252 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_20__SCAN_IN), .A3(P2_DATAWIDTH_REG_21__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_22__SCAN_IN), .ZN(n20201) );
  NOR4_X1 U23253 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_15__SCAN_IN), .A3(P2_DATAWIDTH_REG_16__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_17__SCAN_IN), .ZN(n20200) );
  NOR4_X1 U23254 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n20199) );
  NOR4_X1 U23255 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_25__SCAN_IN), .A3(P2_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n20198) );
  NAND4_X1 U23256 ( .A1(n20201), .A2(n20200), .A3(n20199), .A4(n20198), .ZN(
        n20202) );
  NOR4_X1 U23257 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_2__SCAN_IN), .A3(n20203), .A4(n20202), .ZN(n20204) );
  NAND3_X1 U23258 ( .A1(n20206), .A2(n20205), .A3(n20204), .ZN(n20208) );
  NOR2_X1 U23259 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n20208), .ZN(n20210) );
  INV_X1 U23260 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20207) );
  AOI22_X1 U23261 ( .A1(n20210), .A2(n20211), .B1(n20208), .B2(n20207), .ZN(
        P2_U2820) );
  INV_X1 U23262 ( .A(n20208), .ZN(n20216) );
  NOR2_X1 U23263 ( .A1(n20216), .A2(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20209)
         );
  OR4_X1 U23264 ( .A1(n20208), .A2(P2_REIP_REG_0__SCAN_IN), .A3(
        P2_DATAWIDTH_REG_1__SCAN_IN), .A4(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n20214) );
  OAI21_X1 U23265 ( .B1(n20210), .B2(n20209), .A(n20214), .ZN(P2_U2821) );
  INV_X1 U23266 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n21084) );
  NAND2_X1 U23267 ( .A1(n20210), .A2(n21084), .ZN(n20215) );
  OAI21_X1 U23268 ( .B1(n20211), .B2(n21031), .A(n20216), .ZN(n20212) );
  OAI21_X1 U23269 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n20216), .A(n20212), 
        .ZN(n20213) );
  OAI221_X1 U23270 ( .B1(n20215), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n20215), .C2(P2_REIP_REG_0__SCAN_IN), .A(n20213), .ZN(P2_U2822) );
  INV_X1 U23271 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n22023) );
  OAI211_X1 U23272 ( .C1(n20216), .C2(n22023), .A(n20215), .B(n20214), .ZN(
        P2_U2823) );
  NAND2_X1 U23273 ( .A1(n20240), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n20218) );
  OAI211_X1 U23274 ( .C1(n21056), .C2(n20269), .A(n20218), .B(n20217), .ZN(
        n20219) );
  AOI21_X1 U23275 ( .B1(n20220), .B2(n9708), .A(n20219), .ZN(n20230) );
  NOR2_X1 U23276 ( .A1(n20233), .A2(n20221), .ZN(n20222) );
  XNOR2_X1 U23277 ( .A(n20223), .B(n20222), .ZN(n20228) );
  OAI22_X1 U23278 ( .A1(n20225), .A2(n20277), .B1(n20224), .B2(n20276), .ZN(
        n20226) );
  AOI21_X1 U23279 ( .B1(n20228), .B2(n20227), .A(n20226), .ZN(n20229) );
  OAI211_X1 U23280 ( .C1(n20231), .C2(n11305), .A(n20230), .B(n20229), .ZN(
        P2_U2839) );
  NOR2_X1 U23281 ( .A1(n20233), .A2(n20232), .ZN(n20235) );
  XOR2_X1 U23282 ( .A(n20235), .B(n20234), .Z(n20248) );
  AOI21_X1 U23283 ( .B1(n20271), .B2(P2_EBX_REG_14__SCAN_IN), .A(n20355), .ZN(
        n20236) );
  OAI21_X1 U23284 ( .B1(n20269), .B2(n21053), .A(n20236), .ZN(n20239) );
  NOR2_X1 U23285 ( .A1(n20237), .A2(n20273), .ZN(n20238) );
  AOI211_X1 U23286 ( .C1(n20240), .C2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n20239), .B(n20238), .ZN(n20247) );
  INV_X1 U23287 ( .A(n20241), .ZN(n20243) );
  AOI22_X1 U23288 ( .A1(n20245), .A2(n20244), .B1(n20243), .B2(n20242), .ZN(
        n20246) );
  OAI211_X1 U23289 ( .C1(n21006), .C2(n20248), .A(n20247), .B(n20246), .ZN(
        P2_U2841) );
  NAND2_X1 U23290 ( .A1(n20250), .A2(n20249), .ZN(n20253) );
  INV_X1 U23291 ( .A(n20251), .ZN(n20252) );
  XNOR2_X1 U23292 ( .A(n20253), .B(n20252), .ZN(n20266) );
  NAND2_X1 U23293 ( .A1(n20255), .A2(n9708), .ZN(n20258) );
  AOI21_X1 U23294 ( .B1(n20256), .B2(P2_REIP_REG_9__SCAN_IN), .A(n20355), .ZN(
        n20257) );
  OAI211_X1 U23295 ( .C1(n20260), .C2(n20259), .A(n20258), .B(n20257), .ZN(
        n20264) );
  OAI22_X1 U23296 ( .A1(n20262), .A2(n20276), .B1(n20277), .B2(n20261), .ZN(
        n20263) );
  AOI211_X1 U23297 ( .C1(P2_EBX_REG_9__SCAN_IN), .C2(n20271), .A(n20264), .B(
        n20263), .ZN(n20265) );
  OAI21_X1 U23298 ( .B1(n20266), .B2(n21006), .A(n20265), .ZN(P2_U2846) );
  XOR2_X1 U23299 ( .A(n20268), .B(n20267), .Z(n20282) );
  NOR2_X1 U23300 ( .A1(n20269), .A2(n21042), .ZN(n20270) );
  AOI211_X1 U23301 ( .C1(P2_EBX_REG_7__SCAN_IN), .C2(n20271), .A(n20355), .B(
        n20270), .ZN(n20272) );
  OAI21_X1 U23302 ( .B1(n20274), .B2(n20273), .A(n20272), .ZN(n20280) );
  OAI22_X1 U23303 ( .A1(n20278), .A2(n20277), .B1(n20276), .B2(n20275), .ZN(
        n20279) );
  AOI211_X1 U23304 ( .C1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .C2(n20240), .A(
        n20280), .B(n20279), .ZN(n20281) );
  OAI21_X1 U23305 ( .B1(n20282), .B2(n21006), .A(n20281), .ZN(P2_U2848) );
  INV_X1 U23306 ( .A(n20283), .ZN(n20284) );
  AOI22_X1 U23307 ( .A1(n20285), .A2(n20284), .B1(P2_EAX_REG_8__SCAN_IN), .B2(
        n20303), .ZN(n20286) );
  OAI21_X1 U23308 ( .B1(n20287), .B2(n20311), .A(n20286), .ZN(P2_U2911) );
  AOI22_X1 U23309 ( .A1(n20288), .A2(n20304), .B1(P2_EAX_REG_3__SCAN_IN), .B2(
        n20303), .ZN(n20294) );
  AOI21_X1 U23310 ( .B1(n20291), .B2(n20290), .A(n20289), .ZN(n20292) );
  OR2_X1 U23311 ( .A1(n20292), .A2(n20298), .ZN(n20293) );
  OAI211_X1 U23312 ( .C1(n20408), .C2(n20311), .A(n20294), .B(n20293), .ZN(
        P2_U2916) );
  AOI22_X1 U23313 ( .A1(n20304), .A2(n20295), .B1(P2_EAX_REG_1__SCAN_IN), .B2(
        n20303), .ZN(n20301) );
  AOI21_X1 U23314 ( .B1(n20305), .B2(n20297), .A(n20296), .ZN(n20299) );
  OR2_X1 U23315 ( .A1(n20299), .A2(n20298), .ZN(n20300) );
  OAI211_X1 U23316 ( .C1(n20393), .C2(n20311), .A(n20301), .B(n20300), .ZN(
        P2_U2918) );
  INV_X1 U23317 ( .A(n20302), .ZN(n20308) );
  AOI22_X1 U23318 ( .A1(n20304), .A2(n20308), .B1(P2_EAX_REG_0__SCAN_IN), .B2(
        n20303), .ZN(n20310) );
  INV_X1 U23319 ( .A(n20305), .ZN(n20307) );
  OAI211_X1 U23320 ( .C1(n21111), .C2(n20308), .A(n20307), .B(n20306), .ZN(
        n20309) );
  OAI211_X1 U23321 ( .C1(n20381), .C2(n20311), .A(n20310), .B(n20309), .ZN(
        P2_U2919) );
  NOR2_X1 U23322 ( .A1(n20347), .A2(n20312), .ZN(P2_U2920) );
  AOI22_X1 U23323 ( .A1(n20313), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n20344), 
        .B2(P2_UWORD_REG_14__SCAN_IN), .ZN(n20314) );
  OAI21_X1 U23324 ( .B1(n22204), .B2(n20347), .A(n20314), .ZN(P2_U2921) );
  AOI22_X1 U23325 ( .A1(n20340), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n20344), 
        .B2(P2_LWORD_REG_15__SCAN_IN), .ZN(n20315) );
  OAI21_X1 U23326 ( .B1(n20316), .B2(n20343), .A(n20315), .ZN(P2_U2936) );
  INV_X1 U23327 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n20318) );
  AOI22_X1 U23328 ( .A1(n20340), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n20344), 
        .B2(P2_LWORD_REG_14__SCAN_IN), .ZN(n20317) );
  OAI21_X1 U23329 ( .B1(n20318), .B2(n20343), .A(n20317), .ZN(P2_U2937) );
  AOI22_X1 U23330 ( .A1(n20340), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n20344), 
        .B2(P2_LWORD_REG_13__SCAN_IN), .ZN(n20319) );
  OAI21_X1 U23331 ( .B1(n20320), .B2(n20343), .A(n20319), .ZN(P2_U2938) );
  AOI22_X1 U23332 ( .A1(n20340), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n20344), 
        .B2(P2_LWORD_REG_12__SCAN_IN), .ZN(n20321) );
  OAI21_X1 U23333 ( .B1(n22072), .B2(n20343), .A(n20321), .ZN(P2_U2939) );
  AOI22_X1 U23334 ( .A1(n20340), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n20344), 
        .B2(P2_LWORD_REG_11__SCAN_IN), .ZN(n20322) );
  OAI21_X1 U23335 ( .B1(n20323), .B2(n20343), .A(n20322), .ZN(P2_U2940) );
  AOI22_X1 U23336 ( .A1(n20340), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n20344), 
        .B2(P2_LWORD_REG_10__SCAN_IN), .ZN(n20324) );
  OAI21_X1 U23337 ( .B1(n22102), .B2(n20343), .A(n20324), .ZN(P2_U2941) );
  AOI22_X1 U23338 ( .A1(n20340), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n20344), 
        .B2(P2_LWORD_REG_9__SCAN_IN), .ZN(n20325) );
  OAI21_X1 U23339 ( .B1(n20326), .B2(n20343), .A(n20325), .ZN(P2_U2942) );
  INV_X1 U23340 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n20328) );
  AOI22_X1 U23341 ( .A1(n20340), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n20344), 
        .B2(P2_LWORD_REG_8__SCAN_IN), .ZN(n20327) );
  OAI21_X1 U23342 ( .B1(n20328), .B2(n20343), .A(n20327), .ZN(P2_U2943) );
  AOI22_X1 U23343 ( .A1(n20340), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n20344), 
        .B2(P2_LWORD_REG_7__SCAN_IN), .ZN(n20329) );
  OAI21_X1 U23344 ( .B1(n20330), .B2(n20343), .A(n20329), .ZN(P2_U2944) );
  AOI22_X1 U23345 ( .A1(n20340), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n20344), 
        .B2(P2_LWORD_REG_6__SCAN_IN), .ZN(n20331) );
  OAI21_X1 U23346 ( .B1(n20332), .B2(n20343), .A(n20331), .ZN(P2_U2945) );
  INV_X1 U23347 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n20334) );
  AOI22_X1 U23348 ( .A1(n20340), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n20344), 
        .B2(P2_LWORD_REG_5__SCAN_IN), .ZN(n20333) );
  OAI21_X1 U23349 ( .B1(n20334), .B2(n20343), .A(n20333), .ZN(P2_U2946) );
  AOI22_X1 U23350 ( .A1(n20340), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n20344), 
        .B2(P2_LWORD_REG_4__SCAN_IN), .ZN(n20335) );
  OAI21_X1 U23351 ( .B1(n16511), .B2(n20343), .A(n20335), .ZN(P2_U2947) );
  INV_X1 U23352 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n20337) );
  AOI22_X1 U23353 ( .A1(n20340), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(n20344), 
        .B2(P2_LWORD_REG_3__SCAN_IN), .ZN(n20336) );
  OAI21_X1 U23354 ( .B1(n20337), .B2(n20343), .A(n20336), .ZN(P2_U2948) );
  AOI22_X1 U23355 ( .A1(n20340), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(n20344), 
        .B2(P2_LWORD_REG_2__SCAN_IN), .ZN(n20338) );
  OAI21_X1 U23356 ( .B1(n20339), .B2(n20343), .A(n20338), .ZN(P2_U2949) );
  INV_X1 U23357 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n20342) );
  AOI22_X1 U23358 ( .A1(n20340), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(n20344), 
        .B2(P2_LWORD_REG_1__SCAN_IN), .ZN(n20341) );
  OAI21_X1 U23359 ( .B1(n20342), .B2(n20343), .A(n20341), .ZN(P2_U2950) );
  INV_X1 U23360 ( .A(n20343), .ZN(n20345) );
  AOI22_X1 U23361 ( .A1(n20345), .A2(P2_EAX_REG_0__SCAN_IN), .B1(n20344), .B2(
        P2_LWORD_REG_0__SCAN_IN), .ZN(n20346) );
  OAI21_X1 U23362 ( .B1(n22173), .B2(n20347), .A(n20346), .ZN(P2_U2951) );
  AOI22_X1 U23363 ( .A1(n20352), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(
        P2_EAX_REG_30__SCAN_IN), .B2(n20348), .ZN(n20351) );
  NAND2_X1 U23364 ( .A1(n20350), .A2(n20349), .ZN(n20353) );
  NAND2_X1 U23365 ( .A1(n20351), .A2(n20353), .ZN(P2_U2966) );
  AOI22_X1 U23366 ( .A1(n20352), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(
        P2_EAX_REG_14__SCAN_IN), .B2(n20348), .ZN(n20354) );
  NAND2_X1 U23367 ( .A1(n20354), .A2(n20353), .ZN(P2_U2981) );
  AOI22_X1 U23368 ( .A1(n20356), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        P2_REIP_REG_4__SCAN_IN), .B2(n20355), .ZN(n20366) );
  NAND2_X1 U23369 ( .A1(n20358), .A2(n20357), .ZN(n20361) );
  NAND2_X1 U23370 ( .A1(n20359), .A2(n11457), .ZN(n20360) );
  OAI211_X1 U23371 ( .C1(n20363), .C2(n20362), .A(n20361), .B(n20360), .ZN(
        n20364) );
  INV_X1 U23372 ( .A(n20364), .ZN(n20365) );
  OAI211_X1 U23373 ( .C1(n20368), .C2(n20367), .A(n20366), .B(n20365), .ZN(
        P2_U3010) );
  NAND2_X1 U23374 ( .A1(n20436), .A2(BUF2_REG_16__SCAN_IN), .ZN(n20372) );
  NAND2_X1 U23375 ( .A1(n20437), .A2(BUF1_REG_16__SCAN_IN), .ZN(n20371) );
  NAND2_X1 U23376 ( .A1(n20436), .A2(BUF2_REG_24__SCAN_IN), .ZN(n20375) );
  NAND2_X1 U23377 ( .A1(n20437), .A2(BUF1_REG_24__SCAN_IN), .ZN(n20374) );
  NOR2_X1 U23378 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20483), .ZN(
        n20448) );
  OR2_X1 U23379 ( .A1(n20441), .A2(n9731), .ZN(n20876) );
  AOI22_X1 U23380 ( .A1(n20995), .A2(n20952), .B1(n20442), .B2(n20949), .ZN(
        n20388) );
  INV_X1 U23381 ( .A(n20477), .ZN(n20377) );
  OAI21_X1 U23382 ( .B1(n20377), .B2(n20995), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n20378) );
  NAND2_X1 U23383 ( .A1(n20378), .A2(n20880), .ZN(n20386) );
  NOR2_X1 U23384 ( .A1(n20386), .A2(n20991), .ZN(n20379) );
  AOI211_X1 U23385 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n20382), .A(
        P2_STATE2_REG_3__SCAN_IN), .B(n20379), .ZN(n20380) );
  OAI21_X1 U23386 ( .B1(n20380), .B2(n20442), .A(n20941), .ZN(n20445) );
  NOR2_X2 U23387 ( .A1(n20811), .A2(n20381), .ZN(n20950) );
  NOR2_X1 U23388 ( .A1(n20991), .A2(n20442), .ZN(n20385) );
  INV_X1 U23389 ( .A(n20382), .ZN(n20383) );
  OAI21_X1 U23390 ( .B1(n20383), .B2(n20442), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20384) );
  AOI22_X1 U23391 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20445), .B1(
        n20950), .B2(n20444), .ZN(n20387) );
  OAI211_X1 U23392 ( .C1(n20894), .C2(n20477), .A(n20388), .B(n20387), .ZN(
        P2_U3048) );
  NAND2_X1 U23393 ( .A1(n20436), .A2(BUF2_REG_17__SCAN_IN), .ZN(n20390) );
  NAND2_X1 U23394 ( .A1(n20437), .A2(BUF1_REG_17__SCAN_IN), .ZN(n20389) );
  NAND2_X1 U23395 ( .A1(n20436), .A2(BUF2_REG_25__SCAN_IN), .ZN(n20392) );
  NAND2_X1 U23396 ( .A1(n20437), .A2(BUF1_REG_25__SCAN_IN), .ZN(n20391) );
  AOI22_X1 U23397 ( .A1(n20995), .A2(n20848), .B1(n20442), .B2(n20957), .ZN(
        n20395) );
  NOR2_X2 U23398 ( .A1(n20811), .A2(n20393), .ZN(n20958) );
  AOI22_X1 U23399 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20445), .B1(
        n20958), .B2(n20444), .ZN(n20394) );
  OAI211_X1 U23400 ( .C1(n20899), .C2(n20477), .A(n20395), .B(n20394), .ZN(
        P2_U3049) );
  NAND2_X1 U23401 ( .A1(n20436), .A2(BUF2_REG_18__SCAN_IN), .ZN(n20397) );
  NAND2_X1 U23402 ( .A1(n20437), .A2(BUF1_REG_18__SCAN_IN), .ZN(n20396) );
  NAND2_X1 U23403 ( .A1(n20436), .A2(BUF2_REG_26__SCAN_IN), .ZN(n20399) );
  NAND2_X1 U23404 ( .A1(n20437), .A2(BUF1_REG_26__SCAN_IN), .ZN(n20398) );
  OR2_X1 U23405 ( .A1(n20441), .A2(n20400), .ZN(n20900) );
  AOI22_X1 U23406 ( .A1(n20995), .A2(n20851), .B1(n20442), .B2(n20964), .ZN(
        n20403) );
  NOR2_X2 U23407 ( .A1(n20811), .A2(n20401), .ZN(n20965) );
  AOI22_X1 U23408 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20445), .B1(
        n20965), .B2(n20444), .ZN(n20402) );
  OAI211_X1 U23409 ( .C1(n20901), .C2(n20477), .A(n20403), .B(n20402), .ZN(
        P2_U3050) );
  NAND2_X1 U23410 ( .A1(n20436), .A2(BUF2_REG_19__SCAN_IN), .ZN(n20405) );
  NAND2_X1 U23411 ( .A1(n20437), .A2(BUF1_REG_19__SCAN_IN), .ZN(n20404) );
  NAND2_X1 U23412 ( .A1(n20436), .A2(BUF2_REG_27__SCAN_IN), .ZN(n20407) );
  NAND2_X1 U23413 ( .A1(n20437), .A2(BUF1_REG_27__SCAN_IN), .ZN(n20406) );
  OR2_X1 U23414 ( .A1(n20441), .A2(n10895), .ZN(n20905) );
  AOI22_X1 U23415 ( .A1(n20995), .A2(n20854), .B1(n20442), .B2(n20970), .ZN(
        n20410) );
  NOR2_X2 U23416 ( .A1(n20811), .A2(n20408), .ZN(n20971) );
  AOI22_X1 U23417 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20445), .B1(
        n20971), .B2(n20444), .ZN(n20409) );
  OAI211_X1 U23418 ( .C1(n20906), .C2(n20477), .A(n20410), .B(n20409), .ZN(
        P2_U3051) );
  NAND2_X1 U23419 ( .A1(n20436), .A2(BUF2_REG_20__SCAN_IN), .ZN(n20412) );
  NAND2_X1 U23420 ( .A1(n20437), .A2(BUF1_REG_20__SCAN_IN), .ZN(n20411) );
  NAND2_X1 U23421 ( .A1(n20436), .A2(BUF2_REG_28__SCAN_IN), .ZN(n20414) );
  NAND2_X1 U23422 ( .A1(n20437), .A2(BUF1_REG_28__SCAN_IN), .ZN(n20413) );
  OR2_X1 U23423 ( .A1(n20441), .A2(n20415), .ZN(n20910) );
  AOI22_X1 U23424 ( .A1(n20995), .A2(n20857), .B1(n20442), .B2(n21919), .ZN(
        n20418) );
  NOR2_X2 U23425 ( .A1(n20811), .A2(n20416), .ZN(n21920) );
  AOI22_X1 U23426 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20445), .B1(
        n21920), .B2(n20444), .ZN(n20417) );
  OAI211_X1 U23427 ( .C1(n20914), .C2(n20477), .A(n20418), .B(n20417), .ZN(
        P2_U3052) );
  NAND2_X1 U23428 ( .A1(n20436), .A2(BUF2_REG_21__SCAN_IN), .ZN(n20420) );
  NAND2_X1 U23429 ( .A1(n20437), .A2(BUF1_REG_21__SCAN_IN), .ZN(n20419) );
  NAND2_X1 U23430 ( .A1(n20436), .A2(BUF2_REG_29__SCAN_IN), .ZN(n20422) );
  NAND2_X1 U23431 ( .A1(n20437), .A2(BUF1_REG_29__SCAN_IN), .ZN(n20421) );
  AOI22_X1 U23432 ( .A1(n20995), .A2(n20860), .B1(n20442), .B2(n20978), .ZN(
        n20426) );
  INV_X1 U23433 ( .A(n20423), .ZN(n20424) );
  NOR2_X2 U23434 ( .A1(n20811), .A2(n20424), .ZN(n20979) );
  AOI22_X1 U23435 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20445), .B1(
        n20979), .B2(n20444), .ZN(n20425) );
  OAI211_X1 U23436 ( .C1(n20916), .C2(n20477), .A(n20426), .B(n20425), .ZN(
        P2_U3053) );
  NAND2_X1 U23437 ( .A1(n20436), .A2(BUF2_REG_22__SCAN_IN), .ZN(n20428) );
  NAND2_X1 U23438 ( .A1(n20437), .A2(BUF1_REG_22__SCAN_IN), .ZN(n20427) );
  NAND2_X1 U23439 ( .A1(n20436), .A2(BUF2_REG_30__SCAN_IN), .ZN(n20430) );
  NAND2_X1 U23440 ( .A1(n20437), .A2(BUF1_REG_30__SCAN_IN), .ZN(n20429) );
  OR2_X1 U23441 ( .A1(n20441), .A2(n10900), .ZN(n20920) );
  AOI22_X1 U23442 ( .A1(n20995), .A2(n20863), .B1(n20442), .B2(n20984), .ZN(
        n20433) );
  NOR2_X2 U23443 ( .A1(n20811), .A2(n20431), .ZN(n20985) );
  AOI22_X1 U23444 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20445), .B1(
        n20985), .B2(n20444), .ZN(n20432) );
  OAI211_X1 U23445 ( .C1(n20921), .C2(n20477), .A(n20433), .B(n20432), .ZN(
        P2_U3054) );
  NAND2_X1 U23446 ( .A1(n20436), .A2(BUF2_REG_23__SCAN_IN), .ZN(n20435) );
  NAND2_X1 U23447 ( .A1(n20437), .A2(BUF1_REG_23__SCAN_IN), .ZN(n20434) );
  NAND2_X1 U23448 ( .A1(n20436), .A2(BUF2_REG_31__SCAN_IN), .ZN(n20439) );
  NAND2_X1 U23449 ( .A1(n20437), .A2(BUF1_REG_31__SCAN_IN), .ZN(n20438) );
  AOI22_X1 U23450 ( .A1(n20995), .A2(n20868), .B1(n20442), .B2(n20990), .ZN(
        n20447) );
  NOR2_X2 U23451 ( .A1(n20811), .A2(n20443), .ZN(n20992) );
  AOI22_X1 U23452 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20445), .B1(
        n20992), .B2(n20444), .ZN(n20446) );
  OAI211_X1 U23453 ( .C1(n20927), .C2(n20477), .A(n20447), .B(n20446), .ZN(
        P2_U3055) );
  INV_X1 U23454 ( .A(n20448), .ZN(n20454) );
  INV_X1 U23455 ( .A(n20449), .ZN(n20450) );
  OR2_X1 U23456 ( .A1(n20838), .A2(n20483), .ZN(n20452) );
  NAND3_X1 U23457 ( .A1(n20450), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(n20452), 
        .ZN(n20453) );
  INV_X1 U23458 ( .A(n20453), .ZN(n20451) );
  OAI22_X1 U23459 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n20454), .B1(n20451), 
        .B2(n20945), .ZN(n20473) );
  AOI22_X1 U23460 ( .A1(n20473), .A2(n20950), .B1(n20949), .B2(n20472), .ZN(
        n20459) );
  NAND3_X1 U23461 ( .A1(n21090), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n21099), 
        .ZN(n20577) );
  NAND2_X1 U23462 ( .A1(n21100), .A2(n20453), .ZN(n20455) );
  OAI21_X1 U23463 ( .B1(n20577), .B2(n20455), .A(n20454), .ZN(n20456) );
  OAI211_X1 U23464 ( .C1(n20472), .C2(n21106), .A(n20456), .B(n20941), .ZN(
        n20474) );
  AOI22_X1 U23465 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20474), .B1(
        n20502), .B2(n20951), .ZN(n20458) );
  OAI211_X1 U23466 ( .C1(n20877), .C2(n20477), .A(n20459), .B(n20458), .ZN(
        P2_U3056) );
  AOI22_X1 U23467 ( .A1(n20473), .A2(n20958), .B1(n20957), .B2(n20472), .ZN(
        n20461) );
  AOI22_X1 U23468 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20474), .B1(
        n20502), .B2(n20960), .ZN(n20460) );
  OAI211_X1 U23469 ( .C1(n20963), .C2(n20477), .A(n20461), .B(n20460), .ZN(
        P2_U3057) );
  AOI22_X1 U23470 ( .A1(n20473), .A2(n20965), .B1(n20964), .B2(n20472), .ZN(
        n20463) );
  AOI22_X1 U23471 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20474), .B1(
        n20502), .B2(n20966), .ZN(n20462) );
  OAI211_X1 U23472 ( .C1(n20969), .C2(n20477), .A(n20463), .B(n20462), .ZN(
        P2_U3058) );
  AOI22_X1 U23473 ( .A1(n20473), .A2(n20971), .B1(n20970), .B2(n20472), .ZN(
        n20465) );
  AOI22_X1 U23474 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20474), .B1(
        n20502), .B2(n20972), .ZN(n20464) );
  OAI211_X1 U23475 ( .C1(n20975), .C2(n20477), .A(n20465), .B(n20464), .ZN(
        P2_U3059) );
  AOI22_X1 U23476 ( .A1(n20473), .A2(n21920), .B1(n21919), .B2(n20472), .ZN(
        n20467) );
  AOI22_X1 U23477 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20474), .B1(
        n20502), .B2(n21922), .ZN(n20466) );
  OAI211_X1 U23478 ( .C1(n21928), .C2(n20477), .A(n20467), .B(n20466), .ZN(
        P2_U3060) );
  AOI22_X1 U23479 ( .A1(n20473), .A2(n20979), .B1(n20978), .B2(n20472), .ZN(
        n20469) );
  AOI22_X1 U23480 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20474), .B1(
        n20502), .B2(n20980), .ZN(n20468) );
  OAI211_X1 U23481 ( .C1(n20983), .C2(n20477), .A(n20469), .B(n20468), .ZN(
        P2_U3061) );
  AOI22_X1 U23482 ( .A1(n20473), .A2(n20985), .B1(n20984), .B2(n20472), .ZN(
        n20471) );
  AOI22_X1 U23483 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20474), .B1(
        n20502), .B2(n20986), .ZN(n20470) );
  OAI211_X1 U23484 ( .C1(n20989), .C2(n20477), .A(n20471), .B(n20470), .ZN(
        P2_U3062) );
  AOI22_X1 U23485 ( .A1(n20473), .A2(n20992), .B1(n20990), .B2(n20472), .ZN(
        n20476) );
  AOI22_X1 U23486 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20474), .B1(
        n20502), .B2(n20994), .ZN(n20475) );
  OAI211_X1 U23487 ( .C1(n21000), .C2(n20477), .A(n20476), .B(n20475), .ZN(
        P2_U3063) );
  NOR2_X1 U23488 ( .A1(n20874), .A2(n20483), .ZN(n20500) );
  INV_X1 U23489 ( .A(n20500), .ZN(n20478) );
  AND2_X1 U23490 ( .A1(n20481), .A2(n20478), .ZN(n20480) );
  INV_X1 U23491 ( .A(n20479), .ZN(n20751) );
  OAI22_X1 U23492 ( .A1(n20480), .A2(n20945), .B1(n20751), .B2(n20483), .ZN(
        n20501) );
  AOI22_X1 U23493 ( .A1(n20501), .A2(n20950), .B1(n20949), .B2(n20500), .ZN(
        n20487) );
  AOI21_X1 U23494 ( .B1(n20481), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n20485) );
  INV_X1 U23495 ( .A(n20882), .ZN(n20808) );
  OAI21_X1 U23496 ( .B1(n20502), .B2(n20531), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n20482) );
  OAI21_X1 U23497 ( .B1(n20808), .B2(n20483), .A(n20482), .ZN(n20484) );
  OAI211_X1 U23498 ( .C1(n20485), .C2(n20500), .A(n20941), .B(n20484), .ZN(
        n20503) );
  AOI22_X1 U23499 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20503), .B1(
        n20502), .B2(n20952), .ZN(n20486) );
  OAI211_X1 U23500 ( .C1(n20894), .C2(n20540), .A(n20487), .B(n20486), .ZN(
        P2_U3064) );
  AOI22_X1 U23501 ( .A1(n20501), .A2(n20958), .B1(n20957), .B2(n20500), .ZN(
        n20489) );
  AOI22_X1 U23502 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20503), .B1(
        n20502), .B2(n20848), .ZN(n20488) );
  OAI211_X1 U23503 ( .C1(n20899), .C2(n20540), .A(n20489), .B(n20488), .ZN(
        P2_U3065) );
  AOI22_X1 U23504 ( .A1(n20501), .A2(n20965), .B1(n20964), .B2(n20500), .ZN(
        n20491) );
  AOI22_X1 U23505 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20503), .B1(
        n20502), .B2(n20851), .ZN(n20490) );
  OAI211_X1 U23506 ( .C1(n20901), .C2(n20540), .A(n20491), .B(n20490), .ZN(
        P2_U3066) );
  AOI22_X1 U23507 ( .A1(n20501), .A2(n20971), .B1(n20970), .B2(n20500), .ZN(
        n20493) );
  AOI22_X1 U23508 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20503), .B1(
        n20502), .B2(n20854), .ZN(n20492) );
  OAI211_X1 U23509 ( .C1(n20906), .C2(n20540), .A(n20493), .B(n20492), .ZN(
        P2_U3067) );
  AOI22_X1 U23510 ( .A1(n20501), .A2(n21920), .B1(n21919), .B2(n20500), .ZN(
        n20495) );
  AOI22_X1 U23511 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20503), .B1(
        n20502), .B2(n20857), .ZN(n20494) );
  OAI211_X1 U23512 ( .C1(n20914), .C2(n20540), .A(n20495), .B(n20494), .ZN(
        P2_U3068) );
  AOI22_X1 U23513 ( .A1(n20501), .A2(n20979), .B1(n20978), .B2(n20500), .ZN(
        n20497) );
  AOI22_X1 U23514 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20503), .B1(
        n20502), .B2(n20860), .ZN(n20496) );
  OAI211_X1 U23515 ( .C1(n20916), .C2(n20540), .A(n20497), .B(n20496), .ZN(
        P2_U3069) );
  AOI22_X1 U23516 ( .A1(n20501), .A2(n20985), .B1(n20984), .B2(n20500), .ZN(
        n20499) );
  AOI22_X1 U23517 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20503), .B1(
        n20502), .B2(n20863), .ZN(n20498) );
  OAI211_X1 U23518 ( .C1(n20921), .C2(n20540), .A(n20499), .B(n20498), .ZN(
        P2_U3070) );
  AOI22_X1 U23519 ( .A1(n20501), .A2(n20992), .B1(n20990), .B2(n20500), .ZN(
        n20505) );
  AOI22_X1 U23520 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20503), .B1(
        n20502), .B2(n20868), .ZN(n20504) );
  OAI211_X1 U23521 ( .C1(n20927), .C2(n20540), .A(n20505), .B(n20504), .ZN(
        P2_U3071) );
  NAND2_X1 U23522 ( .A1(n20782), .A2(n20508), .ZN(n20534) );
  INV_X1 U23523 ( .A(n20534), .ZN(n20530) );
  AOI22_X1 U23524 ( .A1(n20531), .A2(n20952), .B1(n20949), .B2(n20530), .ZN(
        n20517) );
  INV_X1 U23525 ( .A(n20506), .ZN(n20507) );
  NAND2_X1 U23526 ( .A1(n20672), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n21087) );
  OAI21_X1 U23527 ( .B1(n20507), .B2(n21087), .A(n20880), .ZN(n20515) );
  AND2_X1 U23528 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20508), .ZN(
        n20512) );
  INV_X1 U23529 ( .A(n20509), .ZN(n20510) );
  OAI211_X1 U23530 ( .C1(n20510), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n20883), 
        .B(n20534), .ZN(n20511) );
  OAI211_X1 U23531 ( .C1(n20515), .C2(n20512), .A(n20941), .B(n20511), .ZN(
        n20537) );
  INV_X1 U23532 ( .A(n20512), .ZN(n20514) );
  OAI21_X1 U23533 ( .B1(n20509), .B2(n20530), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20513) );
  AOI22_X1 U23534 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20537), .B1(
        n20950), .B2(n20536), .ZN(n20516) );
  OAI211_X1 U23535 ( .C1(n20894), .C2(n20547), .A(n20517), .B(n20516), .ZN(
        P2_U3072) );
  OAI22_X1 U23536 ( .A1(n20547), .A2(n20899), .B1(n20895), .B2(n20534), .ZN(
        n20518) );
  INV_X1 U23537 ( .A(n20518), .ZN(n20520) );
  AOI22_X1 U23538 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20537), .B1(
        n20958), .B2(n20536), .ZN(n20519) );
  OAI211_X1 U23539 ( .C1(n20963), .C2(n20540), .A(n20520), .B(n20519), .ZN(
        P2_U3073) );
  AOI22_X1 U23540 ( .A1(n20531), .A2(n20851), .B1(n20964), .B2(n20530), .ZN(
        n20522) );
  AOI22_X1 U23541 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20537), .B1(
        n20965), .B2(n20536), .ZN(n20521) );
  OAI211_X1 U23542 ( .C1(n20901), .C2(n20547), .A(n20522), .B(n20521), .ZN(
        P2_U3074) );
  OAI22_X1 U23543 ( .A1(n20547), .A2(n20906), .B1(n20905), .B2(n20534), .ZN(
        n20523) );
  INV_X1 U23544 ( .A(n20523), .ZN(n20525) );
  AOI22_X1 U23545 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20537), .B1(
        n20971), .B2(n20536), .ZN(n20524) );
  OAI211_X1 U23546 ( .C1(n20975), .C2(n20540), .A(n20525), .B(n20524), .ZN(
        P2_U3075) );
  AOI22_X1 U23547 ( .A1(n20531), .A2(n20857), .B1(n21919), .B2(n20530), .ZN(
        n20527) );
  AOI22_X1 U23548 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20537), .B1(
        n21920), .B2(n20536), .ZN(n20526) );
  OAI211_X1 U23549 ( .C1(n20914), .C2(n20547), .A(n20527), .B(n20526), .ZN(
        P2_U3076) );
  AOI22_X1 U23550 ( .A1(n20531), .A2(n20860), .B1(n20978), .B2(n20530), .ZN(
        n20529) );
  AOI22_X1 U23551 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20537), .B1(
        n20979), .B2(n20536), .ZN(n20528) );
  OAI211_X1 U23552 ( .C1(n20916), .C2(n20547), .A(n20529), .B(n20528), .ZN(
        P2_U3077) );
  AOI22_X1 U23553 ( .A1(n20531), .A2(n20863), .B1(n20984), .B2(n20530), .ZN(
        n20533) );
  AOI22_X1 U23554 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20537), .B1(
        n20985), .B2(n20536), .ZN(n20532) );
  OAI211_X1 U23555 ( .C1(n20921), .C2(n20547), .A(n20533), .B(n20532), .ZN(
        P2_U3078) );
  OAI22_X1 U23556 ( .A1(n20547), .A2(n20927), .B1(n20926), .B2(n20534), .ZN(
        n20535) );
  INV_X1 U23557 ( .A(n20535), .ZN(n20539) );
  AOI22_X1 U23558 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20537), .B1(
        n20992), .B2(n20536), .ZN(n20538) );
  OAI211_X1 U23559 ( .C1(n21000), .C2(n20540), .A(n20539), .B(n20538), .ZN(
        P2_U3079) );
  OR2_X1 U23560 ( .A1(n21100), .A2(n20672), .ZN(n20574) );
  NOR2_X1 U23561 ( .A1(n20574), .A2(n21111), .ZN(n20541) );
  NAND2_X1 U23562 ( .A1(n20808), .A2(n21096), .ZN(n20551) );
  INV_X1 U23563 ( .A(n20542), .ZN(n20545) );
  NAND2_X1 U23564 ( .A1(n21096), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n20639) );
  NOR2_X1 U23565 ( .A1(n20639), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20579) );
  INV_X1 U23566 ( .A(n20579), .ZN(n20582) );
  OAI21_X1 U23567 ( .B1(n20543), .B2(n20568), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20544) );
  AOI22_X1 U23568 ( .A1(n20569), .A2(n20950), .B1(n20949), .B2(n20568), .ZN(
        n20555) );
  AOI21_X1 U23569 ( .B1(n20546), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n20553) );
  INV_X1 U23570 ( .A(n20807), .ZN(n20550) );
  INV_X1 U23571 ( .A(n20605), .ZN(n20548) );
  OAI21_X1 U23572 ( .B1(n20570), .B2(n20548), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n20549) );
  OAI21_X1 U23573 ( .B1(n20551), .B2(n20550), .A(n20549), .ZN(n20552) );
  OAI211_X1 U23574 ( .C1(n20568), .C2(n20553), .A(n20552), .B(n20941), .ZN(
        n20571) );
  AOI22_X1 U23575 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20571), .B1(
        n20570), .B2(n20952), .ZN(n20554) );
  OAI211_X1 U23576 ( .C1(n20894), .C2(n20605), .A(n20555), .B(n20554), .ZN(
        P2_U3080) );
  AOI22_X1 U23577 ( .A1(n20569), .A2(n20958), .B1(n20957), .B2(n20568), .ZN(
        n20557) );
  AOI22_X1 U23578 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20571), .B1(
        n20570), .B2(n20848), .ZN(n20556) );
  OAI211_X1 U23579 ( .C1(n20899), .C2(n20605), .A(n20557), .B(n20556), .ZN(
        P2_U3081) );
  AOI22_X1 U23580 ( .A1(n20569), .A2(n20965), .B1(n20964), .B2(n20568), .ZN(
        n20559) );
  AOI22_X1 U23581 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20571), .B1(
        n20570), .B2(n20851), .ZN(n20558) );
  OAI211_X1 U23582 ( .C1(n20901), .C2(n20605), .A(n20559), .B(n20558), .ZN(
        P2_U3082) );
  AOI22_X1 U23583 ( .A1(n20569), .A2(n20971), .B1(n20970), .B2(n20568), .ZN(
        n20561) );
  AOI22_X1 U23584 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20571), .B1(
        n20570), .B2(n20854), .ZN(n20560) );
  OAI211_X1 U23585 ( .C1(n20906), .C2(n20605), .A(n20561), .B(n20560), .ZN(
        P2_U3083) );
  AOI22_X1 U23586 ( .A1(n20569), .A2(n21920), .B1(n21919), .B2(n20568), .ZN(
        n20563) );
  AOI22_X1 U23587 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20571), .B1(
        n20570), .B2(n20857), .ZN(n20562) );
  OAI211_X1 U23588 ( .C1(n20914), .C2(n20605), .A(n20563), .B(n20562), .ZN(
        P2_U3084) );
  AOI22_X1 U23589 ( .A1(n20569), .A2(n20979), .B1(n20978), .B2(n20568), .ZN(
        n20565) );
  AOI22_X1 U23590 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20571), .B1(
        n20570), .B2(n20860), .ZN(n20564) );
  OAI211_X1 U23591 ( .C1(n20916), .C2(n20605), .A(n20565), .B(n20564), .ZN(
        P2_U3085) );
  AOI22_X1 U23592 ( .A1(n20569), .A2(n20985), .B1(n20984), .B2(n20568), .ZN(
        n20567) );
  AOI22_X1 U23593 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20571), .B1(
        n20570), .B2(n20863), .ZN(n20566) );
  OAI211_X1 U23594 ( .C1(n20921), .C2(n20605), .A(n20567), .B(n20566), .ZN(
        P2_U3086) );
  AOI22_X1 U23595 ( .A1(n20569), .A2(n20992), .B1(n20990), .B2(n20568), .ZN(
        n20573) );
  AOI22_X1 U23596 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20571), .B1(
        n20570), .B2(n20868), .ZN(n20572) );
  OAI211_X1 U23597 ( .C1(n20927), .C2(n20605), .A(n20573), .B(n20572), .ZN(
        P2_U3087) );
  NOR2_X1 U23598 ( .A1(n20574), .A2(n20673), .ZN(n20575) );
  NOR2_X1 U23599 ( .A1(n20838), .A2(n20639), .ZN(n20614) );
  OAI22_X1 U23600 ( .A1(n20620), .A2(n20894), .B1(n20604), .B2(n20876), .ZN(
        n20576) );
  INV_X1 U23601 ( .A(n20576), .ZN(n20585) );
  OAI21_X1 U23602 ( .B1(n20577), .B2(n21100), .A(n20880), .ZN(n20583) );
  OAI211_X1 U23603 ( .C1(n11086), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n20883), 
        .B(n20604), .ZN(n20578) );
  OAI211_X1 U23604 ( .C1(n20583), .C2(n20579), .A(n20941), .B(n20578), .ZN(
        n20608) );
  OAI21_X1 U23605 ( .B1(n20580), .B2(n20614), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20581) );
  AOI22_X1 U23606 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20608), .B1(
        n20950), .B2(n20607), .ZN(n20584) );
  OAI211_X1 U23607 ( .C1(n20877), .C2(n20605), .A(n20585), .B(n20584), .ZN(
        P2_U3088) );
  OAI22_X1 U23608 ( .A1(n20620), .A2(n20899), .B1(n20604), .B2(n20895), .ZN(
        n20586) );
  INV_X1 U23609 ( .A(n20586), .ZN(n20588) );
  AOI22_X1 U23610 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20608), .B1(
        n20958), .B2(n20607), .ZN(n20587) );
  OAI211_X1 U23611 ( .C1(n20963), .C2(n20605), .A(n20588), .B(n20587), .ZN(
        P2_U3089) );
  OAI22_X1 U23612 ( .A1(n20605), .A2(n20969), .B1(n20604), .B2(n20900), .ZN(
        n20589) );
  INV_X1 U23613 ( .A(n20589), .ZN(n20591) );
  AOI22_X1 U23614 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20608), .B1(
        n20965), .B2(n20607), .ZN(n20590) );
  OAI211_X1 U23615 ( .C1(n20901), .C2(n20620), .A(n20591), .B(n20590), .ZN(
        P2_U3090) );
  OAI22_X1 U23616 ( .A1(n20605), .A2(n20975), .B1(n20604), .B2(n20905), .ZN(
        n20592) );
  INV_X1 U23617 ( .A(n20592), .ZN(n20594) );
  AOI22_X1 U23618 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20608), .B1(
        n20971), .B2(n20607), .ZN(n20593) );
  OAI211_X1 U23619 ( .C1(n20906), .C2(n20620), .A(n20594), .B(n20593), .ZN(
        P2_U3091) );
  OAI22_X1 U23620 ( .A1(n20620), .A2(n20914), .B1(n20604), .B2(n20910), .ZN(
        n20595) );
  INV_X1 U23621 ( .A(n20595), .ZN(n20597) );
  AOI22_X1 U23622 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20608), .B1(
        n21920), .B2(n20607), .ZN(n20596) );
  OAI211_X1 U23623 ( .C1(n21928), .C2(n20605), .A(n20597), .B(n20596), .ZN(
        P2_U3092) );
  OAI22_X1 U23624 ( .A1(n20605), .A2(n20983), .B1(n20604), .B2(n20915), .ZN(
        n20598) );
  INV_X1 U23625 ( .A(n20598), .ZN(n20600) );
  AOI22_X1 U23626 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20608), .B1(
        n20979), .B2(n20607), .ZN(n20599) );
  OAI211_X1 U23627 ( .C1(n20916), .C2(n20620), .A(n20600), .B(n20599), .ZN(
        P2_U3093) );
  OAI22_X1 U23628 ( .A1(n20620), .A2(n20921), .B1(n20604), .B2(n20920), .ZN(
        n20601) );
  INV_X1 U23629 ( .A(n20601), .ZN(n20603) );
  AOI22_X1 U23630 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20608), .B1(
        n20985), .B2(n20607), .ZN(n20602) );
  OAI211_X1 U23631 ( .C1(n20989), .C2(n20605), .A(n20603), .B(n20602), .ZN(
        P2_U3094) );
  OAI22_X1 U23632 ( .A1(n20605), .A2(n21000), .B1(n20604), .B2(n20926), .ZN(
        n20606) );
  INV_X1 U23633 ( .A(n20606), .ZN(n20610) );
  AOI22_X1 U23634 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20608), .B1(
        n20992), .B2(n20607), .ZN(n20609) );
  OAI211_X1 U23635 ( .C1(n20927), .C2(n20620), .A(n20610), .B(n20609), .ZN(
        P2_U3095) );
  NOR2_X1 U23636 ( .A1(n20874), .A2(n20639), .ZN(n20633) );
  OAI21_X1 U23637 ( .B1(n20611), .B2(n20633), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20612) );
  AOI22_X1 U23638 ( .A1(n20634), .A2(n20950), .B1(n20949), .B2(n20633), .ZN(
        n20619) );
  NOR2_X1 U23639 ( .A1(n21100), .A2(n21099), .ZN(n20613) );
  AOI21_X1 U23640 ( .B1(n20670), .B2(n20620), .A(n20842), .ZN(n20615) );
  NOR2_X1 U23641 ( .A1(n20615), .A2(n20614), .ZN(n20616) );
  AOI211_X1 U23642 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n11050), .A(
        P2_STATE2_REG_3__SCAN_IN), .B(n20616), .ZN(n20617) );
  OAI21_X1 U23643 ( .B1(n20617), .B2(n20633), .A(n20941), .ZN(n20636) );
  AOI22_X1 U23644 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20636), .B1(
        n20662), .B2(n20951), .ZN(n20618) );
  OAI211_X1 U23645 ( .C1(n20877), .C2(n20620), .A(n20619), .B(n20618), .ZN(
        P2_U3096) );
  AOI22_X1 U23646 ( .A1(n20634), .A2(n20958), .B1(n20957), .B2(n20633), .ZN(
        n20622) );
  AOI22_X1 U23647 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20636), .B1(
        n20635), .B2(n20848), .ZN(n20621) );
  OAI211_X1 U23648 ( .C1(n20899), .C2(n20670), .A(n20622), .B(n20621), .ZN(
        P2_U3097) );
  AOI22_X1 U23649 ( .A1(n20634), .A2(n20965), .B1(n20964), .B2(n20633), .ZN(
        n20624) );
  AOI22_X1 U23650 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20636), .B1(
        n20635), .B2(n20851), .ZN(n20623) );
  OAI211_X1 U23651 ( .C1(n20901), .C2(n20670), .A(n20624), .B(n20623), .ZN(
        P2_U3098) );
  AOI22_X1 U23652 ( .A1(n20634), .A2(n20971), .B1(n20970), .B2(n20633), .ZN(
        n20626) );
  AOI22_X1 U23653 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20636), .B1(
        n20635), .B2(n20854), .ZN(n20625) );
  OAI211_X1 U23654 ( .C1(n20906), .C2(n20670), .A(n20626), .B(n20625), .ZN(
        P2_U3099) );
  AOI22_X1 U23655 ( .A1(n20634), .A2(n21920), .B1(n21919), .B2(n20633), .ZN(
        n20628) );
  AOI22_X1 U23656 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20636), .B1(
        n20635), .B2(n20857), .ZN(n20627) );
  OAI211_X1 U23657 ( .C1(n20914), .C2(n20670), .A(n20628), .B(n20627), .ZN(
        P2_U3100) );
  AOI22_X1 U23658 ( .A1(n20634), .A2(n20979), .B1(n20978), .B2(n20633), .ZN(
        n20630) );
  AOI22_X1 U23659 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20636), .B1(
        n20635), .B2(n20860), .ZN(n20629) );
  OAI211_X1 U23660 ( .C1(n20916), .C2(n20670), .A(n20630), .B(n20629), .ZN(
        P2_U3101) );
  AOI22_X1 U23661 ( .A1(n20634), .A2(n20985), .B1(n20984), .B2(n20633), .ZN(
        n20632) );
  AOI22_X1 U23662 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20636), .B1(
        n20635), .B2(n20863), .ZN(n20631) );
  OAI211_X1 U23663 ( .C1(n20921), .C2(n20670), .A(n20632), .B(n20631), .ZN(
        P2_U3102) );
  AOI22_X1 U23664 ( .A1(n20634), .A2(n20992), .B1(n20990), .B2(n20633), .ZN(
        n20638) );
  AOI22_X1 U23665 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20636), .B1(
        n20635), .B2(n20868), .ZN(n20637) );
  OAI211_X1 U23666 ( .C1(n20927), .C2(n20670), .A(n20638), .B(n20637), .ZN(
        P2_U3103) );
  INV_X1 U23667 ( .A(n20639), .ZN(n20640) );
  NAND2_X1 U23668 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20640), .ZN(
        n20645) );
  OAI21_X1 U23669 ( .B1(n21091), .B2(n20842), .A(n20645), .ZN(n20644) );
  NAND2_X1 U23670 ( .A1(n20782), .A2(n20640), .ZN(n20678) );
  OAI211_X1 U23671 ( .C1(n20681), .C2(n21106), .A(n20647), .B(n20941), .ZN(
        n20642) );
  INV_X1 U23672 ( .A(n20642), .ZN(n20643) );
  INV_X1 U23673 ( .A(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n20650) );
  OAI21_X1 U23674 ( .B1(n20645), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n20945), 
        .ZN(n20646) );
  AOI22_X1 U23675 ( .A1(n20665), .A2(n20950), .B1(n20681), .B2(n20949), .ZN(
        n20649) );
  AOI22_X1 U23676 ( .A1(n20662), .A2(n20952), .B1(n20666), .B2(n20951), .ZN(
        n20648) );
  OAI211_X1 U23677 ( .C1(n20655), .C2(n20650), .A(n20649), .B(n20648), .ZN(
        P2_U3104) );
  AOI22_X1 U23678 ( .A1(n20665), .A2(n20958), .B1(n20681), .B2(n20957), .ZN(
        n20652) );
  AOI22_X1 U23679 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20667), .B1(
        n20662), .B2(n20848), .ZN(n20651) );
  OAI211_X1 U23680 ( .C1(n20899), .C2(n20706), .A(n20652), .B(n20651), .ZN(
        P2_U3105) );
  INV_X1 U23681 ( .A(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n22025) );
  AOI22_X1 U23682 ( .A1(n20665), .A2(n20965), .B1(n20681), .B2(n20964), .ZN(
        n20654) );
  AOI22_X1 U23683 ( .A1(n20662), .A2(n20851), .B1(n20666), .B2(n20966), .ZN(
        n20653) );
  OAI211_X1 U23684 ( .C1(n20655), .C2(n22025), .A(n20654), .B(n20653), .ZN(
        P2_U3106) );
  AOI22_X1 U23685 ( .A1(n20665), .A2(n20971), .B1(n20681), .B2(n20970), .ZN(
        n20657) );
  AOI22_X1 U23686 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20667), .B1(
        n20666), .B2(n20972), .ZN(n20656) );
  OAI211_X1 U23687 ( .C1(n20975), .C2(n20670), .A(n20657), .B(n20656), .ZN(
        P2_U3107) );
  AOI22_X1 U23688 ( .A1(n20665), .A2(n21920), .B1(n20681), .B2(n21919), .ZN(
        n20659) );
  AOI22_X1 U23689 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20667), .B1(
        n20662), .B2(n20857), .ZN(n20658) );
  OAI211_X1 U23690 ( .C1(n20914), .C2(n20706), .A(n20659), .B(n20658), .ZN(
        P2_U3108) );
  AOI22_X1 U23691 ( .A1(n20665), .A2(n20979), .B1(n20681), .B2(n20978), .ZN(
        n20661) );
  AOI22_X1 U23692 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20667), .B1(
        n20666), .B2(n20980), .ZN(n20660) );
  OAI211_X1 U23693 ( .C1(n20983), .C2(n20670), .A(n20661), .B(n20660), .ZN(
        P2_U3109) );
  AOI22_X1 U23694 ( .A1(n20665), .A2(n20985), .B1(n20681), .B2(n20984), .ZN(
        n20664) );
  AOI22_X1 U23695 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20667), .B1(
        n20662), .B2(n20863), .ZN(n20663) );
  OAI211_X1 U23696 ( .C1(n20921), .C2(n20706), .A(n20664), .B(n20663), .ZN(
        P2_U3110) );
  AOI22_X1 U23697 ( .A1(n20665), .A2(n20992), .B1(n20681), .B2(n20990), .ZN(
        n20669) );
  AOI22_X1 U23698 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20667), .B1(
        n20666), .B2(n20994), .ZN(n20668) );
  OAI211_X1 U23699 ( .C1(n21000), .C2(n20670), .A(n20669), .B(n20668), .ZN(
        P2_U3111) );
  NAND2_X1 U23700 ( .A1(n22183), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20781) );
  NOR2_X1 U23701 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20781), .ZN(
        n20717) );
  AND2_X1 U23702 ( .A1(n20717), .A2(n21114), .ZN(n20682) );
  INV_X1 U23703 ( .A(n20682), .ZN(n20705) );
  OAI22_X1 U23704 ( .A1(n20706), .A2(n20877), .B1(n20705), .B2(n20876), .ZN(
        n20674) );
  INV_X1 U23705 ( .A(n20674), .ZN(n20686) );
  AOI21_X1 U23706 ( .B1(n20743), .B2(n20706), .A(n20842), .ZN(n20675) );
  NOR2_X1 U23707 ( .A1(n20675), .A2(n20883), .ZN(n20680) );
  AOI21_X1 U23708 ( .B1(n20676), .B2(n21106), .A(n20880), .ZN(n20677) );
  AOI21_X1 U23709 ( .B1(n20680), .B2(n20678), .A(n20677), .ZN(n20679) );
  OAI21_X1 U23710 ( .B1(n20682), .B2(n20681), .A(n20680), .ZN(n20684) );
  OAI21_X1 U23711 ( .B1(n20676), .B2(n20682), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20683) );
  AOI22_X1 U23712 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20709), .B1(
        n20950), .B2(n20708), .ZN(n20685) );
  OAI211_X1 U23713 ( .C1(n20894), .C2(n20743), .A(n20686), .B(n20685), .ZN(
        P2_U3112) );
  OAI22_X1 U23714 ( .A1(n20706), .A2(n20963), .B1(n20705), .B2(n20895), .ZN(
        n20687) );
  INV_X1 U23715 ( .A(n20687), .ZN(n20689) );
  AOI22_X1 U23716 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20709), .B1(
        n20958), .B2(n20708), .ZN(n20688) );
  OAI211_X1 U23717 ( .C1(n20899), .C2(n20743), .A(n20689), .B(n20688), .ZN(
        P2_U3113) );
  OAI22_X1 U23718 ( .A1(n20706), .A2(n20969), .B1(n20705), .B2(n20900), .ZN(
        n20690) );
  INV_X1 U23719 ( .A(n20690), .ZN(n20692) );
  AOI22_X1 U23720 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20709), .B1(
        n20965), .B2(n20708), .ZN(n20691) );
  OAI211_X1 U23721 ( .C1(n20901), .C2(n20743), .A(n20692), .B(n20691), .ZN(
        P2_U3114) );
  OAI22_X1 U23722 ( .A1(n20706), .A2(n20975), .B1(n20705), .B2(n20905), .ZN(
        n20693) );
  INV_X1 U23723 ( .A(n20693), .ZN(n20695) );
  AOI22_X1 U23724 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20709), .B1(
        n20971), .B2(n20708), .ZN(n20694) );
  OAI211_X1 U23725 ( .C1(n20906), .C2(n20743), .A(n20695), .B(n20694), .ZN(
        P2_U3115) );
  OAI22_X1 U23726 ( .A1(n20706), .A2(n21928), .B1(n20705), .B2(n20910), .ZN(
        n20696) );
  INV_X1 U23727 ( .A(n20696), .ZN(n20698) );
  AOI22_X1 U23728 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20709), .B1(
        n21920), .B2(n20708), .ZN(n20697) );
  OAI211_X1 U23729 ( .C1(n20914), .C2(n20743), .A(n20698), .B(n20697), .ZN(
        P2_U3116) );
  OAI22_X1 U23730 ( .A1(n20706), .A2(n20983), .B1(n20705), .B2(n20915), .ZN(
        n20699) );
  INV_X1 U23731 ( .A(n20699), .ZN(n20701) );
  AOI22_X1 U23732 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20709), .B1(
        n20979), .B2(n20708), .ZN(n20700) );
  OAI211_X1 U23733 ( .C1(n20916), .C2(n20743), .A(n20701), .B(n20700), .ZN(
        P2_U3117) );
  OAI22_X1 U23734 ( .A1(n20706), .A2(n20989), .B1(n20705), .B2(n20920), .ZN(
        n20702) );
  INV_X1 U23735 ( .A(n20702), .ZN(n20704) );
  AOI22_X1 U23736 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20709), .B1(
        n20985), .B2(n20708), .ZN(n20703) );
  OAI211_X1 U23737 ( .C1(n20921), .C2(n20743), .A(n20704), .B(n20703), .ZN(
        P2_U3118) );
  OAI22_X1 U23738 ( .A1(n20706), .A2(n21000), .B1(n20705), .B2(n20926), .ZN(
        n20707) );
  INV_X1 U23739 ( .A(n20707), .ZN(n20711) );
  AOI22_X1 U23740 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20709), .B1(
        n20992), .B2(n20708), .ZN(n20710) );
  OAI211_X1 U23741 ( .C1(n20927), .C2(n20743), .A(n20711), .B(n20710), .ZN(
        P2_U3119) );
  NOR2_X1 U23742 ( .A1(n20838), .A2(n20781), .ZN(n20752) );
  INV_X1 U23743 ( .A(n20752), .ZN(n20742) );
  OAI22_X1 U23744 ( .A1(n20743), .A2(n20877), .B1(n20742), .B2(n20876), .ZN(
        n20712) );
  INV_X1 U23745 ( .A(n20712), .ZN(n20723) );
  INV_X1 U23746 ( .A(n20713), .ZN(n20714) );
  OAI21_X1 U23747 ( .B1(n20714), .B2(n20842), .A(n20880), .ZN(n20721) );
  OAI21_X1 U23748 ( .B1(n20718), .B2(n20945), .A(n21106), .ZN(n20715) );
  AOI21_X1 U23749 ( .B1(n20715), .B2(n20742), .A(n20811), .ZN(n20716) );
  INV_X1 U23750 ( .A(n20717), .ZN(n20720) );
  OAI21_X1 U23751 ( .B1(n20718), .B2(n20752), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20719) );
  AOI22_X1 U23752 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20746), .B1(
        n20950), .B2(n20745), .ZN(n20722) );
  OAI211_X1 U23753 ( .C1(n20894), .C2(n20758), .A(n20723), .B(n20722), .ZN(
        P2_U3120) );
  OAI22_X1 U23754 ( .A1(n20758), .A2(n20899), .B1(n20742), .B2(n20895), .ZN(
        n20724) );
  INV_X1 U23755 ( .A(n20724), .ZN(n20726) );
  AOI22_X1 U23756 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20746), .B1(
        n20958), .B2(n20745), .ZN(n20725) );
  OAI211_X1 U23757 ( .C1(n20963), .C2(n20743), .A(n20726), .B(n20725), .ZN(
        P2_U3121) );
  OAI22_X1 U23758 ( .A1(n20758), .A2(n20901), .B1(n20742), .B2(n20900), .ZN(
        n20727) );
  INV_X1 U23759 ( .A(n20727), .ZN(n20729) );
  AOI22_X1 U23760 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20746), .B1(
        n20965), .B2(n20745), .ZN(n20728) );
  OAI211_X1 U23761 ( .C1(n20969), .C2(n20743), .A(n20729), .B(n20728), .ZN(
        P2_U3122) );
  OAI22_X1 U23762 ( .A1(n20743), .A2(n20975), .B1(n20742), .B2(n20905), .ZN(
        n20730) );
  INV_X1 U23763 ( .A(n20730), .ZN(n20732) );
  AOI22_X1 U23764 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20746), .B1(
        n20971), .B2(n20745), .ZN(n20731) );
  OAI211_X1 U23765 ( .C1(n20906), .C2(n20758), .A(n20732), .B(n20731), .ZN(
        P2_U3123) );
  OAI22_X1 U23766 ( .A1(n20743), .A2(n21928), .B1(n20742), .B2(n20910), .ZN(
        n20733) );
  INV_X1 U23767 ( .A(n20733), .ZN(n20735) );
  AOI22_X1 U23768 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20746), .B1(
        n21920), .B2(n20745), .ZN(n20734) );
  OAI211_X1 U23769 ( .C1(n20914), .C2(n20758), .A(n20735), .B(n20734), .ZN(
        P2_U3124) );
  OAI22_X1 U23770 ( .A1(n20758), .A2(n20916), .B1(n20742), .B2(n20915), .ZN(
        n20736) );
  INV_X1 U23771 ( .A(n20736), .ZN(n20738) );
  AOI22_X1 U23772 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20746), .B1(
        n20979), .B2(n20745), .ZN(n20737) );
  OAI211_X1 U23773 ( .C1(n20983), .C2(n20743), .A(n20738), .B(n20737), .ZN(
        P2_U3125) );
  OAI22_X1 U23774 ( .A1(n20758), .A2(n20921), .B1(n20742), .B2(n20920), .ZN(
        n20739) );
  INV_X1 U23775 ( .A(n20739), .ZN(n20741) );
  AOI22_X1 U23776 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20746), .B1(
        n20985), .B2(n20745), .ZN(n20740) );
  OAI211_X1 U23777 ( .C1(n20989), .C2(n20743), .A(n20741), .B(n20740), .ZN(
        P2_U3126) );
  OAI22_X1 U23778 ( .A1(n20743), .A2(n21000), .B1(n20742), .B2(n20926), .ZN(
        n20744) );
  INV_X1 U23779 ( .A(n20744), .ZN(n20748) );
  AOI22_X1 U23780 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20746), .B1(
        n20992), .B2(n20745), .ZN(n20747) );
  OAI211_X1 U23781 ( .C1(n20927), .C2(n20758), .A(n20748), .B(n20747), .ZN(
        P2_U3127) );
  INV_X1 U23782 ( .A(n20754), .ZN(n20749) );
  NOR2_X1 U23783 ( .A1(n20874), .A2(n20781), .ZN(n20773) );
  OAI21_X1 U23784 ( .B1(n20749), .B2(n20773), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20750) );
  AOI22_X1 U23785 ( .A1(n20774), .A2(n20950), .B1(n20949), .B2(n20773), .ZN(
        n20760) );
  AOI21_X1 U23786 ( .B1(n20758), .B2(n21927), .A(n20842), .ZN(n20753) );
  NOR2_X1 U23787 ( .A1(n20753), .A2(n20752), .ZN(n20755) );
  MUX2_X1 U23788 ( .A(n20755), .B(n20754), .S(P2_STATE2_REG_2__SCAN_IN), .Z(
        n20756) );
  NOR2_X1 U23789 ( .A1(n20756), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20757) );
  AOI22_X1 U23790 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20776), .B1(
        n20775), .B2(n20952), .ZN(n20759) );
  OAI211_X1 U23791 ( .C1(n20894), .C2(n21927), .A(n20760), .B(n20759), .ZN(
        P2_U3128) );
  AOI22_X1 U23792 ( .A1(n20774), .A2(n20958), .B1(n20957), .B2(n20773), .ZN(
        n20762) );
  AOI22_X1 U23793 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20776), .B1(
        n20775), .B2(n20848), .ZN(n20761) );
  OAI211_X1 U23794 ( .C1(n20899), .C2(n21927), .A(n20762), .B(n20761), .ZN(
        P2_U3129) );
  AOI22_X1 U23795 ( .A1(n20774), .A2(n20965), .B1(n20964), .B2(n20773), .ZN(
        n20764) );
  AOI22_X1 U23796 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20776), .B1(
        n20775), .B2(n20851), .ZN(n20763) );
  OAI211_X1 U23797 ( .C1(n20901), .C2(n21927), .A(n20764), .B(n20763), .ZN(
        P2_U3130) );
  AOI22_X1 U23798 ( .A1(n20774), .A2(n20971), .B1(n20970), .B2(n20773), .ZN(
        n20766) );
  AOI22_X1 U23799 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20776), .B1(
        n20775), .B2(n20854), .ZN(n20765) );
  OAI211_X1 U23800 ( .C1(n20906), .C2(n21927), .A(n20766), .B(n20765), .ZN(
        P2_U3131) );
  AOI22_X1 U23801 ( .A1(n20774), .A2(n21920), .B1(n21919), .B2(n20773), .ZN(
        n20768) );
  AOI22_X1 U23802 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20776), .B1(
        n20775), .B2(n20857), .ZN(n20767) );
  OAI211_X1 U23803 ( .C1(n20914), .C2(n21927), .A(n20768), .B(n20767), .ZN(
        P2_U3132) );
  AOI22_X1 U23804 ( .A1(n20774), .A2(n20979), .B1(n20978), .B2(n20773), .ZN(
        n20770) );
  AOI22_X1 U23805 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20776), .B1(
        n20775), .B2(n20860), .ZN(n20769) );
  OAI211_X1 U23806 ( .C1(n20916), .C2(n21927), .A(n20770), .B(n20769), .ZN(
        P2_U3133) );
  AOI22_X1 U23807 ( .A1(n20774), .A2(n20985), .B1(n20984), .B2(n20773), .ZN(
        n20772) );
  AOI22_X1 U23808 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20776), .B1(
        n20775), .B2(n20863), .ZN(n20771) );
  OAI211_X1 U23809 ( .C1(n20921), .C2(n21927), .A(n20772), .B(n20771), .ZN(
        P2_U3134) );
  AOI22_X1 U23810 ( .A1(n20774), .A2(n20992), .B1(n20990), .B2(n20773), .ZN(
        n20778) );
  AOI22_X1 U23811 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20776), .B1(
        n20775), .B2(n20868), .ZN(n20777) );
  OAI211_X1 U23812 ( .C1(n20927), .C2(n21927), .A(n20778), .B(n20777), .ZN(
        P2_U3135) );
  INV_X1 U23813 ( .A(n20781), .ZN(n20785) );
  NAND2_X1 U23814 ( .A1(n20782), .A2(n20785), .ZN(n20788) );
  NAND2_X1 U23815 ( .A1(n20788), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n20783) );
  NAND2_X1 U23816 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20785), .ZN(
        n20787) );
  OAI21_X1 U23817 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n20787), .A(n20945), 
        .ZN(n20786) );
  INV_X1 U23818 ( .A(n20788), .ZN(n21918) );
  AOI22_X1 U23819 ( .A1(n21921), .A2(n20950), .B1(n20949), .B2(n21918), .ZN(
        n20793) );
  OAI21_X1 U23820 ( .B1(n21092), .B2(n21087), .A(n20787), .ZN(n20791) );
  NAND2_X1 U23821 ( .A1(n20788), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20789) );
  NAND4_X1 U23822 ( .A1(n20791), .A2(n20941), .A3(n20790), .A4(n20789), .ZN(
        n21924) );
  INV_X1 U23823 ( .A(n21927), .ZN(n20800) );
  AOI22_X1 U23824 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n21924), .B1(
        n20800), .B2(n20952), .ZN(n20792) );
  OAI211_X1 U23825 ( .C1(n20894), .C2(n20835), .A(n20793), .B(n20792), .ZN(
        P2_U3136) );
  AOI22_X1 U23826 ( .A1(n21921), .A2(n20958), .B1(n20957), .B2(n21918), .ZN(
        n20795) );
  AOI22_X1 U23827 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n21924), .B1(
        n20800), .B2(n20848), .ZN(n20794) );
  OAI211_X1 U23828 ( .C1(n20899), .C2(n20835), .A(n20795), .B(n20794), .ZN(
        P2_U3137) );
  AOI22_X1 U23829 ( .A1(n21921), .A2(n20965), .B1(n20964), .B2(n21918), .ZN(
        n20797) );
  AOI22_X1 U23830 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n21924), .B1(
        n20800), .B2(n20851), .ZN(n20796) );
  OAI211_X1 U23831 ( .C1(n20901), .C2(n20835), .A(n20797), .B(n20796), .ZN(
        P2_U3138) );
  AOI22_X1 U23832 ( .A1(n21921), .A2(n20971), .B1(n20970), .B2(n21918), .ZN(
        n20799) );
  AOI22_X1 U23833 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n21924), .B1(
        n20800), .B2(n20854), .ZN(n20798) );
  OAI211_X1 U23834 ( .C1(n20906), .C2(n20835), .A(n20799), .B(n20798), .ZN(
        P2_U3139) );
  AOI22_X1 U23835 ( .A1(n21921), .A2(n20979), .B1(n20978), .B2(n21918), .ZN(
        n20802) );
  AOI22_X1 U23836 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n21924), .B1(
        n20800), .B2(n20860), .ZN(n20801) );
  OAI211_X1 U23837 ( .C1(n20916), .C2(n20835), .A(n20802), .B(n20801), .ZN(
        P2_U3141) );
  AOI22_X1 U23838 ( .A1(n21921), .A2(n20985), .B1(n20984), .B2(n21918), .ZN(
        n20804) );
  INV_X1 U23839 ( .A(n20835), .ZN(n21923) );
  AOI22_X1 U23840 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n21924), .B1(
        n21923), .B2(n20986), .ZN(n20803) );
  OAI211_X1 U23841 ( .C1(n20989), .C2(n21927), .A(n20804), .B(n20803), .ZN(
        P2_U3142) );
  AOI22_X1 U23842 ( .A1(n21921), .A2(n20992), .B1(n20990), .B2(n21918), .ZN(
        n20806) );
  AOI22_X1 U23843 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n21924), .B1(
        n21923), .B2(n20994), .ZN(n20805) );
  OAI211_X1 U23844 ( .C1(n21000), .C2(n21927), .A(n20806), .B(n20805), .ZN(
        P2_U3143) );
  INV_X1 U23845 ( .A(n20936), .ZN(n20875) );
  NOR3_X2 U23846 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n20875), .ZN(n20830) );
  NOR3_X1 U23847 ( .A1(n11052), .A2(n20830), .A3(n20945), .ZN(n20812) );
  NAND3_X1 U23848 ( .A1(n20808), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        n20807), .ZN(n20813) );
  INV_X1 U23849 ( .A(n20813), .ZN(n20809) );
  AOI21_X1 U23850 ( .B1(n20809), .B2(n21106), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20810) );
  AOI22_X1 U23851 ( .A1(n20831), .A2(n20950), .B1(n20949), .B2(n20830), .ZN(
        n20817) );
  OAI21_X1 U23852 ( .B1(n20869), .B2(n21923), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n20814) );
  AOI211_X1 U23853 ( .C1(n20814), .C2(n20813), .A(n20812), .B(n20811), .ZN(
        n20815) );
  AOI22_X1 U23854 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20832), .B1(
        n20869), .B2(n20951), .ZN(n20816) );
  OAI211_X1 U23855 ( .C1(n20877), .C2(n20835), .A(n20817), .B(n20816), .ZN(
        P2_U3144) );
  AOI22_X1 U23856 ( .A1(n20831), .A2(n20958), .B1(n20957), .B2(n20830), .ZN(
        n20819) );
  AOI22_X1 U23857 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20832), .B1(
        n20869), .B2(n20960), .ZN(n20818) );
  OAI211_X1 U23858 ( .C1(n20963), .C2(n20835), .A(n20819), .B(n20818), .ZN(
        P2_U3145) );
  AOI22_X1 U23859 ( .A1(n20831), .A2(n20965), .B1(n20964), .B2(n20830), .ZN(
        n20821) );
  AOI22_X1 U23860 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20832), .B1(
        n20869), .B2(n20966), .ZN(n20820) );
  OAI211_X1 U23861 ( .C1(n20969), .C2(n20835), .A(n20821), .B(n20820), .ZN(
        P2_U3146) );
  AOI22_X1 U23862 ( .A1(n20831), .A2(n20971), .B1(n20970), .B2(n20830), .ZN(
        n20823) );
  AOI22_X1 U23863 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20832), .B1(
        n20869), .B2(n20972), .ZN(n20822) );
  OAI211_X1 U23864 ( .C1(n20975), .C2(n20835), .A(n20823), .B(n20822), .ZN(
        P2_U3147) );
  AOI22_X1 U23865 ( .A1(n20831), .A2(n21920), .B1(n21919), .B2(n20830), .ZN(
        n20825) );
  AOI22_X1 U23866 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20832), .B1(
        n20869), .B2(n21922), .ZN(n20824) );
  OAI211_X1 U23867 ( .C1(n21928), .C2(n20835), .A(n20825), .B(n20824), .ZN(
        P2_U3148) );
  AOI22_X1 U23868 ( .A1(n20831), .A2(n20979), .B1(n20978), .B2(n20830), .ZN(
        n20827) );
  AOI22_X1 U23869 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20832), .B1(
        n20869), .B2(n20980), .ZN(n20826) );
  OAI211_X1 U23870 ( .C1(n20983), .C2(n20835), .A(n20827), .B(n20826), .ZN(
        P2_U3149) );
  AOI22_X1 U23871 ( .A1(n20831), .A2(n20985), .B1(n20984), .B2(n20830), .ZN(
        n20829) );
  AOI22_X1 U23872 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20832), .B1(
        n20869), .B2(n20986), .ZN(n20828) );
  OAI211_X1 U23873 ( .C1(n20989), .C2(n20835), .A(n20829), .B(n20828), .ZN(
        P2_U3150) );
  AOI22_X1 U23874 ( .A1(n20831), .A2(n20992), .B1(n20990), .B2(n20830), .ZN(
        n20834) );
  AOI22_X1 U23875 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20832), .B1(
        n20869), .B2(n20994), .ZN(n20833) );
  OAI211_X1 U23876 ( .C1(n21000), .C2(n20835), .A(n20834), .B(n20833), .ZN(
        P2_U3151) );
  NAND2_X1 U23877 ( .A1(n20837), .A2(n20936), .ZN(n20841) );
  NOR2_X1 U23878 ( .A1(n20838), .A2(n20875), .ZN(n20866) );
  OAI21_X1 U23879 ( .B1(n20839), .B2(n20866), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20840) );
  OAI21_X1 U23880 ( .B1(n20841), .B2(n20883), .A(n20840), .ZN(n20867) );
  AOI22_X1 U23881 ( .A1(n20867), .A2(n20950), .B1(n20949), .B2(n20866), .ZN(
        n20847) );
  AOI21_X1 U23882 ( .B1(n11087), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n20845) );
  OAI21_X1 U23883 ( .B1(n20843), .B2(n20842), .A(n20841), .ZN(n20844) );
  OAI211_X1 U23884 ( .C1(n20866), .C2(n20845), .A(n20844), .B(n20941), .ZN(
        n20870) );
  AOI22_X1 U23885 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20870), .B1(
        n20869), .B2(n20952), .ZN(n20846) );
  OAI211_X1 U23886 ( .C1(n20894), .C2(n20933), .A(n20847), .B(n20846), .ZN(
        P2_U3152) );
  AOI22_X1 U23887 ( .A1(n20867), .A2(n20958), .B1(n20957), .B2(n20866), .ZN(
        n20850) );
  AOI22_X1 U23888 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20870), .B1(
        n20869), .B2(n20848), .ZN(n20849) );
  OAI211_X1 U23889 ( .C1(n20899), .C2(n20933), .A(n20850), .B(n20849), .ZN(
        P2_U3153) );
  AOI22_X1 U23890 ( .A1(n20867), .A2(n20965), .B1(n20964), .B2(n20866), .ZN(
        n20853) );
  AOI22_X1 U23891 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20870), .B1(
        n20869), .B2(n20851), .ZN(n20852) );
  OAI211_X1 U23892 ( .C1(n20901), .C2(n20933), .A(n20853), .B(n20852), .ZN(
        P2_U3154) );
  AOI22_X1 U23893 ( .A1(n20867), .A2(n20971), .B1(n20970), .B2(n20866), .ZN(
        n20856) );
  AOI22_X1 U23894 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20870), .B1(
        n20869), .B2(n20854), .ZN(n20855) );
  OAI211_X1 U23895 ( .C1(n20906), .C2(n20933), .A(n20856), .B(n20855), .ZN(
        P2_U3155) );
  AOI22_X1 U23896 ( .A1(n20867), .A2(n21920), .B1(n21919), .B2(n20866), .ZN(
        n20859) );
  AOI22_X1 U23897 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20870), .B1(
        n20869), .B2(n20857), .ZN(n20858) );
  OAI211_X1 U23898 ( .C1(n20914), .C2(n20933), .A(n20859), .B(n20858), .ZN(
        P2_U3156) );
  AOI22_X1 U23899 ( .A1(n20867), .A2(n20979), .B1(n20978), .B2(n20866), .ZN(
        n20862) );
  AOI22_X1 U23900 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20870), .B1(
        n20869), .B2(n20860), .ZN(n20861) );
  OAI211_X1 U23901 ( .C1(n20916), .C2(n20933), .A(n20862), .B(n20861), .ZN(
        P2_U3157) );
  AOI22_X1 U23902 ( .A1(n20867), .A2(n20985), .B1(n20984), .B2(n20866), .ZN(
        n20865) );
  AOI22_X1 U23903 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20870), .B1(
        n20869), .B2(n20863), .ZN(n20864) );
  OAI211_X1 U23904 ( .C1(n20921), .C2(n20933), .A(n20865), .B(n20864), .ZN(
        P2_U3158) );
  AOI22_X1 U23905 ( .A1(n20867), .A2(n20992), .B1(n20990), .B2(n20866), .ZN(
        n20872) );
  AOI22_X1 U23906 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20870), .B1(
        n20869), .B2(n20868), .ZN(n20871) );
  OAI211_X1 U23907 ( .C1(n20927), .C2(n20933), .A(n20872), .B(n20871), .ZN(
        P2_U3159) );
  NOR2_X1 U23908 ( .A1(n20875), .A2(n20874), .ZN(n20887) );
  OAI22_X1 U23909 ( .A1(n20933), .A2(n20877), .B1(n20876), .B2(n20925), .ZN(
        n20878) );
  INV_X1 U23910 ( .A(n20878), .ZN(n20893) );
  INV_X1 U23911 ( .A(n20933), .ZN(n20879) );
  INV_X1 U23912 ( .A(n20999), .ZN(n20953) );
  OAI21_X1 U23913 ( .B1(n20879), .B2(n20953), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n20881) );
  NAND2_X1 U23914 ( .A1(n20881), .A2(n20880), .ZN(n20891) );
  AND2_X1 U23915 ( .A1(n20882), .A2(n20936), .ZN(n20886) );
  OAI211_X1 U23916 ( .C1(n20884), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n20883), 
        .B(n20925), .ZN(n20885) );
  OAI211_X1 U23917 ( .C1(n20891), .C2(n20886), .A(n20941), .B(n20885), .ZN(
        n20930) );
  INV_X1 U23918 ( .A(n20886), .ZN(n20890) );
  OAI21_X1 U23919 ( .B1(n20888), .B2(n20887), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20889) );
  AOI22_X1 U23920 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20930), .B1(
        n20950), .B2(n20929), .ZN(n20892) );
  OAI211_X1 U23921 ( .C1(n20894), .C2(n20999), .A(n20893), .B(n20892), .ZN(
        P2_U3160) );
  OAI22_X1 U23922 ( .A1(n20933), .A2(n20963), .B1(n20895), .B2(n20925), .ZN(
        n20896) );
  INV_X1 U23923 ( .A(n20896), .ZN(n20898) );
  AOI22_X1 U23924 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20930), .B1(
        n20958), .B2(n20929), .ZN(n20897) );
  OAI211_X1 U23925 ( .C1(n20899), .C2(n20999), .A(n20898), .B(n20897), .ZN(
        P2_U3161) );
  OAI22_X1 U23926 ( .A1(n20999), .A2(n20901), .B1(n20900), .B2(n20925), .ZN(
        n20902) );
  INV_X1 U23927 ( .A(n20902), .ZN(n20904) );
  AOI22_X1 U23928 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20930), .B1(
        n20965), .B2(n20929), .ZN(n20903) );
  OAI211_X1 U23929 ( .C1(n20969), .C2(n20933), .A(n20904), .B(n20903), .ZN(
        P2_U3162) );
  OAI22_X1 U23930 ( .A1(n20999), .A2(n20906), .B1(n20905), .B2(n20925), .ZN(
        n20907) );
  INV_X1 U23931 ( .A(n20907), .ZN(n20909) );
  AOI22_X1 U23932 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20930), .B1(
        n20971), .B2(n20929), .ZN(n20908) );
  OAI211_X1 U23933 ( .C1(n20975), .C2(n20933), .A(n20909), .B(n20908), .ZN(
        P2_U3163) );
  OAI22_X1 U23934 ( .A1(n20933), .A2(n21928), .B1(n20910), .B2(n20925), .ZN(
        n20911) );
  INV_X1 U23935 ( .A(n20911), .ZN(n20913) );
  AOI22_X1 U23936 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20930), .B1(
        n21920), .B2(n20929), .ZN(n20912) );
  OAI211_X1 U23937 ( .C1(n20914), .C2(n20999), .A(n20913), .B(n20912), .ZN(
        P2_U3164) );
  OAI22_X1 U23938 ( .A1(n20999), .A2(n20916), .B1(n20915), .B2(n20925), .ZN(
        n20917) );
  INV_X1 U23939 ( .A(n20917), .ZN(n20919) );
  AOI22_X1 U23940 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20930), .B1(
        n20979), .B2(n20929), .ZN(n20918) );
  OAI211_X1 U23941 ( .C1(n20983), .C2(n20933), .A(n20919), .B(n20918), .ZN(
        P2_U3165) );
  OAI22_X1 U23942 ( .A1(n20999), .A2(n20921), .B1(n20920), .B2(n20925), .ZN(
        n20922) );
  INV_X1 U23943 ( .A(n20922), .ZN(n20924) );
  AOI22_X1 U23944 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20930), .B1(
        n20985), .B2(n20929), .ZN(n20923) );
  OAI211_X1 U23945 ( .C1(n20989), .C2(n20933), .A(n20924), .B(n20923), .ZN(
        P2_U3166) );
  OAI22_X1 U23946 ( .A1(n20999), .A2(n20927), .B1(n20926), .B2(n20925), .ZN(
        n20928) );
  INV_X1 U23947 ( .A(n20928), .ZN(n20932) );
  AOI22_X1 U23948 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20930), .B1(
        n20992), .B2(n20929), .ZN(n20931) );
  OAI211_X1 U23949 ( .C1(n21000), .C2(n20933), .A(n20932), .B(n20931), .ZN(
        P2_U3167) );
  INV_X1 U23950 ( .A(n21087), .ZN(n20934) );
  NAND2_X1 U23951 ( .A1(n20935), .A2(n20934), .ZN(n20937) );
  NAND2_X1 U23952 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20936), .ZN(
        n20946) );
  NAND2_X1 U23953 ( .A1(n20937), .A2(n20946), .ZN(n20944) );
  NAND2_X1 U23954 ( .A1(n20938), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n20939) );
  OAI211_X1 U23955 ( .C1(n20991), .C2(n21106), .A(n20948), .B(n20941), .ZN(
        n20942) );
  INV_X1 U23956 ( .A(n20942), .ZN(n20943) );
  INV_X1 U23957 ( .A(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n20956) );
  OAI21_X1 U23958 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n20946), .A(n20945), 
        .ZN(n20947) );
  AND2_X1 U23959 ( .A1(n20948), .A2(n20947), .ZN(n20993) );
  AOI22_X1 U23960 ( .A1(n20993), .A2(n20950), .B1(n20991), .B2(n20949), .ZN(
        n20955) );
  AOI22_X1 U23961 ( .A1(n20953), .A2(n20952), .B1(n20995), .B2(n20951), .ZN(
        n20954) );
  OAI211_X1 U23962 ( .C1(n20959), .C2(n20956), .A(n20955), .B(n20954), .ZN(
        P2_U3168) );
  AOI22_X1 U23963 ( .A1(n20993), .A2(n20958), .B1(n20991), .B2(n20957), .ZN(
        n20962) );
  AOI22_X1 U23964 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20996), .B1(
        n20995), .B2(n20960), .ZN(n20961) );
  OAI211_X1 U23965 ( .C1(n20963), .C2(n20999), .A(n20962), .B(n20961), .ZN(
        P2_U3169) );
  AOI22_X1 U23966 ( .A1(n20993), .A2(n20965), .B1(n20991), .B2(n20964), .ZN(
        n20968) );
  AOI22_X1 U23967 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20996), .B1(
        n20995), .B2(n20966), .ZN(n20967) );
  OAI211_X1 U23968 ( .C1(n20969), .C2(n20999), .A(n20968), .B(n20967), .ZN(
        P2_U3170) );
  AOI22_X1 U23969 ( .A1(n20993), .A2(n20971), .B1(n20991), .B2(n20970), .ZN(
        n20974) );
  AOI22_X1 U23970 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20996), .B1(
        n20995), .B2(n20972), .ZN(n20973) );
  OAI211_X1 U23971 ( .C1(n20975), .C2(n20999), .A(n20974), .B(n20973), .ZN(
        P2_U3171) );
  AOI22_X1 U23972 ( .A1(n20993), .A2(n21920), .B1(n20991), .B2(n21919), .ZN(
        n20977) );
  AOI22_X1 U23973 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20996), .B1(
        n20995), .B2(n21922), .ZN(n20976) );
  OAI211_X1 U23974 ( .C1(n21928), .C2(n20999), .A(n20977), .B(n20976), .ZN(
        P2_U3172) );
  AOI22_X1 U23975 ( .A1(n20993), .A2(n20979), .B1(n20991), .B2(n20978), .ZN(
        n20982) );
  AOI22_X1 U23976 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20996), .B1(
        n20995), .B2(n20980), .ZN(n20981) );
  OAI211_X1 U23977 ( .C1(n20983), .C2(n20999), .A(n20982), .B(n20981), .ZN(
        P2_U3173) );
  AOI22_X1 U23978 ( .A1(n20993), .A2(n20985), .B1(n20991), .B2(n20984), .ZN(
        n20988) );
  AOI22_X1 U23979 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20996), .B1(
        n20995), .B2(n20986), .ZN(n20987) );
  OAI211_X1 U23980 ( .C1(n20989), .C2(n20999), .A(n20988), .B(n20987), .ZN(
        P2_U3174) );
  AOI22_X1 U23981 ( .A1(n20993), .A2(n20992), .B1(n20991), .B2(n20990), .ZN(
        n20998) );
  AOI22_X1 U23982 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20996), .B1(
        n20995), .B2(n20994), .ZN(n20997) );
  OAI211_X1 U23983 ( .C1(n21000), .C2(n20999), .A(n20998), .B(n20997), .ZN(
        P2_U3175) );
  NOR3_X1 U23984 ( .A1(n21126), .A2(P2_STATE2_REG_3__SCAN_IN), .A3(n21132), 
        .ZN(n21001) );
  OAI21_X1 U23985 ( .B1(n10671), .B2(n21001), .A(n21002), .ZN(n21008) );
  INV_X1 U23986 ( .A(n21002), .ZN(n21005) );
  INV_X1 U23987 ( .A(n21003), .ZN(n21004) );
  OAI21_X1 U23988 ( .B1(n21005), .B2(n21004), .A(n21126), .ZN(n21007) );
  OAI221_X1 U23989 ( .B1(P2_STATE2_REG_1__SCAN_IN), .B2(n21008), .C1(n11279), 
        .C2(n21007), .A(n21006), .ZN(P2_U3177) );
  AND2_X1 U23990 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n21009), .ZN(
        P2_U3179) );
  AND2_X1 U23991 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n21009), .ZN(
        P2_U3180) );
  AND2_X1 U23992 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n21009), .ZN(
        P2_U3181) );
  AND2_X1 U23993 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n21009), .ZN(
        P2_U3182) );
  AND2_X1 U23994 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n21009), .ZN(
        P2_U3183) );
  AND2_X1 U23995 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n21009), .ZN(
        P2_U3184) );
  AND2_X1 U23996 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n21009), .ZN(
        P2_U3185) );
  AND2_X1 U23997 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n21009), .ZN(
        P2_U3186) );
  INV_X1 U23998 ( .A(P2_DATAWIDTH_REG_23__SCAN_IN), .ZN(n22081) );
  NOR2_X1 U23999 ( .A1(n22081), .A2(n21085), .ZN(P2_U3187) );
  AND2_X1 U24000 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n21009), .ZN(
        P2_U3188) );
  AND2_X1 U24001 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n21009), .ZN(
        P2_U3189) );
  AND2_X1 U24002 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n21009), .ZN(
        P2_U3190) );
  NOR2_X1 U24003 ( .A1(n22071), .A2(n21085), .ZN(P2_U3191) );
  AND2_X1 U24004 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n21009), .ZN(
        P2_U3192) );
  AND2_X1 U24005 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n21009), .ZN(
        P2_U3193) );
  AND2_X1 U24006 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n21009), .ZN(
        P2_U3194) );
  AND2_X1 U24007 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n21009), .ZN(
        P2_U3195) );
  AND2_X1 U24008 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n21009), .ZN(
        P2_U3196) );
  AND2_X1 U24009 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n21009), .ZN(
        P2_U3197) );
  AND2_X1 U24010 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n21009), .ZN(
        P2_U3198) );
  AND2_X1 U24011 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n21009), .ZN(
        P2_U3199) );
  AND2_X1 U24012 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n21009), .ZN(
        P2_U3200) );
  AND2_X1 U24013 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n21009), .ZN(P2_U3201) );
  AND2_X1 U24014 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n21009), .ZN(P2_U3202) );
  AND2_X1 U24015 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n21009), .ZN(P2_U3203) );
  AND2_X1 U24016 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n21009), .ZN(P2_U3204) );
  NOR2_X1 U24017 ( .A1(n22137), .A2(n21085), .ZN(P2_U3205) );
  AND2_X1 U24018 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n21009), .ZN(P2_U3206) );
  AND2_X1 U24019 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n21009), .ZN(P2_U3207) );
  AND2_X1 U24020 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n21009), .ZN(P2_U3208) );
  NOR3_X1 U24021 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(P2_STATE_REG_1__SCAN_IN), 
        .A3(n21010), .ZN(n21029) );
  INV_X1 U24022 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n21016) );
  NOR2_X1 U24023 ( .A1(n21011), .A2(n21016), .ZN(n21012) );
  NAND2_X1 U24024 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n21126), .ZN(n21024) );
  AOI21_X1 U24025 ( .B1(n21012), .B2(n21024), .A(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n21015) );
  AOI211_X1 U24026 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(n21020), .A(
        n21013), .B(n21140), .ZN(n21014) );
  OR3_X1 U24027 ( .A1(n21029), .A2(n21015), .A3(n21014), .ZN(P2_U3209) );
  AOI21_X1 U24028 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n21020), .A(n21030), 
        .ZN(n21022) );
  NOR3_X1 U24029 ( .A1(n21022), .A2(n21016), .A3(n21011), .ZN(n21017) );
  NOR2_X1 U24030 ( .A1(n21017), .A2(n21129), .ZN(n21018) );
  OAI211_X1 U24031 ( .C1(n21020), .C2(n21019), .A(n21018), .B(n21024), .ZN(
        P2_U3210) );
  NOR2_X1 U24032 ( .A1(n21021), .A2(n21030), .ZN(n21023) );
  AOI21_X1 U24033 ( .B1(n21126), .B2(n21023), .A(n21022), .ZN(n21028) );
  OAI22_X1 U24034 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(n21025), .B1(NA), 
        .B2(n21024), .ZN(n21026) );
  OAI211_X1 U24035 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n21026), .ZN(n21027) );
  OAI21_X1 U24036 ( .B1(n21029), .B2(n21028), .A(n21027), .ZN(P2_U3211) );
  NAND2_X2 U24037 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n21140), .ZN(n21077) );
  OAI222_X1 U24038 ( .A1(n21080), .A2(n21034), .B1(n21032), .B2(n21140), .C1(
        n21031), .C2(n21077), .ZN(P2_U3212) );
  OAI222_X1 U24039 ( .A1(n21077), .A2(n21034), .B1(n21033), .B2(n21140), .C1(
        n21035), .C2(n21080), .ZN(P2_U3213) );
  OAI222_X1 U24040 ( .A1(n21080), .A2(n21036), .B1(n22020), .B2(n21140), .C1(
        n21035), .C2(n21077), .ZN(P2_U3214) );
  OAI222_X1 U24041 ( .A1(n21080), .A2(n21038), .B1(n21037), .B2(n21140), .C1(
        n21036), .C2(n21077), .ZN(P2_U3215) );
  OAI222_X1 U24042 ( .A1(n21080), .A2(n21040), .B1(n21039), .B2(n21140), .C1(
        n21038), .C2(n21077), .ZN(P2_U3216) );
  OAI222_X1 U24043 ( .A1(n21080), .A2(n21042), .B1(n21041), .B2(n21140), .C1(
        n21040), .C2(n21077), .ZN(P2_U3217) );
  OAI222_X1 U24044 ( .A1(n21080), .A2(n21044), .B1(n21043), .B2(n21140), .C1(
        n21042), .C2(n21077), .ZN(P2_U3218) );
  OAI222_X1 U24045 ( .A1(n21080), .A2(n21046), .B1(n21045), .B2(n21140), .C1(
        n21044), .C2(n21077), .ZN(P2_U3219) );
  OAI222_X1 U24046 ( .A1(n21080), .A2(n22182), .B1(n21047), .B2(n21140), .C1(
        n21046), .C2(n21077), .ZN(P2_U3220) );
  OAI222_X1 U24047 ( .A1(n21080), .A2(n16694), .B1(n21048), .B2(n21140), .C1(
        n22182), .C2(n21077), .ZN(P2_U3221) );
  OAI222_X1 U24048 ( .A1(n21080), .A2(n21050), .B1(n21049), .B2(n21140), .C1(
        n16694), .C2(n21077), .ZN(P2_U3222) );
  OAI222_X1 U24049 ( .A1(n21080), .A2(n16144), .B1(n21051), .B2(n21140), .C1(
        n21050), .C2(n21077), .ZN(P2_U3223) );
  OAI222_X1 U24050 ( .A1(n21080), .A2(n21053), .B1(n21052), .B2(n21140), .C1(
        n16144), .C2(n21077), .ZN(P2_U3224) );
  OAI222_X1 U24051 ( .A1(n21080), .A2(n21055), .B1(n21054), .B2(n21140), .C1(
        n21053), .C2(n21077), .ZN(P2_U3225) );
  OAI222_X1 U24052 ( .A1(n21080), .A2(n21056), .B1(n22066), .B2(n21140), .C1(
        n21055), .C2(n21077), .ZN(P2_U3226) );
  OAI222_X1 U24053 ( .A1(n21080), .A2(n21058), .B1(n21057), .B2(n21140), .C1(
        n21056), .C2(n21077), .ZN(P2_U3227) );
  OAI222_X1 U24054 ( .A1(n21080), .A2(n16618), .B1(n21059), .B2(n21140), .C1(
        n21058), .C2(n21077), .ZN(P2_U3228) );
  OAI222_X1 U24055 ( .A1(n21080), .A2(n21061), .B1(n21060), .B2(n21140), .C1(
        n16618), .C2(n21077), .ZN(P2_U3229) );
  OAI222_X1 U24056 ( .A1(n21080), .A2(n16606), .B1(n21062), .B2(n21140), .C1(
        n21061), .C2(n21077), .ZN(P2_U3230) );
  OAI222_X1 U24057 ( .A1(n21080), .A2(n21064), .B1(n21063), .B2(n21140), .C1(
        n16606), .C2(n21077), .ZN(P2_U3231) );
  OAI222_X1 U24058 ( .A1(n21080), .A2(n16581), .B1(n21065), .B2(n21140), .C1(
        n21064), .C2(n21077), .ZN(P2_U3232) );
  INV_X1 U24059 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n21067) );
  OAI222_X1 U24060 ( .A1(n21080), .A2(n21067), .B1(n21066), .B2(n21140), .C1(
        n16581), .C2(n21077), .ZN(P2_U3233) );
  OAI222_X1 U24061 ( .A1(n21080), .A2(n11681), .B1(n21068), .B2(n21140), .C1(
        n21067), .C2(n21077), .ZN(P2_U3234) );
  OAI222_X1 U24062 ( .A1(n21080), .A2(n21070), .B1(n21069), .B2(n21140), .C1(
        n11681), .C2(n21077), .ZN(P2_U3235) );
  OAI222_X1 U24063 ( .A1(n21080), .A2(n21072), .B1(n21071), .B2(n21140), .C1(
        n21070), .C2(n21077), .ZN(P2_U3236) );
  OAI222_X1 U24064 ( .A1(n21080), .A2(n21074), .B1(n22117), .B2(n21140), .C1(
        n21072), .C2(n21077), .ZN(P2_U3237) );
  OAI222_X1 U24065 ( .A1(n21077), .A2(n21074), .B1(n21073), .B2(n21140), .C1(
        n16528), .C2(n21080), .ZN(P2_U3238) );
  OAI222_X1 U24066 ( .A1(n21080), .A2(n21076), .B1(n21075), .B2(n21140), .C1(
        n16528), .C2(n21077), .ZN(P2_U3239) );
  OAI222_X1 U24067 ( .A1(n21080), .A2(n21078), .B1(n22233), .B2(n21140), .C1(
        n21076), .C2(n21077), .ZN(P2_U3240) );
  OAI222_X1 U24068 ( .A1(n21080), .A2(n15932), .B1(n21079), .B2(n21140), .C1(
        n21078), .C2(n21077), .ZN(P2_U3241) );
  AOI22_X1 U24069 ( .A1(n21140), .A2(n22023), .B1(n22104), .B2(n21141), .ZN(
        P2_U3585) );
  MUX2_X1 U24070 ( .A(P2_BYTEENABLE_REG_2__SCAN_IN), .B(P2_BE_N_REG_2__SCAN_IN), .S(n21141), .Z(P2_U3586) );
  MUX2_X1 U24071 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .B(P2_BE_N_REG_1__SCAN_IN), .S(n21141), .Z(P2_U3587) );
  OAI22_X1 U24072 ( .A1(n21141), .A2(P2_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P2_BE_N_REG_0__SCAN_IN), .B2(n21140), .ZN(n21081) );
  INV_X1 U24073 ( .A(n21081), .ZN(P2_U3588) );
  OAI21_X1 U24074 ( .B1(n21085), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n21083), 
        .ZN(n21082) );
  INV_X1 U24075 ( .A(n21082), .ZN(P2_U3591) );
  OAI21_X1 U24076 ( .B1(n21085), .B2(n21084), .A(n21083), .ZN(P2_U3592) );
  OR2_X1 U24077 ( .A1(n21087), .A2(n21086), .ZN(n21088) );
  NAND2_X1 U24078 ( .A1(n21088), .A2(n21110), .ZN(n21097) );
  OAI22_X1 U24079 ( .A1(n21090), .A2(n21097), .B1(n21106), .B2(n21089), .ZN(
        n21094) );
  AOI21_X1 U24080 ( .B1(n21092), .B2(n21091), .A(n21098), .ZN(n21093) );
  OAI21_X1 U24081 ( .B1(n21094), .B2(n21093), .A(n21112), .ZN(n21095) );
  OAI21_X1 U24082 ( .B1(n21112), .B2(n21096), .A(n21095), .ZN(P2_U3602) );
  INV_X1 U24083 ( .A(n21097), .ZN(n21102) );
  NOR2_X1 U24084 ( .A1(n21099), .A2(n21098), .ZN(n21101) );
  MUX2_X1 U24085 ( .A(n21102), .B(n21101), .S(n21100), .Z(n21103) );
  AOI21_X1 U24086 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n21104), .A(n21103), 
        .ZN(n21105) );
  AOI22_X1 U24087 ( .A1(n21115), .A2(n22183), .B1(n21105), .B2(n21112), .ZN(
        P2_U3603) );
  OAI22_X1 U24088 ( .A1(n21108), .A2(n21107), .B1(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n21106), .ZN(n21109) );
  AOI21_X1 U24089 ( .B1(n21111), .B2(n21110), .A(n21109), .ZN(n21113) );
  AOI22_X1 U24090 ( .A1(n21115), .A2(n21114), .B1(n21113), .B2(n21112), .ZN(
        P2_U3605) );
  AOI22_X1 U24091 ( .A1(n21140), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n21116), 
        .B2(n21141), .ZN(P2_U3608) );
  INV_X1 U24092 ( .A(n21117), .ZN(n21124) );
  NAND2_X1 U24093 ( .A1(n21119), .A2(n21118), .ZN(n21120) );
  AND2_X1 U24094 ( .A1(n21121), .A2(n21120), .ZN(n21123) );
  NAND2_X1 U24095 ( .A1(n21124), .A2(P2_MORE_REG_SCAN_IN), .ZN(n21122) );
  OAI21_X1 U24096 ( .B1(n21124), .B2(n21123), .A(n21122), .ZN(P2_U3609) );
  OAI22_X1 U24097 ( .A1(n10671), .A2(P2_STATE2_REG_3__SCAN_IN), .B1(n21126), 
        .B2(n21125), .ZN(n21127) );
  NOR2_X1 U24098 ( .A1(n21128), .A2(n21127), .ZN(n21139) );
  NOR3_X1 U24099 ( .A1(n21129), .A2(n9969), .A3(n21132), .ZN(n21131) );
  AOI21_X1 U24100 ( .B1(n21129), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n10922), 
        .ZN(n21130) );
  MUX2_X1 U24101 ( .A(n21131), .B(n21130), .S(n9735), .Z(n21136) );
  AOI21_X1 U24102 ( .B1(n21133), .B2(P2_STATE2_REG_2__SCAN_IN), .A(n21132), 
        .ZN(n21134) );
  NOR3_X1 U24103 ( .A1(n21136), .A2(n21135), .A3(n21134), .ZN(n21138) );
  NAND2_X1 U24104 ( .A1(n21139), .A2(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n21137) );
  OAI21_X1 U24105 ( .B1(n21139), .B2(n21138), .A(n21137), .ZN(P2_U3610) );
  OAI22_X1 U24106 ( .A1(n21141), .A2(P2_MEMORYFETCH_REG_SCAN_IN), .B1(
        P2_M_IO_N_REG_SCAN_IN), .B2(n21140), .ZN(n21142) );
  INV_X1 U24107 ( .A(n21142), .ZN(P2_U3611) );
  INV_X1 U24108 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n22171) );
  AOI21_X1 U24109 ( .B1(n21151), .B2(n22171), .A(n21915), .ZN(P1_U2802) );
  NAND2_X1 U24110 ( .A1(n21819), .A2(n21871), .ZN(n21149) );
  INV_X1 U24111 ( .A(n21145), .ZN(n21147) );
  OAI21_X1 U24112 ( .B1(n21147), .B2(n21146), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n21148) );
  OAI21_X1 U24113 ( .B1(n21149), .B2(n21908), .A(n21148), .ZN(P1_U2803) );
  NOR2_X1 U24114 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n21152) );
  OAI21_X1 U24115 ( .B1(n21152), .B2(P1_D_C_N_REG_SCAN_IN), .A(n21916), .ZN(
        n21150) );
  OAI21_X1 U24116 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n21916), .A(n21150), 
        .ZN(P1_U2804) );
  NOR2_X1 U24117 ( .A1(n21915), .A2(n21151), .ZN(n21895) );
  OAI21_X1 U24118 ( .B1(BS16), .B2(n21152), .A(n21895), .ZN(n21893) );
  OAI21_X1 U24119 ( .B1(n21895), .B2(n21905), .A(n21893), .ZN(P1_U2805) );
  OAI21_X1 U24120 ( .B1(n21154), .B2(n22052), .A(n21153), .ZN(P1_U2806) );
  NOR4_X1 U24121 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_21__SCAN_IN), .A3(P1_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_23__SCAN_IN), .ZN(n21158) );
  NOR4_X1 U24122 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_17__SCAN_IN), .A3(P1_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_19__SCAN_IN), .ZN(n21157) );
  NOR4_X1 U24123 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n21156) );
  NOR4_X1 U24124 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_27__SCAN_IN), .ZN(n21155) );
  NAND4_X1 U24125 ( .A1(n21158), .A2(n21157), .A3(n21156), .A4(n21155), .ZN(
        n21164) );
  NOR4_X1 U24126 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_5__SCAN_IN), .A3(P1_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_7__SCAN_IN), .ZN(n21162) );
  AOI211_X1 U24127 ( .C1(P1_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A(P1_DATAWIDTH_REG_2__SCAN_IN), .B(
        P1_DATAWIDTH_REG_3__SCAN_IN), .ZN(n21161) );
  NOR4_X1 U24128 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_13__SCAN_IN), .A3(P1_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_15__SCAN_IN), .ZN(n21160) );
  NOR4_X1 U24129 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_9__SCAN_IN), .A3(P1_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_11__SCAN_IN), .ZN(n21159) );
  NAND4_X1 U24130 ( .A1(n21162), .A2(n21161), .A3(n21160), .A4(n21159), .ZN(
        n21163) );
  NOR2_X1 U24131 ( .A1(n21164), .A2(n21163), .ZN(n21902) );
  INV_X1 U24132 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n21166) );
  NOR3_X1 U24133 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n21167) );
  OAI21_X1 U24134 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n21167), .A(n21902), .ZN(
        n21165) );
  OAI21_X1 U24135 ( .B1(n21902), .B2(n21166), .A(n21165), .ZN(P1_U2807) );
  INV_X1 U24136 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n21894) );
  AOI21_X1 U24137 ( .B1(n21896), .B2(n21894), .A(n21167), .ZN(n21169) );
  INV_X1 U24138 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n21168) );
  INV_X1 U24139 ( .A(n21902), .ZN(n21898) );
  AOI22_X1 U24140 ( .A1(n21902), .A2(n21169), .B1(n21168), .B2(n21898), .ZN(
        P1_U2808) );
  NAND2_X1 U24141 ( .A1(n21182), .A2(n21170), .ZN(n21216) );
  OAI21_X1 U24142 ( .B1(n21171), .B2(n21216), .A(n21217), .ZN(n21191) );
  AOI22_X1 U24143 ( .A1(n21223), .A2(P1_EBX_REG_9__SCAN_IN), .B1(n21259), .B2(
        n21172), .ZN(n21181) );
  INV_X1 U24144 ( .A(n21173), .ZN(n21179) );
  AOI22_X1 U24145 ( .A1(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n21233), .B1(
        n21175), .B2(n21174), .ZN(n21176) );
  OAI211_X1 U24146 ( .C1(n21177), .C2(P1_REIP_REG_9__SCAN_IN), .A(n21176), .B(
        n21235), .ZN(n21178) );
  AOI21_X1 U24147 ( .B1(n21179), .B2(n21212), .A(n21178), .ZN(n21180) );
  OAI211_X1 U24148 ( .C1(n21878), .C2(n21191), .A(n21181), .B(n21180), .ZN(
        P1_U2831) );
  NAND2_X1 U24149 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .ZN(n21193) );
  NAND2_X1 U24150 ( .A1(n21251), .A2(n21182), .ZN(n21219) );
  NOR2_X1 U24151 ( .A1(n21193), .A2(n21219), .ZN(n21201) );
  AOI21_X1 U24152 ( .B1(P1_REIP_REG_7__SCAN_IN), .B2(n21201), .A(
        P1_REIP_REG_8__SCAN_IN), .ZN(n21192) );
  AOI22_X1 U24153 ( .A1(n21223), .A2(P1_EBX_REG_8__SCAN_IN), .B1(n21259), .B2(
        n21183), .ZN(n21190) );
  INV_X1 U24154 ( .A(n21184), .ZN(n21188) );
  AOI21_X1 U24155 ( .B1(n21233), .B2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n21221), .ZN(n21185) );
  OAI21_X1 U24156 ( .B1(n21263), .B2(n21186), .A(n21185), .ZN(n21187) );
  AOI21_X1 U24157 ( .B1(n21188), .B2(n21212), .A(n21187), .ZN(n21189) );
  OAI211_X1 U24158 ( .C1(n21192), .C2(n21191), .A(n21190), .B(n21189), .ZN(
        P1_U2832) );
  OAI21_X1 U24159 ( .B1(n21193), .B2(n21216), .A(n21217), .ZN(n21215) );
  OAI21_X1 U24160 ( .B1(n21253), .B2(n21194), .A(n21235), .ZN(n21198) );
  OAI22_X1 U24161 ( .A1(n21263), .A2(n21196), .B1(n21195), .B2(n21256), .ZN(
        n21197) );
  AOI211_X1 U24162 ( .C1(n21259), .C2(n21199), .A(n21198), .B(n21197), .ZN(
        n21203) );
  AOI22_X1 U24163 ( .A1(n21204), .A2(n21201), .B1(n21200), .B2(n21212), .ZN(
        n21202) );
  OAI211_X1 U24164 ( .C1(n21204), .C2(n21215), .A(n21203), .B(n21202), .ZN(
        P1_U2833) );
  AOI22_X1 U24165 ( .A1(n21223), .A2(P1_EBX_REG_6__SCAN_IN), .B1(n21259), .B2(
        n21205), .ZN(n21214) );
  OAI21_X1 U24166 ( .B1(n21263), .B2(n21206), .A(n21235), .ZN(n21210) );
  NOR2_X1 U24167 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(n21219), .ZN(n21207) );
  AOI22_X1 U24168 ( .A1(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n21233), .B1(
        P1_REIP_REG_5__SCAN_IN), .B2(n21207), .ZN(n21208) );
  INV_X1 U24169 ( .A(n21208), .ZN(n21209) );
  AOI211_X1 U24170 ( .C1(n21212), .C2(n21211), .A(n21210), .B(n21209), .ZN(
        n21213) );
  OAI211_X1 U24171 ( .C1(n13596), .C2(n21215), .A(n21214), .B(n21213), .ZN(
        P1_U2834) );
  NAND2_X1 U24172 ( .A1(n21217), .A2(n21216), .ZN(n21246) );
  OAI22_X1 U24173 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(n21219), .B1(n21218), 
        .B2(n21263), .ZN(n21220) );
  AOI211_X1 U24174 ( .C1(n21233), .C2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n21221), .B(n21220), .ZN(n21229) );
  AOI22_X1 U24175 ( .A1(n21223), .A2(P1_EBX_REG_5__SCAN_IN), .B1(n21259), .B2(
        n21222), .ZN(n21224) );
  OAI21_X1 U24176 ( .B1(n21226), .B2(n21225), .A(n21224), .ZN(n21227) );
  INV_X1 U24177 ( .A(n21227), .ZN(n21228) );
  OAI211_X1 U24178 ( .C1(n15836), .C2(n21246), .A(n21229), .B(n21228), .ZN(
        P1_U2835) );
  NAND4_X1 U24179 ( .A1(n21251), .A2(P1_REIP_REG_3__SCAN_IN), .A3(
        P1_REIP_REG_1__SCAN_IN), .A4(P1_REIP_REG_2__SCAN_IN), .ZN(n21248) );
  INV_X1 U24180 ( .A(n21230), .ZN(n21244) );
  INV_X1 U24181 ( .A(n21231), .ZN(n21242) );
  AND2_X1 U24182 ( .A1(n21259), .A2(n21232), .ZN(n21238) );
  NAND2_X1 U24183 ( .A1(n21233), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n21234) );
  OAI211_X1 U24184 ( .C1(n21256), .C2(n21236), .A(n21235), .B(n21234), .ZN(
        n21237) );
  AOI211_X1 U24185 ( .C1(n21240), .C2(n21239), .A(n21238), .B(n21237), .ZN(
        n21241) );
  OAI21_X1 U24186 ( .B1(n21263), .B2(n21242), .A(n21241), .ZN(n21243) );
  AOI21_X1 U24187 ( .B1(n21244), .B2(n21265), .A(n21243), .ZN(n21245) );
  OAI221_X1 U24188 ( .B1(P1_REIP_REG_4__SCAN_IN), .B2(n21248), .C1(n21247), 
        .C2(n21246), .A(n21245), .ZN(P1_U2836) );
  NAND3_X1 U24189 ( .A1(n21251), .A2(P1_REIP_REG_1__SCAN_IN), .A3(
        P1_REIP_REG_2__SCAN_IN), .ZN(n21269) );
  AOI221_X1 U24190 ( .B1(n21896), .B2(n21251), .C1(n21250), .C2(n21251), .A(
        n21249), .ZN(n21268) );
  NOR2_X1 U24191 ( .A1(n9922), .A2(n21252), .ZN(n21258) );
  OAI22_X1 U24192 ( .A1(n21256), .A2(n21255), .B1(n21254), .B2(n21253), .ZN(
        n21257) );
  AOI211_X1 U24193 ( .C1(n21260), .C2(n21259), .A(n21258), .B(n21257), .ZN(
        n21261) );
  OAI21_X1 U24194 ( .B1(n21263), .B2(n21262), .A(n21261), .ZN(n21264) );
  AOI21_X1 U24195 ( .B1(n21266), .B2(n21265), .A(n21264), .ZN(n21267) );
  OAI221_X1 U24196 ( .B1(P1_REIP_REG_3__SCAN_IN), .B2(n21269), .C1(n22140), 
        .C2(n21268), .A(n21267), .ZN(P1_U2837) );
  INV_X1 U24197 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n22087) );
  INV_X1 U24198 ( .A(n21270), .ZN(n21271) );
  AOI22_X1 U24199 ( .A1(n21271), .A2(P1_EAX_REG_25__SCAN_IN), .B1(
        P1_UWORD_REG_9__SCAN_IN), .B2(n21299), .ZN(n21272) );
  OAI21_X1 U24200 ( .B1(n22087), .B2(n21285), .A(n21272), .ZN(P1_U2911) );
  AOI22_X1 U24201 ( .A1(P1_EAX_REG_15__SCAN_IN), .A2(n21283), .B1(n21298), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n21273) );
  OAI21_X1 U24202 ( .B1(n21274), .B2(n21281), .A(n21273), .ZN(P1_U2921) );
  INV_X1 U24203 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n21276) );
  AOI22_X1 U24204 ( .A1(P1_LWORD_REG_14__SCAN_IN), .A2(n21299), .B1(n21298), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n21275) );
  OAI21_X1 U24205 ( .B1(n21276), .B2(n21301), .A(n21275), .ZN(P1_U2922) );
  AOI22_X1 U24206 ( .A1(P1_LWORD_REG_13__SCAN_IN), .A2(n21299), .B1(n21298), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n21277) );
  OAI21_X1 U24207 ( .B1(n22101), .B2(n21301), .A(n21277), .ZN(P1_U2923) );
  INV_X1 U24208 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n21279) );
  AOI22_X1 U24209 ( .A1(P1_LWORD_REG_12__SCAN_IN), .A2(n21299), .B1(n21298), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n21278) );
  OAI21_X1 U24210 ( .B1(n21279), .B2(n21301), .A(n21278), .ZN(P1_U2924) );
  INV_X1 U24211 ( .A(P1_LWORD_REG_11__SCAN_IN), .ZN(n22004) );
  AOI22_X1 U24212 ( .A1(P1_EAX_REG_11__SCAN_IN), .A2(n21283), .B1(n21298), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n21280) );
  OAI21_X1 U24213 ( .B1(n22004), .B2(n21281), .A(n21280), .ZN(P1_U2925) );
  AOI22_X1 U24214 ( .A1(P1_LWORD_REG_10__SCAN_IN), .A2(n21299), .B1(n21298), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n21282) );
  OAI21_X1 U24215 ( .B1(n15289), .B2(n21301), .A(n21282), .ZN(P1_U2926) );
  AOI22_X1 U24216 ( .A1(P1_EAX_REG_9__SCAN_IN), .A2(n21283), .B1(
        P1_LWORD_REG_9__SCAN_IN), .B2(n21299), .ZN(n21284) );
  OAI21_X1 U24217 ( .B1(n22210), .B2(n21285), .A(n21284), .ZN(P1_U2927) );
  AOI22_X1 U24218 ( .A1(P1_LWORD_REG_8__SCAN_IN), .A2(n21299), .B1(n21298), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n21286) );
  OAI21_X1 U24219 ( .B1(n21287), .B2(n21301), .A(n21286), .ZN(P1_U2928) );
  AOI22_X1 U24220 ( .A1(P1_LWORD_REG_7__SCAN_IN), .A2(n21299), .B1(n21298), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n21288) );
  OAI21_X1 U24221 ( .B1(n15294), .B2(n21301), .A(n21288), .ZN(P1_U2929) );
  AOI22_X1 U24222 ( .A1(P1_LWORD_REG_6__SCAN_IN), .A2(n21299), .B1(n21298), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n21289) );
  OAI21_X1 U24223 ( .B1(n12726), .B2(n21301), .A(n21289), .ZN(P1_U2930) );
  AOI22_X1 U24224 ( .A1(P1_LWORD_REG_5__SCAN_IN), .A2(n21299), .B1(n21298), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n21290) );
  OAI21_X1 U24225 ( .B1(n22197), .B2(n21301), .A(n21290), .ZN(P1_U2931) );
  AOI22_X1 U24226 ( .A1(P1_LWORD_REG_4__SCAN_IN), .A2(n21299), .B1(n21298), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n21291) );
  OAI21_X1 U24227 ( .B1(n21292), .B2(n21301), .A(n21291), .ZN(P1_U2932) );
  AOI22_X1 U24228 ( .A1(P1_LWORD_REG_3__SCAN_IN), .A2(n21299), .B1(n21298), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n21293) );
  OAI21_X1 U24229 ( .B1(n15297), .B2(n21301), .A(n21293), .ZN(P1_U2933) );
  AOI22_X1 U24230 ( .A1(P1_LWORD_REG_2__SCAN_IN), .A2(n21299), .B1(n21298), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n21294) );
  OAI21_X1 U24231 ( .B1(n21295), .B2(n21301), .A(n21294), .ZN(P1_U2934) );
  AOI22_X1 U24232 ( .A1(P1_LWORD_REG_1__SCAN_IN), .A2(n21299), .B1(n21298), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n21296) );
  OAI21_X1 U24233 ( .B1(n21297), .B2(n21301), .A(n21296), .ZN(P1_U2935) );
  AOI22_X1 U24234 ( .A1(P1_LWORD_REG_0__SCAN_IN), .A2(n21299), .B1(n21298), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n21300) );
  OAI21_X1 U24235 ( .B1(n22214), .B2(n21301), .A(n21300), .ZN(P1_U2936) );
  AOI22_X1 U24236 ( .A1(n21322), .A2(P1_EAX_REG_25__SCAN_IN), .B1(
        P1_UWORD_REG_9__SCAN_IN), .B2(n15346), .ZN(n21304) );
  INV_X1 U24237 ( .A(n21302), .ZN(n21303) );
  NAND2_X1 U24238 ( .A1(n21311), .A2(n21303), .ZN(n21313) );
  NAND2_X1 U24239 ( .A1(n21304), .A2(n21313), .ZN(P1_U2946) );
  AOI22_X1 U24240 ( .A1(n21322), .A2(P1_EAX_REG_27__SCAN_IN), .B1(
        P1_UWORD_REG_11__SCAN_IN), .B2(n21321), .ZN(n21307) );
  INV_X1 U24241 ( .A(n21305), .ZN(n21306) );
  NAND2_X1 U24242 ( .A1(n21311), .A2(n21306), .ZN(n21317) );
  NAND2_X1 U24243 ( .A1(n21307), .A2(n21317), .ZN(P1_U2948) );
  AOI22_X1 U24244 ( .A1(n21322), .A2(P1_EAX_REG_28__SCAN_IN), .B1(
        P1_UWORD_REG_12__SCAN_IN), .B2(n21321), .ZN(n21309) );
  NAND2_X1 U24245 ( .A1(n21311), .A2(n21308), .ZN(n21319) );
  NAND2_X1 U24246 ( .A1(n21309), .A2(n21319), .ZN(P1_U2949) );
  AOI22_X1 U24247 ( .A1(n21322), .A2(P1_EAX_REG_30__SCAN_IN), .B1(
        P1_UWORD_REG_14__SCAN_IN), .B2(n21321), .ZN(n21312) );
  NAND2_X1 U24248 ( .A1(n21311), .A2(n21310), .ZN(n21323) );
  NAND2_X1 U24249 ( .A1(n21312), .A2(n21323), .ZN(P1_U2951) );
  AOI22_X1 U24250 ( .A1(n21322), .A2(P1_EAX_REG_9__SCAN_IN), .B1(
        P1_LWORD_REG_9__SCAN_IN), .B2(n21321), .ZN(n21314) );
  NAND2_X1 U24251 ( .A1(n21314), .A2(n21313), .ZN(P1_U2961) );
  AOI22_X1 U24252 ( .A1(n21322), .A2(P1_EAX_REG_10__SCAN_IN), .B1(
        P1_LWORD_REG_10__SCAN_IN), .B2(n21321), .ZN(n21316) );
  NAND2_X1 U24253 ( .A1(n21316), .A2(n21315), .ZN(P1_U2962) );
  AOI22_X1 U24254 ( .A1(n21322), .A2(P1_EAX_REG_11__SCAN_IN), .B1(
        P1_LWORD_REG_11__SCAN_IN), .B2(n21321), .ZN(n21318) );
  NAND2_X1 U24255 ( .A1(n21318), .A2(n21317), .ZN(P1_U2963) );
  AOI22_X1 U24256 ( .A1(n21322), .A2(P1_EAX_REG_12__SCAN_IN), .B1(
        P1_LWORD_REG_12__SCAN_IN), .B2(n21321), .ZN(n21320) );
  NAND2_X1 U24257 ( .A1(n21320), .A2(n21319), .ZN(P1_U2964) );
  AOI22_X1 U24258 ( .A1(n21322), .A2(P1_EAX_REG_14__SCAN_IN), .B1(
        P1_LWORD_REG_14__SCAN_IN), .B2(n21321), .ZN(n21324) );
  NAND2_X1 U24259 ( .A1(n21324), .A2(n21323), .ZN(P1_U2966) );
  NOR2_X1 U24260 ( .A1(n21326), .A2(n21325), .ZN(P1_U3032) );
  NAND2_X1 U24261 ( .A1(n21328), .A2(n21327), .ZN(n21369) );
  NAND2_X1 U24262 ( .A1(n21329), .A2(n21328), .ZN(n21370) );
  AOI22_X1 U24263 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n21372), .B1(DATAI_16_), 
        .B2(n21371), .ZN(n21739) );
  INV_X1 U24264 ( .A(n21330), .ZN(n21331) );
  INV_X1 U24265 ( .A(n21823), .ZN(n21736) );
  NOR2_X2 U24266 ( .A1(n21374), .A2(n21334), .ZN(n21811) );
  NAND2_X1 U24267 ( .A1(n21636), .A2(n21586), .ZN(n21437) );
  OR2_X1 U24268 ( .A1(n21698), .A2(n21437), .ZN(n21339) );
  AOI22_X1 U24269 ( .A1(n21865), .A2(n21736), .B1(n21811), .B2(n21375), .ZN(
        n21348) );
  INV_X1 U24270 ( .A(n21637), .ZN(n21335) );
  NOR2_X1 U24271 ( .A1(n21335), .A2(n21587), .ZN(n21344) );
  NAND2_X1 U24272 ( .A1(n21343), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n21773) );
  AND2_X1 U24273 ( .A1(n21773), .A2(n21336), .ZN(n21639) );
  NAND2_X1 U24274 ( .A1(n21401), .A2(n21819), .ZN(n21337) );
  NAND2_X1 U24275 ( .A1(n21819), .A2(n21905), .ZN(n21699) );
  OAI21_X1 U24276 ( .B1(n21337), .B2(n21865), .A(n21699), .ZN(n21342) );
  INV_X1 U24277 ( .A(n13896), .ZN(n21338) );
  NAND2_X1 U24278 ( .A1(n10664), .A2(n21702), .ZN(n21345) );
  AOI22_X1 U24279 ( .A1(n21342), .A2(n21345), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n21339), .ZN(n21340) );
  NOR2_X2 U24280 ( .A1(n21476), .A2(n21341), .ZN(n21812) );
  INV_X1 U24281 ( .A(n21342), .ZN(n21346) );
  INV_X1 U24282 ( .A(n21344), .ZN(n21472) );
  AOI22_X1 U24283 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n21378), .B1(
        n21812), .B2(n21377), .ZN(n21347) );
  OAI211_X1 U24284 ( .C1(n21739), .C2(n21401), .A(n21348), .B(n21347), .ZN(
        P1_U3033) );
  AOI22_X1 U24285 ( .A1(DATAI_17_), .A2(n21371), .B1(BUF1_REG_17__SCAN_IN), 
        .B2(n21372), .ZN(n21743) );
  AOI22_X1 U24286 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n21372), .B1(DATAI_25_), 
        .B2(n21371), .ZN(n21829) );
  INV_X1 U24287 ( .A(n21829), .ZN(n21740) );
  NOR2_X2 U24288 ( .A1(n21374), .A2(n12289), .ZN(n21824) );
  AOI22_X1 U24289 ( .A1(n21865), .A2(n21740), .B1(n21824), .B2(n21375), .ZN(
        n21351) );
  NOR2_X2 U24290 ( .A1(n21476), .A2(n21349), .ZN(n21825) );
  AOI22_X1 U24291 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n21378), .B1(
        n21825), .B2(n21377), .ZN(n21350) );
  OAI211_X1 U24292 ( .C1(n21743), .C2(n21401), .A(n21351), .B(n21350), .ZN(
        P1_U3034) );
  AOI22_X1 U24293 ( .A1(DATAI_18_), .A2(n21371), .B1(BUF1_REG_18__SCAN_IN), 
        .B2(n21372), .ZN(n21747) );
  AOI22_X1 U24294 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n21372), .B1(DATAI_26_), 
        .B2(n21371), .ZN(n21835) );
  INV_X1 U24295 ( .A(n21835), .ZN(n21744) );
  NOR2_X2 U24296 ( .A1(n21374), .A2(n13350), .ZN(n21830) );
  AOI22_X1 U24297 ( .A1(n21865), .A2(n21744), .B1(n21830), .B2(n21375), .ZN(
        n21354) );
  NOR2_X2 U24298 ( .A1(n21476), .A2(n21352), .ZN(n21831) );
  AOI22_X1 U24299 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n21378), .B1(
        n21831), .B2(n21377), .ZN(n21353) );
  OAI211_X1 U24300 ( .C1(n21747), .C2(n21401), .A(n21354), .B(n21353), .ZN(
        P1_U3035) );
  AOI22_X1 U24301 ( .A1(DATAI_19_), .A2(n21371), .B1(BUF1_REG_19__SCAN_IN), 
        .B2(n21372), .ZN(n21751) );
  AOI22_X1 U24302 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n21372), .B1(DATAI_27_), 
        .B2(n21371), .ZN(n21841) );
  INV_X1 U24303 ( .A(n21841), .ZN(n21748) );
  NOR2_X2 U24304 ( .A1(n21374), .A2(n12300), .ZN(n21836) );
  AOI22_X1 U24305 ( .A1(n21865), .A2(n21748), .B1(n21836), .B2(n21375), .ZN(
        n21357) );
  NOR2_X2 U24306 ( .A1(n21476), .A2(n21355), .ZN(n21837) );
  AOI22_X1 U24307 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n21378), .B1(
        n21837), .B2(n21377), .ZN(n21356) );
  OAI211_X1 U24308 ( .C1(n21751), .C2(n21401), .A(n21357), .B(n21356), .ZN(
        P1_U3036) );
  AOI22_X1 U24309 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n21372), .B1(DATAI_28_), 
        .B2(n21371), .ZN(n21847) );
  NOR2_X2 U24310 ( .A1(n21374), .A2(n12296), .ZN(n21842) );
  AOI22_X1 U24311 ( .A1(n21865), .A2(n21752), .B1(n21842), .B2(n21375), .ZN(
        n21360) );
  NOR2_X2 U24312 ( .A1(n21476), .A2(n21358), .ZN(n21843) );
  AOI22_X1 U24313 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n21378), .B1(
        n21843), .B2(n21377), .ZN(n21359) );
  OAI211_X1 U24314 ( .C1(n21755), .C2(n21401), .A(n21360), .B(n21359), .ZN(
        P1_U3037) );
  AOI22_X1 U24315 ( .A1(DATAI_21_), .A2(n21371), .B1(BUF1_REG_21__SCAN_IN), 
        .B2(n21372), .ZN(n21759) );
  INV_X1 U24316 ( .A(n21853), .ZN(n21756) );
  NOR2_X2 U24317 ( .A1(n21374), .A2(n21361), .ZN(n21848) );
  AOI22_X1 U24318 ( .A1(n21865), .A2(n21756), .B1(n21848), .B2(n21375), .ZN(
        n21364) );
  NOR2_X2 U24319 ( .A1(n21476), .A2(n21362), .ZN(n21849) );
  AOI22_X1 U24320 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n21378), .B1(
        n21849), .B2(n21377), .ZN(n21363) );
  OAI211_X1 U24321 ( .C1(n21759), .C2(n21401), .A(n21364), .B(n21363), .ZN(
        P1_U3038) );
  AOI22_X1 U24322 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n21372), .B1(DATAI_22_), 
        .B2(n21371), .ZN(n21763) );
  AOI22_X1 U24323 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n21372), .B1(DATAI_30_), 
        .B2(n21371), .ZN(n21859) );
  INV_X1 U24324 ( .A(n21859), .ZN(n21760) );
  NOR2_X2 U24325 ( .A1(n21374), .A2(n21365), .ZN(n21854) );
  AOI22_X1 U24326 ( .A1(n21865), .A2(n21760), .B1(n21854), .B2(n21375), .ZN(
        n21368) );
  NOR2_X2 U24327 ( .A1(n21476), .A2(n21366), .ZN(n21855) );
  AOI22_X1 U24328 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n21378), .B1(
        n21855), .B2(n21377), .ZN(n21367) );
  OAI211_X1 U24329 ( .C1(n21763), .C2(n21401), .A(n21368), .B(n21367), .ZN(
        P1_U3039) );
  INV_X1 U24330 ( .A(DATAI_23_), .ZN(n22174) );
  OAI22_X1 U24331 ( .A1(n22174), .A2(n21370), .B1(n16442), .B2(n21369), .ZN(
        n21864) );
  INV_X1 U24332 ( .A(n21864), .ZN(n21771) );
  AOI22_X1 U24333 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n21372), .B1(DATAI_31_), 
        .B2(n21371), .ZN(n21870) );
  INV_X1 U24334 ( .A(n21870), .ZN(n21766) );
  NOR2_X2 U24335 ( .A1(n21374), .A2(n21373), .ZN(n21861) );
  AOI22_X1 U24336 ( .A1(n21865), .A2(n21766), .B1(n21861), .B2(n21375), .ZN(
        n21380) );
  NOR2_X2 U24337 ( .A1(n21476), .A2(n21376), .ZN(n21863) );
  AOI22_X1 U24338 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n21378), .B1(
        n21863), .B2(n21377), .ZN(n21379) );
  OAI211_X1 U24339 ( .C1(n21771), .C2(n21401), .A(n21380), .B(n21379), .ZN(
        P1_U3040) );
  INV_X1 U24340 ( .A(n21381), .ZN(n21730) );
  NOR3_X2 U24341 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n21729), .A3(
        n21437), .ZN(n21402) );
  AOI21_X1 U24342 ( .B1(n10664), .B2(n21730), .A(n21402), .ZN(n21384) );
  NOR2_X1 U24343 ( .A1(n21437), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n21386) );
  INV_X1 U24344 ( .A(n21386), .ZN(n21382) );
  OAI22_X1 U24345 ( .A1(n21384), .A2(n21810), .B1(n21382), .B2(n12682), .ZN(
        n21403) );
  AOI22_X1 U24346 ( .A1(n21812), .A2(n21403), .B1(n21811), .B2(n21402), .ZN(
        n21388) );
  AOI21_X1 U24347 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n21729), .A(n21476), 
        .ZN(n21817) );
  INV_X1 U24348 ( .A(n21436), .ZN(n21383) );
  NOR2_X1 U24349 ( .A1(n21383), .A2(n21810), .ZN(n21440) );
  INV_X1 U24350 ( .A(n21699), .ZN(n21733) );
  OAI21_X1 U24351 ( .B1(n21440), .B2(n21733), .A(n21384), .ZN(n21385) );
  OAI211_X1 U24352 ( .C1(n21819), .C2(n21386), .A(n21817), .B(n21385), .ZN(
        n21405) );
  INV_X1 U24353 ( .A(n21401), .ZN(n21404) );
  AOI22_X1 U24354 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n21405), .B1(
        n21404), .B2(n21736), .ZN(n21387) );
  OAI211_X1 U24355 ( .C1(n21739), .C2(n21428), .A(n21388), .B(n21387), .ZN(
        P1_U3041) );
  AOI22_X1 U24356 ( .A1(n21825), .A2(n21403), .B1(n21824), .B2(n21402), .ZN(
        n21390) );
  AOI22_X1 U24357 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n21405), .B1(
        n21404), .B2(n21740), .ZN(n21389) );
  OAI211_X1 U24358 ( .C1(n21743), .C2(n21428), .A(n21390), .B(n21389), .ZN(
        P1_U3042) );
  AOI22_X1 U24359 ( .A1(n21831), .A2(n21403), .B1(n21830), .B2(n21402), .ZN(
        n21392) );
  INV_X1 U24360 ( .A(n21747), .ZN(n21832) );
  AOI22_X1 U24361 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n21405), .B1(
        n21430), .B2(n21832), .ZN(n21391) );
  OAI211_X1 U24362 ( .C1(n21835), .C2(n21401), .A(n21392), .B(n21391), .ZN(
        P1_U3043) );
  AOI22_X1 U24363 ( .A1(n21837), .A2(n21403), .B1(n21836), .B2(n21402), .ZN(
        n21394) );
  AOI22_X1 U24364 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n21405), .B1(
        n21404), .B2(n21748), .ZN(n21393) );
  OAI211_X1 U24365 ( .C1(n21751), .C2(n21428), .A(n21394), .B(n21393), .ZN(
        P1_U3044) );
  AOI22_X1 U24366 ( .A1(n21843), .A2(n21403), .B1(n21842), .B2(n21402), .ZN(
        n21396) );
  INV_X1 U24367 ( .A(n21755), .ZN(n21844) );
  AOI22_X1 U24368 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n21405), .B1(
        n21430), .B2(n21844), .ZN(n21395) );
  OAI211_X1 U24369 ( .C1(n21847), .C2(n21401), .A(n21396), .B(n21395), .ZN(
        P1_U3045) );
  AOI22_X1 U24370 ( .A1(n21849), .A2(n21403), .B1(n21848), .B2(n21402), .ZN(
        n21398) );
  INV_X1 U24371 ( .A(n21759), .ZN(n21850) );
  AOI22_X1 U24372 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n21405), .B1(
        n21430), .B2(n21850), .ZN(n21397) );
  OAI211_X1 U24373 ( .C1(n21853), .C2(n21401), .A(n21398), .B(n21397), .ZN(
        P1_U3046) );
  AOI22_X1 U24374 ( .A1(n21855), .A2(n21403), .B1(n21854), .B2(n21402), .ZN(
        n21400) );
  INV_X1 U24375 ( .A(n21763), .ZN(n21856) );
  AOI22_X1 U24376 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n21405), .B1(
        n21430), .B2(n21856), .ZN(n21399) );
  OAI211_X1 U24377 ( .C1(n21859), .C2(n21401), .A(n21400), .B(n21399), .ZN(
        P1_U3047) );
  AOI22_X1 U24378 ( .A1(n21863), .A2(n21403), .B1(n21861), .B2(n21402), .ZN(
        n21407) );
  AOI22_X1 U24379 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n21405), .B1(
        n21404), .B2(n21766), .ZN(n21406) );
  OAI211_X1 U24380 ( .C1(n21771), .C2(n21428), .A(n21407), .B(n21406), .ZN(
        P1_U3048) );
  NAND2_X1 U24381 ( .A1(n15884), .A2(n9734), .ZN(n21523) );
  INV_X1 U24382 ( .A(n21739), .ZN(n21820) );
  NOR3_X2 U24383 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21808), .A3(
        n21437), .ZN(n21429) );
  AOI22_X1 U24384 ( .A1(n21463), .A2(n21820), .B1(n21811), .B2(n21429), .ZN(
        n21415) );
  AOI21_X1 U24385 ( .B1(n21461), .B2(n21428), .A(n21905), .ZN(n21408) );
  NOR2_X1 U24386 ( .A1(n21408), .A2(n21810), .ZN(n21411) );
  NAND2_X1 U24387 ( .A1(n10664), .A2(n21778), .ZN(n21412) );
  INV_X1 U24388 ( .A(n21429), .ZN(n21409) );
  AOI22_X1 U24389 ( .A1(n21411), .A2(n21412), .B1(n21409), .B2(
        P1_STATE2_REG_3__SCAN_IN), .ZN(n21410) );
  OR2_X1 U24390 ( .A1(n21637), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n21530) );
  NAND2_X1 U24391 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n21530), .ZN(n21527) );
  NAND3_X1 U24392 ( .A1(n21639), .A2(n21410), .A3(n21527), .ZN(n21432) );
  INV_X1 U24393 ( .A(n21411), .ZN(n21413) );
  AOI22_X1 U24394 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n21432), .B1(
        n21812), .B2(n21431), .ZN(n21414) );
  OAI211_X1 U24395 ( .C1(n21823), .C2(n21428), .A(n21415), .B(n21414), .ZN(
        P1_U3049) );
  INV_X1 U24396 ( .A(n21743), .ZN(n21826) );
  AOI22_X1 U24397 ( .A1(n21463), .A2(n21826), .B1(n21824), .B2(n21429), .ZN(
        n21417) );
  AOI22_X1 U24398 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n21432), .B1(
        n21825), .B2(n21431), .ZN(n21416) );
  OAI211_X1 U24399 ( .C1(n21829), .C2(n21428), .A(n21417), .B(n21416), .ZN(
        P1_U3050) );
  AOI22_X1 U24400 ( .A1(n21463), .A2(n21832), .B1(n21830), .B2(n21429), .ZN(
        n21419) );
  AOI22_X1 U24401 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n21432), .B1(
        n21831), .B2(n21431), .ZN(n21418) );
  OAI211_X1 U24402 ( .C1(n21835), .C2(n21428), .A(n21419), .B(n21418), .ZN(
        P1_U3051) );
  INV_X1 U24403 ( .A(n21751), .ZN(n21838) );
  AOI22_X1 U24404 ( .A1(n21463), .A2(n21838), .B1(n21836), .B2(n21429), .ZN(
        n21421) );
  AOI22_X1 U24405 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n21432), .B1(
        n21837), .B2(n21431), .ZN(n21420) );
  OAI211_X1 U24406 ( .C1(n21841), .C2(n21428), .A(n21421), .B(n21420), .ZN(
        P1_U3052) );
  AOI22_X1 U24407 ( .A1(n21463), .A2(n21844), .B1(n21842), .B2(n21429), .ZN(
        n21423) );
  AOI22_X1 U24408 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n21432), .B1(
        n21843), .B2(n21431), .ZN(n21422) );
  OAI211_X1 U24409 ( .C1(n21847), .C2(n21428), .A(n21423), .B(n21422), .ZN(
        P1_U3053) );
  AOI22_X1 U24410 ( .A1(n21430), .A2(n21756), .B1(n21848), .B2(n21429), .ZN(
        n21425) );
  AOI22_X1 U24411 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n21432), .B1(
        n21849), .B2(n21431), .ZN(n21424) );
  OAI211_X1 U24412 ( .C1(n21759), .C2(n21461), .A(n21425), .B(n21424), .ZN(
        P1_U3054) );
  AOI22_X1 U24413 ( .A1(n21463), .A2(n21856), .B1(n21854), .B2(n21429), .ZN(
        n21427) );
  AOI22_X1 U24414 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n21432), .B1(
        n21855), .B2(n21431), .ZN(n21426) );
  OAI211_X1 U24415 ( .C1(n21859), .C2(n21428), .A(n21427), .B(n21426), .ZN(
        P1_U3055) );
  AOI22_X1 U24416 ( .A1(n21430), .A2(n21766), .B1(n21861), .B2(n21429), .ZN(
        n21434) );
  AOI22_X1 U24417 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n21432), .B1(
        n21863), .B2(n21431), .ZN(n21433) );
  OAI211_X1 U24418 ( .C1(n21771), .C2(n21461), .A(n21434), .B(n21433), .ZN(
        P1_U3056) );
  INV_X1 U24419 ( .A(n21666), .ZN(n21435) );
  NOR2_X1 U24420 ( .A1(n21804), .A2(n21437), .ZN(n21462) );
  AOI22_X1 U24421 ( .A1(n21463), .A2(n21736), .B1(n21811), .B2(n21462), .ZN(
        n21448) );
  NOR2_X1 U24422 ( .A1(n21808), .A2(n21437), .ZN(n21443) );
  INV_X1 U24423 ( .A(n21438), .ZN(n21439) );
  AND2_X1 U24424 ( .A1(n21439), .A2(n12709), .ZN(n21805) );
  AOI21_X1 U24425 ( .B1(n10664), .B2(n21805), .A(n21462), .ZN(n21442) );
  NAND2_X1 U24426 ( .A1(n21442), .A2(n21444), .ZN(n21441) );
  OAI211_X1 U24427 ( .C1(n21819), .C2(n21443), .A(n21817), .B(n21441), .ZN(
        n21465) );
  INV_X1 U24428 ( .A(n21442), .ZN(n21445) );
  AOI22_X1 U24429 ( .A1(n21445), .A2(n21444), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n21443), .ZN(n21446) );
  AOI22_X1 U24430 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n21465), .B1(
        n21812), .B2(n21464), .ZN(n21447) );
  OAI211_X1 U24431 ( .C1(n21739), .C2(n21468), .A(n21448), .B(n21447), .ZN(
        P1_U3057) );
  AOI22_X1 U24432 ( .A1(n21463), .A2(n21740), .B1(n21824), .B2(n21462), .ZN(
        n21450) );
  AOI22_X1 U24433 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n21465), .B1(
        n21825), .B2(n21464), .ZN(n21449) );
  OAI211_X1 U24434 ( .C1(n21743), .C2(n21468), .A(n21450), .B(n21449), .ZN(
        P1_U3058) );
  AOI22_X1 U24435 ( .A1(n21463), .A2(n21744), .B1(n21830), .B2(n21462), .ZN(
        n21452) );
  AOI22_X1 U24436 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n21465), .B1(
        n21831), .B2(n21464), .ZN(n21451) );
  OAI211_X1 U24437 ( .C1(n21747), .C2(n21468), .A(n21452), .B(n21451), .ZN(
        P1_U3059) );
  AOI22_X1 U24438 ( .A1(n21463), .A2(n21748), .B1(n21836), .B2(n21462), .ZN(
        n21454) );
  AOI22_X1 U24439 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n21465), .B1(
        n21837), .B2(n21464), .ZN(n21453) );
  OAI211_X1 U24440 ( .C1(n21751), .C2(n21468), .A(n21454), .B(n21453), .ZN(
        P1_U3060) );
  AOI22_X1 U24441 ( .A1(n21463), .A2(n21752), .B1(n21842), .B2(n21462), .ZN(
        n21456) );
  AOI22_X1 U24442 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n21465), .B1(
        n21843), .B2(n21464), .ZN(n21455) );
  OAI211_X1 U24443 ( .C1(n21755), .C2(n21468), .A(n21456), .B(n21455), .ZN(
        P1_U3061) );
  AOI22_X1 U24444 ( .A1(n21494), .A2(n21850), .B1(n21848), .B2(n21462), .ZN(
        n21458) );
  AOI22_X1 U24445 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n21465), .B1(
        n21849), .B2(n21464), .ZN(n21457) );
  OAI211_X1 U24446 ( .C1(n21853), .C2(n21461), .A(n21458), .B(n21457), .ZN(
        P1_U3062) );
  AOI22_X1 U24447 ( .A1(n21494), .A2(n21856), .B1(n21854), .B2(n21462), .ZN(
        n21460) );
  AOI22_X1 U24448 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n21465), .B1(
        n21855), .B2(n21464), .ZN(n21459) );
  OAI211_X1 U24449 ( .C1(n21859), .C2(n21461), .A(n21460), .B(n21459), .ZN(
        P1_U3063) );
  AOI22_X1 U24450 ( .A1(n21463), .A2(n21766), .B1(n21861), .B2(n21462), .ZN(
        n21467) );
  AOI22_X1 U24451 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n21465), .B1(
        n21863), .B2(n21464), .ZN(n21466) );
  OAI211_X1 U24452 ( .C1(n21771), .C2(n21468), .A(n21467), .B(n21466), .ZN(
        P1_U3064) );
  NOR2_X1 U24453 ( .A1(n13896), .A2(n21470), .ZN(n21555) );
  NAND3_X1 U24454 ( .A1(n21555), .A2(n21819), .A3(n21702), .ZN(n21471) );
  AOI22_X1 U24455 ( .A1(n21812), .A2(n21493), .B1(n21811), .B2(n10676), .ZN(
        n21480) );
  INV_X1 U24456 ( .A(n21555), .ZN(n21475) );
  INV_X1 U24457 ( .A(n21522), .ZN(n21473) );
  OAI21_X1 U24458 ( .B1(n21494), .B2(n21473), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n21474) );
  OAI21_X1 U24459 ( .B1(n21778), .B2(n21475), .A(n21474), .ZN(n21478) );
  INV_X1 U24460 ( .A(n21642), .ZN(n21477) );
  AOI22_X1 U24461 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n21495), .B1(
        n21494), .B2(n21736), .ZN(n21479) );
  OAI211_X1 U24462 ( .C1(n21739), .C2(n21522), .A(n21480), .B(n21479), .ZN(
        P1_U3065) );
  AOI22_X1 U24463 ( .A1(n21825), .A2(n21493), .B1(n21824), .B2(n10676), .ZN(
        n21482) );
  AOI22_X1 U24464 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n21495), .B1(
        n21494), .B2(n21740), .ZN(n21481) );
  OAI211_X1 U24465 ( .C1(n21743), .C2(n21522), .A(n21482), .B(n21481), .ZN(
        P1_U3066) );
  AOI22_X1 U24466 ( .A1(n21831), .A2(n21493), .B1(n21830), .B2(n10676), .ZN(
        n21484) );
  AOI22_X1 U24467 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n21495), .B1(
        n21494), .B2(n21744), .ZN(n21483) );
  OAI211_X1 U24468 ( .C1(n21747), .C2(n21522), .A(n21484), .B(n21483), .ZN(
        P1_U3067) );
  AOI22_X1 U24469 ( .A1(n21837), .A2(n21493), .B1(n21836), .B2(n10676), .ZN(
        n21486) );
  AOI22_X1 U24470 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n21495), .B1(
        n21494), .B2(n21748), .ZN(n21485) );
  OAI211_X1 U24471 ( .C1(n21751), .C2(n21522), .A(n21486), .B(n21485), .ZN(
        P1_U3068) );
  AOI22_X1 U24472 ( .A1(n21843), .A2(n21493), .B1(n21842), .B2(n10676), .ZN(
        n21488) );
  AOI22_X1 U24473 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n21495), .B1(
        n21494), .B2(n21752), .ZN(n21487) );
  OAI211_X1 U24474 ( .C1(n21755), .C2(n21522), .A(n21488), .B(n21487), .ZN(
        P1_U3069) );
  AOI22_X1 U24475 ( .A1(n21849), .A2(n21493), .B1(n21848), .B2(n10676), .ZN(
        n21490) );
  AOI22_X1 U24476 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n21495), .B1(
        n21494), .B2(n21756), .ZN(n21489) );
  OAI211_X1 U24477 ( .C1(n21759), .C2(n21522), .A(n21490), .B(n21489), .ZN(
        P1_U3070) );
  AOI22_X1 U24478 ( .A1(n21855), .A2(n21493), .B1(n21854), .B2(n10676), .ZN(
        n21492) );
  AOI22_X1 U24479 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n21495), .B1(
        n21494), .B2(n21760), .ZN(n21491) );
  OAI211_X1 U24480 ( .C1(n21763), .C2(n21522), .A(n21492), .B(n21491), .ZN(
        P1_U3071) );
  AOI22_X1 U24481 ( .A1(n21863), .A2(n21493), .B1(n21861), .B2(n10676), .ZN(
        n21497) );
  AOI22_X1 U24482 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n21495), .B1(
        n21494), .B2(n21766), .ZN(n21496) );
  OAI211_X1 U24483 ( .C1(n21771), .C2(n21522), .A(n21497), .B(n21496), .ZN(
        P1_U3072) );
  NOR2_X1 U24484 ( .A1(n21524), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n21501) );
  INV_X1 U24485 ( .A(n21501), .ZN(n21498) );
  NOR2_X1 U24486 ( .A1(n21729), .A2(n21498), .ZN(n21517) );
  AOI21_X1 U24487 ( .B1(n21555), .B2(n21730), .A(n21517), .ZN(n21499) );
  OAI22_X1 U24488 ( .A1(n21499), .A2(n21810), .B1(n21498), .B2(n12682), .ZN(
        n21518) );
  AOI22_X1 U24489 ( .A1(n21812), .A2(n21518), .B1(n21811), .B2(n21517), .ZN(
        n21504) );
  NOR2_X1 U24490 ( .A1(n21561), .A2(n21810), .ZN(n21558) );
  OAI21_X1 U24491 ( .B1(n21558), .B2(n21733), .A(n21499), .ZN(n21500) );
  OAI211_X1 U24492 ( .C1(n21819), .C2(n21501), .A(n21817), .B(n21500), .ZN(
        n21519) );
  NAND2_X1 U24493 ( .A1(n21561), .A2(n21728), .ZN(n21553) );
  AOI22_X1 U24494 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n21519), .B1(
        n21541), .B2(n21820), .ZN(n21503) );
  OAI211_X1 U24495 ( .C1(n21823), .C2(n21522), .A(n21504), .B(n21503), .ZN(
        P1_U3073) );
  AOI22_X1 U24496 ( .A1(n21825), .A2(n21518), .B1(n21824), .B2(n21517), .ZN(
        n21506) );
  AOI22_X1 U24497 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n21519), .B1(
        n21541), .B2(n21826), .ZN(n21505) );
  OAI211_X1 U24498 ( .C1(n21829), .C2(n21522), .A(n21506), .B(n21505), .ZN(
        P1_U3074) );
  AOI22_X1 U24499 ( .A1(n21831), .A2(n21518), .B1(n21830), .B2(n21517), .ZN(
        n21508) );
  AOI22_X1 U24500 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n21519), .B1(
        n21541), .B2(n21832), .ZN(n21507) );
  OAI211_X1 U24501 ( .C1(n21835), .C2(n21522), .A(n21508), .B(n21507), .ZN(
        P1_U3075) );
  AOI22_X1 U24502 ( .A1(n21837), .A2(n21518), .B1(n21836), .B2(n21517), .ZN(
        n21510) );
  AOI22_X1 U24503 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n21519), .B1(
        n21541), .B2(n21838), .ZN(n21509) );
  OAI211_X1 U24504 ( .C1(n21841), .C2(n21522), .A(n21510), .B(n21509), .ZN(
        P1_U3076) );
  AOI22_X1 U24505 ( .A1(n21843), .A2(n21518), .B1(n21842), .B2(n21517), .ZN(
        n21512) );
  AOI22_X1 U24506 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n21519), .B1(
        n21541), .B2(n21844), .ZN(n21511) );
  OAI211_X1 U24507 ( .C1(n21847), .C2(n21522), .A(n21512), .B(n21511), .ZN(
        P1_U3077) );
  AOI22_X1 U24508 ( .A1(n21849), .A2(n21518), .B1(n21848), .B2(n21517), .ZN(
        n21514) );
  AOI22_X1 U24509 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n21519), .B1(
        n21541), .B2(n21850), .ZN(n21513) );
  OAI211_X1 U24510 ( .C1(n21853), .C2(n21522), .A(n21514), .B(n21513), .ZN(
        P1_U3078) );
  AOI22_X1 U24511 ( .A1(n21855), .A2(n21518), .B1(n21854), .B2(n21517), .ZN(
        n21516) );
  AOI22_X1 U24512 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n21519), .B1(
        n21541), .B2(n21856), .ZN(n21515) );
  OAI211_X1 U24513 ( .C1(n21859), .C2(n21522), .A(n21516), .B(n21515), .ZN(
        P1_U3079) );
  AOI22_X1 U24514 ( .A1(n21863), .A2(n21518), .B1(n21861), .B2(n21517), .ZN(
        n21521) );
  AOI22_X1 U24515 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n21519), .B1(
        n21541), .B2(n21864), .ZN(n21520) );
  OAI211_X1 U24516 ( .C1(n21870), .C2(n21522), .A(n21521), .B(n21520), .ZN(
        P1_U3080) );
  NOR2_X1 U24517 ( .A1(n21808), .A2(n21524), .ZN(n21560) );
  NAND2_X1 U24518 ( .A1(n21729), .A2(n21560), .ZN(n21526) );
  AOI22_X1 U24519 ( .A1(n21541), .A2(n21736), .B1(n21811), .B2(n21548), .ZN(
        n21534) );
  NAND2_X1 U24520 ( .A1(n21583), .A2(n21553), .ZN(n21525) );
  AOI21_X1 U24521 ( .B1(n21525), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n21810), 
        .ZN(n21529) );
  NAND2_X1 U24522 ( .A1(n21555), .A2(n21778), .ZN(n21531) );
  AOI22_X1 U24523 ( .A1(n21529), .A2(n21531), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n21526), .ZN(n21528) );
  NAND3_X1 U24524 ( .A1(n21781), .A2(n21528), .A3(n21527), .ZN(n21550) );
  INV_X1 U24525 ( .A(n21529), .ZN(n21532) );
  AOI22_X1 U24526 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n21550), .B1(
        n21812), .B2(n21549), .ZN(n21533) );
  OAI211_X1 U24527 ( .C1(n21739), .C2(n21583), .A(n21534), .B(n21533), .ZN(
        P1_U3081) );
  AOI22_X1 U24528 ( .A1(n21541), .A2(n21740), .B1(n21824), .B2(n21548), .ZN(
        n21536) );
  AOI22_X1 U24529 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n21550), .B1(
        n21825), .B2(n21549), .ZN(n21535) );
  OAI211_X1 U24530 ( .C1(n21743), .C2(n21583), .A(n21536), .B(n21535), .ZN(
        P1_U3082) );
  AOI22_X1 U24531 ( .A1(n21541), .A2(n21744), .B1(n21830), .B2(n21548), .ZN(
        n21538) );
  AOI22_X1 U24532 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n21550), .B1(
        n21831), .B2(n21549), .ZN(n21537) );
  OAI211_X1 U24533 ( .C1(n21747), .C2(n21583), .A(n21538), .B(n21537), .ZN(
        P1_U3083) );
  AOI22_X1 U24534 ( .A1(n21541), .A2(n21748), .B1(n21836), .B2(n21548), .ZN(
        n21540) );
  AOI22_X1 U24535 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n21550), .B1(
        n21837), .B2(n21549), .ZN(n21539) );
  OAI211_X1 U24536 ( .C1(n21751), .C2(n21583), .A(n21540), .B(n21539), .ZN(
        P1_U3084) );
  AOI22_X1 U24537 ( .A1(n21541), .A2(n21752), .B1(n21842), .B2(n21548), .ZN(
        n21543) );
  AOI22_X1 U24538 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n21550), .B1(
        n21843), .B2(n21549), .ZN(n21542) );
  OAI211_X1 U24539 ( .C1(n21755), .C2(n21583), .A(n21543), .B(n21542), .ZN(
        P1_U3085) );
  AOI22_X1 U24540 ( .A1(n21574), .A2(n21850), .B1(n21848), .B2(n21548), .ZN(
        n21545) );
  AOI22_X1 U24541 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n21550), .B1(
        n21849), .B2(n21549), .ZN(n21544) );
  OAI211_X1 U24542 ( .C1(n21853), .C2(n21553), .A(n21545), .B(n21544), .ZN(
        P1_U3086) );
  AOI22_X1 U24543 ( .A1(n21574), .A2(n21856), .B1(n21854), .B2(n21548), .ZN(
        n21547) );
  AOI22_X1 U24544 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n21550), .B1(
        n21855), .B2(n21549), .ZN(n21546) );
  OAI211_X1 U24545 ( .C1(n21859), .C2(n21553), .A(n21547), .B(n21546), .ZN(
        P1_U3087) );
  AOI22_X1 U24546 ( .A1(n21574), .A2(n21864), .B1(n21861), .B2(n21548), .ZN(
        n21552) );
  AOI22_X1 U24547 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n21550), .B1(
        n21863), .B2(n21549), .ZN(n21551) );
  OAI211_X1 U24548 ( .C1(n21870), .C2(n21553), .A(n21552), .B(n21551), .ZN(
        P1_U3088) );
  INV_X1 U24549 ( .A(n21554), .ZN(n21578) );
  AOI21_X1 U24550 ( .B1(n21555), .B2(n21805), .A(n21578), .ZN(n21557) );
  INV_X1 U24551 ( .A(n21560), .ZN(n21556) );
  OAI22_X1 U24552 ( .A1(n21557), .A2(n21810), .B1(n21556), .B2(n12682), .ZN(
        n21579) );
  AOI22_X1 U24553 ( .A1(n21812), .A2(n21579), .B1(n21578), .B2(n21811), .ZN(
        n21563) );
  OAI21_X1 U24554 ( .B1(n21815), .B2(n21558), .A(n21557), .ZN(n21559) );
  OAI211_X1 U24555 ( .C1(n21819), .C2(n21560), .A(n21817), .B(n21559), .ZN(
        n21580) );
  NAND2_X1 U24556 ( .A1(n21561), .A2(n21666), .ZN(n21577) );
  AOI22_X1 U24557 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n21580), .B1(
        n21607), .B2(n21820), .ZN(n21562) );
  OAI211_X1 U24558 ( .C1(n21823), .C2(n21583), .A(n21563), .B(n21562), .ZN(
        P1_U3089) );
  AOI22_X1 U24559 ( .A1(n21825), .A2(n21579), .B1(n21578), .B2(n21824), .ZN(
        n21565) );
  AOI22_X1 U24560 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n21580), .B1(
        n21607), .B2(n21826), .ZN(n21564) );
  OAI211_X1 U24561 ( .C1(n21829), .C2(n21583), .A(n21565), .B(n21564), .ZN(
        P1_U3090) );
  AOI22_X1 U24562 ( .A1(n21831), .A2(n21579), .B1(n21578), .B2(n21830), .ZN(
        n21567) );
  AOI22_X1 U24563 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n21580), .B1(
        n21574), .B2(n21744), .ZN(n21566) );
  OAI211_X1 U24564 ( .C1(n21747), .C2(n21577), .A(n21567), .B(n21566), .ZN(
        P1_U3091) );
  AOI22_X1 U24565 ( .A1(n21837), .A2(n21579), .B1(n21578), .B2(n21836), .ZN(
        n21569) );
  AOI22_X1 U24566 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n21580), .B1(
        n21607), .B2(n21838), .ZN(n21568) );
  OAI211_X1 U24567 ( .C1(n21841), .C2(n21583), .A(n21569), .B(n21568), .ZN(
        P1_U3092) );
  AOI22_X1 U24568 ( .A1(n21843), .A2(n21579), .B1(n21578), .B2(n21842), .ZN(
        n21571) );
  AOI22_X1 U24569 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n21580), .B1(
        n21574), .B2(n21752), .ZN(n21570) );
  OAI211_X1 U24570 ( .C1(n21755), .C2(n21577), .A(n21571), .B(n21570), .ZN(
        P1_U3093) );
  AOI22_X1 U24571 ( .A1(n21849), .A2(n21579), .B1(n21578), .B2(n21848), .ZN(
        n21573) );
  AOI22_X1 U24572 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n21580), .B1(
        n21607), .B2(n21850), .ZN(n21572) );
  OAI211_X1 U24573 ( .C1(n21853), .C2(n21583), .A(n21573), .B(n21572), .ZN(
        P1_U3094) );
  AOI22_X1 U24574 ( .A1(n21855), .A2(n21579), .B1(n21578), .B2(n21854), .ZN(
        n21576) );
  AOI22_X1 U24575 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n21580), .B1(
        n21574), .B2(n21760), .ZN(n21575) );
  OAI211_X1 U24576 ( .C1(n21763), .C2(n21577), .A(n21576), .B(n21575), .ZN(
        P1_U3095) );
  AOI22_X1 U24577 ( .A1(n21863), .A2(n21579), .B1(n21578), .B2(n21861), .ZN(
        n21582) );
  AOI22_X1 U24578 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n21580), .B1(
        n21607), .B2(n21864), .ZN(n21581) );
  OAI211_X1 U24579 ( .C1(n21870), .C2(n21583), .A(n21582), .B(n21581), .ZN(
        P1_U3096) );
  AND2_X1 U24580 ( .A1(n21585), .A2(n13896), .ZN(n21669) );
  NAND2_X1 U24581 ( .A1(n21586), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n21668) );
  AOI21_X1 U24582 ( .B1(n21669), .B2(n21702), .A(n10679), .ZN(n21589) );
  NAND2_X1 U24583 ( .A1(n21587), .A2(n21637), .ZN(n21706) );
  OAI22_X1 U24584 ( .A1(n21589), .A2(n21810), .B1(n21642), .B2(n21706), .ZN(
        n21606) );
  AOI22_X1 U24585 ( .A1(n21812), .A2(n21606), .B1(n10679), .B2(n21811), .ZN(
        n21593) );
  INV_X1 U24586 ( .A(n21634), .ZN(n21588) );
  OAI21_X1 U24587 ( .B1(n21588), .B2(n21607), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n21590) );
  NAND2_X1 U24588 ( .A1(n21590), .A2(n21589), .ZN(n21591) );
  AOI22_X1 U24589 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n21608), .B1(
        n21607), .B2(n21736), .ZN(n21592) );
  OAI211_X1 U24590 ( .C1(n21739), .C2(n21634), .A(n21593), .B(n21592), .ZN(
        P1_U3097) );
  AOI22_X1 U24591 ( .A1(n21825), .A2(n21606), .B1(n10679), .B2(n21824), .ZN(
        n21595) );
  AOI22_X1 U24592 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n21608), .B1(
        n21607), .B2(n21740), .ZN(n21594) );
  OAI211_X1 U24593 ( .C1(n21743), .C2(n21634), .A(n21595), .B(n21594), .ZN(
        P1_U3098) );
  AOI22_X1 U24594 ( .A1(n21831), .A2(n21606), .B1(n10679), .B2(n21830), .ZN(
        n21597) );
  AOI22_X1 U24595 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n21608), .B1(
        n21607), .B2(n21744), .ZN(n21596) );
  OAI211_X1 U24596 ( .C1(n21747), .C2(n21634), .A(n21597), .B(n21596), .ZN(
        P1_U3099) );
  AOI22_X1 U24597 ( .A1(n21837), .A2(n21606), .B1(n10679), .B2(n21836), .ZN(
        n21599) );
  AOI22_X1 U24598 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n21608), .B1(
        n21607), .B2(n21748), .ZN(n21598) );
  OAI211_X1 U24599 ( .C1(n21751), .C2(n21634), .A(n21599), .B(n21598), .ZN(
        P1_U3100) );
  AOI22_X1 U24600 ( .A1(n21843), .A2(n21606), .B1(n10679), .B2(n21842), .ZN(
        n21601) );
  AOI22_X1 U24601 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n21608), .B1(
        n21607), .B2(n21752), .ZN(n21600) );
  OAI211_X1 U24602 ( .C1(n21755), .C2(n21634), .A(n21601), .B(n21600), .ZN(
        P1_U3101) );
  AOI22_X1 U24603 ( .A1(n21849), .A2(n21606), .B1(n10679), .B2(n21848), .ZN(
        n21603) );
  AOI22_X1 U24604 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n21608), .B1(
        n21607), .B2(n21756), .ZN(n21602) );
  OAI211_X1 U24605 ( .C1(n21759), .C2(n21634), .A(n21603), .B(n21602), .ZN(
        P1_U3102) );
  AOI22_X1 U24606 ( .A1(n21855), .A2(n21606), .B1(n10679), .B2(n21854), .ZN(
        n21605) );
  AOI22_X1 U24607 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n21608), .B1(
        n21607), .B2(n21760), .ZN(n21604) );
  OAI211_X1 U24608 ( .C1(n21763), .C2(n21634), .A(n21605), .B(n21604), .ZN(
        P1_U3103) );
  AOI22_X1 U24609 ( .A1(n21863), .A2(n21606), .B1(n10679), .B2(n21861), .ZN(
        n21610) );
  AOI22_X1 U24610 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n21608), .B1(
        n21607), .B2(n21766), .ZN(n21609) );
  OAI211_X1 U24611 ( .C1(n21771), .C2(n21634), .A(n21610), .B(n21609), .ZN(
        P1_U3104) );
  NOR2_X1 U24612 ( .A1(n21668), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n21614) );
  INV_X1 U24613 ( .A(n21614), .ZN(n21611) );
  NOR2_X1 U24614 ( .A1(n21729), .A2(n21611), .ZN(n21629) );
  AOI21_X1 U24615 ( .B1(n21669), .B2(n21730), .A(n21629), .ZN(n21612) );
  OAI22_X1 U24616 ( .A1(n21612), .A2(n21810), .B1(n21611), .B2(n12682), .ZN(
        n21630) );
  AOI22_X1 U24617 ( .A1(n21812), .A2(n21630), .B1(n21811), .B2(n21629), .ZN(
        n21616) );
  NOR2_X1 U24618 ( .A1(n21667), .A2(n21810), .ZN(n21672) );
  OAI21_X1 U24619 ( .B1(n21672), .B2(n21733), .A(n21612), .ZN(n21613) );
  OAI211_X1 U24620 ( .C1(n21819), .C2(n21614), .A(n21817), .B(n21613), .ZN(
        n21631) );
  AOI22_X1 U24621 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n21631), .B1(
        n21655), .B2(n21820), .ZN(n21615) );
  OAI211_X1 U24622 ( .C1(n21823), .C2(n21634), .A(n21616), .B(n21615), .ZN(
        P1_U3105) );
  AOI22_X1 U24623 ( .A1(n21825), .A2(n21630), .B1(n21824), .B2(n21629), .ZN(
        n21618) );
  AOI22_X1 U24624 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n21631), .B1(
        n21655), .B2(n21826), .ZN(n21617) );
  OAI211_X1 U24625 ( .C1(n21829), .C2(n21634), .A(n21618), .B(n21617), .ZN(
        P1_U3106) );
  AOI22_X1 U24626 ( .A1(n21831), .A2(n21630), .B1(n21830), .B2(n21629), .ZN(
        n21620) );
  AOI22_X1 U24627 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n21631), .B1(
        n21655), .B2(n21832), .ZN(n21619) );
  OAI211_X1 U24628 ( .C1(n21835), .C2(n21634), .A(n21620), .B(n21619), .ZN(
        P1_U3107) );
  AOI22_X1 U24629 ( .A1(n21837), .A2(n21630), .B1(n21836), .B2(n21629), .ZN(
        n21622) );
  AOI22_X1 U24630 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n21631), .B1(
        n21655), .B2(n21838), .ZN(n21621) );
  OAI211_X1 U24631 ( .C1(n21841), .C2(n21634), .A(n21622), .B(n21621), .ZN(
        P1_U3108) );
  AOI22_X1 U24632 ( .A1(n21843), .A2(n21630), .B1(n21842), .B2(n21629), .ZN(
        n21624) );
  AOI22_X1 U24633 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n21631), .B1(
        n21655), .B2(n21844), .ZN(n21623) );
  OAI211_X1 U24634 ( .C1(n21847), .C2(n21634), .A(n21624), .B(n21623), .ZN(
        P1_U3109) );
  AOI22_X1 U24635 ( .A1(n21849), .A2(n21630), .B1(n21848), .B2(n21629), .ZN(
        n21626) );
  AOI22_X1 U24636 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n21631), .B1(
        n21655), .B2(n21850), .ZN(n21625) );
  OAI211_X1 U24637 ( .C1(n21853), .C2(n21634), .A(n21626), .B(n21625), .ZN(
        P1_U3110) );
  AOI22_X1 U24638 ( .A1(n21855), .A2(n21630), .B1(n21854), .B2(n21629), .ZN(
        n21628) );
  AOI22_X1 U24639 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n21631), .B1(
        n21655), .B2(n21856), .ZN(n21627) );
  OAI211_X1 U24640 ( .C1(n21859), .C2(n21634), .A(n21628), .B(n21627), .ZN(
        P1_U3111) );
  AOI22_X1 U24641 ( .A1(n21863), .A2(n21630), .B1(n21861), .B2(n21629), .ZN(
        n21633) );
  AOI22_X1 U24642 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n21631), .B1(
        n21655), .B2(n21864), .ZN(n21632) );
  OAI211_X1 U24643 ( .C1(n21870), .C2(n21634), .A(n21633), .B(n21632), .ZN(
        P1_U3112) );
  NOR2_X1 U24644 ( .A1(n21808), .A2(n21668), .ZN(n21674) );
  INV_X1 U24645 ( .A(n21674), .ZN(n21670) );
  NOR2_X1 U24646 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21670), .ZN(
        n21660) );
  AOI22_X1 U24647 ( .A1(n21687), .A2(n21820), .B1(n21811), .B2(n21660), .ZN(
        n21646) );
  OAI21_X1 U24648 ( .B1(n21687), .B2(n21655), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n21635) );
  NAND2_X1 U24649 ( .A1(n21635), .A2(n21819), .ZN(n21644) );
  AND2_X1 U24650 ( .A1(n21669), .A2(n21778), .ZN(n21641) );
  OR2_X1 U24651 ( .A1(n21637), .A2(n21636), .ZN(n21774) );
  NAND2_X1 U24652 ( .A1(n21774), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n21780) );
  OAI21_X1 U24653 ( .B1(n21704), .B2(n21660), .A(n21780), .ZN(n21638) );
  INV_X1 U24654 ( .A(n21638), .ZN(n21640) );
  INV_X1 U24655 ( .A(n21641), .ZN(n21643) );
  AOI22_X1 U24656 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n21662), .B1(
        n21812), .B2(n21661), .ZN(n21645) );
  OAI211_X1 U24657 ( .C1(n21823), .C2(n21665), .A(n21646), .B(n21645), .ZN(
        P1_U3113) );
  AOI22_X1 U24658 ( .A1(n21655), .A2(n21740), .B1(n21824), .B2(n21660), .ZN(
        n21648) );
  AOI22_X1 U24659 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n21662), .B1(
        n21825), .B2(n21661), .ZN(n21647) );
  OAI211_X1 U24660 ( .C1(n21743), .C2(n21696), .A(n21648), .B(n21647), .ZN(
        P1_U3114) );
  AOI22_X1 U24661 ( .A1(n21655), .A2(n21744), .B1(n21830), .B2(n21660), .ZN(
        n21650) );
  AOI22_X1 U24662 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n21662), .B1(
        n21831), .B2(n21661), .ZN(n21649) );
  OAI211_X1 U24663 ( .C1(n21747), .C2(n21696), .A(n21650), .B(n21649), .ZN(
        P1_U3115) );
  AOI22_X1 U24664 ( .A1(n21687), .A2(n21838), .B1(n21836), .B2(n21660), .ZN(
        n21652) );
  AOI22_X1 U24665 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n21662), .B1(
        n21837), .B2(n21661), .ZN(n21651) );
  OAI211_X1 U24666 ( .C1(n21841), .C2(n21665), .A(n21652), .B(n21651), .ZN(
        P1_U3116) );
  AOI22_X1 U24667 ( .A1(n21687), .A2(n21844), .B1(n21842), .B2(n21660), .ZN(
        n21654) );
  AOI22_X1 U24668 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n21662), .B1(
        n21843), .B2(n21661), .ZN(n21653) );
  OAI211_X1 U24669 ( .C1(n21847), .C2(n21665), .A(n21654), .B(n21653), .ZN(
        P1_U3117) );
  AOI22_X1 U24670 ( .A1(n21655), .A2(n21756), .B1(n21848), .B2(n21660), .ZN(
        n21657) );
  AOI22_X1 U24671 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n21662), .B1(
        n21849), .B2(n21661), .ZN(n21656) );
  OAI211_X1 U24672 ( .C1(n21759), .C2(n21696), .A(n21657), .B(n21656), .ZN(
        P1_U3118) );
  AOI22_X1 U24673 ( .A1(n21687), .A2(n21856), .B1(n21854), .B2(n21660), .ZN(
        n21659) );
  AOI22_X1 U24674 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n21662), .B1(
        n21855), .B2(n21661), .ZN(n21658) );
  OAI211_X1 U24675 ( .C1(n21859), .C2(n21665), .A(n21659), .B(n21658), .ZN(
        P1_U3119) );
  AOI22_X1 U24676 ( .A1(n21687), .A2(n21864), .B1(n21861), .B2(n21660), .ZN(
        n21664) );
  AOI22_X1 U24677 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n21662), .B1(
        n21863), .B2(n21661), .ZN(n21663) );
  OAI211_X1 U24678 ( .C1(n21870), .C2(n21665), .A(n21664), .B(n21663), .ZN(
        P1_U3120) );
  NOR2_X1 U24679 ( .A1(n21804), .A2(n21668), .ZN(n21690) );
  AOI21_X1 U24680 ( .B1(n21669), .B2(n21805), .A(n21690), .ZN(n21671) );
  OAI22_X1 U24681 ( .A1(n21671), .A2(n21810), .B1(n21670), .B2(n12682), .ZN(
        n21691) );
  AOI22_X1 U24682 ( .A1(n21812), .A2(n21691), .B1(n21811), .B2(n21690), .ZN(
        n21676) );
  OAI21_X1 U24683 ( .B1(n21815), .B2(n21672), .A(n21671), .ZN(n21673) );
  OAI211_X1 U24684 ( .C1(n21819), .C2(n21674), .A(n21817), .B(n21673), .ZN(
        n21693) );
  AOI22_X1 U24685 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n21693), .B1(
        n21687), .B2(n21736), .ZN(n21675) );
  OAI211_X1 U24686 ( .C1(n21739), .C2(n21727), .A(n21676), .B(n21675), .ZN(
        P1_U3121) );
  AOI22_X1 U24687 ( .A1(n21825), .A2(n21691), .B1(n21824), .B2(n21690), .ZN(
        n21678) );
  INV_X1 U24688 ( .A(n21727), .ZN(n21692) );
  AOI22_X1 U24689 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n21693), .B1(
        n21692), .B2(n21826), .ZN(n21677) );
  OAI211_X1 U24690 ( .C1(n21829), .C2(n21696), .A(n21678), .B(n21677), .ZN(
        P1_U3122) );
  AOI22_X1 U24691 ( .A1(n21831), .A2(n21691), .B1(n21830), .B2(n21690), .ZN(
        n21680) );
  AOI22_X1 U24692 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n21693), .B1(
        n21692), .B2(n21832), .ZN(n21679) );
  OAI211_X1 U24693 ( .C1(n21835), .C2(n21696), .A(n21680), .B(n21679), .ZN(
        P1_U3123) );
  AOI22_X1 U24694 ( .A1(n21837), .A2(n21691), .B1(n21836), .B2(n21690), .ZN(
        n21682) );
  AOI22_X1 U24695 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n21693), .B1(
        n21687), .B2(n21748), .ZN(n21681) );
  OAI211_X1 U24696 ( .C1(n21751), .C2(n21727), .A(n21682), .B(n21681), .ZN(
        P1_U3124) );
  AOI22_X1 U24697 ( .A1(n21843), .A2(n21691), .B1(n21842), .B2(n21690), .ZN(
        n21684) );
  AOI22_X1 U24698 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n21693), .B1(
        n21687), .B2(n21752), .ZN(n21683) );
  OAI211_X1 U24699 ( .C1(n21755), .C2(n21727), .A(n21684), .B(n21683), .ZN(
        P1_U3125) );
  AOI22_X1 U24700 ( .A1(n21849), .A2(n21691), .B1(n21848), .B2(n21690), .ZN(
        n21686) );
  AOI22_X1 U24701 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n21693), .B1(
        n21692), .B2(n21850), .ZN(n21685) );
  OAI211_X1 U24702 ( .C1(n21853), .C2(n21696), .A(n21686), .B(n21685), .ZN(
        P1_U3126) );
  AOI22_X1 U24703 ( .A1(n21855), .A2(n21691), .B1(n21854), .B2(n21690), .ZN(
        n21689) );
  AOI22_X1 U24704 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n21693), .B1(
        n21687), .B2(n21760), .ZN(n21688) );
  OAI211_X1 U24705 ( .C1(n21763), .C2(n21727), .A(n21689), .B(n21688), .ZN(
        P1_U3127) );
  AOI22_X1 U24706 ( .A1(n21863), .A2(n21691), .B1(n21861), .B2(n21690), .ZN(
        n21695) );
  AOI22_X1 U24707 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n21693), .B1(
        n21692), .B2(n21864), .ZN(n21694) );
  OAI211_X1 U24708 ( .C1(n21870), .C2(n21696), .A(n21695), .B(n21694), .ZN(
        P1_U3128) );
  NAND2_X1 U24709 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n21807) );
  AOI22_X1 U24710 ( .A1(n21767), .A2(n21820), .B1(n21811), .B2(n10675), .ZN(
        n21710) );
  NAND2_X1 U24711 ( .A1(n21727), .A2(n21819), .ZN(n21700) );
  OAI21_X1 U24712 ( .B1(n21700), .B2(n21767), .A(n21699), .ZN(n21705) );
  NAND2_X1 U24713 ( .A1(n21806), .A2(n21702), .ZN(n21707) );
  AOI22_X1 U24714 ( .A1(n21705), .A2(n21707), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n21706), .ZN(n21703) );
  INV_X1 U24715 ( .A(n21705), .ZN(n21708) );
  AOI22_X1 U24716 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n21724), .B1(
        n21812), .B2(n21723), .ZN(n21709) );
  OAI211_X1 U24717 ( .C1(n21823), .C2(n21727), .A(n21710), .B(n21709), .ZN(
        P1_U3129) );
  AOI22_X1 U24718 ( .A1(n21767), .A2(n21826), .B1(n21824), .B2(n10675), .ZN(
        n21712) );
  AOI22_X1 U24719 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n21724), .B1(
        n21825), .B2(n21723), .ZN(n21711) );
  OAI211_X1 U24720 ( .C1(n21829), .C2(n21727), .A(n21712), .B(n21711), .ZN(
        P1_U3130) );
  AOI22_X1 U24721 ( .A1(n21767), .A2(n21832), .B1(n21830), .B2(n10675), .ZN(
        n21714) );
  AOI22_X1 U24722 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n21724), .B1(
        n21831), .B2(n21723), .ZN(n21713) );
  OAI211_X1 U24723 ( .C1(n21835), .C2(n21727), .A(n21714), .B(n21713), .ZN(
        P1_U3131) );
  AOI22_X1 U24724 ( .A1(n21767), .A2(n21838), .B1(n21836), .B2(n10675), .ZN(
        n21716) );
  AOI22_X1 U24725 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n21724), .B1(
        n21837), .B2(n21723), .ZN(n21715) );
  OAI211_X1 U24726 ( .C1(n21841), .C2(n21727), .A(n21716), .B(n21715), .ZN(
        P1_U3132) );
  AOI22_X1 U24727 ( .A1(n21767), .A2(n21844), .B1(n21842), .B2(n10675), .ZN(
        n21718) );
  AOI22_X1 U24728 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n21724), .B1(
        n21843), .B2(n21723), .ZN(n21717) );
  OAI211_X1 U24729 ( .C1(n21847), .C2(n21727), .A(n21718), .B(n21717), .ZN(
        P1_U3133) );
  AOI22_X1 U24730 ( .A1(n21767), .A2(n21850), .B1(n21848), .B2(n10675), .ZN(
        n21720) );
  AOI22_X1 U24731 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n21724), .B1(
        n21849), .B2(n21723), .ZN(n21719) );
  OAI211_X1 U24732 ( .C1(n21853), .C2(n21727), .A(n21720), .B(n21719), .ZN(
        P1_U3134) );
  AOI22_X1 U24733 ( .A1(n21767), .A2(n21856), .B1(n21854), .B2(n10675), .ZN(
        n21722) );
  AOI22_X1 U24734 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n21724), .B1(
        n21855), .B2(n21723), .ZN(n21721) );
  OAI211_X1 U24735 ( .C1(n21859), .C2(n21727), .A(n21722), .B(n21721), .ZN(
        P1_U3135) );
  AOI22_X1 U24736 ( .A1(n21767), .A2(n21864), .B1(n21861), .B2(n10675), .ZN(
        n21726) );
  AOI22_X1 U24737 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n21724), .B1(
        n21863), .B2(n21723), .ZN(n21725) );
  OAI211_X1 U24738 ( .C1(n21870), .C2(n21727), .A(n21726), .B(n21725), .ZN(
        P1_U3136) );
  NOR3_X2 U24739 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n21729), .A3(
        n21807), .ZN(n21764) );
  AOI21_X1 U24740 ( .B1(n21806), .B2(n21730), .A(n21764), .ZN(n21732) );
  NOR2_X1 U24741 ( .A1(n21807), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n21735) );
  INV_X1 U24742 ( .A(n21735), .ZN(n21731) );
  OAI22_X1 U24743 ( .A1(n21732), .A2(n21810), .B1(n21731), .B2(n12682), .ZN(
        n21765) );
  AOI22_X1 U24744 ( .A1(n21812), .A2(n21765), .B1(n21811), .B2(n21764), .ZN(
        n21738) );
  NOR2_X1 U24745 ( .A1(n21776), .A2(n21810), .ZN(n21814) );
  OAI21_X1 U24746 ( .B1(n21814), .B2(n21733), .A(n21732), .ZN(n21734) );
  OAI211_X1 U24747 ( .C1(n21819), .C2(n21735), .A(n21817), .B(n21734), .ZN(
        n21768) );
  AOI22_X1 U24748 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n21768), .B1(
        n21767), .B2(n21736), .ZN(n21737) );
  OAI211_X1 U24749 ( .C1(n21739), .C2(n21803), .A(n21738), .B(n21737), .ZN(
        P1_U3137) );
  AOI22_X1 U24750 ( .A1(n21825), .A2(n21765), .B1(n21824), .B2(n21764), .ZN(
        n21742) );
  AOI22_X1 U24751 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n21768), .B1(
        n21767), .B2(n21740), .ZN(n21741) );
  OAI211_X1 U24752 ( .C1(n21743), .C2(n21803), .A(n21742), .B(n21741), .ZN(
        P1_U3138) );
  AOI22_X1 U24753 ( .A1(n21831), .A2(n21765), .B1(n21830), .B2(n21764), .ZN(
        n21746) );
  AOI22_X1 U24754 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n21768), .B1(
        n21767), .B2(n21744), .ZN(n21745) );
  OAI211_X1 U24755 ( .C1(n21747), .C2(n21803), .A(n21746), .B(n21745), .ZN(
        P1_U3139) );
  AOI22_X1 U24756 ( .A1(n21837), .A2(n21765), .B1(n21836), .B2(n21764), .ZN(
        n21750) );
  AOI22_X1 U24757 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n21768), .B1(
        n21767), .B2(n21748), .ZN(n21749) );
  OAI211_X1 U24758 ( .C1(n21751), .C2(n21803), .A(n21750), .B(n21749), .ZN(
        P1_U3140) );
  AOI22_X1 U24759 ( .A1(n21843), .A2(n21765), .B1(n21842), .B2(n21764), .ZN(
        n21754) );
  AOI22_X1 U24760 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n21768), .B1(
        n21767), .B2(n21752), .ZN(n21753) );
  OAI211_X1 U24761 ( .C1(n21755), .C2(n21803), .A(n21754), .B(n21753), .ZN(
        P1_U3141) );
  AOI22_X1 U24762 ( .A1(n21849), .A2(n21765), .B1(n21848), .B2(n21764), .ZN(
        n21758) );
  AOI22_X1 U24763 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n21768), .B1(
        n21767), .B2(n21756), .ZN(n21757) );
  OAI211_X1 U24764 ( .C1(n21759), .C2(n21803), .A(n21758), .B(n21757), .ZN(
        P1_U3142) );
  AOI22_X1 U24765 ( .A1(n21855), .A2(n21765), .B1(n21854), .B2(n21764), .ZN(
        n21762) );
  AOI22_X1 U24766 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n21768), .B1(
        n21767), .B2(n21760), .ZN(n21761) );
  OAI211_X1 U24767 ( .C1(n21763), .C2(n21803), .A(n21762), .B(n21761), .ZN(
        P1_U3143) );
  AOI22_X1 U24768 ( .A1(n21863), .A2(n21765), .B1(n21861), .B2(n21764), .ZN(
        n21770) );
  AOI22_X1 U24769 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n21768), .B1(
        n21767), .B2(n21766), .ZN(n21769) );
  OAI211_X1 U24770 ( .C1(n21771), .C2(n21803), .A(n21770), .B(n21769), .ZN(
        P1_U3144) );
  NAND3_X1 U24771 ( .A1(n21806), .A2(n21778), .A3(n21819), .ZN(n21772) );
  NOR3_X2 U24772 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21808), .A3(
        n21807), .ZN(n21797) );
  AOI22_X1 U24773 ( .A1(n21812), .A2(n21798), .B1(n21811), .B2(n21797), .ZN(
        n21784) );
  AOI21_X1 U24774 ( .B1(n21869), .B2(n21803), .A(n21905), .ZN(n21777) );
  AOI21_X1 U24775 ( .B1(n21806), .B2(n21778), .A(n21777), .ZN(n21779) );
  NOR2_X1 U24776 ( .A1(n21779), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n21782) );
  AOI22_X1 U24777 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n21800), .B1(
        n21799), .B2(n21820), .ZN(n21783) );
  OAI211_X1 U24778 ( .C1(n21823), .C2(n21803), .A(n21784), .B(n21783), .ZN(
        P1_U3145) );
  AOI22_X1 U24779 ( .A1(n21825), .A2(n21798), .B1(n21824), .B2(n21797), .ZN(
        n21786) );
  AOI22_X1 U24780 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n21800), .B1(
        n21799), .B2(n21826), .ZN(n21785) );
  OAI211_X1 U24781 ( .C1(n21829), .C2(n21803), .A(n21786), .B(n21785), .ZN(
        P1_U3146) );
  AOI22_X1 U24782 ( .A1(n21831), .A2(n21798), .B1(n21830), .B2(n21797), .ZN(
        n21788) );
  AOI22_X1 U24783 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n21800), .B1(
        n21799), .B2(n21832), .ZN(n21787) );
  OAI211_X1 U24784 ( .C1(n21835), .C2(n21803), .A(n21788), .B(n21787), .ZN(
        P1_U3147) );
  AOI22_X1 U24785 ( .A1(n21837), .A2(n21798), .B1(n21836), .B2(n21797), .ZN(
        n21790) );
  AOI22_X1 U24786 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n21800), .B1(
        n21799), .B2(n21838), .ZN(n21789) );
  OAI211_X1 U24787 ( .C1(n21841), .C2(n21803), .A(n21790), .B(n21789), .ZN(
        P1_U3148) );
  AOI22_X1 U24788 ( .A1(n21843), .A2(n21798), .B1(n21842), .B2(n21797), .ZN(
        n21792) );
  AOI22_X1 U24789 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n21800), .B1(
        n21799), .B2(n21844), .ZN(n21791) );
  OAI211_X1 U24790 ( .C1(n21847), .C2(n21803), .A(n21792), .B(n21791), .ZN(
        P1_U3149) );
  AOI22_X1 U24791 ( .A1(n21849), .A2(n21798), .B1(n21848), .B2(n21797), .ZN(
        n21794) );
  AOI22_X1 U24792 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n21800), .B1(
        n21799), .B2(n21850), .ZN(n21793) );
  OAI211_X1 U24793 ( .C1(n21853), .C2(n21803), .A(n21794), .B(n21793), .ZN(
        P1_U3150) );
  AOI22_X1 U24794 ( .A1(n21855), .A2(n21798), .B1(n21854), .B2(n21797), .ZN(
        n21796) );
  AOI22_X1 U24795 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n21800), .B1(
        n21799), .B2(n21856), .ZN(n21795) );
  OAI211_X1 U24796 ( .C1(n21859), .C2(n21803), .A(n21796), .B(n21795), .ZN(
        P1_U3151) );
  AOI22_X1 U24797 ( .A1(n21863), .A2(n21798), .B1(n21861), .B2(n21797), .ZN(
        n21802) );
  AOI22_X1 U24798 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n21800), .B1(
        n21799), .B2(n21864), .ZN(n21801) );
  OAI211_X1 U24799 ( .C1(n21870), .C2(n21803), .A(n21802), .B(n21801), .ZN(
        P1_U3152) );
  NOR2_X1 U24800 ( .A1(n21804), .A2(n21807), .ZN(n21860) );
  AOI21_X1 U24801 ( .B1(n21806), .B2(n21805), .A(n21860), .ZN(n21813) );
  NOR2_X1 U24802 ( .A1(n21808), .A2(n21807), .ZN(n21818) );
  INV_X1 U24803 ( .A(n21818), .ZN(n21809) );
  OAI22_X1 U24804 ( .A1(n21813), .A2(n21810), .B1(n21809), .B2(n12682), .ZN(
        n21862) );
  AOI22_X1 U24805 ( .A1(n21812), .A2(n21862), .B1(n21811), .B2(n21860), .ZN(
        n21822) );
  OAI21_X1 U24806 ( .B1(n21815), .B2(n21814), .A(n21813), .ZN(n21816) );
  OAI211_X1 U24807 ( .C1(n21819), .C2(n21818), .A(n21817), .B(n21816), .ZN(
        n21866) );
  AOI22_X1 U24808 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n21866), .B1(
        n21865), .B2(n21820), .ZN(n21821) );
  OAI211_X1 U24809 ( .C1(n21823), .C2(n21869), .A(n21822), .B(n21821), .ZN(
        P1_U3153) );
  AOI22_X1 U24810 ( .A1(n21825), .A2(n21862), .B1(n21824), .B2(n21860), .ZN(
        n21828) );
  AOI22_X1 U24811 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n21866), .B1(
        n21865), .B2(n21826), .ZN(n21827) );
  OAI211_X1 U24812 ( .C1(n21829), .C2(n21869), .A(n21828), .B(n21827), .ZN(
        P1_U3154) );
  AOI22_X1 U24813 ( .A1(n21831), .A2(n21862), .B1(n21830), .B2(n21860), .ZN(
        n21834) );
  AOI22_X1 U24814 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n21866), .B1(
        n21865), .B2(n21832), .ZN(n21833) );
  OAI211_X1 U24815 ( .C1(n21835), .C2(n21869), .A(n21834), .B(n21833), .ZN(
        P1_U3155) );
  AOI22_X1 U24816 ( .A1(n21837), .A2(n21862), .B1(n21836), .B2(n21860), .ZN(
        n21840) );
  AOI22_X1 U24817 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n21866), .B1(
        n21865), .B2(n21838), .ZN(n21839) );
  OAI211_X1 U24818 ( .C1(n21841), .C2(n21869), .A(n21840), .B(n21839), .ZN(
        P1_U3156) );
  AOI22_X1 U24819 ( .A1(n21843), .A2(n21862), .B1(n21842), .B2(n21860), .ZN(
        n21846) );
  AOI22_X1 U24820 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n21866), .B1(
        n21865), .B2(n21844), .ZN(n21845) );
  OAI211_X1 U24821 ( .C1(n21847), .C2(n21869), .A(n21846), .B(n21845), .ZN(
        P1_U3157) );
  AOI22_X1 U24822 ( .A1(n21849), .A2(n21862), .B1(n21848), .B2(n21860), .ZN(
        n21852) );
  AOI22_X1 U24823 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n21866), .B1(
        n21865), .B2(n21850), .ZN(n21851) );
  OAI211_X1 U24824 ( .C1(n21853), .C2(n21869), .A(n21852), .B(n21851), .ZN(
        P1_U3158) );
  AOI22_X1 U24825 ( .A1(n21855), .A2(n21862), .B1(n21854), .B2(n21860), .ZN(
        n21858) );
  AOI22_X1 U24826 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n21866), .B1(
        n21865), .B2(n21856), .ZN(n21857) );
  OAI211_X1 U24827 ( .C1(n21859), .C2(n21869), .A(n21858), .B(n21857), .ZN(
        P1_U3159) );
  AOI22_X1 U24828 ( .A1(n21863), .A2(n21862), .B1(n21861), .B2(n21860), .ZN(
        n21868) );
  AOI22_X1 U24829 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n21866), .B1(
        n21865), .B2(n21864), .ZN(n21867) );
  OAI211_X1 U24830 ( .C1(n21870), .C2(n21869), .A(n21868), .B(n21867), .ZN(
        P1_U3160) );
  NOR2_X1 U24831 ( .A1(n21908), .A2(n21871), .ZN(n21874) );
  INV_X1 U24832 ( .A(n21872), .ZN(n21873) );
  OAI21_X1 U24833 ( .B1(n21874), .B2(n12682), .A(n21873), .ZN(P1_U3163) );
  AND2_X1 U24834 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n21875), .ZN(
        P1_U3164) );
  AND2_X1 U24835 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n21875), .ZN(
        P1_U3165) );
  AND2_X1 U24836 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n21875), .ZN(
        P1_U3166) );
  AND2_X1 U24837 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n21875), .ZN(
        P1_U3167) );
  AND2_X1 U24838 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n21875), .ZN(
        P1_U3168) );
  AND2_X1 U24839 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n21875), .ZN(
        P1_U3169) );
  AND2_X1 U24840 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n21875), .ZN(
        P1_U3170) );
  AND2_X1 U24841 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n21875), .ZN(
        P1_U3171) );
  AND2_X1 U24842 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n21875), .ZN(
        P1_U3172) );
  AND2_X1 U24843 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n21875), .ZN(
        P1_U3173) );
  AND2_X1 U24844 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n21875), .ZN(
        P1_U3174) );
  AND2_X1 U24845 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n21875), .ZN(
        P1_U3175) );
  AND2_X1 U24846 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n21875), .ZN(
        P1_U3176) );
  AND2_X1 U24847 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n21875), .ZN(
        P1_U3177) );
  AND2_X1 U24848 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n21875), .ZN(
        P1_U3178) );
  AND2_X1 U24849 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n21875), .ZN(
        P1_U3179) );
  AND2_X1 U24850 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n21875), .ZN(
        P1_U3180) );
  AND2_X1 U24851 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n21875), .ZN(
        P1_U3181) );
  AND2_X1 U24852 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n21875), .ZN(
        P1_U3182) );
  AND2_X1 U24853 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n21875), .ZN(
        P1_U3183) );
  AND2_X1 U24854 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n21875), .ZN(
        P1_U3184) );
  AND2_X1 U24855 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n21875), .ZN(
        P1_U3185) );
  AND2_X1 U24856 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n21875), .ZN(P1_U3186) );
  AND2_X1 U24857 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n21875), .ZN(P1_U3187) );
  AND2_X1 U24858 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n21875), .ZN(P1_U3188) );
  AND2_X1 U24859 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n21875), .ZN(P1_U3189) );
  AND2_X1 U24860 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n21875), .ZN(P1_U3190) );
  AND2_X1 U24861 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n21875), .ZN(P1_U3191) );
  AND2_X1 U24862 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n21875), .ZN(P1_U3192) );
  AND2_X1 U24863 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n21875), .ZN(P1_U3193) );
  INV_X1 U24864 ( .A(n21876), .ZN(n21886) );
  AOI22_X1 U24865 ( .A1(n21886), .A2(P1_REIP_REG_8__SCAN_IN), .B1(n21916), 
        .B2(P1_ADDRESS_REG_7__SCAN_IN), .ZN(n21877) );
  OAI21_X1 U24866 ( .B1(n21878), .B2(n13610), .A(n21877), .ZN(P1_U3204) );
  AOI22_X1 U24867 ( .A1(n21886), .A2(P1_REIP_REG_12__SCAN_IN), .B1(n21916), 
        .B2(P1_ADDRESS_REG_11__SCAN_IN), .ZN(n21879) );
  OAI21_X1 U24868 ( .B1(n21880), .B2(n13610), .A(n21879), .ZN(P1_U3208) );
  AOI22_X1 U24869 ( .A1(n21886), .A2(P1_REIP_REG_20__SCAN_IN), .B1(n21916), 
        .B2(P1_ADDRESS_REG_19__SCAN_IN), .ZN(n21881) );
  OAI21_X1 U24870 ( .B1(n21882), .B2(n13610), .A(n21881), .ZN(P1_U3216) );
  AOI22_X1 U24871 ( .A1(n21886), .A2(P1_REIP_REG_22__SCAN_IN), .B1(n21916), 
        .B2(P1_ADDRESS_REG_21__SCAN_IN), .ZN(n21883) );
  OAI21_X1 U24872 ( .B1(n21884), .B2(n13610), .A(n21883), .ZN(P1_U3218) );
  AOI22_X1 U24873 ( .A1(n21886), .A2(P1_REIP_REG_24__SCAN_IN), .B1(n21916), 
        .B2(P1_ADDRESS_REG_23__SCAN_IN), .ZN(n21885) );
  OAI21_X1 U24874 ( .B1(n22130), .B2(n13610), .A(n21885), .ZN(P1_U3220) );
  AOI22_X1 U24875 ( .A1(n21886), .A2(P1_REIP_REG_26__SCAN_IN), .B1(n21916), 
        .B2(P1_ADDRESS_REG_25__SCAN_IN), .ZN(n21887) );
  OAI21_X1 U24876 ( .B1(n21888), .B2(n13610), .A(n21887), .ZN(P1_U3222) );
  OAI22_X1 U24877 ( .A1(n21916), .A2(P1_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P1_BE_N_REG_3__SCAN_IN), .B2(n21915), .ZN(n21889) );
  INV_X1 U24878 ( .A(n21889), .ZN(P1_U3458) );
  OAI22_X1 U24879 ( .A1(n21916), .A2(P1_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P1_BE_N_REG_2__SCAN_IN), .B2(n21915), .ZN(n21890) );
  INV_X1 U24880 ( .A(n21890), .ZN(P1_U3459) );
  OAI22_X1 U24881 ( .A1(n21916), .A2(P1_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P1_BE_N_REG_1__SCAN_IN), .B2(n21915), .ZN(n21891) );
  INV_X1 U24882 ( .A(n21891), .ZN(P1_U3460) );
  INV_X1 U24883 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n21901) );
  INV_X1 U24884 ( .A(P1_BE_N_REG_0__SCAN_IN), .ZN(n22022) );
  AOI22_X1 U24885 ( .A1(n21915), .A2(n21901), .B1(n22022), .B2(n21916), .ZN(
        P1_U3461) );
  OAI21_X1 U24886 ( .B1(P1_DATAWIDTH_REG_0__SCAN_IN), .B2(n21895), .A(n21893), 
        .ZN(n21892) );
  INV_X1 U24887 ( .A(n21892), .ZN(P1_U3464) );
  OAI21_X1 U24888 ( .B1(n21895), .B2(n21894), .A(n21893), .ZN(P1_U3465) );
  AOI21_X1 U24889 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n21897) );
  AOI22_X1 U24890 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .B1(n21897), .B2(n21896), .ZN(n21899) );
  INV_X1 U24891 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n21993) );
  AOI22_X1 U24892 ( .A1(n21902), .A2(n21899), .B1(n21993), .B2(n21898), .ZN(
        P1_U3481) );
  OAI21_X1 U24893 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(P1_REIP_REG_0__SCAN_IN), 
        .A(n21902), .ZN(n21900) );
  OAI21_X1 U24894 ( .B1(n21902), .B2(n21901), .A(n21900), .ZN(P1_U3482) );
  INV_X1 U24895 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n21903) );
  AOI22_X1 U24896 ( .A1(n21915), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n21903), 
        .B2(n21916), .ZN(P1_U3483) );
  AOI211_X1 U24897 ( .C1(n21906), .C2(n21905), .A(n12682), .B(n21904), .ZN(
        n21909) );
  OAI21_X1 U24898 ( .B1(n21909), .B2(n21908), .A(n21907), .ZN(n21914) );
  AOI211_X1 U24899 ( .C1(n21299), .C2(n21912), .A(n21911), .B(n21910), .ZN(
        n21913) );
  MUX2_X1 U24900 ( .A(n21914), .B(P1_REQUESTPENDING_REG_SCAN_IN), .S(n21913), 
        .Z(P1_U3485) );
  OAI22_X1 U24901 ( .A1(n21916), .A2(P1_MEMORYFETCH_REG_SCAN_IN), .B1(
        P1_M_IO_N_REG_SCAN_IN), .B2(n21915), .ZN(n21917) );
  INV_X1 U24902 ( .A(n21917), .ZN(P1_U3486) );
  AOI22_X1 U24903 ( .A1(n21921), .A2(n21920), .B1(n21919), .B2(n21918), .ZN(
        n21926) );
  AOI22_X1 U24904 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n21924), .B1(
        n21923), .B2(n21922), .ZN(n21925) );
  OAI211_X1 U24905 ( .C1(n21928), .C2(n21927), .A(n21926), .B(n21925), .ZN(
        n22235) );
  NOR4_X1 U24906 ( .A1(P1_M_IO_N_REG_SCAN_IN), .A2(DATAI_23_), .A3(
        P2_DATAO_REG_0__SCAN_IN), .A4(n22185), .ZN(n21929) );
  NAND3_X1 U24907 ( .A1(P1_ADS_N_REG_SCAN_IN), .A2(n21929), .A3(n22170), .ZN(
        n21939) );
  NAND4_X1 U24908 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(
        P3_EAX_REG_17__SCAN_IN), .A3(n22201), .A4(n22204), .ZN(n21933) );
  NAND4_X1 U24909 ( .A1(P1_EAX_REG_5__SCAN_IN), .A2(BUF2_REG_15__SCAN_IN), 
        .A3(P3_ADDRESS_REG_24__SCAN_IN), .A4(n22194), .ZN(n21932) );
  NAND4_X1 U24910 ( .A1(P1_EAX_REG_13__SCAN_IN), .A2(P2_EAX_REG_10__SCAN_IN), 
        .A3(P3_EBX_REG_23__SCAN_IN), .A4(n22120), .ZN(n21931) );
  NAND4_X1 U24911 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(P1_EBX_REG_25__SCAN_IN), .A4(
        n22114), .ZN(n21930) );
  NOR4_X1 U24912 ( .A1(n21933), .A2(n21932), .A3(n21931), .A4(n21930), .ZN(
        n21937) );
  NAND4_X1 U24913 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_25__SCAN_IN), .A3(n22213), .A4(n22210), .ZN(n21935)
         );
  NAND4_X1 U24914 ( .A1(n22214), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A3(
        P1_INSTQUEUE_REG_3__3__SCAN_IN), .A4(P2_UWORD_REG_4__SCAN_IN), .ZN(
        n21934) );
  NOR2_X1 U24915 ( .A1(n21935), .A2(n21934), .ZN(n21936) );
  NAND2_X1 U24916 ( .A1(n21937), .A2(n21936), .ZN(n21938) );
  NOR4_X1 U24917 ( .A1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A3(n21939), .A4(n21938), .ZN(
        n21974) );
  INV_X1 U24918 ( .A(BS16), .ZN(n22063) );
  NAND4_X1 U24919 ( .A1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(P2_EAX_REG_12__SCAN_IN), .A4(
        n22063), .ZN(n21943) );
  NAND4_X1 U24920 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n22052), .A3(
        n22056), .A4(n22048), .ZN(n21942) );
  NAND4_X1 U24921 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_23__SCAN_IN), .A3(n22088), .A4(n22085), .ZN(n21941)
         );
  NAND4_X1 U24922 ( .A1(DATAI_31_), .A2(P2_DATAWIDTH_REG_19__SCAN_IN), .A3(
        P3_LWORD_REG_7__SCAN_IN), .A4(n22079), .ZN(n21940) );
  NOR4_X1 U24923 ( .A1(n21943), .A2(n21942), .A3(n21941), .A4(n21940), .ZN(
        n21973) );
  NAND4_X1 U24924 ( .A1(P3_BYTEENABLE_REG_0__SCAN_IN), .A2(
        P1_BE_N_REG_0__SCAN_IN), .A3(n13609), .A4(n22023), .ZN(n21947) );
  INV_X1 U24925 ( .A(DATAI_28_), .ZN(n22005) );
  NAND4_X1 U24926 ( .A1(P1_LWORD_REG_11__SCAN_IN), .A2(n22005), .A3(n10077), 
        .A4(n13665), .ZN(n21946) );
  NAND4_X1 U24927 ( .A1(P3_EAX_REG_27__SCAN_IN), .A2(n22042), .A3(n12212), 
        .A4(n22049), .ZN(n21945) );
  NAND4_X1 U24928 ( .A1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_INSTQUEUE_REG_1__6__SCAN_IN), .A3(n16511), .A4(n15264), .ZN(n21944)
         );
  NOR4_X1 U24929 ( .A1(n21947), .A2(n21946), .A3(n21945), .A4(n21944), .ZN(
        n21972) );
  NOR4_X1 U24930 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_12__2__SCAN_IN), .A3(P2_INSTQUEUE_REG_8__2__SCAN_IN), 
        .A4(n22025), .ZN(n21951) );
  NOR4_X1 U24931 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n10988), .A3(
        n22054), .A4(n14469), .ZN(n21950) );
  NOR4_X1 U24932 ( .A1(P2_REIP_REG_10__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(n22020), .A4(n22186), .ZN(n21949) );
  NOR4_X1 U24933 ( .A1(P2_ADDRESS_REG_14__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .A3(n22183), .A4(n22117), .ZN(
        n21948) );
  NAND4_X1 U24934 ( .A1(n21951), .A2(n21950), .A3(n21949), .A4(n21948), .ZN(
        n21970) );
  NOR2_X1 U24935 ( .A1(n22123), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n21956) );
  NOR4_X1 U24936 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_11__SCAN_IN), .A3(n22087), .A4(n21952), .ZN(n21955)
         );
  INV_X1 U24937 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n22062) );
  NOR4_X1 U24938 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_5__3__SCAN_IN), .A3(P2_INSTQUEUE_REG_12__7__SCAN_IN), 
        .A4(n22062), .ZN(n21954) );
  INV_X1 U24939 ( .A(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n22069) );
  INV_X1 U24940 ( .A(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n21991) );
  NOR4_X1 U24941 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_11__6__SCAN_IN), .A3(n22069), .A4(n21991), .ZN(n21953) );
  NAND4_X1 U24942 ( .A1(n21956), .A2(n21955), .A3(n21954), .A4(n21953), .ZN(
        n21969) );
  NOR4_X1 U24943 ( .A1(BUF1_REG_17__SCAN_IN), .A2(P1_UWORD_REG_8__SCAN_IN), 
        .A3(n21976), .A4(n21977), .ZN(n21962) );
  NOR4_X1 U24944 ( .A1(P1_BYTEENABLE_REG_2__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A3(P3_DATAO_REG_10__SCAN_IN), 
        .A4(n11299), .ZN(n21961) );
  NOR4_X1 U24945 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(
        P3_INSTQUEUE_REG_8__3__SCAN_IN), .A3(n21979), .A4(n21957), .ZN(n21958)
         );
  AND4_X1 U24946 ( .A1(n21959), .A2(P1_STATE_REG_1__SCAN_IN), .A3(n21958), 
        .A4(BUF2_REG_0__SCAN_IN), .ZN(n21960) );
  NAND4_X1 U24947 ( .A1(n21962), .A2(n21961), .A3(n21960), .A4(
        P3_ADDRESS_REG_5__SCAN_IN), .ZN(n21968) );
  NOR4_X1 U24948 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(
        P3_ADDRESS_REG_19__SCAN_IN), .A3(n22149), .A4(n22146), .ZN(n21966) );
  NOR4_X1 U24949 ( .A1(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTQUEUE_REG_13__2__SCAN_IN), .A3(P3_EAX_REG_12__SCAN_IN), .A4(
        n22104), .ZN(n21965) );
  NOR4_X1 U24950 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(
        P3_INSTQUEUE_REG_9__2__SCAN_IN), .A3(n21982), .A4(n22140), .ZN(n21964)
         );
  NOR4_X1 U24951 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n22151), .A3(n22154), 
        .A4(n22132), .ZN(n21963) );
  NAND4_X1 U24952 ( .A1(n21966), .A2(n21965), .A3(n21964), .A4(n21963), .ZN(
        n21967) );
  NOR4_X1 U24953 ( .A1(n21970), .A2(n21969), .A3(n21968), .A4(n21967), .ZN(
        n21971) );
  NAND4_X1 U24954 ( .A1(n21974), .A2(n21973), .A3(n21972), .A4(n21971), .ZN(
        n22232) );
  AOI22_X1 U24955 ( .A1(n21977), .A2(keyinput30), .B1(keyinput75), .B2(n21976), 
        .ZN(n21975) );
  OAI221_X1 U24956 ( .B1(n21977), .B2(keyinput30), .C1(n21976), .C2(keyinput75), .A(n21975), .ZN(n21989) );
  AOI22_X1 U24957 ( .A1(n21980), .A2(keyinput35), .B1(n21979), .B2(keyinput109), .ZN(n21978) );
  OAI221_X1 U24958 ( .B1(n21980), .B2(keyinput35), .C1(n21979), .C2(
        keyinput109), .A(n21978), .ZN(n21988) );
  INV_X1 U24959 ( .A(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n21983) );
  AOI22_X1 U24960 ( .A1(n21983), .A2(keyinput18), .B1(keyinput23), .B2(n21982), 
        .ZN(n21981) );
  OAI221_X1 U24961 ( .B1(n21983), .B2(keyinput18), .C1(n21982), .C2(keyinput23), .A(n21981), .ZN(n21987) );
  XNOR2_X1 U24962 ( .A(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B(keyinput95), .ZN(
        n21985) );
  XNOR2_X1 U24963 ( .A(keyinput54), .B(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n21984) );
  NAND2_X1 U24964 ( .A1(n21985), .A2(n21984), .ZN(n21986) );
  NOR4_X1 U24965 ( .A1(n21989), .A2(n21988), .A3(n21987), .A4(n21986), .ZN(
        n22034) );
  AOI22_X1 U24966 ( .A1(n16479), .A2(keyinput119), .B1(n21991), .B2(keyinput46), .ZN(n21990) );
  OAI221_X1 U24967 ( .B1(n16479), .B2(keyinput119), .C1(n21991), .C2(
        keyinput46), .A(n21990), .ZN(n22002) );
  AOI22_X1 U24968 ( .A1(n21994), .A2(keyinput69), .B1(keyinput43), .B2(n21993), 
        .ZN(n21992) );
  OAI221_X1 U24969 ( .B1(n21994), .B2(keyinput69), .C1(n21993), .C2(keyinput43), .A(n21992), .ZN(n22001) );
  INV_X1 U24970 ( .A(P3_DATAO_REG_10__SCAN_IN), .ZN(n21996) );
  AOI22_X1 U24971 ( .A1(n15485), .A2(keyinput6), .B1(keyinput121), .B2(n21996), 
        .ZN(n21995) );
  OAI221_X1 U24972 ( .B1(n15485), .B2(keyinput6), .C1(n21996), .C2(keyinput121), .A(n21995), .ZN(n22000) );
  INV_X1 U24973 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n21998) );
  AOI22_X1 U24974 ( .A1(n11299), .A2(keyinput70), .B1(n21998), .B2(keyinput3), 
        .ZN(n21997) );
  OAI221_X1 U24975 ( .B1(n11299), .B2(keyinput70), .C1(n21998), .C2(keyinput3), 
        .A(n21997), .ZN(n21999) );
  NOR4_X1 U24976 ( .A1(n22002), .A2(n22001), .A3(n22000), .A4(n21999), .ZN(
        n22033) );
  AOI22_X1 U24977 ( .A1(n22005), .A2(keyinput5), .B1(keyinput92), .B2(n22004), 
        .ZN(n22003) );
  OAI221_X1 U24978 ( .B1(n22005), .B2(keyinput5), .C1(n22004), .C2(keyinput92), 
        .A(n22003), .ZN(n22009) );
  XOR2_X1 U24979 ( .A(P1_STATE_REG_1__SCAN_IN), .B(keyinput50), .Z(n22008) );
  XNOR2_X1 U24980 ( .A(n22006), .B(keyinput55), .ZN(n22007) );
  OR3_X1 U24981 ( .A1(n22009), .A2(n22008), .A3(n22007), .ZN(n22015) );
  AOI22_X1 U24982 ( .A1(n21959), .A2(keyinput80), .B1(keyinput65), .B2(n22011), 
        .ZN(n22010) );
  OAI221_X1 U24983 ( .B1(n21959), .B2(keyinput80), .C1(n22011), .C2(keyinput65), .A(n22010), .ZN(n22014) );
  AOI22_X1 U24984 ( .A1(n10077), .A2(keyinput42), .B1(keyinput56), .B2(n13665), 
        .ZN(n22012) );
  OAI221_X1 U24985 ( .B1(n10077), .B2(keyinput42), .C1(n13665), .C2(keyinput56), .A(n22012), .ZN(n22013) );
  NOR3_X1 U24986 ( .A1(n22015), .A2(n22014), .A3(n22013), .ZN(n22032) );
  INV_X1 U24987 ( .A(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n22018) );
  AOI22_X1 U24988 ( .A1(n22018), .A2(keyinput21), .B1(keyinput19), .B2(n22017), 
        .ZN(n22016) );
  OAI221_X1 U24989 ( .B1(n22018), .B2(keyinput21), .C1(n22017), .C2(keyinput19), .A(n22016), .ZN(n22030) );
  AOI22_X1 U24990 ( .A1(n22020), .A2(keyinput104), .B1(keyinput106), .B2(
        n13609), .ZN(n22019) );
  OAI221_X1 U24991 ( .B1(n22020), .B2(keyinput104), .C1(n13609), .C2(
        keyinput106), .A(n22019), .ZN(n22029) );
  AOI22_X1 U24992 ( .A1(n22023), .A2(keyinput90), .B1(keyinput118), .B2(n22022), .ZN(n22021) );
  OAI221_X1 U24993 ( .B1(n22023), .B2(keyinput90), .C1(n22022), .C2(
        keyinput118), .A(n22021), .ZN(n22028) );
  AOI22_X1 U24994 ( .A1(n22026), .A2(keyinput59), .B1(n22025), .B2(keyinput102), .ZN(n22024) );
  OAI221_X1 U24995 ( .B1(n22026), .B2(keyinput59), .C1(n22025), .C2(
        keyinput102), .A(n22024), .ZN(n22027) );
  NOR4_X1 U24996 ( .A1(n22030), .A2(n22029), .A3(n22028), .A4(n22027), .ZN(
        n22031) );
  NAND4_X1 U24997 ( .A1(n22034), .A2(n22033), .A3(n22032), .A4(n22031), .ZN(
        n22230) );
  AOI22_X1 U24998 ( .A1(n11738), .A2(keyinput116), .B1(keyinput82), .B2(n22036), .ZN(n22035) );
  OAI221_X1 U24999 ( .B1(n11738), .B2(keyinput116), .C1(n22036), .C2(
        keyinput82), .A(n22035), .ZN(n22046) );
  AOI22_X1 U25000 ( .A1(n16511), .A2(keyinput61), .B1(keyinput49), .B2(n15264), 
        .ZN(n22037) );
  OAI221_X1 U25001 ( .B1(n16511), .B2(keyinput61), .C1(n15264), .C2(keyinput49), .A(n22037), .ZN(n22045) );
  INV_X1 U25002 ( .A(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n22039) );
  AOI22_X1 U25003 ( .A1(n22039), .A2(keyinput107), .B1(keyinput84), .B2(n12212), .ZN(n22038) );
  OAI221_X1 U25004 ( .B1(n22039), .B2(keyinput107), .C1(n12212), .C2(
        keyinput84), .A(n22038), .ZN(n22044) );
  AOI22_X1 U25005 ( .A1(n22042), .A2(keyinput37), .B1(keyinput89), .B2(n22041), 
        .ZN(n22040) );
  OAI221_X1 U25006 ( .B1(n22042), .B2(keyinput37), .C1(n22041), .C2(keyinput89), .A(n22040), .ZN(n22043) );
  NOR4_X1 U25007 ( .A1(n22046), .A2(n22045), .A3(n22044), .A4(n22043), .ZN(
        n22096) );
  AOI22_X1 U25008 ( .A1(n22049), .A2(keyinput1), .B1(keyinput22), .B2(n22048), 
        .ZN(n22047) );
  OAI221_X1 U25009 ( .B1(n22049), .B2(keyinput1), .C1(n22048), .C2(keyinput22), 
        .A(n22047), .ZN(n22060) );
  INV_X1 U25010 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n22051) );
  AOI22_X1 U25011 ( .A1(n22052), .A2(keyinput44), .B1(n22051), .B2(keyinput33), 
        .ZN(n22050) );
  OAI221_X1 U25012 ( .B1(n22052), .B2(keyinput44), .C1(n22051), .C2(keyinput33), .A(n22050), .ZN(n22059) );
  AOI22_X1 U25013 ( .A1(n13270), .A2(keyinput41), .B1(n22054), .B2(keyinput16), 
        .ZN(n22053) );
  OAI221_X1 U25014 ( .B1(n13270), .B2(keyinput41), .C1(n22054), .C2(keyinput16), .A(n22053), .ZN(n22058) );
  AOI22_X1 U25015 ( .A1(n22056), .A2(keyinput87), .B1(n14469), .B2(keyinput68), 
        .ZN(n22055) );
  OAI221_X1 U25016 ( .B1(n22056), .B2(keyinput87), .C1(n14469), .C2(keyinput68), .A(n22055), .ZN(n22057) );
  NOR4_X1 U25017 ( .A1(n22060), .A2(n22059), .A3(n22058), .A4(n22057), .ZN(
        n22095) );
  AOI22_X1 U25018 ( .A1(n22063), .A2(keyinput124), .B1(n22062), .B2(keyinput2), 
        .ZN(n22061) );
  OAI221_X1 U25019 ( .B1(n22063), .B2(keyinput124), .C1(n22062), .C2(keyinput2), .A(n22061), .ZN(n22076) );
  AOI22_X1 U25020 ( .A1(n22066), .A2(keyinput100), .B1(n22065), .B2(
        keyinput122), .ZN(n22064) );
  OAI221_X1 U25021 ( .B1(n22066), .B2(keyinput100), .C1(n22065), .C2(
        keyinput122), .A(n22064), .ZN(n22075) );
  INV_X1 U25022 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n22068) );
  AOI22_X1 U25023 ( .A1(n22069), .A2(keyinput71), .B1(keyinput83), .B2(n22068), 
        .ZN(n22067) );
  OAI221_X1 U25024 ( .B1(n22069), .B2(keyinput71), .C1(n22068), .C2(keyinput83), .A(n22067), .ZN(n22074) );
  AOI22_X1 U25025 ( .A1(n22072), .A2(keyinput36), .B1(keyinput31), .B2(n22071), 
        .ZN(n22070) );
  OAI221_X1 U25026 ( .B1(n22072), .B2(keyinput36), .C1(n22071), .C2(keyinput31), .A(n22070), .ZN(n22073) );
  NOR4_X1 U25027 ( .A1(n22076), .A2(n22075), .A3(n22074), .A4(n22073), .ZN(
        n22094) );
  INV_X1 U25028 ( .A(DATAI_31_), .ZN(n22078) );
  AOI22_X1 U25029 ( .A1(n22079), .A2(keyinput108), .B1(n22078), .B2(keyinput10), .ZN(n22077) );
  OAI221_X1 U25030 ( .B1(n22079), .B2(keyinput108), .C1(n22078), .C2(
        keyinput10), .A(n22077), .ZN(n22092) );
  AOI22_X1 U25031 ( .A1(n22082), .A2(keyinput97), .B1(keyinput7), .B2(n22081), 
        .ZN(n22080) );
  OAI221_X1 U25032 ( .B1(n22082), .B2(keyinput97), .C1(n22081), .C2(keyinput7), 
        .A(n22080), .ZN(n22091) );
  AOI22_X1 U25033 ( .A1(n22085), .A2(keyinput117), .B1(n22084), .B2(keyinput98), .ZN(n22083) );
  OAI221_X1 U25034 ( .B1(n22085), .B2(keyinput117), .C1(n22084), .C2(
        keyinput98), .A(n22083), .ZN(n22090) );
  AOI22_X1 U25035 ( .A1(n22088), .A2(keyinput110), .B1(keyinput91), .B2(n22087), .ZN(n22086) );
  OAI221_X1 U25036 ( .B1(n22088), .B2(keyinput110), .C1(n22087), .C2(
        keyinput91), .A(n22086), .ZN(n22089) );
  NOR4_X1 U25037 ( .A1(n22092), .A2(n22091), .A3(n22090), .A4(n22089), .ZN(
        n22093) );
  NAND4_X1 U25038 ( .A1(n22096), .A2(n22095), .A3(n22094), .A4(n22093), .ZN(
        n22229) );
  AOI22_X1 U25039 ( .A1(n22099), .A2(keyinput26), .B1(keyinput96), .B2(n22098), 
        .ZN(n22097) );
  OAI221_X1 U25040 ( .B1(n22099), .B2(keyinput26), .C1(n22098), .C2(keyinput96), .A(n22097), .ZN(n22112) );
  AOI22_X1 U25041 ( .A1(n22102), .A2(keyinput11), .B1(keyinput105), .B2(n22101), .ZN(n22100) );
  OAI221_X1 U25042 ( .B1(n22102), .B2(keyinput11), .C1(n22101), .C2(
        keyinput105), .A(n22100), .ZN(n22111) );
  AOI22_X1 U25043 ( .A1(n22105), .A2(keyinput72), .B1(keyinput86), .B2(n22104), 
        .ZN(n22103) );
  OAI221_X1 U25044 ( .B1(n22105), .B2(keyinput72), .C1(n22104), .C2(keyinput86), .A(n22103), .ZN(n22110) );
  AOI22_X1 U25045 ( .A1(n22108), .A2(keyinput40), .B1(n22107), .B2(keyinput85), 
        .ZN(n22106) );
  OAI221_X1 U25046 ( .B1(n22108), .B2(keyinput40), .C1(n22107), .C2(keyinput85), .A(n22106), .ZN(n22109) );
  NOR4_X1 U25047 ( .A1(n22112), .A2(n22111), .A3(n22110), .A4(n22109), .ZN(
        n22163) );
  INV_X1 U25048 ( .A(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n22115) );
  AOI22_X1 U25049 ( .A1(n22115), .A2(keyinput74), .B1(keyinput76), .B2(n22114), 
        .ZN(n22113) );
  OAI221_X1 U25050 ( .B1(n22115), .B2(keyinput74), .C1(n22114), .C2(keyinput76), .A(n22113), .ZN(n22128) );
  AOI22_X1 U25051 ( .A1(n22118), .A2(keyinput39), .B1(keyinput77), .B2(n22117), 
        .ZN(n22116) );
  OAI221_X1 U25052 ( .B1(n22118), .B2(keyinput39), .C1(n22117), .C2(keyinput77), .A(n22116), .ZN(n22127) );
  AOI22_X1 U25053 ( .A1(n22121), .A2(keyinput58), .B1(keyinput38), .B2(n22120), 
        .ZN(n22119) );
  OAI221_X1 U25054 ( .B1(n22121), .B2(keyinput58), .C1(n22120), .C2(keyinput38), .A(n22119), .ZN(n22126) );
  INV_X1 U25055 ( .A(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n22124) );
  AOI22_X1 U25056 ( .A1(n22124), .A2(keyinput111), .B1(keyinput67), .B2(n22123), .ZN(n22122) );
  OAI221_X1 U25057 ( .B1(n22124), .B2(keyinput111), .C1(n22123), .C2(
        keyinput67), .A(n22122), .ZN(n22125) );
  NOR4_X1 U25058 ( .A1(n22128), .A2(n22127), .A3(n22126), .A4(n22125), .ZN(
        n22162) );
  INV_X1 U25059 ( .A(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n22131) );
  AOI22_X1 U25060 ( .A1(n22131), .A2(keyinput73), .B1(keyinput63), .B2(n22130), 
        .ZN(n22129) );
  OAI221_X1 U25061 ( .B1(n22131), .B2(keyinput73), .C1(n22130), .C2(keyinput63), .A(n22129), .ZN(n22135) );
  XNOR2_X1 U25062 ( .A(n22132), .B(keyinput24), .ZN(n22134) );
  XOR2_X1 U25063 ( .A(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B(keyinput103), .Z(
        n22133) );
  OR3_X1 U25064 ( .A1(n22135), .A2(n22134), .A3(n22133), .ZN(n22143) );
  AOI22_X1 U25065 ( .A1(n10988), .A2(keyinput88), .B1(keyinput57), .B2(n22137), 
        .ZN(n22136) );
  OAI221_X1 U25066 ( .B1(n10988), .B2(keyinput88), .C1(n22137), .C2(keyinput57), .A(n22136), .ZN(n22142) );
  AOI22_X1 U25067 ( .A1(n22140), .A2(keyinput101), .B1(keyinput126), .B2(
        n22139), .ZN(n22138) );
  OAI221_X1 U25068 ( .B1(n22140), .B2(keyinput101), .C1(n22139), .C2(
        keyinput126), .A(n22138), .ZN(n22141) );
  NOR3_X1 U25069 ( .A1(n22143), .A2(n22142), .A3(n22141), .ZN(n22161) );
  AOI22_X1 U25070 ( .A1(n22146), .A2(keyinput17), .B1(n22145), .B2(keyinput28), 
        .ZN(n22144) );
  OAI221_X1 U25071 ( .B1(n22146), .B2(keyinput17), .C1(n22145), .C2(keyinput28), .A(n22144), .ZN(n22159) );
  AOI22_X1 U25072 ( .A1(n22149), .A2(keyinput53), .B1(n22148), .B2(keyinput81), 
        .ZN(n22147) );
  OAI221_X1 U25073 ( .B1(n22149), .B2(keyinput53), .C1(n22148), .C2(keyinput81), .A(n22147), .ZN(n22158) );
  INV_X1 U25074 ( .A(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n22152) );
  AOI22_X1 U25075 ( .A1(n22152), .A2(keyinput32), .B1(keyinput79), .B2(n22151), 
        .ZN(n22150) );
  OAI221_X1 U25076 ( .B1(n22152), .B2(keyinput32), .C1(n22151), .C2(keyinput79), .A(n22150), .ZN(n22157) );
  AOI22_X1 U25077 ( .A1(n22155), .A2(keyinput12), .B1(n22154), .B2(keyinput125), .ZN(n22153) );
  OAI221_X1 U25078 ( .B1(n22155), .B2(keyinput12), .C1(n22154), .C2(
        keyinput125), .A(n22153), .ZN(n22156) );
  NOR4_X1 U25079 ( .A1(n22159), .A2(n22158), .A3(n22157), .A4(n22156), .ZN(
        n22160) );
  NAND4_X1 U25080 ( .A1(n22163), .A2(n22162), .A3(n22161), .A4(n22160), .ZN(
        n22228) );
  AOI22_X1 U25081 ( .A1(n11761), .A2(keyinput15), .B1(keyinput8), .B2(n22165), 
        .ZN(n22164) );
  OAI221_X1 U25082 ( .B1(n11761), .B2(keyinput15), .C1(n22165), .C2(keyinput8), 
        .A(n22164), .ZN(n22178) );
  AOI22_X1 U25083 ( .A1(n22168), .A2(keyinput120), .B1(keyinput127), .B2(
        n22167), .ZN(n22166) );
  OAI221_X1 U25084 ( .B1(n22168), .B2(keyinput120), .C1(n22167), .C2(
        keyinput127), .A(n22166), .ZN(n22177) );
  AOI22_X1 U25085 ( .A1(n22171), .A2(keyinput94), .B1(n22170), .B2(keyinput113), .ZN(n22169) );
  OAI221_X1 U25086 ( .B1(n22171), .B2(keyinput94), .C1(n22170), .C2(
        keyinput113), .A(n22169), .ZN(n22176) );
  AOI22_X1 U25087 ( .A1(n22174), .A2(keyinput112), .B1(keyinput78), .B2(n22173), .ZN(n22172) );
  OAI221_X1 U25088 ( .B1(n22174), .B2(keyinput112), .C1(n22173), .C2(
        keyinput78), .A(n22172), .ZN(n22175) );
  NOR4_X1 U25089 ( .A1(n22178), .A2(n22177), .A3(n22176), .A4(n22175), .ZN(
        n22226) );
  AOI22_X1 U25090 ( .A1(keyinput115), .A2(n22180), .B1(keyinput14), .B2(n22233), .ZN(n22179) );
  OAI21_X1 U25091 ( .B1(n22180), .B2(keyinput115), .A(n22179), .ZN(n22192) );
  AOI22_X1 U25092 ( .A1(n22183), .A2(keyinput64), .B1(keyinput9), .B2(n22182), 
        .ZN(n22181) );
  OAI221_X1 U25093 ( .B1(n22183), .B2(keyinput64), .C1(n22182), .C2(keyinput9), 
        .A(n22181), .ZN(n22191) );
  AOI22_X1 U25094 ( .A1(n22186), .A2(keyinput45), .B1(n22185), .B2(keyinput27), 
        .ZN(n22184) );
  OAI221_X1 U25095 ( .B1(n22186), .B2(keyinput45), .C1(n22185), .C2(keyinput27), .A(n22184), .ZN(n22190) );
  AOI22_X1 U25096 ( .A1(n22188), .A2(keyinput52), .B1(n11556), .B2(keyinput66), 
        .ZN(n22187) );
  OAI221_X1 U25097 ( .B1(n22188), .B2(keyinput52), .C1(n11556), .C2(keyinput66), .A(n22187), .ZN(n22189) );
  NOR4_X1 U25098 ( .A1(n22192), .A2(n22191), .A3(n22190), .A4(n22189), .ZN(
        n22225) );
  AOI22_X1 U25099 ( .A1(n22195), .A2(keyinput13), .B1(n22194), .B2(keyinput0), 
        .ZN(n22193) );
  OAI221_X1 U25100 ( .B1(n22195), .B2(keyinput13), .C1(n22194), .C2(keyinput0), 
        .A(n22193), .ZN(n22208) );
  AOI22_X1 U25101 ( .A1(n22198), .A2(keyinput25), .B1(n22197), .B2(keyinput20), 
        .ZN(n22196) );
  OAI221_X1 U25102 ( .B1(n22198), .B2(keyinput25), .C1(n22197), .C2(keyinput20), .A(n22196), .ZN(n22207) );
  AOI22_X1 U25103 ( .A1(n22201), .A2(keyinput51), .B1(keyinput62), .B2(n22200), 
        .ZN(n22199) );
  OAI221_X1 U25104 ( .B1(n22201), .B2(keyinput51), .C1(n22200), .C2(keyinput62), .A(n22199), .ZN(n22206) );
  AOI22_X1 U25105 ( .A1(n22204), .A2(keyinput93), .B1(n22203), .B2(keyinput48), 
        .ZN(n22202) );
  OAI221_X1 U25106 ( .B1(n22204), .B2(keyinput93), .C1(n22203), .C2(keyinput48), .A(n22202), .ZN(n22205) );
  NOR4_X1 U25107 ( .A1(n22208), .A2(n22207), .A3(n22206), .A4(n22205), .ZN(
        n22224) );
  AOI22_X1 U25108 ( .A1(n22210), .A2(keyinput47), .B1(keyinput114), .B2(n13754), .ZN(n22209) );
  OAI221_X1 U25109 ( .B1(n22210), .B2(keyinput47), .C1(n13754), .C2(
        keyinput114), .A(n22209), .ZN(n22222) );
  AOI22_X1 U25110 ( .A1(n22213), .A2(keyinput123), .B1(keyinput60), .B2(n22212), .ZN(n22211) );
  OAI221_X1 U25111 ( .B1(n22213), .B2(keyinput123), .C1(n22212), .C2(
        keyinput60), .A(n22211), .ZN(n22221) );
  XOR2_X1 U25112 ( .A(n22214), .B(keyinput29), .Z(n22219) );
  XOR2_X1 U25113 ( .A(n22215), .B(keyinput99), .Z(n22218) );
  XNOR2_X1 U25114 ( .A(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B(keyinput4), .ZN(
        n22217) );
  XNOR2_X1 U25115 ( .A(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B(keyinput34), .ZN(
        n22216) );
  NAND4_X1 U25116 ( .A1(n22219), .A2(n22218), .A3(n22217), .A4(n22216), .ZN(
        n22220) );
  NOR3_X1 U25117 ( .A1(n22222), .A2(n22221), .A3(n22220), .ZN(n22223) );
  NAND4_X1 U25118 ( .A1(n22226), .A2(n22225), .A3(n22224), .A4(n22223), .ZN(
        n22227) );
  NOR4_X1 U25119 ( .A1(n22230), .A2(n22229), .A3(n22228), .A4(n22227), .ZN(
        n22231) );
  OAI221_X1 U25120 ( .B1(keyinput14), .B2(n22233), .C1(keyinput14), .C2(n22232), .A(n22231), .ZN(n22234) );
  XNOR2_X1 U25121 ( .A(n22235), .B(n22234), .ZN(P2_U3140) );
  NOR2_X2 U11188 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n17149) );
  CLKBUF_X1 U11198 ( .A(n12295), .Z(n12618) );
  CLKBUF_X1 U11200 ( .A(n13385), .Z(n9713) );
  CLKBUF_X1 U11209 ( .A(n12306), .Z(n15907) );
  CLKBUF_X1 U11247 ( .A(n13825), .Z(n9734) );
  CLKBUF_X1 U11248 ( .A(n10899), .Z(n11476) );
  CLKBUF_X1 U11252 ( .A(n10970), .Z(n10973) );
  CLKBUF_X1 U11282 ( .A(n10898), .Z(n9735) );
  NOR2_X1 U11318 ( .A1(n18582), .A2(n18561), .ZN(n17574) );
  INV_X2 U12033 ( .A(n20171), .ZN(n19535) );
  AND2_X1 U12138 ( .A1(n17576), .A2(n17459), .ZN(n22236) );
endmodule

