

module b15_C_gen_AntiSAT_k_256_6 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput_f0, keyinput_f1, 
        keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, 
        keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, 
        keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, 
        keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, 
        keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, 
        keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, 
        keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, 
        keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, 
        keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, 
        keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, 
        keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, 
        keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, 
        keyinput_f62, keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66, 
        keyinput_f67, keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71, 
        keyinput_f72, keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76, 
        keyinput_f77, keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81, 
        keyinput_f82, keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86, 
        keyinput_f87, keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91, 
        keyinput_f92, keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96, 
        keyinput_f97, keyinput_f98, keyinput_f99, keyinput_f100, keyinput_f101, 
        keyinput_f102, keyinput_f103, keyinput_f104, keyinput_f105, 
        keyinput_f106, keyinput_f107, keyinput_f108, keyinput_f109, 
        keyinput_f110, keyinput_f111, keyinput_f112, keyinput_f113, 
        keyinput_f114, keyinput_f115, keyinput_f116, keyinput_f117, 
        keyinput_f118, keyinput_f119, keyinput_f120, keyinput_f121, 
        keyinput_f122, keyinput_f123, keyinput_f124, keyinput_f125, 
        keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, keyinput_g2, 
        keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, 
        keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, 
        keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, 
        keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, 
        keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, 
        keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, 
        keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, 
        keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, 
        keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, 
        keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, 
        keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, 
        keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, 
        keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, keyinput_g67, 
        keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, keyinput_g72, 
        keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, keyinput_g77, 
        keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, keyinput_g82, 
        keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, keyinput_g87, 
        keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, keyinput_g92, 
        keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, keyinput_g97, 
        keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101, 
        keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105, 
        keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109, 
        keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113, 
        keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117, 
        keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121, 
        keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125, 
        keyinput_g126, keyinput_g127, U3445, U3446, U3447, U3448, U3213, U3212, 
        U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, U3203, U3202, 
        U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, U3193, U3192, 
        U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, U3183, U3182, 
        U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, U3175, U3174, 
        U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, U3165, U3164, 
        U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, U3155, U3154, 
        U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, U3146, U3145, 
        U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, U3136, U3135, 
        U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, U3126, U3125, 
        U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, U3116, U3115, 
        U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, U3106, U3105, 
        U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, U3096, U3095, 
        U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, U3086, U3085, 
        U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, U3076, U3075, 
        U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, U3066, U3065, 
        U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, U3056, U3055, 
        U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, U3046, U3045, 
        U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, U3036, U3035, 
        U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, U3026, U3025, 
        U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, U3460, U3461, 
        U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, U3015, U3014, 
        U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, U3005, U3004, 
        U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, U2995, U2994, 
        U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, U2985, U2984, 
        U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, U2975, U2974, 
        U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, U2965, U2964, 
        U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, U2955, U2954, 
        U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, U2945, U2944, 
        U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, U2935, U2934, 
        U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, U2925, U2924, 
        U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, U2915, U2914, 
        U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, U2905, U2904, 
        U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, U2895, U2894, 
        U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, U2885, U2884, 
        U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, U2875, U2874, 
        U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, U2865, U2864, 
        U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, U2855, U2854, 
        U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, U2845, U2844, 
        U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, U2835, U2834, 
        U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, U2825, U2824, 
        U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, U2815, U2814, 
        U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, U2805, U2804, 
        U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, U2795, U3468, 
        U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, U3473, U2790, 
        U2789, U3474, U2788 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput_f0, keyinput_f1,
         keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6,
         keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11,
         keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16,
         keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21,
         keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26,
         keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31,
         keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36,
         keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41,
         keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46,
         keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51,
         keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56,
         keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61,
         keyinput_f62, keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66,
         keyinput_f67, keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71,
         keyinput_f72, keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76,
         keyinput_f77, keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81,
         keyinput_f82, keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86,
         keyinput_f87, keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91,
         keyinput_f92, keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96,
         keyinput_f97, keyinput_f98, keyinput_f99, keyinput_f100,
         keyinput_f101, keyinput_f102, keyinput_f103, keyinput_f104,
         keyinput_f105, keyinput_f106, keyinput_f107, keyinput_f108,
         keyinput_f109, keyinput_f110, keyinput_f111, keyinput_f112,
         keyinput_f113, keyinput_f114, keyinput_f115, keyinput_f116,
         keyinput_f117, keyinput_f118, keyinput_f119, keyinput_f120,
         keyinput_f121, keyinput_f122, keyinput_f123, keyinput_f124,
         keyinput_f125, keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1,
         keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6,
         keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11,
         keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16,
         keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21,
         keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26,
         keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31,
         keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36,
         keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41,
         keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46,
         keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51,
         keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56,
         keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61,
         keyinput_g62, keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66,
         keyinput_g67, keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71,
         keyinput_g72, keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76,
         keyinput_g77, keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81,
         keyinput_g82, keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86,
         keyinput_g87, keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91,
         keyinput_g92, keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96,
         keyinput_g97, keyinput_g98, keyinput_g99, keyinput_g100,
         keyinput_g101, keyinput_g102, keyinput_g103, keyinput_g104,
         keyinput_g105, keyinput_g106, keyinput_g107, keyinput_g108,
         keyinput_g109, keyinput_g110, keyinput_g111, keyinput_g112,
         keyinput_g113, keyinput_g114, keyinput_g115, keyinput_g116,
         keyinput_g117, keyinput_g118, keyinput_g119, keyinput_g120,
         keyinput_g121, keyinput_g122, keyinput_g123, keyinput_g124,
         keyinput_g125, keyinput_g126, keyinput_g127;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170,
         n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180,
         n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190,
         n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200,
         n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210,
         n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220,
         n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230,
         n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240,
         n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250,
         n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260,
         n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270,
         n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280,
         n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290,
         n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300,
         n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310,
         n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320,
         n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330,
         n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340,
         n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350,
         n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360,
         n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370,
         n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380,
         n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390,
         n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400,
         n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410,
         n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420,
         n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430,
         n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440,
         n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450,
         n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460,
         n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470,
         n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480,
         n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490,
         n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500,
         n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510,
         n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520,
         n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530,
         n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540,
         n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550,
         n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560,
         n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570,
         n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580,
         n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590,
         n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600,
         n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610,
         n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620,
         n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630,
         n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640,
         n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650,
         n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660,
         n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670,
         n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680,
         n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690,
         n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700,
         n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710,
         n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720,
         n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730,
         n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740,
         n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750,
         n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760,
         n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770,
         n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780,
         n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790,
         n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800,
         n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810,
         n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820,
         n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830,
         n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840,
         n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850,
         n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860,
         n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870,
         n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880,
         n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890,
         n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900,
         n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910,
         n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920,
         n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930,
         n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940,
         n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950,
         n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960,
         n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970,
         n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980,
         n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990,
         n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000,
         n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010,
         n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020,
         n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030,
         n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040,
         n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050,
         n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060,
         n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070,
         n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080,
         n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090,
         n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100,
         n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110,
         n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120,
         n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130,
         n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140,
         n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150,
         n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160,
         n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170,
         n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180,
         n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190,
         n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200,
         n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210,
         n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220,
         n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230,
         n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240,
         n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250,
         n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260,
         n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270,
         n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280,
         n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290,
         n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300,
         n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310,
         n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320,
         n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330,
         n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340,
         n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350,
         n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360,
         n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370,
         n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380,
         n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390,
         n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400,
         n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410,
         n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420,
         n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430,
         n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440,
         n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450,
         n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460,
         n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470,
         n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480,
         n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490,
         n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500,
         n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510,
         n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520,
         n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530,
         n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540,
         n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550,
         n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560,
         n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570,
         n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580,
         n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590,
         n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600,
         n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610,
         n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620,
         n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630,
         n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640,
         n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650,
         n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660,
         n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670,
         n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680,
         n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690,
         n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700,
         n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710,
         n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720,
         n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730,
         n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740,
         n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750,
         n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760,
         n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770,
         n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780,
         n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790,
         n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
         n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
         n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
         n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
         n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
         n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
         n4852, n4853, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6488, n6489, n6490, n6491, n6492, n6493,
         n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503,
         n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513,
         n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523,
         n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533,
         n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543,
         n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553,
         n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563,
         n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573,
         n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583,
         n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593,
         n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603,
         n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613,
         n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623,
         n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633,
         n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643,
         n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653,
         n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663,
         n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673,
         n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683,
         n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693,
         n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703,
         n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713,
         n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723,
         n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733,
         n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743,
         n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753,
         n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763,
         n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773,
         n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783,
         n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793,
         n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803,
         n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813,
         n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823,
         n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833,
         n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843,
         n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853,
         n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863,
         n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873,
         n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883,
         n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893,
         n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903,
         n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913,
         n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923,
         n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933,
         n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943,
         n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953,
         n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963,
         n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973,
         n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983,
         n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993,
         n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003,
         n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013,
         n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023,
         n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033,
         n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043,
         n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7052;

  CLKBUF_X2 U3609 ( .A(n4233), .Z(n4376) );
  CLKBUF_X2 U3610 ( .A(n3176), .Z(n4413) );
  CLKBUF_X2 U3611 ( .A(n3412), .Z(n3375) );
  CLKBUF_X2 U3612 ( .A(n3446), .Z(n4404) );
  CLKBUF_X2 U3613 ( .A(n3380), .Z(n4405) );
  CLKBUF_X1 U3614 ( .A(n4731), .Z(n3162) );
  AND4_X1 U3615 ( .A1(n3301), .A2(n3300), .A3(n3299), .A4(n3298), .ZN(n3312)
         );
  AND4_X1 U3616 ( .A1(n3241), .A2(n3240), .A3(n3239), .A4(n3238), .ZN(n3186)
         );
  AND2_X1 U3617 ( .A1(n4636), .A2(n3193), .ZN(n3419) );
  AND2_X2 U3618 ( .A1(n3198), .A2(n4524), .ZN(n3176) );
  INV_X1 U3620 ( .A(n7052), .ZN(n3161) );
  CLKBUF_X2 U3621 ( .A(n3419), .Z(n4417) );
  AND4_X1 U3622 ( .A1(n3280), .A2(n3279), .A3(n3278), .A4(n3277), .ZN(n3281)
         );
  AND2_X1 U3623 ( .A1(n3315), .A2(n3314), .ZN(n4239) );
  NAND2_X1 U3624 ( .A1(n3282), .A2(n3281), .ZN(n3287) );
  NAND2_X1 U3625 ( .A1(n4755), .A2(n4298), .ZN(n4784) );
  INV_X1 U3626 ( .A(n3178), .ZN(n4293) );
  BUF_X1 U3627 ( .A(n4303), .Z(n3175) );
  INV_X1 U3628 ( .A(n4387), .ZN(n4388) );
  INV_X1 U3629 ( .A(n4388), .ZN(n5452) );
  INV_X1 U3630 ( .A(n5907), .ZN(n4770) );
  NAND4_X2 U3631 ( .A1(n3313), .A2(n3312), .A3(n3311), .A4(n3310), .ZN(n5907)
         );
  NAND2_X1 U3632 ( .A1(n4391), .A2(n4390), .ZN(n5469) );
  INV_X1 U3633 ( .A(n5802), .ZN(n5885) );
  OAI211_X2 U3634 ( .C1(n4510), .C2(n3351), .A(n4519), .B(n4380), .ZN(n3352)
         );
  INV_X4 U3636 ( .A(n5203), .ZN(n3685) );
  NAND2_X1 U3637 ( .A1(n4274), .A2(n3500), .ZN(n4233) );
  INV_X1 U3638 ( .A(n4274), .ZN(n4731) );
  NAND2_X2 U3639 ( .A1(n3348), .A2(n5203), .ZN(n4567) );
  AND2_X2 U3640 ( .A1(n4239), .A2(n3318), .ZN(n3337) );
  NAND2_X2 U3641 ( .A1(n3186), .A2(n3188), .ZN(n4235) );
  AND4_X2 U3642 ( .A1(n3245), .A2(n3244), .A3(n3243), .A4(n3242), .ZN(n3188)
         );
  AND4_X4 U3643 ( .A1(n3227), .A2(n3226), .A3(n3225), .A4(n3224), .ZN(n5203)
         );
  NAND2_X1 U3645 ( .A1(n3556), .A2(n3555), .ZN(n3558) );
  XNOR2_X2 U3646 ( .A(n3392), .B(n3391), .ZN(n3491) );
  NAND2_X1 U3647 ( .A1(n4274), .A2(n3500), .ZN(n3163) );
  NAND2_X1 U3648 ( .A1(n4274), .A2(n3500), .ZN(n3164) );
  XNOR2_X2 U3649 ( .A(n3517), .B(n3516), .ZN(n3771) );
  INV_X2 U3650 ( .A(n3492), .ZN(n3516) );
  NAND2_X2 U3651 ( .A1(n3548), .A2(n3549), .ZN(n3584) );
  AND2_X4 U3652 ( .A1(n3200), .A2(n4524), .ZN(n3413) );
  NAND2_X2 U3653 ( .A1(n3207), .A2(n3206), .ZN(n3348) );
  AND4_X2 U3654 ( .A1(n3197), .A2(n3196), .A3(n3195), .A4(n3194), .ZN(n3207)
         );
  AND2_X2 U3655 ( .A1(n3201), .A2(n4631), .ZN(n3401) );
  NAND2_X2 U3656 ( .A1(n3655), .A2(n3654), .ZN(n5477) );
  BUF_X2 U3657 ( .A(n3395), .Z(n3437) );
  AOI21_X2 U3658 ( .B1(n3463), .B2(n3507), .A(n3624), .ZN(n3492) );
  NOR2_X1 U3659 ( .A1(n4618), .A2(n4623), .ZN(n4624) );
  INV_X1 U3661 ( .A(n3500), .ZN(n4675) );
  AND4_X1 U3662 ( .A1(n3260), .A2(n3259), .A3(n3258), .A4(n3257), .ZN(n3179)
         );
  AND4_X1 U3663 ( .A1(n3276), .A2(n3275), .A3(n3274), .A4(n3273), .ZN(n3282)
         );
  CLKBUF_X2 U3664 ( .A(n3374), .Z(n4402) );
  BUF_X2 U3665 ( .A(n3439), .Z(n4418) );
  CLKBUF_X2 U3666 ( .A(n3272), .Z(n3374) );
  BUF_X2 U3667 ( .A(n3403), .Z(n3414) );
  CLKBUF_X1 U3668 ( .A(n3468), .Z(n4645) );
  AND2_X2 U3669 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4630) );
  NOR2_X1 U3670 ( .A1(n5468), .A2(n4392), .ZN(n4393) );
  NOR2_X1 U3671 ( .A1(n5469), .A2(n5470), .ZN(n5468) );
  CLKBUF_X1 U3672 ( .A(n3661), .Z(n5513) );
  NOR2_X1 U3673 ( .A1(n5245), .A2(n5244), .ZN(n4439) );
  XNOR2_X1 U3674 ( .A(n5245), .B(n5244), .ZN(n5425) );
  CLKBUF_X1 U3675 ( .A(n5426), .Z(n5446) );
  OR2_X1 U3676 ( .A1(n5321), .A2(n4186), .ZN(n4187) );
  OR2_X1 U3677 ( .A1(n5365), .A2(n5366), .ZN(n5363) );
  NAND2_X1 U3678 ( .A1(n5370), .A2(n5368), .ZN(n5365) );
  CLKBUF_X1 U3679 ( .A(n5177), .Z(n5626) );
  NAND2_X1 U3680 ( .A1(n5633), .A2(n3641), .ZN(n5634) );
  CLKBUF_X1 U3681 ( .A(n5052), .Z(n5113) );
  NAND2_X1 U3682 ( .A1(n4377), .A2(n5250), .ZN(n4379) );
  AND2_X1 U3683 ( .A1(n5255), .A2(n5254), .ZN(n5486) );
  AND2_X1 U3684 ( .A1(n5110), .A2(n5112), .ZN(n5053) );
  AND2_X1 U3685 ( .A1(n3640), .A2(n5111), .ZN(n5632) );
  OR2_X1 U3686 ( .A1(n3863), .A2(n3862), .ZN(n3876) );
  AND2_X1 U3687 ( .A1(n3637), .A2(n5080), .ZN(n5112) );
  CLKBUF_X1 U3688 ( .A(n4799), .Z(n4817) );
  INV_X1 U3689 ( .A(n3636), .ZN(n5092) );
  INV_X1 U3690 ( .A(n3636), .ZN(n4387) );
  NOR2_X2 U3691 ( .A1(n5374), .A2(n4350), .ZN(n5356) );
  AND2_X1 U3692 ( .A1(n3623), .A2(n3603), .ZN(n3820) );
  AND2_X1 U3693 ( .A1(n4624), .A2(n4734), .ZN(n4735) );
  NAND2_X1 U3694 ( .A1(n3490), .A2(n3489), .ZN(n3533) );
  AND2_X1 U3695 ( .A1(n4697), .A2(n3526), .ZN(n5994) );
  OR2_X1 U3696 ( .A1(n6068), .A2(n3625), .ZN(n3503) );
  NAND2_X1 U3697 ( .A1(n3524), .A2(n3523), .ZN(n4698) );
  XNOR2_X1 U3698 ( .A(n3534), .B(n4689), .ZN(n4665) );
  INV_X1 U3699 ( .A(n6068), .ZN(n3165) );
  NAND2_X2 U3700 ( .A1(n5905), .A2(n4616), .ZN(n5413) );
  INV_X2 U3701 ( .A(n4500), .ZN(n4575) );
  AND2_X1 U3702 ( .A1(n3466), .A2(n3493), .ZN(n3467) );
  NAND2_X1 U3703 ( .A1(n3486), .A2(n3485), .ZN(n4689) );
  INV_X2 U3705 ( .A(n4501), .ZN(n4600) );
  INV_X2 U3706 ( .A(n5889), .ZN(n3166) );
  CLKBUF_X1 U3707 ( .A(n4517), .Z(n6071) );
  OR2_X1 U3708 ( .A1(n3777), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3504) );
  CLKBUF_X1 U3709 ( .A(n3777), .Z(n6624) );
  XNOR2_X1 U3710 ( .A(n3396), .B(n3437), .ZN(n4517) );
  NAND2_X1 U3711 ( .A1(n4243), .A2(n3341), .ZN(n3433) );
  OAI211_X1 U3712 ( .C1(n3469), .C2(n3664), .A(n3362), .B(n3361), .ZN(n3394)
         );
  CLKBUF_X2 U3713 ( .A(n3359), .Z(n3469) );
  AND2_X1 U3714 ( .A1(n3340), .A2(n3339), .ZN(n3341) );
  OAI21_X1 U3715 ( .B1(n3359), .B2(n6510), .A(n3325), .ZN(n3432) );
  NAND2_X1 U3716 ( .A1(n3350), .A2(n3349), .ZN(n4380) );
  CLKBUF_X1 U3717 ( .A(n4219), .Z(n4521) );
  AND2_X1 U3718 ( .A1(n3321), .A2(n4520), .ZN(n3329) );
  AND2_X1 U3719 ( .A1(n3266), .A2(n3330), .ZN(n3271) );
  NAND2_X1 U3720 ( .A1(n3269), .A2(n3268), .ZN(n3270) );
  AOI21_X1 U3721 ( .B1(n3319), .B2(n4235), .A(n3256), .ZN(n3266) );
  NAND2_X1 U3722 ( .A1(n4567), .A2(n4765), .ZN(n3319) );
  INV_X2 U3723 ( .A(n3317), .ZN(n4765) );
  INV_X2 U3724 ( .A(n4235), .ZN(n4680) );
  CLKBUF_X1 U3725 ( .A(n3317), .Z(n3389) );
  NAND2_X1 U3726 ( .A1(n3237), .A2(n3236), .ZN(n3317) );
  AND4_X1 U3727 ( .A1(n3291), .A2(n3290), .A3(n3289), .A4(n3288), .ZN(n3292)
         );
  AND4_X1 U3728 ( .A1(n3297), .A2(n3296), .A3(n3295), .A4(n3294), .ZN(n3313)
         );
  AND4_X1 U3729 ( .A1(n3309), .A2(n3308), .A3(n3307), .A4(n3306), .ZN(n3310)
         );
  AND4_X1 U3730 ( .A1(n3305), .A2(n3304), .A3(n3303), .A4(n3302), .ZN(n3311)
         );
  AND4_X1 U3731 ( .A1(n3211), .A2(n3210), .A3(n3209), .A4(n3208), .ZN(n3227)
         );
  NAND2_X2 U3732 ( .A1(STATE_REG_2__SCAN_IN), .A2(n7048), .ZN(n6602) );
  AND4_X1 U3733 ( .A1(n3215), .A2(n3214), .A3(n3213), .A4(n3212), .ZN(n3226)
         );
  AND4_X1 U3734 ( .A1(n3223), .A2(n3222), .A3(n3221), .A4(n3220), .ZN(n3224)
         );
  AND4_X1 U3735 ( .A1(n3231), .A2(n3230), .A3(n3229), .A4(n3228), .ZN(n3237)
         );
  AND4_X1 U3736 ( .A1(n3235), .A2(n3234), .A3(n3233), .A4(n3232), .ZN(n3236)
         );
  AND4_X1 U3737 ( .A1(n3265), .A2(n3264), .A3(n3263), .A4(n3262), .ZN(n3185)
         );
  BUF_X2 U3738 ( .A(n3413), .Z(n4415) );
  BUF_X2 U3739 ( .A(n3382), .Z(n4412) );
  BUF_X2 U3740 ( .A(n3420), .Z(n4169) );
  BUF_X2 U3741 ( .A(n3381), .Z(n4403) );
  BUF_X2 U3742 ( .A(n3261), .Z(n3380) );
  BUF_X2 U3743 ( .A(n3440), .Z(n4414) );
  INV_X2 U3744 ( .A(n6447), .ZN(n3167) );
  CLKBUF_X2 U3745 ( .A(n3401), .Z(n3445) );
  INV_X2 U3746 ( .A(n7047), .ZN(n7048) );
  AND2_X1 U3747 ( .A1(n3191), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3199)
         );
  AND2_X2 U3748 ( .A1(n4631), .A2(n4525), .ZN(n3412) );
  NOR2_X1 U3749 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3193) );
  AND2_X1 U3750 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4636) );
  INV_X1 U3751 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3668) );
  NAND2_X1 U3752 ( .A1(n3271), .A2(n3270), .ZN(n4203) );
  AND2_X2 U3753 ( .A1(n5217), .A2(n5307), .ZN(n5296) );
  AND2_X2 U3754 ( .A1(n4525), .A2(n4630), .ZN(n3168) );
  OR2_X4 U3755 ( .A1(n5104), .A2(n4327), .ZN(n5209) );
  AND2_X1 U3756 ( .A1(n3198), .A2(n3201), .ZN(n3169) );
  OR2_X4 U3757 ( .A1(n4784), .A2(n4819), .ZN(n4881) );
  NAND4_X1 U3758 ( .A1(n3313), .A2(n3312), .A3(n3311), .A4(n3310), .ZN(n3170)
         );
  NAND4_X1 U3759 ( .A1(n3313), .A2(n3312), .A3(n3311), .A4(n3310), .ZN(n3171)
         );
  AND2_X1 U3760 ( .A1(n4631), .A2(n4525), .ZN(n3172) );
  AND2_X4 U3761 ( .A1(n3198), .A2(n3201), .ZN(n3402) );
  AND2_X2 U3762 ( .A1(n5356), .A2(n5355), .ZN(n5358) );
  BUF_X4 U3763 ( .A(n3771), .Z(n4666) );
  OR2_X2 U3764 ( .A1(n4976), .A2(n4975), .ZN(n4978) );
  NAND2_X2 U3765 ( .A1(n3370), .A2(n3369), .ZN(n4652) );
  XNOR2_X2 U3766 ( .A(n3607), .B(n4789), .ZN(n4783) );
  OR2_X2 U3767 ( .A1(n5337), .A2(n5338), .ZN(n5340) );
  AND2_X2 U3768 ( .A1(n4911), .A2(n4910), .ZN(n4923) );
  NOR2_X4 U3769 ( .A1(n4881), .A2(n4882), .ZN(n4911) );
  OR2_X1 U3770 ( .A1(n3170), .A2(n4274), .ZN(n5002) );
  AND2_X1 U3771 ( .A1(n4636), .A2(n3193), .ZN(n3173) );
  AND2_X1 U3772 ( .A1(n4636), .A2(n3193), .ZN(n3174) );
  NOR2_X2 U3773 ( .A1(n3287), .A2(n3190), .ZN(n3293) );
  NAND2_X1 U3774 ( .A1(n4292), .A2(n4233), .ZN(n4303) );
  AND2_X4 U3775 ( .A1(n3171), .A2(n4274), .ZN(n3178) );
  NAND2_X4 U3776 ( .A1(n3293), .A2(n3292), .ZN(n4274) );
  NOR2_X4 U3777 ( .A1(n5049), .A2(n5050), .ZN(n5106) );
  OR2_X4 U3778 ( .A1(n4978), .A2(n4961), .ZN(n5049) );
  NAND2_X1 U3779 ( .A1(n4675), .A2(n3170), .ZN(n4292) );
  AOI21_X2 U3780 ( .B1(n3328), .B2(n3327), .A(n3181), .ZN(n4243) );
  INV_X1 U3781 ( .A(n4246), .ZN(n3327) );
  INV_X1 U3782 ( .A(n5002), .ZN(n4610) );
  NOR2_X2 U3783 ( .A1(n5320), .A2(n5319), .ZN(n5321) );
  OAI21_X1 U3784 ( .B1(n4203), .B2(n4274), .A(n4770), .ZN(n3326) );
  CLKBUF_X1 U3785 ( .A(n3401), .Z(n4407) );
  NAND2_X1 U3786 ( .A1(n5202), .A2(n3320), .ZN(n4204) );
  INV_X1 U3787 ( .A(n3319), .ZN(n3320) );
  INV_X1 U3788 ( .A(n5202), .ZN(n3256) );
  NAND2_X1 U3789 ( .A1(n3319), .A2(n4794), .ZN(n3268) );
  OR2_X1 U3790 ( .A1(n3426), .A2(n3425), .ZN(n3628) );
  INV_X1 U3791 ( .A(n5336), .ZN(n4122) );
  NAND2_X1 U3792 ( .A1(n4919), .A2(n3770), .ZN(n3823) );
  BUF_X1 U3793 ( .A(n4280), .Z(n4359) );
  INV_X1 U3794 ( .A(n4359), .ZN(n4346) );
  NOR2_X1 U3795 ( .A1(n3336), .A2(n3335), .ZN(n3340) );
  OR2_X1 U3796 ( .A1(n4495), .A2(READY_N), .ZN(n4497) );
  CLKBUF_X1 U3797 ( .A(n5196), .Z(n5197) );
  OR2_X1 U3798 ( .A1(n5452), .A2(n5673), .ZN(n4390) );
  INV_X1 U3799 ( .A(n5026), .ZN(n4289) );
  INV_X1 U3800 ( .A(n4518), .ZN(n3350) );
  AND2_X1 U3801 ( .A1(n4223), .A2(n4222), .ZN(n4384) );
  INV_X1 U3802 ( .A(n6135), .ZN(n6227) );
  OR2_X1 U3803 ( .A1(n6647), .A2(n4441), .ZN(n5820) );
  AND2_X1 U3804 ( .A1(n4453), .A2(n4446), .ZN(n5866) );
  INV_X1 U3805 ( .A(n5905), .ZN(n5900) );
  XNOR2_X1 U3806 ( .A(n4439), .B(n4438), .ZN(n5383) );
  INV_X1 U3807 ( .A(n6058), .ZN(n6041) );
  NAND2_X1 U3808 ( .A1(n3506), .A2(n3505), .ZN(n3510) );
  AND2_X1 U3809 ( .A1(n3678), .A2(n3679), .ZN(n3676) );
  INV_X1 U3810 ( .A(n3601), .ZN(n3599) );
  INV_X1 U3811 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3664) );
  INV_X1 U3812 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3468) );
  AND2_X1 U3813 ( .A1(n5002), .A2(n3686), .ZN(n3706) );
  AND2_X1 U3814 ( .A1(n4731), .A2(n5907), .ZN(n3487) );
  NAND2_X1 U3815 ( .A1(n3822), .A2(n3821), .ZN(n4799) );
  INV_X1 U3816 ( .A(n4801), .ZN(n3821) );
  NAND2_X1 U3817 ( .A1(n4387), .A2(n5427), .ZN(n3660) );
  NAND2_X1 U3818 ( .A1(n3634), .A2(n3633), .ZN(n4906) );
  INV_X1 U3819 ( .A(n4367), .ZN(n4361) );
  NOR2_X1 U3820 ( .A1(n4234), .A2(n3685), .ZN(n3343) );
  NAND2_X1 U3821 ( .A1(n3267), .A2(n3348), .ZN(n3269) );
  AND2_X1 U3822 ( .A1(n4274), .A2(n3685), .ZN(n3673) );
  OR2_X1 U3823 ( .A1(n3453), .A2(n3452), .ZN(n3520) );
  OR2_X1 U3824 ( .A1(n3388), .A2(n3387), .ZN(n3390) );
  INV_X1 U3825 ( .A(n3390), .ZN(n3499) );
  NOR2_X1 U3826 ( .A1(n3474), .A2(n6544), .ZN(n3709) );
  OR2_X1 U3827 ( .A1(n6068), .A2(n4687), .ZN(n6075) );
  INV_X1 U3828 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6521) );
  CLKBUF_X1 U3829 ( .A(n3487), .Z(n4490) );
  MUX2_X1 U3830 ( .A(n4280), .B(n4233), .S(EBX_REG_1__SCAN_IN), .Z(n4276) );
  NAND2_X1 U3831 ( .A1(n5820), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5008) );
  INV_X1 U3832 ( .A(n4615), .ZN(n4576) );
  AND2_X1 U3833 ( .A1(n4163), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4434)
         );
  INV_X1 U3834 ( .A(n5268), .ZN(n4143) );
  NOR2_X1 U3835 ( .A1(n4102), .A2(n4101), .ZN(n4103) );
  CLKBUF_X1 U3837 ( .A(n5332), .Z(n5333) );
  NAND2_X1 U3838 ( .A1(n4043), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4102)
         );
  AND2_X1 U3839 ( .A1(n5345), .A2(n5344), .ZN(n5352) );
  AND2_X1 U3840 ( .A1(n4064), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4063)
         );
  NOR2_X1 U3841 ( .A1(n3975), .A2(n3974), .ZN(n3976) );
  CLKBUF_X1 U3842 ( .A(n5290), .Z(n5291) );
  NOR2_X1 U3843 ( .A1(n3952), .A2(n5760), .ZN(n3953) );
  NAND2_X1 U3844 ( .A1(n3953), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3975)
         );
  NOR2_X1 U3845 ( .A1(n3909), .A2(n3893), .ZN(n3923) );
  OR2_X1 U3847 ( .A1(n3892), .A2(n5128), .ZN(n3909) );
  AND2_X1 U3849 ( .A1(n3857), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3858)
         );
  NOR2_X1 U3850 ( .A1(n3735), .A2(n5786), .ZN(n3824) );
  OR2_X1 U3851 ( .A1(n6634), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6644) );
  NOR2_X1 U3852 ( .A1(n3793), .A2(n5863), .ZN(n3798) );
  NAND2_X1 U3853 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3793) );
  AND2_X1 U3854 ( .A1(n4570), .A2(n6537), .ZN(n5546) );
  NAND2_X1 U3855 ( .A1(n4374), .A2(n4373), .ZN(n5232) );
  NOR2_X2 U3856 ( .A1(n5340), .A2(n5270), .ZN(n5324) );
  CLKBUF_X1 U3857 ( .A(n4196), .Z(n4197) );
  NAND2_X1 U3858 ( .A1(n4388), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n4389) );
  NAND2_X1 U3859 ( .A1(n4923), .A2(n4922), .ZN(n4976) );
  CLKBUF_X1 U3860 ( .A(n4906), .Z(n4907) );
  AND2_X1 U3861 ( .A1(n4283), .A2(n4282), .ZN(n5027) );
  OR2_X1 U3862 ( .A1(n4384), .A2(n4571), .ZN(n5064) );
  NAND2_X1 U3863 ( .A1(n3437), .A2(n3436), .ZN(n3777) );
  NAND2_X1 U3864 ( .A1(n3504), .A2(n3507), .ZN(n3506) );
  XNOR2_X1 U3865 ( .A(n3515), .B(n3514), .ZN(n3517) );
  NAND2_X1 U3866 ( .A1(n4652), .A2(n3373), .ZN(n4532) );
  INV_X1 U3867 ( .A(n6617), .ZN(n6620) );
  CLKBUF_X1 U3868 ( .A(n4665), .Z(n6070) );
  AND2_X1 U3869 ( .A1(n4666), .A2(n6253), .ZN(n6076) );
  INV_X1 U3870 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n4656) );
  NOR2_X1 U3871 ( .A1(n5851), .A2(n4457), .ZN(n5776) );
  AND2_X1 U3872 ( .A1(n5820), .A2(STATE2_REG_3__SCAN_IN), .ZN(n5849) );
  INV_X1 U3873 ( .A(n5851), .ZN(n5845) );
  INV_X1 U3874 ( .A(n5849), .ZN(n5886) );
  INV_X1 U3875 ( .A(n5862), .ZN(n5879) );
  AND2_X1 U3876 ( .A1(n4572), .A2(n6537), .ZN(n5892) );
  NAND2_X1 U3877 ( .A1(n4615), .A2(n4614), .ZN(n5905) );
  NOR2_X1 U3878 ( .A1(n6536), .A2(n5937), .ZN(n5952) );
  INV_X1 U3880 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n5990) );
  INV_X1 U3881 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n5863) );
  INV_X1 U3882 ( .A(n6010), .ZN(n5972) );
  NAND2_X1 U3883 ( .A1(n5989), .A2(n6011), .ZN(n6005) );
  INV_X1 U3884 ( .A(n5989), .ZN(n6012) );
  AND2_X1 U3885 ( .A1(n5546), .A2(n6526), .ZN(n6010) );
  OR2_X1 U3886 ( .A1(n4384), .A2(n4383), .ZN(n6058) );
  INV_X1 U3887 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6509) );
  CLKBUF_X1 U3888 ( .A(n4532), .Z(n4533) );
  INV_X1 U3889 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6403) );
  INV_X1 U3890 ( .A(n6156), .ZN(n6132) );
  INV_X1 U3891 ( .A(n6220), .ZN(n6187) );
  OR2_X1 U3892 ( .A1(n6232), .A2(n6231), .ZN(n6250) );
  INV_X1 U3893 ( .A(n6331), .ZN(n6356) );
  AND2_X1 U3894 ( .A1(n6448), .A2(n6398), .ZN(n6480) );
  INV_X1 U3895 ( .A(n6484), .ZN(n6502) );
  CLKBUF_X1 U3896 ( .A(n6598), .Z(n6606) );
  OAI21_X1 U3897 ( .B1(n5316), .B2(n5881), .A(n4466), .ZN(n4467) );
  NAND2_X1 U3898 ( .A1(n3623), .A2(n3627), .ZN(n3643) );
  AND2_X2 U3899 ( .A1(n4631), .A2(n4524), .ZN(n3446) );
  NOR2_X2 U3900 ( .A1(n4740), .A2(n4739), .ZN(n4738) );
  OAI221_X2 U3901 ( .B1(n6576), .B2(n6785), .C1(STATE_REG_1__SCAN_IN), .C2(
        n6785), .A(n7047), .ZN(n6608) );
  CLKBUF_X1 U3902 ( .A(n6433), .Z(n3180) );
  AND2_X1 U3903 ( .A1(n5907), .A2(n4235), .ZN(n3181) );
  NOR2_X2 U3904 ( .A1(n4828), .A2(n6070), .ZN(n3182) );
  INV_X1 U3905 ( .A(n4047), .ZN(n3790) );
  NAND2_X1 U3906 ( .A1(n4735), .A2(n4775), .ZN(n4774) );
  OR2_X1 U3907 ( .A1(n4388), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n3183)
         );
  AND2_X1 U3908 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6615), .ZN(n3184) );
  NOR2_X1 U3909 ( .A1(n5079), .A2(n5083), .ZN(n3187) );
  OR2_X1 U3910 ( .A1(n5228), .A2(n6447), .ZN(n3189) );
  NAND4_X1 U3911 ( .A1(n3286), .A2(n3285), .A3(n3284), .A4(n3283), .ZN(n3190)
         );
  AND2_X2 U3912 ( .A1(n3200), .A2(n3199), .ZN(n3440) );
  INV_X1 U3913 ( .A(n4236), .ZN(n3349) );
  INV_X1 U3914 ( .A(n5202), .ZN(n5381) );
  OR2_X1 U3915 ( .A1(n3690), .A2(n3692), .ZN(n3667) );
  OAI21_X1 U3916 ( .B1(n3338), .B2(n4675), .A(n4274), .ZN(n3339) );
  OR2_X1 U3917 ( .A1(n3681), .A2(n3680), .ZN(n3682) );
  INV_X1 U3918 ( .A(n3316), .ZN(n4205) );
  OR2_X1 U3919 ( .A1(n3409), .A2(n3408), .ZN(n3519) );
  INV_X1 U3920 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n6510) );
  NAND2_X1 U3921 ( .A1(n3323), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3359) );
  AND2_X2 U3922 ( .A1(n3668), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3200)
         );
  NAND2_X1 U3923 ( .A1(n3389), .A2(n5907), .ZN(n3474) );
  INV_X1 U3924 ( .A(n5199), .ZN(n3956) );
  AND2_X1 U3925 ( .A1(n3598), .A2(n3597), .ZN(n3601) );
  NOR2_X1 U3926 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5617) );
  NAND2_X1 U3927 ( .A1(n3178), .A2(n3164), .ZN(n4280) );
  OR2_X1 U3928 ( .A1(n3691), .A2(n3163), .ZN(n4520) );
  AND2_X1 U3929 ( .A1(n3474), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3713) );
  OR2_X1 U3930 ( .A1(n4303), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4275)
         );
  NOR2_X1 U3931 ( .A1(n4293), .A2(n4376), .ZN(n4367) );
  XNOR2_X1 U3932 ( .A(n3623), .B(n3613), .ZN(n3769) );
  AND2_X1 U3933 ( .A1(n5053), .A2(n5055), .ZN(n3638) );
  OR2_X1 U3934 ( .A1(n3797), .A2(n3891), .ZN(n3805) );
  AND2_X1 U3935 ( .A1(n4680), .A2(n3500), .ZN(n3720) );
  NOR2_X1 U3936 ( .A1(n4388), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n4392)
         );
  AND2_X1 U3937 ( .A1(n5452), .A2(n3647), .ZN(n3649) );
  INV_X1 U3938 ( .A(n4627), .ZN(n4288) );
  NAND2_X1 U3939 ( .A1(n3432), .A2(n3433), .ZN(n3395) );
  NAND2_X1 U3940 ( .A1(n6257), .A2(n6544), .ZN(n3486) );
  AND4_X1 U3941 ( .A1(n3205), .A2(n3204), .A3(n3203), .A4(n3202), .ZN(n3206)
         );
  AND2_X1 U3942 ( .A1(n3709), .A2(n3673), .ZN(n3694) );
  AOI21_X1 U3943 ( .B1(n3769), .B2(n3902), .A(n3768), .ZN(n4816) );
  AND2_X1 U3944 ( .A1(PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n4162), .ZN(n4163)
         );
  AND2_X1 U3945 ( .A1(n4063), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4043)
         );
  AND2_X1 U3946 ( .A1(n5635), .A2(n5632), .ZN(n3641) );
  AOI21_X1 U3947 ( .B1(n3165), .B2(n3902), .A(n3790), .ZN(n4621) );
  NAND2_X1 U3948 ( .A1(n4289), .A2(n4288), .ZN(n4740) );
  NAND2_X1 U3949 ( .A1(n5028), .A2(n5027), .ZN(n5026) );
  NAND2_X1 U3950 ( .A1(n3473), .A2(n3472), .ZN(n4892) );
  INV_X1 U3951 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6517) );
  AOI21_X1 U3952 ( .B1(n6650), .B2(n5545), .A(n6620), .ZN(n4674) );
  NAND2_X1 U3953 ( .A1(n5324), .A2(n5323), .ZN(n4371) );
  NOR2_X1 U3954 ( .A1(n3840), .A2(n5779), .ZN(n3857) );
  NOR2_X1 U3955 ( .A1(n3814), .A2(n5980), .ZN(n3764) );
  OR2_X1 U3956 ( .A1(n5008), .A2(n4987), .ZN(n5862) );
  OR2_X1 U3957 ( .A1(n5008), .A2(n4448), .ZN(n5851) );
  NAND2_X1 U3958 ( .A1(n5358), .A2(n5348), .ZN(n5337) );
  INV_X1 U3959 ( .A(n3891), .ZN(n3902) );
  NAND2_X1 U3960 ( .A1(n3661), .A2(n5510), .ZN(n5437) );
  NOR2_X1 U3961 ( .A1(n4095), .A2(n4039), .ZN(n4064) );
  AOI21_X1 U3962 ( .B1(n3820), .B2(n3902), .A(n3819), .ZN(n4801) );
  CLKBUF_X1 U3963 ( .A(n4735), .Z(n4776) );
  NAND2_X1 U3964 ( .A1(n5475), .A2(n4389), .ZN(n5612) );
  NAND2_X1 U3965 ( .A1(n3560), .A2(n3559), .ZN(n4750) );
  NAND2_X1 U3966 ( .A1(n3346), .A2(n3345), .ZN(n4519) );
  NOR2_X1 U3967 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4674), .ZN(n6135) );
  AND2_X1 U3968 ( .A1(n6070), .A2(n6068), .ZN(n6222) );
  NAND2_X1 U3969 ( .A1(n3508), .A2(n3507), .ZN(n3509) );
  OR2_X1 U3970 ( .A1(n6613), .A2(n4674), .ZN(n4795) );
  NAND2_X1 U3971 ( .A1(n3716), .A2(n3715), .ZN(n4570) );
  NAND2_X1 U3973 ( .A1(n3858), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3892)
         );
  AND2_X1 U3974 ( .A1(n5820), .A2(n4444), .ZN(n5804) );
  NOR2_X1 U3975 ( .A1(n3807), .A2(n5990), .ZN(n3815) );
  AND2_X1 U3976 ( .A1(n5820), .A2(n4992), .ZN(n5802) );
  INV_X1 U3977 ( .A(n5378), .ZN(n5888) );
  AND2_X1 U3978 ( .A1(n5905), .A2(n5204), .ZN(n5901) );
  AND2_X1 U3979 ( .A1(n5905), .A2(n3349), .ZN(n5897) );
  NAND2_X1 U3980 ( .A1(n5321), .A2(n4186), .ZN(n5245) );
  AND2_X1 U3981 ( .A1(n5605), .A2(n3167), .ZN(n5606) );
  NAND2_X1 U3982 ( .A1(n3976), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n4095)
         );
  OR2_X1 U3983 ( .A1(n5120), .A2(n5139), .ZN(n5151) );
  INV_X1 U3984 ( .A(n6005), .ZN(n5983) );
  OAI22_X1 U3985 ( .A1(n5460), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .B1(n5454), .B2(n5453), .ZN(n5455) );
  OAI21_X1 U3986 ( .B1(n4398), .B2(n4397), .A(n4396), .ZN(n4399) );
  NOR2_X1 U3987 ( .A1(n5689), .A2(n4248), .ZN(n5674) );
  INV_X1 U3988 ( .A(n5064), .ZN(n6048) );
  INV_X1 U3989 ( .A(n6033), .ZN(n6060) );
  INV_X1 U3990 ( .A(n6129), .ZN(n6119) );
  INV_X1 U3991 ( .A(n6102), .ZN(n6101) );
  AND2_X1 U3992 ( .A1(n4666), .A2(n6409), .ZN(n6398) );
  AND2_X1 U3993 ( .A1(n4726), .A2(n6076), .ZN(n6249) );
  AND2_X1 U3994 ( .A1(n6222), .A2(n6221), .ZN(n6254) );
  AND2_X1 U3995 ( .A1(n6222), .A2(n6398), .ZN(n6312) );
  NAND2_X2 U3996 ( .A1(n3510), .A2(n3509), .ZN(n6409) );
  NAND2_X1 U3997 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n4570), .ZN(n6617) );
  NAND2_X1 U3998 ( .A1(n5546), .A2(n4479), .ZN(n4495) );
  INV_X1 U3999 ( .A(n4467), .ZN(n4468) );
  INV_X1 U4000 ( .A(n5866), .ZN(n5881) );
  INV_X1 U4001 ( .A(n5804), .ZN(n5830) );
  OR2_X1 U4002 ( .A1(n5278), .A2(n5351), .ZN(n5463) );
  OR2_X1 U4003 ( .A1(n4497), .A2(n3162), .ZN(n4615) );
  INV_X1 U4004 ( .A(n5568), .ZN(n5450) );
  OR2_X1 U4005 ( .A1(n6010), .A2(n4189), .ZN(n5989) );
  OR2_X1 U4006 ( .A1(n5316), .A2(n6058), .ZN(n4385) );
  AOI21_X1 U4007 ( .B1(n5588), .B2(n6041), .A(n4399), .ZN(n4400) );
  OR2_X1 U4008 ( .A1(n4384), .A2(n4228), .ZN(n6033) );
  OR2_X1 U4009 ( .A1(n4384), .A2(n6511), .ZN(n6064) );
  NAND2_X1 U4010 ( .A1(n6101), .A2(n6409), .ZN(n6129) );
  NAND2_X1 U4011 ( .A1(n6101), .A2(n6253), .ZN(n6156) );
  OR2_X1 U4012 ( .A1(n4829), .A2(n6070), .ZN(n4957) );
  NAND2_X1 U4013 ( .A1(n6254), .A2(n6253), .ZN(n6318) );
  INV_X1 U4014 ( .A(n6480), .ZN(n6507) );
  INV_X1 U4015 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6615) );
  OAI211_X1 U4016 ( .C1(n4473), .C2(n6033), .A(n4386), .B(n4385), .ZN(U2987)
         );
  AND2_X2 U4017 ( .A1(n3468), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3198)
         );
  AND2_X4 U4018 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4524) );
  INV_X1 U4019 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3191) );
  NOR2_X4 U4020 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4631) );
  AND2_X2 U4021 ( .A1(n3199), .A2(n4631), .ZN(n3381) );
  AOI22_X1 U4022 ( .A1(n3176), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3381), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3197) );
  INV_X1 U4023 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3192) );
  AND2_X2 U4024 ( .A1(n3192), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3201)
         );
  AOI22_X1 U4025 ( .A1(n3402), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3401), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3196) );
  AND2_X2 U4026 ( .A1(n3201), .A2(n4630), .ZN(n3439) );
  AOI22_X1 U4027 ( .A1(n3439), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3419), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3195) );
  AND2_X4 U4028 ( .A1(n4630), .A2(n4524), .ZN(n3447) );
  AOI22_X1 U4029 ( .A1(n3440), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3194) );
  NOR2_X4 U4030 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4525) );
  AND2_X2 U4031 ( .A1(n3198), .A2(n4525), .ZN(n3382) );
  AND2_X2 U4032 ( .A1(n3199), .A2(n4630), .ZN(n3420) );
  AOI22_X1 U4033 ( .A1(n3382), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3420), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3205) );
  AND2_X2 U4034 ( .A1(n3200), .A2(n4525), .ZN(n3272) );
  AOI22_X1 U4035 ( .A1(n3272), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3172), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3204) );
  AND2_X2 U4036 ( .A1(n4525), .A2(n4630), .ZN(n3403) );
  AOI22_X1 U4037 ( .A1(n3413), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3168), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3203) );
  AND2_X2 U4038 ( .A1(n3201), .A2(n3200), .ZN(n3261) );
  AOI22_X1 U4039 ( .A1(n3261), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3446), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3202) );
  NAND2_X1 U4040 ( .A1(n3439), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3211)
         );
  NAND2_X1 U4041 ( .A1(n3402), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3210) );
  NAND2_X1 U4042 ( .A1(n3401), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3209) );
  NAND2_X1 U4043 ( .A1(n3174), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3208) );
  NAND2_X1 U4044 ( .A1(n3382), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3215) );
  NAND2_X1 U4045 ( .A1(n3420), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3214)
         );
  NAND2_X1 U4046 ( .A1(n3261), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3213) );
  NAND2_X1 U4047 ( .A1(n3446), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3212) );
  NAND2_X1 U4048 ( .A1(n3381), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3219) );
  NAND2_X1 U4049 ( .A1(n3440), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3218)
         );
  NAND2_X1 U4050 ( .A1(n3413), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3217)
         );
  NAND2_X1 U4051 ( .A1(n3168), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3216)
         );
  NAND2_X1 U4052 ( .A1(n3176), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3223) );
  NAND2_X1 U4053 ( .A1(n3272), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3222) );
  NAND2_X1 U4054 ( .A1(n3172), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3221) );
  NAND2_X1 U4055 ( .A1(n3447), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3220)
         );
  AOI22_X1 U4056 ( .A1(n3420), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3261), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3231) );
  AOI22_X1 U4057 ( .A1(n3381), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3413), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3230) );
  AOI22_X1 U4058 ( .A1(n3440), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3168), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3229) );
  AOI22_X1 U4059 ( .A1(n3382), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3446), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3228) );
  AOI22_X1 U4060 ( .A1(n3402), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3401), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3235) );
  AOI22_X1 U4061 ( .A1(n3176), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3272), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3234) );
  AOI22_X1 U4062 ( .A1(n3439), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3419), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3233) );
  AOI22_X1 U4063 ( .A1(n3412), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3232) );
  AOI22_X1 U4064 ( .A1(n3402), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3272), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3241) );
  AOI22_X1 U4065 ( .A1(n3401), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3446), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3240) );
  AOI22_X1 U4066 ( .A1(n3382), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3412), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3239) );
  AOI22_X1 U4067 ( .A1(n3439), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3419), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3238) );
  AOI22_X1 U4068 ( .A1(n3381), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3261), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3245) );
  AOI22_X1 U4069 ( .A1(n3420), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3413), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3244) );
  AOI22_X1 U4070 ( .A1(n3440), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3243) );
  AOI22_X1 U4071 ( .A1(n3176), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3403), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3242) );
  AOI22_X1 U4072 ( .A1(n3402), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3401), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3249) );
  AOI22_X1 U4073 ( .A1(n3176), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3374), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3248) );
  AOI22_X1 U4074 ( .A1(n3439), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3419), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3247) );
  AOI22_X1 U4075 ( .A1(n3412), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3246) );
  NAND4_X1 U4076 ( .A1(n3249), .A2(n3248), .A3(n3247), .A4(n3246), .ZN(n3255)
         );
  AOI22_X1 U4077 ( .A1(n3420), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3380), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3253) );
  AOI22_X1 U4078 ( .A1(n3381), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3413), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3252) );
  AOI22_X1 U4079 ( .A1(n3440), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3403), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3251) );
  AOI22_X1 U4080 ( .A1(n3382), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3446), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3250) );
  NAND4_X1 U4081 ( .A1(n3253), .A2(n3252), .A3(n3251), .A4(n3250), .ZN(n3254)
         );
  OR2_X2 U4082 ( .A1(n3255), .A2(n3254), .ZN(n5202) );
  INV_X2 U4083 ( .A(n3348), .ZN(n4794) );
  NAND2_X2 U4084 ( .A1(n3685), .A2(n4794), .ZN(n3316) );
  AOI22_X1 U4085 ( .A1(n3402), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3401), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3260) );
  AOI22_X1 U4086 ( .A1(n3176), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3374), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3259) );
  AOI22_X1 U4087 ( .A1(n3439), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3174), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3258) );
  AOI22_X1 U4088 ( .A1(n3412), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3257) );
  AOI22_X1 U4089 ( .A1(n3420), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3261), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3265) );
  AOI22_X1 U4090 ( .A1(n3381), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3413), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3264) );
  AOI22_X1 U4091 ( .A1(n3440), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3403), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3263) );
  AOI22_X1 U4092 ( .A1(n3382), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3446), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3262) );
  NAND2_X2 U4093 ( .A1(n3179), .A2(n3185), .ZN(n3500) );
  NAND2_X1 U4094 ( .A1(n3316), .A2(n3500), .ZN(n3330) );
  NAND2_X1 U4095 ( .A1(n4567), .A2(n4680), .ZN(n3267) );
  NAND2_X1 U4096 ( .A1(n3439), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3276)
         );
  NAND2_X1 U4097 ( .A1(n3169), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3275) );
  NAND2_X1 U4098 ( .A1(n3272), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3274) );
  NAND2_X1 U4099 ( .A1(n3173), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3273) );
  NAND2_X1 U4100 ( .A1(n3176), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3280) );
  NAND2_X1 U4101 ( .A1(n3403), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3279)
         );
  NAND2_X1 U4102 ( .A1(n3172), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3278) );
  NAND2_X1 U4103 ( .A1(n3446), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3277) );
  NAND2_X1 U4104 ( .A1(n3440), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3286)
         );
  NAND2_X1 U4105 ( .A1(n3413), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3285)
         );
  NAND2_X1 U4106 ( .A1(n3401), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3284) );
  NAND2_X1 U4107 ( .A1(n3447), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3283)
         );
  NAND2_X1 U4108 ( .A1(n3381), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3291) );
  NAND2_X1 U4109 ( .A1(n3382), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3290) );
  NAND2_X1 U4110 ( .A1(n3420), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3289)
         );
  NAND2_X1 U4111 ( .A1(n3380), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3288) );
  NAND2_X1 U4112 ( .A1(n3380), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3297) );
  NAND2_X1 U4113 ( .A1(n3439), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3296)
         );
  NAND2_X1 U4114 ( .A1(n3402), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3295) );
  NAND2_X1 U4115 ( .A1(n3374), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3294) );
  NAND2_X1 U4116 ( .A1(n3445), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3301) );
  NAND2_X1 U4117 ( .A1(n3440), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3300)
         );
  NAND2_X1 U4118 ( .A1(n3420), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3299)
         );
  NAND2_X1 U4119 ( .A1(n3413), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3298)
         );
  NAND2_X1 U4120 ( .A1(n3381), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3305) );
  NAND2_X1 U4121 ( .A1(n3382), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3304) );
  NAND2_X1 U4122 ( .A1(n3446), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3303) );
  NAND2_X1 U4123 ( .A1(n3168), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3302)
         );
  NAND2_X1 U4124 ( .A1(n3176), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3309) );
  NAND2_X1 U4125 ( .A1(n3412), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3308) );
  NAND2_X1 U4126 ( .A1(n3447), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3307)
         );
  NAND2_X1 U4127 ( .A1(n3419), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3306) );
  NAND2_X1 U4128 ( .A1(n4205), .A2(n4765), .ZN(n3315) );
  AND2_X1 U4129 ( .A1(n4567), .A2(n5202), .ZN(n3314) );
  NAND2_X1 U4130 ( .A1(n3316), .A2(n3389), .ZN(n3318) );
  NAND2_X1 U4131 ( .A1(STATE_REG_1__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n6568) );
  OAI21_X1 U4132 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .A(
        n6568), .ZN(n4210) );
  NAND2_X1 U4133 ( .A1(n3162), .A2(n4210), .ZN(n3344) );
  INV_X1 U4134 ( .A(n3720), .ZN(n4234) );
  AOI21_X1 U4135 ( .B1(n5203), .B2(n3344), .A(n4234), .ZN(n3322) );
  NAND2_X1 U4136 ( .A1(n4204), .A2(n3487), .ZN(n3321) );
  NAND2_X1 U4137 ( .A1(n4765), .A2(n3685), .ZN(n3691) );
  NAND4_X1 U4138 ( .A1(n3326), .A2(n3337), .A3(n3322), .A4(n3329), .ZN(n3323)
         );
  AND2_X1 U4139 ( .A1(n4656), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3717) );
  INV_X1 U4140 ( .A(n3717), .ZN(n3354) );
  NAND2_X1 U4141 ( .A1(n6615), .A2(n4656), .ZN(n6634) );
  INV_X1 U4142 ( .A(n6644), .ZN(n3353) );
  MUX2_X1 U4143 ( .A(n3354), .B(n3353), .S(n6509), .Z(n3324) );
  INV_X1 U4144 ( .A(n3324), .ZN(n3325) );
  INV_X1 U4145 ( .A(n3326), .ZN(n3328) );
  NOR2_X1 U4146 ( .A1(n3691), .A2(n3162), .ZN(n4246) );
  INV_X1 U4147 ( .A(n3329), .ZN(n3336) );
  NAND2_X1 U4148 ( .A1(n3330), .A2(n3487), .ZN(n3334) );
  INV_X1 U4149 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6544) );
  OR2_X1 U4150 ( .A1(n6634), .A2(n6544), .ZN(n6551) );
  INV_X1 U4151 ( .A(n6551), .ZN(n3333) );
  NAND2_X1 U4152 ( .A1(n3389), .A2(n5202), .ZN(n3718) );
  INV_X1 U4153 ( .A(n3718), .ZN(n3332) );
  NOR2_X1 U4154 ( .A1(n3500), .A2(n3348), .ZN(n3331) );
  NAND3_X1 U4155 ( .A1(n3332), .A2(n3331), .A3(n4680), .ZN(n4638) );
  NAND3_X1 U4156 ( .A1(n3334), .A2(n3333), .A3(n4638), .ZN(n3335) );
  INV_X1 U4157 ( .A(n3337), .ZN(n3338) );
  INV_X1 U4158 ( .A(n4204), .ZN(n3342) );
  NAND2_X1 U4159 ( .A1(n3343), .A2(n3342), .ZN(n4219) );
  OR2_X2 U4160 ( .A1(n4219), .A2(n4770), .ZN(n4510) );
  INV_X1 U4161 ( .A(n3344), .ZN(n3351) );
  INV_X1 U4162 ( .A(n4203), .ZN(n3346) );
  NOR2_X1 U4163 ( .A1(n3691), .A2(n5002), .ZN(n3345) );
  NOR2_X1 U4164 ( .A1(n3685), .A2(n3500), .ZN(n3347) );
  NAND3_X1 U4165 ( .A1(n4610), .A2(n4680), .A3(n3347), .ZN(n4518) );
  NAND2_X1 U4166 ( .A1(n3348), .A2(n5202), .ZN(n4236) );
  NAND2_X1 U4167 ( .A1(n3352), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3361) );
  INV_X1 U4168 ( .A(n3361), .ZN(n3358) );
  XNOR2_X1 U4169 ( .A(n6509), .B(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6294)
         );
  NAND2_X1 U4170 ( .A1(n3353), .A2(n6294), .ZN(n3356) );
  NAND2_X1 U4171 ( .A1(n3354), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3355) );
  NAND2_X1 U4172 ( .A1(n3356), .A2(n3355), .ZN(n3360) );
  OR2_X1 U4173 ( .A1(n3360), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3357)
         );
  NAND2_X1 U4174 ( .A1(n3358), .A2(n3357), .ZN(n3393) );
  NAND2_X1 U4175 ( .A1(n3395), .A2(n3393), .ZN(n3363) );
  INV_X1 U4176 ( .A(n3360), .ZN(n3362) );
  NAND2_X1 U4177 ( .A1(n3363), .A2(n3394), .ZN(n3372) );
  INV_X1 U4178 ( .A(n3372), .ZN(n3370) );
  INV_X1 U4179 ( .A(n3469), .ZN(n3368) );
  AND2_X1 U4180 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n3364) );
  NAND2_X1 U4181 ( .A1(n3364), .A2(n6521), .ZN(n4668) );
  INV_X1 U4182 ( .A(n3364), .ZN(n3365) );
  NAND2_X1 U4183 ( .A1(n3365), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3366) );
  AND2_X1 U4184 ( .A1(n4668), .A2(n3366), .ZN(n4897) );
  OAI22_X1 U4185 ( .A1(n4897), .A2(n6644), .B1(n3717), .B2(n6521), .ZN(n3367)
         );
  AOI21_X2 U4186 ( .B1(n3368), .B2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n3367), 
        .ZN(n3371) );
  INV_X1 U4187 ( .A(n3371), .ZN(n3369) );
  NAND2_X1 U4188 ( .A1(n3372), .A2(n3371), .ZN(n3373) );
  AOI22_X1 U4189 ( .A1(n3402), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4407), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3379) );
  AOI22_X1 U4190 ( .A1(n4413), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4402), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3378) );
  AOI22_X1 U4191 ( .A1(n4418), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4417), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3377) );
  INV_X1 U4192 ( .A(n3447), .ZN(n4637) );
  INV_X2 U4193 ( .A(n4637), .ZN(n4406) );
  AOI22_X1 U4194 ( .A1(n3375), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4406), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3376) );
  NAND4_X1 U4195 ( .A1(n3379), .A2(n3378), .A3(n3377), .A4(n3376), .ZN(n3388)
         );
  AOI22_X1 U4196 ( .A1(n4169), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4405), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3386) );
  AOI22_X1 U4197 ( .A1(n4403), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n4415), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3385) );
  AOI22_X1 U4198 ( .A1(n4414), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3168), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3384) );
  AOI22_X1 U4199 ( .A1(n4412), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4404), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3383) );
  NAND4_X1 U4200 ( .A1(n3386), .A2(n3385), .A3(n3384), .A4(n3383), .ZN(n3387)
         );
  NAND2_X1 U4201 ( .A1(n4765), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3431) );
  OAI22_X2 U4202 ( .A1(n4532), .A2(STATE2_REG_0__SCAN_IN), .B1(n3499), .B2(
        n3431), .ZN(n3392) );
  NOR2_X1 U4203 ( .A1(n5907), .A2(n6544), .ZN(n3428) );
  AOI22_X1 U4204 ( .A1(n3709), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3428), 
        .B2(n3390), .ZN(n3391) );
  NAND2_X1 U4205 ( .A1(n3394), .A2(n3393), .ZN(n3396) );
  INV_X1 U4206 ( .A(n3431), .ZN(n3410) );
  AOI22_X1 U4207 ( .A1(n4413), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4403), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3400) );
  AOI22_X1 U4208 ( .A1(n4414), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4402), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3399) );
  AOI22_X1 U4209 ( .A1(n4406), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n4417), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3398) );
  AOI22_X1 U4210 ( .A1(n4169), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4404), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3397) );
  NAND4_X1 U4211 ( .A1(n3400), .A2(n3399), .A3(n3398), .A4(n3397), .ZN(n3409)
         );
  AOI22_X1 U4212 ( .A1(n4412), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n4418), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3407) );
  AOI22_X1 U4213 ( .A1(n4407), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n4415), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3406) );
  BUF_X1 U4214 ( .A(n3402), .Z(n4416) );
  AOI22_X1 U4215 ( .A1(n3402), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3412), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3405) );
  AOI22_X1 U4216 ( .A1(n4405), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3403), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3404) );
  NAND4_X1 U4217 ( .A1(n3407), .A2(n3406), .A3(n3405), .A4(n3404), .ZN(n3408)
         );
  NAND2_X1 U4218 ( .A1(n3410), .A2(n3519), .ZN(n3411) );
  OAI21_X2 U4219 ( .B1(n4517), .B2(STATE2_REG_0__SCAN_IN), .A(n3411), .ZN(
        n3515) );
  AOI22_X1 U4220 ( .A1(n4414), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4405), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3418) );
  AOI22_X1 U4221 ( .A1(n4402), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3445), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3417) );
  AOI22_X1 U4222 ( .A1(n4403), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3412), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3416) );
  AOI22_X1 U4223 ( .A1(n3413), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3403), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3415) );
  NAND4_X1 U4224 ( .A1(n3418), .A2(n3417), .A3(n3416), .A4(n3415), .ZN(n3426)
         );
  AOI22_X1 U4225 ( .A1(n3176), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4412), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3424) );
  AOI22_X1 U4226 ( .A1(n4418), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4417), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3423) );
  AOI22_X1 U4227 ( .A1(n4169), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4404), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3422) );
  AOI22_X1 U4228 ( .A1(n3402), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3421) );
  NAND4_X1 U4229 ( .A1(n3424), .A2(n3423), .A3(n3422), .A4(n3421), .ZN(n3425)
         );
  INV_X1 U4230 ( .A(n3709), .ZN(n3612) );
  INV_X1 U4231 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3427) );
  OR2_X1 U4232 ( .A1(n3612), .A2(n3427), .ZN(n3430) );
  NAND2_X1 U4233 ( .A1(n3428), .A2(n3519), .ZN(n3429) );
  OAI211_X1 U4234 ( .C1(n3431), .C2(n3628), .A(n3430), .B(n3429), .ZN(n3514)
         );
  NAND2_X1 U4235 ( .A1(n3515), .A2(n3514), .ZN(n3495) );
  INV_X1 U4236 ( .A(n3432), .ZN(n3435) );
  INV_X1 U4237 ( .A(n3433), .ZN(n3434) );
  NAND2_X1 U4238 ( .A1(n3435), .A2(n3434), .ZN(n3436) );
  NAND2_X1 U4239 ( .A1(n4765), .A2(n3628), .ZN(n3462) );
  INV_X1 U4240 ( .A(n3628), .ZN(n3438) );
  NAND2_X1 U4241 ( .A1(n4765), .A2(n3438), .ZN(n3454) );
  AOI22_X1 U4242 ( .A1(n4412), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4418), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3444) );
  AOI22_X1 U4243 ( .A1(INSTQUEUE_REG_6__0__SCAN_IN), .A2(n3402), .B1(n4402), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3443) );
  AOI22_X1 U4244 ( .A1(n4403), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n4414), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3442) );
  AOI22_X1 U4245 ( .A1(n3176), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3413), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3441) );
  NAND4_X1 U4246 ( .A1(n3444), .A2(n3443), .A3(n3442), .A4(n3441), .ZN(n3453)
         );
  AOI22_X1 U4247 ( .A1(INSTQUEUE_REG_2__0__SCAN_IN), .A2(n3445), .B1(n3168), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3451) );
  AOI22_X1 U4248 ( .A1(n4405), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3375), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3450) );
  AOI22_X1 U4249 ( .A1(INSTQUEUE_REG_15__0__SCAN_IN), .A2(n4169), .B1(n4404), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3449) );
  AOI22_X1 U4250 ( .A1(n3447), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n4417), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3448) );
  NAND4_X1 U4251 ( .A1(n3451), .A2(n3450), .A3(n3449), .A4(n3448), .ZN(n3452)
         );
  MUX2_X1 U4252 ( .A(n3462), .B(n3454), .S(n3520), .Z(n3455) );
  INV_X1 U4253 ( .A(n3455), .ZN(n3456) );
  NAND2_X1 U4254 ( .A1(n3456), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3505) );
  NAND2_X1 U4255 ( .A1(n3504), .A2(n3505), .ZN(n3463) );
  INV_X1 U4256 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3457) );
  OR2_X1 U4257 ( .A1(n3612), .A2(n3457), .ZN(n3461) );
  INV_X1 U4258 ( .A(n3520), .ZN(n3458) );
  OAI211_X1 U4259 ( .C1(n3458), .C2(n3170), .A(n3462), .B(
        STATE2_REG_0__SCAN_IN), .ZN(n3459) );
  INV_X1 U4260 ( .A(n3459), .ZN(n3460) );
  NAND2_X1 U4261 ( .A1(n3461), .A2(n3460), .ZN(n3507) );
  NOR2_X1 U4262 ( .A1(n3462), .A2(n6544), .ZN(n3624) );
  NAND2_X1 U4263 ( .A1(n3495), .A2(n3492), .ZN(n3466) );
  INV_X1 U4264 ( .A(n3515), .ZN(n3465) );
  INV_X1 U4265 ( .A(n3514), .ZN(n3464) );
  NAND2_X1 U4266 ( .A1(n3465), .A2(n3464), .ZN(n3493) );
  NAND2_X2 U4267 ( .A1(n3491), .A2(n3467), .ZN(n3534) );
  OR2_X1 U4268 ( .A1(n3469), .A2(n4645), .ZN(n3473) );
  NAND3_X1 U4269 ( .A1(n6403), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6186) );
  NOR2_X1 U4270 ( .A1(n6509), .A2(n6186), .ZN(n6215) );
  OR2_X1 U4271 ( .A1(n6215), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3470)
         );
  NAND3_X1 U4272 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n6452) );
  NOR2_X1 U4273 ( .A1(n6509), .A2(n6452), .ZN(n6500) );
  INV_X1 U4274 ( .A(n6500), .ZN(n6440) );
  NAND2_X1 U4275 ( .A1(n3470), .A2(n6440), .ZN(n6223) );
  OAI22_X1 U4276 ( .A1(n6223), .A2(n6644), .B1(n3717), .B2(n6403), .ZN(n3471)
         );
  INV_X1 U4277 ( .A(n3471), .ZN(n3472) );
  XNOR2_X2 U4278 ( .A(n4652), .B(n4892), .ZN(n6257) );
  AOI22_X1 U4279 ( .A1(n3402), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4407), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3478) );
  AOI22_X1 U4280 ( .A1(n4413), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4402), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3477) );
  AOI22_X1 U4281 ( .A1(n4418), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4417), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3476) );
  AOI22_X1 U4282 ( .A1(n3375), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n4406), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3475) );
  NAND4_X1 U4283 ( .A1(n3478), .A2(n3477), .A3(n3476), .A4(n3475), .ZN(n3484)
         );
  AOI22_X1 U4284 ( .A1(n4169), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4405), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3482) );
  AOI22_X1 U4285 ( .A1(n4403), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n4415), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3481) );
  AOI22_X1 U4286 ( .A1(n4414), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3414), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3480) );
  AOI22_X1 U4287 ( .A1(n4412), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4404), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3479) );
  NAND4_X1 U4288 ( .A1(n3482), .A2(n3481), .A3(n3480), .A4(n3479), .ZN(n3483)
         );
  OR2_X1 U4289 ( .A1(n3484), .A2(n3483), .ZN(n3488) );
  AOI22_X1 U4290 ( .A1(n3709), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3713), 
        .B2(n3488), .ZN(n3485) );
  NAND2_X1 U4291 ( .A1(n4665), .A2(n3673), .ZN(n3490) );
  NAND2_X1 U4292 ( .A1(n3520), .A2(n3519), .ZN(n3518) );
  NAND2_X1 U4293 ( .A1(n3518), .A2(n3499), .ZN(n3498) );
  NAND2_X1 U4294 ( .A1(n3498), .A2(n3488), .ZN(n3575) );
  OAI211_X1 U4295 ( .C1(n3488), .C2(n3498), .A(n3575), .B(n4490), .ZN(n3489)
         );
  XNOR2_X1 U4296 ( .A(n3533), .B(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4706)
         );
  INV_X1 U4297 ( .A(n4706), .ZN(n3532) );
  INV_X1 U4298 ( .A(n3491), .ZN(n3496) );
  NAND2_X1 U4299 ( .A1(n3493), .A2(n3516), .ZN(n3494) );
  NAND3_X1 U4300 ( .A1(n3496), .A2(n3495), .A3(n3494), .ZN(n3497) );
  NAND2_X2 U4301 ( .A1(n3497), .A2(n3534), .ZN(n6068) );
  INV_X1 U4302 ( .A(n3673), .ZN(n3625) );
  OAI21_X1 U4303 ( .B1(n3499), .B2(n3518), .A(n3498), .ZN(n3501) );
  NAND2_X1 U4304 ( .A1(n4770), .A2(n3500), .ZN(n3511) );
  INV_X1 U4305 ( .A(n3511), .ZN(n4245) );
  AOI21_X1 U4306 ( .B1(n3501), .B2(n4490), .A(n4245), .ZN(n3502) );
  NAND2_X1 U4307 ( .A1(n3503), .A2(n3502), .ZN(n3527) );
  NAND2_X1 U4308 ( .A1(n3527), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n5991)
         );
  INV_X1 U4309 ( .A(n3505), .ZN(n3508) );
  INV_X1 U4310 ( .A(n4490), .ZN(n6649) );
  OAI21_X1 U4311 ( .B1(n6649), .B2(n3520), .A(n3511), .ZN(n3512) );
  INV_X1 U4312 ( .A(n3512), .ZN(n3513) );
  OAI21_X1 U4313 ( .B1(n6409), .B2(n3625), .A(n3513), .ZN(n6006) );
  NAND2_X1 U4314 ( .A1(n6006), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3525)
         );
  XNOR2_X1 U4315 ( .A(n3525), .B(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4699)
         );
  NAND2_X1 U4316 ( .A1(n4666), .A2(n3673), .ZN(n3524) );
  OAI21_X1 U4317 ( .B1(n3520), .B2(n3519), .A(n3518), .ZN(n3521) );
  OAI211_X1 U4318 ( .C1(n3521), .C2(n6649), .A(n3720), .B(n3685), .ZN(n3522)
         );
  INV_X1 U4319 ( .A(n3522), .ZN(n3523) );
  NAND2_X1 U4320 ( .A1(n4699), .A2(n4698), .ZN(n4697) );
  INV_X1 U4321 ( .A(n3525), .ZN(n6007) );
  NAND2_X1 U4322 ( .A1(n6007), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n3526)
         );
  NAND2_X1 U4323 ( .A1(n5991), .A2(n5994), .ZN(n3530) );
  INV_X1 U4324 ( .A(n3527), .ZN(n3529) );
  INV_X1 U4325 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3528) );
  NAND2_X1 U4326 ( .A1(n3529), .A2(n3528), .ZN(n5992) );
  NAND2_X1 U4327 ( .A1(n3530), .A2(n5992), .ZN(n4705) );
  INV_X1 U4328 ( .A(n4705), .ZN(n3531) );
  NAND2_X1 U4329 ( .A1(n3532), .A2(n3531), .ZN(n4744) );
  NAND2_X1 U4330 ( .A1(n3533), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4743)
         );
  INV_X1 U4331 ( .A(n3534), .ZN(n3535) );
  NAND2_X1 U4332 ( .A1(n3535), .A2(n4689), .ZN(n3551) );
  INV_X1 U4333 ( .A(n3551), .ZN(n3548) );
  NAND2_X1 U4334 ( .A1(n3709), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3547) );
  AOI22_X1 U4335 ( .A1(n3402), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n4407), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3539) );
  AOI22_X1 U4336 ( .A1(n4413), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4402), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3538) );
  AOI22_X1 U4337 ( .A1(n4418), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4417), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3537) );
  AOI22_X1 U4338 ( .A1(n3375), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n4406), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3536) );
  NAND4_X1 U4339 ( .A1(n3539), .A2(n3538), .A3(n3537), .A4(n3536), .ZN(n3545)
         );
  AOI22_X1 U4340 ( .A1(n4169), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4405), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3543) );
  AOI22_X1 U4341 ( .A1(n4403), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n4415), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3542) );
  AOI22_X1 U4342 ( .A1(n4414), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3414), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3541) );
  AOI22_X1 U4343 ( .A1(n4412), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4404), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3540) );
  NAND4_X1 U4344 ( .A1(n3543), .A2(n3542), .A3(n3541), .A4(n3540), .ZN(n3544)
         );
  OR2_X1 U4345 ( .A1(n3545), .A2(n3544), .ZN(n3573) );
  NAND2_X1 U4346 ( .A1(n3713), .A2(n3573), .ZN(n3546) );
  NAND2_X1 U4347 ( .A1(n3547), .A2(n3546), .ZN(n3549) );
  INV_X1 U4348 ( .A(n3549), .ZN(n3550) );
  NAND2_X1 U4349 ( .A1(n3551), .A2(n3550), .ZN(n3552) );
  NAND2_X1 U4350 ( .A1(n3584), .A2(n3552), .ZN(n3797) );
  INV_X1 U4351 ( .A(n3797), .ZN(n3553) );
  NAND2_X1 U4352 ( .A1(n3553), .A2(n3673), .ZN(n3556) );
  XNOR2_X1 U4353 ( .A(n3575), .B(n3573), .ZN(n3554) );
  NAND2_X1 U4354 ( .A1(n3554), .A2(n4490), .ZN(n3555) );
  NAND2_X1 U4355 ( .A1(n3558), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3559)
         );
  AND2_X1 U4356 ( .A1(n4743), .A2(n3559), .ZN(n3557) );
  NAND2_X1 U4357 ( .A1(n4744), .A2(n3557), .ZN(n4751) );
  INV_X1 U4358 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6027) );
  XNOR2_X2 U4359 ( .A(n3558), .B(n6027), .ZN(n4746) );
  INV_X1 U4360 ( .A(n4746), .ZN(n3560) );
  NAND2_X1 U4361 ( .A1(n3709), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3572) );
  AOI22_X1 U4362 ( .A1(n4413), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4403), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3564) );
  AOI22_X1 U4363 ( .A1(n4412), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4402), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3563) );
  AOI22_X1 U4364 ( .A1(n4418), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4417), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3562) );
  AOI22_X1 U4365 ( .A1(n3402), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4406), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3561) );
  NAND4_X1 U4366 ( .A1(n3564), .A2(n3563), .A3(n3562), .A4(n3561), .ZN(n3570)
         );
  AOI22_X1 U4367 ( .A1(n4414), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4169), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3568) );
  AOI22_X1 U4368 ( .A1(n4407), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n4415), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3567) );
  AOI22_X1 U4369 ( .A1(n3375), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n4404), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3566) );
  AOI22_X1 U4370 ( .A1(n4405), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3414), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3565) );
  NAND4_X1 U4371 ( .A1(n3568), .A2(n3567), .A3(n3566), .A4(n3565), .ZN(n3569)
         );
  OR2_X1 U4372 ( .A1(n3570), .A2(n3569), .ZN(n3576) );
  NAND2_X1 U4373 ( .A1(n3713), .A2(n3576), .ZN(n3571) );
  NAND2_X1 U4374 ( .A1(n3572), .A2(n3571), .ZN(n3585) );
  XNOR2_X1 U4375 ( .A(n3584), .B(n3585), .ZN(n3806) );
  NAND2_X1 U4376 ( .A1(n3806), .A2(n3673), .ZN(n3579) );
  INV_X1 U4377 ( .A(n3573), .ZN(n3574) );
  NOR2_X1 U4378 ( .A1(n3575), .A2(n3574), .ZN(n3577) );
  NAND2_X1 U4379 ( .A1(n3577), .A2(n3576), .ZN(n3614) );
  OAI211_X1 U4380 ( .C1(n3577), .C2(n3576), .A(n3614), .B(n4490), .ZN(n3578)
         );
  NAND2_X1 U4381 ( .A1(n3579), .A2(n3578), .ZN(n3581) );
  INV_X1 U4382 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3580) );
  XNOR2_X1 U4383 ( .A(n3581), .B(n3580), .ZN(n4752) );
  NAND3_X1 U4384 ( .A1(n4751), .A2(n4750), .A3(n4752), .ZN(n3583) );
  NAND2_X1 U4385 ( .A1(n3581), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3582)
         );
  NAND2_X1 U4386 ( .A1(n3583), .A2(n3582), .ZN(n4781) );
  INV_X1 U4387 ( .A(n3584), .ZN(n3586) );
  NAND2_X1 U4388 ( .A1(n3586), .A2(n3585), .ZN(n3602) );
  INV_X1 U4389 ( .A(n3602), .ZN(n3600) );
  NAND2_X1 U4390 ( .A1(n3709), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3598) );
  AOI22_X1 U4391 ( .A1(n3402), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4407), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3590) );
  AOI22_X1 U4392 ( .A1(n4413), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4402), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3589) );
  AOI22_X1 U4393 ( .A1(n4418), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4417), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3588) );
  AOI22_X1 U4394 ( .A1(n3375), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n4406), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3587) );
  NAND4_X1 U4395 ( .A1(n3590), .A2(n3589), .A3(n3588), .A4(n3587), .ZN(n3596)
         );
  AOI22_X1 U4396 ( .A1(n4169), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4405), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3594) );
  AOI22_X1 U4397 ( .A1(n4403), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n4415), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3593) );
  AOI22_X1 U4398 ( .A1(n4414), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3414), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3592) );
  AOI22_X1 U4399 ( .A1(n4412), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4404), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3591) );
  NAND4_X1 U4400 ( .A1(n3594), .A2(n3593), .A3(n3592), .A4(n3591), .ZN(n3595)
         );
  OR2_X1 U4401 ( .A1(n3596), .A2(n3595), .ZN(n3615) );
  NAND2_X1 U4402 ( .A1(n3713), .A2(n3615), .ZN(n3597) );
  NAND2_X2 U4403 ( .A1(n3600), .A2(n3599), .ZN(n3623) );
  NAND2_X1 U4404 ( .A1(n3602), .A2(n3601), .ZN(n3603) );
  NAND2_X1 U4405 ( .A1(n3820), .A2(n3673), .ZN(n3606) );
  XNOR2_X1 U4406 ( .A(n3614), .B(n3615), .ZN(n3604) );
  NAND2_X1 U4407 ( .A1(n3604), .A2(n4490), .ZN(n3605) );
  NAND2_X1 U4408 ( .A1(n3606), .A2(n3605), .ZN(n3607) );
  INV_X1 U4409 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4789) );
  NAND2_X1 U4410 ( .A1(n4781), .A2(n4783), .ZN(n3609) );
  NAND2_X1 U4411 ( .A1(n3607), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3608)
         );
  NAND2_X1 U4412 ( .A1(n3609), .A2(n3608), .ZN(n4885) );
  INV_X1 U4413 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3611) );
  NAND2_X1 U4414 ( .A1(n3713), .A2(n3628), .ZN(n3610) );
  OAI21_X1 U4415 ( .B1(n3612), .B2(n3611), .A(n3610), .ZN(n3613) );
  NAND2_X1 U4416 ( .A1(n3769), .A2(n3673), .ZN(n3619) );
  INV_X1 U4417 ( .A(n3614), .ZN(n3616) );
  NAND2_X1 U4418 ( .A1(n3616), .A2(n3615), .ZN(n3630) );
  XNOR2_X1 U4419 ( .A(n3630), .B(n3628), .ZN(n3617) );
  NAND2_X1 U4420 ( .A1(n3617), .A2(n4490), .ZN(n3618) );
  NAND2_X1 U4421 ( .A1(n3619), .A2(n3618), .ZN(n3620) );
  INV_X1 U4422 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4879) );
  XNOR2_X1 U4423 ( .A(n3620), .B(n4879), .ZN(n4886) );
  NAND2_X1 U4424 ( .A1(n4885), .A2(n4886), .ZN(n3622) );
  NAND2_X1 U4425 ( .A1(n3620), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3621)
         );
  NAND2_X1 U4426 ( .A1(n3622), .A2(n3621), .ZN(n4869) );
  INV_X1 U4427 ( .A(n3624), .ZN(n3626) );
  NOR2_X1 U4428 ( .A1(n3626), .A2(n3625), .ZN(n3627) );
  NAND2_X1 U4429 ( .A1(n4490), .A2(n3628), .ZN(n3629) );
  OR2_X1 U4430 ( .A1(n3630), .A2(n3629), .ZN(n3631) );
  NAND2_X1 U4431 ( .A1(n3643), .A2(n3631), .ZN(n3632) );
  INV_X1 U4432 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4878) );
  XNOR2_X1 U4433 ( .A(n3632), .B(n4878), .ZN(n4870) );
  NAND2_X1 U4434 ( .A1(n4869), .A2(n4870), .ZN(n3634) );
  NAND2_X1 U4435 ( .A1(n3632), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3633)
         );
  INV_X1 U4436 ( .A(n4906), .ZN(n3635) );
  INV_X1 U4437 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6017) );
  NOR2_X1 U4438 ( .A1(n3643), .A2(n6017), .ZN(n5079) );
  AND2_X1 U4439 ( .A1(n4388), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5083)
         );
  NAND2_X1 U4440 ( .A1(n3635), .A2(n3187), .ZN(n5052) );
  INV_X1 U4441 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5119) );
  NAND2_X1 U4442 ( .A1(n5092), .A2(n5119), .ZN(n5110) );
  INV_X1 U4443 ( .A(n3643), .ZN(n3636) );
  INV_X1 U4444 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n6018) );
  AND2_X1 U4445 ( .A1(n4387), .A2(n6018), .ZN(n5082) );
  INV_X1 U4446 ( .A(n5082), .ZN(n3637) );
  NAND2_X1 U4447 ( .A1(n4387), .A2(n6017), .ZN(n5080) );
  INV_X1 U4448 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n3639) );
  NAND2_X1 U4449 ( .A1(n5092), .A2(n3639), .ZN(n5055) );
  NAND2_X1 U4450 ( .A1(n5052), .A2(n3638), .ZN(n5633) );
  XNOR2_X1 U4451 ( .A(n5092), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5635)
         );
  NOR2_X1 U4452 ( .A1(n4387), .A2(n3639), .ZN(n5057) );
  INV_X1 U4453 ( .A(n5057), .ZN(n3640) );
  NAND2_X1 U4454 ( .A1(n4388), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5111) );
  INV_X1 U4455 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5095) );
  NAND2_X1 U4456 ( .A1(n5452), .A2(n5095), .ZN(n3642) );
  NAND2_X1 U4457 ( .A1(n5634), .A2(n3642), .ZN(n5091) );
  NAND2_X1 U4458 ( .A1(n4388), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n3644) );
  NAND2_X1 U4459 ( .A1(n5091), .A2(n3644), .ZN(n3646) );
  INV_X1 U4460 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5102) );
  NAND2_X1 U4461 ( .A1(n5452), .A2(n5102), .ZN(n3645) );
  NAND2_X1 U4462 ( .A1(n3646), .A2(n3645), .ZN(n5160) );
  INV_X1 U4463 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n3647) );
  NAND2_X1 U4464 ( .A1(n4388), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n3648) );
  OAI21_X2 U4465 ( .B1(n5160), .B2(n3649), .A(n3648), .ZN(n5177) );
  INV_X1 U4466 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5627) );
  NAND2_X1 U4467 ( .A1(n5452), .A2(n5627), .ZN(n3650) );
  NAND2_X1 U4468 ( .A1(n5177), .A2(n3650), .ZN(n5619) );
  INV_X1 U4469 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5622) );
  AND2_X1 U4470 ( .A1(n5617), .A2(n5622), .ZN(n3651) );
  NAND2_X1 U4471 ( .A1(n5619), .A2(n3651), .ZN(n3652) );
  NAND2_X1 U4472 ( .A1(n3652), .A2(n4388), .ZN(n3655) );
  INV_X1 U4473 ( .A(n5619), .ZN(n3653) );
  AND2_X1 U4474 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4252) );
  NAND2_X1 U4475 ( .A1(n3653), .A2(n4252), .ZN(n3654) );
  NOR2_X1 U4476 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n4397) );
  NOR2_X1 U4477 ( .A1(INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5666) );
  INV_X1 U4478 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5525) );
  INV_X1 U4479 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5531) );
  AND4_X1 U4480 ( .A1(n4397), .A2(n5666), .A3(n5525), .A4(n5531), .ZN(n3656)
         );
  NOR2_X1 U4481 ( .A1(n5092), .A2(n3656), .ZN(n3659) );
  AND2_X1 U4482 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5667) );
  AND2_X1 U4483 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4249) );
  NAND2_X1 U4484 ( .A1(n5667), .A2(n4249), .ZN(n5523) );
  NAND2_X1 U4485 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4260) );
  NOR2_X1 U4486 ( .A1(n5523), .A2(n4260), .ZN(n4268) );
  INV_X1 U4487 ( .A(n4268), .ZN(n3657) );
  NAND2_X1 U4488 ( .A1(n5092), .A2(n3657), .ZN(n3658) );
  OAI21_X1 U4489 ( .B1(n5477), .B2(n3659), .A(n3658), .ZN(n5426) );
  XNOR2_X1 U4490 ( .A(n5092), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5447)
         );
  NAND2_X1 U4491 ( .A1(n5426), .A2(n5447), .ZN(n4196) );
  INV_X1 U4492 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5427) );
  AND2_X2 U4493 ( .A1(n4196), .A2(n3660), .ZN(n3661) );
  NOR2_X1 U4494 ( .A1(n4387), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5511)
         );
  NOR2_X1 U4495 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5503) );
  NAND2_X1 U4496 ( .A1(n5511), .A2(n5503), .ZN(n4198) );
  AND2_X1 U4497 ( .A1(n4387), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5510)
         );
  NAND2_X1 U4498 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4269) );
  NOR2_X2 U4499 ( .A1(n5437), .A2(n4269), .ZN(n4195) );
  INV_X1 U4500 ( .A(n4195), .ZN(n3662) );
  OAI21_X1 U4501 ( .B1(n5513), .B2(n4198), .A(n3662), .ZN(n3663) );
  XNOR2_X1 U4502 ( .A(n3663), .B(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5501)
         );
  INV_X1 U4503 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n5722) );
  NAND2_X1 U4504 ( .A1(n6517), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3666) );
  NAND2_X1 U4505 ( .A1(n3664), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3665) );
  NAND2_X1 U4506 ( .A1(n3666), .A2(n3665), .ZN(n3690) );
  NAND2_X1 U4507 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n6509), .ZN(n3692) );
  NAND2_X1 U4508 ( .A1(n3667), .A2(n3666), .ZN(n3684) );
  NAND2_X1 U4509 ( .A1(n6521), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3671) );
  NAND2_X1 U4510 ( .A1(n3668), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3669) );
  NAND2_X1 U4511 ( .A1(n3671), .A2(n3669), .ZN(n3683) );
  INV_X1 U4512 ( .A(n3683), .ZN(n3670) );
  NAND2_X1 U4513 ( .A1(n3684), .A2(n3670), .ZN(n3672) );
  NAND2_X1 U4514 ( .A1(n3672), .A2(n3671), .ZN(n3678) );
  XNOR2_X1 U4515 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3679) );
  AOI21_X1 U4516 ( .B1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n6403), .A(n3676), 
        .ZN(n3674) );
  OAI222_X1 U4517 ( .A1(n5722), .A2(n3674), .B1(n5722), .B2(
        INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .C1(n3674), .C2(
        INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n4216) );
  NAND2_X1 U4518 ( .A1(n4216), .A2(n3694), .ZN(n3716) );
  NAND2_X1 U4519 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n3674), .ZN(n3675) );
  NOR2_X1 U4520 ( .A1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n3675), .ZN(n3681)
         );
  INV_X1 U4521 ( .A(n3676), .ZN(n3677) );
  OAI21_X1 U4522 ( .B1(n3679), .B2(n3678), .A(n3677), .ZN(n3680) );
  AOI22_X1 U4523 ( .A1(n3694), .A2(n3682), .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n6544), .ZN(n3711) );
  INV_X1 U4524 ( .A(n3682), .ZN(n4211) );
  XNOR2_X1 U4525 ( .A(n3684), .B(n3683), .ZN(n4214) );
  NAND2_X1 U4526 ( .A1(n4214), .A2(n3713), .ZN(n3707) );
  NAND2_X1 U4527 ( .A1(n3162), .A2(n3685), .ZN(n3686) );
  INV_X1 U4528 ( .A(n4214), .ZN(n3687) );
  NAND2_X1 U4529 ( .A1(n3709), .A2(n3687), .ZN(n3688) );
  AND3_X1 U4530 ( .A1(n3706), .A2(n3688), .A3(n3707), .ZN(n3705) );
  AOI21_X1 U4531 ( .B1(n3713), .B2(n4274), .A(n5203), .ZN(n3699) );
  INV_X1 U4532 ( .A(n3692), .ZN(n3689) );
  XNOR2_X1 U4533 ( .A(n3690), .B(n3689), .ZN(n4212) );
  NAND2_X1 U4534 ( .A1(n4212), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3696) );
  INV_X1 U4535 ( .A(n3691), .ZN(n4201) );
  OAI21_X1 U4536 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6509), .A(n3692), 
        .ZN(n3697) );
  OAI21_X1 U4537 ( .B1(n4201), .B2(n3697), .A(n5907), .ZN(n3693) );
  AOI22_X1 U4538 ( .A1(n3699), .A2(n3696), .B1(n3693), .B2(n3706), .ZN(n3703)
         );
  INV_X1 U4539 ( .A(n3694), .ZN(n3695) );
  OAI21_X1 U4540 ( .B1(n3699), .B2(n3696), .A(n3695), .ZN(n3702) );
  INV_X1 U4541 ( .A(n3713), .ZN(n3698) );
  NOR2_X1 U4542 ( .A1(n3698), .A2(n3697), .ZN(n3701) );
  NAND2_X1 U4543 ( .A1(n3699), .A2(n4212), .ZN(n3700) );
  AOI222_X1 U4544 ( .A1(n3703), .A2(n3702), .B1(n3703), .B2(n3701), .C1(n3702), 
        .C2(n3700), .ZN(n3704) );
  OAI22_X1 U4545 ( .A1(n3707), .A2(n3706), .B1(n3705), .B2(n3704), .ZN(n3708)
         );
  OAI21_X1 U4546 ( .B1(n3709), .B2(n4211), .A(n3708), .ZN(n3710) );
  NAND2_X1 U4547 ( .A1(n3711), .A2(n3710), .ZN(n3712) );
  AOI21_X1 U4548 ( .B1(n3713), .B2(n4216), .A(n3712), .ZN(n3714) );
  INV_X1 U4549 ( .A(n3714), .ZN(n3715) );
  NAND2_X1 U4550 ( .A1(n3717), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6550) );
  INV_X1 U4551 ( .A(n6550), .ZN(n6537) );
  OR2_X1 U4552 ( .A1(n3316), .A2(n3718), .ZN(n4229) );
  NAND2_X1 U4553 ( .A1(n4229), .A2(n4770), .ZN(n3719) );
  AND3_X1 U4554 ( .A1(n4239), .A2(n3720), .A3(n3719), .ZN(n4225) );
  AND2_X1 U4555 ( .A1(n4225), .A2(n4201), .ZN(n6526) );
  NAND2_X1 U4556 ( .A1(n3798), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3807)
         );
  NAND2_X1 U4557 ( .A1(n3815), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3814)
         );
  INV_X1 U4558 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n5980) );
  NAND2_X1 U4559 ( .A1(n3764), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3735)
         );
  INV_X1 U4560 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n5786) );
  XNOR2_X1 U4561 ( .A(n3824), .B(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n5086)
         );
  NOR2_X1 U4562 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n3993) );
  AOI22_X1 U4563 ( .A1(n4412), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4415), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3724) );
  AOI22_X1 U4564 ( .A1(n4418), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3414), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3723) );
  AOI22_X1 U4565 ( .A1(n4403), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4404), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3722) );
  AOI22_X1 U4566 ( .A1(n4413), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4417), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3721) );
  NAND4_X1 U4567 ( .A1(n3724), .A2(n3723), .A3(n3722), .A4(n3721), .ZN(n3730)
         );
  AOI22_X1 U4568 ( .A1(n4169), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4405), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3728) );
  AOI22_X1 U4569 ( .A1(n4416), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4407), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3727) );
  AOI22_X1 U4570 ( .A1(n4414), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3375), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3726) );
  AOI22_X1 U4571 ( .A1(n4402), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4406), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3725) );
  NAND4_X1 U4572 ( .A1(n3728), .A2(n3727), .A3(n3726), .A4(n3725), .ZN(n3729)
         );
  NAND2_X1 U4573 ( .A1(n4794), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3891) );
  OAI21_X1 U4574 ( .B1(n3730), .B2(n3729), .A(n3902), .ZN(n3733) );
  INV_X2 U4575 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6443) );
  OR2_X1 U4576 ( .A1(n5202), .A2(n6443), .ZN(n4049) );
  NAND2_X1 U4577 ( .A1(n4430), .A2(EAX_REG_10__SCAN_IN), .ZN(n3732) );
  NAND2_X1 U4578 ( .A1(n6443), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4047) );
  NAND2_X1 U4579 ( .A1(n3790), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3731)
         );
  NAND3_X1 U4580 ( .A1(n3733), .A2(n3732), .A3(n3731), .ZN(n3734) );
  AOI21_X1 U4581 ( .B1(n5086), .B2(n3993), .A(n3734), .ZN(n4918) );
  XNOR2_X1 U4582 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .B(n3735), .ZN(n5790) );
  INV_X1 U4583 ( .A(n5790), .ZN(n5014) );
  AOI22_X1 U4584 ( .A1(n4403), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n4418), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3739) );
  AOI22_X1 U4585 ( .A1(n4414), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4407), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3738) );
  AOI22_X1 U4586 ( .A1(n4169), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n3375), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3737) );
  AOI22_X1 U4587 ( .A1(n4413), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4417), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3736) );
  NAND4_X1 U4588 ( .A1(n3739), .A2(n3738), .A3(n3737), .A4(n3736), .ZN(n3745)
         );
  AOI22_X1 U4589 ( .A1(n4405), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4415), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3743) );
  AOI22_X1 U4590 ( .A1(n3402), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3414), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3742) );
  AOI22_X1 U4591 ( .A1(n4402), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4404), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3741) );
  AOI22_X1 U4592 ( .A1(n4412), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4406), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3740) );
  NAND4_X1 U4593 ( .A1(n3743), .A2(n3742), .A3(n3741), .A4(n3740), .ZN(n3744)
         );
  OAI21_X1 U4594 ( .B1(n3745), .B2(n3744), .A(n3902), .ZN(n3748) );
  NAND2_X1 U4595 ( .A1(n4430), .A2(EAX_REG_9__SCAN_IN), .ZN(n3747) );
  NAND2_X1 U4596 ( .A1(n3790), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3746)
         );
  NAND3_X1 U4597 ( .A1(n3748), .A2(n3747), .A3(n3746), .ZN(n3749) );
  AOI21_X1 U4598 ( .B1(n5014), .B2(n3993), .A(n3749), .ZN(n4968) );
  NOR2_X1 U4599 ( .A1(n4918), .A2(n4968), .ZN(n3763) );
  AOI22_X1 U4600 ( .A1(INSTQUEUE_REG_12__0__SCAN_IN), .A2(n4414), .B1(n4407), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3753) );
  AOI22_X1 U4601 ( .A1(INSTQUEUE_REG_0__0__SCAN_IN), .A2(n4169), .B1(n4405), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3752) );
  AOI22_X1 U4602 ( .A1(INSTQUEUE_REG_6__0__SCAN_IN), .A2(n4412), .B1(n4415), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3751) );
  AOI22_X1 U4603 ( .A1(n4403), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3414), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3750) );
  NAND4_X1 U4604 ( .A1(n3753), .A2(n3752), .A3(n3751), .A4(n3750), .ZN(n3759)
         );
  AOI22_X1 U4605 ( .A1(n4413), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3375), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3757) );
  AOI22_X1 U4606 ( .A1(n4402), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4404), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3756) );
  AOI22_X1 U4607 ( .A1(n4418), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4417), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3755) );
  AOI22_X1 U4608 ( .A1(n4416), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4406), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3754) );
  NAND4_X1 U4609 ( .A1(n3757), .A2(n3756), .A3(n3755), .A4(n3754), .ZN(n3758)
         );
  NOR2_X1 U4610 ( .A1(n3759), .A2(n3758), .ZN(n3762) );
  XNOR2_X1 U4611 ( .A(n3764), .B(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n5801) );
  NAND2_X1 U4612 ( .A1(n5801), .A2(n3993), .ZN(n3761) );
  AOI22_X1 U4613 ( .A1(n4430), .A2(EAX_REG_8__SCAN_IN), .B1(n3790), .B2(
        PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3760) );
  OAI211_X1 U4614 ( .C1(n3762), .C2(n3891), .A(n3761), .B(n3760), .ZN(n5019)
         );
  AND2_X1 U4615 ( .A1(n3763), .A2(n5019), .ZN(n4919) );
  AOI21_X1 U4616 ( .B1(n3814), .B2(n5980), .A(n3764), .ZN(n3765) );
  INV_X1 U4617 ( .A(n3765), .ZN(n5974) );
  NAND2_X1 U4618 ( .A1(n5974), .A2(n3993), .ZN(n3767) );
  AOI22_X1 U4619 ( .A1(n4430), .A2(EAX_REG_7__SCAN_IN), .B1(n3790), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3766) );
  NAND2_X1 U4620 ( .A1(n3767), .A2(n3766), .ZN(n3768) );
  INV_X1 U4621 ( .A(n4816), .ZN(n3770) );
  NAND2_X1 U4622 ( .A1(n3771), .A2(n3902), .ZN(n3775) );
  AOI22_X1 U4623 ( .A1(n4430), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n6443), .ZN(n3773) );
  AND2_X1 U4624 ( .A1(n3349), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3784) );
  NAND2_X1 U4625 ( .A1(n3784), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3772) );
  AND2_X1 U4626 ( .A1(n3773), .A2(n3772), .ZN(n3774) );
  NAND2_X1 U4627 ( .A1(n3775), .A2(n3774), .ZN(n4566) );
  AND2_X1 U4628 ( .A1(n4794), .A2(n5202), .ZN(n3776) );
  AOI21_X1 U4629 ( .B1(n6409), .B2(n3776), .A(n6443), .ZN(n4605) );
  OR2_X1 U4630 ( .A1(n6624), .A2(n3891), .ZN(n3781) );
  INV_X1 U4631 ( .A(n3784), .ZN(n3802) );
  NOR2_X1 U4632 ( .A1(n3802), .A2(n6510), .ZN(n3779) );
  INV_X1 U4633 ( .A(EAX_REG_0__SCAN_IN), .ZN(n5967) );
  INV_X1 U4634 ( .A(PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n5887) );
  OAI22_X1 U4635 ( .A1(n4049), .A2(n5967), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5887), .ZN(n3778) );
  NOR2_X1 U4636 ( .A1(n3779), .A2(n3778), .ZN(n3780) );
  NAND2_X1 U4637 ( .A1(n3781), .A2(n3780), .ZN(n3782) );
  NAND2_X1 U4638 ( .A1(n4605), .A2(n3782), .ZN(n4608) );
  INV_X1 U4639 ( .A(n3782), .ZN(n4606) );
  INV_X1 U4640 ( .A(n3993), .ZN(n4435) );
  INV_X1 U4641 ( .A(n4435), .ZN(n4183) );
  NAND2_X1 U4642 ( .A1(n4606), .A2(n4183), .ZN(n3783) );
  NAND2_X1 U4643 ( .A1(n4608), .A2(n3783), .ZN(n4565) );
  NAND2_X1 U4644 ( .A1(n4566), .A2(n4565), .ZN(n4619) );
  NAND2_X1 U4645 ( .A1(n3784), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3789) );
  INV_X2 U4646 ( .A(n4049), .ZN(n4430) );
  INV_X1 U4647 ( .A(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3786) );
  OAI21_X1 U4648 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n3793), .ZN(n5998) );
  NAND2_X1 U4649 ( .A1(n4183), .A2(n5998), .ZN(n3785) );
  OAI21_X1 U4650 ( .B1(n4047), .B2(n3786), .A(n3785), .ZN(n3787) );
  AOI21_X1 U4651 ( .B1(n4430), .B2(EAX_REG_2__SCAN_IN), .A(n3787), .ZN(n3788)
         );
  AND2_X1 U4652 ( .A1(n3789), .A2(n3788), .ZN(n4620) );
  OAI21_X1 U4653 ( .B1(n4619), .B2(n4620), .A(n4621), .ZN(n3792) );
  NAND2_X1 U4654 ( .A1(n4619), .A2(n4620), .ZN(n3791) );
  NAND2_X1 U4655 ( .A1(n3792), .A2(n3791), .ZN(n4618) );
  AOI21_X1 U4656 ( .B1(n5863), .B2(n3793), .A(n3798), .ZN(n5860) );
  OAI22_X1 U4657 ( .A1(n5860), .A2(n4435), .B1(n4047), .B2(n5863), .ZN(n3794)
         );
  AOI21_X1 U4658 ( .B1(n4430), .B2(EAX_REG_3__SCAN_IN), .A(n3794), .ZN(n3795)
         );
  OAI21_X1 U4659 ( .B1(n4645), .B2(n3802), .A(n3795), .ZN(n3796) );
  AOI21_X1 U4660 ( .B1(n4665), .B2(n3902), .A(n3796), .ZN(n4623) );
  OAI21_X1 U4661 ( .B1(n3798), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n3807), 
        .ZN(n5859) );
  INV_X1 U4662 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3799) );
  AOI21_X1 U4663 ( .B1(STATEBS16_REG_SCAN_IN), .B2(n3799), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3800) );
  AOI21_X1 U4664 ( .B1(n4430), .B2(EAX_REG_4__SCAN_IN), .A(n3800), .ZN(n3801)
         );
  OAI21_X1 U4665 ( .B1(n5722), .B2(n3802), .A(n3801), .ZN(n3803) );
  OAI21_X1 U4666 ( .B1(n5859), .B2(n4435), .A(n3803), .ZN(n3804) );
  NAND2_X1 U4667 ( .A1(n3805), .A2(n3804), .ZN(n4734) );
  NAND2_X1 U4668 ( .A1(n3806), .A2(n3902), .ZN(n3813) );
  INV_X1 U4669 ( .A(n3807), .ZN(n3809) );
  INV_X1 U4670 ( .A(n3815), .ZN(n3808) );
  OAI21_X1 U4671 ( .B1(PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n3809), .A(n3808), 
        .ZN(n5982) );
  NAND2_X1 U4672 ( .A1(n5982), .A2(n3993), .ZN(n3810) );
  OAI21_X1 U4673 ( .B1(n5990), .B2(n4047), .A(n3810), .ZN(n3811) );
  AOI21_X1 U4674 ( .B1(n4430), .B2(EAX_REG_5__SCAN_IN), .A(n3811), .ZN(n3812)
         );
  NAND2_X1 U4675 ( .A1(n3813), .A2(n3812), .ZN(n4775) );
  INV_X1 U4676 ( .A(n4774), .ZN(n3822) );
  INV_X1 U4677 ( .A(EAX_REG_6__SCAN_IN), .ZN(n3818) );
  OAI21_X1 U4678 ( .B1(n3815), .B2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n3814), 
        .ZN(n5836) );
  NAND2_X1 U4679 ( .A1(n5836), .A2(n3993), .ZN(n3817) );
  NAND2_X1 U4680 ( .A1(n3790), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3816)
         );
  OAI211_X1 U4681 ( .C1(n4049), .C2(n3818), .A(n3817), .B(n3816), .ZN(n3819)
         );
  NOR2_X1 U4682 ( .A1(n3823), .A2(n4799), .ZN(n4959) );
  NAND2_X1 U4683 ( .A1(n3824), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3840)
         );
  INV_X1 U4684 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n5779) );
  INV_X1 U4685 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5074) );
  XNOR2_X1 U4686 ( .A(n3857), .B(n5074), .ZN(n5071) );
  NAND2_X1 U4687 ( .A1(n5071), .A2(n3993), .ZN(n3827) );
  INV_X1 U4688 ( .A(EAX_REG_12__SCAN_IN), .ZN(n5041) );
  INV_X1 U4689 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6852) );
  OAI21_X1 U4690 ( .B1(n6852), .B2(PHYADDRPOINTER_REG_12__SCAN_IN), .A(n6443), 
        .ZN(n3825) );
  OAI21_X1 U4691 ( .B1(n4049), .B2(n5041), .A(n3825), .ZN(n3826) );
  NAND2_X1 U4692 ( .A1(n3827), .A2(n3826), .ZN(n3839) );
  AOI22_X1 U4693 ( .A1(n4416), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4402), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3831) );
  AOI22_X1 U4694 ( .A1(n4414), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4169), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3830) );
  AOI22_X1 U4695 ( .A1(n4405), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4407), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3829) );
  AOI22_X1 U4696 ( .A1(n4418), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4417), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3828) );
  NAND4_X1 U4697 ( .A1(n3831), .A2(n3830), .A3(n3829), .A4(n3828), .ZN(n3837)
         );
  AOI22_X1 U4698 ( .A1(n4403), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3375), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3835) );
  AOI22_X1 U4699 ( .A1(n4415), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3414), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3834) );
  AOI22_X1 U4700 ( .A1(n4412), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n4404), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3833) );
  AOI22_X1 U4701 ( .A1(n4413), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4406), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3832) );
  NAND4_X1 U4702 ( .A1(n3835), .A2(n3834), .A3(n3833), .A4(n3832), .ZN(n3836)
         );
  OAI21_X1 U4703 ( .B1(n3837), .B2(n3836), .A(n3902), .ZN(n3838) );
  NAND2_X1 U4704 ( .A1(n3839), .A2(n3838), .ZN(n4960) );
  XNOR2_X1 U4705 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .B(n3840), .ZN(n5968)
         );
  INV_X1 U4706 ( .A(n5968), .ZN(n3855) );
  AOI22_X1 U4707 ( .A1(n4405), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4415), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3844) );
  AOI22_X1 U4708 ( .A1(n4416), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3414), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3843) );
  AOI22_X1 U4709 ( .A1(n4418), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4417), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3842) );
  AOI22_X1 U4710 ( .A1(n4404), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4406), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3841) );
  NAND4_X1 U4711 ( .A1(n3844), .A2(n3843), .A3(n3842), .A4(n3841), .ZN(n3850)
         );
  AOI22_X1 U4712 ( .A1(n4413), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4407), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3848) );
  AOI22_X1 U4713 ( .A1(n4412), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4169), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3847) );
  AOI22_X1 U4714 ( .A1(n4403), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4402), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3846) );
  AOI22_X1 U4715 ( .A1(n4414), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3375), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3845) );
  NAND4_X1 U4716 ( .A1(n3848), .A2(n3847), .A3(n3846), .A4(n3845), .ZN(n3849)
         );
  OAI21_X1 U4717 ( .B1(n3850), .B2(n3849), .A(n3902), .ZN(n3853) );
  NAND2_X1 U4718 ( .A1(n4430), .A2(EAX_REG_11__SCAN_IN), .ZN(n3852) );
  NAND2_X1 U4719 ( .A1(n3790), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3851)
         );
  NAND3_X1 U4720 ( .A1(n3853), .A2(n3852), .A3(n3851), .ZN(n3854) );
  AOI21_X1 U4721 ( .B1(n3855), .B2(n3993), .A(n3854), .ZN(n4974) );
  INV_X1 U4722 ( .A(n4974), .ZN(n4958) );
  AND2_X1 U4723 ( .A1(n4960), .A2(n4958), .ZN(n3856) );
  NAND2_X1 U4724 ( .A1(n4959), .A2(n3856), .ZN(n3863) );
  INV_X1 U4725 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3860) );
  OAI21_X1 U4726 ( .B1(PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n3858), .A(n3892), 
        .ZN(n5775) );
  NAND2_X1 U4727 ( .A1(n5775), .A2(n3993), .ZN(n3859) );
  OAI21_X1 U4728 ( .B1(n3860), .B2(n4047), .A(n3859), .ZN(n3861) );
  AOI21_X1 U4729 ( .B1(n4430), .B2(EAX_REG_13__SCAN_IN), .A(n3861), .ZN(n3862)
         );
  NAND2_X1 U4730 ( .A1(n3863), .A2(n3862), .ZN(n3864) );
  AND2_X2 U4731 ( .A1(n3876), .A2(n3864), .ZN(n5038) );
  AOI22_X1 U4732 ( .A1(n4413), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4418), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3868) );
  AOI22_X1 U4733 ( .A1(n4169), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n4405), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3867) );
  AOI22_X1 U4734 ( .A1(n4402), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4407), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3866) );
  AOI22_X1 U4735 ( .A1(n4403), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n4404), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3865) );
  NAND4_X1 U4736 ( .A1(n3868), .A2(n3867), .A3(n3866), .A4(n3865), .ZN(n3874)
         );
  AOI22_X1 U4737 ( .A1(n4412), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4415), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3872) );
  AOI22_X1 U4738 ( .A1(n4414), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3375), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3871) );
  AOI22_X1 U4739 ( .A1(n4416), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3414), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3870) );
  AOI22_X1 U4740 ( .A1(n4406), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n4417), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3869) );
  NAND4_X1 U4741 ( .A1(n3872), .A2(n3871), .A3(n3870), .A4(n3869), .ZN(n3873)
         );
  OR2_X1 U4742 ( .A1(n3874), .A2(n3873), .ZN(n3875) );
  AND2_X1 U4743 ( .A1(n3902), .A2(n3875), .ZN(n5037) );
  NAND2_X1 U4744 ( .A1(n5038), .A2(n5037), .ZN(n5036) );
  NAND2_X1 U4745 ( .A1(n5036), .A2(n3876), .ZN(n5122) );
  AOI22_X1 U4746 ( .A1(n4403), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4405), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3880) );
  AOI22_X1 U4747 ( .A1(n4169), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n4415), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3879) );
  AOI22_X1 U4748 ( .A1(n4406), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n4417), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3878) );
  AOI22_X1 U4749 ( .A1(n4413), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3414), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3877) );
  NAND4_X1 U4750 ( .A1(n3880), .A2(n3879), .A3(n3878), .A4(n3877), .ZN(n3886)
         );
  AOI22_X1 U4751 ( .A1(n4412), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4418), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3884) );
  AOI22_X1 U4752 ( .A1(n4416), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4402), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3883) );
  AOI22_X1 U4753 ( .A1(n4414), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3375), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3882) );
  AOI22_X1 U4754 ( .A1(n4407), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n4404), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3881) );
  NAND4_X1 U4755 ( .A1(n3884), .A2(n3883), .A3(n3882), .A4(n3881), .ZN(n3885)
         );
  NOR2_X1 U4756 ( .A1(n3886), .A2(n3885), .ZN(n3890) );
  XNOR2_X1 U4757 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .B(n3892), .ZN(n5193)
         );
  INV_X1 U4758 ( .A(n5193), .ZN(n3887) );
  AOI22_X1 U4759 ( .A1(n3790), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .B1(n4183), 
        .B2(n3887), .ZN(n3889) );
  NAND2_X1 U4760 ( .A1(n4430), .A2(EAX_REG_14__SCAN_IN), .ZN(n3888) );
  OAI211_X1 U4761 ( .C1(n3891), .C2(n3890), .A(n3889), .B(n3888), .ZN(n5121)
         );
  NAND2_X1 U4762 ( .A1(n5122), .A2(n5121), .ZN(n5120) );
  INV_X1 U4763 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5128) );
  INV_X1 U4764 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3893) );
  XNOR2_X1 U4765 ( .A(n3909), .B(n3893), .ZN(n5162) );
  AOI22_X1 U4766 ( .A1(n4416), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4402), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3897) );
  AOI22_X1 U4767 ( .A1(n4412), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4404), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3896) );
  AOI22_X1 U4768 ( .A1(n4407), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n4417), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3895) );
  AOI22_X1 U4769 ( .A1(n4414), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4406), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3894) );
  NAND4_X1 U4770 ( .A1(n3897), .A2(n3896), .A3(n3895), .A4(n3894), .ZN(n3904)
         );
  AOI22_X1 U4771 ( .A1(n4413), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4405), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3901) );
  AOI22_X1 U4772 ( .A1(n4403), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n4415), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3900) );
  AOI22_X1 U4773 ( .A1(n4418), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3375), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3899) );
  AOI22_X1 U4774 ( .A1(n4169), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3414), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3898) );
  NAND4_X1 U4775 ( .A1(n3901), .A2(n3900), .A3(n3899), .A4(n3898), .ZN(n3903)
         );
  OAI21_X1 U4776 ( .B1(n3904), .B2(n3903), .A(n3902), .ZN(n3907) );
  NAND2_X1 U4777 ( .A1(n4430), .A2(EAX_REG_15__SCAN_IN), .ZN(n3906) );
  NAND2_X1 U4778 ( .A1(n3790), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3905)
         );
  NAND3_X1 U4779 ( .A1(n3907), .A2(n3906), .A3(n3905), .ZN(n3908) );
  AOI21_X1 U4780 ( .B1(n5162), .B2(n4183), .A(n3908), .ZN(n5139) );
  XOR2_X1 U4781 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .B(n3923), .Z(n5225) );
  INV_X1 U4782 ( .A(n5225), .ZN(n5171) );
  INV_X1 U4783 ( .A(n4229), .ZN(n6622) );
  NAND2_X1 U4784 ( .A1(n6622), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4432) );
  AOI22_X1 U4785 ( .A1(n4413), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4418), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3913) );
  AOI22_X1 U4786 ( .A1(n4403), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3445), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3912) );
  AOI22_X1 U4787 ( .A1(INSTQUEUE_REG_12__0__SCAN_IN), .A2(n4405), .B1(n4415), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3911) );
  AOI22_X1 U4788 ( .A1(n3375), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n3414), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3910) );
  NAND4_X1 U4789 ( .A1(n3913), .A2(n3912), .A3(n3911), .A4(n3910), .ZN(n3919)
         );
  AOI22_X1 U4790 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n4414), .B1(n4169), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3917) );
  AOI22_X1 U4791 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n4412), .B1(n4402), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3916) );
  AOI22_X1 U4792 ( .A1(n4406), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n4417), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3915) );
  AOI22_X1 U4793 ( .A1(n4416), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4404), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3914) );
  NAND4_X1 U4794 ( .A1(n3917), .A2(n3916), .A3(n3915), .A4(n3914), .ZN(n3918)
         );
  NOR2_X1 U4795 ( .A1(n3919), .A2(n3918), .ZN(n3921) );
  AOI22_X1 U4796 ( .A1(n4430), .A2(EAX_REG_16__SCAN_IN), .B1(n3790), .B2(
        PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3920) );
  OAI21_X1 U4797 ( .B1(n4432), .B2(n3921), .A(n3920), .ZN(n3922) );
  AOI21_X1 U4798 ( .B1(n5171), .B2(n4183), .A(n3922), .ZN(n5150) );
  NOR2_X2 U4799 ( .A1(n5151), .A2(n5150), .ZN(n5152) );
  NAND2_X1 U4800 ( .A1(n3923), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3952)
         );
  XNOR2_X1 U4801 ( .A(n3952), .B(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5758)
         );
  AOI22_X1 U4802 ( .A1(n4430), .A2(EAX_REG_17__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n6443), .ZN(n3937) );
  AOI22_X1 U4803 ( .A1(n4169), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n4405), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3927) );
  AOI22_X1 U4804 ( .A1(n4402), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3375), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3926) );
  AOI22_X1 U4805 ( .A1(n4415), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3414), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3925) );
  AOI22_X1 U4806 ( .A1(n4418), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n4406), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3924) );
  NAND4_X1 U4807 ( .A1(n3927), .A2(n3926), .A3(n3925), .A4(n3924), .ZN(n3935)
         );
  AOI22_X1 U4808 ( .A1(n4413), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4416), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3933) );
  AOI22_X1 U4809 ( .A1(n4403), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n4407), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3932) );
  AOI22_X1 U4810 ( .A1(n4414), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4404), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3931) );
  NAND2_X1 U4811 ( .A1(n4412), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3929) );
  AOI21_X1 U4812 ( .B1(n4417), .B2(INSTQUEUE_REG_9__1__SCAN_IN), .A(n4183), 
        .ZN(n3928) );
  AND2_X1 U4813 ( .A1(n3929), .A2(n3928), .ZN(n3930) );
  NAND4_X1 U4814 ( .A1(n3933), .A2(n3932), .A3(n3931), .A4(n3930), .ZN(n3934)
         );
  NAND2_X1 U4815 ( .A1(n4432), .A2(n4435), .ZN(n4094) );
  OAI21_X1 U4816 ( .B1(n3935), .B2(n3934), .A(n4094), .ZN(n3936) );
  AOI22_X1 U4817 ( .A1(n5758), .A2(n4183), .B1(n3937), .B2(n3936), .ZN(n5208)
         );
  NAND2_X1 U4818 ( .A1(n5152), .A2(n5208), .ZN(n5198) );
  INV_X1 U4819 ( .A(n5198), .ZN(n3957) );
  AOI22_X1 U4820 ( .A1(n4414), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4169), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3941) );
  AOI22_X1 U4821 ( .A1(n4416), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3445), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3940) );
  AOI22_X1 U4822 ( .A1(n4403), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4406), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3939) );
  AOI22_X1 U4823 ( .A1(n4415), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3414), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3938) );
  NAND4_X1 U4824 ( .A1(n3941), .A2(n3940), .A3(n3939), .A4(n3938), .ZN(n3947)
         );
  AOI22_X1 U4825 ( .A1(n4405), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4402), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3945) );
  AOI22_X1 U4826 ( .A1(n4418), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3375), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3944) );
  AOI22_X1 U4827 ( .A1(n4412), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4404), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3943) );
  AOI22_X1 U4828 ( .A1(n4413), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4417), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3942) );
  NAND4_X1 U4829 ( .A1(n3945), .A2(n3944), .A3(n3943), .A4(n3942), .ZN(n3946)
         );
  NOR2_X1 U4830 ( .A1(n3947), .A2(n3946), .ZN(n3951) );
  NAND2_X1 U4831 ( .A1(n6443), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3948)
         );
  NAND2_X1 U4832 ( .A1(n4435), .A2(n3948), .ZN(n3949) );
  AOI21_X1 U4833 ( .B1(n4430), .B2(EAX_REG_18__SCAN_IN), .A(n3949), .ZN(n3950)
         );
  OAI21_X1 U4834 ( .B1(n4432), .B2(n3951), .A(n3950), .ZN(n3955) );
  INV_X1 U4835 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5760) );
  OAI21_X1 U4836 ( .B1(PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n3953), .A(n3975), 
        .ZN(n5743) );
  OR2_X1 U4837 ( .A1(n4435), .A2(n5743), .ZN(n3954) );
  NAND2_X1 U4838 ( .A1(n3955), .A2(n3954), .ZN(n5199) );
  NAND2_X1 U4839 ( .A1(n3957), .A2(n3956), .ZN(n5196) );
  AOI22_X1 U4840 ( .A1(n4412), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4405), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3961) );
  AOI22_X1 U4841 ( .A1(n4413), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4418), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3960) );
  AOI22_X1 U4842 ( .A1(n4403), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3375), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3959) );
  AOI22_X1 U4843 ( .A1(n4415), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4404), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3958) );
  NAND4_X1 U4844 ( .A1(n3961), .A2(n3960), .A3(n3959), .A4(n3958), .ZN(n3969)
         );
  AOI22_X1 U4845 ( .A1(n4416), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3401), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3967) );
  AOI22_X1 U4846 ( .A1(n4414), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3414), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3966) );
  AOI22_X1 U4847 ( .A1(n4402), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4406), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3965) );
  NAND2_X1 U4848 ( .A1(n4169), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3963) );
  AOI21_X1 U4849 ( .B1(n4417), .B2(INSTQUEUE_REG_9__3__SCAN_IN), .A(n4183), 
        .ZN(n3962) );
  AND2_X1 U4850 ( .A1(n3963), .A2(n3962), .ZN(n3964) );
  NAND4_X1 U4851 ( .A1(n3967), .A2(n3966), .A3(n3965), .A4(n3964), .ZN(n3968)
         );
  OAI21_X1 U4852 ( .B1(n3969), .B2(n3968), .A(n4094), .ZN(n3971) );
  AOI22_X1 U4853 ( .A1(n4430), .A2(EAX_REG_19__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n6443), .ZN(n3970) );
  NAND2_X1 U4854 ( .A1(n3971), .A2(n3970), .ZN(n3973) );
  XNOR2_X1 U4855 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .B(n3975), .ZN(n5478)
         );
  NAND2_X1 U4856 ( .A1(n5478), .A2(n4183), .ZN(n3972) );
  NAND2_X1 U4857 ( .A1(n3973), .A2(n3972), .ZN(n5306) );
  NOR2_X2 U4858 ( .A1(n5196), .A2(n5306), .ZN(n5290) );
  INV_X1 U4859 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3974) );
  OR2_X1 U4860 ( .A1(n3976), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n3977)
         );
  NAND2_X1 U4861 ( .A1(n3977), .A2(n4095), .ZN(n5616) );
  INV_X1 U4862 ( .A(n5616), .ZN(n3994) );
  INV_X1 U4863 ( .A(n4432), .ZN(n4180) );
  AOI22_X1 U4864 ( .A1(n4403), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4416), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3981) );
  AOI22_X1 U4865 ( .A1(n4402), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4415), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3980) );
  AOI22_X1 U4866 ( .A1(n4418), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n4417), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3979) );
  AOI22_X1 U4867 ( .A1(n4169), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3414), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3978) );
  NAND4_X1 U4868 ( .A1(n3981), .A2(n3980), .A3(n3979), .A4(n3978), .ZN(n3987)
         );
  AOI22_X1 U4869 ( .A1(n4412), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4407), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3985) );
  AOI22_X1 U4870 ( .A1(n4413), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3375), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3984) );
  AOI22_X1 U4871 ( .A1(n4405), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4404), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3983) );
  AOI22_X1 U4872 ( .A1(n4414), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4406), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3982) );
  NAND4_X1 U4873 ( .A1(n3985), .A2(n3984), .A3(n3983), .A4(n3982), .ZN(n3986)
         );
  OR2_X1 U4874 ( .A1(n3987), .A2(n3986), .ZN(n3991) );
  INV_X1 U4875 ( .A(EAX_REG_20__SCAN_IN), .ZN(n3989) );
  NAND2_X1 U4876 ( .A1(n6443), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n3988)
         );
  OAI211_X1 U4877 ( .C1(n4049), .C2(n3989), .A(n4435), .B(n3988), .ZN(n3990)
         );
  AOI21_X1 U4878 ( .B1(n4180), .B2(n3991), .A(n3990), .ZN(n3992) );
  AOI21_X1 U4879 ( .B1(n3994), .B2(n3993), .A(n3992), .ZN(n5289) );
  AND2_X2 U4880 ( .A1(n5290), .A2(n5289), .ZN(n5275) );
  AOI22_X1 U4881 ( .A1(n4416), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4418), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3998) );
  AOI22_X1 U4882 ( .A1(n4413), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4407), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3997) );
  AOI22_X1 U4883 ( .A1(n4403), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3375), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3996) );
  AOI22_X1 U4884 ( .A1(n4402), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4406), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3995) );
  NAND4_X1 U4885 ( .A1(n3998), .A2(n3997), .A3(n3996), .A4(n3995), .ZN(n4004)
         );
  AOI22_X1 U4886 ( .A1(n4169), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n4405), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n4002) );
  AOI22_X1 U4887 ( .A1(n4414), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3414), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4001) );
  AOI22_X1 U4888 ( .A1(n4412), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4404), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4000) );
  AOI22_X1 U4889 ( .A1(n4415), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4417), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3999) );
  NAND4_X1 U4890 ( .A1(n4002), .A2(n4001), .A3(n4000), .A4(n3999), .ZN(n4003)
         );
  NOR2_X1 U4891 ( .A1(n4004), .A2(n4003), .ZN(n4106) );
  AOI22_X1 U4892 ( .A1(n4169), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n4405), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4008) );
  AOI22_X1 U4893 ( .A1(n4413), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4415), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4007) );
  AOI22_X1 U4894 ( .A1(n3375), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n4417), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n4006) );
  AOI22_X1 U4895 ( .A1(n4412), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3414), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4005) );
  NAND4_X1 U4896 ( .A1(n4008), .A2(n4007), .A3(n4006), .A4(n4005), .ZN(n4014)
         );
  AOI22_X1 U4897 ( .A1(n4416), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4418), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4012) );
  AOI22_X1 U4898 ( .A1(n4403), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n4402), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n4011) );
  AOI22_X1 U4899 ( .A1(n4407), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n4406), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4010) );
  AOI22_X1 U4900 ( .A1(n4414), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4404), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4009) );
  NAND4_X1 U4901 ( .A1(n4012), .A2(n4011), .A3(n4010), .A4(n4009), .ZN(n4013)
         );
  NOR2_X1 U4902 ( .A1(n4014), .A2(n4013), .ZN(n4055) );
  AOI22_X1 U4903 ( .A1(INSTQUEUE_REG_2__0__SCAN_IN), .A2(n4169), .B1(n4405), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n4018) );
  AOI22_X1 U4904 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n4416), .B1(n4418), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4017) );
  AOI22_X1 U4905 ( .A1(n4413), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3375), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4016) );
  AOI22_X1 U4906 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n4404), .B1(n3414), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4015) );
  NAND4_X1 U4907 ( .A1(n4018), .A2(n4017), .A3(n4016), .A4(n4015), .ZN(n4024)
         );
  AOI22_X1 U4908 ( .A1(INSTQUEUE_REG_6__0__SCAN_IN), .A2(n4403), .B1(n4407), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4022) );
  AOI22_X1 U4909 ( .A1(n4414), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4402), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n4021) );
  AOI22_X1 U4910 ( .A1(n4412), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4415), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4020) );
  AOI22_X1 U4911 ( .A1(n4406), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n4417), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4019) );
  NAND4_X1 U4912 ( .A1(n4022), .A2(n4021), .A3(n4020), .A4(n4019), .ZN(n4023)
         );
  NOR2_X1 U4913 ( .A1(n4024), .A2(n4023), .ZN(n4054) );
  OR2_X1 U4914 ( .A1(n4055), .A2(n4054), .ZN(n4045) );
  AOI22_X1 U4915 ( .A1(n4416), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4169), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4028) );
  AOI22_X1 U4916 ( .A1(n4414), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4415), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4027) );
  AOI22_X1 U4917 ( .A1(n4412), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3375), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4026) );
  AOI22_X1 U4918 ( .A1(n4413), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3414), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4025) );
  NAND4_X1 U4919 ( .A1(n4028), .A2(n4027), .A3(n4026), .A4(n4025), .ZN(n4034)
         );
  AOI22_X1 U4920 ( .A1(n4405), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4402), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4032) );
  AOI22_X1 U4921 ( .A1(n4407), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n4404), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4031) );
  AOI22_X1 U4922 ( .A1(n4403), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4417), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n4030) );
  AOI22_X1 U4923 ( .A1(n4418), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n4406), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4029) );
  NAND4_X1 U4924 ( .A1(n4032), .A2(n4031), .A3(n4030), .A4(n4029), .ZN(n4033)
         );
  OR2_X1 U4925 ( .A1(n4034), .A2(n4033), .ZN(n4044) );
  INV_X1 U4926 ( .A(n4044), .ZN(n4035) );
  OR2_X1 U4927 ( .A1(n4045), .A2(n4035), .ZN(n4105) );
  XOR2_X1 U4928 ( .A(n4106), .B(n4105), .Z(n4036) );
  NAND2_X1 U4929 ( .A1(n4036), .A2(n4180), .ZN(n4042) );
  NAND2_X1 U4930 ( .A1(n6443), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4037)
         );
  NAND2_X1 U4931 ( .A1(n4435), .A2(n4037), .ZN(n4038) );
  AOI21_X1 U4932 ( .B1(n4430), .B2(EAX_REG_25__SCAN_IN), .A(n4038), .ZN(n4041)
         );
  INV_X1 U4933 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n4039) );
  XNOR2_X1 U4934 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .B(n4102), .ZN(n5566)
         );
  AND2_X1 U4935 ( .A1(n5566), .A2(n4183), .ZN(n4040) );
  AOI21_X1 U4936 ( .B1(n4042), .B2(n4041), .A(n4040), .ZN(n5346) );
  XNOR2_X1 U4937 ( .A(n4043), .B(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5575)
         );
  NAND2_X1 U4938 ( .A1(n5575), .A2(n4183), .ZN(n4053) );
  XNOR2_X1 U4939 ( .A(n4045), .B(n4044), .ZN(n4051) );
  INV_X1 U4940 ( .A(EAX_REG_24__SCAN_IN), .ZN(n4048) );
  INV_X1 U4941 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4046) );
  OAI22_X1 U4942 ( .A1(n4049), .A2(n4048), .B1(n4047), .B2(n4046), .ZN(n4050)
         );
  AOI21_X1 U4943 ( .B1(n4051), .B2(n4180), .A(n4050), .ZN(n4052) );
  AND2_X1 U4944 ( .A1(n4053), .A2(n4052), .ZN(n5354) );
  INV_X1 U4945 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5462) );
  XNOR2_X1 U4946 ( .A(n4063), .B(n5462), .ZN(n5466) );
  NAND2_X1 U4947 ( .A1(n5466), .A2(n4183), .ZN(n4062) );
  XOR2_X1 U4948 ( .A(n4055), .B(n4054), .Z(n4056) );
  NAND2_X1 U4949 ( .A1(n4056), .A2(n4180), .ZN(n4060) );
  NAND2_X1 U4950 ( .A1(n6443), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4057)
         );
  NAND2_X1 U4951 ( .A1(n4435), .A2(n4057), .ZN(n4058) );
  AOI21_X1 U4952 ( .B1(n4430), .B2(EAX_REG_23__SCAN_IN), .A(n4058), .ZN(n4059)
         );
  NAND2_X1 U4953 ( .A1(n4060), .A2(n4059), .ZN(n4061) );
  NAND2_X1 U4954 ( .A1(n4062), .A2(n4061), .ZN(n5276) );
  INV_X1 U4955 ( .A(n4063), .ZN(n4066) );
  OR2_X1 U4956 ( .A1(n4064), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4065)
         );
  NAND2_X1 U4957 ( .A1(n4066), .A2(n4065), .ZN(n5610) );
  AOI22_X1 U4958 ( .A1(n4414), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4405), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4070) );
  AOI22_X1 U4959 ( .A1(n4416), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4418), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4069) );
  AOI22_X1 U4960 ( .A1(n4415), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3375), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4068) );
  AOI22_X1 U4961 ( .A1(n4407), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4406), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4067) );
  NAND4_X1 U4962 ( .A1(n4070), .A2(n4069), .A3(n4068), .A4(n4067), .ZN(n4076)
         );
  AOI22_X1 U4963 ( .A1(n4403), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4412), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4074) );
  AOI22_X1 U4964 ( .A1(n4413), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3414), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4073) );
  AOI22_X1 U4965 ( .A1(n4169), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n4404), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4072) );
  AOI22_X1 U4966 ( .A1(n4402), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4417), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n4071) );
  NAND4_X1 U4967 ( .A1(n4074), .A2(n4073), .A3(n4072), .A4(n4071), .ZN(n4075)
         );
  NOR2_X1 U4968 ( .A1(n4076), .A2(n4075), .ZN(n4079) );
  OAI21_X1 U4969 ( .B1(PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n6852), .A(n6443), 
        .ZN(n4078) );
  NAND2_X1 U4970 ( .A1(n4430), .A2(EAX_REG_22__SCAN_IN), .ZN(n4077) );
  OAI211_X1 U4971 ( .C1(n4432), .C2(n4079), .A(n4078), .B(n4077), .ZN(n4080)
         );
  OAI21_X1 U4972 ( .B1(n5610), .B2(n4435), .A(n4080), .ZN(n5366) );
  OR2_X1 U4973 ( .A1(n5276), .A2(n5366), .ZN(n5277) );
  NOR2_X1 U4974 ( .A1(n5354), .A2(n5277), .ZN(n5344) );
  AND2_X1 U4975 ( .A1(n5346), .A2(n5344), .ZN(n4099) );
  AOI22_X1 U4976 ( .A1(n4414), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4405), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4086) );
  AOI22_X1 U4977 ( .A1(n4413), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3445), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4085) );
  AOI22_X1 U4978 ( .A1(n4402), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3375), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4084) );
  NAND2_X1 U4979 ( .A1(n4412), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4082) );
  AOI21_X1 U4980 ( .B1(n4417), .B2(INSTQUEUE_REG_9__5__SCAN_IN), .A(n4183), 
        .ZN(n4081) );
  AND2_X1 U4981 ( .A1(n4082), .A2(n4081), .ZN(n4083) );
  NAND4_X1 U4982 ( .A1(n4086), .A2(n4085), .A3(n4084), .A4(n4083), .ZN(n4092)
         );
  AOI22_X1 U4983 ( .A1(n4416), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4418), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4090) );
  AOI22_X1 U4984 ( .A1(n4415), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3414), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4089) );
  AOI22_X1 U4985 ( .A1(n4169), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n4404), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4088) );
  AOI22_X1 U4986 ( .A1(n4403), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4406), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4087) );
  NAND4_X1 U4987 ( .A1(n4090), .A2(n4089), .A3(n4088), .A4(n4087), .ZN(n4091)
         );
  OR2_X1 U4988 ( .A1(n4092), .A2(n4091), .ZN(n4093) );
  NAND2_X1 U4989 ( .A1(n4094), .A2(n4093), .ZN(n4098) );
  AOI22_X1 U4990 ( .A1(n4430), .A2(EAX_REG_21__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n6443), .ZN(n4097) );
  XNOR2_X1 U4991 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .B(n4095), .ZN(n5592)
         );
  AND2_X1 U4992 ( .A1(n5592), .A2(n4183), .ZN(n4096) );
  AOI21_X1 U4993 ( .B1(n4098), .B2(n4097), .A(n4096), .ZN(n5368) );
  AND2_X1 U4994 ( .A1(n4099), .A2(n5368), .ZN(n4100) );
  NAND2_X1 U4995 ( .A1(n5275), .A2(n4100), .ZN(n5332) );
  INV_X1 U4996 ( .A(n5332), .ZN(n4123) );
  INV_X1 U4997 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4101) );
  OR2_X1 U4998 ( .A1(n4103), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4104)
         );
  NAND2_X1 U4999 ( .A1(n4103), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4161)
         );
  NAND2_X1 U5000 ( .A1(n4104), .A2(n4161), .ZN(n5604) );
  NOR2_X1 U5001 ( .A1(n4106), .A2(n4105), .ZN(n4125) );
  AOI22_X1 U5002 ( .A1(n4416), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4407), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4110) );
  AOI22_X1 U5003 ( .A1(n4413), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4402), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4109) );
  AOI22_X1 U5004 ( .A1(n4418), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n4417), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4108) );
  AOI22_X1 U5005 ( .A1(n3375), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4406), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4107) );
  NAND4_X1 U5006 ( .A1(n4110), .A2(n4109), .A3(n4108), .A4(n4107), .ZN(n4116)
         );
  AOI22_X1 U5007 ( .A1(n4169), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n4405), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n4114) );
  AOI22_X1 U5008 ( .A1(n4403), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4415), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4113) );
  AOI22_X1 U5009 ( .A1(n4414), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3414), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4112) );
  AOI22_X1 U5010 ( .A1(n4412), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4404), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4111) );
  NAND4_X1 U5011 ( .A1(n4114), .A2(n4113), .A3(n4112), .A4(n4111), .ZN(n4115)
         );
  OR2_X1 U5012 ( .A1(n4116), .A2(n4115), .ZN(n4124) );
  XNOR2_X1 U5013 ( .A(n4125), .B(n4124), .ZN(n4120) );
  NAND2_X1 U5014 ( .A1(n6443), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4117)
         );
  NAND2_X1 U5015 ( .A1(n4435), .A2(n4117), .ZN(n4118) );
  AOI21_X1 U5016 ( .B1(n4430), .B2(EAX_REG_26__SCAN_IN), .A(n4118), .ZN(n4119)
         );
  OAI21_X1 U5017 ( .B1(n4120), .B2(n4432), .A(n4119), .ZN(n4121) );
  OAI21_X1 U5018 ( .B1(n5604), .B2(n4435), .A(n4121), .ZN(n5336) );
  NAND2_X1 U5019 ( .A1(n4123), .A2(n4122), .ZN(n5266) );
  INV_X1 U5020 ( .A(n5266), .ZN(n4144) );
  NAND2_X1 U5021 ( .A1(n4125), .A2(n4124), .ZN(n4145) );
  AOI22_X1 U5022 ( .A1(n4413), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4418), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4129) );
  AOI22_X1 U5023 ( .A1(n4412), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4169), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4128) );
  AOI22_X1 U5024 ( .A1(n4403), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n4407), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4127) );
  AOI22_X1 U5025 ( .A1(n4405), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3412), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4126) );
  NAND4_X1 U5026 ( .A1(n4129), .A2(n4128), .A3(n4127), .A4(n4126), .ZN(n4135)
         );
  AOI22_X1 U5027 ( .A1(n4414), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4415), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4133) );
  AOI22_X1 U5028 ( .A1(n4416), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3414), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4132) );
  AOI22_X1 U5029 ( .A1(n4402), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4404), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4131) );
  AOI22_X1 U5030 ( .A1(n4406), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n4417), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4130) );
  NAND4_X1 U5031 ( .A1(n4133), .A2(n4132), .A3(n4131), .A4(n4130), .ZN(n4134)
         );
  NOR2_X1 U5032 ( .A1(n4135), .A2(n4134), .ZN(n4146) );
  XOR2_X1 U5033 ( .A(n4145), .B(n4146), .Z(n4136) );
  NAND2_X1 U5034 ( .A1(n4136), .A2(n4180), .ZN(n4140) );
  NAND2_X1 U5035 ( .A1(n6443), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4137)
         );
  NAND2_X1 U5036 ( .A1(n4435), .A2(n4137), .ZN(n4138) );
  AOI21_X1 U5037 ( .B1(n4430), .B2(EAX_REG_27__SCAN_IN), .A(n4138), .ZN(n4139)
         );
  NAND2_X1 U5038 ( .A1(n4140), .A2(n4139), .ZN(n4142) );
  XNOR2_X1 U5039 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .B(n4161), .ZN(n5271)
         );
  NAND2_X1 U5040 ( .A1(n4183), .A2(n5271), .ZN(n4141) );
  NAND2_X1 U5041 ( .A1(n4142), .A2(n4141), .ZN(n5268) );
  NAND2_X1 U5042 ( .A1(n4144), .A2(n4143), .ZN(n5320) );
  NOR2_X1 U5043 ( .A1(n4146), .A2(n4145), .ZN(n4168) );
  AOI22_X1 U5044 ( .A1(n4416), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3401), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4150) );
  AOI22_X1 U5045 ( .A1(n4413), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4402), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4149) );
  AOI22_X1 U5046 ( .A1(n4418), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n4417), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4148) );
  AOI22_X1 U5047 ( .A1(n3375), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n4406), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4147) );
  NAND4_X1 U5048 ( .A1(n4150), .A2(n4149), .A3(n4148), .A4(n4147), .ZN(n4156)
         );
  AOI22_X1 U5049 ( .A1(n4169), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n4405), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n4154) );
  AOI22_X1 U5050 ( .A1(n4403), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4415), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4153) );
  AOI22_X1 U5051 ( .A1(n4414), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3414), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4152) );
  AOI22_X1 U5052 ( .A1(n4412), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4404), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4151) );
  NAND4_X1 U5053 ( .A1(n4154), .A2(n4153), .A3(n4152), .A4(n4151), .ZN(n4155)
         );
  OR2_X1 U5054 ( .A1(n4156), .A2(n4155), .ZN(n4167) );
  XNOR2_X1 U5055 ( .A(n4168), .B(n4167), .ZN(n4160) );
  NAND2_X1 U5056 ( .A1(n6443), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4157)
         );
  NAND2_X1 U5057 ( .A1(n4435), .A2(n4157), .ZN(n4158) );
  AOI21_X1 U5058 ( .B1(n4430), .B2(EAX_REG_28__SCAN_IN), .A(n4158), .ZN(n4159)
         );
  OAI21_X1 U5059 ( .B1(n4160), .B2(n4432), .A(n4159), .ZN(n4166) );
  INV_X1 U5060 ( .A(n4161), .ZN(n4162) );
  NOR2_X1 U5061 ( .A1(n4163), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4164)
         );
  NOR2_X1 U5062 ( .A1(n4434), .A2(n4164), .ZN(n5432) );
  NAND2_X1 U5063 ( .A1(n5432), .A2(n4183), .ZN(n4165) );
  NAND2_X1 U5064 ( .A1(n4166), .A2(n4165), .ZN(n5319) );
  NAND2_X1 U5065 ( .A1(n4168), .A2(n4167), .ZN(n4425) );
  AOI22_X1 U5066 ( .A1(n4169), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n4405), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n4173) );
  AOI22_X1 U5067 ( .A1(n4402), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3412), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4172) );
  AOI22_X1 U5068 ( .A1(n4404), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3414), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4171) );
  AOI22_X1 U5069 ( .A1(n3401), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4406), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4170) );
  NAND4_X1 U5070 ( .A1(n4173), .A2(n4172), .A3(n4171), .A4(n4170), .ZN(n4179)
         );
  AOI22_X1 U5071 ( .A1(n4403), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4416), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n4177) );
  AOI22_X1 U5072 ( .A1(n4413), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4414), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4176) );
  AOI22_X1 U5073 ( .A1(n4412), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4415), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4175) );
  AOI22_X1 U5074 ( .A1(n4418), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n4417), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4174) );
  NAND4_X1 U5075 ( .A1(n4177), .A2(n4176), .A3(n4175), .A4(n4174), .ZN(n4178)
         );
  NOR2_X1 U5076 ( .A1(n4179), .A2(n4178), .ZN(n4426) );
  XOR2_X1 U5077 ( .A(n4425), .B(n4426), .Z(n4181) );
  NAND2_X1 U5078 ( .A1(n4181), .A2(n4180), .ZN(n4185) );
  INV_X1 U5079 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4192) );
  NOR2_X1 U5080 ( .A1(n4192), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4182) );
  AOI211_X1 U5081 ( .C1(n4430), .C2(EAX_REG_29__SCAN_IN), .A(n4183), .B(n4182), 
        .ZN(n4184) );
  XOR2_X1 U5082 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .B(n4434), .Z(n5236) );
  AOI22_X1 U5083 ( .A1(n4185), .A2(n4184), .B1(n4183), .B2(n5236), .ZN(n4186)
         );
  NAND2_X1 U5084 ( .A1(n5245), .A2(n4187), .ZN(n5228) );
  NAND3_X1 U5085 ( .A1(n6544), .A2(STATEBS16_REG_SCAN_IN), .A3(
        STATE2_REG_1__SCAN_IN), .ZN(n6556) );
  INV_X1 U5086 ( .A(n6556), .ZN(n4188) );
  NOR2_X2 U5087 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6405) );
  NAND2_X1 U5088 ( .A1(n4188), .A2(n6405), .ZN(n6447) );
  INV_X1 U5089 ( .A(n6405), .ZN(n6643) );
  AOI21_X1 U5090 ( .B1(n6643), .B2(n6644), .A(STATE2_REG_0__SCAN_IN), .ZN(
        n4189) );
  NAND2_X1 U5091 ( .A1(n6544), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4191) );
  NAND2_X1 U5092 ( .A1(n6852), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4190) );
  NAND2_X1 U5093 ( .A1(n4191), .A2(n4190), .ZN(n6011) );
  NOR2_X1 U5094 ( .A1(STATE2_REG_0__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6558) );
  INV_X1 U5095 ( .A(n6558), .ZN(n6549) );
  OR2_X1 U5096 ( .A1(n6634), .A2(n6549), .ZN(n6015) );
  INV_X2 U5097 ( .A(n6015), .ZN(n6054) );
  NAND2_X1 U5098 ( .A1(n6054), .A2(REIP_REG_29__SCAN_IN), .ZN(n5496) );
  OAI21_X1 U5099 ( .B1(n5989), .B2(n4192), .A(n5496), .ZN(n4193) );
  AOI21_X1 U5100 ( .B1(n5983), .B2(n5236), .A(n4193), .ZN(n4194) );
  OAI211_X1 U5101 ( .C1(n5501), .C2(n5972), .A(n3189), .B(n4194), .ZN(U2957)
         );
  NAND2_X1 U5102 ( .A1(n4195), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5419) );
  INV_X1 U5103 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5421) );
  NOR2_X1 U5104 ( .A1(n4198), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5418)
         );
  NAND2_X1 U5105 ( .A1(n5418), .A2(n5421), .ZN(n4199) );
  OAI22_X2 U5106 ( .A1(n5419), .A2(n5421), .B1(n4197), .B2(n4199), .ZN(n4200)
         );
  XNOR2_X1 U5107 ( .A(n4200), .B(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4473)
         );
  NAND2_X1 U5108 ( .A1(n4201), .A2(n4770), .ZN(n4202) );
  NOR2_X1 U5109 ( .A1(n4203), .A2(n4202), .ZN(n4484) );
  INV_X1 U5110 ( .A(n4484), .ZN(n4480) );
  NAND2_X1 U5111 ( .A1(n4204), .A2(n5907), .ZN(n4206) );
  MUX2_X1 U5112 ( .A(n4206), .B(n6649), .S(n4205), .Z(n4232) );
  NAND2_X1 U5113 ( .A1(n4232), .A2(n4225), .ZN(n4207) );
  NAND2_X1 U5114 ( .A1(n4480), .A2(n4207), .ZN(n4231) );
  NAND2_X1 U5115 ( .A1(n6622), .A2(n4274), .ZN(n4208) );
  OR2_X1 U5116 ( .A1(n4570), .A2(n4208), .ZN(n4209) );
  NAND2_X1 U5117 ( .A1(n4231), .A2(n4209), .ZN(n4508) );
  OR2_X1 U5118 ( .A1(n4210), .A2(STATE_REG_0__SCAN_IN), .ZN(n6566) );
  NAND2_X1 U5119 ( .A1(n4274), .A2(n6566), .ZN(n4217) );
  AND2_X1 U5120 ( .A1(n4212), .A2(n4211), .ZN(n4213) );
  AND2_X1 U5121 ( .A1(n4214), .A2(n4213), .ZN(n4215) );
  OR2_X1 U5122 ( .A1(n4216), .A2(n4215), .ZN(n4440) );
  NOR2_X1 U5123 ( .A1(READY_N), .A2(n4440), .ZN(n4505) );
  AND3_X1 U5124 ( .A1(n4217), .A2(n4505), .A3(n4235), .ZN(n4218) );
  OAI21_X1 U5125 ( .B1(n4508), .B2(n4218), .A(n6537), .ZN(n4223) );
  NAND2_X1 U5126 ( .A1(n3162), .A2(n6566), .ZN(n4447) );
  INV_X1 U5127 ( .A(n4447), .ZN(n4220) );
  OR3_X1 U5128 ( .A1(n4521), .A2(n4220), .A3(READY_N), .ZN(n4509) );
  NAND3_X1 U5129 ( .A1(n4509), .A2(n3170), .A3(n4236), .ZN(n4221) );
  NAND3_X1 U5130 ( .A1(n5546), .A2(n4680), .A3(n4221), .ZN(n4222) );
  NOR2_X1 U5131 ( .A1(n4380), .A2(n4765), .ZN(n4224) );
  NOR2_X1 U5132 ( .A1(n6526), .A2(n4224), .ZN(n4227) );
  AND2_X1 U5133 ( .A1(n4225), .A2(n4610), .ZN(n4504) );
  INV_X1 U5134 ( .A(n4504), .ZN(n4534) );
  OR2_X1 U5135 ( .A1(n4510), .A2(n3162), .ZN(n4226) );
  AND4_X1 U5136 ( .A1(n4227), .A2(n4519), .A3(n4534), .A4(n4226), .ZN(n4228)
         );
  NAND2_X1 U5137 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5099) );
  NOR2_X1 U5138 ( .A1(n5095), .A2(n5099), .ZN(n5103) );
  NAND2_X1 U5139 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n5103), .ZN(n5179) );
  NAND2_X1 U5140 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5183) );
  NOR2_X1 U5141 ( .A1(n5179), .A2(n5183), .ZN(n4258) );
  NOR2_X1 U5142 ( .A1(n4229), .A2(n4770), .ZN(n4230) );
  NAND2_X1 U5143 ( .A1(n4231), .A2(n4230), .ZN(n4571) );
  NOR2_X1 U5144 ( .A1(n4879), .A2(n4878), .ZN(n4914) );
  NAND3_X1 U5145 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A3(n4914), .ZN(n5060) );
  AOI21_X1 U5146 ( .B1(INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .A(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n6047) );
  NAND2_X1 U5147 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6036) );
  NOR2_X1 U5148 ( .A1(n6047), .A2(n6036), .ZN(n4757) );
  NAND3_X1 U5149 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_6__SCAN_IN), .A3(n4757), .ZN(n4877) );
  NOR2_X1 U5150 ( .A1(n5060), .A2(n4877), .ZN(n4251) );
  NAND2_X1 U5151 ( .A1(n6048), .A2(n4251), .ZN(n5098) );
  NAND2_X1 U5152 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4711) );
  NOR2_X1 U5153 ( .A1(n4711), .A2(n6036), .ZN(n4761) );
  NAND3_X1 U5154 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_6__SCAN_IN), .A3(n4761), .ZN(n4872) );
  NOR2_X1 U5155 ( .A1(n4872), .A2(n5060), .ZN(n5094) );
  INV_X1 U5156 ( .A(n4638), .ZN(n4244) );
  INV_X1 U5157 ( .A(n4232), .ZN(n4241) );
  NAND2_X1 U5158 ( .A1(n4770), .A2(n4274), .ZN(n5007) );
  NOR2_X1 U5159 ( .A1(n5007), .A2(n4235), .ZN(n4512) );
  OAI21_X1 U5160 ( .B1(n4512), .B2(n3175), .A(n4234), .ZN(n4238) );
  NAND2_X1 U5161 ( .A1(n4236), .A2(n4235), .ZN(n4237) );
  OAI211_X1 U5162 ( .C1(n4239), .C2(n4376), .A(n4238), .B(n4237), .ZN(n4240)
         );
  NOR2_X1 U5163 ( .A1(n4241), .A2(n4240), .ZN(n4242) );
  NAND2_X1 U5164 ( .A1(n4243), .A2(n4242), .ZN(n4523) );
  AOI211_X1 U5165 ( .C1(n4246), .C2(n4245), .A(n4244), .B(n4523), .ZN(n4247)
         );
  NOR2_X1 U5166 ( .A1(n4384), .A2(n4247), .ZN(n4257) );
  NAND2_X1 U5167 ( .A1(n4257), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5097)
         );
  NAND2_X1 U5168 ( .A1(n4484), .A2(n4274), .ZN(n6511) );
  NAND2_X1 U5169 ( .A1(n5097), .A2(n6064), .ZN(n6049) );
  NAND2_X1 U5170 ( .A1(n5094), .A2(n6049), .ZN(n5063) );
  NAND2_X1 U5171 ( .A1(n5098), .A2(n5063), .ZN(n5697) );
  NAND2_X1 U5172 ( .A1(n4258), .A2(n5697), .ZN(n5689) );
  INV_X1 U5173 ( .A(n4252), .ZN(n4248) );
  NAND2_X1 U5174 ( .A1(n5674), .A2(n5667), .ZN(n5661) );
  NOR2_X1 U5175 ( .A1(n5661), .A2(n4249), .ZN(n4395) );
  OR2_X1 U5176 ( .A1(n4257), .A2(n6048), .ZN(n5100) );
  INV_X1 U5177 ( .A(n5100), .ZN(n4250) );
  NAND2_X1 U5178 ( .A1(n4250), .A2(n6064), .ZN(n5664) );
  NAND2_X1 U5179 ( .A1(n4258), .A2(n4251), .ZN(n5663) );
  INV_X1 U5180 ( .A(n5663), .ZN(n4253) );
  NAND3_X1 U5181 ( .A1(n4253), .A2(n5667), .A3(n4252), .ZN(n4254) );
  AND2_X1 U5182 ( .A1(n5664), .A2(n4254), .ZN(n4259) );
  INV_X1 U5183 ( .A(n6064), .ZN(n4255) );
  NOR2_X1 U5184 ( .A1(n4257), .A2(n4255), .ZN(n4871) );
  INV_X1 U5185 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6065) );
  NAND2_X1 U5186 ( .A1(n4384), .A2(n6015), .ZN(n6063) );
  INV_X1 U5187 ( .A(n6063), .ZN(n4256) );
  AOI21_X1 U5188 ( .B1(n6065), .B2(n4257), .A(n4256), .ZN(n4875) );
  OAI221_X1 U5189 ( .B1(n5094), .B2(n4871), .C1(n4258), .C2(n4871), .A(n4875), 
        .ZN(n5662) );
  OR2_X1 U5190 ( .A1(n4259), .A2(n5662), .ZN(n5655) );
  OR2_X1 U5191 ( .A1(n4395), .A2(n5655), .ZN(n5537) );
  OAI21_X1 U5192 ( .B1(n6049), .B2(n6048), .A(n4260), .ZN(n4261) );
  INV_X1 U5193 ( .A(n4261), .ZN(n4262) );
  NOR2_X1 U5194 ( .A1(n5537), .A2(n4262), .ZN(n5654) );
  INV_X1 U5195 ( .A(n5664), .ZN(n5181) );
  NAND2_X1 U5196 ( .A1(n5654), .A2(n5181), .ZN(n4267) );
  NAND2_X1 U5197 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5518) );
  INV_X1 U5198 ( .A(n5518), .ZN(n4263) );
  NAND2_X1 U5199 ( .A1(n5654), .A2(n4263), .ZN(n4264) );
  AND2_X1 U5200 ( .A1(n4267), .A2(n4264), .ZN(n5645) );
  AND2_X1 U5201 ( .A1(n4267), .A2(n4269), .ZN(n4265) );
  NOR2_X1 U5202 ( .A1(n5645), .A2(n4265), .ZN(n5492) );
  INV_X1 U5203 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5494) );
  AOI21_X1 U5204 ( .B1(n5664), .B2(n5494), .A(n5421), .ZN(n4266) );
  NAND2_X1 U5205 ( .A1(n5492), .A2(n4266), .ZN(n5487) );
  NAND3_X1 U5206 ( .A1(n5487), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .A3(n4267), .ZN(n4273) );
  NAND2_X1 U5207 ( .A1(n6054), .A2(REIP_REG_31__SCAN_IN), .ZN(n4471) );
  AND2_X1 U5208 ( .A1(n5674), .A2(n4268), .ZN(n5648) );
  NAND3_X1 U5209 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .A3(n5648), .ZN(n5504) );
  INV_X1 U5210 ( .A(n4269), .ZN(n5502) );
  NAND2_X1 U5211 ( .A1(n5502), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4270) );
  NOR2_X1 U5212 ( .A1(n5504), .A2(n4270), .ZN(n5488) );
  INV_X1 U5213 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4271) );
  NAND3_X1 U5214 ( .A1(n5488), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(n4271), .ZN(n4272) );
  AND3_X1 U5215 ( .A1(n4273), .A2(n4471), .A3(n4272), .ZN(n4386) );
  NAND2_X2 U5216 ( .A1(n4276), .A2(n4275), .ZN(n4279) );
  INV_X1 U5217 ( .A(n3177), .ZN(n4277) );
  INV_X1 U5218 ( .A(EBX_REG_0__SCAN_IN), .ZN(n4278) );
  OAI22_X1 U5219 ( .A1(n4292), .A2(n4278), .B1(n4233), .B2(EBX_REG_0__SCAN_IN), 
        .ZN(n4603) );
  XNOR2_X1 U5220 ( .A(n4279), .B(n4603), .ZN(n4573) );
  AOI21_X2 U5221 ( .B1(n4573), .B2(n3178), .A(n4279), .ZN(n5028) );
  INV_X1 U5222 ( .A(EBX_REG_2__SCAN_IN), .ZN(n5891) );
  NAND2_X1 U5223 ( .A1(n4346), .A2(n5891), .ZN(n4283) );
  NAND2_X1 U5224 ( .A1(n4376), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4281)
         );
  OAI211_X1 U5225 ( .C1(n4293), .C2(EBX_REG_2__SCAN_IN), .A(n3177), .B(n4281), 
        .ZN(n4282) );
  INV_X1 U5226 ( .A(EBX_REG_3__SCAN_IN), .ZN(n5861) );
  NAND2_X1 U5227 ( .A1(n4367), .A2(n5861), .ZN(n4287) );
  INV_X1 U5228 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4717) );
  NAND2_X1 U5229 ( .A1(n3177), .A2(n4717), .ZN(n4285) );
  NAND2_X1 U5230 ( .A1(n3178), .A2(n5861), .ZN(n4284) );
  NAND3_X1 U5231 ( .A1(n4285), .A2(n4376), .A3(n4284), .ZN(n4286) );
  AND2_X1 U5232 ( .A1(n4287), .A2(n4286), .ZN(n4627) );
  NAND2_X1 U5233 ( .A1(n4376), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4290)
         );
  OAI211_X1 U5234 ( .C1(n4293), .C2(EBX_REG_4__SCAN_IN), .A(n3177), .B(n4290), 
        .ZN(n4291) );
  OAI21_X1 U5235 ( .B1(n4359), .B2(EBX_REG_4__SCAN_IN), .A(n4291), .ZN(n4739)
         );
  MUX2_X1 U5236 ( .A(n4361), .B(n3177), .S(EBX_REG_5__SCAN_IN), .Z(n4296) );
  NAND2_X1 U5237 ( .A1(n4277), .A2(n4293), .ZN(n4343) );
  NAND2_X1 U5238 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n4293), .ZN(n4294)
         );
  AND2_X1 U5239 ( .A1(n4343), .A2(n4294), .ZN(n4295) );
  NAND2_X1 U5240 ( .A1(n4296), .A2(n4295), .ZN(n4756) );
  AND2_X2 U5241 ( .A1(n4738), .A2(n4756), .ZN(n4755) );
  MUX2_X1 U5242 ( .A(n4359), .B(n4376), .S(EBX_REG_6__SCAN_IN), .Z(n4297) );
  OAI21_X1 U5243 ( .B1(INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n3175), .A(n4297), 
        .ZN(n4787) );
  INV_X1 U5244 ( .A(n4787), .ZN(n4298) );
  INV_X1 U5245 ( .A(EBX_REG_7__SCAN_IN), .ZN(n5813) );
  NAND2_X1 U5246 ( .A1(n4367), .A2(n5813), .ZN(n4302) );
  NAND2_X1 U5247 ( .A1(n3177), .A2(n4879), .ZN(n4300) );
  NAND2_X1 U5248 ( .A1(n3178), .A2(n5813), .ZN(n4299) );
  NAND3_X1 U5249 ( .A1(n4300), .A2(n4376), .A3(n4299), .ZN(n4301) );
  AND2_X1 U5250 ( .A1(n4302), .A2(n4301), .ZN(n4819) );
  MUX2_X1 U5251 ( .A(n4359), .B(n4376), .S(EBX_REG_8__SCAN_IN), .Z(n4304) );
  OAI21_X1 U5252 ( .B1(INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n3175), .A(n4304), 
        .ZN(n4882) );
  OR2_X1 U5253 ( .A1(n4361), .A2(EBX_REG_9__SCAN_IN), .ZN(n4308) );
  NAND2_X1 U5254 ( .A1(n3177), .A2(n6017), .ZN(n4306) );
  INV_X1 U5255 ( .A(EBX_REG_9__SCAN_IN), .ZN(n4969) );
  NAND2_X1 U5256 ( .A1(n3178), .A2(n4969), .ZN(n4305) );
  NAND3_X1 U5257 ( .A1(n4306), .A2(n4376), .A3(n4305), .ZN(n4307) );
  NAND2_X1 U5258 ( .A1(n4308), .A2(n4307), .ZN(n4910) );
  INV_X1 U5259 ( .A(EBX_REG_10__SCAN_IN), .ZN(n4997) );
  NAND2_X1 U5260 ( .A1(n4346), .A2(n4997), .ZN(n4311) );
  NAND2_X1 U5261 ( .A1(n4376), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n4309) );
  OAI211_X1 U5262 ( .C1(n4293), .C2(EBX_REG_10__SCAN_IN), .A(n3177), .B(n4309), 
        .ZN(n4310) );
  AND2_X1 U5263 ( .A1(n4311), .A2(n4310), .ZN(n4922) );
  MUX2_X1 U5264 ( .A(n4361), .B(n3177), .S(EBX_REG_11__SCAN_IN), .Z(n4313) );
  NAND2_X1 U5265 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n4293), .ZN(n4312) );
  AND3_X1 U5266 ( .A1(n4313), .A2(n4343), .A3(n4312), .ZN(n4975) );
  NAND2_X1 U5267 ( .A1(n4376), .A2(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n4314) );
  OAI211_X1 U5268 ( .C1(n4293), .C2(EBX_REG_12__SCAN_IN), .A(n3177), .B(n4314), 
        .ZN(n4315) );
  OAI21_X1 U5269 ( .B1(n4359), .B2(EBX_REG_12__SCAN_IN), .A(n4315), .ZN(n4961)
         );
  MUX2_X1 U5270 ( .A(n4361), .B(n3177), .S(EBX_REG_13__SCAN_IN), .Z(n4317) );
  NAND2_X1 U5271 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n4293), .ZN(n4316) );
  AND3_X1 U5272 ( .A1(n4317), .A2(n4343), .A3(n4316), .ZN(n5050) );
  INV_X1 U5273 ( .A(EBX_REG_14__SCAN_IN), .ZN(n5129) );
  NAND2_X1 U5274 ( .A1(n4346), .A2(n5129), .ZN(n4320) );
  NAND2_X1 U5275 ( .A1(n4376), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n4318) );
  OAI211_X1 U5276 ( .C1(n4293), .C2(EBX_REG_14__SCAN_IN), .A(n3177), .B(n4318), 
        .ZN(n4319) );
  AND2_X1 U5277 ( .A1(n4320), .A2(n4319), .ZN(n5105) );
  NAND2_X2 U5278 ( .A1(n5106), .A2(n5105), .ZN(n5104) );
  MUX2_X1 U5279 ( .A(n4361), .B(n3177), .S(EBX_REG_15__SCAN_IN), .Z(n4323) );
  NAND2_X1 U5280 ( .A1(n4293), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n4321) );
  AND2_X1 U5281 ( .A1(n4343), .A2(n4321), .ZN(n4322) );
  NAND2_X1 U5282 ( .A1(n4323), .A2(n4322), .ZN(n5146) );
  INV_X1 U5283 ( .A(EBX_REG_16__SCAN_IN), .ZN(n5167) );
  NAND2_X1 U5284 ( .A1(n4346), .A2(n5167), .ZN(n4326) );
  NAND2_X1 U5285 ( .A1(n4376), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n4324) );
  OAI211_X1 U5286 ( .C1(n4293), .C2(EBX_REG_16__SCAN_IN), .A(n3177), .B(n4324), 
        .ZN(n4325) );
  AND2_X1 U5287 ( .A1(n4326), .A2(n4325), .ZN(n5154) );
  NAND2_X1 U5288 ( .A1(n5146), .A2(n5154), .ZN(n4327) );
  MUX2_X1 U5289 ( .A(n4361), .B(n3177), .S(EBX_REG_17__SCAN_IN), .Z(n4329) );
  NAND2_X1 U5290 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n4293), .ZN(n4328) );
  AND3_X1 U5291 ( .A1(n4329), .A2(n4343), .A3(n4328), .ZN(n5210) );
  NOR2_X4 U5292 ( .A1(n5209), .A2(n5210), .ZN(n5217) );
  INV_X1 U5293 ( .A(EBX_REG_19__SCAN_IN), .ZN(n5312) );
  NAND2_X1 U5294 ( .A1(n4346), .A2(n5312), .ZN(n4332) );
  NAND2_X1 U5295 ( .A1(n4376), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n4330) );
  OAI211_X1 U5296 ( .C1(n4293), .C2(EBX_REG_19__SCAN_IN), .A(n3177), .B(n4330), 
        .ZN(n4331) );
  AND2_X1 U5297 ( .A1(n4332), .A2(n4331), .ZN(n5307) );
  OR2_X1 U5298 ( .A1(n3175), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n4334)
         );
  INV_X1 U5299 ( .A(EBX_REG_20__SCAN_IN), .ZN(n5376) );
  NAND2_X1 U5300 ( .A1(n3178), .A2(n5376), .ZN(n4333) );
  NAND2_X1 U5301 ( .A1(n4334), .A2(n4333), .ZN(n5299) );
  OR2_X1 U5302 ( .A1(n3175), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4335)
         );
  INV_X1 U5303 ( .A(EBX_REG_18__SCAN_IN), .ZN(n5220) );
  NAND2_X1 U5304 ( .A1(n3178), .A2(n5220), .ZN(n5214) );
  AND2_X1 U5305 ( .A1(n4335), .A2(n5214), .ZN(n5297) );
  NAND2_X1 U5306 ( .A1(n5297), .A2(n5299), .ZN(n4338) );
  INV_X1 U5307 ( .A(n5297), .ZN(n4336) );
  NAND2_X1 U5308 ( .A1(n4336), .A2(n4376), .ZN(n4337) );
  OAI211_X1 U5309 ( .C1(n5299), .C2(n4376), .A(n4338), .B(n4337), .ZN(n4339)
         );
  INV_X1 U5310 ( .A(n4339), .ZN(n4340) );
  NAND2_X1 U5311 ( .A1(n5296), .A2(n4340), .ZN(n5372) );
  MUX2_X1 U5312 ( .A(n4359), .B(n4376), .S(EBX_REG_21__SCAN_IN), .Z(n4341) );
  OAI21_X1 U5313 ( .B1(INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n3175), .A(n4341), 
        .ZN(n5371) );
  OR2_X2 U5314 ( .A1(n5372), .A2(n5371), .ZN(n5374) );
  MUX2_X1 U5315 ( .A(n4361), .B(n3177), .S(EBX_REG_22__SCAN_IN), .Z(n4345) );
  NAND2_X1 U5316 ( .A1(n4293), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4342) );
  AND2_X1 U5317 ( .A1(n4343), .A2(n4342), .ZN(n4344) );
  NAND2_X1 U5318 ( .A1(n4345), .A2(n4344), .ZN(n5281) );
  INV_X1 U5319 ( .A(EBX_REG_23__SCAN_IN), .ZN(n5360) );
  NAND2_X1 U5320 ( .A1(n4346), .A2(n5360), .ZN(n4349) );
  NAND2_X1 U5321 ( .A1(n4376), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4347) );
  OAI211_X1 U5322 ( .C1(n4293), .C2(EBX_REG_23__SCAN_IN), .A(n3177), .B(n4347), 
        .ZN(n4348) );
  AND2_X1 U5323 ( .A1(n4349), .A2(n4348), .ZN(n5280) );
  NAND2_X1 U5324 ( .A1(n5281), .A2(n5280), .ZN(n4350) );
  MUX2_X1 U5325 ( .A(n4361), .B(n3177), .S(EBX_REG_24__SCAN_IN), .Z(n4352) );
  NAND2_X1 U5326 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n4293), .ZN(n4351) );
  NAND2_X1 U5327 ( .A1(n4352), .A2(n4351), .ZN(n5355) );
  MUX2_X1 U5328 ( .A(n4359), .B(n4376), .S(EBX_REG_25__SCAN_IN), .Z(n4354) );
  OR2_X1 U5329 ( .A1(n3175), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n4353)
         );
  AND2_X1 U5330 ( .A1(n4354), .A2(n4353), .ZN(n5348) );
  INV_X1 U5331 ( .A(EBX_REG_26__SCAN_IN), .ZN(n5341) );
  NAND2_X1 U5332 ( .A1(n4367), .A2(n5341), .ZN(n4358) );
  INV_X1 U5333 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5521) );
  NAND2_X1 U5334 ( .A1(n3177), .A2(n5521), .ZN(n4356) );
  NAND2_X1 U5335 ( .A1(n3178), .A2(n5341), .ZN(n4355) );
  NAND3_X1 U5336 ( .A1(n4356), .A2(n4376), .A3(n4355), .ZN(n4357) );
  AND2_X1 U5337 ( .A1(n4358), .A2(n4357), .ZN(n5338) );
  MUX2_X1 U5338 ( .A(n4359), .B(n4376), .S(EBX_REG_27__SCAN_IN), .Z(n4360) );
  OAI21_X1 U5339 ( .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n3175), .A(n4360), 
        .ZN(n5270) );
  OR2_X1 U5340 ( .A1(n4361), .A2(EBX_REG_28__SCAN_IN), .ZN(n4366) );
  INV_X1 U5341 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4362) );
  NAND2_X1 U5342 ( .A1(n3177), .A2(n4362), .ZN(n4364) );
  INV_X1 U5343 ( .A(EBX_REG_28__SCAN_IN), .ZN(n5327) );
  NAND2_X1 U5344 ( .A1(n3178), .A2(n5327), .ZN(n4363) );
  NAND3_X1 U5345 ( .A1(n4364), .A2(n4376), .A3(n4363), .ZN(n4365) );
  NAND2_X1 U5346 ( .A1(n4366), .A2(n4365), .ZN(n5323) );
  INV_X1 U5347 ( .A(n5326), .ZN(n5247) );
  INV_X1 U5348 ( .A(EBX_REG_29__SCAN_IN), .ZN(n4368) );
  AND2_X1 U5349 ( .A1(n4367), .A2(n4368), .ZN(n5230) );
  NAND2_X1 U5350 ( .A1(n5247), .A2(n5230), .ZN(n4374) );
  OR2_X1 U5351 ( .A1(n3175), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4370)
         );
  NAND2_X1 U5352 ( .A1(n3178), .A2(n4368), .ZN(n4369) );
  NAND2_X1 U5353 ( .A1(n4370), .A2(n4369), .ZN(n5229) );
  OR2_X2 U5354 ( .A1(n4371), .A2(n5229), .ZN(n5253) );
  INV_X1 U5355 ( .A(n4233), .ZN(n5298) );
  NOR2_X2 U5356 ( .A1(n5253), .A2(n5298), .ZN(n4372) );
  INV_X1 U5357 ( .A(n4372), .ZN(n4373) );
  AND2_X1 U5358 ( .A1(n4293), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4375)
         );
  AOI21_X1 U5359 ( .B1(n3175), .B2(EBX_REG_30__SCAN_IN), .A(n4375), .ZN(n5252)
         );
  NAND2_X1 U5360 ( .A1(n5232), .A2(n5252), .ZN(n4377) );
  NAND2_X1 U5361 ( .A1(n5253), .A2(n4376), .ZN(n5250) );
  OAI22_X1 U5362 ( .A1(n3175), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        EBX_REG_31__SCAN_IN), .B2(n4293), .ZN(n4378) );
  OR2_X1 U5364 ( .A1(n4521), .A2(n6649), .ZN(n6540) );
  INV_X1 U5365 ( .A(n4380), .ZN(n4381) );
  NAND2_X1 U5366 ( .A1(n4381), .A2(n4765), .ZN(n4382) );
  AND2_X1 U5367 ( .A1(n6540), .A2(n4382), .ZN(n4383) );
  XNOR2_X1 U5368 ( .A(n5092), .B(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5476)
         );
  NAND2_X1 U5369 ( .A1(n5477), .A2(n5476), .ZN(n5475) );
  INV_X1 U5370 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5680) );
  NAND2_X1 U5371 ( .A1(n5612), .A2(n3183), .ZN(n4391) );
  INV_X1 U5372 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5673) );
  XNOR2_X1 U5373 ( .A(n4388), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5470)
         );
  INV_X1 U5374 ( .A(n4393), .ZN(n5454) );
  XNOR2_X1 U5375 ( .A(n5452), .B(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4394)
         );
  XNOR2_X1 U5376 ( .A(n5454), .B(n4394), .ZN(n5607) );
  NAND2_X1 U5377 ( .A1(n5607), .A2(n6060), .ZN(n4401) );
  XNOR2_X1 U5378 ( .A(n5374), .B(n5281), .ZN(n5588) );
  AOI21_X1 U5379 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n5655), .A(n4395), 
        .ZN(n4398) );
  NAND2_X1 U5380 ( .A1(n6054), .A2(REIP_REG_22__SCAN_IN), .ZN(n4396) );
  NAND2_X1 U5381 ( .A1(n4401), .A2(n4400), .ZN(U2996) );
  AOI22_X1 U5382 ( .A1(n4403), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4402), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4411) );
  AOI22_X1 U5383 ( .A1(n3412), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3414), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4410) );
  AOI22_X1 U5384 ( .A1(n4405), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4404), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4409) );
  AOI22_X1 U5385 ( .A1(n4407), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n4406), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4408) );
  NAND4_X1 U5386 ( .A1(n4411), .A2(n4410), .A3(n4409), .A4(n4408), .ZN(n4424)
         );
  AOI22_X1 U5387 ( .A1(n4413), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4412), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4422) );
  AOI22_X1 U5388 ( .A1(n4414), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4169), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4421) );
  AOI22_X1 U5389 ( .A1(n4416), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4415), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4420) );
  AOI22_X1 U5390 ( .A1(n4418), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n4417), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4419) );
  NAND4_X1 U5391 ( .A1(n4422), .A2(n4421), .A3(n4420), .A4(n4419), .ZN(n4423)
         );
  NOR2_X1 U5392 ( .A1(n4424), .A2(n4423), .ZN(n4428) );
  NOR2_X1 U5393 ( .A1(n4426), .A2(n4425), .ZN(n4427) );
  XOR2_X1 U5394 ( .A(n4428), .B(n4427), .Z(n4433) );
  INV_X1 U5395 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5257) );
  OAI21_X1 U5396 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5257), .A(n4435), .ZN(
        n4429) );
  AOI21_X1 U5397 ( .B1(n4430), .B2(EAX_REG_30__SCAN_IN), .A(n4429), .ZN(n4431)
         );
  OAI21_X1 U5398 ( .B1(n4433), .B2(n4432), .A(n4431), .ZN(n4437) );
  NAND2_X1 U5399 ( .A1(n4434), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4442)
         );
  XNOR2_X1 U5400 ( .A(n4442), .B(n5257), .ZN(n5416) );
  OR2_X1 U5401 ( .A1(n5416), .A2(n4435), .ZN(n4436) );
  NAND2_X1 U5402 ( .A1(n4437), .A2(n4436), .ZN(n5244) );
  AOI22_X1 U5403 ( .A1(n4430), .A2(EAX_REG_31__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n3790), .ZN(n4438) );
  INV_X1 U5404 ( .A(n4510), .ZN(n4479) );
  INV_X1 U5405 ( .A(n4440), .ZN(n4485) );
  NAND3_X1 U5406 ( .A1(n4485), .A2(n6537), .A3(n4484), .ZN(n4476) );
  NAND2_X1 U5407 ( .A1(n4495), .A2(n4476), .ZN(n6647) );
  NOR3_X1 U5408 ( .A1(STATEBS16_REG_SCAN_IN), .A2(n6549), .A3(n4656), .ZN(
        n6552) );
  NAND2_X1 U5409 ( .A1(n4656), .A2(n6443), .ZN(n6650) );
  NOR3_X1 U5410 ( .A1(n6615), .A2(n6544), .A3(n6650), .ZN(n6542) );
  OR3_X1 U5411 ( .A1(n6552), .A2(n6542), .A3(n6054), .ZN(n4441) );
  NOR2_X1 U5412 ( .A1(n4442), .A2(n5257), .ZN(n4443) );
  XNOR2_X1 U5413 ( .A(n4443), .B(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4991)
         );
  NOR2_X1 U5414 ( .A1(n4991), .A2(n4656), .ZN(n4444) );
  NAND2_X1 U5415 ( .A1(n5383), .A2(n5804), .ZN(n4469) );
  INV_X1 U5416 ( .A(EBX_REG_31__SCAN_IN), .ZN(n4445) );
  NOR2_X1 U5417 ( .A1(n5008), .A2(n4445), .ZN(n4453) );
  NOR2_X1 U5418 ( .A1(READY_N), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4983) );
  NOR2_X1 U5419 ( .A1(n4293), .A2(n4983), .ZN(n4446) );
  NAND3_X1 U5420 ( .A1(n4447), .A2(n4983), .A3(n5907), .ZN(n4448) );
  INV_X1 U5421 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6811) );
  AND2_X1 U5422 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n4462) );
  INV_X1 U5423 ( .A(REIP_REG_23__SCAN_IN), .ZN(n6842) );
  INV_X1 U5424 ( .A(REIP_REG_22__SCAN_IN), .ZN(n6871) );
  INV_X1 U5425 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6972) );
  NOR3_X1 U5426 ( .A1(n6842), .A2(n6871), .A3(n6972), .ZN(n4450) );
  NAND3_X1 U5427 ( .A1(REIP_REG_20__SCAN_IN), .A2(REIP_REG_19__SCAN_IN), .A3(
        REIP_REG_18__SCAN_IN), .ZN(n4460) );
  INV_X1 U5428 ( .A(REIP_REG_15__SCAN_IN), .ZN(n6596) );
  NAND3_X1 U5429 ( .A1(REIP_REG_14__SCAN_IN), .A2(REIP_REG_13__SCAN_IN), .A3(
        REIP_REG_12__SCAN_IN), .ZN(n5144) );
  NOR2_X1 U5430 ( .A1(n6596), .A2(n5144), .ZN(n4458) );
  INV_X1 U5431 ( .A(n5820), .ZN(n5844) );
  INV_X1 U5432 ( .A(REIP_REG_8__SCAN_IN), .ZN(n6586) );
  INV_X1 U5433 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6583) );
  INV_X1 U5434 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6581) );
  NAND3_X1 U5435 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_3__SCAN_IN), .A3(
        REIP_REG_2__SCAN_IN), .ZN(n5850) );
  NOR2_X1 U5436 ( .A1(n6581), .A2(n5850), .ZN(n5822) );
  NAND2_X1 U5437 ( .A1(REIP_REG_5__SCAN_IN), .A2(n5822), .ZN(n5819) );
  NOR2_X1 U5438 ( .A1(n6583), .A2(n5819), .ZN(n5810) );
  NAND2_X1 U5439 ( .A1(REIP_REG_7__SCAN_IN), .A2(n5810), .ZN(n5795) );
  NOR2_X1 U5440 ( .A1(n6586), .A2(n5795), .ZN(n5796) );
  NAND2_X1 U5441 ( .A1(REIP_REG_9__SCAN_IN), .A2(n5796), .ZN(n4457) );
  NAND2_X1 U5442 ( .A1(REIP_REG_11__SCAN_IN), .A2(REIP_REG_10__SCAN_IN), .ZN(
        n4449) );
  NOR3_X1 U5443 ( .A1(n5844), .A2(n4457), .A3(n4449), .ZN(n5125) );
  NAND4_X1 U5444 ( .A1(n4458), .A2(REIP_REG_17__SCAN_IN), .A3(
        REIP_REG_16__SCAN_IN), .A4(n5125), .ZN(n5309) );
  NOR2_X1 U5445 ( .A1(n4460), .A2(n5309), .ZN(n5295) );
  NOR2_X1 U5446 ( .A1(n5844), .A2(n5845), .ZN(n5876) );
  AOI21_X1 U5447 ( .B1(n4450), .B2(n5295), .A(n5876), .ZN(n5577) );
  NAND3_X1 U5448 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_26__SCAN_IN), .A3(
        REIP_REG_25__SCAN_IN), .ZN(n4461) );
  INV_X1 U5449 ( .A(n4461), .ZN(n4451) );
  NOR2_X1 U5450 ( .A1(n5851), .A2(n4451), .ZN(n4452) );
  NOR2_X1 U5451 ( .A1(n5577), .A2(n4452), .ZN(n5560) );
  OAI21_X1 U5452 ( .B1(n4462), .B2(n5851), .A(n5560), .ZN(n5235) );
  AOI21_X1 U5453 ( .B1(n5845), .B2(n6811), .A(n5235), .ZN(n5256) );
  OAI21_X1 U5454 ( .B1(REIP_REG_30__SCAN_IN), .B2(n5851), .A(n5256), .ZN(n4465) );
  INV_X1 U5455 ( .A(n4453), .ZN(n4456) );
  INV_X1 U5456 ( .A(n6566), .ZN(n4454) );
  NAND2_X1 U5457 ( .A1(n4454), .A2(n4983), .ZN(n6541) );
  NAND2_X1 U5458 ( .A1(n4490), .A2(n6541), .ZN(n4986) );
  INV_X1 U5459 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4455) );
  OAI22_X1 U5460 ( .A1(n4456), .A2(n4986), .B1(n4455), .B2(n5886), .ZN(n4464)
         );
  NAND3_X1 U5461 ( .A1(n5776), .A2(REIP_REG_11__SCAN_IN), .A3(
        REIP_REG_10__SCAN_IN), .ZN(n5766) );
  INV_X1 U5462 ( .A(n4458), .ZN(n4459) );
  NOR2_X1 U5463 ( .A1(n5766), .A2(n4459), .ZN(n5755) );
  NAND3_X1 U5464 ( .A1(n5755), .A2(REIP_REG_17__SCAN_IN), .A3(
        REIP_REG_16__SCAN_IN), .ZN(n5749) );
  NOR2_X1 U5465 ( .A1(n5749), .A2(n4460), .ZN(n5595) );
  NAND4_X1 U5466 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .A4(n5595), .ZN(n5569) );
  NOR2_X1 U5467 ( .A1(n5569), .A2(n4461), .ZN(n5555) );
  NAND2_X1 U5468 ( .A1(n5555), .A2(n4462), .ZN(n5265) );
  INV_X1 U5469 ( .A(REIP_REG_30__SCAN_IN), .ZN(n5415) );
  NOR4_X1 U5470 ( .A1(n5265), .A2(REIP_REG_31__SCAN_IN), .A3(n5415), .A4(n6811), .ZN(n4463) );
  AOI211_X1 U5471 ( .C1(REIP_REG_31__SCAN_IN), .C2(n4465), .A(n4464), .B(n4463), .ZN(n4466) );
  NAND2_X1 U5472 ( .A1(n4469), .A2(n4468), .ZN(U2796) );
  NAND2_X1 U5473 ( .A1(n6012), .A2(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4470)
         );
  OAI211_X1 U5474 ( .C1(n6005), .C2(n4991), .A(n4471), .B(n4470), .ZN(n4472)
         );
  AOI21_X1 U5475 ( .B1(n5383), .B2(n3167), .A(n4472), .ZN(n4475) );
  OR2_X2 U5476 ( .A1(n4473), .A2(n5972), .ZN(n4474) );
  NAND2_X1 U5477 ( .A1(n4475), .A2(n4474), .ZN(U2955) );
  INV_X1 U5478 ( .A(n4476), .ZN(n4478) );
  INV_X1 U5479 ( .A(MEMORYFETCH_REG_SCAN_IN), .ZN(n6656) );
  AND2_X1 U5480 ( .A1(n6405), .A2(n4656), .ZN(n4988) );
  INV_X1 U5481 ( .A(n4988), .ZN(n4477) );
  OAI211_X1 U5482 ( .C1(n4478), .C2(n6656), .A(n4495), .B(n4477), .ZN(U2788)
         );
  INV_X1 U5483 ( .A(n4571), .ZN(n4483) );
  NOR3_X1 U5484 ( .A1(n6526), .A2(n4504), .A3(n4479), .ZN(n4481) );
  OAI22_X1 U5485 ( .A1(n4481), .A2(n4570), .B1(n4485), .B2(n4480), .ZN(n4482)
         );
  AOI21_X1 U5486 ( .B1(n4483), .B2(n4570), .A(n4482), .ZN(n6530) );
  NAND2_X1 U5487 ( .A1(n4485), .A2(n4484), .ZN(n4486) );
  NAND2_X1 U5488 ( .A1(n4486), .A2(n4510), .ZN(n4488) );
  OR2_X1 U5489 ( .A1(n4570), .A2(n4610), .ZN(n4487) );
  NAND2_X1 U5490 ( .A1(n4488), .A2(n4487), .ZN(n5723) );
  INV_X1 U5491 ( .A(n5007), .ZN(n4489) );
  OR2_X1 U5492 ( .A1(n4490), .A2(n4489), .ZN(n4493) );
  AOI21_X1 U5493 ( .B1(n4493), .B2(n6566), .A(READY_N), .ZN(n6648) );
  NOR2_X1 U5494 ( .A1(n5723), .A2(n6648), .ZN(n6527) );
  OR2_X1 U5495 ( .A1(n6527), .A2(n6550), .ZN(n5727) );
  NAND2_X1 U5496 ( .A1(n5727), .A2(MORE_REG_SCAN_IN), .ZN(n4491) );
  OAI21_X1 U5497 ( .B1(n6530), .B2(n5727), .A(n4491), .ZN(U3471) );
  INV_X1 U5498 ( .A(n6647), .ZN(n4494) );
  OAI21_X1 U5499 ( .B1(n4988), .B2(READREQUEST_REG_SCAN_IN), .A(n4494), .ZN(
        n4492) );
  OAI21_X1 U5500 ( .B1(n4494), .B2(n4493), .A(n4492), .ZN(U3474) );
  INV_X1 U5501 ( .A(LWORD_REG_15__SCAN_IN), .ZN(n4499) );
  INV_X1 U5502 ( .A(n6540), .ZN(n4496) );
  NAND2_X1 U5503 ( .A1(n5546), .A2(n4496), .ZN(n4501) );
  NAND2_X1 U5504 ( .A1(n4497), .A2(n4501), .ZN(n4500) );
  INV_X1 U5505 ( .A(DATAI_15_), .ZN(n6993) );
  INV_X1 U5506 ( .A(EAX_REG_15__SCAN_IN), .ZN(n4498) );
  OAI222_X1 U5507 ( .A1(n4499), .A2(n4500), .B1(n4615), .B2(n6993), .C1(n4498), 
        .C2(n4501), .ZN(U2954) );
  AOI22_X1 U5508 ( .A1(n4575), .A2(LWORD_REG_12__SCAN_IN), .B1(
        EAX_REG_12__SCAN_IN), .B2(n4600), .ZN(n4503) );
  INV_X1 U5509 ( .A(DATAI_12_), .ZN(n4502) );
  OR2_X1 U5510 ( .A1(n4615), .A2(n4502), .ZN(n4563) );
  NAND2_X1 U5511 ( .A1(n4503), .A2(n4563), .ZN(U2951) );
  NAND2_X1 U5512 ( .A1(n6544), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6613) );
  NAND2_X1 U5513 ( .A1(n4570), .A2(n4504), .ZN(n4507) );
  INV_X1 U5514 ( .A(n4519), .ZN(n4654) );
  NAND2_X1 U5515 ( .A1(n4654), .A2(n4505), .ZN(n4506) );
  NAND2_X1 U5516 ( .A1(n4507), .A2(n4506), .ZN(n4613) );
  NOR2_X1 U5517 ( .A1(n4508), .A2(n4613), .ZN(n4516) );
  OAI21_X1 U5518 ( .B1(n6511), .B2(READY_N), .A(n4509), .ZN(n4514) );
  NAND2_X1 U5519 ( .A1(n4510), .A2(n6566), .ZN(n4511) );
  AND2_X1 U5520 ( .A1(n4570), .A2(n4511), .ZN(n4513) );
  AOI21_X1 U5521 ( .B1(n4514), .B2(n4513), .A(n4512), .ZN(n4515) );
  NAND2_X1 U5522 ( .A1(n4516), .A2(n4515), .ZN(n6515) );
  NAND2_X1 U5523 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), 
        .ZN(n5545) );
  NOR2_X1 U5524 ( .A1(n6544), .A2(n5545), .ZN(n4659) );
  AOI22_X1 U5525 ( .A1(n6515), .A2(n6537), .B1(FLUSH_REG_SCAN_IN), .B2(n4659), 
        .ZN(n5718) );
  NAND2_X1 U5526 ( .A1(n6613), .A2(n5718), .ZN(n6629) );
  INV_X1 U5527 ( .A(n6629), .ZN(n6631) );
  INV_X1 U5528 ( .A(n6071), .ZN(n5009) );
  NAND4_X1 U5529 ( .A1(n4521), .A2(n4520), .A3(n4519), .A4(n4518), .ZN(n4522)
         );
  NOR2_X1 U5530 ( .A1(n4523), .A2(n4522), .ZN(n6623) );
  INV_X1 U5531 ( .A(n6623), .ZN(n4644) );
  NAND2_X1 U5532 ( .A1(n5009), .A2(n4644), .ZN(n4527) );
  CLKBUF_X1 U5533 ( .A(n4524), .Z(n4632) );
  INV_X1 U5534 ( .A(n4632), .ZN(n4531) );
  INV_X1 U5535 ( .A(n4525), .ZN(n4651) );
  NAND3_X1 U5536 ( .A1(n6622), .A2(n4531), .A3(n4651), .ZN(n4526) );
  OAI211_X1 U5537 ( .C1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C2(n6511), .A(n4527), .B(n4526), .ZN(n6514) );
  INV_X1 U5538 ( .A(n6634), .ZN(n6621) );
  NOR2_X1 U5539 ( .A1(n4656), .A2(n6065), .ZN(n6627) );
  INV_X1 U5540 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4696) );
  AOI22_X1 U5541 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B1(n4271), .B2(n4696), .ZN(n4542)
         );
  INV_X1 U5542 ( .A(n4542), .ZN(n4528) );
  NOR2_X1 U5543 ( .A1(n4632), .A2(n6617), .ZN(n4543) );
  AOI222_X1 U5544 ( .A1(n6514), .A2(n6621), .B1(n6627), .B2(n4528), .C1(n4651), 
        .C2(n4543), .ZN(n4530) );
  NAND2_X1 U5545 ( .A1(n6631), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4529) );
  OAI21_X1 U5546 ( .B1(n6631), .B2(n4530), .A(n4529), .ZN(U3460) );
  NOR3_X1 U5547 ( .A1(n4531), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n6617), 
        .ZN(n4541) );
  NAND2_X1 U5548 ( .A1(n4571), .A2(n4534), .ZN(n4635) );
  XNOR2_X1 U5549 ( .A(n4632), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4537)
         );
  XNOR2_X1 U5550 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4535) );
  OAI22_X1 U5551 ( .A1(n6511), .A2(n4535), .B1(n4638), .B2(n4537), .ZN(n4536)
         );
  AOI21_X1 U5552 ( .B1(n4635), .B2(n4537), .A(n4536), .ZN(n4538) );
  OAI21_X1 U5553 ( .B1(n4533), .B2(n6623), .A(n4538), .ZN(n4646) );
  INV_X1 U5554 ( .A(n4646), .ZN(n4539) );
  NOR2_X1 U5555 ( .A1(n4539), .A2(n6634), .ZN(n4540) );
  AOI211_X1 U5556 ( .C1(n6627), .C2(n4542), .A(n4541), .B(n4540), .ZN(n4545)
         );
  OAI21_X1 U5557 ( .B1(n6631), .B2(n4543), .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), 
        .ZN(n4544) );
  OAI21_X1 U5558 ( .B1(n4545), .B2(n6631), .A(n4544), .ZN(U3459) );
  AOI22_X1 U5559 ( .A1(n4575), .A2(LWORD_REG_13__SCAN_IN), .B1(
        EAX_REG_13__SCAN_IN), .B2(n4600), .ZN(n4546) );
  NAND2_X1 U5560 ( .A1(n4576), .A2(DATAI_13_), .ZN(n4560) );
  NAND2_X1 U5561 ( .A1(n4546), .A2(n4560), .ZN(U2952) );
  AOI22_X1 U5562 ( .A1(n4575), .A2(LWORD_REG_4__SCAN_IN), .B1(n4600), .B2(
        EAX_REG_4__SCAN_IN), .ZN(n4547) );
  NAND2_X1 U5563 ( .A1(n4576), .A2(DATAI_4_), .ZN(n4598) );
  NAND2_X1 U5564 ( .A1(n4547), .A2(n4598), .ZN(U2943) );
  AOI22_X1 U5565 ( .A1(n4575), .A2(LWORD_REG_5__SCAN_IN), .B1(
        EAX_REG_5__SCAN_IN), .B2(n4600), .ZN(n4548) );
  NAND2_X1 U5566 ( .A1(n4576), .A2(DATAI_5_), .ZN(n4596) );
  NAND2_X1 U5567 ( .A1(n4548), .A2(n4596), .ZN(U2944) );
  AOI22_X1 U5568 ( .A1(n4575), .A2(LWORD_REG_8__SCAN_IN), .B1(
        EAX_REG_8__SCAN_IN), .B2(n4600), .ZN(n4549) );
  NAND2_X1 U5569 ( .A1(n4576), .A2(DATAI_8_), .ZN(n4592) );
  NAND2_X1 U5570 ( .A1(n4549), .A2(n4592), .ZN(U2947) );
  AOI22_X1 U5571 ( .A1(n4575), .A2(LWORD_REG_7__SCAN_IN), .B1(
        EAX_REG_7__SCAN_IN), .B2(n4600), .ZN(n4550) );
  NAND2_X1 U5572 ( .A1(n4576), .A2(DATAI_7_), .ZN(n4594) );
  NAND2_X1 U5573 ( .A1(n4550), .A2(n4594), .ZN(U2946) );
  AOI22_X1 U5574 ( .A1(n4575), .A2(LWORD_REG_9__SCAN_IN), .B1(
        EAX_REG_9__SCAN_IN), .B2(n4600), .ZN(n4551) );
  NAND2_X1 U5575 ( .A1(n4576), .A2(DATAI_9_), .ZN(n4584) );
  NAND2_X1 U5576 ( .A1(n4551), .A2(n4584), .ZN(U2948) );
  AOI22_X1 U5577 ( .A1(n4575), .A2(LWORD_REG_11__SCAN_IN), .B1(
        EAX_REG_11__SCAN_IN), .B2(n4600), .ZN(n4552) );
  NAND2_X1 U5578 ( .A1(n4576), .A2(DATAI_11_), .ZN(n4586) );
  NAND2_X1 U5579 ( .A1(n4552), .A2(n4586), .ZN(U2950) );
  AOI22_X1 U5580 ( .A1(n4575), .A2(LWORD_REG_6__SCAN_IN), .B1(
        EAX_REG_6__SCAN_IN), .B2(n4600), .ZN(n4553) );
  NAND2_X1 U5581 ( .A1(n4576), .A2(DATAI_6_), .ZN(n4601) );
  NAND2_X1 U5582 ( .A1(n4553), .A2(n4601), .ZN(U2945) );
  AOI22_X1 U5583 ( .A1(n4575), .A2(LWORD_REG_3__SCAN_IN), .B1(
        EAX_REG_3__SCAN_IN), .B2(n4600), .ZN(n4554) );
  NAND2_X1 U5584 ( .A1(n4576), .A2(DATAI_3_), .ZN(n4590) );
  NAND2_X1 U5585 ( .A1(n4554), .A2(n4590), .ZN(U2942) );
  AOI22_X1 U5586 ( .A1(n4575), .A2(LWORD_REG_10__SCAN_IN), .B1(
        EAX_REG_10__SCAN_IN), .B2(n4600), .ZN(n4555) );
  NAND2_X1 U5587 ( .A1(n4576), .A2(DATAI_10_), .ZN(n4588) );
  NAND2_X1 U5588 ( .A1(n4555), .A2(n4588), .ZN(U2949) );
  AOI22_X1 U5589 ( .A1(n4575), .A2(LWORD_REG_2__SCAN_IN), .B1(
        EAX_REG_2__SCAN_IN), .B2(n4600), .ZN(n4556) );
  NAND2_X1 U5590 ( .A1(n4576), .A2(DATAI_2_), .ZN(n4582) );
  NAND2_X1 U5591 ( .A1(n4556), .A2(n4582), .ZN(U2941) );
  AOI22_X1 U5592 ( .A1(n4575), .A2(UWORD_REG_14__SCAN_IN), .B1(
        EAX_REG_30__SCAN_IN), .B2(n4600), .ZN(n4557) );
  NAND2_X1 U5593 ( .A1(n4576), .A2(DATAI_14_), .ZN(n4558) );
  NAND2_X1 U5594 ( .A1(n4557), .A2(n4558), .ZN(U2938) );
  AOI22_X1 U5595 ( .A1(n4575), .A2(LWORD_REG_14__SCAN_IN), .B1(
        EAX_REG_14__SCAN_IN), .B2(n4600), .ZN(n4559) );
  NAND2_X1 U5596 ( .A1(n4559), .A2(n4558), .ZN(U2953) );
  AOI22_X1 U5597 ( .A1(n4575), .A2(UWORD_REG_13__SCAN_IN), .B1(
        EAX_REG_29__SCAN_IN), .B2(n4600), .ZN(n4561) );
  NAND2_X1 U5598 ( .A1(n4561), .A2(n4560), .ZN(U2937) );
  AOI22_X1 U5599 ( .A1(n4575), .A2(LWORD_REG_0__SCAN_IN), .B1(
        EAX_REG_0__SCAN_IN), .B2(n4600), .ZN(n4562) );
  NAND2_X1 U5600 ( .A1(n4576), .A2(DATAI_0_), .ZN(n4578) );
  NAND2_X1 U5601 ( .A1(n4562), .A2(n4578), .ZN(U2939) );
  AOI22_X1 U5602 ( .A1(n4575), .A2(UWORD_REG_12__SCAN_IN), .B1(
        EAX_REG_28__SCAN_IN), .B2(n4600), .ZN(n4564) );
  NAND2_X1 U5603 ( .A1(n4564), .A2(n4563), .ZN(U2936) );
  OAI21_X1 U5604 ( .B1(n4566), .B2(n4565), .A(n4619), .ZN(n6000) );
  NAND4_X1 U5605 ( .A1(n4765), .A2(n5381), .A3(n4675), .A4(n4680), .ZN(n4568)
         );
  NOR2_X1 U5606 ( .A1(n4568), .A2(n4567), .ZN(n4611) );
  NAND2_X1 U5607 ( .A1(n4611), .A2(n3178), .ZN(n4569) );
  OAI21_X1 U5608 ( .B1(n4571), .B2(n4570), .A(n4569), .ZN(n4572) );
  AND2_X1 U5609 ( .A1(n5892), .A2(n5202), .ZN(n5889) );
  NAND2_X1 U5610 ( .A1(n5892), .A2(n5381), .ZN(n5378) );
  XNOR2_X1 U5611 ( .A(n4573), .B(n3178), .ZN(n4700) );
  INV_X1 U5612 ( .A(n5892), .ZN(n5379) );
  AOI22_X1 U5613 ( .A1(n5888), .A2(n4700), .B1(EBX_REG_1__SCAN_IN), .B2(n5379), 
        .ZN(n4574) );
  OAI21_X1 U5614 ( .B1(n6000), .B2(n3166), .A(n4574), .ZN(U2858) );
  AOI22_X1 U5615 ( .A1(n4575), .A2(LWORD_REG_1__SCAN_IN), .B1(
        EAX_REG_1__SCAN_IN), .B2(n4600), .ZN(n4577) );
  NAND2_X1 U5616 ( .A1(n4576), .A2(DATAI_1_), .ZN(n4580) );
  NAND2_X1 U5617 ( .A1(n4577), .A2(n4580), .ZN(U2940) );
  AOI22_X1 U5618 ( .A1(n4575), .A2(UWORD_REG_0__SCAN_IN), .B1(
        EAX_REG_16__SCAN_IN), .B2(n4600), .ZN(n4579) );
  NAND2_X1 U5619 ( .A1(n4579), .A2(n4578), .ZN(U2924) );
  AOI22_X1 U5620 ( .A1(n4575), .A2(UWORD_REG_1__SCAN_IN), .B1(
        EAX_REG_17__SCAN_IN), .B2(n4600), .ZN(n4581) );
  NAND2_X1 U5621 ( .A1(n4581), .A2(n4580), .ZN(U2925) );
  AOI22_X1 U5622 ( .A1(n4575), .A2(UWORD_REG_2__SCAN_IN), .B1(
        EAX_REG_18__SCAN_IN), .B2(n4600), .ZN(n4583) );
  NAND2_X1 U5623 ( .A1(n4583), .A2(n4582), .ZN(U2926) );
  AOI22_X1 U5624 ( .A1(n4575), .A2(UWORD_REG_9__SCAN_IN), .B1(
        EAX_REG_25__SCAN_IN), .B2(n4600), .ZN(n4585) );
  NAND2_X1 U5625 ( .A1(n4585), .A2(n4584), .ZN(U2933) );
  AOI22_X1 U5626 ( .A1(n4575), .A2(UWORD_REG_11__SCAN_IN), .B1(
        EAX_REG_27__SCAN_IN), .B2(n4600), .ZN(n4587) );
  NAND2_X1 U5627 ( .A1(n4587), .A2(n4586), .ZN(U2935) );
  AOI22_X1 U5628 ( .A1(n4575), .A2(UWORD_REG_10__SCAN_IN), .B1(
        EAX_REG_26__SCAN_IN), .B2(n4600), .ZN(n4589) );
  NAND2_X1 U5629 ( .A1(n4589), .A2(n4588), .ZN(U2934) );
  AOI22_X1 U5630 ( .A1(n4575), .A2(UWORD_REG_3__SCAN_IN), .B1(
        EAX_REG_19__SCAN_IN), .B2(n4600), .ZN(n4591) );
  NAND2_X1 U5631 ( .A1(n4591), .A2(n4590), .ZN(U2927) );
  AOI22_X1 U5632 ( .A1(n4575), .A2(UWORD_REG_8__SCAN_IN), .B1(
        EAX_REG_24__SCAN_IN), .B2(n4600), .ZN(n4593) );
  NAND2_X1 U5633 ( .A1(n4593), .A2(n4592), .ZN(U2932) );
  AOI22_X1 U5634 ( .A1(n4575), .A2(UWORD_REG_7__SCAN_IN), .B1(
        EAX_REG_23__SCAN_IN), .B2(n4600), .ZN(n4595) );
  NAND2_X1 U5635 ( .A1(n4595), .A2(n4594), .ZN(U2931) );
  AOI22_X1 U5636 ( .A1(n4575), .A2(UWORD_REG_5__SCAN_IN), .B1(
        EAX_REG_21__SCAN_IN), .B2(n4600), .ZN(n4597) );
  NAND2_X1 U5637 ( .A1(n4597), .A2(n4596), .ZN(U2929) );
  AOI22_X1 U5638 ( .A1(n4575), .A2(UWORD_REG_4__SCAN_IN), .B1(
        EAX_REG_20__SCAN_IN), .B2(n4600), .ZN(n4599) );
  NAND2_X1 U5639 ( .A1(n4599), .A2(n4598), .ZN(U2928) );
  AOI22_X1 U5640 ( .A1(n4575), .A2(UWORD_REG_6__SCAN_IN), .B1(
        EAX_REG_22__SCAN_IN), .B2(n4600), .ZN(n4602) );
  NAND2_X1 U5641 ( .A1(n4602), .A2(n4601), .ZN(U2930) );
  NOR2_X1 U5642 ( .A1(n3175), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4604)
         );
  OR2_X1 U5643 ( .A1(n4604), .A2(n4603), .ZN(n6057) );
  INV_X1 U5644 ( .A(n4605), .ZN(n4607) );
  NAND2_X1 U5645 ( .A1(n4607), .A2(n4606), .ZN(n4609) );
  AND2_X1 U5646 ( .A1(n4609), .A2(n4608), .ZN(n6009) );
  INV_X1 U5647 ( .A(n6009), .ZN(n5906) );
  OAI222_X1 U5648 ( .A1(n6057), .A2(n5378), .B1(n4278), .B2(n5892), .C1(n5906), 
        .C2(n3166), .ZN(U2859) );
  AND2_X1 U5649 ( .A1(n4611), .A2(n4610), .ZN(n4612) );
  OAI21_X1 U5650 ( .B1(n4613), .B2(n4612), .A(n6537), .ZN(n4614) );
  NAND2_X1 U5651 ( .A1(n3316), .A2(n5202), .ZN(n4616) );
  INV_X1 U5652 ( .A(n4616), .ZN(n4617) );
  NAND2_X1 U5653 ( .A1(n5905), .A2(n4617), .ZN(n5904) );
  INV_X1 U5654 ( .A(DATAI_1_), .ZN(n6839) );
  INV_X1 U5655 ( .A(EAX_REG_1__SCAN_IN), .ZN(n5963) );
  OAI222_X1 U5656 ( .A1(n6000), .A2(n5413), .B1(n5904), .B2(n6839), .C1(n5905), 
        .C2(n5963), .ZN(U2890) );
  NAND3_X1 U5657 ( .A1(n4621), .A2(n4620), .A3(n4619), .ZN(n4622) );
  AND2_X1 U5658 ( .A1(n4618), .A2(n4622), .ZN(n5995) );
  INV_X1 U5659 ( .A(n5995), .ZN(n5035) );
  INV_X1 U5660 ( .A(DATAI_2_), .ZN(n4679) );
  INV_X1 U5661 ( .A(EAX_REG_2__SCAN_IN), .ZN(n5961) );
  OAI222_X1 U5662 ( .A1(n5035), .A2(n5413), .B1(n5904), .B2(n4679), .C1(n5905), 
        .C2(n5961), .ZN(U2889) );
  AND2_X1 U5663 ( .A1(n4618), .A2(n4623), .ZN(n4626) );
  CLKBUF_X1 U5664 ( .A(n4624), .Z(n4625) );
  OR2_X1 U5665 ( .A1(n4626), .A2(n4625), .ZN(n4707) );
  NAND2_X1 U5666 ( .A1(n5026), .A2(n4627), .ZN(n4628) );
  NAND2_X1 U5667 ( .A1(n4740), .A2(n4628), .ZN(n4713) );
  INV_X1 U5668 ( .A(n4713), .ZN(n5865) );
  AOI22_X1 U5669 ( .A1(n5888), .A2(n5865), .B1(EBX_REG_3__SCAN_IN), .B2(n5379), 
        .ZN(n4629) );
  OAI21_X1 U5670 ( .B1(n4707), .B2(n3166), .A(n4629), .ZN(U2856) );
  INV_X1 U5671 ( .A(DATAI_3_), .ZN(n6990) );
  INV_X1 U5672 ( .A(EAX_REG_3__SCAN_IN), .ZN(n5959) );
  OAI222_X1 U5673 ( .A1(n4707), .A2(n5413), .B1(n5904), .B2(n6990), .C1(n5905), 
        .C2(n5959), .ZN(U2888) );
  INV_X1 U5674 ( .A(FLUSH_REG_SCAN_IN), .ZN(n5728) );
  NAND2_X1 U5675 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n5728), .ZN(n4650) );
  INV_X1 U5676 ( .A(n4630), .ZN(n4649) );
  INV_X1 U5677 ( .A(n4631), .ZN(n4633) );
  MUX2_X1 U5678 ( .A(n4633), .B(n4645), .S(n4632), .Z(n4634) );
  NAND3_X1 U5679 ( .A1(n4635), .A2(n4649), .A3(n4634), .ZN(n4642) );
  XNOR2_X1 U5680 ( .A(n4636), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4639)
         );
  OAI21_X1 U5681 ( .B1(n4413), .B2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(n4637), 
        .ZN(n6616) );
  OAI22_X1 U5682 ( .A1(n6511), .A2(n4639), .B1(n4638), .B2(n6616), .ZN(n4640)
         );
  INV_X1 U5683 ( .A(n4640), .ZN(n4641) );
  NAND2_X1 U5684 ( .A1(n4642), .A2(n4641), .ZN(n4643) );
  AOI21_X1 U5685 ( .B1(n6257), .B2(n4644), .A(n4643), .ZN(n6618) );
  MUX2_X1 U5686 ( .A(n4645), .B(n6618), .S(n6515), .Z(n6525) );
  INV_X1 U5687 ( .A(n6525), .ZN(n4647) );
  MUX2_X1 U5688 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n4646), .S(n6515), 
        .Z(n6520) );
  NAND3_X1 U5689 ( .A1(n4647), .A2(n6520), .A3(n4656), .ZN(n4648) );
  OAI21_X1 U5690 ( .B1(n4650), .B2(n4649), .A(n4648), .ZN(n6533) );
  NAND2_X1 U5691 ( .A1(n6533), .A2(n4651), .ZN(n4662) );
  INV_X1 U5692 ( .A(n4892), .ZN(n6332) );
  NOR2_X1 U5693 ( .A1(n4652), .A2(n6332), .ZN(n4653) );
  XNOR2_X1 U5694 ( .A(n4653), .B(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n5846)
         );
  NAND2_X1 U5695 ( .A1(n4654), .A2(n4656), .ZN(n4655) );
  NOR2_X1 U5696 ( .A1(n5846), .A2(n4655), .ZN(n5720) );
  MUX2_X1 U5697 ( .A(FLUSH_REG_SCAN_IN), .B(n6515), .S(n4656), .Z(n4657) );
  NOR2_X1 U5698 ( .A1(n4657), .A2(n5722), .ZN(n4658) );
  NOR2_X1 U5699 ( .A1(n5720), .A2(n4658), .ZN(n6531) );
  AND3_X1 U5700 ( .A1(n4662), .A2(n6531), .A3(n5728), .ZN(n4660) );
  INV_X1 U5701 ( .A(n4659), .ZN(n6612) );
  OAI21_X1 U5702 ( .B1(n4660), .B2(n6612), .A(n6227), .ZN(n6066) );
  INV_X1 U5703 ( .A(n5545), .ZN(n4661) );
  AND3_X1 U5704 ( .A1(n4662), .A2(n6531), .A3(n4661), .ZN(n6543) );
  OAI22_X1 U5705 ( .A1(n6409), .A2(n6643), .B1(n6624), .B2(n3184), .ZN(n4663)
         );
  OAI21_X1 U5706 ( .B1(n6543), .B2(n4663), .A(n6066), .ZN(n4664) );
  OAI21_X1 U5707 ( .B1(n6066), .B2(n6509), .A(n4664), .ZN(U3465) );
  INV_X1 U5708 ( .A(n6222), .ZN(n4688) );
  NAND2_X1 U5709 ( .A1(n4666), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5542) );
  OAI21_X1 U5710 ( .B1(n4688), .B2(n5542), .A(n6405), .ZN(n4672) );
  NAND2_X1 U5711 ( .A1(n4533), .A2(n5009), .ZN(n4825) );
  INV_X1 U5712 ( .A(n4825), .ZN(n4667) );
  NAND2_X1 U5713 ( .A1(n4667), .A2(n6257), .ZN(n6296) );
  OR2_X1 U5714 ( .A1(n6296), .A2(n6624), .ZN(n4669) );
  INV_X1 U5715 ( .A(n4668), .ZN(n4826) );
  NAND2_X1 U5716 ( .A1(n4826), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6319) );
  NAND2_X1 U5717 ( .A1(n4669), .A2(n6319), .ZN(n4673) );
  INV_X1 U5718 ( .A(n4673), .ZN(n4670) );
  NAND3_X1 U5719 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n6521), .ZN(n6288) );
  OAI22_X1 U5720 ( .A1(n4672), .A2(n4670), .B1(n6288), .B2(n6443), .ZN(n6323)
         );
  INV_X1 U5721 ( .A(n6323), .ZN(n4815) );
  NOR2_X2 U5722 ( .A1(n6990), .A2(n6227), .ZN(n6472) );
  INV_X1 U5723 ( .A(n6472), .ZN(n4934) );
  OAI21_X1 U5724 ( .B1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n6615), .A(n6135), 
        .ZN(n6451) );
  AOI21_X1 U5725 ( .B1(n6288), .B2(n6643), .A(n6451), .ZN(n4671) );
  OAI21_X1 U5726 ( .B1(n4673), .B2(n4672), .A(n4671), .ZN(n6324) );
  NAND2_X1 U5727 ( .A1(n6324), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n4678)
         );
  AND2_X1 U5728 ( .A1(n3167), .A2(DATAI_27_), .ZN(n6474) );
  NOR2_X2 U5729 ( .A1(n4795), .A2(n4675), .ZN(n6473) );
  INV_X1 U5730 ( .A(n6473), .ZN(n4838) );
  AND2_X1 U5731 ( .A1(n3167), .A2(DATAI_19_), .ZN(n6380) );
  INV_X1 U5732 ( .A(n6380), .ZN(n6477) );
  INV_X1 U5733 ( .A(n6409), .ZN(n6253) );
  NAND2_X1 U5734 ( .A1(n6222), .A2(n6076), .ZN(n6331) );
  OAI22_X1 U5735 ( .A1(n4838), .A2(n6319), .B1(n6477), .B2(n6331), .ZN(n4676)
         );
  AOI21_X1 U5736 ( .B1(n6474), .B2(n6312), .A(n4676), .ZN(n4677) );
  OAI211_X1 U5737 ( .C1(n4815), .C2(n4934), .A(n4678), .B(n4677), .ZN(U3111)
         );
  NOR2_X2 U5738 ( .A1(n4679), .A2(n6227), .ZN(n6466) );
  INV_X1 U5739 ( .A(n6466), .ZN(n4942) );
  NAND2_X1 U5740 ( .A1(n6324), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n4683)
         );
  AND2_X1 U5741 ( .A1(n3167), .A2(DATAI_26_), .ZN(n6468) );
  NOR2_X2 U5742 ( .A1(n4795), .A2(n4680), .ZN(n6467) );
  INV_X1 U5743 ( .A(n6467), .ZN(n4850) );
  AND2_X1 U5744 ( .A1(n3167), .A2(DATAI_18_), .ZN(n6376) );
  INV_X1 U5745 ( .A(n6376), .ZN(n6471) );
  OAI22_X1 U5746 ( .A1(n4850), .A2(n6319), .B1(n6471), .B2(n6331), .ZN(n4681)
         );
  AOI21_X1 U5747 ( .B1(n6468), .B2(n6312), .A(n4681), .ZN(n4682) );
  OAI211_X1 U5748 ( .C1(n4815), .C2(n4942), .A(n4683), .B(n4682), .ZN(U3110)
         );
  INV_X1 U5749 ( .A(DATAI_7_), .ZN(n6961) );
  NOR2_X2 U5750 ( .A1(n6961), .A2(n6227), .ZN(n6499) );
  INV_X1 U5751 ( .A(n6499), .ZN(n4946) );
  NAND2_X1 U5752 ( .A1(n6324), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n4686)
         );
  AND2_X1 U5753 ( .A1(n3167), .A2(DATAI_31_), .ZN(n6435) );
  NOR2_X2 U5754 ( .A1(n4795), .A2(n5381), .ZN(n6501) );
  INV_X1 U5755 ( .A(n6501), .ZN(n4830) );
  AND2_X1 U5756 ( .A1(n3167), .A2(DATAI_23_), .ZN(n6503) );
  INV_X1 U5757 ( .A(n6503), .ZN(n6439) );
  OAI22_X1 U5758 ( .A1(n4830), .A2(n6319), .B1(n6439), .B2(n6331), .ZN(n4684)
         );
  AOI21_X1 U5759 ( .B1(n6435), .B2(n6312), .A(n4684), .ZN(n4685) );
  OAI211_X1 U5760 ( .C1(n4815), .C2(n4946), .A(n4686), .B(n4685), .ZN(U3115)
         );
  INV_X1 U5761 ( .A(n4689), .ZN(n4687) );
  NOR2_X1 U5762 ( .A1(n6075), .A2(n4666), .ZN(n6368) );
  NAND2_X1 U5763 ( .A1(n6368), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6408) );
  NAND2_X1 U5764 ( .A1(n6408), .A2(n4688), .ZN(n4823) );
  INV_X1 U5765 ( .A(n4823), .ZN(n4691) );
  OR2_X1 U5766 ( .A1(n6068), .A2(n4689), .ZN(n4891) );
  INV_X1 U5767 ( .A(n4891), .ZN(n4726) );
  INV_X1 U5768 ( .A(n5542), .ZN(n4690) );
  NAND2_X1 U5769 ( .A1(n4726), .A2(n4690), .ZN(n4720) );
  AOI21_X1 U5770 ( .B1(n4691), .B2(n4720), .A(n6643), .ZN(n4694) );
  INV_X1 U5771 ( .A(n6070), .ZN(n4692) );
  NAND2_X1 U5772 ( .A1(n6405), .A2(n6852), .ZN(n6289) );
  INV_X1 U5773 ( .A(n6257), .ZN(n6399) );
  OAI22_X1 U5774 ( .A1(n4692), .A2(n6289), .B1(n6399), .B2(n3184), .ZN(n4693)
         );
  OAI21_X1 U5775 ( .B1(n4694), .B2(n4693), .A(n6066), .ZN(n4695) );
  OAI21_X1 U5776 ( .B1(n6066), .B2(n6403), .A(n4695), .ZN(U3462) );
  AOI211_X1 U5777 ( .C1(n6065), .C2(n6064), .A(INSTADDRPOINTER_REG_1__SCAN_IN), 
        .B(n5181), .ZN(n4704) );
  NAND2_X1 U5778 ( .A1(n5100), .A2(n6065), .ZN(n6056) );
  AOI21_X1 U5779 ( .B1(n6063), .B2(n6056), .A(n4696), .ZN(n4703) );
  OAI21_X1 U5780 ( .B1(n4699), .B2(n4698), .A(n4697), .ZN(n5999) );
  AOI22_X1 U5781 ( .A1(n6041), .A2(n4700), .B1(n6054), .B2(REIP_REG_1__SCAN_IN), .ZN(n4701) );
  OAI21_X1 U5782 ( .B1(n5999), .B2(n6033), .A(n4701), .ZN(n4702) );
  OR3_X1 U5783 ( .A1(n4704), .A2(n4703), .A3(n4702), .ZN(U3017) );
  XNOR2_X1 U5784 ( .A(n4706), .B(n4705), .ZN(n4719) );
  INV_X1 U5785 ( .A(n4707), .ZN(n5869) );
  NAND2_X1 U5786 ( .A1(n5983), .A2(n5860), .ZN(n4708) );
  NAND2_X1 U5787 ( .A1(n6054), .A2(REIP_REG_3__SCAN_IN), .ZN(n4712) );
  OAI211_X1 U5788 ( .C1(n5989), .C2(n5863), .A(n4708), .B(n4712), .ZN(n4709)
         );
  AOI21_X1 U5789 ( .B1(n5869), .B2(n3167), .A(n4709), .ZN(n4710) );
  OAI21_X1 U5790 ( .B1(n4719), .B2(n5972), .A(n4710), .ZN(U2983) );
  INV_X1 U5791 ( .A(n4711), .ZN(n4714) );
  AOI21_X1 U5792 ( .B1(n4714), .B2(n6049), .A(n6048), .ZN(n4876) );
  NOR2_X1 U5793 ( .A1(n6047), .A2(n4876), .ZN(n6037) );
  OAI21_X1 U5794 ( .B1(n6058), .B2(n4713), .A(n4712), .ZN(n4716) );
  OAI21_X1 U5795 ( .B1(n4871), .B2(n4714), .A(n4875), .ZN(n6042) );
  AOI21_X1 U5796 ( .B1(n6048), .B2(n6047), .A(n6042), .ZN(n6028) );
  NOR2_X1 U5797 ( .A1(n6028), .A2(n4717), .ZN(n4715) );
  AOI211_X1 U5798 ( .C1(n6037), .C2(n4717), .A(n4716), .B(n4715), .ZN(n4718)
         );
  OAI21_X1 U5799 ( .B1(n4719), .B2(n6033), .A(n4718), .ZN(U3015) );
  INV_X1 U5800 ( .A(n6215), .ZN(n4798) );
  NAND2_X1 U5801 ( .A1(n6405), .A2(n4720), .ZN(n4724) );
  INV_X1 U5802 ( .A(n4533), .ZN(n5024) );
  NAND2_X1 U5803 ( .A1(n5024), .A2(n5009), .ZN(n6441) );
  OR2_X1 U5804 ( .A1(n6257), .A2(n6441), .ZN(n6188) );
  INV_X1 U5805 ( .A(n6188), .ZN(n4721) );
  INV_X1 U5806 ( .A(n6624), .ZN(n6256) );
  AOI21_X1 U5807 ( .B1(n4721), .B2(n6256), .A(n6215), .ZN(n4725) );
  INV_X1 U5808 ( .A(n4725), .ZN(n4723) );
  AOI21_X1 U5809 ( .B1(n6186), .B2(n6643), .A(n6451), .ZN(n4722) );
  OAI21_X1 U5810 ( .B1(n4724), .B2(n4723), .A(n4722), .ZN(n6217) );
  OAI22_X1 U5811 ( .A1(n4725), .A2(n4724), .B1(n6443), .B2(n6186), .ZN(n6216)
         );
  AOI22_X1 U5812 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n6217), .B1(n6499), 
        .B2(n6216), .ZN(n4728) );
  NAND2_X1 U5813 ( .A1(n4726), .A2(n6398), .ZN(n6220) );
  AOI22_X1 U5814 ( .A1(n6187), .A2(n6435), .B1(n6249), .B2(n6503), .ZN(n4727)
         );
  OAI211_X1 U5815 ( .C1(n4830), .C2(n4798), .A(n4728), .B(n4727), .ZN(U3083)
         );
  AOI22_X1 U5816 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n6217), .B1(n6472), 
        .B2(n6216), .ZN(n4730) );
  AOI22_X1 U5817 ( .A1(n6187), .A2(n6474), .B1(n6249), .B2(n6380), .ZN(n4729)
         );
  OAI211_X1 U5818 ( .C1(n4838), .C2(n4798), .A(n4730), .B(n4729), .ZN(U3079)
         );
  NOR2_X2 U5819 ( .A1(n4795), .A2(n3162), .ZN(n6461) );
  INV_X1 U5820 ( .A(n6461), .ZN(n4842) );
  NOR2_X2 U5821 ( .A1(n6839), .A2(n6227), .ZN(n6460) );
  AOI22_X1 U5822 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n6217), .B1(n6460), 
        .B2(n6216), .ZN(n4733) );
  AND2_X1 U5823 ( .A1(n3167), .A2(DATAI_25_), .ZN(n6462) );
  AND2_X1 U5824 ( .A1(n3167), .A2(DATAI_17_), .ZN(n6372) );
  AOI22_X1 U5825 ( .A1(n6187), .A2(n6462), .B1(n6249), .B2(n6372), .ZN(n4732)
         );
  OAI211_X1 U5826 ( .C1(n4842), .C2(n4798), .A(n4733), .B(n4732), .ZN(U3077)
         );
  INV_X1 U5827 ( .A(n4734), .ZN(n4737) );
  INV_X1 U5828 ( .A(n4625), .ZN(n4736) );
  AOI21_X1 U5829 ( .B1(n4737), .B2(n4736), .A(n4776), .ZN(n5856) );
  INV_X1 U5830 ( .A(n5856), .ZN(n4764) );
  AND2_X1 U5831 ( .A1(n4740), .A2(n4739), .ZN(n4741) );
  NOR2_X1 U5832 ( .A1(n4738), .A2(n4741), .ZN(n6030) );
  AOI22_X1 U5833 ( .A1(n5888), .A2(n6030), .B1(EBX_REG_4__SCAN_IN), .B2(n5379), 
        .ZN(n4742) );
  OAI21_X1 U5834 ( .B1(n4764), .B2(n3166), .A(n4742), .ZN(U2855) );
  NAND2_X1 U5835 ( .A1(n4744), .A2(n4743), .ZN(n4745) );
  XNOR2_X1 U5836 ( .A(n4746), .B(n4745), .ZN(n6034) );
  NOR2_X1 U5837 ( .A1(n6015), .A2(n6581), .ZN(n6029) );
  AOI21_X1 U5838 ( .B1(n6012), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n6029), 
        .ZN(n4747) );
  OAI21_X1 U5839 ( .B1(n5859), .B2(n6005), .A(n4747), .ZN(n4748) );
  AOI21_X1 U5840 ( .B1(n5856), .B2(n3167), .A(n4748), .ZN(n4749) );
  OAI21_X1 U5841 ( .B1(n5972), .B2(n6034), .A(n4749), .ZN(U2982) );
  AND2_X1 U5842 ( .A1(n4751), .A2(n4750), .ZN(n4753) );
  XNOR2_X1 U5843 ( .A(n4753), .B(n4752), .ZN(n5981) );
  INV_X1 U5844 ( .A(n6049), .ZN(n4754) );
  NOR2_X1 U5845 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n4754), .ZN(n4762)
         );
  INV_X1 U5846 ( .A(n4755), .ZN(n4786) );
  OAI21_X1 U5847 ( .B1(n4738), .B2(n4756), .A(n4786), .ZN(n5837) );
  NAND2_X1 U5848 ( .A1(n6054), .A2(REIP_REG_5__SCAN_IN), .ZN(n5987) );
  OAI21_X1 U5849 ( .B1(n5837), .B2(n6058), .A(n5987), .ZN(n4760) );
  NAND2_X1 U5850 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n4757), .ZN(n4788)
         );
  AOI21_X1 U5851 ( .B1(n4788), .B2(n5664), .A(n6042), .ZN(n4790) );
  AOI21_X1 U5852 ( .B1(n6048), .B2(n4757), .A(INSTADDRPOINTER_REG_5__SCAN_IN), 
        .ZN(n4758) );
  NOR2_X1 U5853 ( .A1(n4790), .A2(n4758), .ZN(n4759) );
  AOI211_X1 U5854 ( .C1(n4762), .C2(n4761), .A(n4760), .B(n4759), .ZN(n4763)
         );
  OAI21_X1 U5855 ( .B1(n6033), .B2(n5981), .A(n4763), .ZN(U3013) );
  INV_X1 U5856 ( .A(EAX_REG_4__SCAN_IN), .ZN(n5957) );
  INV_X1 U5857 ( .A(DATAI_4_), .ZN(n6978) );
  OAI222_X1 U5858 ( .A1(n5413), .A2(n4764), .B1(n5905), .B2(n5957), .C1(n5904), 
        .C2(n6978), .ZN(U2887) );
  NOR2_X2 U5859 ( .A1(n4795), .A2(n4765), .ZN(n6479) );
  INV_X1 U5860 ( .A(n6479), .ZN(n4858) );
  NOR2_X2 U5861 ( .A1(n6978), .A2(n6227), .ZN(n6478) );
  AOI22_X1 U5862 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n6217), .B1(n6478), 
        .B2(n6216), .ZN(n4767) );
  AND2_X1 U5863 ( .A1(n3167), .A2(DATAI_28_), .ZN(n6481) );
  AND2_X1 U5864 ( .A1(n3167), .A2(DATAI_20_), .ZN(n6384) );
  AOI22_X1 U5865 ( .A1(n6187), .A2(n6481), .B1(n6249), .B2(n6384), .ZN(n4766)
         );
  OAI211_X1 U5866 ( .C1(n4858), .C2(n4798), .A(n4767), .B(n4766), .ZN(U3080)
         );
  INV_X1 U5868 ( .A(DATAI_5_), .ZN(n4778) );
  NOR2_X2 U5869 ( .A1(n4778), .A2(n6227), .ZN(n6486) );
  AOI22_X1 U5870 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n6217), .B1(n6486), 
        .B2(n6216), .ZN(n4769) );
  AND2_X1 U5871 ( .A1(n3167), .A2(DATAI_29_), .ZN(n6424) );
  AND2_X1 U5872 ( .A1(n3167), .A2(DATAI_21_), .ZN(n6488) );
  AOI22_X1 U5873 ( .A1(n6187), .A2(n6424), .B1(n6249), .B2(n6488), .ZN(n4768)
         );
  OAI211_X1 U5874 ( .C1(n7052), .C2(n4798), .A(n4769), .B(n4768), .ZN(U3081)
         );
  INV_X1 U5875 ( .A(DATAI_0_), .ZN(n7023) );
  NOR2_X2 U5876 ( .A1(n7023), .A2(n6227), .ZN(n6445) );
  INV_X1 U5877 ( .A(n6445), .ZN(n4900) );
  NAND2_X1 U5878 ( .A1(n6324), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n4773)
         );
  AND2_X1 U5879 ( .A1(n3167), .A2(DATAI_24_), .ZN(n6412) );
  NOR2_X2 U5880 ( .A1(n4795), .A2(n4770), .ZN(n6446) );
  INV_X1 U5881 ( .A(n6446), .ZN(n4846) );
  AND2_X1 U5882 ( .A1(n3167), .A2(DATAI_16_), .ZN(n6456) );
  INV_X1 U5883 ( .A(n6456), .ZN(n6415) );
  OAI22_X1 U5884 ( .A1(n4846), .A2(n6319), .B1(n6415), .B2(n6331), .ZN(n4771)
         );
  AOI21_X1 U5885 ( .B1(n6412), .B2(n6312), .A(n4771), .ZN(n4772) );
  OAI211_X1 U5886 ( .C1(n4815), .C2(n4900), .A(n4773), .B(n4772), .ZN(U3108)
         );
  OR2_X1 U5887 ( .A1(n4776), .A2(n4775), .ZN(n4777) );
  AND2_X1 U5888 ( .A1(n4774), .A2(n4777), .ZN(n5985) );
  INV_X1 U5889 ( .A(n5985), .ZN(n4780) );
  INV_X1 U5890 ( .A(EAX_REG_5__SCAN_IN), .ZN(n5955) );
  OAI222_X1 U5891 ( .A1(n4780), .A2(n5413), .B1(n5904), .B2(n4778), .C1(n5905), 
        .C2(n5955), .ZN(U2886) );
  INV_X1 U5892 ( .A(EBX_REG_5__SCAN_IN), .ZN(n4779) );
  OAI222_X1 U5893 ( .A1(n4780), .A2(n3166), .B1(n4779), .B2(n5892), .C1(n5378), 
        .C2(n5837), .ZN(U2854) );
  CLKBUF_X1 U5894 ( .A(n4781), .Z(n4782) );
  XNOR2_X1 U5895 ( .A(n4783), .B(n4782), .ZN(n4808) );
  INV_X1 U5896 ( .A(n4784), .ZN(n4785) );
  AOI21_X1 U5897 ( .B1(n4787), .B2(n4786), .A(n4785), .ZN(n5834) );
  NOR2_X1 U5898 ( .A1(n6015), .A2(n6583), .ZN(n4803) );
  OAI33_X1 U5900 ( .A1(1'b0), .A2(n4790), .A3(n4789), .B1(
        INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n4876), .B3(n4788), .ZN(n4792) );
  AOI211_X1 U5901 ( .C1(n6041), .C2(n5834), .A(n4803), .B(n4792), .ZN(n4793)
         );
  OAI21_X1 U5902 ( .B1(n6033), .B2(n4808), .A(n4793), .ZN(U3012) );
  NOR2_X2 U5903 ( .A1(n4795), .A2(n4794), .ZN(n6493) );
  INV_X1 U5904 ( .A(n6493), .ZN(n4863) );
  INV_X1 U5905 ( .A(DATAI_6_), .ZN(n7008) );
  NOR2_X2 U5906 ( .A1(n7008), .A2(n6227), .ZN(n6492) );
  AOI22_X1 U5907 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n6217), .B1(n6492), 
        .B2(n6216), .ZN(n4797) );
  AND2_X1 U5908 ( .A1(n3167), .A2(DATAI_30_), .ZN(n6428) );
  AND2_X1 U5909 ( .A1(n3167), .A2(DATAI_22_), .ZN(n6494) );
  AOI22_X1 U5910 ( .A1(n6187), .A2(n6428), .B1(n6249), .B2(n6494), .ZN(n4796)
         );
  OAI211_X1 U5911 ( .C1(n4863), .C2(n4798), .A(n4797), .B(n4796), .ZN(U3082)
         );
  INV_X1 U5912 ( .A(n4817), .ZN(n4800) );
  AOI21_X1 U5913 ( .B1(n4801), .B2(n4774), .A(n4800), .ZN(n4806) );
  INV_X1 U5914 ( .A(n4806), .ZN(n5831) );
  AOI22_X1 U5915 ( .A1(n5834), .A2(n5888), .B1(EBX_REG_6__SCAN_IN), .B2(n5379), 
        .ZN(n4802) );
  OAI21_X1 U5916 ( .B1(n5831), .B2(n3166), .A(n4802), .ZN(U2853) );
  AOI21_X1 U5917 ( .B1(n6012), .B2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n4803), 
        .ZN(n4804) );
  OAI21_X1 U5918 ( .B1(n5836), .B2(n6005), .A(n4804), .ZN(n4805) );
  AOI21_X1 U5919 ( .B1(n4806), .B2(n3167), .A(n4805), .ZN(n4807) );
  OAI21_X1 U5920 ( .B1(n5972), .B2(n4808), .A(n4807), .ZN(U2980) );
  OAI222_X1 U5921 ( .A1(n5831), .A2(n5413), .B1(n5904), .B2(n7008), .C1(n5905), 
        .C2(n3818), .ZN(U2885) );
  INV_X1 U5922 ( .A(n6478), .ZN(n4951) );
  NAND2_X1 U5923 ( .A1(n6324), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n4811)
         );
  INV_X1 U5924 ( .A(n6384), .ZN(n6485) );
  OAI22_X1 U5925 ( .A1(n4858), .A2(n6319), .B1(n6485), .B2(n6331), .ZN(n4809)
         );
  AOI21_X1 U5926 ( .B1(n6481), .B2(n6312), .A(n4809), .ZN(n4810) );
  OAI211_X1 U5927 ( .C1(n4815), .C2(n4951), .A(n4811), .B(n4810), .ZN(U3112)
         );
  INV_X1 U5928 ( .A(n6486), .ZN(n4938) );
  NAND2_X1 U5929 ( .A1(n6324), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n4814)
         );
  INV_X1 U5930 ( .A(n6488), .ZN(n6427) );
  OAI22_X1 U5931 ( .A1(n7052), .A2(n6319), .B1(n6427), .B2(n6331), .ZN(n4812)
         );
  AOI21_X1 U5932 ( .B1(n6424), .B2(n6312), .A(n4812), .ZN(n4813) );
  OAI211_X1 U5933 ( .C1(n4815), .C2(n4938), .A(n4814), .B(n4813), .ZN(U3113)
         );
  AND2_X1 U5934 ( .A1(n4817), .A2(n4816), .ZN(n4818) );
  NOR2_X1 U5935 ( .A1(n4817), .A2(n4816), .ZN(n5018) );
  OR2_X1 U5936 ( .A1(n4818), .A2(n5018), .ZN(n5975) );
  NAND2_X1 U5937 ( .A1(n4784), .A2(n4819), .ZN(n4820) );
  NAND2_X1 U5938 ( .A1(n4881), .A2(n4820), .ZN(n5811) );
  OAI22_X1 U5939 ( .A1(n5811), .A2(n5378), .B1(n5813), .B2(n5892), .ZN(n4821)
         );
  INV_X1 U5940 ( .A(n4821), .ZN(n4822) );
  OAI21_X1 U5941 ( .B1(n5975), .B2(n3166), .A(n4822), .ZN(U2852) );
  NOR3_X1 U5942 ( .A1(n4823), .A2(n3165), .A3(n5542), .ZN(n4824) );
  NOR2_X1 U5943 ( .A1(n4824), .A2(n6643), .ZN(n4832) );
  OR2_X1 U5944 ( .A1(n6257), .A2(n4825), .ZN(n6133) );
  NAND2_X1 U5945 ( .A1(n4826), .A2(n6403), .ZN(n4862) );
  OAI21_X1 U5946 ( .B1(n6133), .B2(n6624), .A(n4862), .ZN(n4835) );
  NAND3_X1 U5947 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n6403), .A3(n6521), .ZN(n6130) );
  INV_X1 U5948 ( .A(n6130), .ZN(n4827) );
  AOI22_X1 U5949 ( .A1(n4832), .A2(n4835), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4827), .ZN(n4868) );
  NAND2_X1 U5950 ( .A1(n6398), .A2(n6068), .ZN(n4828) );
  NAND2_X1 U5951 ( .A1(n6076), .A2(n6068), .ZN(n4829) );
  OAI22_X1 U5952 ( .A1(n4830), .A2(n4862), .B1(n4957), .B2(n6439), .ZN(n4831)
         );
  AOI21_X1 U5953 ( .B1(n6435), .B2(n3182), .A(n4831), .ZN(n4837) );
  INV_X1 U5954 ( .A(n4832), .ZN(n4834) );
  AOI21_X1 U5955 ( .B1(n6130), .B2(n6643), .A(n6451), .ZN(n4833) );
  OAI21_X1 U5956 ( .B1(n4835), .B2(n4834), .A(n4833), .ZN(n4865) );
  NAND2_X1 U5957 ( .A1(n4865), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4836) );
  OAI211_X1 U5958 ( .C1(n4868), .C2(n4946), .A(n4837), .B(n4836), .ZN(U3051)
         );
  OAI22_X1 U5959 ( .A1(n4838), .A2(n4862), .B1(n4957), .B2(n6477), .ZN(n4839)
         );
  AOI21_X1 U5960 ( .B1(n6474), .B2(n3182), .A(n4839), .ZN(n4841) );
  NAND2_X1 U5961 ( .A1(n4865), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4840) );
  OAI211_X1 U5962 ( .C1(n4868), .C2(n4934), .A(n4841), .B(n4840), .ZN(U3047)
         );
  INV_X1 U5963 ( .A(n6460), .ZN(n4930) );
  INV_X1 U5964 ( .A(n6372), .ZN(n6465) );
  OAI22_X1 U5965 ( .A1(n4842), .A2(n4862), .B1(n4957), .B2(n6465), .ZN(n4843)
         );
  AOI21_X1 U5966 ( .B1(n6462), .B2(n3182), .A(n4843), .ZN(n4845) );
  NAND2_X1 U5967 ( .A1(n4865), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4844) );
  OAI211_X1 U5968 ( .C1(n4868), .C2(n4930), .A(n4845), .B(n4844), .ZN(U3045)
         );
  OAI22_X1 U5969 ( .A1(n4846), .A2(n4862), .B1(n4957), .B2(n6415), .ZN(n4847)
         );
  AOI21_X1 U5970 ( .B1(n6412), .B2(n3182), .A(n4847), .ZN(n4849) );
  NAND2_X1 U5971 ( .A1(n4865), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4848) );
  OAI211_X1 U5972 ( .C1(n4868), .C2(n4900), .A(n4849), .B(n4848), .ZN(U3044)
         );
  OAI22_X1 U5973 ( .A1(n4850), .A2(n4862), .B1(n4957), .B2(n6471), .ZN(n4851)
         );
  AOI21_X1 U5974 ( .B1(n6468), .B2(n3182), .A(n4851), .ZN(n4853) );
  NAND2_X1 U5975 ( .A1(n4865), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4852) );
  OAI211_X1 U5976 ( .C1(n4868), .C2(n4942), .A(n4853), .B(n4852), .ZN(U3046)
         );
  OAI22_X1 U5977 ( .A1(n7052), .A2(n4862), .B1(n4957), .B2(n6427), .ZN(n4855)
         );
  AOI21_X1 U5978 ( .B1(n6424), .B2(n3182), .A(n4855), .ZN(n4857) );
  NAND2_X1 U5979 ( .A1(n4865), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4856) );
  OAI211_X1 U5980 ( .C1(n4868), .C2(n4938), .A(n4857), .B(n4856), .ZN(U3049)
         );
  OAI22_X1 U5981 ( .A1(n4858), .A2(n4862), .B1(n4957), .B2(n6485), .ZN(n4859)
         );
  AOI21_X1 U5982 ( .B1(n6481), .B2(n3182), .A(n4859), .ZN(n4861) );
  NAND2_X1 U5983 ( .A1(n4865), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4860) );
  OAI211_X1 U5984 ( .C1(n4868), .C2(n4951), .A(n4861), .B(n4860), .ZN(U3048)
         );
  INV_X1 U5985 ( .A(n6492), .ZN(n4926) );
  INV_X1 U5986 ( .A(n6494), .ZN(n6431) );
  OAI22_X1 U5987 ( .A1(n4863), .A2(n4862), .B1(n4957), .B2(n6431), .ZN(n4864)
         );
  AOI21_X1 U5988 ( .B1(n6428), .B2(n3182), .A(n4864), .ZN(n4867) );
  NAND2_X1 U5989 ( .A1(n4865), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4866) );
  OAI211_X1 U5990 ( .C1(n4868), .C2(n4926), .A(n4867), .B(n4866), .ZN(U3050)
         );
  INV_X1 U5991 ( .A(EAX_REG_7__SCAN_IN), .ZN(n5951) );
  OAI222_X1 U5992 ( .A1(n5975), .A2(n5413), .B1(n5904), .B2(n6961), .C1(n5905), 
        .C2(n5951), .ZN(U2884) );
  XNOR2_X1 U5993 ( .A(n4869), .B(n4870), .ZN(n5047) );
  INV_X1 U5994 ( .A(n4871), .ZN(n4873) );
  AOI22_X1 U5995 ( .A1(n6048), .A2(n4877), .B1(n4873), .B2(n4872), .ZN(n4874)
         );
  NAND2_X1 U5996 ( .A1(n4875), .A2(n4874), .ZN(n5062) );
  NOR2_X1 U5997 ( .A1(n4877), .A2(n4876), .ZN(n4913) );
  AOI21_X1 U5998 ( .B1(n4879), .B2(n4878), .A(n4914), .ZN(n4880) );
  AOI22_X1 U5999 ( .A1(INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n5062), .B1(n4913), 
        .B2(n4880), .ZN(n4884) );
  AOI21_X1 U6000 ( .B1(n4882), .B2(n4881), .A(n4911), .ZN(n5799) );
  NOR2_X1 U6001 ( .A1(n6015), .A2(n6586), .ZN(n5043) );
  AOI21_X1 U6002 ( .B1(n5799), .B2(n6041), .A(n5043), .ZN(n4883) );
  OAI211_X1 U6003 ( .C1(n5047), .C2(n6033), .A(n4884), .B(n4883), .ZN(U3010)
         );
  INV_X1 U6004 ( .A(n4913), .ZN(n4890) );
  XOR2_X1 U6005 ( .A(n4885), .B(n4886), .Z(n5977) );
  NAND2_X1 U6006 ( .A1(n5977), .A2(n6060), .ZN(n4889) );
  NAND2_X1 U6007 ( .A1(n6054), .A2(REIP_REG_7__SCAN_IN), .ZN(n5978) );
  OAI21_X1 U6008 ( .B1(n5811), .B2(n6058), .A(n5978), .ZN(n4887) );
  AOI21_X1 U6009 ( .B1(n5062), .B2(INSTADDRPOINTER_REG_7__SCAN_IN), .A(n4887), 
        .ZN(n4888) );
  OAI211_X1 U6010 ( .C1(INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n4890), .A(n4889), 
        .B(n4888), .ZN(U3011) );
  NOR2_X1 U6011 ( .A1(n4891), .A2(n4666), .ZN(n4896) );
  INV_X1 U6012 ( .A(n4896), .ZN(n6157) );
  OAI21_X1 U6013 ( .B1(n6157), .B2(n6852), .A(n6405), .ZN(n6164) );
  INV_X1 U6014 ( .A(n6289), .ZN(n6449) );
  NOR2_X1 U6015 ( .A1(n4533), .A2(n5009), .ZN(n6360) );
  INV_X1 U6016 ( .A(n6360), .ZN(n6333) );
  OAI22_X1 U6017 ( .A1(n4957), .A2(n6449), .B1(n4892), .B2(n6333), .ZN(n4895)
         );
  NAND2_X1 U6018 ( .A1(n6517), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6362) );
  OR2_X1 U6019 ( .A1(n6362), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6162)
         );
  NOR2_X1 U6020 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6162), .ZN(n4954)
         );
  INV_X1 U6021 ( .A(n4954), .ZN(n4893) );
  AND2_X1 U6022 ( .A1(n4897), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6402) );
  INV_X1 U6023 ( .A(n6294), .ZN(n6401) );
  AND2_X1 U6024 ( .A1(n6223), .A2(n6401), .ZN(n6072) );
  OAI21_X1 U6025 ( .B1(n6072), .B2(n6443), .A(n6135), .ZN(n6078) );
  AOI211_X1 U6026 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4893), .A(n6402), .B(
        n6078), .ZN(n4894) );
  OAI21_X1 U6027 ( .B1(n6164), .B2(n4895), .A(n4894), .ZN(n4950) );
  INV_X1 U6028 ( .A(n4950), .ZN(n4905) );
  INV_X1 U6029 ( .A(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4904) );
  INV_X1 U6030 ( .A(n6412), .ZN(n6459) );
  NOR2_X1 U6031 ( .A1(n4957), .A2(n6459), .ZN(n4902) );
  NAND2_X1 U6032 ( .A1(n4896), .A2(n6409), .ZN(n6184) );
  AND2_X1 U6033 ( .A1(n6360), .A2(n6405), .ZN(n6328) );
  NAND2_X1 U6034 ( .A1(n6328), .A2(n6399), .ZN(n4899) );
  NOR2_X1 U6035 ( .A1(n4897), .A2(n6443), .ZN(n6226) );
  NAND2_X1 U6036 ( .A1(n6072), .A2(n6226), .ZN(n4898) );
  AND2_X1 U6037 ( .A1(n4899), .A2(n4898), .ZN(n4952) );
  OAI22_X1 U6038 ( .A1(n6184), .A2(n6415), .B1(n4952), .B2(n4900), .ZN(n4901)
         );
  AOI211_X1 U6039 ( .C1(n6446), .C2(n4954), .A(n4902), .B(n4901), .ZN(n4903)
         );
  OAI21_X1 U6040 ( .B1(n4905), .B2(n4904), .A(n4903), .ZN(U3052) );
  XNOR2_X1 U6041 ( .A(n5092), .B(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n4908)
         );
  XNOR2_X1 U6042 ( .A(n4907), .B(n4908), .ZN(n5017) );
  INV_X1 U6043 ( .A(n5062), .ZN(n4909) );
  OAI21_X1 U6044 ( .B1(n5181), .B2(n4914), .A(n4909), .ZN(n6021) );
  NOR2_X1 U6045 ( .A1(n4911), .A2(n4910), .ZN(n4912) );
  OR2_X1 U6046 ( .A1(n4923), .A2(n4912), .ZN(n5785) );
  NOR2_X1 U6047 ( .A1(n5785), .A2(n6058), .ZN(n4916) );
  NAND2_X1 U6048 ( .A1(n4914), .A2(n4913), .ZN(n6026) );
  NAND2_X1 U6049 ( .A1(n6054), .A2(REIP_REG_9__SCAN_IN), .ZN(n5013) );
  OAI21_X1 U6050 ( .B1(INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n6026), .A(n5013), 
        .ZN(n4915) );
  AOI211_X1 U6051 ( .C1(n6021), .C2(INSTADDRPOINTER_REG_9__SCAN_IN), .A(n4916), 
        .B(n4915), .ZN(n4917) );
  OAI21_X1 U6052 ( .B1(n5017), .B2(n6033), .A(n4917), .ZN(U3009) );
  NAND2_X1 U6053 ( .A1(n5018), .A2(n5019), .ZN(n4967) );
  NOR2_X1 U6054 ( .A1(n4967), .A2(n4968), .ZN(n4966) );
  INV_X1 U6055 ( .A(n4918), .ZN(n4920) );
  NAND2_X1 U6056 ( .A1(n5018), .A2(n4919), .ZN(n4973) );
  OAI21_X1 U6057 ( .B1(n4966), .B2(n4920), .A(n4973), .ZN(n5090) );
  INV_X1 U6058 ( .A(n5904), .ZN(n5142) );
  AOI22_X1 U6059 ( .A1(n5142), .A2(DATAI_10_), .B1(EAX_REG_10__SCAN_IN), .B2(
        n5900), .ZN(n4921) );
  OAI21_X1 U6060 ( .B1(n5090), .B2(n5413), .A(n4921), .ZN(U2881) );
  OAI21_X1 U6061 ( .B1(n4923), .B2(n4922), .A(n4976), .ZN(n4924) );
  INV_X1 U6062 ( .A(n4924), .ZN(n6020) );
  AOI22_X1 U6063 ( .A1(n6020), .A2(n5888), .B1(EBX_REG_10__SCAN_IN), .B2(n5379), .ZN(n4925) );
  OAI21_X1 U6064 ( .B1(n5090), .B2(n3166), .A(n4925), .ZN(U2849) );
  INV_X1 U6065 ( .A(n6428), .ZN(n6497) );
  NAND2_X1 U6066 ( .A1(n4950), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4929) );
  OAI22_X1 U6067 ( .A1(n6184), .A2(n6431), .B1(n4952), .B2(n4926), .ZN(n4927)
         );
  AOI21_X1 U6068 ( .B1(n4954), .B2(n6493), .A(n4927), .ZN(n4928) );
  OAI211_X1 U6069 ( .C1(n4957), .C2(n6497), .A(n4929), .B(n4928), .ZN(U3058)
         );
  INV_X1 U6070 ( .A(n6462), .ZN(n6375) );
  NAND2_X1 U6071 ( .A1(n4950), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4933) );
  OAI22_X1 U6072 ( .A1(n6184), .A2(n6465), .B1(n4952), .B2(n4930), .ZN(n4931)
         );
  AOI21_X1 U6073 ( .B1(n4954), .B2(n6461), .A(n4931), .ZN(n4932) );
  OAI211_X1 U6074 ( .C1(n4957), .C2(n6375), .A(n4933), .B(n4932), .ZN(U3053)
         );
  INV_X1 U6075 ( .A(n6474), .ZN(n6383) );
  NAND2_X1 U6076 ( .A1(n4950), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4937) );
  OAI22_X1 U6077 ( .A1(n6184), .A2(n6477), .B1(n4952), .B2(n4934), .ZN(n4935)
         );
  AOI21_X1 U6078 ( .B1(n4954), .B2(n6473), .A(n4935), .ZN(n4936) );
  OAI211_X1 U6079 ( .C1(n4957), .C2(n6383), .A(n4937), .B(n4936), .ZN(U3055)
         );
  INV_X1 U6080 ( .A(n6424), .ZN(n6491) );
  NAND2_X1 U6081 ( .A1(n4950), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4941) );
  OAI22_X1 U6082 ( .A1(n6184), .A2(n6427), .B1(n4952), .B2(n4938), .ZN(n4939)
         );
  AOI21_X1 U6083 ( .B1(n4954), .B2(n3161), .A(n4939), .ZN(n4940) );
  OAI211_X1 U6084 ( .C1(n4957), .C2(n6491), .A(n4941), .B(n4940), .ZN(U3057)
         );
  INV_X1 U6085 ( .A(n6468), .ZN(n6379) );
  NAND2_X1 U6086 ( .A1(n4950), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4945) );
  OAI22_X1 U6087 ( .A1(n6184), .A2(n6471), .B1(n4952), .B2(n4942), .ZN(n4943)
         );
  AOI21_X1 U6088 ( .B1(n4954), .B2(n6467), .A(n4943), .ZN(n4944) );
  OAI211_X1 U6089 ( .C1(n4957), .C2(n6379), .A(n4945), .B(n4944), .ZN(U3054)
         );
  INV_X1 U6090 ( .A(n6435), .ZN(n6508) );
  NAND2_X1 U6091 ( .A1(n4950), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4949) );
  OAI22_X1 U6092 ( .A1(n6184), .A2(n6439), .B1(n4952), .B2(n4946), .ZN(n4947)
         );
  AOI21_X1 U6093 ( .B1(n4954), .B2(n6501), .A(n4947), .ZN(n4948) );
  OAI211_X1 U6094 ( .C1(n4957), .C2(n6508), .A(n4949), .B(n4948), .ZN(U3059)
         );
  INV_X1 U6095 ( .A(n6481), .ZN(n6387) );
  NAND2_X1 U6096 ( .A1(n4950), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4956) );
  OAI22_X1 U6097 ( .A1(n6184), .A2(n6485), .B1(n4952), .B2(n4951), .ZN(n4953)
         );
  AOI21_X1 U6098 ( .B1(n4954), .B2(n6479), .A(n4953), .ZN(n4955) );
  OAI211_X1 U6099 ( .C1(n4957), .C2(n6387), .A(n4956), .B(n4955), .ZN(U3056)
         );
  AND2_X1 U6100 ( .A1(n4959), .A2(n4958), .ZN(n4972) );
  XOR2_X1 U6101 ( .A(n4960), .B(n4972), .Z(n5076) );
  INV_X1 U6102 ( .A(n5076), .ZN(n5042) );
  NAND2_X1 U6103 ( .A1(n4978), .A2(n4961), .ZN(n4962) );
  NAND2_X1 U6104 ( .A1(n5049), .A2(n4962), .ZN(n5066) );
  INV_X1 U6105 ( .A(EBX_REG_12__SCAN_IN), .ZN(n4963) );
  OAI22_X1 U6106 ( .A1(n5066), .A2(n5378), .B1(n4963), .B2(n5892), .ZN(n4964)
         );
  INV_X1 U6107 ( .A(n4964), .ZN(n4965) );
  OAI21_X1 U6108 ( .B1(n5042), .B2(n3166), .A(n4965), .ZN(U2847) );
  AOI21_X1 U6109 ( .B1(n4968), .B2(n4967), .A(n4966), .ZN(n5789) );
  OAI22_X1 U6110 ( .A1(n5785), .A2(n5378), .B1(n4969), .B2(n5892), .ZN(n4970)
         );
  AOI21_X1 U6111 ( .B1(n5789), .B2(n5889), .A(n4970), .ZN(n4971) );
  INV_X1 U6112 ( .A(n4971), .ZN(U2850) );
  AOI21_X1 U6113 ( .B1(n4974), .B2(n4973), .A(n4972), .ZN(n5969) );
  INV_X1 U6114 ( .A(n5969), .ZN(n4982) );
  INV_X1 U6115 ( .A(EBX_REG_11__SCAN_IN), .ZN(n4979) );
  NAND2_X1 U6116 ( .A1(n4976), .A2(n4975), .ZN(n4977) );
  NAND2_X1 U6117 ( .A1(n4978), .A2(n4977), .ZN(n5778) );
  OAI222_X1 U6118 ( .A1(n4982), .A2(n3166), .B1(n4979), .B2(n5892), .C1(n5378), 
        .C2(n5778), .ZN(U2848) );
  INV_X1 U6119 ( .A(EAX_REG_11__SCAN_IN), .ZN(n4981) );
  INV_X1 U6120 ( .A(DATAI_11_), .ZN(n4980) );
  OAI222_X1 U6121 ( .A1(n4982), .A2(n5413), .B1(n5905), .B2(n4981), .C1(n5904), 
        .C2(n4980), .ZN(U2880) );
  NOR2_X1 U6122 ( .A1(n5876), .A2(n5125), .ZN(n5777) );
  NOR2_X1 U6123 ( .A1(REIP_REG_12__SCAN_IN), .A2(n5766), .ZN(n5772) );
  INV_X1 U6124 ( .A(n4983), .ZN(n4984) );
  NAND3_X1 U6125 ( .A1(n5907), .A2(n4445), .A3(n4984), .ZN(n4985) );
  AND2_X1 U6126 ( .A1(n4986), .A2(n4985), .ZN(n4987) );
  AOI22_X1 U6127 ( .A1(EBX_REG_12__SCAN_IN), .A2(n5879), .B1(
        PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n5849), .ZN(n4989) );
  NAND2_X1 U6128 ( .A1(n5820), .A2(n4988), .ZN(n5825) );
  OAI211_X1 U6129 ( .C1(n5881), .C2(n5066), .A(n4989), .B(n5825), .ZN(n4990)
         );
  AOI211_X1 U6130 ( .C1(n5777), .C2(REIP_REG_12__SCAN_IN), .A(n5772), .B(n4990), .ZN(n4994) );
  AND2_X1 U6131 ( .A1(n4991), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4992) );
  NAND2_X1 U6132 ( .A1(n5802), .A2(n5071), .ZN(n4993) );
  OAI211_X1 U6133 ( .C1(n5042), .C2(n5830), .A(n4994), .B(n4993), .ZN(U2815)
         );
  OAI221_X1 U6134 ( .B1(n5851), .B2(REIP_REG_9__SCAN_IN), .C1(n5851), .C2(
        n5796), .A(n5820), .ZN(n5000) );
  INV_X1 U6135 ( .A(n5825), .ZN(n5848) );
  AOI21_X1 U6136 ( .B1(n5849), .B2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n5848), 
        .ZN(n4995) );
  OAI21_X1 U6137 ( .B1(n5086), .B2(n5885), .A(n4995), .ZN(n4999) );
  INV_X1 U6138 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6589) );
  AOI22_X1 U6139 ( .A1(n5866), .A2(n6020), .B1(n5776), .B2(n6589), .ZN(n4996)
         );
  OAI21_X1 U6140 ( .B1(n4997), .B2(n5862), .A(n4996), .ZN(n4998) );
  AOI211_X1 U6141 ( .C1(REIP_REG_10__SCAN_IN), .C2(n5000), .A(n4999), .B(n4998), .ZN(n5001) );
  OAI21_X1 U6142 ( .B1(n5090), .B2(n5830), .A(n5001), .ZN(U2817) );
  OAI21_X1 U6143 ( .B1(n5002), .B2(n5008), .A(n5830), .ZN(n5883) );
  INV_X1 U6144 ( .A(n5883), .ZN(n5034) );
  INV_X1 U6145 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6577) );
  INV_X1 U6146 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n5003) );
  NOR2_X1 U6147 ( .A1(n5886), .A2(n5003), .ZN(n5006) );
  AOI22_X1 U6148 ( .A1(EBX_REG_1__SCAN_IN), .A2(n5879), .B1(n5844), .B2(
        REIP_REG_1__SCAN_IN), .ZN(n5004) );
  OAI21_X1 U6149 ( .B1(n5885), .B2(PHYADDRPOINTER_REG_1__SCAN_IN), .A(n5004), 
        .ZN(n5005) );
  AOI211_X1 U6150 ( .C1(n6577), .C2(n5845), .A(n5006), .B(n5005), .ZN(n5011)
         );
  OR2_X1 U6151 ( .A1(n5008), .A2(n5007), .ZN(n5877) );
  INV_X1 U6152 ( .A(n5877), .ZN(n5025) );
  AOI22_X1 U6153 ( .A1(n5866), .A2(n4573), .B1(n5009), .B2(n5025), .ZN(n5010)
         );
  OAI211_X1 U6154 ( .C1(n6000), .C2(n5034), .A(n5011), .B(n5010), .ZN(U2826)
         );
  NAND2_X1 U6155 ( .A1(n6012), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n5012)
         );
  OAI211_X1 U6156 ( .C1(n6005), .C2(n5014), .A(n5013), .B(n5012), .ZN(n5015)
         );
  AOI21_X1 U6157 ( .B1(n5789), .B2(n3167), .A(n5015), .ZN(n5016) );
  OAI21_X1 U6158 ( .B1(n5017), .B2(n5972), .A(n5016), .ZN(U2977) );
  XOR2_X1 U6159 ( .A(n5019), .B(n5018), .Z(n5805) );
  INV_X1 U6160 ( .A(n5805), .ZN(n5021) );
  AOI22_X1 U6161 ( .A1(n5799), .A2(n5888), .B1(EBX_REG_8__SCAN_IN), .B2(n5379), 
        .ZN(n5020) );
  OAI21_X1 U6162 ( .B1(n5021), .B2(n3166), .A(n5020), .ZN(U2851) );
  NOR2_X1 U6163 ( .A1(n5862), .A2(n5891), .ZN(n5023) );
  OAI22_X1 U6164 ( .A1(n5998), .A2(n5885), .B1(n5886), .B2(n3786), .ZN(n5022)
         );
  AOI211_X1 U6165 ( .C1(n5025), .C2(n5024), .A(n5023), .B(n5022), .ZN(n5033)
         );
  OAI21_X1 U6166 ( .B1(n5028), .B2(n5027), .A(n5026), .ZN(n5029) );
  INV_X1 U6167 ( .A(n5029), .ZN(n6040) );
  INV_X1 U6168 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6578) );
  OAI21_X1 U6169 ( .B1(n5851), .B2(n6577), .A(n6578), .ZN(n5031) );
  AOI211_X1 U6170 ( .C1(n5845), .C2(n6577), .A(n5844), .B(n6578), .ZN(n5872)
         );
  INV_X1 U6171 ( .A(n5872), .ZN(n5030) );
  AOI22_X1 U6172 ( .A1(n5866), .A2(n6040), .B1(n5031), .B2(n5030), .ZN(n5032)
         );
  OAI211_X1 U6173 ( .C1(n5035), .C2(n5034), .A(n5033), .B(n5032), .ZN(U2825)
         );
  OAI21_X1 U6174 ( .B1(n5038), .B2(n5037), .A(n5036), .ZN(n5765) );
  AOI22_X1 U6175 ( .A1(n5142), .A2(DATAI_13_), .B1(EAX_REG_13__SCAN_IN), .B2(
        n5900), .ZN(n5039) );
  OAI21_X1 U6176 ( .B1(n5765), .B2(n5413), .A(n5039), .ZN(U2878) );
  INV_X1 U6177 ( .A(n5413), .ZN(n5898) );
  AOI222_X1 U6178 ( .A1(n5805), .A2(n5898), .B1(DATAI_8_), .B2(n5142), .C1(
        EAX_REG_8__SCAN_IN), .C2(n5900), .ZN(n5040) );
  INV_X1 U6179 ( .A(n5040), .ZN(U2883) );
  OAI222_X1 U6180 ( .A1(n5904), .A2(n4502), .B1(n5413), .B2(n5042), .C1(n5041), 
        .C2(n5905), .ZN(U2879) );
  AOI21_X1 U6181 ( .B1(n6012), .B2(PHYADDRPOINTER_REG_8__SCAN_IN), .A(n5043), 
        .ZN(n5044) );
  OAI21_X1 U6182 ( .B1(n5801), .B2(n6005), .A(n5044), .ZN(n5045) );
  AOI21_X1 U6183 ( .B1(n5805), .B2(n3167), .A(n5045), .ZN(n5046) );
  OAI21_X1 U6184 ( .B1(n5972), .B2(n5047), .A(n5046), .ZN(U2978) );
  AOI222_X1 U6185 ( .A1(n5789), .A2(n5898), .B1(EAX_REG_9__SCAN_IN), .B2(n5900), .C1(DATAI_9_), .C2(n5142), .ZN(n5048) );
  INV_X1 U6186 ( .A(n5048), .ZN(U2882) );
  INV_X1 U6187 ( .A(EBX_REG_13__SCAN_IN), .ZN(n5051) );
  AOI21_X1 U6188 ( .B1(n5050), .B2(n5049), .A(n5106), .ZN(n5767) );
  INV_X1 U6189 ( .A(n5767), .ZN(n5710) );
  OAI222_X1 U6190 ( .A1(n5765), .A2(n3166), .B1(n5051), .B2(n5892), .C1(n5378), 
        .C2(n5710), .ZN(U2846) );
  NAND2_X1 U6191 ( .A1(n5113), .A2(n5053), .ZN(n5054) );
  NAND2_X1 U6192 ( .A1(n5054), .A2(n5111), .ZN(n5059) );
  INV_X1 U6193 ( .A(n5055), .ZN(n5056) );
  NOR2_X1 U6194 ( .A1(n5057), .A2(n5056), .ZN(n5058) );
  XNOR2_X1 U6195 ( .A(n5059), .B(n5058), .ZN(n5078) );
  INV_X1 U6196 ( .A(n5099), .ZN(n5096) );
  AND2_X1 U6197 ( .A1(n5664), .A2(n5060), .ZN(n5061) );
  NOR2_X1 U6198 ( .A1(n5062), .A2(n5061), .ZN(n5180) );
  OAI221_X1 U6199 ( .B1(n5096), .B2(n5064), .C1(n5096), .C2(n5063), .A(n5180), 
        .ZN(n5069) );
  INV_X1 U6200 ( .A(n5697), .ZN(n5065) );
  OAI21_X1 U6201 ( .B1(n5065), .B2(n5119), .A(n3639), .ZN(n5068) );
  NAND2_X1 U6202 ( .A1(n6054), .A2(REIP_REG_12__SCAN_IN), .ZN(n5072) );
  OAI21_X1 U6203 ( .B1(n5066), .B2(n6058), .A(n5072), .ZN(n5067) );
  AOI21_X1 U6204 ( .B1(n5069), .B2(n5068), .A(n5067), .ZN(n5070) );
  OAI21_X1 U6205 ( .B1(n5078), .B2(n6033), .A(n5070), .ZN(U3006) );
  NAND2_X1 U6206 ( .A1(n5983), .A2(n5071), .ZN(n5073) );
  OAI211_X1 U6207 ( .C1(n5989), .C2(n5074), .A(n5073), .B(n5072), .ZN(n5075)
         );
  AOI21_X1 U6208 ( .B1(n5076), .B2(n3167), .A(n5075), .ZN(n5077) );
  OAI21_X1 U6209 ( .B1(n5078), .B2(n5972), .A(n5077), .ZN(U2974) );
  OR2_X1 U6210 ( .A1(n4907), .A2(n5079), .ZN(n5081) );
  NAND2_X1 U6211 ( .A1(n5081), .A2(n5080), .ZN(n5085) );
  NOR2_X1 U6212 ( .A1(n5083), .A2(n5082), .ZN(n5084) );
  XNOR2_X1 U6213 ( .A(n5085), .B(n5084), .ZN(n6022) );
  NAND2_X1 U6214 ( .A1(n6022), .A2(n6010), .ZN(n5089) );
  NOR2_X1 U6215 ( .A1(n6015), .A2(n6589), .ZN(n6019) );
  NOR2_X1 U6216 ( .A1(n6005), .A2(n5086), .ZN(n5087) );
  AOI211_X1 U6217 ( .C1(n6012), .C2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n6019), 
        .B(n5087), .ZN(n5088) );
  OAI211_X1 U6218 ( .C1(n6447), .C2(n5090), .A(n5089), .B(n5088), .ZN(U2976)
         );
  XNOR2_X1 U6219 ( .A(n5092), .B(n5102), .ZN(n5093) );
  XNOR2_X1 U6220 ( .A(n5091), .B(n5093), .ZN(n5195) );
  INV_X1 U6221 ( .A(n5094), .ZN(n5708) );
  NAND2_X1 U6222 ( .A1(n5096), .A2(n5095), .ZN(n5707) );
  AOI221_X1 U6223 ( .B1(n5708), .B2(n5098), .C1(n5097), .C2(n5098), .A(n5707), 
        .ZN(n5712) );
  AOI21_X1 U6224 ( .B1(n5100), .B2(n5099), .A(n5712), .ZN(n5101) );
  OAI211_X1 U6225 ( .C1(n5103), .C2(n6064), .A(n5180), .B(n5101), .ZN(n5714)
         );
  OAI222_X1 U6226 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n5103), .B1(
        INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n5697), .C1(n5102), .C2(n5714), 
        .ZN(n5109) );
  OAI21_X1 U6227 ( .B1(n5106), .B2(n5105), .A(n5104), .ZN(n5131) );
  INV_X1 U6228 ( .A(n5131), .ZN(n5123) );
  NAND2_X1 U6229 ( .A1(n6054), .A2(REIP_REG_14__SCAN_IN), .ZN(n5189) );
  INV_X1 U6230 ( .A(n5189), .ZN(n5107) );
  AOI21_X1 U6231 ( .B1(n5123), .B2(n6041), .A(n5107), .ZN(n5108) );
  OAI211_X1 U6232 ( .C1(n5195), .C2(n6033), .A(n5109), .B(n5108), .ZN(U3004)
         );
  NAND2_X1 U6233 ( .A1(n5111), .A2(n5110), .ZN(n5115) );
  AND2_X1 U6234 ( .A1(n5113), .A2(n5112), .ZN(n5114) );
  XOR2_X1 U6235 ( .A(n5115), .B(n5114), .Z(n5973) );
  OR2_X1 U6236 ( .A1(n5973), .A2(n6033), .ZN(n5118) );
  OAI22_X1 U6237 ( .A1(n5778), .A2(n6058), .B1(n6015), .B2(n6590), .ZN(n5116)
         );
  AOI21_X1 U6238 ( .B1(n5697), .B2(n5119), .A(n5116), .ZN(n5117) );
  OAI211_X1 U6239 ( .C1(n5180), .C2(n5119), .A(n5118), .B(n5117), .ZN(U3007)
         );
  OAI21_X1 U6240 ( .B1(n5122), .B2(n5121), .A(n5138), .ZN(n5190) );
  AOI22_X1 U6241 ( .A1(n5123), .A2(n5888), .B1(EBX_REG_14__SCAN_IN), .B2(n5379), .ZN(n5124) );
  OAI21_X1 U6242 ( .B1(n5190), .B2(n3166), .A(n5124), .ZN(U2845) );
  INV_X1 U6243 ( .A(n5144), .ZN(n5126) );
  AOI21_X1 U6244 ( .B1(n5126), .B2(n5125), .A(n5876), .ZN(n5170) );
  NAND2_X1 U6245 ( .A1(REIP_REG_13__SCAN_IN), .A2(REIP_REG_12__SCAN_IN), .ZN(
        n5127) );
  INV_X1 U6246 ( .A(REIP_REG_14__SCAN_IN), .ZN(n6595) );
  OAI21_X1 U6247 ( .B1(n5766), .B2(n5127), .A(n6595), .ZN(n5134) );
  OAI22_X1 U6248 ( .A1(n5129), .A2(n5862), .B1(n5128), .B2(n5886), .ZN(n5133)
         );
  AOI21_X1 U6249 ( .B1(n5193), .B2(n5802), .A(n5848), .ZN(n5130) );
  OAI21_X1 U6250 ( .B1(n5131), .B2(n5881), .A(n5130), .ZN(n5132) );
  AOI211_X1 U6251 ( .C1(n5170), .C2(n5134), .A(n5133), .B(n5132), .ZN(n5135)
         );
  OAI21_X1 U6252 ( .B1(n5190), .B2(n5830), .A(n5135), .ZN(U2813) );
  INV_X1 U6253 ( .A(EAX_REG_14__SCAN_IN), .ZN(n5137) );
  INV_X1 U6254 ( .A(DATAI_14_), .ZN(n5136) );
  OAI222_X1 U6255 ( .A1(n5190), .A2(n5413), .B1(n5905), .B2(n5137), .C1(n5136), 
        .C2(n5904), .ZN(U2877) );
  INV_X1 U6256 ( .A(n5138), .ZN(n5141) );
  INV_X1 U6257 ( .A(n5139), .ZN(n5140) );
  OAI21_X1 U6258 ( .B1(n5141), .B2(n5140), .A(n5151), .ZN(n5176) );
  AOI22_X1 U6259 ( .A1(n5142), .A2(DATAI_15_), .B1(EAX_REG_15__SCAN_IN), .B2(
        n5900), .ZN(n5143) );
  OAI21_X1 U6260 ( .B1(n5176), .B2(n5413), .A(n5143), .ZN(U2876) );
  NOR3_X1 U6261 ( .A1(REIP_REG_15__SCAN_IN), .A2(n5766), .A3(n5144), .ZN(n5169) );
  AOI22_X1 U6262 ( .A1(EBX_REG_15__SCAN_IN), .A2(n5879), .B1(
        REIP_REG_15__SCAN_IN), .B2(n5170), .ZN(n5145) );
  OAI211_X1 U6263 ( .C1(n5886), .C2(n3893), .A(n5145), .B(n5825), .ZN(n5148)
         );
  INV_X1 U6264 ( .A(n5146), .ZN(n5156) );
  XNOR2_X1 U6265 ( .A(n5104), .B(n5156), .ZN(n5699) );
  OAI22_X1 U6266 ( .A1(n5699), .A2(n5881), .B1(n5162), .B2(n5885), .ZN(n5147)
         );
  NOR3_X1 U6267 ( .A1(n5169), .A2(n5148), .A3(n5147), .ZN(n5149) );
  OAI21_X1 U6268 ( .B1(n5176), .B2(n5830), .A(n5149), .ZN(U2812) );
  AND2_X1 U6269 ( .A1(n5151), .A2(n5150), .ZN(n5153) );
  OR2_X1 U6270 ( .A1(n5153), .A2(n5207), .ZN(n5896) );
  INV_X1 U6271 ( .A(n5154), .ZN(n5155) );
  OAI21_X1 U6272 ( .B1(n5104), .B2(n5156), .A(n5155), .ZN(n5157) );
  NAND2_X1 U6273 ( .A1(n5157), .A2(n5209), .ZN(n5186) );
  OAI22_X1 U6274 ( .A1(n5186), .A2(n5378), .B1(n5167), .B2(n5892), .ZN(n5158)
         );
  INV_X1 U6275 ( .A(n5158), .ZN(n5159) );
  OAI21_X1 U6276 ( .B1(n5896), .B2(n3166), .A(n5159), .ZN(U2843) );
  XNOR2_X1 U6277 ( .A(n5452), .B(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5161)
         );
  XNOR2_X1 U6278 ( .A(n5160), .B(n5161), .ZN(n5703) );
  NAND2_X1 U6279 ( .A1(n5703), .A2(n6010), .ZN(n5165) );
  NOR2_X1 U6280 ( .A1(n6015), .A2(n6596), .ZN(n5700) );
  NOR2_X1 U6281 ( .A1(n6005), .A2(n5162), .ZN(n5163) );
  AOI211_X1 U6282 ( .C1(n6012), .C2(PHYADDRPOINTER_REG_15__SCAN_IN), .A(n5700), 
        .B(n5163), .ZN(n5164) );
  OAI211_X1 U6283 ( .C1(n6447), .C2(n5176), .A(n5165), .B(n5164), .ZN(U2971)
         );
  INV_X1 U6284 ( .A(REIP_REG_16__SCAN_IN), .ZN(n6746) );
  AOI22_X1 U6285 ( .A1(PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n5849), .B1(n5755), 
        .B2(n6746), .ZN(n5166) );
  OAI211_X1 U6286 ( .C1(n5862), .C2(n5167), .A(n5166), .B(n5825), .ZN(n5168)
         );
  AOI221_X1 U6287 ( .B1(n5170), .B2(REIP_REG_16__SCAN_IN), .C1(n5169), .C2(
        REIP_REG_16__SCAN_IN), .A(n5168), .ZN(n5174) );
  OAI22_X1 U6288 ( .A1(n5186), .A2(n5881), .B1(n5885), .B2(n5171), .ZN(n5172)
         );
  INV_X1 U6289 ( .A(n5172), .ZN(n5173) );
  OAI211_X1 U6290 ( .C1(n5896), .C2(n5830), .A(n5174), .B(n5173), .ZN(U2811)
         );
  INV_X1 U6291 ( .A(EBX_REG_15__SCAN_IN), .ZN(n5175) );
  OAI222_X1 U6292 ( .A1(n5176), .A2(n3166), .B1(n5175), .B2(n5892), .C1(n5378), 
        .C2(n5699), .ZN(U2844) );
  MUX2_X1 U6293 ( .A(n5627), .B(INSTADDRPOINTER_REG_16__SCAN_IN), .S(n5452), 
        .Z(n5178) );
  XNOR2_X1 U6294 ( .A(n5626), .B(n5178), .ZN(n5227) );
  INV_X1 U6295 ( .A(n5179), .ZN(n5698) );
  OAI21_X1 U6296 ( .B1(n5181), .B2(n5698), .A(n5180), .ZN(n5702) );
  OAI211_X1 U6297 ( .C1(INSTADDRPOINTER_REG_15__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .A(n5697), .B(n5698), .ZN(n5182) );
  INV_X1 U6298 ( .A(n5182), .ZN(n5184) );
  NAND2_X1 U6299 ( .A1(n5184), .A2(n5183), .ZN(n5185) );
  NAND2_X1 U6300 ( .A1(n6054), .A2(REIP_REG_16__SCAN_IN), .ZN(n5221) );
  OAI211_X1 U6301 ( .C1(n6058), .C2(n5186), .A(n5185), .B(n5221), .ZN(n5187)
         );
  AOI21_X1 U6302 ( .B1(n5702), .B2(INSTADDRPOINTER_REG_16__SCAN_IN), .A(n5187), 
        .ZN(n5188) );
  OAI21_X1 U6303 ( .B1(n5227), .B2(n6033), .A(n5188), .ZN(U3002) );
  OAI21_X1 U6304 ( .B1(n5989), .B2(n5128), .A(n5189), .ZN(n5192) );
  NOR2_X1 U6305 ( .A1(n5190), .A2(n6447), .ZN(n5191) );
  AOI211_X1 U6306 ( .C1(n5983), .C2(n5193), .A(n5192), .B(n5191), .ZN(n5194)
         );
  OAI21_X1 U6307 ( .B1(n5972), .B2(n5195), .A(n5194), .ZN(U2972) );
  NAND2_X1 U6308 ( .A1(n5200), .A2(n5199), .ZN(n5201) );
  AND2_X1 U6309 ( .A1(n5197), .A2(n5201), .ZN(n5748) );
  INV_X1 U6310 ( .A(n5748), .ZN(n5219) );
  AND2_X1 U6311 ( .A1(n5203), .A2(n5202), .ZN(n5204) );
  AOI22_X1 U6312 ( .A1(n5901), .A2(DATAI_2_), .B1(n5900), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n5206) );
  NAND2_X1 U6313 ( .A1(n5897), .A2(DATAI_18_), .ZN(n5205) );
  OAI211_X1 U6314 ( .C1(n5219), .C2(n5413), .A(n5206), .B(n5205), .ZN(U2873)
         );
  XOR2_X1 U6315 ( .A(n5208), .B(n5207), .Z(n5893) );
  INV_X1 U6316 ( .A(n5893), .ZN(n5213) );
  INV_X1 U6317 ( .A(EBX_REG_17__SCAN_IN), .ZN(n5212) );
  AOI21_X1 U6318 ( .B1(n5210), .B2(n5209), .A(n5217), .ZN(n5211) );
  INV_X1 U6319 ( .A(n5211), .ZN(n5764) );
  OAI222_X1 U6320 ( .A1(n5213), .A2(n3166), .B1(n5212), .B2(n5892), .C1(n5764), 
        .C2(n5378), .ZN(U2842) );
  INV_X1 U6321 ( .A(n5214), .ZN(n5215) );
  MUX2_X1 U6322 ( .A(n5297), .B(n5215), .S(n5298), .Z(n5216) );
  NAND2_X1 U6323 ( .A1(n5217), .A2(n5216), .ZN(n5308) );
  OR2_X1 U6324 ( .A1(n5217), .A2(n5216), .ZN(n5218) );
  NAND2_X1 U6325 ( .A1(n5308), .A2(n5218), .ZN(n5746) );
  OAI222_X1 U6326 ( .A1(n5746), .A2(n5378), .B1(n5220), .B2(n5892), .C1(n5219), 
        .C2(n3166), .ZN(U2841) );
  INV_X1 U6327 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5222) );
  OAI21_X1 U6328 ( .B1(n5989), .B2(n5222), .A(n5221), .ZN(n5224) );
  NOR2_X1 U6329 ( .A1(n5896), .A2(n6447), .ZN(n5223) );
  AOI211_X1 U6330 ( .C1(n5983), .C2(n5225), .A(n5224), .B(n5223), .ZN(n5226)
         );
  OAI21_X1 U6331 ( .B1(n5227), .B2(n5972), .A(n5226), .ZN(U2970) );
  INV_X1 U6332 ( .A(n5229), .ZN(n5231) );
  AOI211_X1 U6333 ( .C1(n5231), .C2(n4376), .A(n5230), .B(n5247), .ZN(n5233)
         );
  NOR2_X1 U6334 ( .A1(n5233), .A2(n5232), .ZN(n5493) );
  AOI22_X1 U6335 ( .A1(n5493), .A2(n5888), .B1(EBX_REG_29__SCAN_IN), .B2(n5379), .ZN(n5234) );
  OAI21_X1 U6336 ( .B1(n5228), .B2(n3166), .A(n5234), .ZN(U2830) );
  NOR2_X1 U6337 ( .A1(n5265), .A2(REIP_REG_29__SCAN_IN), .ZN(n5240) );
  INV_X1 U6338 ( .A(n5235), .ZN(n5552) );
  AOI22_X1 U6339 ( .A1(PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n5849), .B1(n5802), 
        .B2(n5236), .ZN(n5238) );
  NAND2_X1 U6340 ( .A1(n5879), .A2(EBX_REG_29__SCAN_IN), .ZN(n5237) );
  OAI211_X1 U6341 ( .C1(n5552), .C2(n6811), .A(n5238), .B(n5237), .ZN(n5239)
         );
  AOI211_X1 U6342 ( .C1(n5493), .C2(n5866), .A(n5240), .B(n5239), .ZN(n5241)
         );
  OAI21_X1 U6343 ( .B1(n5228), .B2(n5830), .A(n5241), .ZN(U2798) );
  AOI22_X1 U6344 ( .A1(n5897), .A2(DATAI_29_), .B1(n5900), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n5243) );
  NAND2_X1 U6345 ( .A1(n5901), .A2(DATAI_13_), .ZN(n5242) );
  OAI211_X1 U6346 ( .C1(n5228), .C2(n5413), .A(n5243), .B(n5242), .ZN(U2862)
         );
  NAND2_X1 U6347 ( .A1(REIP_REG_29__SCAN_IN), .A2(n5415), .ZN(n5264) );
  INV_X1 U6348 ( .A(n5425), .ZN(n5246) );
  NAND2_X1 U6349 ( .A1(n5246), .A2(n5804), .ZN(n5263) );
  INV_X1 U6350 ( .A(n5252), .ZN(n5249) );
  NAND2_X1 U6351 ( .A1(n5253), .A2(n5247), .ZN(n5248) );
  NAND3_X1 U6352 ( .A1(n5250), .A2(n5249), .A3(n5248), .ZN(n5255) );
  NAND2_X1 U6353 ( .A1(n5326), .A2(n5298), .ZN(n5251) );
  NAND3_X1 U6354 ( .A1(n5253), .A2(n5252), .A3(n5251), .ZN(n5254) );
  INV_X1 U6355 ( .A(EBX_REG_30__SCAN_IN), .ZN(n5318) );
  NOR2_X1 U6356 ( .A1(n5256), .A2(n5415), .ZN(n5259) );
  OAI22_X1 U6357 ( .A1(n5257), .A2(n5886), .B1(n5416), .B2(n5885), .ZN(n5258)
         );
  NOR2_X1 U6358 ( .A1(n5259), .A2(n5258), .ZN(n5260) );
  OAI21_X1 U6359 ( .B1(n5862), .B2(n5318), .A(n5260), .ZN(n5261) );
  AOI21_X1 U6360 ( .B1(n5486), .B2(n5866), .A(n5261), .ZN(n5262) );
  OAI211_X1 U6361 ( .C1(n5265), .C2(n5264), .A(n5263), .B(n5262), .ZN(U2797)
         );
  INV_X1 U6362 ( .A(n5320), .ZN(n5267) );
  AOI21_X1 U6363 ( .B1(n5268), .B2(n5334), .A(n5267), .ZN(n5442) );
  INV_X1 U6364 ( .A(n5442), .ZN(n5392) );
  INV_X1 U6365 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6875) );
  AOI22_X1 U6366 ( .A1(EBX_REG_27__SCAN_IN), .A2(n5879), .B1(
        PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n5849), .ZN(n5269) );
  OAI21_X1 U6367 ( .B1(n5560), .B2(n6875), .A(n5269), .ZN(n5273) );
  AOI21_X1 U6368 ( .B1(n5270), .B2(n5340), .A(n5324), .ZN(n5640) );
  INV_X1 U6369 ( .A(n5640), .ZN(n5330) );
  INV_X1 U6370 ( .A(n5271), .ZN(n5440) );
  OAI22_X1 U6371 ( .A1(n5330), .A2(n5881), .B1(n5440), .B2(n5885), .ZN(n5272)
         );
  AOI211_X1 U6372 ( .C1(n6875), .C2(n5555), .A(n5273), .B(n5272), .ZN(n5274)
         );
  OAI21_X1 U6373 ( .B1(n5392), .B2(n5830), .A(n5274), .ZN(U2800) );
  AND2_X1 U6374 ( .A1(n5363), .A2(n5276), .ZN(n5278) );
  NOR2_X1 U6375 ( .A1(n5365), .A2(n5277), .ZN(n5351) );
  INV_X1 U6376 ( .A(n5595), .ZN(n5584) );
  NAND2_X1 U6377 ( .A1(REIP_REG_22__SCAN_IN), .A2(REIP_REG_21__SCAN_IN), .ZN(
        n5279) );
  OAI21_X1 U6378 ( .B1(n5584), .B2(n5279), .A(n6842), .ZN(n5287) );
  INV_X1 U6379 ( .A(n5374), .ZN(n5282) );
  AOI21_X1 U6380 ( .B1(n5282), .B2(n5281), .A(n5280), .ZN(n5283) );
  OR2_X1 U6381 ( .A1(n5283), .A2(n5356), .ZN(n5535) );
  OAI22_X1 U6382 ( .A1(n5360), .A2(n5862), .B1(n5462), .B2(n5886), .ZN(n5284)
         );
  AOI21_X1 U6383 ( .B1(n5466), .B2(n5802), .A(n5284), .ZN(n5285) );
  OAI21_X1 U6384 ( .B1(n5535), .B2(n5881), .A(n5285), .ZN(n5286) );
  AOI21_X1 U6385 ( .B1(n5287), .B2(n5577), .A(n5286), .ZN(n5288) );
  OAI21_X1 U6386 ( .B1(n5463), .B2(n5830), .A(n5288), .ZN(U2804) );
  INV_X1 U6387 ( .A(n5289), .ZN(n5293) );
  INV_X1 U6388 ( .A(n5291), .ZN(n5292) );
  AOI21_X1 U6389 ( .B1(n5293), .B2(n5292), .A(n5370), .ZN(n5613) );
  INV_X1 U6390 ( .A(n5613), .ZN(n5410) );
  NAND2_X1 U6391 ( .A1(REIP_REG_19__SCAN_IN), .A2(REIP_REG_18__SCAN_IN), .ZN(
        n5294) );
  INV_X1 U6392 ( .A(REIP_REG_20__SCAN_IN), .ZN(n6600) );
  OAI21_X1 U6393 ( .B1(n5749), .B2(n5294), .A(n6600), .ZN(n5304) );
  NOR2_X1 U6394 ( .A1(n5876), .A2(n5295), .ZN(n5593) );
  MUX2_X1 U6395 ( .A(n5298), .B(n5297), .S(n5296), .Z(n5300) );
  XNOR2_X1 U6396 ( .A(n5300), .B(n5299), .ZN(n5669) );
  INV_X1 U6397 ( .A(n5669), .ZN(n5377) );
  OAI22_X1 U6398 ( .A1(n5376), .A2(n5862), .B1(n5616), .B2(n5885), .ZN(n5301)
         );
  AOI21_X1 U6399 ( .B1(n5849), .B2(PHYADDRPOINTER_REG_20__SCAN_IN), .A(n5301), 
        .ZN(n5302) );
  OAI21_X1 U6400 ( .B1(n5377), .B2(n5881), .A(n5302), .ZN(n5303) );
  AOI21_X1 U6401 ( .B1(n5304), .B2(n5593), .A(n5303), .ZN(n5305) );
  OAI21_X1 U6402 ( .B1(n5410), .B2(n5830), .A(n5305), .ZN(U2807) );
  AOI21_X1 U6403 ( .B1(n5306), .B2(n5197), .A(n5291), .ZN(n5482) );
  INV_X1 U6404 ( .A(n5482), .ZN(n5414) );
  XNOR2_X1 U6405 ( .A(n5308), .B(n5307), .ZN(n5676) );
  AOI21_X1 U6406 ( .B1(n5849), .B2(PHYADDRPOINTER_REG_19__SCAN_IN), .A(n5848), 
        .ZN(n5311) );
  INV_X1 U6407 ( .A(n5309), .ZN(n5757) );
  AOI21_X1 U6408 ( .B1(REIP_REG_18__SCAN_IN), .B2(n5757), .A(n5876), .ZN(n5750) );
  AOI22_X1 U6409 ( .A1(n5478), .A2(n5802), .B1(REIP_REG_19__SCAN_IN), .B2(
        n5750), .ZN(n5310) );
  OAI211_X1 U6410 ( .C1(n5312), .C2(n5862), .A(n5311), .B(n5310), .ZN(n5314)
         );
  INV_X1 U6411 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6854) );
  NOR3_X1 U6412 ( .A1(REIP_REG_19__SCAN_IN), .A2(n5749), .A3(n6854), .ZN(n5313) );
  AOI211_X1 U6413 ( .C1(n5676), .C2(n5866), .A(n5314), .B(n5313), .ZN(n5315)
         );
  OAI21_X1 U6414 ( .B1(n5414), .B2(n5830), .A(n5315), .ZN(U2808) );
  OAI22_X1 U6415 ( .A1(n5316), .A2(n5378), .B1(n4445), .B2(n5892), .ZN(U2828)
         );
  INV_X1 U6416 ( .A(n5486), .ZN(n5317) );
  OAI222_X1 U6417 ( .A1(n3166), .A2(n5425), .B1(n5318), .B2(n5892), .C1(n5317), 
        .C2(n5378), .ZN(U2829) );
  AND2_X1 U6418 ( .A1(n5320), .A2(n5319), .ZN(n5322) );
  OR2_X1 U6419 ( .A1(n5322), .A2(n5321), .ZN(n5431) );
  OR2_X1 U6420 ( .A1(n5324), .A2(n5323), .ZN(n5325) );
  NAND2_X1 U6421 ( .A1(n5326), .A2(n5325), .ZN(n5558) );
  OAI22_X1 U6422 ( .A1(n5558), .A2(n5378), .B1(n5327), .B2(n5892), .ZN(n5328)
         );
  INV_X1 U6423 ( .A(n5328), .ZN(n5329) );
  OAI21_X1 U6424 ( .B1(n5431), .B2(n3166), .A(n5329), .ZN(U2831) );
  INV_X1 U6425 ( .A(EBX_REG_27__SCAN_IN), .ZN(n5331) );
  OAI222_X1 U6426 ( .A1(n3166), .A2(n5392), .B1(n5331), .B2(n5892), .C1(n5330), 
        .C2(n5378), .ZN(U2832) );
  INV_X1 U6427 ( .A(n5334), .ZN(n5335) );
  AOI21_X1 U6428 ( .B1(n5336), .B2(n5333), .A(n5335), .ZN(n5601) );
  INV_X1 U6429 ( .A(n5601), .ZN(n5395) );
  NAND2_X1 U6430 ( .A1(n5337), .A2(n5338), .ZN(n5339) );
  NAND2_X1 U6431 ( .A1(n5340), .A2(n5339), .ZN(n5559) );
  OAI22_X1 U6432 ( .A1(n5559), .A2(n5378), .B1(n5341), .B2(n5892), .ZN(n5342)
         );
  INV_X1 U6433 ( .A(n5342), .ZN(n5343) );
  OAI21_X1 U6434 ( .B1(n5395), .B2(n3166), .A(n5343), .ZN(U2833) );
  AND2_X1 U6435 ( .A1(n5370), .A2(n5368), .ZN(n5345) );
  OR2_X1 U6436 ( .A1(n5352), .A2(n5346), .ZN(n5347) );
  AND2_X1 U6437 ( .A1(n5333), .A2(n5347), .ZN(n5568) );
  INV_X1 U6438 ( .A(EBX_REG_25__SCAN_IN), .ZN(n5350) );
  OR2_X1 U6439 ( .A1(n5358), .A2(n5348), .ZN(n5349) );
  NAND2_X1 U6440 ( .A1(n5337), .A2(n5349), .ZN(n5649) );
  OAI222_X1 U6441 ( .A1(n5450), .A2(n3166), .B1(n5350), .B2(n5892), .C1(n5378), 
        .C2(n5649), .ZN(U2834) );
  INV_X1 U6442 ( .A(n5351), .ZN(n5353) );
  AOI21_X1 U6443 ( .B1(n5354), .B2(n5353), .A(n5352), .ZN(n5458) );
  INV_X1 U6444 ( .A(n5458), .ZN(n5579) );
  INV_X1 U6445 ( .A(EBX_REG_24__SCAN_IN), .ZN(n5359) );
  NOR2_X1 U6446 ( .A1(n5356), .A2(n5355), .ZN(n5357) );
  OR2_X1 U6447 ( .A1(n5358), .A2(n5357), .ZN(n5583) );
  OAI222_X1 U6448 ( .A1(n3166), .A2(n5579), .B1(n5892), .B2(n5359), .C1(n5583), 
        .C2(n5378), .ZN(U2835) );
  OAI22_X1 U6449 ( .A1(n5535), .A2(n5378), .B1(n5360), .B2(n5892), .ZN(n5361)
         );
  INV_X1 U6450 ( .A(n5361), .ZN(n5362) );
  OAI21_X1 U6451 ( .B1(n5463), .B2(n3166), .A(n5362), .ZN(U2836) );
  INV_X1 U6452 ( .A(n5363), .ZN(n5364) );
  AOI21_X1 U6453 ( .B1(n5366), .B2(n5365), .A(n5364), .ZN(n5605) );
  INV_X1 U6454 ( .A(n5605), .ZN(n5404) );
  AOI22_X1 U6455 ( .A1(n5588), .A2(n5888), .B1(EBX_REG_22__SCAN_IN), .B2(n5379), .ZN(n5367) );
  OAI21_X1 U6456 ( .B1(n5404), .B2(n3166), .A(n5367), .ZN(U2837) );
  INV_X1 U6457 ( .A(n5368), .ZN(n5369) );
  XNOR2_X1 U6458 ( .A(n5370), .B(n5369), .ZN(n5594) );
  INV_X1 U6459 ( .A(n5594), .ZN(n5407) );
  NAND2_X1 U6460 ( .A1(n5372), .A2(n5371), .ZN(n5373) );
  AND2_X1 U6461 ( .A1(n5374), .A2(n5373), .ZN(n5657) );
  AOI22_X1 U6462 ( .A1(n5657), .A2(n5888), .B1(EBX_REG_21__SCAN_IN), .B2(n5379), .ZN(n5375) );
  OAI21_X1 U6463 ( .B1(n5407), .B2(n3166), .A(n5375), .ZN(U2838) );
  OAI222_X1 U6464 ( .A1(n5378), .A2(n5377), .B1(n5376), .B2(n5892), .C1(n3166), 
        .C2(n5410), .ZN(U2839) );
  AOI22_X1 U6465 ( .A1(n5676), .A2(n5888), .B1(EBX_REG_19__SCAN_IN), .B2(n5379), .ZN(n5380) );
  OAI21_X1 U6466 ( .B1(n5414), .B2(n3166), .A(n5380), .ZN(U2840) );
  AND2_X1 U6467 ( .A1(n5905), .A2(n5381), .ZN(n5382) );
  NAND2_X1 U6468 ( .A1(n5383), .A2(n5382), .ZN(n5385) );
  AOI22_X1 U6469 ( .A1(n5897), .A2(DATAI_31_), .B1(n5900), .B2(
        EAX_REG_31__SCAN_IN), .ZN(n5384) );
  NAND2_X1 U6470 ( .A1(n5385), .A2(n5384), .ZN(U2860) );
  AOI22_X1 U6471 ( .A1(n5897), .A2(DATAI_30_), .B1(n5900), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n5387) );
  NAND2_X1 U6472 ( .A1(n5901), .A2(DATAI_14_), .ZN(n5386) );
  OAI211_X1 U6473 ( .C1(n5425), .C2(n5413), .A(n5387), .B(n5386), .ZN(U2861)
         );
  AOI22_X1 U6474 ( .A1(n5901), .A2(DATAI_12_), .B1(n5900), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n5389) );
  NAND2_X1 U6475 ( .A1(n5897), .A2(DATAI_28_), .ZN(n5388) );
  OAI211_X1 U6476 ( .C1(n5431), .C2(n5413), .A(n5389), .B(n5388), .ZN(U2863)
         );
  AOI22_X1 U6477 ( .A1(n5897), .A2(DATAI_27_), .B1(n5900), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n5391) );
  NAND2_X1 U6478 ( .A1(n5901), .A2(DATAI_11_), .ZN(n5390) );
  OAI211_X1 U6479 ( .C1(n5392), .C2(n5413), .A(n5391), .B(n5390), .ZN(U2864)
         );
  AOI22_X1 U6480 ( .A1(n5901), .A2(DATAI_10_), .B1(n5900), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n5394) );
  NAND2_X1 U6481 ( .A1(n5897), .A2(DATAI_26_), .ZN(n5393) );
  OAI211_X1 U6482 ( .C1(n5395), .C2(n5413), .A(n5394), .B(n5393), .ZN(U2865)
         );
  AOI22_X1 U6483 ( .A1(n5901), .A2(DATAI_9_), .B1(n5900), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n5397) );
  NAND2_X1 U6484 ( .A1(n5897), .A2(DATAI_25_), .ZN(n5396) );
  OAI211_X1 U6485 ( .C1(n5450), .C2(n5413), .A(n5397), .B(n5396), .ZN(U2866)
         );
  AOI22_X1 U6486 ( .A1(n5901), .A2(DATAI_8_), .B1(n5900), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n5399) );
  NAND2_X1 U6487 ( .A1(n5897), .A2(DATAI_24_), .ZN(n5398) );
  OAI211_X1 U6488 ( .C1(n5579), .C2(n5413), .A(n5399), .B(n5398), .ZN(U2867)
         );
  AOI22_X1 U6489 ( .A1(n5897), .A2(DATAI_23_), .B1(n5900), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n5401) );
  NAND2_X1 U6490 ( .A1(n5901), .A2(DATAI_7_), .ZN(n5400) );
  OAI211_X1 U6491 ( .C1(n5463), .C2(n5413), .A(n5401), .B(n5400), .ZN(U2868)
         );
  AOI22_X1 U6492 ( .A1(n5901), .A2(DATAI_6_), .B1(n5900), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n5403) );
  NAND2_X1 U6493 ( .A1(n5897), .A2(DATAI_22_), .ZN(n5402) );
  OAI211_X1 U6494 ( .C1(n5404), .C2(n5413), .A(n5403), .B(n5402), .ZN(U2869)
         );
  AOI22_X1 U6495 ( .A1(n5901), .A2(DATAI_5_), .B1(n5900), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n5406) );
  NAND2_X1 U6496 ( .A1(n5897), .A2(DATAI_21_), .ZN(n5405) );
  OAI211_X1 U6497 ( .C1(n5407), .C2(n5413), .A(n5406), .B(n5405), .ZN(U2870)
         );
  AOI22_X1 U6498 ( .A1(n5901), .A2(DATAI_4_), .B1(n5900), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n5409) );
  NAND2_X1 U6499 ( .A1(n5897), .A2(DATAI_20_), .ZN(n5408) );
  OAI211_X1 U6500 ( .C1(n5410), .C2(n5413), .A(n5409), .B(n5408), .ZN(U2871)
         );
  AOI22_X1 U6501 ( .A1(n5897), .A2(DATAI_19_), .B1(n5900), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n5412) );
  NAND2_X1 U6502 ( .A1(n5901), .A2(DATAI_3_), .ZN(n5411) );
  OAI211_X1 U6503 ( .C1(n5414), .C2(n5413), .A(n5412), .B(n5411), .ZN(U2872)
         );
  NOR2_X1 U6504 ( .A1(n6015), .A2(n5415), .ZN(n5485) );
  NOR2_X1 U6505 ( .A1(n6005), .A2(n5416), .ZN(n5417) );
  AOI211_X1 U6506 ( .C1(n6012), .C2(PHYADDRPOINTER_REG_30__SCAN_IN), .A(n5485), 
        .B(n5417), .ZN(n5424) );
  INV_X1 U6507 ( .A(n5418), .ZN(n5420) );
  OAI21_X1 U6508 ( .B1(n5513), .B2(n5420), .A(n5419), .ZN(n5422) );
  XNOR2_X1 U6509 ( .A(n5422), .B(n5421), .ZN(n5484) );
  NAND2_X1 U6510 ( .A1(n5484), .A2(n6010), .ZN(n5423) );
  OAI211_X1 U6511 ( .C1(n5425), .C2(n6447), .A(n5424), .B(n5423), .ZN(U2956)
         );
  NAND3_X1 U6512 ( .A1(n5513), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .A3(n5452), .ZN(n5429) );
  AND2_X1 U6513 ( .A1(n5511), .A2(n5427), .ZN(n5428) );
  NAND2_X1 U6514 ( .A1(n5446), .A2(n5428), .ZN(n5436) );
  AOI22_X1 U6515 ( .A1(n5429), .A2(n5436), .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n5521), .ZN(n5430) );
  XNOR2_X1 U6516 ( .A(n5430), .B(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5509)
         );
  INV_X1 U6517 ( .A(n5431), .ZN(n5554) );
  INV_X1 U6518 ( .A(n5432), .ZN(n5548) );
  NAND2_X1 U6519 ( .A1(n6054), .A2(REIP_REG_28__SCAN_IN), .ZN(n5505) );
  NAND2_X1 U6520 ( .A1(n6012), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5433)
         );
  OAI211_X1 U6521 ( .C1(n6005), .C2(n5548), .A(n5505), .B(n5433), .ZN(n5434)
         );
  AOI21_X1 U6522 ( .B1(n5554), .B2(n3167), .A(n5434), .ZN(n5435) );
  OAI21_X1 U6523 ( .B1(n5972), .B2(n5509), .A(n5435), .ZN(U2958) );
  NAND2_X1 U6524 ( .A1(n5437), .A2(n5436), .ZN(n5438) );
  XNOR2_X1 U6525 ( .A(n5438), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5639)
         );
  AOI22_X1 U6526 ( .A1(n6012), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .B1(n6054), 
        .B2(REIP_REG_27__SCAN_IN), .ZN(n5439) );
  OAI21_X1 U6527 ( .B1(n5440), .B2(n6005), .A(n5439), .ZN(n5441) );
  AOI21_X1 U6528 ( .B1(n5442), .B2(n3167), .A(n5441), .ZN(n5443) );
  OAI21_X1 U6529 ( .B1(n5639), .B2(n5972), .A(n5443), .ZN(U2959) );
  INV_X1 U6530 ( .A(REIP_REG_25__SCAN_IN), .ZN(n5444) );
  OAI22_X1 U6531 ( .A1(n5989), .A2(n4101), .B1(n6015), .B2(n5444), .ZN(n5445)
         );
  AOI21_X1 U6532 ( .B1(n5983), .B2(n5566), .A(n5445), .ZN(n5449) );
  OAI21_X1 U6533 ( .B1(n5447), .B2(n5446), .A(n4197), .ZN(n5651) );
  NAND2_X1 U6534 ( .A1(n5651), .A2(n6010), .ZN(n5448) );
  OAI211_X1 U6535 ( .C1(n5450), .C2(n6447), .A(n5449), .B(n5448), .ZN(U2961)
         );
  INV_X1 U6536 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5451) );
  NAND3_X1 U6537 ( .A1(n5468), .A2(n4388), .A3(n5451), .ZN(n5460) );
  NAND3_X1 U6538 ( .A1(n5452), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5453) );
  XNOR2_X1 U6539 ( .A(n5455), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5530)
         );
  NAND2_X1 U6540 ( .A1(n6054), .A2(REIP_REG_24__SCAN_IN), .ZN(n5522) );
  NAND2_X1 U6541 ( .A1(n6012), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5456)
         );
  OAI211_X1 U6542 ( .C1(n5575), .C2(n6005), .A(n5522), .B(n5456), .ZN(n5457)
         );
  AOI21_X1 U6543 ( .B1(n5458), .B2(n3167), .A(n5457), .ZN(n5459) );
  OAI21_X1 U6544 ( .B1(n5530), .B2(n5972), .A(n5459), .ZN(U2962) );
  OAI21_X1 U6545 ( .B1(n5475), .B2(n5523), .A(n5460), .ZN(n5461) );
  XNOR2_X1 U6546 ( .A(n5461), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5539)
         );
  NAND2_X1 U6547 ( .A1(n6054), .A2(REIP_REG_23__SCAN_IN), .ZN(n5533) );
  OAI21_X1 U6548 ( .B1(n5989), .B2(n5462), .A(n5533), .ZN(n5465) );
  NOR2_X1 U6549 ( .A1(n5463), .A2(n6447), .ZN(n5464) );
  AOI211_X1 U6550 ( .C1(n5983), .C2(n5466), .A(n5465), .B(n5464), .ZN(n5467)
         );
  OAI21_X1 U6551 ( .B1(n5539), .B2(n5972), .A(n5467), .ZN(U2963) );
  AOI21_X1 U6552 ( .B1(n5470), .B2(n5469), .A(n5468), .ZN(n5656) );
  INV_X1 U6553 ( .A(n5592), .ZN(n5472) );
  AOI22_X1 U6554 ( .A1(n6012), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .B1(n6054), 
        .B2(REIP_REG_21__SCAN_IN), .ZN(n5471) );
  OAI21_X1 U6555 ( .B1(n5472), .B2(n6005), .A(n5471), .ZN(n5473) );
  AOI21_X1 U6556 ( .B1(n5594), .B2(n3167), .A(n5473), .ZN(n5474) );
  OAI21_X1 U6557 ( .B1(n5656), .B2(n5972), .A(n5474), .ZN(U2965) );
  OAI21_X1 U6558 ( .B1(n5477), .B2(n5476), .A(n5475), .ZN(n5675) );
  INV_X1 U6559 ( .A(n5478), .ZN(n5480) );
  AOI22_X1 U6560 ( .A1(n6012), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .B1(n6054), 
        .B2(REIP_REG_19__SCAN_IN), .ZN(n5479) );
  OAI21_X1 U6561 ( .B1(n5480), .B2(n6005), .A(n5479), .ZN(n5481) );
  AOI21_X1 U6562 ( .B1(n5482), .B2(n3167), .A(n5481), .ZN(n5483) );
  OAI21_X1 U6563 ( .B1(n5972), .B2(n5675), .A(n5483), .ZN(U2967) );
  INV_X1 U6564 ( .A(n5484), .ZN(n5491) );
  AOI21_X1 U6565 ( .B1(n5486), .B2(n6041), .A(n5485), .ZN(n5490) );
  OAI21_X1 U6566 ( .B1(INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n5488), .A(n5487), 
        .ZN(n5489) );
  OAI211_X1 U6567 ( .C1(n5491), .C2(n6033), .A(n5490), .B(n5489), .ZN(U2988)
         );
  INV_X1 U6568 ( .A(n5492), .ZN(n5499) );
  INV_X1 U6569 ( .A(n5493), .ZN(n5497) );
  INV_X1 U6570 ( .A(n5504), .ZN(n5644) );
  NAND3_X1 U6571 ( .A1(n5644), .A2(n5502), .A3(n5494), .ZN(n5495) );
  OAI211_X1 U6572 ( .C1(n5497), .C2(n6058), .A(n5496), .B(n5495), .ZN(n5498)
         );
  AOI21_X1 U6573 ( .B1(INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n5499), .A(n5498), 
        .ZN(n5500) );
  OAI21_X1 U6574 ( .B1(n5501), .B2(n6033), .A(n5500), .ZN(U2989) );
  NOR3_X1 U6575 ( .A1(n5504), .A2(n5503), .A3(n5502), .ZN(n5507) );
  OAI21_X1 U6576 ( .B1(n5558), .B2(n6058), .A(n5505), .ZN(n5506) );
  AOI211_X1 U6577 ( .C1(n5645), .C2(INSTADDRPOINTER_REG_28__SCAN_IN), .A(n5507), .B(n5506), .ZN(n5508) );
  OAI21_X1 U6578 ( .B1(n5509), .B2(n6033), .A(n5508), .ZN(U2990) );
  NOR2_X1 U6579 ( .A1(n5511), .A2(n5510), .ZN(n5512) );
  XNOR2_X1 U6580 ( .A(n5513), .B(n5512), .ZN(n5600) );
  NAND2_X1 U6581 ( .A1(n5600), .A2(n6060), .ZN(n5520) );
  OAI21_X1 U6582 ( .B1(INSTADDRPOINTER_REG_26__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .A(n5648), .ZN(n5514) );
  INV_X1 U6583 ( .A(n5514), .ZN(n5517) );
  INV_X1 U6584 ( .A(REIP_REG_26__SCAN_IN), .ZN(n5515) );
  OAI22_X1 U6585 ( .A1(n5559), .A2(n6058), .B1(n6015), .B2(n5515), .ZN(n5516)
         );
  AOI21_X1 U6586 ( .B1(n5518), .B2(n5517), .A(n5516), .ZN(n5519) );
  OAI211_X1 U6587 ( .C1(n5654), .C2(n5521), .A(n5520), .B(n5519), .ZN(U2992)
         );
  INV_X1 U6588 ( .A(n5583), .ZN(n5528) );
  INV_X1 U6589 ( .A(n5522), .ZN(n5527) );
  INV_X1 U6590 ( .A(n5523), .ZN(n5532) );
  NAND3_X1 U6591 ( .A1(n5674), .A2(n5532), .A3(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5524) );
  AOI21_X1 U6592 ( .B1(n5525), .B2(n5524), .A(n5654), .ZN(n5526) );
  AOI211_X1 U6593 ( .C1(n6041), .C2(n5528), .A(n5527), .B(n5526), .ZN(n5529)
         );
  OAI21_X1 U6594 ( .B1(n5530), .B2(n6033), .A(n5529), .ZN(U2994) );
  NAND3_X1 U6595 ( .A1(n5674), .A2(n5532), .A3(n5531), .ZN(n5534) );
  OAI211_X1 U6596 ( .C1(n5535), .C2(n6058), .A(n5534), .B(n5533), .ZN(n5536)
         );
  AOI21_X1 U6597 ( .B1(n5537), .B2(INSTADDRPOINTER_REG_23__SCAN_IN), .A(n5536), 
        .ZN(n5538) );
  OAI21_X1 U6598 ( .B1(n5539), .B2(n6033), .A(n5538), .ZN(U2995) );
  OAI211_X1 U6599 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n4666), .A(n5542), .B(
        n6405), .ZN(n5540) );
  OAI21_X1 U6600 ( .B1(n3184), .B2(n6071), .A(n5540), .ZN(n5541) );
  MUX2_X1 U6601 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n5541), .S(n6066), 
        .Z(U3464) );
  XNOR2_X1 U6602 ( .A(n5542), .B(n6068), .ZN(n5543) );
  OAI22_X1 U6603 ( .A1(n5543), .A2(n6643), .B1(n4533), .B2(n3184), .ZN(n5544)
         );
  MUX2_X1 U6604 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n5544), .S(n6066), 
        .Z(U3463) );
  OR2_X1 U6605 ( .A1(n5545), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6645) );
  INV_X2 U6606 ( .A(n6645), .ZN(n6536) );
  AOI21_X1 U6607 ( .B1(n6511), .B2(n6540), .A(n6566), .ZN(n5547) );
  AND2_X1 U6608 ( .A1(n5547), .A2(n5546), .ZN(n5937) );
  AND2_X1 U6609 ( .A1(n5952), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  INV_X1 U6610 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6741) );
  INV_X1 U6611 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5549) );
  OAI22_X1 U6612 ( .A1(n5549), .A2(n5886), .B1(n5885), .B2(n5548), .ZN(n5550)
         );
  AOI21_X1 U6613 ( .B1(n5879), .B2(EBX_REG_28__SCAN_IN), .A(n5550), .ZN(n5551)
         );
  OAI21_X1 U6614 ( .B1(n5552), .B2(n6741), .A(n5551), .ZN(n5553) );
  AOI21_X1 U6615 ( .B1(n5554), .B2(n5804), .A(n5553), .ZN(n5557) );
  NAND3_X1 U6616 ( .A1(REIP_REG_27__SCAN_IN), .A2(n5555), .A3(n6741), .ZN(
        n5556) );
  OAI211_X1 U6617 ( .C1(n5881), .C2(n5558), .A(n5557), .B(n5556), .ZN(U2799)
         );
  AOI22_X1 U6618 ( .A1(EBX_REG_26__SCAN_IN), .A2(n5879), .B1(
        PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n5849), .ZN(n5564) );
  INV_X1 U6619 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6791) );
  NOR2_X1 U6620 ( .A1(n6791), .A2(n5569), .ZN(n5565) );
  AOI21_X1 U6621 ( .B1(REIP_REG_25__SCAN_IN), .B2(n5565), .A(
        REIP_REG_26__SCAN_IN), .ZN(n5561) );
  OAI22_X1 U6622 ( .A1(n5561), .A2(n5560), .B1(n5559), .B2(n5881), .ZN(n5562)
         );
  AOI21_X1 U6623 ( .B1(n5601), .B2(n5804), .A(n5562), .ZN(n5563) );
  OAI211_X1 U6624 ( .C1(n5604), .C2(n5885), .A(n5564), .B(n5563), .ZN(U2801)
         );
  AOI22_X1 U6625 ( .A1(EBX_REG_25__SCAN_IN), .A2(n5879), .B1(
        PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n5849), .ZN(n5573) );
  AOI22_X1 U6626 ( .A1(n5566), .A2(n5802), .B1(n5565), .B2(n5444), .ZN(n5572)
         );
  NOR2_X1 U6627 ( .A1(n5649), .A2(n5881), .ZN(n5567) );
  AOI21_X1 U6628 ( .B1(n5568), .B2(n5804), .A(n5567), .ZN(n5571) );
  NOR2_X1 U6629 ( .A1(REIP_REG_24__SCAN_IN), .A2(n5569), .ZN(n5580) );
  OAI21_X1 U6630 ( .B1(n5577), .B2(n5580), .A(REIP_REG_25__SCAN_IN), .ZN(n5570) );
  NAND4_X1 U6631 ( .A1(n5573), .A2(n5572), .A3(n5571), .A4(n5570), .ZN(U2802)
         );
  AOI22_X1 U6632 ( .A1(n5879), .A2(EBX_REG_24__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n5849), .ZN(n5574) );
  OAI21_X1 U6633 ( .B1(n5575), .B2(n5885), .A(n5574), .ZN(n5576) );
  AOI21_X1 U6634 ( .B1(n5577), .B2(REIP_REG_24__SCAN_IN), .A(n5576), .ZN(n5578) );
  OAI21_X1 U6635 ( .B1(n5579), .B2(n5830), .A(n5578), .ZN(n5581) );
  NOR2_X1 U6636 ( .A1(n5581), .A2(n5580), .ZN(n5582) );
  OAI21_X1 U6637 ( .B1(n5583), .B2(n5881), .A(n5582), .ZN(U2803) );
  AOI21_X1 U6638 ( .B1(n5595), .B2(n6972), .A(n5593), .ZN(n5591) );
  NOR3_X1 U6639 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6972), .A3(n5584), .ZN(n5587) );
  INV_X1 U6640 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5585) );
  OAI22_X1 U6641 ( .A1(n5585), .A2(n5886), .B1(n5610), .B2(n5885), .ZN(n5586)
         );
  AOI211_X1 U6642 ( .C1(n5879), .C2(EBX_REG_22__SCAN_IN), .A(n5587), .B(n5586), 
        .ZN(n5590) );
  AOI22_X1 U6643 ( .A1(n5605), .A2(n5804), .B1(n5866), .B2(n5588), .ZN(n5589)
         );
  OAI211_X1 U6644 ( .C1(n5591), .C2(n6871), .A(n5590), .B(n5589), .ZN(U2805)
         );
  AOI22_X1 U6645 ( .A1(PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n5849), .B1(n5592), 
        .B2(n5802), .ZN(n5599) );
  AOI22_X1 U6646 ( .A1(EBX_REG_21__SCAN_IN), .A2(n5879), .B1(
        REIP_REG_21__SCAN_IN), .B2(n5593), .ZN(n5598) );
  AOI22_X1 U6647 ( .A1(n5594), .A2(n5804), .B1(n5657), .B2(n5866), .ZN(n5597)
         );
  NAND2_X1 U6648 ( .A1(n5595), .A2(n6972), .ZN(n5596) );
  NAND4_X1 U6649 ( .A1(n5599), .A2(n5598), .A3(n5597), .A4(n5596), .ZN(U2806)
         );
  AOI22_X1 U6650 ( .A1(n6054), .A2(REIP_REG_26__SCAN_IN), .B1(n6012), .B2(
        PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5603) );
  AOI22_X1 U6651 ( .A1(n5601), .A2(n3167), .B1(n6010), .B2(n5600), .ZN(n5602)
         );
  OAI211_X1 U6652 ( .C1(n6005), .C2(n5604), .A(n5603), .B(n5602), .ZN(U2960)
         );
  AOI22_X1 U6653 ( .A1(n6054), .A2(REIP_REG_22__SCAN_IN), .B1(n6012), .B2(
        PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5609) );
  AOI21_X1 U6654 ( .B1(n5607), .B2(n6010), .A(n5606), .ZN(n5608) );
  OAI211_X1 U6655 ( .C1(n6005), .C2(n5610), .A(n5609), .B(n5608), .ZN(U2964)
         );
  AOI22_X1 U6656 ( .A1(n6054), .A2(REIP_REG_20__SCAN_IN), .B1(n6012), .B2(
        PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5615) );
  XNOR2_X1 U6657 ( .A(n3636), .B(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5611)
         );
  XNOR2_X1 U6658 ( .A(n5612), .B(n5611), .ZN(n5670) );
  AOI22_X1 U6659 ( .A1(n6010), .A2(n5670), .B1(n5613), .B2(n3167), .ZN(n5614)
         );
  OAI211_X1 U6660 ( .C1(n6005), .C2(n5616), .A(n5615), .B(n5614), .ZN(U2966)
         );
  AOI22_X1 U6661 ( .A1(n6054), .A2(REIP_REG_18__SCAN_IN), .B1(n6012), .B2(
        PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5625) );
  INV_X1 U6662 ( .A(n5617), .ZN(n5618) );
  NOR2_X1 U6663 ( .A1(n5626), .A2(n5618), .ZN(n5621) );
  INV_X1 U6664 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5695) );
  NOR2_X1 U6665 ( .A1(n5619), .A2(n5695), .ZN(n5620) );
  MUX2_X1 U6666 ( .A(n5621), .B(n5620), .S(n5452), .Z(n5623) );
  XNOR2_X1 U6667 ( .A(n5623), .B(n5622), .ZN(n5684) );
  AOI22_X1 U6668 ( .A1(n5684), .A2(n6010), .B1(n3167), .B2(n5748), .ZN(n5624)
         );
  OAI211_X1 U6669 ( .C1(n6005), .C2(n5743), .A(n5625), .B(n5624), .ZN(U2968)
         );
  MUX2_X1 U6670 ( .A(n5452), .B(n5627), .S(n5626), .Z(n5628) );
  AOI21_X1 U6671 ( .B1(INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n4388), .A(n5628), 
        .ZN(n5629) );
  XNOR2_X1 U6672 ( .A(n5629), .B(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5690)
         );
  AOI22_X1 U6673 ( .A1(n6054), .A2(REIP_REG_17__SCAN_IN), .B1(n6012), .B2(
        PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5631) );
  AOI22_X1 U6674 ( .A1(n5893), .A2(n3167), .B1(n5983), .B2(n5758), .ZN(n5630)
         );
  OAI211_X1 U6675 ( .C1(n5690), .C2(n5972), .A(n5631), .B(n5630), .ZN(U2969)
         );
  AND2_X1 U6676 ( .A1(n5633), .A2(n5632), .ZN(n5636) );
  OAI21_X1 U6677 ( .B1(n5636), .B2(n5635), .A(n5634), .ZN(n5709) );
  OAI22_X1 U6678 ( .A1(n5765), .A2(n6447), .B1(n5775), .B2(n6005), .ZN(n5637)
         );
  AOI21_X1 U6679 ( .B1(n6010), .B2(n5709), .A(n5637), .ZN(n5638) );
  NAND2_X1 U6680 ( .A1(n6054), .A2(REIP_REG_13__SCAN_IN), .ZN(n5715) );
  OAI211_X1 U6681 ( .C1(n3860), .C2(n5989), .A(n5638), .B(n5715), .ZN(U2973)
         );
  INV_X1 U6682 ( .A(n5639), .ZN(n5641) );
  AOI22_X1 U6683 ( .A1(n5641), .A2(n6060), .B1(n6041), .B2(n5640), .ZN(n5647)
         );
  INV_X1 U6684 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5643) );
  NOR2_X1 U6685 ( .A1(n6015), .A2(n6875), .ZN(n5642) );
  AOI221_X1 U6686 ( .B1(n5645), .B2(INSTADDRPOINTER_REG_27__SCAN_IN), .C1(
        n5644), .C2(n5643), .A(n5642), .ZN(n5646) );
  NAND2_X1 U6687 ( .A1(n5647), .A2(n5646), .ZN(U2991) );
  AOI22_X1 U6688 ( .A1(n6054), .A2(REIP_REG_25__SCAN_IN), .B1(n5648), .B2(
        n5427), .ZN(n5653) );
  INV_X1 U6689 ( .A(n5649), .ZN(n5650) );
  AOI22_X1 U6690 ( .A1(n5651), .A2(n6060), .B1(n6041), .B2(n5650), .ZN(n5652)
         );
  OAI211_X1 U6691 ( .C1(n5654), .C2(n5427), .A(n5653), .B(n5652), .ZN(U2993)
         );
  AOI22_X1 U6692 ( .A1(n6054), .A2(REIP_REG_21__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n5655), .ZN(n5660) );
  INV_X1 U6693 ( .A(n5656), .ZN(n5658) );
  AOI22_X1 U6694 ( .A1(n5658), .A2(n6060), .B1(n6041), .B2(n5657), .ZN(n5659)
         );
  OAI211_X1 U6695 ( .C1(INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n5661), .A(n5660), .B(n5659), .ZN(U2997) );
  AOI21_X1 U6696 ( .B1(n6048), .B2(n5663), .A(n5662), .ZN(n5696) );
  OAI21_X1 U6697 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n5689), .A(n5696), 
        .ZN(n5686) );
  AOI21_X1 U6698 ( .B1(n5622), .B2(n5664), .A(n5686), .ZN(n5681) );
  INV_X1 U6699 ( .A(n5674), .ZN(n5665) );
  NOR3_X1 U6700 ( .A1(n5667), .A2(n5666), .A3(n5665), .ZN(n5668) );
  AOI21_X1 U6701 ( .B1(REIP_REG_20__SCAN_IN), .B2(n6054), .A(n5668), .ZN(n5672) );
  AOI22_X1 U6702 ( .A1(n5670), .A2(n6060), .B1(n6041), .B2(n5669), .ZN(n5671)
         );
  OAI211_X1 U6703 ( .C1(n5681), .C2(n5673), .A(n5672), .B(n5671), .ZN(U2998)
         );
  AOI22_X1 U6704 ( .A1(n6054), .A2(REIP_REG_19__SCAN_IN), .B1(n5674), .B2(
        n5680), .ZN(n5679) );
  INV_X1 U6705 ( .A(n5675), .ZN(n5677) );
  AOI22_X1 U6706 ( .A1(n5677), .A2(n6060), .B1(n6041), .B2(n5676), .ZN(n5678)
         );
  OAI211_X1 U6707 ( .C1(n5681), .C2(n5680), .A(n5679), .B(n5678), .ZN(U2999)
         );
  NOR3_X1 U6708 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n5695), .A3(n5689), 
        .ZN(n5683) );
  NOR2_X1 U6709 ( .A1(n6015), .A2(n6854), .ZN(n5682) );
  AOI211_X1 U6710 ( .C1(n5684), .C2(n6060), .A(n5683), .B(n5682), .ZN(n5688)
         );
  INV_X1 U6711 ( .A(n5746), .ZN(n5685) );
  AOI22_X1 U6712 ( .A1(n5686), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .B1(n6041), .B2(n5685), .ZN(n5687) );
  NAND2_X1 U6713 ( .A1(n5688), .A2(n5687), .ZN(U3000) );
  NOR2_X1 U6714 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n5689), .ZN(n5692)
         );
  OAI22_X1 U6715 ( .A1(n5690), .A2(n6033), .B1(n6058), .B2(n5764), .ZN(n5691)
         );
  NOR2_X1 U6716 ( .A1(n5692), .A2(n5691), .ZN(n5694) );
  NAND2_X1 U6717 ( .A1(n6054), .A2(REIP_REG_17__SCAN_IN), .ZN(n5693) );
  OAI211_X1 U6718 ( .C1(n5696), .C2(n5695), .A(n5694), .B(n5693), .ZN(U3001)
         );
  NAND2_X1 U6719 ( .A1(n5698), .A2(n5697), .ZN(n5706) );
  INV_X1 U6720 ( .A(n5699), .ZN(n5701) );
  AOI21_X1 U6721 ( .B1(n5701), .B2(n6041), .A(n5700), .ZN(n5705) );
  AOI22_X1 U6722 ( .A1(n5703), .A2(n6060), .B1(INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n5702), .ZN(n5704) );
  OAI211_X1 U6723 ( .C1(INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n5706), .A(n5705), .B(n5704), .ZN(U3003) );
  OR2_X1 U6724 ( .A1(n5708), .A2(n5707), .ZN(n5717) );
  INV_X1 U6725 ( .A(n5709), .ZN(n5711) );
  OAI22_X1 U6726 ( .A1(n5711), .A2(n6033), .B1(n6058), .B2(n5710), .ZN(n5713)
         );
  AOI211_X1 U6727 ( .C1(n5714), .C2(INSTADDRPOINTER_REG_13__SCAN_IN), .A(n5713), .B(n5712), .ZN(n5716) );
  OAI211_X1 U6728 ( .C1(n5717), .C2(n6064), .A(n5716), .B(n5715), .ZN(U3005)
         );
  INV_X1 U6729 ( .A(n5718), .ZN(n5719) );
  NAND3_X1 U6730 ( .A1(n5720), .A2(n6615), .A3(n5719), .ZN(n5721) );
  OAI21_X1 U6731 ( .B1(n6629), .B2(n5722), .A(n5721), .ZN(U3455) );
  INV_X1 U6732 ( .A(STATE_REG_0__SCAN_IN), .ZN(n6785) );
  NAND2_X1 U6733 ( .A1(n6785), .A2(STATE_REG_1__SCAN_IN), .ZN(n7047) );
  INV_X1 U6734 ( .A(ADS_N_REG_SCAN_IN), .ZN(n7004) );
  INV_X1 U6735 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6576) );
  OAI21_X1 U6736 ( .B1(n7048), .B2(n7004), .A(n6608), .ZN(U2789) );
  OAI21_X1 U6737 ( .B1(n5723), .B2(n6550), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n5724) );
  OAI21_X1 U6738 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6551), .A(n5724), .ZN(
        U2790) );
  INV_X1 U6739 ( .A(D_C_N_REG_SCAN_IN), .ZN(n7018) );
  NOR2_X1 U6740 ( .A1(STATE_REG_0__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n5726) );
  NOR2_X1 U6741 ( .A1(n7048), .A2(n5726), .ZN(n5725) );
  AOI22_X1 U6742 ( .A1(CODEFETCH_REG_SCAN_IN), .A2(n7048), .B1(n7018), .B2(
        n5725), .ZN(U2791) );
  INV_X1 U6743 ( .A(n6608), .ZN(n6611) );
  OAI21_X1 U6744 ( .B1(BS16_N), .B2(n5726), .A(n6611), .ZN(n6609) );
  OAI21_X1 U6745 ( .B1(n6611), .B2(n6852), .A(n6609), .ZN(U2792) );
  INV_X1 U6746 ( .A(n5727), .ZN(n5729) );
  OAI21_X1 U6747 ( .B1(n5729), .B2(n5728), .A(n5972), .ZN(U2793) );
  NOR4_X1 U6748 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(
        DATAWIDTH_REG_20__SCAN_IN), .A3(DATAWIDTH_REG_6__SCAN_IN), .A4(
        DATAWIDTH_REG_21__SCAN_IN), .ZN(n5733) );
  NOR4_X1 U6749 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(DATAWIDTH_REG_18__SCAN_IN), .A3(DATAWIDTH_REG_8__SCAN_IN), .A4(DATAWIDTH_REG_15__SCAN_IN), .ZN(n5732) );
  NOR4_X1 U6750 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(
        DATAWIDTH_REG_29__SCAN_IN), .A3(DATAWIDTH_REG_30__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n5731) );
  NOR4_X1 U6751 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(
        DATAWIDTH_REG_25__SCAN_IN), .A3(DATAWIDTH_REG_26__SCAN_IN), .A4(
        DATAWIDTH_REG_27__SCAN_IN), .ZN(n5730) );
  NAND4_X1 U6752 ( .A1(n5733), .A2(n5732), .A3(n5731), .A4(n5730), .ZN(n5739)
         );
  NOR4_X1 U6753 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(DATAWIDTH_REG_5__SCAN_IN), 
        .A3(DATAWIDTH_REG_3__SCAN_IN), .A4(DATAWIDTH_REG_14__SCAN_IN), .ZN(
        n5737) );
  AOI211_X1 U6754 ( .C1(DATAWIDTH_REG_0__SCAN_IN), .C2(
        DATAWIDTH_REG_1__SCAN_IN), .A(DATAWIDTH_REG_19__SCAN_IN), .B(
        DATAWIDTH_REG_17__SCAN_IN), .ZN(n5736) );
  NOR4_X1 U6755 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(
        DATAWIDTH_REG_23__SCAN_IN), .A3(DATAWIDTH_REG_10__SCAN_IN), .A4(
        DATAWIDTH_REG_11__SCAN_IN), .ZN(n5735) );
  NOR4_X1 U6756 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(DATAWIDTH_REG_16__SCAN_IN), .A3(DATAWIDTH_REG_7__SCAN_IN), .A4(DATAWIDTH_REG_13__SCAN_IN), .ZN(n5734) );
  NAND4_X1 U6757 ( .A1(n5737), .A2(n5736), .A3(n5735), .A4(n5734), .ZN(n5738)
         );
  NOR2_X1 U6758 ( .A1(n5739), .A2(n5738), .ZN(n6641) );
  INV_X1 U6759 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n6992) );
  NOR3_X1 U6760 ( .A1(REIP_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_0__SCAN_IN), 
        .A3(DATAWIDTH_REG_1__SCAN_IN), .ZN(n5741) );
  OAI21_X1 U6761 ( .B1(REIP_REG_1__SCAN_IN), .B2(n5741), .A(n6641), .ZN(n5740)
         );
  OAI21_X1 U6762 ( .B1(n6641), .B2(n6992), .A(n5740), .ZN(U2794) );
  INV_X1 U6763 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n6987) );
  NOR2_X1 U6764 ( .A1(REIP_REG_1__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .ZN(n6637) );
  OAI21_X1 U6765 ( .B1(n5741), .B2(n6637), .A(n6641), .ZN(n5742) );
  OAI21_X1 U6766 ( .B1(n6641), .B2(n6987), .A(n5742), .ZN(U2795) );
  INV_X1 U6767 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5744) );
  OAI22_X1 U6768 ( .A1(n5744), .A2(n5886), .B1(n5743), .B2(n5885), .ZN(n5745)
         );
  AOI211_X1 U6769 ( .C1(n5879), .C2(EBX_REG_18__SCAN_IN), .A(n5848), .B(n5745), 
        .ZN(n5754) );
  NOR2_X1 U6770 ( .A1(n5746), .A2(n5881), .ZN(n5747) );
  AOI21_X1 U6771 ( .B1(n5748), .B2(n5804), .A(n5747), .ZN(n5753) );
  INV_X1 U6772 ( .A(n5749), .ZN(n5751) );
  OAI21_X1 U6773 ( .B1(n5751), .B2(REIP_REG_18__SCAN_IN), .A(n5750), .ZN(n5752) );
  NAND3_X1 U6774 ( .A1(n5754), .A2(n5753), .A3(n5752), .ZN(U2809) );
  AOI21_X1 U6775 ( .B1(n5755), .B2(REIP_REG_16__SCAN_IN), .A(
        REIP_REG_17__SCAN_IN), .ZN(n5756) );
  NOR3_X1 U6776 ( .A1(n5876), .A2(n5757), .A3(n5756), .ZN(n5762) );
  AOI22_X1 U6777 ( .A1(EBX_REG_17__SCAN_IN), .A2(n5879), .B1(n5758), .B2(n5802), .ZN(n5759) );
  OAI211_X1 U6778 ( .C1(n5886), .C2(n5760), .A(n5759), .B(n5825), .ZN(n5761)
         );
  AOI211_X1 U6779 ( .C1(n5893), .C2(n5804), .A(n5762), .B(n5761), .ZN(n5763)
         );
  OAI21_X1 U6780 ( .B1(n5881), .B2(n5764), .A(n5763), .ZN(U2810) );
  INV_X1 U6781 ( .A(n5765), .ZN(n5771) );
  INV_X1 U6782 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6592) );
  NOR3_X1 U6783 ( .A1(REIP_REG_13__SCAN_IN), .A2(n5766), .A3(n6592), .ZN(n5770) );
  AOI22_X1 U6784 ( .A1(EBX_REG_13__SCAN_IN), .A2(n5879), .B1(n5866), .B2(n5767), .ZN(n5768) );
  OAI211_X1 U6785 ( .C1(n5886), .C2(n3860), .A(n5768), .B(n5825), .ZN(n5769)
         );
  AOI211_X1 U6786 ( .C1(n5771), .C2(n5804), .A(n5770), .B(n5769), .ZN(n5774)
         );
  OAI21_X1 U6787 ( .B1(n5777), .B2(n5772), .A(REIP_REG_13__SCAN_IN), .ZN(n5773) );
  OAI211_X1 U6788 ( .C1(n5885), .C2(n5775), .A(n5774), .B(n5773), .ZN(U2814)
         );
  AOI21_X1 U6789 ( .B1(n5776), .B2(REIP_REG_10__SCAN_IN), .A(
        REIP_REG_11__SCAN_IN), .ZN(n5784) );
  INV_X1 U6790 ( .A(n5777), .ZN(n5783) );
  OAI22_X1 U6791 ( .A1(n5779), .A2(n5886), .B1(n5881), .B2(n5778), .ZN(n5780)
         );
  AOI211_X1 U6792 ( .C1(n5879), .C2(EBX_REG_11__SCAN_IN), .A(n5848), .B(n5780), 
        .ZN(n5782) );
  AOI22_X1 U6793 ( .A1(n5969), .A2(n5804), .B1(n5802), .B2(n5968), .ZN(n5781)
         );
  OAI211_X1 U6794 ( .C1(n5784), .C2(n5783), .A(n5782), .B(n5781), .ZN(U2816)
         );
  OAI21_X1 U6795 ( .B1(n5796), .B2(n5851), .A(n5820), .ZN(n5800) );
  AOI22_X1 U6796 ( .A1(EBX_REG_9__SCAN_IN), .A2(n5879), .B1(
        REIP_REG_9__SCAN_IN), .B2(n5800), .ZN(n5794) );
  NOR2_X1 U6797 ( .A1(n5785), .A2(n5881), .ZN(n5788) );
  OAI21_X1 U6798 ( .B1(n5886), .B2(n5786), .A(n5825), .ZN(n5787) );
  AOI211_X1 U6799 ( .C1(n5789), .C2(n5804), .A(n5788), .B(n5787), .ZN(n5793)
         );
  INV_X1 U6800 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6587) );
  NAND3_X1 U6801 ( .A1(n5845), .A2(n5796), .A3(n6587), .ZN(n5792) );
  NAND2_X1 U6802 ( .A1(n5790), .A2(n5802), .ZN(n5791) );
  NAND4_X1 U6803 ( .A1(n5794), .A2(n5793), .A3(n5792), .A4(n5791), .ZN(U2818)
         );
  INV_X1 U6804 ( .A(n5795), .ZN(n5798) );
  NOR2_X1 U6805 ( .A1(n5796), .A2(n5851), .ZN(n5797) );
  AOI22_X1 U6806 ( .A1(n5866), .A2(n5799), .B1(n5798), .B2(n5797), .ZN(n5809)
         );
  AOI22_X1 U6807 ( .A1(EBX_REG_8__SCAN_IN), .A2(n5879), .B1(
        PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n5849), .ZN(n5808) );
  AOI21_X1 U6808 ( .B1(REIP_REG_8__SCAN_IN), .B2(n5800), .A(n5848), .ZN(n5807)
         );
  INV_X1 U6809 ( .A(n5801), .ZN(n5803) );
  AOI22_X1 U6810 ( .A1(n5805), .A2(n5804), .B1(n5803), .B2(n5802), .ZN(n5806)
         );
  NAND4_X1 U6811 ( .A1(n5809), .A2(n5808), .A3(n5807), .A4(n5806), .ZN(U2819)
         );
  INV_X1 U6812 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6584) );
  NAND3_X1 U6813 ( .A1(n5845), .A2(n5810), .A3(n6584), .ZN(n5817) );
  INV_X1 U6814 ( .A(n5811), .ZN(n5815) );
  NAND2_X1 U6815 ( .A1(n5849), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n5812)
         );
  OAI211_X1 U6816 ( .C1(n5862), .C2(n5813), .A(n5812), .B(n5825), .ZN(n5814)
         );
  AOI21_X1 U6817 ( .B1(n5815), .B2(n5866), .A(n5814), .ZN(n5816) );
  OAI211_X1 U6818 ( .C1(n5975), .C2(n5830), .A(n5817), .B(n5816), .ZN(n5818)
         );
  INV_X1 U6819 ( .A(n5818), .ZN(n5824) );
  INV_X1 U6820 ( .A(n5819), .ZN(n5821) );
  OAI21_X1 U6821 ( .B1(n5851), .B2(n5821), .A(n5820), .ZN(n5840) );
  INV_X1 U6822 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6582) );
  NAND2_X1 U6823 ( .A1(n5845), .A2(n5822), .ZN(n5839) );
  NOR3_X1 U6824 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6582), .A3(n5839), .ZN(n5833)
         );
  OAI21_X1 U6825 ( .B1(n5840), .B2(n5833), .A(REIP_REG_7__SCAN_IN), .ZN(n5823)
         );
  OAI211_X1 U6826 ( .C1(n5885), .C2(n5974), .A(n5824), .B(n5823), .ZN(U2820)
         );
  INV_X1 U6827 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n5827) );
  NAND2_X1 U6828 ( .A1(n5879), .A2(EBX_REG_6__SCAN_IN), .ZN(n5826) );
  OAI211_X1 U6829 ( .C1(n5886), .C2(n5827), .A(n5826), .B(n5825), .ZN(n5828)
         );
  AOI21_X1 U6830 ( .B1(REIP_REG_6__SCAN_IN), .B2(n5840), .A(n5828), .ZN(n5829)
         );
  OAI21_X1 U6831 ( .B1(n5831), .B2(n5830), .A(n5829), .ZN(n5832) );
  AOI211_X1 U6832 ( .C1(n5834), .C2(n5866), .A(n5833), .B(n5832), .ZN(n5835)
         );
  OAI21_X1 U6833 ( .B1(n5836), .B2(n5885), .A(n5835), .ZN(U2821) );
  OAI22_X1 U6834 ( .A1(n5990), .A2(n5886), .B1(n5881), .B2(n5837), .ZN(n5838)
         );
  AOI211_X1 U6835 ( .C1(n5879), .C2(EBX_REG_5__SCAN_IN), .A(n5848), .B(n5838), 
        .ZN(n5843) );
  NAND2_X1 U6836 ( .A1(n6582), .A2(n5839), .ZN(n5841) );
  AOI22_X1 U6837 ( .A1(n5841), .A2(n5840), .B1(n5985), .B2(n5883), .ZN(n5842)
         );
  OAI211_X1 U6838 ( .C1(n5982), .C2(n5885), .A(n5843), .B(n5842), .ZN(U2822)
         );
  AOI21_X1 U6839 ( .B1(n5845), .B2(n5850), .A(n5844), .ZN(n5870) );
  OAI22_X1 U6840 ( .A1(n6581), .A2(n5870), .B1(n5846), .B2(n5877), .ZN(n5847)
         );
  AOI211_X1 U6841 ( .C1(n5849), .C2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n5848), 
        .B(n5847), .ZN(n5858) );
  INV_X1 U6842 ( .A(EBX_REG_4__SCAN_IN), .ZN(n5854) );
  NAND2_X1 U6843 ( .A1(n5866), .A2(n6030), .ZN(n5853) );
  OR3_X1 U6844 ( .A1(n5851), .A2(REIP_REG_4__SCAN_IN), .A3(n5850), .ZN(n5852)
         );
  OAI211_X1 U6845 ( .C1(n5854), .C2(n5862), .A(n5853), .B(n5852), .ZN(n5855)
         );
  AOI21_X1 U6846 ( .B1(n5856), .B2(n5883), .A(n5855), .ZN(n5857) );
  OAI211_X1 U6847 ( .C1(n5859), .C2(n5885), .A(n5858), .B(n5857), .ZN(U2823)
         );
  INV_X1 U6848 ( .A(n5860), .ZN(n5875) );
  OAI22_X1 U6849 ( .A1(n5886), .A2(n5863), .B1(n5862), .B2(n5861), .ZN(n5864)
         );
  AOI21_X1 U6850 ( .B1(n5866), .B2(n5865), .A(n5864), .ZN(n5867) );
  OAI21_X1 U6851 ( .B1(n6399), .B2(n5877), .A(n5867), .ZN(n5868) );
  AOI21_X1 U6852 ( .B1(n5869), .B2(n5883), .A(n5868), .ZN(n5874) );
  INV_X1 U6853 ( .A(n5870), .ZN(n5871) );
  OAI21_X1 U6854 ( .B1(REIP_REG_3__SCAN_IN), .B2(n5872), .A(n5871), .ZN(n5873)
         );
  OAI211_X1 U6855 ( .C1(n5885), .C2(n5875), .A(n5874), .B(n5873), .ZN(U2824)
         );
  INV_X1 U6856 ( .A(REIP_REG_0__SCAN_IN), .ZN(n6016) );
  OAI22_X1 U6857 ( .A1(n5877), .A2(n6624), .B1(n5876), .B2(n6016), .ZN(n5878)
         );
  AOI21_X1 U6858 ( .B1(n5879), .B2(EBX_REG_0__SCAN_IN), .A(n5878), .ZN(n5880)
         );
  OAI21_X1 U6859 ( .B1(n5881), .B2(n6057), .A(n5880), .ZN(n5882) );
  AOI21_X1 U6860 ( .B1(n6009), .B2(n5883), .A(n5882), .ZN(n5884) );
  OAI221_X1 U6861 ( .B1(n5887), .B2(n5886), .C1(n5887), .C2(n5885), .A(n5884), 
        .ZN(U2827) );
  AOI22_X1 U6862 ( .A1(n5995), .A2(n5889), .B1(n5888), .B2(n6040), .ZN(n5890)
         );
  OAI21_X1 U6863 ( .B1(n5892), .B2(n5891), .A(n5890), .ZN(U2857) );
  AOI22_X1 U6864 ( .A1(n5893), .A2(n5898), .B1(n5897), .B2(DATAI_17_), .ZN(
        n5895) );
  AOI22_X1 U6865 ( .A1(n5901), .A2(DATAI_1_), .B1(n5900), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n5894) );
  NAND2_X1 U6866 ( .A1(n5895), .A2(n5894), .ZN(U2874) );
  INV_X1 U6867 ( .A(n5896), .ZN(n5899) );
  AOI22_X1 U6868 ( .A1(n5899), .A2(n5898), .B1(n5897), .B2(DATAI_16_), .ZN(
        n5903) );
  AOI22_X1 U6869 ( .A1(n5901), .A2(DATAI_0_), .B1(n5900), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n5902) );
  NAND2_X1 U6870 ( .A1(n5903), .A2(n5902), .ZN(U2875) );
  OAI222_X1 U6871 ( .A1(n5906), .A2(n5413), .B1(n5905), .B2(n5967), .C1(n5904), 
        .C2(n7023), .ZN(U2891) );
  INV_X1 U6872 ( .A(EAX_REG_30__SCAN_IN), .ZN(n5909) );
  NAND2_X1 U6873 ( .A1(n5937), .A2(n5907), .ZN(n5935) );
  AOI22_X1 U6874 ( .A1(n6536), .A2(UWORD_REG_14__SCAN_IN), .B1(n5964), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n5908) );
  OAI21_X1 U6875 ( .B1(n5909), .B2(n5935), .A(n5908), .ZN(U2893) );
  INV_X1 U6876 ( .A(EAX_REG_29__SCAN_IN), .ZN(n5911) );
  AOI22_X1 U6877 ( .A1(n6536), .A2(UWORD_REG_13__SCAN_IN), .B1(n5964), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n5910) );
  OAI21_X1 U6878 ( .B1(n5911), .B2(n5935), .A(n5910), .ZN(U2894) );
  INV_X1 U6879 ( .A(EAX_REG_28__SCAN_IN), .ZN(n5913) );
  AOI22_X1 U6880 ( .A1(n6536), .A2(UWORD_REG_12__SCAN_IN), .B1(n5952), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n5912) );
  OAI21_X1 U6881 ( .B1(n5913), .B2(n5935), .A(n5912), .ZN(U2895) );
  INV_X1 U6882 ( .A(EAX_REG_27__SCAN_IN), .ZN(n5915) );
  AOI22_X1 U6883 ( .A1(n6536), .A2(UWORD_REG_11__SCAN_IN), .B1(n5952), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n5914) );
  OAI21_X1 U6884 ( .B1(n5915), .B2(n5935), .A(n5914), .ZN(U2896) );
  INV_X1 U6885 ( .A(EAX_REG_26__SCAN_IN), .ZN(n5917) );
  AOI22_X1 U6886 ( .A1(n6536), .A2(UWORD_REG_10__SCAN_IN), .B1(n5952), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n5916) );
  OAI21_X1 U6887 ( .B1(n5917), .B2(n5935), .A(n5916), .ZN(U2897) );
  INV_X1 U6888 ( .A(EAX_REG_25__SCAN_IN), .ZN(n5919) );
  AOI22_X1 U6889 ( .A1(n6536), .A2(UWORD_REG_9__SCAN_IN), .B1(n5952), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n5918) );
  OAI21_X1 U6890 ( .B1(n5919), .B2(n5935), .A(n5918), .ZN(U2898) );
  AOI22_X1 U6891 ( .A1(n6536), .A2(UWORD_REG_8__SCAN_IN), .B1(n5952), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n5920) );
  OAI21_X1 U6892 ( .B1(n4048), .B2(n5935), .A(n5920), .ZN(U2899) );
  INV_X1 U6893 ( .A(EAX_REG_23__SCAN_IN), .ZN(n5922) );
  AOI22_X1 U6894 ( .A1(n6536), .A2(UWORD_REG_7__SCAN_IN), .B1(n5964), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n5921) );
  OAI21_X1 U6895 ( .B1(n5922), .B2(n5935), .A(n5921), .ZN(U2900) );
  INV_X1 U6896 ( .A(EAX_REG_22__SCAN_IN), .ZN(n5924) );
  AOI22_X1 U6897 ( .A1(n6536), .A2(UWORD_REG_6__SCAN_IN), .B1(n5964), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n5923) );
  OAI21_X1 U6898 ( .B1(n5924), .B2(n5935), .A(n5923), .ZN(U2901) );
  INV_X1 U6899 ( .A(EAX_REG_21__SCAN_IN), .ZN(n5926) );
  AOI22_X1 U6900 ( .A1(n6536), .A2(UWORD_REG_5__SCAN_IN), .B1(n5964), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n5925) );
  OAI21_X1 U6901 ( .B1(n5926), .B2(n5935), .A(n5925), .ZN(U2902) );
  AOI22_X1 U6902 ( .A1(n6536), .A2(UWORD_REG_4__SCAN_IN), .B1(n5964), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n5927) );
  OAI21_X1 U6903 ( .B1(n3989), .B2(n5935), .A(n5927), .ZN(U2903) );
  INV_X1 U6904 ( .A(EAX_REG_19__SCAN_IN), .ZN(n5929) );
  AOI22_X1 U6905 ( .A1(n6536), .A2(UWORD_REG_3__SCAN_IN), .B1(n5964), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n5928) );
  OAI21_X1 U6906 ( .B1(n5929), .B2(n5935), .A(n5928), .ZN(U2904) );
  INV_X1 U6907 ( .A(EAX_REG_18__SCAN_IN), .ZN(n5931) );
  AOI22_X1 U6908 ( .A1(n6536), .A2(UWORD_REG_2__SCAN_IN), .B1(n5964), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n5930) );
  OAI21_X1 U6909 ( .B1(n5931), .B2(n5935), .A(n5930), .ZN(U2905) );
  INV_X1 U6910 ( .A(EAX_REG_17__SCAN_IN), .ZN(n5933) );
  AOI22_X1 U6911 ( .A1(n6536), .A2(UWORD_REG_1__SCAN_IN), .B1(n5964), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n5932) );
  OAI21_X1 U6912 ( .B1(n5933), .B2(n5935), .A(n5932), .ZN(U2906) );
  INV_X1 U6913 ( .A(EAX_REG_16__SCAN_IN), .ZN(n5936) );
  AOI22_X1 U6914 ( .A1(n6536), .A2(UWORD_REG_0__SCAN_IN), .B1(n5964), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n5934) );
  OAI21_X1 U6915 ( .B1(n5936), .B2(n5935), .A(n5934), .ZN(U2907) );
  INV_X1 U6916 ( .A(n5937), .ZN(n5966) );
  AOI22_X1 U6917 ( .A1(n6536), .A2(LWORD_REG_15__SCAN_IN), .B1(n5964), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n5938) );
  OAI21_X1 U6918 ( .B1(n4498), .B2(n5966), .A(n5938), .ZN(U2908) );
  AOI22_X1 U6919 ( .A1(n6536), .A2(LWORD_REG_14__SCAN_IN), .B1(n5964), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n5939) );
  OAI21_X1 U6920 ( .B1(n5137), .B2(n5966), .A(n5939), .ZN(U2909) );
  INV_X1 U6921 ( .A(EAX_REG_13__SCAN_IN), .ZN(n5941) );
  AOI22_X1 U6922 ( .A1(n6536), .A2(LWORD_REG_13__SCAN_IN), .B1(n5964), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n5940) );
  OAI21_X1 U6923 ( .B1(n5941), .B2(n5966), .A(n5940), .ZN(U2910) );
  AOI22_X1 U6924 ( .A1(n6536), .A2(LWORD_REG_12__SCAN_IN), .B1(n5964), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n5942) );
  OAI21_X1 U6925 ( .B1(n5041), .B2(n5966), .A(n5942), .ZN(U2911) );
  AOI22_X1 U6926 ( .A1(n6536), .A2(LWORD_REG_11__SCAN_IN), .B1(n5964), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n5943) );
  OAI21_X1 U6927 ( .B1(n4981), .B2(n5966), .A(n5943), .ZN(U2912) );
  INV_X1 U6928 ( .A(EAX_REG_10__SCAN_IN), .ZN(n5945) );
  AOI22_X1 U6929 ( .A1(n6536), .A2(LWORD_REG_10__SCAN_IN), .B1(n5952), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n5944) );
  OAI21_X1 U6930 ( .B1(n5945), .B2(n5966), .A(n5944), .ZN(U2913) );
  INV_X1 U6931 ( .A(EAX_REG_9__SCAN_IN), .ZN(n5947) );
  AOI22_X1 U6932 ( .A1(n6536), .A2(LWORD_REG_9__SCAN_IN), .B1(n5952), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n5946) );
  OAI21_X1 U6933 ( .B1(n5947), .B2(n5966), .A(n5946), .ZN(U2914) );
  INV_X1 U6934 ( .A(EAX_REG_8__SCAN_IN), .ZN(n5949) );
  AOI22_X1 U6935 ( .A1(n6536), .A2(LWORD_REG_8__SCAN_IN), .B1(n5952), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n5948) );
  OAI21_X1 U6936 ( .B1(n5949), .B2(n5966), .A(n5948), .ZN(U2915) );
  AOI22_X1 U6937 ( .A1(n6536), .A2(LWORD_REG_7__SCAN_IN), .B1(n5952), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n5950) );
  OAI21_X1 U6938 ( .B1(n5951), .B2(n5966), .A(n5950), .ZN(U2916) );
  AOI22_X1 U6939 ( .A1(n6536), .A2(LWORD_REG_6__SCAN_IN), .B1(n5952), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n5953) );
  OAI21_X1 U6940 ( .B1(n3818), .B2(n5966), .A(n5953), .ZN(U2917) );
  AOI22_X1 U6941 ( .A1(n6536), .A2(LWORD_REG_5__SCAN_IN), .B1(n5964), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n5954) );
  OAI21_X1 U6942 ( .B1(n5955), .B2(n5966), .A(n5954), .ZN(U2918) );
  AOI22_X1 U6943 ( .A1(n6536), .A2(LWORD_REG_4__SCAN_IN), .B1(n5964), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n5956) );
  OAI21_X1 U6944 ( .B1(n5957), .B2(n5966), .A(n5956), .ZN(U2919) );
  AOI22_X1 U6945 ( .A1(n6536), .A2(LWORD_REG_3__SCAN_IN), .B1(n5964), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n5958) );
  OAI21_X1 U6946 ( .B1(n5959), .B2(n5966), .A(n5958), .ZN(U2920) );
  AOI22_X1 U6947 ( .A1(n6536), .A2(LWORD_REG_2__SCAN_IN), .B1(n5964), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n5960) );
  OAI21_X1 U6948 ( .B1(n5961), .B2(n5966), .A(n5960), .ZN(U2921) );
  AOI22_X1 U6949 ( .A1(n6536), .A2(LWORD_REG_1__SCAN_IN), .B1(n5964), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n5962) );
  OAI21_X1 U6950 ( .B1(n5963), .B2(n5966), .A(n5962), .ZN(U2922) );
  AOI22_X1 U6951 ( .A1(n6536), .A2(LWORD_REG_0__SCAN_IN), .B1(n5964), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n5965) );
  OAI21_X1 U6952 ( .B1(n5967), .B2(n5966), .A(n5965), .ZN(U2923) );
  AOI22_X1 U6953 ( .A1(n6054), .A2(REIP_REG_11__SCAN_IN), .B1(n6012), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n5971) );
  AOI22_X1 U6954 ( .A1(n5969), .A2(n3167), .B1(n5983), .B2(n5968), .ZN(n5970)
         );
  OAI211_X1 U6955 ( .C1(n5973), .C2(n5972), .A(n5971), .B(n5970), .ZN(U2975)
         );
  OAI22_X1 U6956 ( .A1(n5975), .A2(n6447), .B1(n5974), .B2(n6005), .ZN(n5976)
         );
  AOI21_X1 U6957 ( .B1(n5977), .B2(n6010), .A(n5976), .ZN(n5979) );
  OAI211_X1 U6958 ( .C1(n5980), .C2(n5989), .A(n5979), .B(n5978), .ZN(U2979)
         );
  INV_X1 U6959 ( .A(n5981), .ZN(n5986) );
  INV_X1 U6960 ( .A(n5982), .ZN(n5984) );
  AOI222_X1 U6961 ( .A1(n5986), .A2(n6010), .B1(n5985), .B2(n3167), .C1(n5984), 
        .C2(n5983), .ZN(n5988) );
  OAI211_X1 U6962 ( .C1(n5990), .C2(n5989), .A(n5988), .B(n5987), .ZN(U2981)
         );
  AOI22_X1 U6963 ( .A1(n6054), .A2(REIP_REG_2__SCAN_IN), .B1(n6012), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n5997) );
  NAND2_X1 U6964 ( .A1(n5992), .A2(n5991), .ZN(n5993) );
  XOR2_X1 U6965 ( .A(n5994), .B(n5993), .Z(n6046) );
  AOI22_X1 U6966 ( .A1(n6046), .A2(n6010), .B1(n3167), .B2(n5995), .ZN(n5996)
         );
  OAI211_X1 U6967 ( .C1(n6005), .C2(n5998), .A(n5997), .B(n5996), .ZN(U2984)
         );
  AOI22_X1 U6968 ( .A1(n6054), .A2(REIP_REG_1__SCAN_IN), .B1(n6012), .B2(
        PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n6004) );
  INV_X1 U6969 ( .A(n5999), .ZN(n6002) );
  INV_X1 U6970 ( .A(n6000), .ZN(n6001) );
  AOI22_X1 U6971 ( .A1(n6010), .A2(n6002), .B1(n6001), .B2(n3167), .ZN(n6003)
         );
  OAI211_X1 U6972 ( .C1(PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n6005), .A(n6004), 
        .B(n6003), .ZN(U2985) );
  INV_X1 U6973 ( .A(n6006), .ZN(n6008) );
  AOI21_X1 U6974 ( .B1(n6008), .B2(n6065), .A(n6007), .ZN(n6061) );
  AOI22_X1 U6975 ( .A1(n6010), .A2(n6061), .B1(n3167), .B2(n6009), .ZN(n6014)
         );
  OAI21_X1 U6976 ( .B1(n6012), .B2(n6011), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n6013) );
  OAI211_X1 U6977 ( .C1(n6016), .C2(n6015), .A(n6014), .B(n6013), .ZN(U2986)
         );
  AOI22_X1 U6978 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n6018), .B1(
        INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n6017), .ZN(n6025) );
  AOI21_X1 U6979 ( .B1(n6020), .B2(n6041), .A(n6019), .ZN(n6024) );
  AOI22_X1 U6980 ( .A1(n6022), .A2(n6060), .B1(INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n6021), .ZN(n6023) );
  OAI211_X1 U6981 ( .C1(n6026), .C2(n6025), .A(n6024), .B(n6023), .ZN(U3008)
         );
  OR2_X1 U6982 ( .A1(n6028), .A2(n6027), .ZN(n6032) );
  AOI21_X1 U6983 ( .B1(n6041), .B2(n6030), .A(n6029), .ZN(n6031) );
  OAI211_X1 U6984 ( .C1(n6034), .C2(n6033), .A(n6032), .B(n6031), .ZN(n6035)
         );
  INV_X1 U6985 ( .A(n6035), .ZN(n6039) );
  OAI211_X1 U6986 ( .C1(INSTADDRPOINTER_REG_3__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A(n6037), .B(n6036), .ZN(n6038) );
  NAND2_X1 U6987 ( .A1(n6039), .A2(n6038), .ZN(U3014) );
  AOI22_X1 U6988 ( .A1(n6041), .A2(n6040), .B1(n6054), .B2(REIP_REG_2__SCAN_IN), .ZN(n6053) );
  NAND3_X1 U6989 ( .A1(n6048), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6044) );
  INV_X1 U6990 ( .A(n6042), .ZN(n6043) );
  NAND2_X1 U6991 ( .A1(n6044), .A2(n6043), .ZN(n6045) );
  AOI22_X1 U6992 ( .A1(n6046), .A2(n6060), .B1(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .B2(n6045), .ZN(n6052) );
  NAND2_X1 U6993 ( .A1(n6048), .A2(n6047), .ZN(n6051) );
  NAND3_X1 U6994 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n3528), .A3(n6049), 
        .ZN(n6050) );
  NAND4_X1 U6995 ( .A1(n6053), .A2(n6052), .A3(n6051), .A4(n6050), .ZN(U3016)
         );
  NAND2_X1 U6996 ( .A1(n6054), .A2(REIP_REG_0__SCAN_IN), .ZN(n6055) );
  OAI211_X1 U6997 ( .C1(n6058), .C2(n6057), .A(n6056), .B(n6055), .ZN(n6059)
         );
  AOI21_X1 U6998 ( .B1(n6061), .B2(n6060), .A(n6059), .ZN(n6062) );
  OAI221_X1 U6999 ( .B1(n6065), .B2(n6064), .C1(n6065), .C2(n6063), .A(n6062), 
        .ZN(U3018) );
  INV_X1 U7000 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6067) );
  NOR2_X1 U7001 ( .A1(n6067), .A2(n6066), .ZN(U3019) );
  INV_X1 U7002 ( .A(n4666), .ZN(n6221) );
  NAND2_X1 U7003 ( .A1(n6221), .A2(n6068), .ZN(n6069) );
  OR2_X1 U7004 ( .A1(n6070), .A2(n6069), .ZN(n6102) );
  NAND2_X1 U7005 ( .A1(n4533), .A2(n6071), .ZN(n6258) );
  NOR2_X1 U7006 ( .A1(n6257), .A2(n6258), .ZN(n6103) );
  INV_X1 U7007 ( .A(n6103), .ZN(n6074) );
  INV_X1 U7008 ( .A(n6072), .ZN(n6073) );
  INV_X1 U7009 ( .A(n6402), .ZN(n6335) );
  OAI22_X1 U7010 ( .A1(n6074), .A2(n6643), .B1(n6073), .B2(n6335), .ZN(n6096)
         );
  NAND3_X1 U7011 ( .A1(n6403), .A2(n6521), .A3(n6517), .ZN(n6106) );
  NOR2_X1 U7012 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6106), .ZN(n6097)
         );
  AOI22_X1 U7013 ( .A1(n6445), .A2(n6096), .B1(n6446), .B2(n6097), .ZN(n6083)
         );
  INV_X1 U7014 ( .A(n6075), .ZN(n6448) );
  NAND2_X1 U7015 ( .A1(n6448), .A2(n6076), .ZN(n6484) );
  NOR3_X1 U7016 ( .A1(n6119), .A2(n6502), .A3(n6643), .ZN(n6077) );
  NOR2_X1 U7017 ( .A1(n6077), .A2(n6449), .ZN(n6081) );
  INV_X1 U7018 ( .A(n6097), .ZN(n6079) );
  AOI211_X1 U7019 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6079), .A(n6226), .B(
        n6078), .ZN(n6080) );
  OAI21_X1 U7020 ( .B1(n6081), .B2(n6103), .A(n6080), .ZN(n6098) );
  AOI22_X1 U7021 ( .A1(INSTQUEUE_REG_0__0__SCAN_IN), .A2(n6098), .B1(n6412), 
        .B2(n6502), .ZN(n6082) );
  OAI211_X1 U7022 ( .C1(n6415), .C2(n6129), .A(n6083), .B(n6082), .ZN(U3020)
         );
  AOI22_X1 U7023 ( .A1(n6461), .A2(n6097), .B1(n6460), .B2(n6096), .ZN(n6085)
         );
  AOI22_X1 U7024 ( .A1(INSTQUEUE_REG_0__1__SCAN_IN), .A2(n6098), .B1(n6462), 
        .B2(n6502), .ZN(n6084) );
  OAI211_X1 U7025 ( .C1(n6465), .C2(n6129), .A(n6085), .B(n6084), .ZN(U3021)
         );
  AOI22_X1 U7026 ( .A1(n6467), .A2(n6097), .B1(n6466), .B2(n6096), .ZN(n6087)
         );
  AOI22_X1 U7027 ( .A1(INSTQUEUE_REG_0__2__SCAN_IN), .A2(n6098), .B1(n6468), 
        .B2(n6502), .ZN(n6086) );
  OAI211_X1 U7028 ( .C1(n6471), .C2(n6129), .A(n6087), .B(n6086), .ZN(U3022)
         );
  AOI22_X1 U7029 ( .A1(n6473), .A2(n6097), .B1(n6472), .B2(n6096), .ZN(n6089)
         );
  AOI22_X1 U7030 ( .A1(INSTQUEUE_REG_0__3__SCAN_IN), .A2(n6098), .B1(n6474), 
        .B2(n6502), .ZN(n6088) );
  OAI211_X1 U7031 ( .C1(n6477), .C2(n6129), .A(n6089), .B(n6088), .ZN(U3023)
         );
  AOI22_X1 U7032 ( .A1(n6479), .A2(n6097), .B1(n6478), .B2(n6096), .ZN(n6091)
         );
  AOI22_X1 U7033 ( .A1(INSTQUEUE_REG_0__4__SCAN_IN), .A2(n6098), .B1(n6481), 
        .B2(n6502), .ZN(n6090) );
  OAI211_X1 U7034 ( .C1(n6485), .C2(n6129), .A(n6091), .B(n6090), .ZN(U3024)
         );
  AOI22_X1 U7035 ( .A1(n3161), .A2(n6097), .B1(n6486), .B2(n6096), .ZN(n6093)
         );
  AOI22_X1 U7036 ( .A1(INSTQUEUE_REG_0__5__SCAN_IN), .A2(n6098), .B1(n6424), 
        .B2(n6502), .ZN(n6092) );
  OAI211_X1 U7037 ( .C1(n6427), .C2(n6129), .A(n6093), .B(n6092), .ZN(U3025)
         );
  AOI22_X1 U7038 ( .A1(n6493), .A2(n6097), .B1(n6492), .B2(n6096), .ZN(n6095)
         );
  AOI22_X1 U7039 ( .A1(INSTQUEUE_REG_0__6__SCAN_IN), .A2(n6098), .B1(n6428), 
        .B2(n6502), .ZN(n6094) );
  OAI211_X1 U7040 ( .C1(n6431), .C2(n6129), .A(n6095), .B(n6094), .ZN(U3026)
         );
  AOI22_X1 U7041 ( .A1(n6501), .A2(n6097), .B1(n6499), .B2(n6096), .ZN(n6100)
         );
  AOI22_X1 U7042 ( .A1(INSTQUEUE_REG_0__7__SCAN_IN), .A2(n6098), .B1(n6435), 
        .B2(n6502), .ZN(n6099) );
  OAI211_X1 U7043 ( .C1(n6439), .C2(n6129), .A(n6100), .B(n6099), .ZN(U3027)
         );
  NOR2_X1 U7044 ( .A1(n6509), .A2(n6106), .ZN(n6124) );
  AOI22_X1 U7045 ( .A1(n6132), .A2(n6456), .B1(n6446), .B2(n6124), .ZN(n6110)
         );
  OAI21_X1 U7046 ( .B1(n6102), .B2(n6852), .A(n6405), .ZN(n6108) );
  AOI21_X1 U7047 ( .B1(n6103), .B2(n6256), .A(n6124), .ZN(n6107) );
  INV_X1 U7048 ( .A(n6107), .ZN(n6105) );
  AOI21_X1 U7049 ( .B1(n6643), .B2(n6106), .A(n6451), .ZN(n6104) );
  OAI21_X1 U7050 ( .B1(n6108), .B2(n6105), .A(n6104), .ZN(n6126) );
  OAI22_X1 U7051 ( .A1(n6108), .A2(n6107), .B1(n6443), .B2(n6106), .ZN(n6125)
         );
  AOI22_X1 U7052 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n6126), .B1(n6445), 
        .B2(n6125), .ZN(n6109) );
  OAI211_X1 U7053 ( .C1(n6459), .C2(n6129), .A(n6110), .B(n6109), .ZN(U3028)
         );
  AOI22_X1 U7054 ( .A1(n6132), .A2(n6372), .B1(n6461), .B2(n6124), .ZN(n6112)
         );
  AOI22_X1 U7055 ( .A1(INSTQUEUE_REG_1__1__SCAN_IN), .A2(n6126), .B1(n6460), 
        .B2(n6125), .ZN(n6111) );
  OAI211_X1 U7056 ( .C1(n6375), .C2(n6129), .A(n6112), .B(n6111), .ZN(U3029)
         );
  AOI22_X1 U7057 ( .A1(n6468), .A2(n6119), .B1(n6467), .B2(n6124), .ZN(n6114)
         );
  AOI22_X1 U7058 ( .A1(INSTQUEUE_REG_1__2__SCAN_IN), .A2(n6126), .B1(n6466), 
        .B2(n6125), .ZN(n6113) );
  OAI211_X1 U7059 ( .C1(n6156), .C2(n6471), .A(n6114), .B(n6113), .ZN(U3030)
         );
  AOI22_X1 U7060 ( .A1(n6119), .A2(n6474), .B1(n6473), .B2(n6124), .ZN(n6116)
         );
  AOI22_X1 U7061 ( .A1(INSTQUEUE_REG_1__3__SCAN_IN), .A2(n6126), .B1(n6472), 
        .B2(n6125), .ZN(n6115) );
  OAI211_X1 U7062 ( .C1(n6156), .C2(n6477), .A(n6116), .B(n6115), .ZN(U3031)
         );
  AOI22_X1 U7063 ( .A1(n6119), .A2(n6481), .B1(n6479), .B2(n6124), .ZN(n6118)
         );
  AOI22_X1 U7064 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n6126), .B1(n6478), 
        .B2(n6125), .ZN(n6117) );
  OAI211_X1 U7065 ( .C1(n6156), .C2(n6485), .A(n6118), .B(n6117), .ZN(U3032)
         );
  AOI22_X1 U7066 ( .A1(n6119), .A2(n6424), .B1(n3161), .B2(n6124), .ZN(n6121)
         );
  AOI22_X1 U7067 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(n6126), .B1(n6486), 
        .B2(n6125), .ZN(n6120) );
  OAI211_X1 U7068 ( .C1(n6156), .C2(n6427), .A(n6121), .B(n6120), .ZN(U3033)
         );
  AOI22_X1 U7069 ( .A1(n6132), .A2(n6494), .B1(n6493), .B2(n6124), .ZN(n6123)
         );
  AOI22_X1 U7070 ( .A1(INSTQUEUE_REG_1__6__SCAN_IN), .A2(n6126), .B1(n6492), 
        .B2(n6125), .ZN(n6122) );
  OAI211_X1 U7071 ( .C1(n6497), .C2(n6129), .A(n6123), .B(n6122), .ZN(U3034)
         );
  AOI22_X1 U7072 ( .A1(n6132), .A2(n6503), .B1(n6501), .B2(n6124), .ZN(n6128)
         );
  AOI22_X1 U7073 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(n6126), .B1(n6499), 
        .B2(n6125), .ZN(n6127) );
  OAI211_X1 U7074 ( .C1(n6508), .C2(n6129), .A(n6128), .B(n6127), .ZN(U3035)
         );
  NOR2_X1 U7075 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6130), .ZN(n6152)
         );
  NAND3_X1 U7076 ( .A1(n6402), .A2(n6294), .A3(n6403), .ZN(n6131) );
  OAI21_X1 U7077 ( .B1(n6133), .B2(n6643), .A(n6131), .ZN(n6151) );
  AOI22_X1 U7078 ( .A1(n6152), .A2(n6446), .B1(n6445), .B2(n6151), .ZN(n6138)
         );
  OAI21_X1 U7079 ( .B1(n6132), .B2(n3182), .A(n6289), .ZN(n6134) );
  AOI21_X1 U7080 ( .B1(n6134), .B2(n6133), .A(STATE2_REG_3__SCAN_IN), .ZN(
        n6136) );
  OAI21_X1 U7081 ( .B1(n6294), .B2(n6443), .A(n6135), .ZN(n6404) );
  NOR2_X1 U7082 ( .A1(n6226), .A2(n6404), .ZN(n6292) );
  OAI21_X1 U7083 ( .B1(n6136), .B2(n6152), .A(n6292), .ZN(n6153) );
  AOI22_X1 U7084 ( .A1(n6153), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n6456), 
        .B2(n3182), .ZN(n6137) );
  OAI211_X1 U7085 ( .C1(n6459), .C2(n6156), .A(n6138), .B(n6137), .ZN(U3036)
         );
  AOI22_X1 U7086 ( .A1(n6461), .A2(n6152), .B1(n6460), .B2(n6151), .ZN(n6140)
         );
  AOI22_X1 U7087 ( .A1(n6153), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n6372), 
        .B2(n3182), .ZN(n6139) );
  OAI211_X1 U7088 ( .C1(n6156), .C2(n6375), .A(n6140), .B(n6139), .ZN(U3037)
         );
  AOI22_X1 U7089 ( .A1(n6152), .A2(n6467), .B1(n6466), .B2(n6151), .ZN(n6142)
         );
  AOI22_X1 U7090 ( .A1(n6153), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n6376), 
        .B2(n3182), .ZN(n6141) );
  OAI211_X1 U7091 ( .C1(n6156), .C2(n6379), .A(n6142), .B(n6141), .ZN(U3038)
         );
  AOI22_X1 U7092 ( .A1(n6473), .A2(n6152), .B1(n6472), .B2(n6151), .ZN(n6144)
         );
  AOI22_X1 U7093 ( .A1(n6153), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n6380), 
        .B2(n3182), .ZN(n6143) );
  OAI211_X1 U7094 ( .C1(n6156), .C2(n6383), .A(n6144), .B(n6143), .ZN(U3039)
         );
  AOI22_X1 U7095 ( .A1(n6479), .A2(n6152), .B1(n6478), .B2(n6151), .ZN(n6146)
         );
  AOI22_X1 U7096 ( .A1(n6153), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n6384), 
        .B2(n3182), .ZN(n6145) );
  OAI211_X1 U7097 ( .C1(n6156), .C2(n6387), .A(n6146), .B(n6145), .ZN(U3040)
         );
  AOI22_X1 U7098 ( .A1(n3161), .A2(n6152), .B1(n6486), .B2(n6151), .ZN(n6148)
         );
  AOI22_X1 U7099 ( .A1(n6153), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n6488), 
        .B2(n3182), .ZN(n6147) );
  OAI211_X1 U7100 ( .C1(n6156), .C2(n6491), .A(n6148), .B(n6147), .ZN(U3041)
         );
  AOI22_X1 U7101 ( .A1(n6493), .A2(n6152), .B1(n6492), .B2(n6151), .ZN(n6150)
         );
  AOI22_X1 U7102 ( .A1(n6153), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n6494), 
        .B2(n3182), .ZN(n6149) );
  OAI211_X1 U7103 ( .C1(n6156), .C2(n6497), .A(n6150), .B(n6149), .ZN(U3042)
         );
  AOI22_X1 U7104 ( .A1(n6501), .A2(n6152), .B1(n6499), .B2(n6151), .ZN(n6155)
         );
  AOI22_X1 U7105 ( .A1(n6153), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n6503), 
        .B2(n3182), .ZN(n6154) );
  OAI211_X1 U7106 ( .C1(n6156), .C2(n6508), .A(n6155), .B(n6154), .ZN(U3043)
         );
  NOR2_X2 U7107 ( .A1(n6157), .A2(n6409), .ZN(n6209) );
  NOR2_X1 U7108 ( .A1(n6509), .A2(n6162), .ZN(n6179) );
  AOI22_X1 U7109 ( .A1(n6456), .A2(n6209), .B1(n6446), .B2(n6179), .ZN(n6166)
         );
  NAND3_X1 U7110 ( .A1(n6360), .A2(n6332), .A3(n6256), .ZN(n6159) );
  INV_X1 U7111 ( .A(n6179), .ZN(n6158) );
  NAND2_X1 U7112 ( .A1(n6159), .A2(n6158), .ZN(n6161) );
  AOI21_X1 U7113 ( .B1(n6162), .B2(n6643), .A(n6451), .ZN(n6160) );
  OAI21_X1 U7114 ( .B1(n6164), .B2(n6161), .A(n6160), .ZN(n6181) );
  INV_X1 U7115 ( .A(n6161), .ZN(n6163) );
  OAI22_X1 U7116 ( .A1(n6164), .A2(n6163), .B1(n6162), .B2(n6443), .ZN(n6180)
         );
  AOI22_X1 U7117 ( .A1(INSTQUEUE_REG_5__0__SCAN_IN), .A2(n6181), .B1(n6445), 
        .B2(n6180), .ZN(n6165) );
  OAI211_X1 U7118 ( .C1(n6459), .C2(n6184), .A(n6166), .B(n6165), .ZN(U3060)
         );
  AOI22_X1 U7119 ( .A1(n6209), .A2(n6372), .B1(n6461), .B2(n6179), .ZN(n6168)
         );
  AOI22_X1 U7120 ( .A1(INSTQUEUE_REG_5__1__SCAN_IN), .A2(n6181), .B1(n6460), 
        .B2(n6180), .ZN(n6167) );
  OAI211_X1 U7121 ( .C1(n6375), .C2(n6184), .A(n6168), .B(n6167), .ZN(U3061)
         );
  AOI22_X1 U7122 ( .A1(n6376), .A2(n6209), .B1(n6467), .B2(n6179), .ZN(n6170)
         );
  AOI22_X1 U7123 ( .A1(INSTQUEUE_REG_5__2__SCAN_IN), .A2(n6181), .B1(n6466), 
        .B2(n6180), .ZN(n6169) );
  OAI211_X1 U7124 ( .C1(n6379), .C2(n6184), .A(n6170), .B(n6169), .ZN(U3062)
         );
  AOI22_X1 U7125 ( .A1(n6209), .A2(n6380), .B1(n6473), .B2(n6179), .ZN(n6172)
         );
  AOI22_X1 U7126 ( .A1(INSTQUEUE_REG_5__3__SCAN_IN), .A2(n6181), .B1(n6472), 
        .B2(n6180), .ZN(n6171) );
  OAI211_X1 U7127 ( .C1(n6383), .C2(n6184), .A(n6172), .B(n6171), .ZN(U3063)
         );
  AOI22_X1 U7128 ( .A1(n6209), .A2(n6384), .B1(n6479), .B2(n6179), .ZN(n6174)
         );
  AOI22_X1 U7129 ( .A1(INSTQUEUE_REG_5__4__SCAN_IN), .A2(n6181), .B1(n6478), 
        .B2(n6180), .ZN(n6173) );
  OAI211_X1 U7130 ( .C1(n6387), .C2(n6184), .A(n6174), .B(n6173), .ZN(U3064)
         );
  AOI22_X1 U7131 ( .A1(n6209), .A2(n6488), .B1(n3161), .B2(n6179), .ZN(n6176)
         );
  AOI22_X1 U7132 ( .A1(INSTQUEUE_REG_5__5__SCAN_IN), .A2(n6181), .B1(n6486), 
        .B2(n6180), .ZN(n6175) );
  OAI211_X1 U7133 ( .C1(n6491), .C2(n6184), .A(n6176), .B(n6175), .ZN(U3065)
         );
  AOI22_X1 U7134 ( .A1(n6209), .A2(n6494), .B1(n6493), .B2(n6179), .ZN(n6178)
         );
  AOI22_X1 U7135 ( .A1(INSTQUEUE_REG_5__6__SCAN_IN), .A2(n6181), .B1(n6492), 
        .B2(n6180), .ZN(n6177) );
  OAI211_X1 U7136 ( .C1(n6497), .C2(n6184), .A(n6178), .B(n6177), .ZN(U3066)
         );
  AOI22_X1 U7137 ( .A1(n6209), .A2(n6503), .B1(n6501), .B2(n6179), .ZN(n6183)
         );
  AOI22_X1 U7138 ( .A1(INSTQUEUE_REG_5__7__SCAN_IN), .A2(n6181), .B1(n6499), 
        .B2(n6180), .ZN(n6182) );
  OAI211_X1 U7139 ( .C1(n6508), .C2(n6184), .A(n6183), .B(n6182), .ZN(U3067)
         );
  NAND3_X1 U7140 ( .A1(n6226), .A2(n6294), .A3(n6403), .ZN(n6185) );
  OAI21_X1 U7141 ( .B1(n6188), .B2(n6643), .A(n6185), .ZN(n6207) );
  NOR2_X1 U7142 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6186), .ZN(n6208)
         );
  AOI22_X1 U7143 ( .A1(n6445), .A2(n6207), .B1(n6446), .B2(n6208), .ZN(n6194)
         );
  OAI21_X1 U7144 ( .B1(n6209), .B2(n6187), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n6189) );
  NAND3_X1 U7145 ( .A1(n6189), .A2(n6405), .A3(n6188), .ZN(n6192) );
  INV_X1 U7146 ( .A(n6208), .ZN(n6190) );
  AOI211_X1 U7147 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6190), .A(n6402), .B(
        n6404), .ZN(n6191) );
  NAND3_X1 U7148 ( .A1(n6403), .A2(n6192), .A3(n6191), .ZN(n6210) );
  AOI22_X1 U7149 ( .A1(INSTQUEUE_REG_6__0__SCAN_IN), .A2(n6210), .B1(n6412), 
        .B2(n6209), .ZN(n6193) );
  OAI211_X1 U7150 ( .C1(n6415), .C2(n6220), .A(n6194), .B(n6193), .ZN(U3068)
         );
  AOI22_X1 U7151 ( .A1(n6461), .A2(n6208), .B1(n6460), .B2(n6207), .ZN(n6196)
         );
  AOI22_X1 U7152 ( .A1(INSTQUEUE_REG_6__1__SCAN_IN), .A2(n6210), .B1(n6462), 
        .B2(n6209), .ZN(n6195) );
  OAI211_X1 U7153 ( .C1(n6465), .C2(n6220), .A(n6196), .B(n6195), .ZN(U3069)
         );
  AOI22_X1 U7154 ( .A1(n6467), .A2(n6208), .B1(n6466), .B2(n6207), .ZN(n6198)
         );
  AOI22_X1 U7155 ( .A1(INSTQUEUE_REG_6__2__SCAN_IN), .A2(n6210), .B1(n6468), 
        .B2(n6209), .ZN(n6197) );
  OAI211_X1 U7156 ( .C1(n6471), .C2(n6220), .A(n6198), .B(n6197), .ZN(U3070)
         );
  AOI22_X1 U7157 ( .A1(n6473), .A2(n6208), .B1(n6472), .B2(n6207), .ZN(n6200)
         );
  AOI22_X1 U7158 ( .A1(INSTQUEUE_REG_6__3__SCAN_IN), .A2(n6210), .B1(n6474), 
        .B2(n6209), .ZN(n6199) );
  OAI211_X1 U7159 ( .C1(n6477), .C2(n6220), .A(n6200), .B(n6199), .ZN(U3071)
         );
  AOI22_X1 U7160 ( .A1(n6479), .A2(n6208), .B1(n6478), .B2(n6207), .ZN(n6202)
         );
  AOI22_X1 U7161 ( .A1(INSTQUEUE_REG_6__4__SCAN_IN), .A2(n6210), .B1(n6481), 
        .B2(n6209), .ZN(n6201) );
  OAI211_X1 U7162 ( .C1(n6485), .C2(n6220), .A(n6202), .B(n6201), .ZN(U3072)
         );
  AOI22_X1 U7163 ( .A1(n3161), .A2(n6208), .B1(n6486), .B2(n6207), .ZN(n6204)
         );
  AOI22_X1 U7164 ( .A1(INSTQUEUE_REG_6__5__SCAN_IN), .A2(n6210), .B1(n6424), 
        .B2(n6209), .ZN(n6203) );
  OAI211_X1 U7165 ( .C1(n6427), .C2(n6220), .A(n6204), .B(n6203), .ZN(U3073)
         );
  AOI22_X1 U7166 ( .A1(n6493), .A2(n6208), .B1(n6492), .B2(n6207), .ZN(n6206)
         );
  AOI22_X1 U7167 ( .A1(INSTQUEUE_REG_6__6__SCAN_IN), .A2(n6210), .B1(n6428), 
        .B2(n6209), .ZN(n6205) );
  OAI211_X1 U7168 ( .C1(n6431), .C2(n6220), .A(n6206), .B(n6205), .ZN(U3074)
         );
  AOI22_X1 U7169 ( .A1(n6501), .A2(n6208), .B1(n6499), .B2(n6207), .ZN(n6212)
         );
  AOI22_X1 U7170 ( .A1(INSTQUEUE_REG_6__7__SCAN_IN), .A2(n6210), .B1(n6435), 
        .B2(n6209), .ZN(n6211) );
  OAI211_X1 U7171 ( .C1(n6439), .C2(n6220), .A(n6212), .B(n6211), .ZN(U3075)
         );
  AOI22_X1 U7172 ( .A1(n6446), .A2(n6215), .B1(n6456), .B2(n6249), .ZN(n6214)
         );
  AOI22_X1 U7173 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n6217), .B1(n6445), 
        .B2(n6216), .ZN(n6213) );
  OAI211_X1 U7174 ( .C1(n6459), .C2(n6220), .A(n6214), .B(n6213), .ZN(U3076)
         );
  AOI22_X1 U7175 ( .A1(n6467), .A2(n6215), .B1(n6376), .B2(n6249), .ZN(n6219)
         );
  AOI22_X1 U7176 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n6217), .B1(n6466), 
        .B2(n6216), .ZN(n6218) );
  OAI211_X1 U7177 ( .C1(n6379), .C2(n6220), .A(n6219), .B(n6218), .ZN(U3078)
         );
  NAND2_X1 U7178 ( .A1(n6254), .A2(n6409), .ZN(n6277) );
  NOR2_X1 U7179 ( .A1(n6399), .A2(n6258), .ZN(n6229) );
  INV_X1 U7180 ( .A(n6229), .ZN(n6225) );
  INV_X1 U7181 ( .A(n6223), .ZN(n6224) );
  NAND2_X1 U7182 ( .A1(n6224), .A2(n6401), .ZN(n6329) );
  OAI22_X1 U7183 ( .A1(n6225), .A2(n6643), .B1(n6335), .B2(n6329), .ZN(n6247)
         );
  NAND3_X1 U7184 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6521), .A3(n6517), .ZN(n6263) );
  NOR2_X1 U7185 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6263), .ZN(n6248)
         );
  AOI22_X1 U7186 ( .A1(n6445), .A2(n6247), .B1(n6446), .B2(n6248), .ZN(n6234)
         );
  INV_X1 U7187 ( .A(n6226), .ZN(n6400) );
  AOI21_X1 U7188 ( .B1(n6329), .B2(STATE2_REG_2__SCAN_IN), .A(n6227), .ZN(
        n6334) );
  OAI211_X1 U7189 ( .C1(n6615), .C2(n6248), .A(n6400), .B(n6334), .ZN(n6232)
         );
  INV_X1 U7190 ( .A(n6249), .ZN(n6228) );
  NAND3_X1 U7191 ( .A1(n6277), .A2(n6405), .A3(n6228), .ZN(n6230) );
  AOI21_X1 U7192 ( .B1(n6230), .B2(n6289), .A(n6229), .ZN(n6231) );
  AOI22_X1 U7193 ( .A1(n6250), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n6412), 
        .B2(n6249), .ZN(n6233) );
  OAI211_X1 U7194 ( .C1(n6415), .C2(n6277), .A(n6234), .B(n6233), .ZN(U3084)
         );
  AOI22_X1 U7195 ( .A1(n6461), .A2(n6248), .B1(n6460), .B2(n6247), .ZN(n6236)
         );
  AOI22_X1 U7196 ( .A1(n6250), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n6462), 
        .B2(n6249), .ZN(n6235) );
  OAI211_X1 U7197 ( .C1(n6465), .C2(n6277), .A(n6236), .B(n6235), .ZN(U3085)
         );
  AOI22_X1 U7198 ( .A1(n6467), .A2(n6248), .B1(n6466), .B2(n6247), .ZN(n6238)
         );
  AOI22_X1 U7199 ( .A1(n6250), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n6468), 
        .B2(n6249), .ZN(n6237) );
  OAI211_X1 U7200 ( .C1(n6471), .C2(n6277), .A(n6238), .B(n6237), .ZN(U3086)
         );
  AOI22_X1 U7201 ( .A1(n6473), .A2(n6248), .B1(n6472), .B2(n6247), .ZN(n6240)
         );
  AOI22_X1 U7202 ( .A1(n6250), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n6474), 
        .B2(n6249), .ZN(n6239) );
  OAI211_X1 U7203 ( .C1(n6477), .C2(n6277), .A(n6240), .B(n6239), .ZN(U3087)
         );
  AOI22_X1 U7204 ( .A1(n6479), .A2(n6248), .B1(n6478), .B2(n6247), .ZN(n6242)
         );
  AOI22_X1 U7205 ( .A1(n6250), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n6481), 
        .B2(n6249), .ZN(n6241) );
  OAI211_X1 U7206 ( .C1(n6485), .C2(n6277), .A(n6242), .B(n6241), .ZN(U3088)
         );
  AOI22_X1 U7207 ( .A1(n3161), .A2(n6248), .B1(n6486), .B2(n6247), .ZN(n6244)
         );
  AOI22_X1 U7208 ( .A1(n6250), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n6424), 
        .B2(n6249), .ZN(n6243) );
  OAI211_X1 U7209 ( .C1(n6427), .C2(n6277), .A(n6244), .B(n6243), .ZN(U3089)
         );
  AOI22_X1 U7210 ( .A1(n6493), .A2(n6248), .B1(n6492), .B2(n6247), .ZN(n6246)
         );
  AOI22_X1 U7211 ( .A1(n6250), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n6428), 
        .B2(n6249), .ZN(n6245) );
  OAI211_X1 U7212 ( .C1(n6431), .C2(n6277), .A(n6246), .B(n6245), .ZN(U3090)
         );
  AOI22_X1 U7213 ( .A1(n6501), .A2(n6248), .B1(n6499), .B2(n6247), .ZN(n6252)
         );
  AOI22_X1 U7214 ( .A1(n6250), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n6435), 
        .B2(n6249), .ZN(n6251) );
  OAI211_X1 U7215 ( .C1(n6439), .C2(n6277), .A(n6252), .B(n6251), .ZN(U3091)
         );
  INV_X1 U7216 ( .A(n6277), .ZN(n6283) );
  NOR2_X1 U7217 ( .A1(n6509), .A2(n6263), .ZN(n6282) );
  AOI22_X1 U7218 ( .A1(n6412), .A2(n6283), .B1(n6446), .B2(n6282), .ZN(n6267)
         );
  INV_X1 U7219 ( .A(n6254), .ZN(n6255) );
  OAI21_X1 U7220 ( .B1(n6255), .B2(n6852), .A(n6405), .ZN(n6264) );
  NAND2_X1 U7221 ( .A1(n6257), .A2(n6256), .ZN(n6442) );
  OR2_X1 U7222 ( .A1(n6442), .A2(n6258), .ZN(n6260) );
  INV_X1 U7223 ( .A(n6282), .ZN(n6259) );
  AND2_X1 U7224 ( .A1(n6260), .A2(n6259), .ZN(n6265) );
  INV_X1 U7225 ( .A(n6265), .ZN(n6262) );
  AOI21_X1 U7226 ( .B1(n6643), .B2(n6263), .A(n6451), .ZN(n6261) );
  OAI21_X1 U7227 ( .B1(n6264), .B2(n6262), .A(n6261), .ZN(n6285) );
  OAI22_X1 U7228 ( .A1(n6265), .A2(n6264), .B1(n6443), .B2(n6263), .ZN(n6284)
         );
  AOI22_X1 U7229 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n6285), .B1(n6445), 
        .B2(n6284), .ZN(n6266) );
  OAI211_X1 U7230 ( .C1(n6415), .C2(n6318), .A(n6267), .B(n6266), .ZN(U3092)
         );
  AOI22_X1 U7231 ( .A1(n6283), .A2(n6462), .B1(n6461), .B2(n6282), .ZN(n6269)
         );
  AOI22_X1 U7232 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n6285), .B1(n6460), 
        .B2(n6284), .ZN(n6268) );
  OAI211_X1 U7233 ( .C1(n6465), .C2(n6318), .A(n6269), .B(n6268), .ZN(U3093)
         );
  AOI22_X1 U7234 ( .A1(n6468), .A2(n6283), .B1(n6467), .B2(n6282), .ZN(n6271)
         );
  AOI22_X1 U7235 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n6285), .B1(n6466), 
        .B2(n6284), .ZN(n6270) );
  OAI211_X1 U7236 ( .C1(n6471), .C2(n6318), .A(n6271), .B(n6270), .ZN(U3094)
         );
  AOI22_X1 U7237 ( .A1(n6283), .A2(n6474), .B1(n6473), .B2(n6282), .ZN(n6273)
         );
  AOI22_X1 U7238 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n6285), .B1(n6472), 
        .B2(n6284), .ZN(n6272) );
  OAI211_X1 U7239 ( .C1(n6477), .C2(n6318), .A(n6273), .B(n6272), .ZN(U3095)
         );
  INV_X1 U7240 ( .A(n6318), .ZN(n6274) );
  AOI22_X1 U7241 ( .A1(n6274), .A2(n6384), .B1(n6479), .B2(n6282), .ZN(n6276)
         );
  AOI22_X1 U7242 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n6285), .B1(n6478), 
        .B2(n6284), .ZN(n6275) );
  OAI211_X1 U7243 ( .C1(n6387), .C2(n6277), .A(n6276), .B(n6275), .ZN(U3096)
         );
  AOI22_X1 U7244 ( .A1(n6283), .A2(n6424), .B1(n3161), .B2(n6282), .ZN(n6279)
         );
  AOI22_X1 U7245 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n6285), .B1(n6486), 
        .B2(n6284), .ZN(n6278) );
  OAI211_X1 U7246 ( .C1(n6427), .C2(n6318), .A(n6279), .B(n6278), .ZN(U3097)
         );
  AOI22_X1 U7247 ( .A1(n6283), .A2(n6428), .B1(n6493), .B2(n6282), .ZN(n6281)
         );
  AOI22_X1 U7248 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n6285), .B1(n6492), 
        .B2(n6284), .ZN(n6280) );
  OAI211_X1 U7249 ( .C1(n6431), .C2(n6318), .A(n6281), .B(n6280), .ZN(U3098)
         );
  AOI22_X1 U7250 ( .A1(n6283), .A2(n6435), .B1(n6501), .B2(n6282), .ZN(n6287)
         );
  AOI22_X1 U7251 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n6285), .B1(n6499), 
        .B2(n6284), .ZN(n6286) );
  OAI211_X1 U7252 ( .C1(n6439), .C2(n6318), .A(n6287), .B(n6286), .ZN(U3099)
         );
  NOR2_X1 U7253 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6288), .ZN(n6313)
         );
  AOI22_X1 U7254 ( .A1(n6456), .A2(n6312), .B1(n6446), .B2(n6313), .ZN(n6299)
         );
  INV_X1 U7255 ( .A(n6312), .ZN(n6327) );
  NAND3_X1 U7256 ( .A1(n6327), .A2(n6318), .A3(n6405), .ZN(n6290) );
  NAND2_X1 U7257 ( .A1(n6290), .A2(n6289), .ZN(n6293) );
  AOI22_X1 U7258 ( .A1(n6293), .A2(n6296), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6403), .ZN(n6291) );
  OAI211_X1 U7259 ( .C1(n6313), .C2(n6615), .A(n6292), .B(n6291), .ZN(n6315)
         );
  INV_X1 U7260 ( .A(n6293), .ZN(n6297) );
  NAND3_X1 U7261 ( .A1(n6402), .A2(n6294), .A3(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6295) );
  OAI21_X1 U7262 ( .B1(n6297), .B2(n6296), .A(n6295), .ZN(n6314) );
  AOI22_X1 U7263 ( .A1(INSTQUEUE_REG_10__0__SCAN_IN), .A2(n6315), .B1(n6445), 
        .B2(n6314), .ZN(n6298) );
  OAI211_X1 U7264 ( .C1(n6459), .C2(n6318), .A(n6299), .B(n6298), .ZN(U3100)
         );
  AOI22_X1 U7265 ( .A1(n6461), .A2(n6313), .B1(n6312), .B2(n6372), .ZN(n6301)
         );
  AOI22_X1 U7266 ( .A1(INSTQUEUE_REG_10__1__SCAN_IN), .A2(n6315), .B1(n6460), 
        .B2(n6314), .ZN(n6300) );
  OAI211_X1 U7267 ( .C1(n6375), .C2(n6318), .A(n6301), .B(n6300), .ZN(U3101)
         );
  AOI22_X1 U7268 ( .A1(n6376), .A2(n6312), .B1(n6467), .B2(n6313), .ZN(n6303)
         );
  AOI22_X1 U7269 ( .A1(INSTQUEUE_REG_10__2__SCAN_IN), .A2(n6315), .B1(n6466), 
        .B2(n6314), .ZN(n6302) );
  OAI211_X1 U7270 ( .C1(n6379), .C2(n6318), .A(n6303), .B(n6302), .ZN(U3102)
         );
  AOI22_X1 U7271 ( .A1(n6473), .A2(n6313), .B1(n6312), .B2(n6380), .ZN(n6305)
         );
  AOI22_X1 U7272 ( .A1(INSTQUEUE_REG_10__3__SCAN_IN), .A2(n6315), .B1(n6472), 
        .B2(n6314), .ZN(n6304) );
  OAI211_X1 U7273 ( .C1(n6383), .C2(n6318), .A(n6305), .B(n6304), .ZN(U3103)
         );
  AOI22_X1 U7274 ( .A1(n6479), .A2(n6313), .B1(n6312), .B2(n6384), .ZN(n6307)
         );
  AOI22_X1 U7275 ( .A1(INSTQUEUE_REG_10__4__SCAN_IN), .A2(n6315), .B1(n6478), 
        .B2(n6314), .ZN(n6306) );
  OAI211_X1 U7276 ( .C1(n6387), .C2(n6318), .A(n6307), .B(n6306), .ZN(U3104)
         );
  AOI22_X1 U7277 ( .A1(n3161), .A2(n6313), .B1(n6312), .B2(n6488), .ZN(n6309)
         );
  AOI22_X1 U7278 ( .A1(INSTQUEUE_REG_10__5__SCAN_IN), .A2(n6315), .B1(n6486), 
        .B2(n6314), .ZN(n6308) );
  OAI211_X1 U7279 ( .C1(n6491), .C2(n6318), .A(n6309), .B(n6308), .ZN(U3105)
         );
  AOI22_X1 U7280 ( .A1(n6493), .A2(n6313), .B1(n6312), .B2(n6494), .ZN(n6311)
         );
  AOI22_X1 U7281 ( .A1(INSTQUEUE_REG_10__6__SCAN_IN), .A2(n6315), .B1(n6492), 
        .B2(n6314), .ZN(n6310) );
  OAI211_X1 U7282 ( .C1(n6497), .C2(n6318), .A(n6311), .B(n6310), .ZN(U3106)
         );
  AOI22_X1 U7283 ( .A1(n6501), .A2(n6313), .B1(n6312), .B2(n6503), .ZN(n6317)
         );
  AOI22_X1 U7284 ( .A1(INSTQUEUE_REG_10__7__SCAN_IN), .A2(n6315), .B1(n6499), 
        .B2(n6314), .ZN(n6316) );
  OAI211_X1 U7285 ( .C1(n6508), .C2(n6318), .A(n6317), .B(n6316), .ZN(U3107)
         );
  INV_X1 U7286 ( .A(n6319), .ZN(n6322) );
  AOI22_X1 U7287 ( .A1(n6461), .A2(n6322), .B1(n6356), .B2(n6372), .ZN(n6321)
         );
  AOI22_X1 U7288 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6324), .B1(n6460), 
        .B2(n6323), .ZN(n6320) );
  OAI211_X1 U7289 ( .C1(n6375), .C2(n6327), .A(n6321), .B(n6320), .ZN(U3109)
         );
  AOI22_X1 U7290 ( .A1(n6493), .A2(n6322), .B1(n6356), .B2(n6494), .ZN(n6326)
         );
  AOI22_X1 U7291 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6324), .B1(n6492), 
        .B2(n6323), .ZN(n6325) );
  OAI211_X1 U7292 ( .C1(n6497), .C2(n6327), .A(n6326), .B(n6325), .ZN(U3114)
         );
  NAND2_X1 U7293 ( .A1(n6368), .A2(n6409), .ZN(n6397) );
  INV_X1 U7294 ( .A(n6328), .ZN(n6330) );
  OAI22_X1 U7295 ( .A1(n6330), .A2(n6399), .B1(n6329), .B2(n6400), .ZN(n6354)
         );
  NOR2_X1 U7296 ( .A1(n6403), .A2(n6362), .ZN(n6367) );
  AND2_X1 U7297 ( .A1(n6509), .A2(n6367), .ZN(n6355) );
  AOI22_X1 U7298 ( .A1(n6445), .A2(n6354), .B1(n6446), .B2(n6355), .ZN(n6341)
         );
  AOI21_X1 U7299 ( .B1(n6397), .B2(n6331), .A(n6852), .ZN(n6339) );
  OAI21_X1 U7300 ( .B1(n6333), .B2(n6332), .A(n6405), .ZN(n6338) );
  OAI211_X1 U7301 ( .C1(n6615), .C2(n6355), .A(n6335), .B(n6334), .ZN(n6336)
         );
  INV_X1 U7302 ( .A(n6336), .ZN(n6337) );
  OAI21_X1 U7303 ( .B1(n6339), .B2(n6338), .A(n6337), .ZN(n6357) );
  AOI22_X1 U7304 ( .A1(n6357), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n6412), 
        .B2(n6356), .ZN(n6340) );
  OAI211_X1 U7305 ( .C1(n6415), .C2(n6397), .A(n6341), .B(n6340), .ZN(U3116)
         );
  AOI22_X1 U7306 ( .A1(n6461), .A2(n6355), .B1(n6460), .B2(n6354), .ZN(n6343)
         );
  AOI22_X1 U7307 ( .A1(n6357), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n6462), 
        .B2(n6356), .ZN(n6342) );
  OAI211_X1 U7308 ( .C1(n6465), .C2(n6397), .A(n6343), .B(n6342), .ZN(U3117)
         );
  AOI22_X1 U7309 ( .A1(n6467), .A2(n6355), .B1(n6466), .B2(n6354), .ZN(n6345)
         );
  AOI22_X1 U7310 ( .A1(n6357), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n6468), 
        .B2(n6356), .ZN(n6344) );
  OAI211_X1 U7311 ( .C1(n6471), .C2(n6397), .A(n6345), .B(n6344), .ZN(U3118)
         );
  AOI22_X1 U7312 ( .A1(n6473), .A2(n6355), .B1(n6472), .B2(n6354), .ZN(n6347)
         );
  AOI22_X1 U7313 ( .A1(n6357), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n6474), 
        .B2(n6356), .ZN(n6346) );
  OAI211_X1 U7314 ( .C1(n6477), .C2(n6397), .A(n6347), .B(n6346), .ZN(U3119)
         );
  AOI22_X1 U7315 ( .A1(n6479), .A2(n6355), .B1(n6478), .B2(n6354), .ZN(n6349)
         );
  AOI22_X1 U7316 ( .A1(n6357), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n6481), 
        .B2(n6356), .ZN(n6348) );
  OAI211_X1 U7317 ( .C1(n6485), .C2(n6397), .A(n6349), .B(n6348), .ZN(U3120)
         );
  AOI22_X1 U7318 ( .A1(n3161), .A2(n6355), .B1(n6486), .B2(n6354), .ZN(n6351)
         );
  AOI22_X1 U7319 ( .A1(n6357), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n6424), 
        .B2(n6356), .ZN(n6350) );
  OAI211_X1 U7320 ( .C1(n6427), .C2(n6397), .A(n6351), .B(n6350), .ZN(U3121)
         );
  AOI22_X1 U7321 ( .A1(n6493), .A2(n6355), .B1(n6492), .B2(n6354), .ZN(n6353)
         );
  AOI22_X1 U7322 ( .A1(n6357), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n6428), 
        .B2(n6356), .ZN(n6352) );
  OAI211_X1 U7323 ( .C1(n6431), .C2(n6397), .A(n6353), .B(n6352), .ZN(U3122)
         );
  AOI22_X1 U7324 ( .A1(n6501), .A2(n6355), .B1(n6499), .B2(n6354), .ZN(n6359)
         );
  AOI22_X1 U7325 ( .A1(n6357), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n6435), 
        .B2(n6356), .ZN(n6358) );
  OAI211_X1 U7326 ( .C1(n6439), .C2(n6397), .A(n6359), .B(n6358), .ZN(U3123)
         );
  INV_X1 U7327 ( .A(n6442), .ZN(n6361) );
  AND2_X1 U7328 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6367), .ZN(n6393)
         );
  AOI21_X1 U7329 ( .B1(n6361), .B2(n6360), .A(n6393), .ZN(n6364) );
  NAND2_X1 U7330 ( .A1(STATE2_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6363) );
  OAI22_X1 U7331 ( .A1(n6364), .A2(n6643), .B1(n6363), .B2(n6362), .ZN(n6392)
         );
  AOI22_X1 U7332 ( .A1(n6445), .A2(n6392), .B1(n6446), .B2(n6393), .ZN(n6371)
         );
  NAND2_X1 U7333 ( .A1(n6364), .A2(n6408), .ZN(n6366) );
  INV_X1 U7334 ( .A(n6451), .ZN(n6365) );
  OAI221_X1 U7335 ( .B1(n6405), .B2(n6367), .C1(n6643), .C2(n6366), .A(n6365), 
        .ZN(n6394) );
  INV_X1 U7336 ( .A(n6368), .ZN(n6369) );
  NOR2_X2 U7337 ( .A1(n6369), .A2(n6409), .ZN(n6434) );
  AOI22_X1 U7338 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n6394), .B1(n6456), 
        .B2(n6434), .ZN(n6370) );
  OAI211_X1 U7339 ( .C1(n6459), .C2(n6397), .A(n6371), .B(n6370), .ZN(U3124)
         );
  AOI22_X1 U7340 ( .A1(n6461), .A2(n6393), .B1(n6460), .B2(n6392), .ZN(n6374)
         );
  AOI22_X1 U7341 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n6394), .B1(n6372), 
        .B2(n6434), .ZN(n6373) );
  OAI211_X1 U7342 ( .C1(n6375), .C2(n6397), .A(n6374), .B(n6373), .ZN(U3125)
         );
  AOI22_X1 U7343 ( .A1(n6467), .A2(n6393), .B1(n6466), .B2(n6392), .ZN(n6378)
         );
  AOI22_X1 U7344 ( .A1(INSTQUEUE_REG_13__2__SCAN_IN), .A2(n6394), .B1(n6376), 
        .B2(n6434), .ZN(n6377) );
  OAI211_X1 U7345 ( .C1(n6379), .C2(n6397), .A(n6378), .B(n6377), .ZN(U3126)
         );
  AOI22_X1 U7346 ( .A1(n6473), .A2(n6393), .B1(n6472), .B2(n6392), .ZN(n6382)
         );
  AOI22_X1 U7347 ( .A1(INSTQUEUE_REG_13__3__SCAN_IN), .A2(n6394), .B1(n6380), 
        .B2(n6434), .ZN(n6381) );
  OAI211_X1 U7348 ( .C1(n6383), .C2(n6397), .A(n6382), .B(n6381), .ZN(U3127)
         );
  AOI22_X1 U7349 ( .A1(n6479), .A2(n6393), .B1(n6478), .B2(n6392), .ZN(n6386)
         );
  AOI22_X1 U7350 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n6394), .B1(n6384), 
        .B2(n6434), .ZN(n6385) );
  OAI211_X1 U7351 ( .C1(n6387), .C2(n6397), .A(n6386), .B(n6385), .ZN(U3128)
         );
  AOI22_X1 U7352 ( .A1(n3161), .A2(n6393), .B1(n6486), .B2(n6392), .ZN(n6389)
         );
  AOI22_X1 U7353 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(n6394), .B1(n6488), 
        .B2(n6434), .ZN(n6388) );
  OAI211_X1 U7354 ( .C1(n6491), .C2(n6397), .A(n6389), .B(n6388), .ZN(U3129)
         );
  AOI22_X1 U7355 ( .A1(n6493), .A2(n6393), .B1(n6492), .B2(n6392), .ZN(n6391)
         );
  AOI22_X1 U7356 ( .A1(INSTQUEUE_REG_13__6__SCAN_IN), .A2(n6394), .B1(n6494), 
        .B2(n6434), .ZN(n6390) );
  OAI211_X1 U7357 ( .C1(n6497), .C2(n6397), .A(n6391), .B(n6390), .ZN(U3130)
         );
  AOI22_X1 U7358 ( .A1(n6501), .A2(n6393), .B1(n6499), .B2(n6392), .ZN(n6396)
         );
  AOI22_X1 U7359 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n6394), .B1(n6503), 
        .B2(n6434), .ZN(n6395) );
  OAI211_X1 U7360 ( .C1(n6508), .C2(n6397), .A(n6396), .B(n6395), .ZN(U3131)
         );
  OAI33_X1 U7361 ( .A1(n6403), .A2(n6401), .A3(n6400), .B1(n6441), .B2(n6643), 
        .B3(n6399), .ZN(n6433) );
  NOR2_X1 U7362 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6452), .ZN(n6432)
         );
  AOI22_X1 U7363 ( .A1(n6445), .A2(n3180), .B1(n6446), .B2(n6432), .ZN(n6414)
         );
  NOR3_X1 U7364 ( .A1(n6404), .A2(n6403), .A3(n6402), .ZN(n6411) );
  NAND2_X1 U7365 ( .A1(n6405), .A2(n6441), .ZN(n6406) );
  AOI21_X1 U7366 ( .B1(n6480), .B2(STATEBS16_REG_SCAN_IN), .A(n6406), .ZN(
        n6407) );
  OAI21_X1 U7367 ( .B1(n6409), .B2(n6408), .A(n6407), .ZN(n6410) );
  OAI211_X1 U7368 ( .C1(n6432), .C2(n6615), .A(n6411), .B(n6410), .ZN(n6436)
         );
  AOI22_X1 U7369 ( .A1(INSTQUEUE_REG_14__0__SCAN_IN), .A2(n6436), .B1(n6412), 
        .B2(n6434), .ZN(n6413) );
  OAI211_X1 U7370 ( .C1(n6415), .C2(n6507), .A(n6414), .B(n6413), .ZN(U3132)
         );
  AOI22_X1 U7371 ( .A1(n3180), .A2(n6460), .B1(n6461), .B2(n6432), .ZN(n6417)
         );
  AOI22_X1 U7372 ( .A1(INSTQUEUE_REG_14__1__SCAN_IN), .A2(n6436), .B1(n6462), 
        .B2(n6434), .ZN(n6416) );
  OAI211_X1 U7373 ( .C1(n6465), .C2(n6507), .A(n6417), .B(n6416), .ZN(U3133)
         );
  AOI22_X1 U7374 ( .A1(n6467), .A2(n6432), .B1(n6466), .B2(n3180), .ZN(n6419)
         );
  AOI22_X1 U7375 ( .A1(INSTQUEUE_REG_14__2__SCAN_IN), .A2(n6436), .B1(n6468), 
        .B2(n6434), .ZN(n6418) );
  OAI211_X1 U7376 ( .C1(n6471), .C2(n6507), .A(n6419), .B(n6418), .ZN(U3134)
         );
  AOI22_X1 U7377 ( .A1(n3180), .A2(n6472), .B1(n6473), .B2(n6432), .ZN(n6421)
         );
  AOI22_X1 U7378 ( .A1(INSTQUEUE_REG_14__3__SCAN_IN), .A2(n6436), .B1(n6474), 
        .B2(n6434), .ZN(n6420) );
  OAI211_X1 U7379 ( .C1(n6477), .C2(n6507), .A(n6421), .B(n6420), .ZN(U3135)
         );
  AOI22_X1 U7380 ( .A1(n3180), .A2(n6478), .B1(n6479), .B2(n6432), .ZN(n6423)
         );
  AOI22_X1 U7381 ( .A1(INSTQUEUE_REG_14__4__SCAN_IN), .A2(n6436), .B1(n6481), 
        .B2(n6434), .ZN(n6422) );
  OAI211_X1 U7382 ( .C1(n6485), .C2(n6507), .A(n6423), .B(n6422), .ZN(U3136)
         );
  AOI22_X1 U7383 ( .A1(n3180), .A2(n6486), .B1(n3161), .B2(n6432), .ZN(n6426)
         );
  AOI22_X1 U7384 ( .A1(INSTQUEUE_REG_14__5__SCAN_IN), .A2(n6436), .B1(n6424), 
        .B2(n6434), .ZN(n6425) );
  OAI211_X1 U7385 ( .C1(n6427), .C2(n6507), .A(n6426), .B(n6425), .ZN(U3137)
         );
  AOI22_X1 U7386 ( .A1(n3180), .A2(n6492), .B1(n6493), .B2(n6432), .ZN(n6430)
         );
  AOI22_X1 U7387 ( .A1(INSTQUEUE_REG_14__6__SCAN_IN), .A2(n6436), .B1(n6428), 
        .B2(n6434), .ZN(n6429) );
  OAI211_X1 U7388 ( .C1(n6431), .C2(n6507), .A(n6430), .B(n6429), .ZN(U3138)
         );
  AOI22_X1 U7389 ( .A1(n3180), .A2(n6499), .B1(n6501), .B2(n6432), .ZN(n6438)
         );
  AOI22_X1 U7390 ( .A1(INSTQUEUE_REG_14__7__SCAN_IN), .A2(n6436), .B1(n6435), 
        .B2(n6434), .ZN(n6437) );
  OAI211_X1 U7391 ( .C1(n6439), .C2(n6507), .A(n6438), .B(n6437), .ZN(U3139)
         );
  OAI21_X1 U7392 ( .B1(n6442), .B2(n6441), .A(n6440), .ZN(n6454) );
  INV_X1 U7393 ( .A(n6454), .ZN(n6444) );
  OAI22_X1 U7394 ( .A1(n6444), .A2(n6643), .B1(n6452), .B2(n6443), .ZN(n6498)
         );
  AOI22_X1 U7395 ( .A1(n6500), .A2(n6446), .B1(n6445), .B2(n6498), .ZN(n6458)
         );
  AOI21_X1 U7396 ( .B1(n6448), .B2(n4666), .A(n6447), .ZN(n6450) );
  NOR2_X1 U7397 ( .A1(n6450), .A2(n6449), .ZN(n6455) );
  AOI21_X1 U7398 ( .B1(n6452), .B2(n6643), .A(n6451), .ZN(n6453) );
  OAI21_X1 U7399 ( .B1(n6455), .B2(n6454), .A(n6453), .ZN(n6504) );
  AOI22_X1 U7400 ( .A1(INSTQUEUE_REG_15__0__SCAN_IN), .A2(n6504), .B1(n6456), 
        .B2(n6502), .ZN(n6457) );
  OAI211_X1 U7401 ( .C1(n6459), .C2(n6507), .A(n6458), .B(n6457), .ZN(U3140)
         );
  AOI22_X1 U7402 ( .A1(n6461), .A2(n6500), .B1(n6460), .B2(n6498), .ZN(n6464)
         );
  AOI22_X1 U7403 ( .A1(INSTQUEUE_REG_15__1__SCAN_IN), .A2(n6504), .B1(n6462), 
        .B2(n6480), .ZN(n6463) );
  OAI211_X1 U7404 ( .C1(n6465), .C2(n6484), .A(n6464), .B(n6463), .ZN(U3141)
         );
  AOI22_X1 U7405 ( .A1(n6500), .A2(n6467), .B1(n6466), .B2(n6498), .ZN(n6470)
         );
  AOI22_X1 U7406 ( .A1(INSTQUEUE_REG_15__2__SCAN_IN), .A2(n6504), .B1(n6468), 
        .B2(n6480), .ZN(n6469) );
  OAI211_X1 U7407 ( .C1(n6471), .C2(n6484), .A(n6470), .B(n6469), .ZN(U3142)
         );
  AOI22_X1 U7408 ( .A1(n6473), .A2(n6500), .B1(n6472), .B2(n6498), .ZN(n6476)
         );
  AOI22_X1 U7409 ( .A1(INSTQUEUE_REG_15__3__SCAN_IN), .A2(n6504), .B1(n6474), 
        .B2(n6480), .ZN(n6475) );
  OAI211_X1 U7410 ( .C1(n6477), .C2(n6484), .A(n6476), .B(n6475), .ZN(U3143)
         );
  AOI22_X1 U7411 ( .A1(n6479), .A2(n6500), .B1(n6478), .B2(n6498), .ZN(n6483)
         );
  AOI22_X1 U7412 ( .A1(INSTQUEUE_REG_15__4__SCAN_IN), .A2(n6504), .B1(n6481), 
        .B2(n6480), .ZN(n6482) );
  OAI211_X1 U7413 ( .C1(n6485), .C2(n6484), .A(n6483), .B(n6482), .ZN(U3144)
         );
  AOI22_X1 U7414 ( .A1(n3161), .A2(n6500), .B1(n6486), .B2(n6498), .ZN(n6490)
         );
  AOI22_X1 U7415 ( .A1(INSTQUEUE_REG_15__5__SCAN_IN), .A2(n6504), .B1(n6488), 
        .B2(n6502), .ZN(n6489) );
  OAI211_X1 U7416 ( .C1(n6491), .C2(n6507), .A(n6490), .B(n6489), .ZN(U3145)
         );
  AOI22_X1 U7417 ( .A1(n6493), .A2(n6500), .B1(n6492), .B2(n6498), .ZN(n6496)
         );
  AOI22_X1 U7418 ( .A1(INSTQUEUE_REG_15__6__SCAN_IN), .A2(n6504), .B1(n6494), 
        .B2(n6502), .ZN(n6495) );
  OAI211_X1 U7419 ( .C1(n6497), .C2(n6507), .A(n6496), .B(n6495), .ZN(U3146)
         );
  AOI22_X1 U7420 ( .A1(n6501), .A2(n6500), .B1(n6499), .B2(n6498), .ZN(n6506)
         );
  AOI22_X1 U7421 ( .A1(INSTQUEUE_REG_15__7__SCAN_IN), .A2(n6504), .B1(n6503), 
        .B2(n6502), .ZN(n6505) );
  OAI211_X1 U7422 ( .C1(n6508), .C2(n6507), .A(n6506), .B(n6505), .ZN(U3147)
         );
  AOI21_X1 U7423 ( .B1(n6622), .B2(n6510), .A(n6509), .ZN(n6513) );
  INV_X1 U7424 ( .A(n6511), .ZN(n6512) );
  NAND2_X1 U7425 ( .A1(n6512), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n6633) );
  OAI211_X1 U7426 ( .C1(n6624), .C2(n6623), .A(n6513), .B(n6633), .ZN(n6516)
         );
  OAI211_X1 U7427 ( .C1(n6517), .C2(n6516), .A(n6515), .B(n6514), .ZN(n6519)
         );
  NAND2_X1 U7428 ( .A1(n6517), .A2(n6516), .ZN(n6518) );
  NAND2_X1 U7429 ( .A1(n6519), .A2(n6518), .ZN(n6522) );
  AOI21_X1 U7430 ( .B1(n6522), .B2(n6521), .A(n6520), .ZN(n6524) );
  NOR2_X1 U7431 ( .A1(n6522), .A2(n6521), .ZN(n6523) );
  OAI22_X1 U7432 ( .A1(n6524), .A2(n6523), .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n6525), .ZN(n6535) );
  AOI21_X1 U7433 ( .B1(n6525), .B2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6534) );
  INV_X1 U7434 ( .A(n6526), .ZN(n6529) );
  OAI21_X1 U7435 ( .B1(FLUSH_REG_SCAN_IN), .B2(MORE_REG_SCAN_IN), .A(n6527), 
        .ZN(n6528) );
  NAND4_X1 U7436 ( .A1(n6531), .A2(n6530), .A3(n6529), .A4(n6528), .ZN(n6532)
         );
  AOI211_X1 U7437 ( .C1(n6535), .C2(n6534), .A(n6533), .B(n6532), .ZN(n6547)
         );
  INV_X1 U7438 ( .A(READY_N), .ZN(n6789) );
  AOI22_X1 U7439 ( .A1(n6547), .A2(n6537), .B1(READY_N), .B2(n6536), .ZN(n6538) );
  INV_X1 U7440 ( .A(n6538), .ZN(n6539) );
  OAI21_X1 U7441 ( .B1(n6541), .B2(n6540), .A(n6539), .ZN(n6614) );
  OAI21_X1 U7442 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6789), .A(n6614), .ZN(
        n6548) );
  AOI221_X1 U7443 ( .B1(n6543), .B2(STATE2_REG_0__SCAN_IN), .C1(n6548), .C2(
        STATE2_REG_0__SCAN_IN), .A(n6542), .ZN(n6546) );
  OAI211_X1 U7444 ( .C1(n6650), .C2(n6617), .A(n6544), .B(n6614), .ZN(n6545)
         );
  OAI211_X1 U7445 ( .C1(n6547), .C2(n6550), .A(n6546), .B(n6545), .ZN(U3148)
         );
  NAND3_X1 U7446 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6549), .A3(n6548), .ZN(
        n6555) );
  OAI21_X1 U7447 ( .B1(READY_N), .B2(n6551), .A(n6550), .ZN(n6553) );
  AOI21_X1 U7448 ( .B1(n6553), .B2(n6614), .A(n6552), .ZN(n6554) );
  NAND2_X1 U7449 ( .A1(n6555), .A2(n6554), .ZN(U3149) );
  OAI211_X1 U7450 ( .C1(STATE2_REG_2__SCAN_IN), .C2(n6789), .A(n6612), .B(
        n6650), .ZN(n6557) );
  OAI21_X1 U7451 ( .B1(n6558), .B2(n6557), .A(n6556), .ZN(U3150) );
  AND2_X1 U7452 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6608), .ZN(U3151) );
  AND2_X1 U7453 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6608), .ZN(U3152) );
  AND2_X1 U7454 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6608), .ZN(U3153) );
  AND2_X1 U7455 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6608), .ZN(U3154) );
  AND2_X1 U7456 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6608), .ZN(U3155) );
  AND2_X1 U7457 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6608), .ZN(U3156) );
  AND2_X1 U7458 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6608), .ZN(U3157) );
  AND2_X1 U7459 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6608), .ZN(U3158) );
  AND2_X1 U7460 ( .A1(n6608), .A2(DATAWIDTH_REG_23__SCAN_IN), .ZN(U3159) );
  INV_X1 U7461 ( .A(DATAWIDTH_REG_22__SCAN_IN), .ZN(n6768) );
  NOR2_X1 U7462 ( .A1(n6611), .A2(n6768), .ZN(U3160) );
  AND2_X1 U7463 ( .A1(n6608), .A2(DATAWIDTH_REG_21__SCAN_IN), .ZN(U3161) );
  INV_X1 U7464 ( .A(DATAWIDTH_REG_20__SCAN_IN), .ZN(n6971) );
  NOR2_X1 U7465 ( .A1(n6611), .A2(n6971), .ZN(U3162) );
  INV_X1 U7466 ( .A(DATAWIDTH_REG_19__SCAN_IN), .ZN(n6824) );
  NOR2_X1 U7467 ( .A1(n6611), .A2(n6824), .ZN(U3163) );
  INV_X1 U7468 ( .A(DATAWIDTH_REG_18__SCAN_IN), .ZN(n7005) );
  NOR2_X1 U7469 ( .A1(n6611), .A2(n7005), .ZN(U3164) );
  INV_X1 U7470 ( .A(DATAWIDTH_REG_17__SCAN_IN), .ZN(n6772) );
  NOR2_X1 U7471 ( .A1(n6611), .A2(n6772), .ZN(U3165) );
  INV_X1 U7472 ( .A(DATAWIDTH_REG_16__SCAN_IN), .ZN(n6774) );
  NOR2_X1 U7473 ( .A1(n6611), .A2(n6774), .ZN(U3166) );
  INV_X1 U7474 ( .A(DATAWIDTH_REG_15__SCAN_IN), .ZN(n7010) );
  NOR2_X1 U7475 ( .A1(n6611), .A2(n7010), .ZN(U3167) );
  INV_X1 U7476 ( .A(DATAWIDTH_REG_14__SCAN_IN), .ZN(n6800) );
  NOR2_X1 U7477 ( .A1(n6611), .A2(n6800), .ZN(U3168) );
  INV_X1 U7478 ( .A(DATAWIDTH_REG_13__SCAN_IN), .ZN(n6841) );
  NOR2_X1 U7479 ( .A1(n6611), .A2(n6841), .ZN(U3169) );
  INV_X1 U7480 ( .A(DATAWIDTH_REG_12__SCAN_IN), .ZN(n7027) );
  NOR2_X1 U7481 ( .A1(n6611), .A2(n7027), .ZN(U3170) );
  INV_X1 U7482 ( .A(DATAWIDTH_REG_11__SCAN_IN), .ZN(n6820) );
  NOR2_X1 U7483 ( .A1(n6611), .A2(n6820), .ZN(U3171) );
  INV_X1 U7484 ( .A(DATAWIDTH_REG_10__SCAN_IN), .ZN(n6857) );
  NOR2_X1 U7485 ( .A1(n6611), .A2(n6857), .ZN(U3172) );
  AND2_X1 U7486 ( .A1(n6608), .A2(DATAWIDTH_REG_9__SCAN_IN), .ZN(U3173) );
  INV_X1 U7487 ( .A(DATAWIDTH_REG_8__SCAN_IN), .ZN(n7007) );
  NOR2_X1 U7488 ( .A1(n6611), .A2(n7007), .ZN(U3174) );
  AND2_X1 U7489 ( .A1(n6608), .A2(DATAWIDTH_REG_7__SCAN_IN), .ZN(U3175) );
  INV_X1 U7490 ( .A(DATAWIDTH_REG_6__SCAN_IN), .ZN(n6980) );
  NOR2_X1 U7491 ( .A1(n6611), .A2(n6980), .ZN(U3176) );
  INV_X1 U7492 ( .A(DATAWIDTH_REG_5__SCAN_IN), .ZN(n6729) );
  NOR2_X1 U7493 ( .A1(n6611), .A2(n6729), .ZN(U3177) );
  INV_X1 U7494 ( .A(DATAWIDTH_REG_4__SCAN_IN), .ZN(n6996) );
  NOR2_X1 U7495 ( .A1(n6611), .A2(n6996), .ZN(U3178) );
  AND2_X1 U7496 ( .A1(n6608), .A2(DATAWIDTH_REG_3__SCAN_IN), .ZN(U3179) );
  INV_X1 U7497 ( .A(DATAWIDTH_REG_2__SCAN_IN), .ZN(n6735) );
  NOR2_X1 U7498 ( .A1(n6611), .A2(n6735), .ZN(U3180) );
  NAND2_X1 U7499 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n6562) );
  NAND2_X1 U7500 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n6567) );
  NAND2_X1 U7501 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .ZN(n6571) );
  NAND2_X1 U7502 ( .A1(n6567), .A2(n6571), .ZN(n6560) );
  INV_X1 U7503 ( .A(NA_N), .ZN(n6743) );
  INV_X1 U7504 ( .A(n6568), .ZN(n6559) );
  AOI211_X1 U7505 ( .C1(STATE_REG_2__SCAN_IN), .C2(n6743), .A(
        STATE_REG_0__SCAN_IN), .B(n6559), .ZN(n6575) );
  AOI21_X1 U7506 ( .B1(n6568), .B2(n6560), .A(n6575), .ZN(n6561) );
  OAI221_X1 U7507 ( .B1(n7048), .B2(REQUESTPENDING_REG_SCAN_IN), .C1(n7048), 
        .C2(n6562), .A(n6561), .ZN(U3181) );
  AND2_X1 U7508 ( .A1(STATE_REG_0__SCAN_IN), .A2(REQUESTPENDING_REG_SCAN_IN), 
        .ZN(n6564) );
  INV_X1 U7509 ( .A(n6562), .ZN(n6563) );
  OAI21_X1 U7510 ( .B1(n6564), .B2(n6563), .A(n6567), .ZN(n6565) );
  NAND3_X1 U7511 ( .A1(n6566), .A2(n6571), .A3(n6565), .ZN(U3182) );
  AOI221_X1 U7512 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n6789), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6570) );
  OAI211_X1 U7513 ( .C1(n6568), .C2(n6571), .A(STATE_REG_0__SCAN_IN), .B(n6567), .ZN(n6569) );
  AOI21_X1 U7514 ( .B1(HOLD), .B2(n6570), .A(n6569), .ZN(n6574) );
  INV_X1 U7515 ( .A(n6571), .ZN(n6572) );
  NAND4_X1 U7516 ( .A1(REQUESTPENDING_REG_SCAN_IN), .A2(STATE_REG_0__SCAN_IN), 
        .A3(n6572), .A4(n6743), .ZN(n6573) );
  OAI21_X1 U7517 ( .B1(n6575), .B2(n6574), .A(n6573), .ZN(U3183) );
  NAND2_X1 U7518 ( .A1(n7048), .A2(n6576), .ZN(n6598) );
  INV_X1 U7519 ( .A(ADDRESS_REG_0__SCAN_IN), .ZN(n6755) );
  OAI222_X1 U7520 ( .A1(n6598), .A2(n6578), .B1(n6755), .B2(n7048), .C1(n6577), 
        .C2(n6602), .ZN(U3184) );
  INV_X1 U7521 ( .A(ADDRESS_REG_1__SCAN_IN), .ZN(n6876) );
  INV_X1 U7522 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6580) );
  OAI222_X1 U7523 ( .A1(n6602), .A2(n6578), .B1(n6876), .B2(n7048), .C1(n6580), 
        .C2(n6606), .ZN(U3185) );
  INV_X1 U7524 ( .A(ADDRESS_REG_2__SCAN_IN), .ZN(n6579) );
  OAI222_X1 U7525 ( .A1(n6602), .A2(n6580), .B1(n6579), .B2(n7048), .C1(n6581), 
        .C2(n6606), .ZN(U3186) );
  INV_X1 U7526 ( .A(ADDRESS_REG_3__SCAN_IN), .ZN(n6861) );
  OAI222_X1 U7527 ( .A1(n6602), .A2(n6581), .B1(n6861), .B2(n7048), .C1(n6582), 
        .C2(n6598), .ZN(U3187) );
  INV_X1 U7528 ( .A(ADDRESS_REG_4__SCAN_IN), .ZN(n6855) );
  OAI222_X1 U7529 ( .A1(n6602), .A2(n6582), .B1(n6855), .B2(n7048), .C1(n6583), 
        .C2(n6606), .ZN(U3188) );
  INV_X1 U7530 ( .A(ADDRESS_REG_5__SCAN_IN), .ZN(n6813) );
  OAI222_X1 U7531 ( .A1(n6602), .A2(n6583), .B1(n6813), .B2(n7048), .C1(n6584), 
        .C2(n6606), .ZN(U3189) );
  INV_X1 U7532 ( .A(ADDRESS_REG_6__SCAN_IN), .ZN(n6860) );
  OAI222_X1 U7533 ( .A1(n6602), .A2(n6584), .B1(n6860), .B2(n7048), .C1(n6586), 
        .C2(n6598), .ZN(U3190) );
  INV_X1 U7534 ( .A(ADDRESS_REG_7__SCAN_IN), .ZN(n6585) );
  OAI222_X1 U7535 ( .A1(n6602), .A2(n6586), .B1(n6585), .B2(n7048), .C1(n6587), 
        .C2(n6606), .ZN(U3191) );
  INV_X1 U7536 ( .A(ADDRESS_REG_8__SCAN_IN), .ZN(n6588) );
  OAI222_X1 U7537 ( .A1(n6598), .A2(n6589), .B1(n6588), .B2(n7048), .C1(n6587), 
        .C2(n6602), .ZN(U3192) );
  INV_X1 U7538 ( .A(ADDRESS_REG_9__SCAN_IN), .ZN(n6867) );
  INV_X1 U7539 ( .A(REIP_REG_11__SCAN_IN), .ZN(n6590) );
  OAI222_X1 U7540 ( .A1(n6602), .A2(n6589), .B1(n6867), .B2(n7048), .C1(n6590), 
        .C2(n6598), .ZN(U3193) );
  INV_X1 U7541 ( .A(ADDRESS_REG_10__SCAN_IN), .ZN(n6873) );
  OAI222_X1 U7542 ( .A1(n6606), .A2(n6592), .B1(n6873), .B2(n7048), .C1(n6590), 
        .C2(n6602), .ZN(U3194) );
  INV_X1 U7543 ( .A(ADDRESS_REG_11__SCAN_IN), .ZN(n6591) );
  INV_X1 U7544 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6594) );
  OAI222_X1 U7545 ( .A1(n6602), .A2(n6592), .B1(n6591), .B2(n7048), .C1(n6594), 
        .C2(n6598), .ZN(U3195) );
  INV_X1 U7546 ( .A(ADDRESS_REG_12__SCAN_IN), .ZN(n6593) );
  OAI222_X1 U7547 ( .A1(n6602), .A2(n6594), .B1(n6593), .B2(n7048), .C1(n6595), 
        .C2(n6598), .ZN(U3196) );
  INV_X1 U7548 ( .A(ADDRESS_REG_13__SCAN_IN), .ZN(n6731) );
  OAI222_X1 U7549 ( .A1(n6602), .A2(n6595), .B1(n6731), .B2(n7048), .C1(n6596), 
        .C2(n6598), .ZN(U3197) );
  INV_X1 U7550 ( .A(ADDRESS_REG_14__SCAN_IN), .ZN(n6761) );
  OAI222_X1 U7551 ( .A1(n6598), .A2(n6746), .B1(n6761), .B2(n7048), .C1(n6596), 
        .C2(n6602), .ZN(U3198) );
  INV_X1 U7552 ( .A(ADDRESS_REG_15__SCAN_IN), .ZN(n7020) );
  INV_X1 U7553 ( .A(REIP_REG_17__SCAN_IN), .ZN(n6597) );
  OAI222_X1 U7554 ( .A1(n6602), .A2(n6746), .B1(n7020), .B2(n7048), .C1(n6597), 
        .C2(n6606), .ZN(U3199) );
  INV_X1 U7555 ( .A(ADDRESS_REG_16__SCAN_IN), .ZN(n6808) );
  OAI222_X1 U7556 ( .A1(n6598), .A2(n6854), .B1(n6808), .B2(n7048), .C1(n6597), 
        .C2(n6602), .ZN(U3200) );
  INV_X1 U7557 ( .A(ADDRESS_REG_17__SCAN_IN), .ZN(n6823) );
  INV_X1 U7558 ( .A(REIP_REG_19__SCAN_IN), .ZN(n6599) );
  OAI222_X1 U7559 ( .A1(n6602), .A2(n6854), .B1(n6823), .B2(n7048), .C1(n6599), 
        .C2(n6606), .ZN(U3201) );
  INV_X1 U7560 ( .A(ADDRESS_REG_18__SCAN_IN), .ZN(n6788) );
  OAI222_X1 U7561 ( .A1(n6602), .A2(n6599), .B1(n6788), .B2(n7048), .C1(n6600), 
        .C2(n6606), .ZN(U3202) );
  INV_X1 U7562 ( .A(ADDRESS_REG_19__SCAN_IN), .ZN(n6995) );
  OAI222_X1 U7563 ( .A1(n6602), .A2(n6600), .B1(n6995), .B2(n7048), .C1(n6972), 
        .C2(n6606), .ZN(U3203) );
  INV_X1 U7564 ( .A(ADDRESS_REG_20__SCAN_IN), .ZN(n6758) );
  OAI222_X1 U7565 ( .A1(n6602), .A2(n6972), .B1(n6758), .B2(n7048), .C1(n6871), 
        .C2(n6606), .ZN(U3204) );
  INV_X1 U7566 ( .A(ADDRESS_REG_21__SCAN_IN), .ZN(n6770) );
  OAI222_X1 U7567 ( .A1(n6602), .A2(n6871), .B1(n6770), .B2(n7048), .C1(n6842), 
        .C2(n6606), .ZN(U3205) );
  INV_X1 U7568 ( .A(ADDRESS_REG_22__SCAN_IN), .ZN(n6760) );
  OAI222_X1 U7569 ( .A1(n6602), .A2(n6842), .B1(n6760), .B2(n7048), .C1(n6791), 
        .C2(n6606), .ZN(U3206) );
  INV_X1 U7570 ( .A(ADDRESS_REG_23__SCAN_IN), .ZN(n6775) );
  OAI222_X1 U7571 ( .A1(n6606), .A2(n5444), .B1(n6775), .B2(n7048), .C1(n6791), 
        .C2(n6602), .ZN(U3207) );
  INV_X1 U7572 ( .A(ADDRESS_REG_24__SCAN_IN), .ZN(n6601) );
  OAI222_X1 U7573 ( .A1(n6602), .A2(n5444), .B1(n6601), .B2(n7048), .C1(n5515), 
        .C2(n6606), .ZN(U3208) );
  INV_X1 U7574 ( .A(ADDRESS_REG_25__SCAN_IN), .ZN(n6754) );
  OAI222_X1 U7575 ( .A1(n6602), .A2(n5515), .B1(n6754), .B2(n7048), .C1(n6875), 
        .C2(n6606), .ZN(U3209) );
  INV_X1 U7576 ( .A(ADDRESS_REG_26__SCAN_IN), .ZN(n6603) );
  OAI222_X1 U7577 ( .A1(n6602), .A2(n6875), .B1(n6603), .B2(n7048), .C1(n6741), 
        .C2(n6606), .ZN(U3210) );
  INV_X1 U7578 ( .A(ADDRESS_REG_27__SCAN_IN), .ZN(n6604) );
  OAI222_X1 U7579 ( .A1(n6602), .A2(n6741), .B1(n6604), .B2(n7048), .C1(n6811), 
        .C2(n6606), .ZN(U3211) );
  INV_X1 U7580 ( .A(ADDRESS_REG_28__SCAN_IN), .ZN(n6889) );
  OAI222_X1 U7581 ( .A1(n6602), .A2(n6811), .B1(n6889), .B2(n7048), .C1(n5415), 
        .C2(n6606), .ZN(U3212) );
  INV_X1 U7582 ( .A(REIP_REG_31__SCAN_IN), .ZN(n6605) );
  INV_X1 U7583 ( .A(ADDRESS_REG_29__SCAN_IN), .ZN(n6884) );
  OAI222_X1 U7584 ( .A1(n6606), .A2(n6605), .B1(n6884), .B2(n7048), .C1(n5415), 
        .C2(n6602), .ZN(U3213) );
  INV_X1 U7585 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6844) );
  INV_X1 U7586 ( .A(BE_N_REG_2__SCAN_IN), .ZN(n6986) );
  AOI22_X1 U7587 ( .A1(n7048), .A2(n6844), .B1(n6986), .B2(n7047), .ZN(U3446)
         );
  INV_X1 U7588 ( .A(BE_N_REG_1__SCAN_IN), .ZN(n6890) );
  AOI22_X1 U7589 ( .A1(n7048), .A2(n6992), .B1(n6890), .B2(n7047), .ZN(U3447)
         );
  INV_X1 U7590 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6798) );
  INV_X1 U7591 ( .A(BE_N_REG_0__SCAN_IN), .ZN(n6975) );
  AOI22_X1 U7592 ( .A1(n7048), .A2(n6798), .B1(n6975), .B2(n7047), .ZN(U3448)
         );
  INV_X1 U7593 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6636) );
  INV_X1 U7594 ( .A(n6609), .ZN(n6607) );
  AOI21_X1 U7595 ( .B1(n6636), .B2(n6608), .A(n6607), .ZN(U3451) );
  INV_X1 U7596 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6610) );
  OAI21_X1 U7597 ( .B1(n6611), .B2(n6610), .A(n6609), .ZN(U3452) );
  OAI211_X1 U7598 ( .C1(n6615), .C2(n6614), .A(n6613), .B(n6612), .ZN(U3453)
         );
  OAI22_X1 U7599 ( .A1(n6618), .A2(n6634), .B1(n6617), .B2(n6616), .ZN(n6619)
         );
  MUX2_X1 U7600 ( .A(n6619), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n6631), 
        .Z(U3456) );
  AOI21_X1 U7601 ( .B1(n6622), .B2(n6621), .A(n6620), .ZN(n6628) );
  NOR3_X1 U7602 ( .A1(n6624), .A2(n6623), .A3(STATE2_REG_3__SCAN_IN), .ZN(
        n6625) );
  NOR2_X1 U7603 ( .A1(n6625), .A2(STATE2_REG_1__SCAN_IN), .ZN(n6626) );
  OAI22_X1 U7604 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n6628), .B1(n6627), .B2(n6626), .ZN(n6630) );
  AOI22_X1 U7605 ( .A1(n6631), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(n6630), .B2(n6629), .ZN(n6632) );
  OAI21_X1 U7606 ( .B1(n6634), .B2(n6633), .A(n6632), .ZN(U3461) );
  NOR3_X1 U7607 ( .A1(n6636), .A2(REIP_REG_0__SCAN_IN), .A3(
        REIP_REG_1__SCAN_IN), .ZN(n6635) );
  AOI221_X1 U7608 ( .B1(n6637), .B2(n6636), .C1(REIP_REG_1__SCAN_IN), .C2(
        REIP_REG_0__SCAN_IN), .A(n6635), .ZN(n6638) );
  INV_X1 U7609 ( .A(n6641), .ZN(n6639) );
  AOI22_X1 U7610 ( .A1(n6641), .A2(n6638), .B1(n6844), .B2(n6639), .ZN(U3468)
         );
  NOR2_X1 U7611 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .ZN(
        n6640) );
  AOI22_X1 U7612 ( .A1(n6641), .A2(n6640), .B1(n6798), .B2(n6639), .ZN(U3469)
         );
  INV_X1 U7613 ( .A(W_R_N_REG_SCAN_IN), .ZN(n6642) );
  AOI22_X1 U7614 ( .A1(n7048), .A2(READREQUEST_REG_SCAN_IN), .B1(n6642), .B2(
        n7047), .ZN(U3470) );
  OAI211_X1 U7615 ( .C1(READY_N), .C2(n6645), .A(n6644), .B(n6643), .ZN(n6646)
         );
  NOR2_X1 U7616 ( .A1(n6647), .A2(n6646), .ZN(n6655) );
  OAI211_X1 U7617 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n6649), .A(n6648), .B(
        STATE2_REG_2__SCAN_IN), .ZN(n6652) );
  INV_X1 U7618 ( .A(n6650), .ZN(n6651) );
  AOI21_X1 U7619 ( .B1(n6652), .B2(STATE2_REG_0__SCAN_IN), .A(n6651), .ZN(
        n6654) );
  NAND2_X1 U7620 ( .A1(n6655), .A2(REQUESTPENDING_REG_SCAN_IN), .ZN(n6653) );
  OAI21_X1 U7621 ( .B1(n6655), .B2(n6654), .A(n6653), .ZN(U3472) );
  INV_X1 U7622 ( .A(M_IO_N_REG_SCAN_IN), .ZN(n7026) );
  AOI22_X1 U7623 ( .A1(n7048), .A2(n6656), .B1(n7026), .B2(n7047), .ZN(U3473)
         );
  XOR2_X1 U7624 ( .A(ADDRESS_REG_29__SCAN_IN), .B(keyinput_g71), .Z(n6663) );
  AOI22_X1 U7625 ( .A1(ADDRESS_REG_26__SCAN_IN), .A2(keyinput_g74), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(keyinput_g88), .ZN(n6657) );
  OAI221_X1 U7626 ( .B1(ADDRESS_REG_26__SCAN_IN), .B2(keyinput_g74), .C1(
        ADDRESS_REG_12__SCAN_IN), .C2(keyinput_g88), .A(n6657), .ZN(n6662) );
  AOI22_X1 U7627 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(keyinput_g108), .B1(HOLD), .B2(keyinput_g36), .ZN(n6658) );
  OAI221_X1 U7628 ( .B1(DATAWIDTH_REG_4__SCAN_IN), .B2(keyinput_g108), .C1(
        HOLD), .C2(keyinput_g36), .A(n6658), .ZN(n6661) );
  AOI22_X1 U7629 ( .A1(BE_N_REG_1__SCAN_IN), .A2(keyinput_g69), .B1(
        REIP_REG_25__SCAN_IN), .B2(keyinput_g57), .ZN(n6659) );
  OAI221_X1 U7630 ( .B1(BE_N_REG_1__SCAN_IN), .B2(keyinput_g69), .C1(
        REIP_REG_25__SCAN_IN), .C2(keyinput_g57), .A(n6659), .ZN(n6660) );
  NOR4_X1 U7631 ( .A1(n6663), .A2(n6662), .A3(n6661), .A4(n6660), .ZN(n6691)
         );
  AOI22_X1 U7632 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(keyinput_g107), .B1(
        DATAI_11_), .B2(keyinput_g20), .ZN(n6664) );
  OAI221_X1 U7633 ( .B1(DATAWIDTH_REG_3__SCAN_IN), .B2(keyinput_g107), .C1(
        DATAI_11_), .C2(keyinput_g20), .A(n6664), .ZN(n6671) );
  AOI22_X1 U7634 ( .A1(FLUSH_REG_SCAN_IN), .A2(keyinput_g45), .B1(DATAI_23_), 
        .B2(keyinput_g8), .ZN(n6665) );
  OAI221_X1 U7635 ( .B1(FLUSH_REG_SCAN_IN), .B2(keyinput_g45), .C1(DATAI_23_), 
        .C2(keyinput_g8), .A(n6665), .ZN(n6670) );
  AOI22_X1 U7636 ( .A1(W_R_N_REG_SCAN_IN), .A2(keyinput_g46), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(keyinput_g93), .ZN(n6666) );
  OAI221_X1 U7637 ( .B1(W_R_N_REG_SCAN_IN), .B2(keyinput_g46), .C1(
        ADDRESS_REG_7__SCAN_IN), .C2(keyinput_g93), .A(n6666), .ZN(n6669) );
  AOI22_X1 U7638 ( .A1(DATAI_5_), .A2(keyinput_g26), .B1(DATAI_8_), .B2(
        keyinput_g23), .ZN(n6667) );
  OAI221_X1 U7639 ( .B1(DATAI_5_), .B2(keyinput_g26), .C1(DATAI_8_), .C2(
        keyinput_g23), .A(n6667), .ZN(n6668) );
  NOR4_X1 U7640 ( .A1(n6671), .A2(n6670), .A3(n6669), .A4(n6668), .ZN(n6690)
         );
  AOI22_X1 U7641 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(keyinput_g127), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(keyinput_g98), .ZN(n6672) );
  OAI221_X1 U7642 ( .B1(DATAWIDTH_REG_23__SCAN_IN), .B2(keyinput_g127), .C1(
        ADDRESS_REG_2__SCAN_IN), .C2(keyinput_g98), .A(n6672), .ZN(n6679) );
  AOI22_X1 U7643 ( .A1(REQUESTPENDING_REG_SCAN_IN), .A2(keyinput_g42), .B1(
        REIP_REG_19__SCAN_IN), .B2(keyinput_g63), .ZN(n6673) );
  OAI221_X1 U7644 ( .B1(REQUESTPENDING_REG_SCAN_IN), .B2(keyinput_g42), .C1(
        REIP_REG_19__SCAN_IN), .C2(keyinput_g63), .A(n6673), .ZN(n6678) );
  AOI22_X1 U7645 ( .A1(DATAI_15_), .A2(keyinput_g16), .B1(REIP_REG_22__SCAN_IN), .B2(keyinput_g60), .ZN(n6674) );
  OAI221_X1 U7646 ( .B1(DATAI_15_), .B2(keyinput_g16), .C1(
        REIP_REG_22__SCAN_IN), .C2(keyinput_g60), .A(n6674), .ZN(n6677) );
  AOI22_X1 U7647 ( .A1(MEMORYFETCH_REG_SCAN_IN), .A2(keyinput_g32), .B1(
        REIP_REG_17__SCAN_IN), .B2(keyinput_g65), .ZN(n6675) );
  OAI221_X1 U7648 ( .B1(MEMORYFETCH_REG_SCAN_IN), .B2(keyinput_g32), .C1(
        REIP_REG_17__SCAN_IN), .C2(keyinput_g65), .A(n6675), .ZN(n6676) );
  NOR4_X1 U7649 ( .A1(n6679), .A2(n6678), .A3(n6677), .A4(n6676), .ZN(n6689)
         );
  AOI22_X1 U7650 ( .A1(BE_N_REG_2__SCAN_IN), .A2(keyinput_g68), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(keyinput_g73), .ZN(n6680) );
  OAI221_X1 U7651 ( .B1(BE_N_REG_2__SCAN_IN), .B2(keyinput_g68), .C1(
        ADDRESS_REG_27__SCAN_IN), .C2(keyinput_g73), .A(n6680), .ZN(n6687) );
  AOI22_X1 U7652 ( .A1(DATAI_24_), .A2(keyinput_g7), .B1(REIP_REG_21__SCAN_IN), 
        .B2(keyinput_g61), .ZN(n6681) );
  OAI221_X1 U7653 ( .B1(DATAI_24_), .B2(keyinput_g7), .C1(REIP_REG_21__SCAN_IN), .C2(keyinput_g61), .A(n6681), .ZN(n6686) );
  AOI22_X1 U7654 ( .A1(ADDRESS_REG_24__SCAN_IN), .A2(keyinput_g76), .B1(
        REIP_REG_27__SCAN_IN), .B2(keyinput_g55), .ZN(n6682) );
  OAI221_X1 U7655 ( .B1(ADDRESS_REG_24__SCAN_IN), .B2(keyinput_g76), .C1(
        REIP_REG_27__SCAN_IN), .C2(keyinput_g55), .A(n6682), .ZN(n6685) );
  AOI22_X1 U7656 ( .A1(DATAWIDTH_REG_0__SCAN_IN), .A2(keyinput_g104), .B1(
        DATAWIDTH_REG_9__SCAN_IN), .B2(keyinput_g113), .ZN(n6683) );
  OAI221_X1 U7657 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(keyinput_g104), .C1(
        DATAWIDTH_REG_9__SCAN_IN), .C2(keyinput_g113), .A(n6683), .ZN(n6684)
         );
  NOR4_X1 U7658 ( .A1(n6687), .A2(n6686), .A3(n6685), .A4(n6684), .ZN(n6688)
         );
  NAND4_X1 U7659 ( .A1(n6691), .A2(n6690), .A3(n6689), .A4(n6688), .ZN(n6836)
         );
  AOI22_X1 U7660 ( .A1(ADDRESS_REG_15__SCAN_IN), .A2(keyinput_g85), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(keyinput_g89), .ZN(n6692) );
  OAI221_X1 U7661 ( .B1(ADDRESS_REG_15__SCAN_IN), .B2(keyinput_g85), .C1(
        ADDRESS_REG_11__SCAN_IN), .C2(keyinput_g89), .A(n6692), .ZN(n6699) );
  AOI22_X1 U7662 ( .A1(DATAI_25_), .A2(keyinput_g6), .B1(DATAI_29_), .B2(
        keyinput_g2), .ZN(n6693) );
  OAI221_X1 U7663 ( .B1(DATAI_25_), .B2(keyinput_g6), .C1(DATAI_29_), .C2(
        keyinput_g2), .A(n6693), .ZN(n6698) );
  AOI22_X1 U7664 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(keyinput_g111), .B1(
        DATAI_7_), .B2(keyinput_g24), .ZN(n6694) );
  OAI221_X1 U7665 ( .B1(DATAWIDTH_REG_7__SCAN_IN), .B2(keyinput_g111), .C1(
        DATAI_7_), .C2(keyinput_g24), .A(n6694), .ZN(n6697) );
  AOI22_X1 U7666 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(keyinput_g112), .B1(
        BYTEENABLE_REG_1__SCAN_IN), .B2(keyinput_g48), .ZN(n6695) );
  OAI221_X1 U7667 ( .B1(DATAWIDTH_REG_8__SCAN_IN), .B2(keyinput_g112), .C1(
        BYTEENABLE_REG_1__SCAN_IN), .C2(keyinput_g48), .A(n6695), .ZN(n6696)
         );
  NOR4_X1 U7668 ( .A1(n6699), .A2(n6698), .A3(n6697), .A4(n6696), .ZN(n6727)
         );
  AOI22_X1 U7669 ( .A1(DATAI_18_), .A2(keyinput_g13), .B1(DATAI_12_), .B2(
        keyinput_g19), .ZN(n6700) );
  OAI221_X1 U7670 ( .B1(DATAI_18_), .B2(keyinput_g13), .C1(DATAI_12_), .C2(
        keyinput_g19), .A(n6700), .ZN(n6707) );
  AOI22_X1 U7671 ( .A1(ADDRESS_REG_28__SCAN_IN), .A2(keyinput_g72), .B1(BS16_N), .B2(keyinput_g34), .ZN(n6701) );
  OAI221_X1 U7672 ( .B1(ADDRESS_REG_28__SCAN_IN), .B2(keyinput_g72), .C1(
        BS16_N), .C2(keyinput_g34), .A(n6701), .ZN(n6706) );
  AOI22_X1 U7673 ( .A1(DATAI_22_), .A2(keyinput_g9), .B1(DATAI_14_), .B2(
        keyinput_g17), .ZN(n6702) );
  OAI221_X1 U7674 ( .B1(DATAI_22_), .B2(keyinput_g9), .C1(DATAI_14_), .C2(
        keyinput_g17), .A(n6702), .ZN(n6705) );
  AOI22_X1 U7675 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(keyinput_g116), .B1(
        STATE_REG_2__SCAN_IN), .B2(keyinput_g101), .ZN(n6703) );
  OAI221_X1 U7676 ( .B1(DATAWIDTH_REG_12__SCAN_IN), .B2(keyinput_g116), .C1(
        STATE_REG_2__SCAN_IN), .C2(keyinput_g101), .A(n6703), .ZN(n6704) );
  NOR4_X1 U7677 ( .A1(n6707), .A2(n6706), .A3(n6705), .A4(n6704), .ZN(n6726)
         );
  AOI22_X1 U7678 ( .A1(DATAWIDTH_REG_1__SCAN_IN), .A2(keyinput_g105), .B1(
        REIP_REG_20__SCAN_IN), .B2(keyinput_g62), .ZN(n6708) );
  OAI221_X1 U7679 ( .B1(DATAWIDTH_REG_1__SCAN_IN), .B2(keyinput_g105), .C1(
        REIP_REG_20__SCAN_IN), .C2(keyinput_g62), .A(n6708), .ZN(n6715) );
  AOI22_X1 U7680 ( .A1(DATAI_20_), .A2(keyinput_g11), .B1(REIP_REG_26__SCAN_IN), .B2(keyinput_g56), .ZN(n6709) );
  OAI221_X1 U7681 ( .B1(DATAI_20_), .B2(keyinput_g11), .C1(
        REIP_REG_26__SCAN_IN), .C2(keyinput_g56), .A(n6709), .ZN(n6714) );
  AOI22_X1 U7682 ( .A1(REIP_REG_18__SCAN_IN), .A2(keyinput_g64), .B1(DATAI_31_), .B2(keyinput_g0), .ZN(n6710) );
  OAI221_X1 U7683 ( .B1(REIP_REG_18__SCAN_IN), .B2(keyinput_g64), .C1(
        DATAI_31_), .C2(keyinput_g0), .A(n6710), .ZN(n6713) );
  AOI22_X1 U7684 ( .A1(REIP_REG_31__SCAN_IN), .A2(keyinput_g51), .B1(
        STATE_REG_1__SCAN_IN), .B2(keyinput_g102), .ZN(n6711) );
  OAI221_X1 U7685 ( .B1(REIP_REG_31__SCAN_IN), .B2(keyinput_g51), .C1(
        STATE_REG_1__SCAN_IN), .C2(keyinput_g102), .A(n6711), .ZN(n6712) );
  NOR4_X1 U7686 ( .A1(n6715), .A2(n6714), .A3(n6713), .A4(n6712), .ZN(n6725)
         );
  AOI22_X1 U7687 ( .A1(DATAI_2_), .A2(keyinput_g29), .B1(DATAI_19_), .B2(
        keyinput_g12), .ZN(n6716) );
  OAI221_X1 U7688 ( .B1(DATAI_2_), .B2(keyinput_g29), .C1(DATAI_19_), .C2(
        keyinput_g12), .A(n6716), .ZN(n6723) );
  AOI22_X1 U7689 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(keyinput_g114), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(keyinput_g92), .ZN(n6717) );
  OAI221_X1 U7690 ( .B1(DATAWIDTH_REG_10__SCAN_IN), .B2(keyinput_g114), .C1(
        ADDRESS_REG_8__SCAN_IN), .C2(keyinput_g92), .A(n6717), .ZN(n6722) );
  AOI22_X1 U7691 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(keyinput_g110), .B1(
        REIP_REG_30__SCAN_IN), .B2(keyinput_g52), .ZN(n6718) );
  OAI221_X1 U7692 ( .B1(DATAWIDTH_REG_6__SCAN_IN), .B2(keyinput_g110), .C1(
        REIP_REG_30__SCAN_IN), .C2(keyinput_g52), .A(n6718), .ZN(n6721) );
  AOI22_X1 U7693 ( .A1(READREQUEST_REG_SCAN_IN), .A2(keyinput_g37), .B1(n7005), 
        .B2(keyinput_g122), .ZN(n6719) );
  OAI221_X1 U7694 ( .B1(READREQUEST_REG_SCAN_IN), .B2(keyinput_g37), .C1(n7005), .C2(keyinput_g122), .A(n6719), .ZN(n6720) );
  NOR4_X1 U7695 ( .A1(n6723), .A2(n6722), .A3(n6721), .A4(n6720), .ZN(n6724)
         );
  NAND4_X1 U7696 ( .A1(n6727), .A2(n6726), .A3(n6725), .A4(n6724), .ZN(n6835)
         );
  AOI22_X1 U7697 ( .A1(n6839), .A2(keyinput_g30), .B1(keyinput_g109), .B2(
        n6729), .ZN(n6728) );
  OAI221_X1 U7698 ( .B1(n6839), .B2(keyinput_g30), .C1(n6729), .C2(
        keyinput_g109), .A(n6728), .ZN(n6739) );
  INV_X1 U7699 ( .A(DATAI_9_), .ZN(n6732) );
  AOI22_X1 U7700 ( .A1(n6732), .A2(keyinput_g22), .B1(keyinput_g87), .B2(n6731), .ZN(n6730) );
  OAI221_X1 U7701 ( .B1(n6732), .B2(keyinput_g22), .C1(n6731), .C2(
        keyinput_g87), .A(n6730), .ZN(n6738) );
  AOI22_X1 U7702 ( .A1(n6855), .A2(keyinput_g96), .B1(keyinput_g81), .B2(n6995), .ZN(n6733) );
  OAI221_X1 U7703 ( .B1(n6855), .B2(keyinput_g96), .C1(n6995), .C2(
        keyinput_g81), .A(n6733), .ZN(n6737) );
  AOI22_X1 U7704 ( .A1(n6735), .A2(keyinput_g106), .B1(keyinput_g117), .B2(
        n6841), .ZN(n6734) );
  OAI221_X1 U7705 ( .B1(n6735), .B2(keyinput_g106), .C1(n6841), .C2(
        keyinput_g117), .A(n6734), .ZN(n6736) );
  NOR4_X1 U7706 ( .A1(n6739), .A2(n6738), .A3(n6737), .A4(n6736), .ZN(n6783)
         );
  AOI22_X1 U7707 ( .A1(n6741), .A2(keyinput_g54), .B1(keyinput_g97), .B2(n6861), .ZN(n6740) );
  OAI221_X1 U7708 ( .B1(n6741), .B2(keyinput_g54), .C1(n6861), .C2(
        keyinput_g97), .A(n6740), .ZN(n6752) );
  INV_X1 U7709 ( .A(BE_N_REG_3__SCAN_IN), .ZN(n6744) );
  AOI22_X1 U7710 ( .A1(n6744), .A2(keyinput_g67), .B1(keyinput_g33), .B2(n6743), .ZN(n6742) );
  OAI221_X1 U7711 ( .B1(n6744), .B2(keyinput_g67), .C1(n6743), .C2(
        keyinput_g33), .A(n6742), .ZN(n6751) );
  INV_X1 U7712 ( .A(DATAI_28_), .ZN(n6747) );
  AOI22_X1 U7713 ( .A1(n6747), .A2(keyinput_g3), .B1(n6746), .B2(keyinput_g66), 
        .ZN(n6745) );
  OAI221_X1 U7714 ( .B1(n6747), .B2(keyinput_g3), .C1(n6746), .C2(keyinput_g66), .A(n6745), .ZN(n6750) );
  INV_X1 U7715 ( .A(DATAI_21_), .ZN(n6882) );
  AOI22_X1 U7716 ( .A1(n6882), .A2(keyinput_g10), .B1(n6852), .B2(keyinput_g43), .ZN(n6748) );
  OAI221_X1 U7717 ( .B1(n6882), .B2(keyinput_g10), .C1(n6852), .C2(
        keyinput_g43), .A(n6748), .ZN(n6749) );
  NOR4_X1 U7718 ( .A1(n6752), .A2(n6751), .A3(n6750), .A4(n6749), .ZN(n6782)
         );
  AOI22_X1 U7719 ( .A1(n6755), .A2(keyinput_g100), .B1(keyinput_g75), .B2(
        n6754), .ZN(n6753) );
  OAI221_X1 U7720 ( .B1(n6755), .B2(keyinput_g100), .C1(n6754), .C2(
        keyinput_g75), .A(n6753), .ZN(n6765) );
  INV_X1 U7721 ( .A(DATAI_30_), .ZN(n7002) );
  AOI22_X1 U7722 ( .A1(n7002), .A2(keyinput_g1), .B1(keyinput_g27), .B2(n6978), 
        .ZN(n6756) );
  OAI221_X1 U7723 ( .B1(n7002), .B2(keyinput_g1), .C1(n6978), .C2(keyinput_g27), .A(n6756), .ZN(n6764) );
  AOI22_X1 U7724 ( .A1(n6758), .A2(keyinput_g80), .B1(keyinput_g41), .B2(n7018), .ZN(n6757) );
  OAI221_X1 U7725 ( .B1(n6758), .B2(keyinput_g80), .C1(n7018), .C2(
        keyinput_g41), .A(n6757), .ZN(n6763) );
  AOI22_X1 U7726 ( .A1(n6761), .A2(keyinput_g86), .B1(keyinput_g78), .B2(n6760), .ZN(n6759) );
  OAI221_X1 U7727 ( .B1(n6761), .B2(keyinput_g86), .C1(n6760), .C2(
        keyinput_g78), .A(n6759), .ZN(n6762) );
  NOR4_X1 U7728 ( .A1(n6765), .A2(n6764), .A3(n6763), .A4(n6762), .ZN(n6781)
         );
  INV_X1 U7729 ( .A(DATAI_27_), .ZN(n6767) );
  AOI22_X1 U7730 ( .A1(n6768), .A2(keyinput_g126), .B1(n6767), .B2(keyinput_g4), .ZN(n6766) );
  OAI221_X1 U7731 ( .B1(n6768), .B2(keyinput_g126), .C1(n6767), .C2(
        keyinput_g4), .A(n6766), .ZN(n6779) );
  AOI22_X1 U7732 ( .A1(n6770), .A2(keyinput_g79), .B1(keyinput_g124), .B2(
        n6971), .ZN(n6769) );
  OAI221_X1 U7733 ( .B1(n6770), .B2(keyinput_g79), .C1(n6971), .C2(
        keyinput_g124), .A(n6769), .ZN(n6778) );
  AOI22_X1 U7734 ( .A1(n6772), .A2(keyinput_g121), .B1(keyinput_g91), .B2(
        n6867), .ZN(n6771) );
  OAI221_X1 U7735 ( .B1(n6772), .B2(keyinput_g121), .C1(n6867), .C2(
        keyinput_g91), .A(n6771), .ZN(n6777) );
  AOI22_X1 U7736 ( .A1(n6775), .A2(keyinput_g77), .B1(keyinput_g120), .B2(
        n6774), .ZN(n6773) );
  OAI221_X1 U7737 ( .B1(n6775), .B2(keyinput_g77), .C1(n6774), .C2(
        keyinput_g120), .A(n6773), .ZN(n6776) );
  NOR4_X1 U7738 ( .A1(n6779), .A2(n6778), .A3(n6777), .A4(n6776), .ZN(n6780)
         );
  NAND4_X1 U7739 ( .A1(n6783), .A2(n6782), .A3(n6781), .A4(n6780), .ZN(n6834)
         );
  INV_X1 U7740 ( .A(DATAI_17_), .ZN(n6851) );
  AOI22_X1 U7741 ( .A1(n6851), .A2(keyinput_g14), .B1(n6785), .B2(
        keyinput_g103), .ZN(n6784) );
  OAI221_X1 U7742 ( .B1(n6851), .B2(keyinput_g14), .C1(n6785), .C2(
        keyinput_g103), .A(n6784), .ZN(n6795) );
  AOI22_X1 U7743 ( .A1(n7023), .A2(keyinput_g31), .B1(keyinput_g99), .B2(n6876), .ZN(n6786) );
  OAI221_X1 U7744 ( .B1(n7023), .B2(keyinput_g31), .C1(n6876), .C2(
        keyinput_g99), .A(n6786), .ZN(n6794) );
  AOI22_X1 U7745 ( .A1(n6789), .A2(keyinput_g35), .B1(keyinput_g82), .B2(n6788), .ZN(n6787) );
  OAI221_X1 U7746 ( .B1(n6789), .B2(keyinput_g35), .C1(n6788), .C2(
        keyinput_g82), .A(n6787), .ZN(n6793) );
  INV_X1 U7747 ( .A(DATAI_16_), .ZN(n6887) );
  AOI22_X1 U7748 ( .A1(n6887), .A2(keyinput_g15), .B1(n6791), .B2(keyinput_g58), .ZN(n6790) );
  OAI221_X1 U7749 ( .B1(n6887), .B2(keyinput_g15), .C1(n6791), .C2(
        keyinput_g58), .A(n6790), .ZN(n6792) );
  NOR4_X1 U7750 ( .A1(n6795), .A2(n6794), .A3(n6793), .A4(n6792), .ZN(n6832)
         );
  INV_X1 U7751 ( .A(DATAI_13_), .ZN(n6845) );
  INV_X1 U7752 ( .A(MORE_REG_SCAN_IN), .ZN(n6858) );
  AOI22_X1 U7753 ( .A1(n6845), .A2(keyinput_g18), .B1(keyinput_g44), .B2(n6858), .ZN(n6796) );
  OAI221_X1 U7754 ( .B1(n6845), .B2(keyinput_g18), .C1(n6858), .C2(
        keyinput_g44), .A(n6796), .ZN(n6806) );
  AOI22_X1 U7755 ( .A1(n7026), .A2(keyinput_g40), .B1(n6798), .B2(keyinput_g47), .ZN(n6797) );
  OAI221_X1 U7756 ( .B1(n7026), .B2(keyinput_g40), .C1(n6798), .C2(
        keyinput_g47), .A(n6797), .ZN(n6805) );
  AOI22_X1 U7757 ( .A1(n6800), .A2(keyinput_g118), .B1(keyinput_g70), .B2(
        n6975), .ZN(n6799) );
  OAI221_X1 U7758 ( .B1(n6800), .B2(keyinput_g118), .C1(n6975), .C2(
        keyinput_g70), .A(n6799), .ZN(n6804) );
  INV_X1 U7759 ( .A(CODEFETCH_REG_SCAN_IN), .ZN(n6802) );
  AOI22_X1 U7760 ( .A1(n6873), .A2(keyinput_g90), .B1(n6802), .B2(keyinput_g39), .ZN(n6801) );
  OAI221_X1 U7761 ( .B1(n6873), .B2(keyinput_g90), .C1(n6802), .C2(
        keyinput_g39), .A(n6801), .ZN(n6803) );
  NOR4_X1 U7762 ( .A1(n6806), .A2(n6805), .A3(n6804), .A4(n6803), .ZN(n6831)
         );
  AOI22_X1 U7763 ( .A1(n7008), .A2(keyinput_g25), .B1(keyinput_g84), .B2(n6808), .ZN(n6807) );
  OAI221_X1 U7764 ( .B1(n7008), .B2(keyinput_g25), .C1(n6808), .C2(
        keyinput_g84), .A(n6807), .ZN(n6817) );
  AOI22_X1 U7765 ( .A1(n6860), .A2(keyinput_g94), .B1(keyinput_g50), .B2(n6987), .ZN(n6809) );
  OAI221_X1 U7766 ( .B1(n6860), .B2(keyinput_g94), .C1(n6987), .C2(
        keyinput_g50), .A(n6809), .ZN(n6816) );
  AOI22_X1 U7767 ( .A1(n6811), .A2(keyinput_g53), .B1(keyinput_g119), .B2(
        n7010), .ZN(n6810) );
  OAI221_X1 U7768 ( .B1(n6811), .B2(keyinput_g53), .C1(n7010), .C2(
        keyinput_g119), .A(n6810), .ZN(n6815) );
  INV_X1 U7769 ( .A(DATAI_10_), .ZN(n6868) );
  AOI22_X1 U7770 ( .A1(n6813), .A2(keyinput_g95), .B1(n6868), .B2(keyinput_g21), .ZN(n6812) );
  OAI221_X1 U7771 ( .B1(n6813), .B2(keyinput_g95), .C1(n6868), .C2(
        keyinput_g21), .A(n6812), .ZN(n6814) );
  NOR4_X1 U7772 ( .A1(n6817), .A2(n6816), .A3(n6815), .A4(n6814), .ZN(n6830)
         );
  INV_X1 U7773 ( .A(DATAI_26_), .ZN(n7017) );
  AOI22_X1 U7774 ( .A1(n7004), .A2(keyinput_g38), .B1(n7017), .B2(keyinput_g5), 
        .ZN(n6818) );
  OAI221_X1 U7775 ( .B1(n7004), .B2(keyinput_g38), .C1(n7017), .C2(keyinput_g5), .A(n6818), .ZN(n6828) );
  AOI22_X1 U7776 ( .A1(n6820), .A2(keyinput_g115), .B1(n6844), .B2(
        keyinput_g49), .ZN(n6819) );
  OAI221_X1 U7777 ( .B1(n6820), .B2(keyinput_g115), .C1(n6844), .C2(
        keyinput_g49), .A(n6819), .ZN(n6827) );
  AOI22_X1 U7778 ( .A1(n6842), .A2(keyinput_g59), .B1(keyinput_g28), .B2(n6990), .ZN(n6821) );
  OAI221_X1 U7779 ( .B1(n6842), .B2(keyinput_g59), .C1(n6990), .C2(
        keyinput_g28), .A(n6821), .ZN(n6826) );
  AOI22_X1 U7780 ( .A1(n6824), .A2(keyinput_g123), .B1(keyinput_g83), .B2(
        n6823), .ZN(n6822) );
  OAI221_X1 U7781 ( .B1(n6824), .B2(keyinput_g123), .C1(n6823), .C2(
        keyinput_g83), .A(n6822), .ZN(n6825) );
  NOR4_X1 U7782 ( .A1(n6828), .A2(n6827), .A3(n6826), .A4(n6825), .ZN(n6829)
         );
  NAND4_X1 U7783 ( .A1(n6832), .A2(n6831), .A3(n6830), .A4(n6829), .ZN(n6833)
         );
  NOR4_X1 U7784 ( .A1(n6836), .A2(n6835), .A3(n6834), .A4(n6833), .ZN(n7046)
         );
  INV_X1 U7785 ( .A(DATAI_22_), .ZN(n6838) );
  AOI22_X1 U7786 ( .A1(n6839), .A2(keyinput_f30), .B1(n6838), .B2(keyinput_f9), 
        .ZN(n6837) );
  OAI221_X1 U7787 ( .B1(n6839), .B2(keyinput_f30), .C1(n6838), .C2(keyinput_f9), .A(n6837), .ZN(n7042) );
  OAI22_X1 U7788 ( .A1(n6842), .A2(keyinput_f59), .B1(n6841), .B2(
        keyinput_f117), .ZN(n6840) );
  AOI221_X1 U7789 ( .B1(n6842), .B2(keyinput_f59), .C1(keyinput_f117), .C2(
        n6841), .A(n6840), .ZN(n6849) );
  OAI22_X1 U7790 ( .A1(n6845), .A2(keyinput_f18), .B1(n6844), .B2(keyinput_f49), .ZN(n6843) );
  AOI221_X1 U7791 ( .B1(n6845), .B2(keyinput_f18), .C1(keyinput_f49), .C2(
        n6844), .A(n6843), .ZN(n6848) );
  XNOR2_X1 U7792 ( .A(keyinput_f126), .B(DATAWIDTH_REG_22__SCAN_IN), .ZN(n6847) );
  XNOR2_X1 U7793 ( .A(keyinput_f127), .B(DATAWIDTH_REG_23__SCAN_IN), .ZN(n6846) );
  NAND4_X1 U7794 ( .A1(n6849), .A2(n6848), .A3(n6847), .A4(n6846), .ZN(n7041)
         );
  AOI22_X1 U7795 ( .A1(n6852), .A2(keyinput_f43), .B1(keyinput_f14), .B2(n6851), .ZN(n6850) );
  OAI221_X1 U7796 ( .B1(n6852), .B2(keyinput_f43), .C1(n6851), .C2(
        keyinput_f14), .A(n6850), .ZN(n6865) );
  AOI22_X1 U7797 ( .A1(n6855), .A2(keyinput_f96), .B1(n6854), .B2(keyinput_f64), .ZN(n6853) );
  OAI221_X1 U7798 ( .B1(n6855), .B2(keyinput_f96), .C1(n6854), .C2(
        keyinput_f64), .A(n6853), .ZN(n6864) );
  AOI22_X1 U7799 ( .A1(n6858), .A2(keyinput_f44), .B1(keyinput_f114), .B2(
        n6857), .ZN(n6856) );
  OAI221_X1 U7800 ( .B1(n6858), .B2(keyinput_f44), .C1(n6857), .C2(
        keyinput_f114), .A(n6856), .ZN(n6863) );
  AOI22_X1 U7801 ( .A1(n6861), .A2(keyinput_f97), .B1(keyinput_f94), .B2(n6860), .ZN(n6859) );
  OAI221_X1 U7802 ( .B1(n6861), .B2(keyinput_f97), .C1(n6860), .C2(
        keyinput_f94), .A(n6859), .ZN(n6862) );
  NOR4_X1 U7803 ( .A1(n6865), .A2(n6864), .A3(n6863), .A4(n6862), .ZN(n6897)
         );
  AOI22_X1 U7804 ( .A1(n6868), .A2(keyinput_f21), .B1(keyinput_f91), .B2(n6867), .ZN(n6866) );
  OAI221_X1 U7805 ( .B1(n6868), .B2(keyinput_f21), .C1(n6867), .C2(
        keyinput_f91), .A(n6866), .ZN(n6880) );
  INV_X1 U7806 ( .A(keyinput_f34), .ZN(n6870) );
  AOI22_X1 U7807 ( .A1(n6871), .A2(keyinput_f60), .B1(BS16_N), .B2(n6870), 
        .ZN(n6869) );
  OAI221_X1 U7808 ( .B1(n6871), .B2(keyinput_f60), .C1(n6870), .C2(BS16_N), 
        .A(n6869), .ZN(n6879) );
  AOI22_X1 U7809 ( .A1(n5515), .A2(keyinput_f56), .B1(keyinput_f90), .B2(n6873), .ZN(n6872) );
  OAI221_X1 U7810 ( .B1(n5515), .B2(keyinput_f56), .C1(n6873), .C2(
        keyinput_f90), .A(n6872), .ZN(n6878) );
  AOI22_X1 U7811 ( .A1(n6876), .A2(keyinput_f99), .B1(n6875), .B2(keyinput_f55), .ZN(n6874) );
  OAI221_X1 U7812 ( .B1(n6876), .B2(keyinput_f99), .C1(n6875), .C2(
        keyinput_f55), .A(n6874), .ZN(n6877) );
  NOR4_X1 U7813 ( .A1(n6880), .A2(n6879), .A3(n6878), .A4(n6877), .ZN(n6896)
         );
  AOI22_X1 U7814 ( .A1(n6882), .A2(keyinput_f10), .B1(n4980), .B2(keyinput_f20), .ZN(n6881) );
  OAI221_X1 U7815 ( .B1(n6882), .B2(keyinput_f10), .C1(n4980), .C2(
        keyinput_f20), .A(n6881), .ZN(n6894) );
  AOI22_X1 U7816 ( .A1(n6884), .A2(keyinput_f71), .B1(n5415), .B2(keyinput_f52), .ZN(n6883) );
  OAI221_X1 U7817 ( .B1(n6884), .B2(keyinput_f71), .C1(n5415), .C2(
        keyinput_f52), .A(n6883), .ZN(n6893) );
  INV_X1 U7818 ( .A(DATAI_31_), .ZN(n6886) );
  AOI22_X1 U7819 ( .A1(n6887), .A2(keyinput_f15), .B1(n6886), .B2(keyinput_f0), 
        .ZN(n6885) );
  OAI221_X1 U7820 ( .B1(n6887), .B2(keyinput_f15), .C1(n6886), .C2(keyinput_f0), .A(n6885), .ZN(n6892) );
  AOI22_X1 U7821 ( .A1(n6890), .A2(keyinput_f69), .B1(keyinput_f72), .B2(n6889), .ZN(n6888) );
  OAI221_X1 U7822 ( .B1(n6890), .B2(keyinput_f69), .C1(n6889), .C2(
        keyinput_f72), .A(n6888), .ZN(n6891) );
  NOR4_X1 U7823 ( .A1(n6894), .A2(n6893), .A3(n6892), .A4(n6891), .ZN(n6895)
         );
  NAND3_X1 U7824 ( .A1(n6897), .A2(n6896), .A3(n6895), .ZN(n7040) );
  OAI22_X1 U7825 ( .A1(keyinput_f123), .A2(DATAWIDTH_REG_19__SCAN_IN), .B1(
        keyinput_f100), .B2(ADDRESS_REG_0__SCAN_IN), .ZN(n6898) );
  AOI221_X1 U7826 ( .B1(keyinput_f123), .B2(DATAWIDTH_REG_19__SCAN_IN), .C1(
        ADDRESS_REG_0__SCAN_IN), .C2(keyinput_f100), .A(n6898), .ZN(n6904) );
  OAI22_X1 U7827 ( .A1(DATAI_28_), .A2(keyinput_f3), .B1(keyinput_f32), .B2(
        MEMORYFETCH_REG_SCAN_IN), .ZN(n6899) );
  AOI221_X1 U7828 ( .B1(DATAI_28_), .B2(keyinput_f3), .C1(
        MEMORYFETCH_REG_SCAN_IN), .C2(keyinput_f32), .A(n6899), .ZN(n6903) );
  OAI22_X1 U7829 ( .A1(FLUSH_REG_SCAN_IN), .A2(keyinput_f45), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(keyinput_f88), .ZN(n6900) );
  AOI221_X1 U7830 ( .B1(FLUSH_REG_SCAN_IN), .B2(keyinput_f45), .C1(
        keyinput_f88), .C2(ADDRESS_REG_12__SCAN_IN), .A(n6900), .ZN(n6902) );
  XNOR2_X1 U7831 ( .A(DATAI_29_), .B(keyinput_f2), .ZN(n6901) );
  NAND4_X1 U7832 ( .A1(n6904), .A2(n6903), .A3(n6902), .A4(n6901), .ZN(n6932)
         );
  OAI22_X1 U7833 ( .A1(keyinput_f121), .A2(DATAWIDTH_REG_17__SCAN_IN), .B1(
        keyinput_f113), .B2(DATAWIDTH_REG_9__SCAN_IN), .ZN(n6905) );
  AOI221_X1 U7834 ( .B1(keyinput_f121), .B2(DATAWIDTH_REG_17__SCAN_IN), .C1(
        DATAWIDTH_REG_9__SCAN_IN), .C2(keyinput_f113), .A(n6905), .ZN(n6912)
         );
  OAI22_X1 U7835 ( .A1(keyinput_f75), .A2(ADDRESS_REG_25__SCAN_IN), .B1(
        keyinput_f109), .B2(DATAWIDTH_REG_5__SCAN_IN), .ZN(n6906) );
  AOI221_X1 U7836 ( .B1(keyinput_f75), .B2(ADDRESS_REG_25__SCAN_IN), .C1(
        DATAWIDTH_REG_5__SCAN_IN), .C2(keyinput_f109), .A(n6906), .ZN(n6911)
         );
  OAI22_X1 U7837 ( .A1(keyinput_f104), .A2(DATAWIDTH_REG_0__SCAN_IN), .B1(
        keyinput_f80), .B2(ADDRESS_REG_20__SCAN_IN), .ZN(n6907) );
  AOI221_X1 U7838 ( .B1(keyinput_f104), .B2(DATAWIDTH_REG_0__SCAN_IN), .C1(
        ADDRESS_REG_20__SCAN_IN), .C2(keyinput_f80), .A(n6907), .ZN(n6910) );
  OAI22_X1 U7839 ( .A1(REIP_REG_31__SCAN_IN), .A2(keyinput_f51), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(keyinput_f89), .ZN(n6908) );
  AOI221_X1 U7840 ( .B1(REIP_REG_31__SCAN_IN), .B2(keyinput_f51), .C1(
        keyinput_f89), .C2(ADDRESS_REG_11__SCAN_IN), .A(n6908), .ZN(n6909) );
  NAND4_X1 U7841 ( .A1(n6912), .A2(n6911), .A3(n6910), .A4(n6909), .ZN(n6931)
         );
  OAI22_X1 U7842 ( .A1(STATE_REG_0__SCAN_IN), .A2(keyinput_f103), .B1(
        REIP_REG_20__SCAN_IN), .B2(keyinput_f62), .ZN(n6913) );
  AOI221_X1 U7843 ( .B1(STATE_REG_0__SCAN_IN), .B2(keyinput_f103), .C1(
        keyinput_f62), .C2(REIP_REG_20__SCAN_IN), .A(n6913), .ZN(n6920) );
  OAI22_X1 U7844 ( .A1(REIP_REG_29__SCAN_IN), .A2(keyinput_f53), .B1(
        keyinput_f107), .B2(DATAWIDTH_REG_3__SCAN_IN), .ZN(n6914) );
  AOI221_X1 U7845 ( .B1(REIP_REG_29__SCAN_IN), .B2(keyinput_f53), .C1(
        DATAWIDTH_REG_3__SCAN_IN), .C2(keyinput_f107), .A(n6914), .ZN(n6919)
         );
  OAI22_X1 U7846 ( .A1(keyinput_f76), .A2(ADDRESS_REG_24__SCAN_IN), .B1(
        keyinput_f86), .B2(ADDRESS_REG_14__SCAN_IN), .ZN(n6915) );
  AOI221_X1 U7847 ( .B1(keyinput_f76), .B2(ADDRESS_REG_24__SCAN_IN), .C1(
        ADDRESS_REG_14__SCAN_IN), .C2(keyinput_f86), .A(n6915), .ZN(n6918) );
  OAI22_X1 U7848 ( .A1(DATAI_27_), .A2(keyinput_f4), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(keyinput_f82), .ZN(n6916) );
  AOI221_X1 U7849 ( .B1(DATAI_27_), .B2(keyinput_f4), .C1(keyinput_f82), .C2(
        ADDRESS_REG_18__SCAN_IN), .A(n6916), .ZN(n6917) );
  NAND4_X1 U7850 ( .A1(n6920), .A2(n6919), .A3(n6918), .A4(n6917), .ZN(n6930)
         );
  OAI22_X1 U7851 ( .A1(STATE_REG_1__SCAN_IN), .A2(keyinput_f102), .B1(
        keyinput_f6), .B2(DATAI_25_), .ZN(n6921) );
  AOI221_X1 U7852 ( .B1(STATE_REG_1__SCAN_IN), .B2(keyinput_f102), .C1(
        DATAI_25_), .C2(keyinput_f6), .A(n6921), .ZN(n6928) );
  OAI22_X1 U7853 ( .A1(REQUESTPENDING_REG_SCAN_IN), .A2(keyinput_f42), .B1(
        keyinput_f36), .B2(HOLD), .ZN(n6922) );
  AOI221_X1 U7854 ( .B1(REQUESTPENDING_REG_SCAN_IN), .B2(keyinput_f42), .C1(
        HOLD), .C2(keyinput_f36), .A(n6922), .ZN(n6927) );
  OAI22_X1 U7855 ( .A1(REIP_REG_17__SCAN_IN), .A2(keyinput_f65), .B1(
        keyinput_f47), .B2(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6923) );
  AOI221_X1 U7856 ( .B1(REIP_REG_17__SCAN_IN), .B2(keyinput_f65), .C1(
        BYTEENABLE_REG_0__SCAN_IN), .C2(keyinput_f47), .A(n6923), .ZN(n6926)
         );
  OAI22_X1 U7857 ( .A1(STATE_REG_2__SCAN_IN), .A2(keyinput_f101), .B1(
        keyinput_f67), .B2(BE_N_REG_3__SCAN_IN), .ZN(n6924) );
  AOI221_X1 U7858 ( .B1(STATE_REG_2__SCAN_IN), .B2(keyinput_f101), .C1(
        BE_N_REG_3__SCAN_IN), .C2(keyinput_f67), .A(n6924), .ZN(n6925) );
  NAND4_X1 U7859 ( .A1(n6928), .A2(n6927), .A3(n6926), .A4(n6925), .ZN(n6929)
         );
  NOR4_X1 U7860 ( .A1(n6932), .A2(n6931), .A3(n6930), .A4(n6929), .ZN(n7038)
         );
  OAI22_X1 U7861 ( .A1(keyinput_f83), .A2(ADDRESS_REG_17__SCAN_IN), .B1(
        keyinput_f118), .B2(DATAWIDTH_REG_14__SCAN_IN), .ZN(n6933) );
  AOI221_X1 U7862 ( .B1(keyinput_f83), .B2(ADDRESS_REG_17__SCAN_IN), .C1(
        DATAWIDTH_REG_14__SCAN_IN), .C2(keyinput_f118), .A(n6933), .ZN(n6940)
         );
  OAI22_X1 U7863 ( .A1(DATAI_18_), .A2(keyinput_f13), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(keyinput_f79), .ZN(n6934) );
  AOI221_X1 U7864 ( .B1(DATAI_18_), .B2(keyinput_f13), .C1(keyinput_f79), .C2(
        ADDRESS_REG_21__SCAN_IN), .A(n6934), .ZN(n6939) );
  OAI22_X1 U7865 ( .A1(ADDRESS_REG_16__SCAN_IN), .A2(keyinput_f84), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(keyinput_f77), .ZN(n6935) );
  AOI221_X1 U7866 ( .B1(ADDRESS_REG_16__SCAN_IN), .B2(keyinput_f84), .C1(
        keyinput_f77), .C2(ADDRESS_REG_23__SCAN_IN), .A(n6935), .ZN(n6938) );
  OAI22_X1 U7867 ( .A1(DATAI_9_), .A2(keyinput_f22), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(keyinput_f92), .ZN(n6936) );
  AOI221_X1 U7868 ( .B1(DATAI_9_), .B2(keyinput_f22), .C1(keyinput_f92), .C2(
        ADDRESS_REG_8__SCAN_IN), .A(n6936), .ZN(n6937) );
  NAND4_X1 U7869 ( .A1(n6940), .A2(n6939), .A3(n6938), .A4(n6937), .ZN(n6969)
         );
  OAI22_X1 U7870 ( .A1(DATAI_19_), .A2(keyinput_f12), .B1(keyinput_f29), .B2(
        DATAI_2_), .ZN(n6941) );
  AOI221_X1 U7871 ( .B1(DATAI_19_), .B2(keyinput_f12), .C1(DATAI_2_), .C2(
        keyinput_f29), .A(n6941), .ZN(n6948) );
  OAI22_X1 U7872 ( .A1(CODEFETCH_REG_SCAN_IN), .A2(keyinput_f39), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(keyinput_f93), .ZN(n6942) );
  AOI221_X1 U7873 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(keyinput_f39), .C1(
        keyinput_f93), .C2(ADDRESS_REG_7__SCAN_IN), .A(n6942), .ZN(n6947) );
  OAI22_X1 U7874 ( .A1(REIP_REG_24__SCAN_IN), .A2(keyinput_f58), .B1(
        keyinput_f63), .B2(REIP_REG_19__SCAN_IN), .ZN(n6943) );
  AOI221_X1 U7875 ( .B1(REIP_REG_24__SCAN_IN), .B2(keyinput_f58), .C1(
        REIP_REG_19__SCAN_IN), .C2(keyinput_f63), .A(n6943), .ZN(n6946) );
  OAI22_X1 U7876 ( .A1(REIP_REG_28__SCAN_IN), .A2(keyinput_f54), .B1(
        DATAWIDTH_REG_2__SCAN_IN), .B2(keyinput_f106), .ZN(n6944) );
  AOI221_X1 U7877 ( .B1(REIP_REG_28__SCAN_IN), .B2(keyinput_f54), .C1(
        keyinput_f106), .C2(DATAWIDTH_REG_2__SCAN_IN), .A(n6944), .ZN(n6945)
         );
  NAND4_X1 U7878 ( .A1(n6948), .A2(n6947), .A3(n6946), .A4(n6945), .ZN(n6968)
         );
  OAI22_X1 U7879 ( .A1(keyinput_f95), .A2(ADDRESS_REG_5__SCAN_IN), .B1(
        keyinput_f74), .B2(ADDRESS_REG_26__SCAN_IN), .ZN(n6949) );
  AOI221_X1 U7880 ( .B1(keyinput_f95), .B2(ADDRESS_REG_5__SCAN_IN), .C1(
        ADDRESS_REG_26__SCAN_IN), .C2(keyinput_f74), .A(n6949), .ZN(n6956) );
  OAI22_X1 U7881 ( .A1(READY_N), .A2(keyinput_f35), .B1(DATAI_12_), .B2(
        keyinput_f19), .ZN(n6950) );
  AOI221_X1 U7882 ( .B1(READY_N), .B2(keyinput_f35), .C1(keyinput_f19), .C2(
        DATAI_12_), .A(n6950), .ZN(n6955) );
  OAI22_X1 U7883 ( .A1(DATAI_5_), .A2(keyinput_f26), .B1(keyinput_f78), .B2(
        ADDRESS_REG_22__SCAN_IN), .ZN(n6951) );
  AOI221_X1 U7884 ( .B1(DATAI_5_), .B2(keyinput_f26), .C1(
        ADDRESS_REG_22__SCAN_IN), .C2(keyinput_f78), .A(n6951), .ZN(n6954) );
  OAI22_X1 U7885 ( .A1(keyinput_f105), .A2(DATAWIDTH_REG_1__SCAN_IN), .B1(
        keyinput_f120), .B2(DATAWIDTH_REG_16__SCAN_IN), .ZN(n6952) );
  AOI221_X1 U7886 ( .B1(keyinput_f105), .B2(DATAWIDTH_REG_1__SCAN_IN), .C1(
        DATAWIDTH_REG_16__SCAN_IN), .C2(keyinput_f120), .A(n6952), .ZN(n6953)
         );
  NAND4_X1 U7887 ( .A1(n6956), .A2(n6955), .A3(n6954), .A4(n6953), .ZN(n6967)
         );
  OAI22_X1 U7888 ( .A1(keyinput_f46), .A2(W_R_N_REG_SCAN_IN), .B1(
        keyinput_f111), .B2(DATAWIDTH_REG_7__SCAN_IN), .ZN(n6957) );
  AOI221_X1 U7889 ( .B1(keyinput_f46), .B2(W_R_N_REG_SCAN_IN), .C1(
        DATAWIDTH_REG_7__SCAN_IN), .C2(keyinput_f111), .A(n6957), .ZN(n6965)
         );
  OAI22_X1 U7890 ( .A1(keyinput_f98), .A2(ADDRESS_REG_2__SCAN_IN), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(keyinput_f87), .ZN(n6958) );
  AOI221_X1 U7891 ( .B1(keyinput_f98), .B2(ADDRESS_REG_2__SCAN_IN), .C1(
        keyinput_f87), .C2(ADDRESS_REG_13__SCAN_IN), .A(n6958), .ZN(n6964) );
  OAI22_X1 U7892 ( .A1(REIP_REG_16__SCAN_IN), .A2(keyinput_f66), .B1(
        keyinput_f73), .B2(ADDRESS_REG_27__SCAN_IN), .ZN(n6959) );
  AOI221_X1 U7893 ( .B1(REIP_REG_16__SCAN_IN), .B2(keyinput_f66), .C1(
        ADDRESS_REG_27__SCAN_IN), .C2(keyinput_f73), .A(n6959), .ZN(n6963) );
  OAI22_X1 U7894 ( .A1(n6961), .A2(keyinput_f24), .B1(NA_N), .B2(keyinput_f33), 
        .ZN(n6960) );
  AOI221_X1 U7895 ( .B1(n6961), .B2(keyinput_f24), .C1(keyinput_f33), .C2(NA_N), .A(n6960), .ZN(n6962) );
  NAND4_X1 U7896 ( .A1(n6965), .A2(n6964), .A3(n6963), .A4(n6962), .ZN(n6966)
         );
  NOR4_X1 U7897 ( .A1(n6969), .A2(n6968), .A3(n6967), .A4(n6966), .ZN(n7037)
         );
  AOI22_X1 U7898 ( .A1(n6972), .A2(keyinput_f61), .B1(keyinput_f124), .B2(
        n6971), .ZN(n6970) );
  OAI221_X1 U7899 ( .B1(n6972), .B2(keyinput_f61), .C1(n6971), .C2(
        keyinput_f124), .A(n6970), .ZN(n6984) );
  INV_X1 U7900 ( .A(DATAI_20_), .ZN(n6974) );
  AOI22_X1 U7901 ( .A1(n6975), .A2(keyinput_f70), .B1(n6974), .B2(keyinput_f11), .ZN(n6973) );
  OAI221_X1 U7902 ( .B1(n6975), .B2(keyinput_f70), .C1(n6974), .C2(
        keyinput_f11), .A(n6973), .ZN(n6983) );
  INV_X1 U7903 ( .A(READREQUEST_REG_SCAN_IN), .ZN(n6977) );
  AOI22_X1 U7904 ( .A1(n6978), .A2(keyinput_f27), .B1(keyinput_f37), .B2(n6977), .ZN(n6976) );
  OAI221_X1 U7905 ( .B1(n6978), .B2(keyinput_f27), .C1(n6977), .C2(
        keyinput_f37), .A(n6976), .ZN(n6982) );
  AOI22_X1 U7906 ( .A1(n5136), .A2(keyinput_f17), .B1(keyinput_f110), .B2(
        n6980), .ZN(n6979) );
  OAI221_X1 U7907 ( .B1(n5136), .B2(keyinput_f17), .C1(n6980), .C2(
        keyinput_f110), .A(n6979), .ZN(n6981) );
  NOR4_X1 U7908 ( .A1(n6984), .A2(n6983), .A3(n6982), .A4(n6981), .ZN(n7036)
         );
  OAI22_X1 U7909 ( .A1(n6987), .A2(keyinput_f50), .B1(n6986), .B2(keyinput_f68), .ZN(n6985) );
  AOI221_X1 U7910 ( .B1(n6987), .B2(keyinput_f50), .C1(keyinput_f68), .C2(
        n6986), .A(n6985), .ZN(n7000) );
  INV_X1 U7911 ( .A(keyinput_f115), .ZN(n6989) );
  OAI22_X1 U7912 ( .A1(n6990), .A2(keyinput_f28), .B1(n6989), .B2(
        DATAWIDTH_REG_11__SCAN_IN), .ZN(n6988) );
  AOI221_X1 U7913 ( .B1(n6990), .B2(keyinput_f28), .C1(
        DATAWIDTH_REG_11__SCAN_IN), .C2(n6989), .A(n6988), .ZN(n6999) );
  OAI22_X1 U7914 ( .A1(n6993), .A2(keyinput_f16), .B1(n6992), .B2(keyinput_f48), .ZN(n6991) );
  AOI221_X1 U7915 ( .B1(n6993), .B2(keyinput_f16), .C1(keyinput_f48), .C2(
        n6992), .A(n6991), .ZN(n6998) );
  OAI22_X1 U7916 ( .A1(keyinput_f108), .A2(n6996), .B1(n6995), .B2(
        keyinput_f81), .ZN(n6994) );
  AOI221_X1 U7917 ( .B1(n6996), .B2(keyinput_f108), .C1(n6995), .C2(
        keyinput_f81), .A(n6994), .ZN(n6997) );
  NAND4_X1 U7918 ( .A1(n7000), .A2(n6999), .A3(n6998), .A4(n6997), .ZN(n7034)
         );
  OAI22_X1 U7919 ( .A1(n5444), .A2(keyinput_f57), .B1(n7002), .B2(keyinput_f1), 
        .ZN(n7001) );
  AOI221_X1 U7920 ( .B1(n5444), .B2(keyinput_f57), .C1(keyinput_f1), .C2(n7002), .A(n7001), .ZN(n7015) );
  OAI22_X1 U7921 ( .A1(keyinput_f122), .A2(n7005), .B1(n7004), .B2(
        keyinput_f38), .ZN(n7003) );
  AOI221_X1 U7922 ( .B1(n7005), .B2(keyinput_f122), .C1(n7004), .C2(
        keyinput_f38), .A(n7003), .ZN(n7014) );
  OAI22_X1 U7923 ( .A1(n7008), .A2(keyinput_f25), .B1(n7007), .B2(
        keyinput_f112), .ZN(n7006) );
  AOI221_X1 U7924 ( .B1(n7008), .B2(keyinput_f25), .C1(keyinput_f112), .C2(
        n7007), .A(n7006), .ZN(n7013) );
  INV_X1 U7925 ( .A(DATAI_23_), .ZN(n7011) );
  OAI22_X1 U7926 ( .A1(n7011), .A2(keyinput_f8), .B1(n7010), .B2(keyinput_f119), .ZN(n7009) );
  AOI221_X1 U7927 ( .B1(n7011), .B2(keyinput_f8), .C1(keyinput_f119), .C2(
        n7010), .A(n7009), .ZN(n7012) );
  NAND4_X1 U7928 ( .A1(n7015), .A2(n7014), .A3(n7013), .A4(n7012), .ZN(n7033)
         );
  AOI22_X1 U7929 ( .A1(n7018), .A2(keyinput_f41), .B1(n7017), .B2(keyinput_f5), 
        .ZN(n7016) );
  OAI221_X1 U7930 ( .B1(n7018), .B2(keyinput_f41), .C1(n7017), .C2(keyinput_f5), .A(n7016), .ZN(n7032) );
  INV_X1 U7931 ( .A(DATAI_24_), .ZN(n7021) );
  OAI22_X1 U7932 ( .A1(n7021), .A2(keyinput_f7), .B1(n7020), .B2(keyinput_f85), 
        .ZN(n7019) );
  AOI221_X1 U7933 ( .B1(n7021), .B2(keyinput_f7), .C1(keyinput_f85), .C2(n7020), .A(n7019), .ZN(n7030) );
  INV_X1 U7934 ( .A(DATAI_8_), .ZN(n7024) );
  OAI22_X1 U7935 ( .A1(n7024), .A2(keyinput_f23), .B1(n7023), .B2(keyinput_f31), .ZN(n7022) );
  AOI221_X1 U7936 ( .B1(n7024), .B2(keyinput_f23), .C1(keyinput_f31), .C2(
        n7023), .A(n7022), .ZN(n7029) );
  OAI22_X1 U7937 ( .A1(keyinput_f116), .A2(n7027), .B1(n7026), .B2(
        keyinput_f40), .ZN(n7025) );
  AOI221_X1 U7938 ( .B1(n7027), .B2(keyinput_f116), .C1(n7026), .C2(
        keyinput_f40), .A(n7025), .ZN(n7028) );
  NAND3_X1 U7939 ( .A1(n7030), .A2(n7029), .A3(n7028), .ZN(n7031) );
  NOR4_X1 U7940 ( .A1(n7034), .A2(n7033), .A3(n7032), .A4(n7031), .ZN(n7035)
         );
  NAND4_X1 U7941 ( .A1(n7038), .A2(n7037), .A3(n7036), .A4(n7035), .ZN(n7039)
         );
  NOR4_X1 U7942 ( .A1(n7042), .A2(n7041), .A3(n7040), .A4(n7039), .ZN(n7044)
         );
  XOR2_X1 U7943 ( .A(DATAWIDTH_REG_21__SCAN_IN), .B(keyinput_f125), .Z(n7043)
         );
  OAI22_X1 U7944 ( .A1(n7044), .A2(n7043), .B1(keyinput_g125), .B2(
        DATAWIDTH_REG_21__SCAN_IN), .ZN(n7045) );
  AOI211_X1 U7945 ( .C1(DATAWIDTH_REG_21__SCAN_IN), .C2(keyinput_g125), .A(
        n7046), .B(n7045), .ZN(n7050) );
  AOI22_X1 U7946 ( .A1(n7048), .A2(BYTEENABLE_REG_3__SCAN_IN), .B1(
        BE_N_REG_3__SCAN_IN), .B2(n7047), .ZN(n7049) );
  XNOR2_X1 U7947 ( .A(n7050), .B(n7049), .ZN(U3445) );
  CLKBUF_X1 U3608 ( .A(n4292), .Z(n3177) );
  CLKBUF_X1 U3619 ( .A(n5198), .Z(n5200) );
  CLKBUF_X1 U3635 ( .A(n5266), .Z(n5334) );
  BUF_X1 U3644 ( .A(n5275), .Z(n5370) );
  AND4_X1 U3660 ( .A1(n3219), .A2(n3218), .A3(n3217), .A4(n3216), .ZN(n3225)
         );
  CLKBUF_X1 U3704 ( .A(n4371), .Z(n5326) );
  CLKBUF_X1 U3836 ( .A(n5152), .Z(n5207) );
  CLKBUF_X1 U3846 ( .A(n5120), .Z(n5138) );
  CLKBUF_X1 U3848 ( .A(n5952), .Z(n5964) );
  XNOR2_X1 U3879 ( .A(n4379), .B(n4378), .ZN(n5316) );
  OR2_X1 U3972 ( .A1(n4795), .A2(n5203), .ZN(n7052) );
endmodule

