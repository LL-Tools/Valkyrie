

module b21_C_gen_AntiSAT_k_128_1 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2, 
        keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7, 
        keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12, 
        keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17, 
        keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22, 
        keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27, 
        keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32, 
        keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37, 
        keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42, 
        keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47, 
        keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52, 
        keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57, 
        keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62, 
        keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2, keyinput_g3, 
        keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, keyinput_g8, 
        keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, keyinput_g13, 
        keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, keyinput_g18, 
        keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, keyinput_g23, 
        keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, keyinput_g28, 
        keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, keyinput_g33, 
        keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, keyinput_g38, 
        keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, keyinput_g43, 
        keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, keyinput_g48, 
        keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, keyinput_g53, 
        keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, keyinput_g58, 
        keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, keyinput_g63, 
        ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58, 
        ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63, 
        ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51, 
        ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46, 
        U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, 
        P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, 
        P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, 
        P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, 
        P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440, P1_U3441, 
        P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, 
        P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, 
        P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, 
        P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, 
        P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463, P1_U3466, 
        P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484, P1_U3487, 
        P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505, P1_U3508, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289, P1_U3288, 
        P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, 
        P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, 
        P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, 
        P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262, P1_U3261, 
        P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, 
        P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, 
        P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238, P1_U3237, 
        P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, 
        P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, 
        P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, 
        P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084, P1_U3083, 
        P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354, P2_U3353, 
        P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347, P2_U3346, 
        P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340, P2_U3339, 
        P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333, P2_U3332, 
        P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437, P2_U3438, 
        P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, 
        P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, 
        P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, 
        P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, 
        P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, 
        P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, 
        P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502, P2_U3505, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, 
        P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533, P2_U3534, 
        P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, 
        P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, 
        P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294, P2_U3293, 
        P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, 
        P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, 
        P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, 
        P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, 
        P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, 
        P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, 
        P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3552, 
        P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, 
        P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565, P2_U3566, 
        P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572, P2_U3573, 
        P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579, P2_U3580, 
        P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152, P2_U3151, 
        P2_U3966 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2, keyinput_g3,
         keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, keyinput_g8,
         keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, keyinput_g13,
         keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, keyinput_g18,
         keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, keyinput_g23,
         keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, keyinput_g28,
         keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, keyinput_g33,
         keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, keyinput_g38,
         keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, keyinput_g43,
         keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, keyinput_g48,
         keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, keyinput_g53,
         keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, keyinput_g58,
         keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, keyinput_g63;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4306, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316,
         n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326,
         n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336,
         n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346,
         n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356,
         n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366,
         n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376,
         n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386,
         n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396,
         n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406,
         n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416,
         n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426,
         n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436,
         n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446,
         n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456,
         n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466,
         n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476,
         n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486,
         n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496,
         n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506,
         n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516,
         n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526,
         n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536,
         n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546,
         n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556,
         n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
         n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576,
         n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586,
         n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596,
         n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606,
         n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616,
         n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626,
         n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636,
         n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646,
         n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656,
         n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666,
         n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676,
         n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686,
         n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696,
         n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706,
         n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716,
         n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726,
         n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736,
         n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746,
         n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756,
         n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766,
         n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776,
         n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786,
         n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796,
         n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806,
         n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816,
         n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826,
         n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836,
         n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846,
         n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856,
         n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866,
         n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876,
         n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886,
         n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896,
         n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906,
         n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916,
         n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926,
         n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936,
         n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946,
         n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956,
         n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966,
         n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976,
         n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986,
         n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996,
         n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006,
         n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016,
         n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026,
         n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036,
         n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046,
         n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056,
         n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066,
         n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076,
         n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086,
         n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096,
         n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106,
         n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116,
         n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126,
         n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136,
         n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146,
         n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156,
         n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166,
         n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176,
         n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186,
         n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196,
         n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206,
         n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216,
         n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226,
         n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236,
         n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246,
         n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256,
         n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266,
         n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276,
         n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286,
         n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296,
         n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306,
         n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316,
         n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326,
         n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336,
         n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346,
         n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356,
         n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366,
         n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376,
         n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386,
         n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396,
         n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406,
         n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416,
         n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426,
         n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436,
         n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446,
         n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456,
         n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466,
         n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476,
         n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486,
         n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496,
         n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506,
         n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516,
         n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526,
         n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536,
         n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546,
         n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556,
         n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566,
         n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576,
         n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586,
         n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596,
         n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606,
         n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616,
         n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626,
         n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636,
         n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646,
         n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656,
         n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666,
         n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676,
         n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686,
         n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696,
         n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706,
         n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716,
         n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726,
         n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736,
         n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746,
         n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756,
         n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766,
         n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776,
         n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786,
         n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796,
         n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806,
         n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816,
         n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826,
         n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836,
         n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846,
         n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856,
         n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866,
         n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876,
         n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886,
         n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896,
         n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906,
         n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916,
         n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926,
         n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936,
         n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946,
         n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956,
         n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966,
         n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976,
         n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986,
         n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996,
         n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006,
         n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016,
         n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026,
         n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036,
         n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046,
         n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056,
         n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066,
         n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076,
         n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086,
         n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096,
         n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106,
         n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116,
         n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126,
         n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136,
         n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146,
         n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156,
         n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166,
         n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176,
         n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186,
         n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196,
         n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206,
         n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216,
         n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226,
         n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236,
         n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246,
         n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256,
         n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266,
         n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276,
         n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286,
         n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296,
         n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306,
         n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316,
         n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326,
         n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336,
         n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346,
         n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356,
         n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366,
         n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376,
         n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386,
         n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396,
         n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406,
         n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416,
         n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426,
         n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436,
         n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446,
         n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456,
         n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466,
         n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476,
         n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486,
         n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496,
         n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506,
         n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516,
         n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526,
         n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536,
         n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546,
         n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556,
         n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566,
         n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576,
         n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586,
         n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596,
         n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606,
         n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616,
         n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626,
         n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636,
         n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646,
         n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656,
         n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666,
         n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676,
         n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686,
         n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696,
         n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706,
         n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716,
         n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726,
         n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736,
         n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746,
         n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756,
         n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766,
         n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776,
         n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786,
         n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796,
         n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806,
         n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816,
         n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826,
         n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836,
         n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846,
         n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856,
         n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866,
         n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876,
         n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886,
         n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896,
         n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906,
         n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916,
         n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926,
         n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936,
         n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946,
         n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956,
         n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966,
         n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976,
         n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986,
         n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996,
         n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006,
         n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016,
         n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026,
         n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036,
         n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046,
         n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056,
         n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066,
         n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076,
         n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086,
         n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096,
         n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106,
         n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116,
         n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126,
         n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136,
         n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146,
         n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156,
         n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166,
         n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176,
         n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186,
         n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196,
         n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206,
         n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216,
         n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226,
         n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236,
         n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246,
         n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256,
         n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266,
         n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276,
         n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286,
         n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296,
         n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306,
         n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316,
         n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326,
         n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336,
         n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346,
         n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356,
         n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366,
         n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376,
         n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386,
         n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396,
         n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406,
         n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416,
         n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426,
         n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436,
         n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446,
         n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456,
         n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466,
         n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476,
         n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486,
         n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496,
         n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506,
         n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516,
         n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526,
         n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536,
         n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546,
         n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556,
         n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566,
         n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576,
         n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586,
         n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596,
         n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606,
         n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616,
         n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626,
         n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636,
         n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646,
         n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656,
         n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666,
         n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676,
         n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686,
         n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696,
         n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706,
         n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716,
         n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726,
         n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736,
         n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746,
         n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756,
         n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766,
         n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776,
         n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786,
         n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796,
         n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806,
         n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816,
         n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826,
         n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836,
         n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846,
         n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856,
         n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866,
         n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876,
         n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886,
         n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896,
         n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906,
         n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916,
         n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926,
         n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936,
         n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946,
         n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956,
         n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966,
         n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976,
         n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986,
         n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996,
         n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006,
         n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016,
         n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026,
         n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036,
         n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046,
         n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056,
         n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066,
         n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076,
         n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086,
         n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096,
         n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106,
         n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116,
         n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126,
         n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136,
         n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146,
         n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156,
         n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166,
         n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176,
         n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186,
         n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196,
         n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206,
         n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216,
         n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226,
         n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236,
         n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246,
         n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256,
         n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266,
         n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276,
         n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286,
         n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296,
         n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306,
         n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316,
         n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326,
         n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336,
         n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346,
         n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356,
         n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366,
         n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376,
         n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386,
         n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396,
         n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406,
         n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416,
         n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426,
         n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436,
         n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446,
         n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456,
         n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466,
         n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476,
         n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486,
         n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496,
         n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506,
         n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516,
         n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526,
         n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536,
         n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546,
         n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556,
         n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566,
         n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576,
         n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586,
         n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596,
         n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606,
         n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616,
         n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626,
         n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636,
         n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646,
         n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656,
         n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666,
         n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676,
         n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686,
         n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696,
         n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706,
         n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716,
         n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726,
         n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736,
         n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746,
         n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756,
         n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766,
         n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776,
         n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786,
         n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796,
         n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806,
         n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816,
         n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826,
         n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836,
         n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846,
         n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856,
         n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866,
         n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876,
         n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886,
         n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896,
         n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906,
         n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916,
         n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926,
         n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936,
         n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946,
         n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956,
         n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966,
         n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976,
         n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986,
         n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996,
         n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006,
         n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016,
         n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026,
         n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036,
         n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046,
         n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056,
         n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066,
         n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076,
         n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086,
         n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096,
         n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106,
         n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116,
         n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126,
         n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136,
         n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146,
         n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156,
         n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166,
         n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176,
         n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186,
         n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196,
         n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206,
         n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216,
         n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226,
         n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236,
         n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246,
         n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256,
         n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266,
         n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276,
         n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286,
         n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296,
         n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306,
         n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316,
         n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326,
         n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336,
         n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346,
         n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356,
         n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366,
         n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376,
         n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386,
         n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396,
         n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406,
         n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416,
         n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426,
         n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436,
         n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446,
         n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456,
         n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466,
         n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476,
         n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486,
         n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496,
         n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506,
         n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516,
         n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526,
         n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536,
         n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546,
         n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556,
         n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566,
         n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576,
         n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586,
         n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596,
         n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606,
         n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616,
         n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626,
         n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636,
         n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646,
         n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656,
         n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666,
         n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676,
         n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686,
         n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696,
         n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706,
         n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716,
         n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726,
         n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736,
         n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746,
         n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756,
         n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766,
         n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776,
         n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786,
         n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796,
         n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806,
         n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816,
         n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826,
         n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836,
         n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846,
         n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856,
         n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866,
         n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876,
         n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886,
         n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896,
         n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906,
         n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916,
         n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926,
         n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936,
         n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946,
         n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956,
         n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966,
         n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976,
         n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986,
         n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996,
         n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005,
         n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013,
         n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021,
         n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029,
         n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037,
         n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045,
         n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053,
         n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061,
         n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069,
         n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077,
         n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085,
         n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093,
         n10094, n10095, n10096;

  OR3_X1 U4811 ( .A1(n8503), .A2(n8502), .A3(n8501), .ZN(n8561) );
  AOI21_X1 U4812 ( .B1(n8464), .B2(n10034), .A(n4372), .ZN(n4434) );
  BUF_X2 U4813 ( .A(n4413), .Z(n7981) );
  NAND2_X1 U4815 ( .A1(n6124), .A2(n8283), .ZN(n6293) );
  INV_X2 U4816 ( .A(n5698), .ZN(n5750) );
  CLKBUF_X2 U4817 ( .A(n5697), .Z(n4310) );
  CLKBUF_X2 U4818 ( .A(n5005), .Z(n5451) );
  CLKBUF_X2 U4819 ( .A(n5004), .Z(n6280) );
  BUF_X4 U4820 ( .A(n5509), .Z(n4308) );
  NAND2_X1 U4821 ( .A1(n5658), .A2(n5657), .ZN(n8202) );
  XNOR2_X1 U4822 ( .A(n5665), .B(n5661), .ZN(n5666) );
  INV_X4 U4823 ( .A(n6170), .ZN(n5462) );
  INV_X1 U4824 ( .A(n7893), .ZN(n7966) );
  AND3_X1 U4825 ( .A1(n4758), .A2(n4757), .A3(n4756), .ZN(n4937) );
  INV_X1 U4826 ( .A(n6093), .ZN(n5732) );
  NAND2_X1 U4827 ( .A1(n8525), .A2(n8212), .ZN(n8043) );
  BUF_X1 U4828 ( .A(n5715), .Z(n7861) );
  NAND2_X1 U4829 ( .A1(n9921), .A2(n8814), .ZN(n6448) );
  INV_X1 U4830 ( .A(n5017), .ZN(n5311) );
  NOR2_X2 U4831 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n4922) );
  BUF_X2 U4832 ( .A(n5699), .Z(n4312) );
  OR2_X1 U4833 ( .A1(n6123), .A2(n8006), .ZN(n8524) );
  NAND2_X1 U4834 ( .A1(n8573), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5663) );
  NAND2_X1 U4835 ( .A1(n5017), .A2(n6170), .ZN(n5112) );
  AND2_X1 U4836 ( .A1(n9123), .A2(n9102), .ZN(n9100) );
  NAND2_X1 U4837 ( .A1(n5867), .A2(n5866), .ZN(n8550) );
  INV_X2 U4838 ( .A(n5942), .ZN(n6145) );
  NAND2_X1 U4839 ( .A1(n4845), .A2(n4341), .ZN(n6724) );
  MUX2_X1 U4840 ( .A(P1_IR_REG_0__SCAN_IN), .B(n6168), .S(n5017), .Z(n9930) );
  INV_X1 U4841 ( .A(n6279), .ZN(n5489) );
  AOI211_X1 U4842 ( .C1(n9294), .C2(n5550), .A(n9263), .B(n9054), .ZN(n9293)
         );
  INV_X1 U4843 ( .A(n8939), .ZN(n9941) );
  NAND2_X1 U4844 ( .A1(n5464), .A2(n5463), .ZN(n9060) );
  XNOR2_X1 U4846 ( .A(n5502), .B(P1_IR_REG_21__SCAN_IN), .ZN(n8814) );
  NAND4_X1 U4847 ( .A1(n4992), .A2(n4991), .A3(n4990), .A4(n4989), .ZN(n9001)
         );
  INV_X2 U4848 ( .A(n9918), .ZN(n9938) );
  INV_X1 U4849 ( .A(n9920), .ZN(n9911) );
  INV_X2 U4850 ( .A(n8524), .ZN(n7178) );
  BUF_X1 U4851 ( .A(n4987), .Z(n5509) );
  XNOR2_X1 U4852 ( .A(n4955), .B(n4954), .ZN(n5508) );
  AND2_X1 U4853 ( .A1(n5667), .A2(n8579), .ZN(n5699) );
  OR3_X1 U4854 ( .A1(n8800), .A2(n8805), .A3(n8884), .ZN(n4306) );
  MUX2_X2 U4855 ( .A(n8194), .B(n8193), .S(n8425), .Z(n8195) );
  OAI21_X2 U4856 ( .B1(n5034), .B2(n4564), .A(n4565), .ZN(n5062) );
  NAND4_X2 U4857 ( .A1(n4964), .A2(n4963), .A3(n4962), .A4(n4961), .ZN(n6454)
         );
  OAI21_X2 U4858 ( .B1(n6672), .B2(n6671), .A(n5780), .ZN(n6816) );
  OAI21_X2 U4859 ( .B1(n5322), .B2(n5323), .A(n5324), .ZN(n5338) );
  AOI21_X2 U4860 ( .B1(n4566), .B2(n5045), .A(n4385), .ZN(n4565) );
  XNOR2_X2 U4861 ( .A(n5047), .B(n9592), .ZN(n5045) );
  INV_X2 U4862 ( .A(n6864), .ZN(n8939) );
  INV_X1 U4863 ( .A(n8006), .ZN(n6122) );
  AOI21_X2 U4864 ( .B1(n8228), .B2(n8053), .A(n8052), .ZN(n8058) );
  OAI21_X2 U4865 ( .B1(n9176), .B2(n8756), .A(n8897), .ZN(n9163) );
  BUF_X4 U4866 ( .A(n5697), .Z(n4309) );
  AND2_X2 U4867 ( .A1(n8576), .A2(n5666), .ZN(n5697) );
  BUF_X2 U4868 ( .A(n5699), .Z(n4311) );
  AND2_X4 U4869 ( .A1(n7193), .A2(n6450), .ZN(n7146) );
  OAI21_X2 U4870 ( .B1(n7264), .B2(n7912), .A(n7920), .ZN(n7345) );
  AOI21_X2 U4871 ( .B1(n7174), .B2(n8016), .A(n7173), .ZN(n7264) );
  INV_X4 U4872 ( .A(n4520), .ZN(n7733) );
  OAI222_X1 U4873 ( .A1(n7729), .A2(n6180), .B1(n9420), .B2(n6179), .C1(n6328), 
        .C2(P1_U3084), .ZN(P1_U3349) );
  OAI211_X1 U4874 ( .C1(n5060), .C2(n6179), .A(n5023), .B(n5022), .ZN(n6935)
         );
  XNOR2_X1 U4875 ( .A(n4643), .B(n5031), .ZN(n6179) );
  NOR2_X2 U4876 ( .A1(n7033), .A2(n7120), .ZN(n7132) );
  NAND2_X2 U4877 ( .A1(n5787), .A2(n5786), .ZN(n7120) );
  OAI21_X2 U4878 ( .B1(n5222), .B2(n5221), .A(n5220), .ZN(n5242) );
  OAI21_X1 U4879 ( .B1(n4561), .B2(n4330), .A(n8034), .ZN(n4649) );
  NAND2_X1 U4880 ( .A1(n5432), .A2(n5431), .ZN(n9092) );
  NAND2_X1 U4881 ( .A1(n7891), .A2(n6630), .ZN(n4544) );
  NAND2_X1 U4882 ( .A1(n8081), .A2(n6686), .ZN(n6630) );
  NAND2_X1 U4883 ( .A1(n8080), .A2(n6655), .ZN(n7891) );
  BUF_X2 U4884 ( .A(n7146), .Z(n7666) );
  INV_X1 U4885 ( .A(n6627), .ZN(n6655) );
  INV_X1 U4886 ( .A(n6448), .ZN(n7193) );
  CLKBUF_X2 U4887 ( .A(P1_U4006), .Z(n4315) );
  NAND2_X2 U4888 ( .A1(n6122), .A2(n7874), .ZN(n6644) );
  NOR2_X1 U4889 ( .A1(n9067), .A2(n9061), .ZN(n5608) );
  AOI21_X1 U4890 ( .B1(n4467), .B2(n4466), .A(n4926), .ZN(n4465) );
  INV_X1 U4891 ( .A(n8465), .ZN(n8470) );
  AND2_X1 U4892 ( .A1(n4573), .A2(n4576), .ZN(n6158) );
  NAND2_X1 U4893 ( .A1(n6048), .A2(n7776), .ZN(n6052) );
  AND2_X1 U4894 ( .A1(n8787), .A2(n8786), .ZN(n8802) );
  NAND2_X1 U4895 ( .A1(n8271), .A2(n8049), .ZN(n8260) );
  AOI22_X1 U4896 ( .A1(n8790), .A2(n7981), .B1(n5715), .B2(
        P1_DATAO_REG_30__SCAN_IN), .ZN(n9696) );
  NAND2_X1 U4897 ( .A1(n7625), .A2(n7624), .ZN(n7631) );
  NAND2_X1 U4898 ( .A1(n5485), .A2(n5484), .ZN(n9294) );
  OR2_X1 U4899 ( .A1(n9299), .A2(n9087), .ZN(n8821) );
  NAND2_X1 U4900 ( .A1(n6069), .A2(n6068), .ZN(n8476) );
  NAND2_X1 U4901 ( .A1(n6054), .A2(n6053), .ZN(n8483) );
  NAND2_X1 U4902 ( .A1(n8342), .A2(n4834), .ZN(n4833) );
  CLKBUF_X1 U4903 ( .A(n5549), .Z(n9310) );
  NAND2_X1 U4904 ( .A1(n7784), .A2(n5934), .ZN(n7795) );
  XNOR2_X1 U4905 ( .A(n5442), .B(n5441), .ZN(n8587) );
  OAI21_X2 U4906 ( .B1(n7786), .B2(n7564), .A(n7785), .ZN(n7784) );
  NAND2_X1 U4907 ( .A1(n5393), .A2(n5392), .ZN(n9120) );
  NAND2_X1 U4908 ( .A1(n7578), .A2(n8732), .ZN(n9255) );
  NAND2_X1 U4909 ( .A1(n6025), .A2(n6024), .ZN(n8492) );
  NAND2_X1 U4910 ( .A1(n5376), .A2(n5375), .ZN(n9319) );
  NAND2_X1 U4911 ( .A1(n5986), .A2(n5985), .ZN(n8509) );
  NAND2_X1 U4912 ( .A1(n5982), .A2(n5981), .ZN(n8514) );
  NAND2_X1 U4913 ( .A1(n5969), .A2(n5968), .ZN(n8521) );
  NOR2_X1 U4914 ( .A1(n8525), .A2(n8416), .ZN(n4425) );
  NAND2_X1 U4915 ( .A1(n5252), .A2(n5251), .ZN(n9247) );
  NAND2_X1 U4916 ( .A1(n5953), .A2(n5952), .ZN(n8525) );
  NAND2_X1 U4917 ( .A1(n5939), .A2(n5938), .ZN(n8530) );
  INV_X1 U4918 ( .A(n8022), .ZN(n4313) );
  NAND2_X1 U4919 ( .A1(n5889), .A2(n5888), .ZN(n8544) );
  INV_X2 U4920 ( .A(n8422), .ZN(n8463) );
  NAND2_X1 U4921 ( .A1(n5852), .A2(n5851), .ZN(n7416) );
  NAND2_X1 U4922 ( .A1(n6650), .A2(n8426), .ZN(n8422) );
  NAND2_X1 U4923 ( .A1(n4481), .A2(n8944), .ZN(n6854) );
  INV_X2 U4924 ( .A(n10036), .ZN(n4314) );
  NAND2_X1 U4925 ( .A1(n4599), .A2(n5836), .ZN(n7338) );
  OR2_X1 U4926 ( .A1(n8082), .A2(n10008), .ZN(n6568) );
  NAND2_X1 U4927 ( .A1(n5819), .A2(n5818), .ZN(n7389) );
  NAND2_X2 U4928 ( .A1(n9272), .A2(n7200), .ZN(n9918) );
  NAND4_X1 U4929 ( .A1(n5703), .A2(n5702), .A3(n5701), .A4(n5700), .ZN(n8082)
         );
  NAND4_X1 U4930 ( .A1(n5714), .A2(n5713), .A3(n5712), .A4(n5711), .ZN(n8081)
         );
  NAND4_X2 U4931 ( .A1(n5671), .A2(n5670), .A3(n5669), .A4(n5668), .ZN(n8084)
         );
  BUF_X2 U4932 ( .A(n5732), .Z(n6070) );
  NAND2_X2 U4933 ( .A1(n5592), .A2(n6448), .ZN(n7736) );
  NAND4_X1 U4934 ( .A1(n5010), .A2(n5009), .A3(n5008), .A4(n5007), .ZN(n9000)
         );
  AND2_X1 U4935 ( .A1(n5667), .A2(n5666), .ZN(n5698) );
  OAI211_X1 U4936 ( .C1(n6225), .C2(n5731), .A(n5730), .B(n5729), .ZN(n6627)
         );
  AND2_X4 U4937 ( .A1(n6450), .A2(n6448), .ZN(n6865) );
  AND2_X1 U4938 ( .A1(n4949), .A2(n9418), .ZN(n4987) );
  AND2_X1 U4939 ( .A1(n9415), .A2(n9418), .ZN(n5005) );
  OR3_X2 U4940 ( .A1(n5533), .A2(n7503), .A3(n7545), .ZN(n6450) );
  INV_X1 U4941 ( .A(n5666), .ZN(n8579) );
  AND2_X1 U4942 ( .A1(n4949), .A2(n4948), .ZN(n5004) );
  XNOR2_X1 U4943 ( .A(n5642), .B(P2_IR_REG_20__SCAN_IN), .ZN(n8006) );
  OAI21_X1 U4944 ( .B1(n5498), .B2(P1_IR_REG_20__SCAN_IN), .A(n4492), .ZN(
        n5502) );
  XNOR2_X1 U4945 ( .A(n5525), .B(n5524), .ZN(n7545) );
  NAND2_X1 U4946 ( .A1(n5641), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5642) );
  NAND2_X1 U4947 ( .A1(n5657), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5656) );
  OR2_X1 U4948 ( .A1(n4331), .A2(n9410), .ZN(n5525) );
  NAND2_X1 U4949 ( .A1(n4460), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4955) );
  NAND2_X2 U4950 ( .A1(n5462), .A2(P1_U3084), .ZN(n9420) );
  OR2_X2 U4951 ( .A1(n5462), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6195) );
  OAI211_X1 U4952 ( .C1(n6170), .C2(P2_DATAO_REG_0__SCAN_IN), .A(SI_0_), .B(
        n4523), .ZN(n4973) );
  AND2_X1 U4953 ( .A1(n5652), .A2(n5651), .ZN(n5653) );
  NOR2_X1 U4954 ( .A1(n5629), .A2(n5628), .ZN(n5652) );
  INV_X1 U4955 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5647) );
  NOR2_X2 U4956 ( .A1(P1_ADDR_REG_19__SCAN_IN), .A2(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n9651) );
  INV_X1 U4957 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5765) );
  NOR2_X1 U4958 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n5625) );
  INV_X1 U4959 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5644) );
  NOR2_X1 U4960 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n4516) );
  INV_X1 U4961 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6120) );
  INV_X1 U4962 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n4942) );
  INV_X1 U4963 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5832) );
  INV_X1 U4964 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n6100) );
  INV_X1 U4965 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5816) );
  AND2_X1 U4966 ( .A1(P2_ADDR_REG_19__SCAN_IN), .A2(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n9650) );
  INV_X1 U4967 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5885) );
  INV_X1 U4968 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5882) );
  NAND2_X1 U4969 ( .A1(n8344), .A2(n8343), .ZN(n8342) );
  NAND2_X1 U4970 ( .A1(n8576), .A2(n8579), .ZN(n5942) );
  OAI22_X2 U4971 ( .A1(n7489), .A2(n8023), .B1(n8544), .B2(n8071), .ZN(n7490)
         );
  NOR3_X2 U4972 ( .A1(n9740), .A2(n9712), .A3(n4636), .ZN(n4634) );
  INV_X1 U4973 ( .A(n6225), .ZN(n4316) );
  BUF_X2 U4974 ( .A(n5684), .Z(n6225) );
  AOI22_X2 U4975 ( .A1(n8364), .A2(n4376), .B1(n8514), .B2(n8358), .ZN(n8350)
         );
  OAI22_X2 U4976 ( .A1(n8378), .A2(n8381), .B1(n8390), .B2(n8213), .ZN(n8364)
         );
  AOI22_X2 U4977 ( .A1(n8350), .A2(n8215), .B1(n8355), .B2(n8214), .ZN(n8339)
         );
  NOR2_X2 U4978 ( .A1(n8311), .A2(n8488), .ZN(n8294) );
  OR2_X2 U4979 ( .A1(n8327), .A2(n8492), .ZN(n8311) );
  NAND2_X1 U4980 ( .A1(n6041), .A2(n6040), .ZN(n8488) );
  INV_X1 U4981 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5496) );
  INV_X1 U4982 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n5119) );
  NAND2_X1 U4983 ( .A1(n8979), .A2(n9911), .ZN(n5592) );
  NAND2_X1 U4984 ( .A1(n4769), .A2(n4771), .ZN(n4766) );
  AOI21_X1 U4985 ( .B1(n4594), .B2(n4596), .A(n4592), .ZN(n4591) );
  INV_X1 U4986 ( .A(n5118), .ZN(n4592) );
  NAND3_X1 U4987 ( .A1(n6293), .A2(n6123), .A3(n8054), .ZN(n5643) );
  NAND2_X1 U4988 ( .A1(n5636), .A2(n8054), .ZN(n6123) );
  NAND2_X1 U4989 ( .A1(n9255), .A2(n8862), .ZN(n4693) );
  AOI21_X1 U4990 ( .B1(n7925), .B2(n7924), .A(n7923), .ZN(n4553) );
  NAND2_X1 U4991 ( .A1(n4539), .A2(n8002), .ZN(n4536) );
  OAI21_X1 U4992 ( .B1(n4655), .B2(n4653), .A(n4540), .ZN(n4539) );
  NOR2_X1 U4993 ( .A1(n7958), .A2(n7956), .ZN(n4540) );
  OR2_X1 U4994 ( .A1(n4530), .A2(n4532), .ZN(n4526) );
  OAI21_X1 U4995 ( .B1(n9077), .B2(n8780), .A(n8779), .ZN(n8781) );
  AND2_X1 U4996 ( .A1(n4790), .A2(n5441), .ZN(n4789) );
  NAND2_X1 U4997 ( .A1(n5424), .A2(n5423), .ZN(n4790) );
  INV_X1 U4998 ( .A(n4725), .ZN(n4722) );
  NAND2_X1 U4999 ( .A1(n7794), .A2(n4726), .ZN(n4724) );
  NOR2_X1 U5000 ( .A1(n8244), .A2(n4353), .ZN(n4849) );
  NAND2_X1 U5001 ( .A1(n5632), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6101) );
  AND2_X1 U5002 ( .A1(n5644), .A2(n5637), .ZN(n5631) );
  NAND2_X1 U5003 ( .A1(n4498), .A2(n4497), .ZN(n4496) );
  AND2_X1 U5004 ( .A1(n4901), .A2(n4903), .ZN(n4899) );
  INV_X1 U5005 ( .A(n4900), .ZN(n4497) );
  OAI21_X1 U5006 ( .B1(n6932), .B2(n4485), .A(n4486), .ZN(n6955) );
  AOI21_X1 U5007 ( .B1(n6944), .B2(n4487), .A(n4366), .ZN(n4486) );
  OR2_X1 U5008 ( .A1(n9080), .A2(n9092), .ZN(n8894) );
  INV_X1 U5009 ( .A(n9228), .ZN(n4428) );
  NAND2_X1 U5010 ( .A1(n5575), .A2(n4747), .ZN(n4746) );
  NOR2_X1 U5011 ( .A1(n4320), .A2(n4754), .ZN(n4747) );
  OAI21_X1 U5012 ( .B1(n9874), .B2(n5567), .A(n4446), .ZN(n7403) );
  OR2_X1 U5013 ( .A1(n9875), .A2(n8995), .ZN(n4446) );
  NAND2_X1 U5014 ( .A1(n5139), .A2(n5138), .ZN(n5155) );
  AND2_X1 U5015 ( .A1(n5118), .A2(n5111), .ZN(n5116) );
  NAND2_X1 U5016 ( .A1(n5082), .A2(n5081), .ZN(n5085) );
  XNOR2_X1 U5017 ( .A(n7389), .B(n6070), .ZN(n5827) );
  NAND2_X1 U5018 ( .A1(n4703), .A2(n7258), .ZN(n4701) );
  INV_X1 U5019 ( .A(n4705), .ZN(n4703) );
  OAI21_X2 U5020 ( .B1(n7795), .B2(n4721), .A(n4717), .ZN(n7758) );
  AOI21_X1 U5021 ( .B1(n4720), .B2(n4719), .A(n4718), .ZN(n4717) );
  INV_X1 U5022 ( .A(n4723), .ZN(n4719) );
  INV_X1 U5023 ( .A(n7759), .ZN(n4718) );
  NAND2_X1 U5024 ( .A1(n6490), .A2(n4729), .ZN(n4728) );
  INV_X1 U5025 ( .A(n4311), .ZN(n6088) );
  NOR2_X1 U5026 ( .A1(n8471), .A2(n4777), .ZN(n4859) );
  NAND2_X1 U5027 ( .A1(n4379), .A2(n4329), .ZN(n4863) );
  AND2_X1 U5028 ( .A1(n8329), .A2(n8304), .ZN(n8216) );
  NOR2_X1 U5029 ( .A1(n8333), .A2(n4876), .ZN(n4875) );
  NAND2_X1 U5030 ( .A1(n8343), .A2(n4882), .ZN(n4876) );
  NAND2_X1 U5031 ( .A1(n4874), .A2(n4873), .ZN(n8308) );
  NOR2_X1 U5032 ( .A1(n4321), .A2(n8302), .ZN(n4873) );
  NAND2_X1 U5033 ( .A1(n8339), .A2(n4879), .ZN(n4874) );
  NAND2_X1 U5034 ( .A1(n4833), .A2(n4832), .ZN(n8301) );
  AND2_X1 U5035 ( .A1(n4347), .A2(n8302), .ZN(n4832) );
  NOR2_X1 U5036 ( .A1(n8339), .A2(n8343), .ZN(n4881) );
  INV_X1 U5037 ( .A(n6225), .ZN(n6188) );
  CLKBUF_X1 U5038 ( .A(n6122), .Z(n8034) );
  XNOR2_X1 U5039 ( .A(n6101), .B(n6100), .ZN(n5636) );
  XNOR2_X1 U5040 ( .A(n5640), .B(n5644), .ZN(n8054) );
  NAND2_X1 U5041 ( .A1(n6955), .A2(n6954), .ZN(n4910) );
  NOR2_X1 U5042 ( .A1(n7534), .A2(n4913), .ZN(n4912) );
  INV_X1 U5043 ( .A(n7530), .ZN(n4913) );
  XNOR2_X1 U5044 ( .A(n6878), .B(n7673), .ZN(n6882) );
  NAND2_X1 U5045 ( .A1(n6865), .A2(n6449), .ZN(n4520) );
  OR2_X1 U5046 ( .A1(n5433), .A2(n8688), .ZN(n5467) );
  AOI21_X1 U5047 ( .B1(n8809), .B2(n8887), .A(n8808), .ZN(n8816) );
  NAND2_X1 U5048 ( .A1(n4477), .A2(n4306), .ZN(n8809) );
  CLKBUF_X3 U5049 ( .A(n5004), .Z(n5510) );
  NOR2_X1 U5050 ( .A1(n9861), .A2(n4619), .ZN(n9036) );
  AND2_X1 U5051 ( .A1(n9859), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n4619) );
  NAND2_X1 U5052 ( .A1(n8821), .A2(n8880), .ZN(n9077) );
  NOR2_X1 U5053 ( .A1(n4767), .A2(n4454), .ZN(n4453) );
  INV_X1 U5054 ( .A(n5585), .ZN(n4454) );
  NAND2_X1 U5055 ( .A1(n4768), .A2(n4769), .ZN(n4767) );
  INV_X1 U5056 ( .A(n5589), .ZN(n4768) );
  INV_X1 U5057 ( .A(n4776), .ZN(n4773) );
  OR2_X1 U5058 ( .A1(n9152), .A2(n8987), .ZN(n4776) );
  OAI22_X1 U5059 ( .A1(n9174), .A2(n5584), .B1(n9197), .B2(n5548), .ZN(n9160)
         );
  NOR2_X1 U5060 ( .A1(n5578), .A2(n4751), .ZN(n4750) );
  INV_X1 U5061 ( .A(n5576), .ZN(n4751) );
  NAND2_X1 U5062 ( .A1(n7510), .A2(n4356), .ZN(n7578) );
  NAND2_X1 U5063 ( .A1(n7479), .A2(n5572), .ZN(n7506) );
  NAND2_X1 U5064 ( .A1(n7403), .A2(n8913), .ZN(n5569) );
  AND2_X1 U5065 ( .A1(n5135), .A2(n8911), .ZN(n4690) );
  NAND2_X1 U5066 ( .A1(n9883), .A2(n8848), .ZN(n4691) );
  NAND2_X1 U5067 ( .A1(n5052), .A2(n8949), .ZN(n4689) );
  INV_X1 U5068 ( .A(n4456), .ZN(n4455) );
  OAI21_X1 U5069 ( .B1(n4344), .B2(n4457), .A(n8908), .ZN(n4456) );
  INV_X1 U5070 ( .A(n5563), .ZN(n4457) );
  OR2_X1 U5071 ( .A1(n9922), .A2(n5591), .ZN(n9263) );
  NAND2_X1 U5072 ( .A1(n5506), .A2(n5505), .ZN(n9892) );
  XNOR2_X1 U5073 ( .A(n5500), .B(P1_IR_REG_22__SCAN_IN), .ZN(n8979) );
  NAND2_X1 U5074 ( .A1(n5499), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5500) );
  AOI21_X1 U5075 ( .B1(n5498), .B2(n4492), .A(n4490), .ZN(n4489) );
  XNOR2_X1 U5076 ( .A(n5155), .B(n5151), .ZN(n6218) );
  NAND2_X1 U5077 ( .A1(n4545), .A2(n4543), .ZN(n7892) );
  NAND2_X1 U5078 ( .A1(n4544), .A2(n7893), .ZN(n4543) );
  NAND2_X1 U5079 ( .A1(n7870), .A2(n7966), .ZN(n4545) );
  OAI21_X1 U5080 ( .B1(n4525), .B2(n4524), .A(n4369), .ZN(n7916) );
  AOI21_X1 U5081 ( .B1(n7882), .B2(n7881), .A(n4351), .ZN(n4524) );
  INV_X1 U5082 ( .A(n7899), .ZN(n4525) );
  INV_X1 U5083 ( .A(n7916), .ZN(n7914) );
  NAND2_X1 U5084 ( .A1(n4839), .A2(n7900), .ZN(n4652) );
  AOI21_X1 U5085 ( .B1(n8715), .B2(n4328), .A(n4374), .ZN(n4476) );
  AOI21_X1 U5086 ( .B1(n8708), .B2(n8848), .A(n4396), .ZN(n4474) );
  NAND2_X1 U5087 ( .A1(n8001), .A2(n8002), .ZN(n4542) );
  AND2_X1 U5088 ( .A1(n4547), .A2(n4546), .ZN(n7943) );
  NOR2_X1 U5089 ( .A1(n7937), .A2(n7936), .ZN(n4546) );
  NAND2_X1 U5090 ( .A1(n8038), .A2(n4659), .ZN(n4658) );
  INV_X1 U5091 ( .A(n7942), .ZN(n4659) );
  NAND2_X1 U5092 ( .A1(n4654), .A2(n8004), .ZN(n4653) );
  INV_X1 U5093 ( .A(n7955), .ZN(n4654) );
  INV_X1 U5094 ( .A(n4542), .ZN(n4535) );
  NAND2_X1 U5095 ( .A1(n4527), .A2(n4528), .ZN(n7961) );
  AOI21_X1 U5096 ( .B1(n4530), .B2(n4531), .A(n4529), .ZN(n4528) );
  NAND2_X1 U5097 ( .A1(n4536), .A2(n8044), .ZN(n4531) );
  NAND2_X1 U5098 ( .A1(n4558), .A2(n8048), .ZN(n4557) );
  NAND2_X1 U5099 ( .A1(n4559), .A2(n4644), .ZN(n4558) );
  NOR2_X1 U5100 ( .A1(n4645), .A2(n7998), .ZN(n4644) );
  NAND2_X1 U5101 ( .A1(n8291), .A2(n4555), .ZN(n4554) );
  NAND2_X1 U5102 ( .A1(n8492), .A2(n7969), .ZN(n4555) );
  NAND2_X1 U5103 ( .A1(n7968), .A2(n7966), .ZN(n4556) );
  AND2_X1 U5104 ( .A1(n4902), .A2(n8668), .ZN(n4901) );
  OR2_X1 U5105 ( .A1(n4903), .A2(n7656), .ZN(n4902) );
  NOR2_X1 U5106 ( .A1(n7712), .A2(n6170), .ZN(n4759) );
  INV_X1 U5107 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n4758) );
  INV_X1 U5108 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n4756) );
  NOR2_X1 U5109 ( .A1(n9341), .A2(n9219), .ZN(n4631) );
  INV_X1 U5110 ( .A(n5458), .ZN(n4782) );
  INV_X1 U5111 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5501) );
  AND2_X1 U5112 ( .A1(n4800), .A2(n5262), .ZN(n4799) );
  NAND2_X1 U5113 ( .A1(n5241), .A2(n5240), .ZN(n4800) );
  INV_X1 U5114 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n5223) );
  INV_X1 U5115 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n5181) );
  INV_X1 U5116 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n5180) );
  INV_X1 U5117 ( .A(SI_15_), .ZN(n9619) );
  AND2_X1 U5118 ( .A1(n4581), .A2(n4579), .ZN(n4578) );
  OR2_X1 U5119 ( .A1(n7769), .A2(n4584), .ZN(n4581) );
  NAND2_X1 U5120 ( .A1(n4580), .A2(n4582), .ZN(n4579) );
  NAND2_X1 U5121 ( .A1(n4808), .A2(n7966), .ZN(n4807) );
  INV_X1 U5122 ( .A(n8056), .ZN(n4808) );
  INV_X1 U5123 ( .A(n8053), .ZN(n7994) );
  OR2_X1 U5124 ( .A1(n6084), .A2(n6137), .ZN(n6139) );
  NAND2_X1 U5125 ( .A1(n6001), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6015) );
  NOR2_X1 U5126 ( .A1(n8509), .A2(n8514), .ZN(n4672) );
  NAND2_X1 U5127 ( .A1(n4842), .A2(n7900), .ZN(n4841) );
  AND2_X1 U5128 ( .A1(n7900), .A2(n7915), .ZN(n8014) );
  OR2_X1 U5129 ( .A1(n8435), .A2(n8436), .ZN(n4886) );
  CLKBUF_X1 U5130 ( .A(n5636), .Z(n7864) );
  AND2_X1 U5131 ( .A1(n6572), .A2(n6655), .ZN(n6636) );
  INV_X1 U5132 ( .A(n6179), .ZN(n4642) );
  INV_X1 U5133 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n4663) );
  NOR2_X2 U5134 ( .A1(n5950), .A2(P2_IR_REG_18__SCAN_IN), .ZN(n5638) );
  NAND2_X1 U5135 ( .A1(n9651), .A2(n4959), .ZN(n4522) );
  INV_X1 U5136 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4959) );
  NAND2_X1 U5137 ( .A1(n9650), .A2(n4960), .ZN(n4521) );
  INV_X1 U5138 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4960) );
  AND2_X1 U5139 ( .A1(n9921), .A2(n9911), .ZN(n5598) );
  OR2_X1 U5140 ( .A1(n7600), .A2(n4897), .ZN(n4896) );
  INV_X1 U5141 ( .A(n8594), .ZN(n4897) );
  NOR2_X1 U5142 ( .A1(n7601), .A2(n8594), .ZN(n4895) );
  AND2_X1 U5143 ( .A1(n8798), .A2(n8803), .ZN(n8807) );
  INV_X1 U5144 ( .A(n4453), .ZN(n4452) );
  NOR2_X1 U5145 ( .A1(n9183), .A2(n4630), .ZN(n4629) );
  INV_X1 U5146 ( .A(n4631), .ZN(n4630) );
  OR2_X1 U5147 ( .A1(n9183), .A2(n9197), .ZN(n8897) );
  OR2_X1 U5148 ( .A1(n7408), .A2(n9888), .ZN(n8849) );
  OAI21_X1 U5149 ( .B1(n5556), .B2(n4461), .A(n4966), .ZN(n6604) );
  AND2_X1 U5150 ( .A1(n9246), .A2(n9237), .ZN(n9231) );
  NOR2_X2 U5151 ( .A1(n9262), .A2(n9247), .ZN(n9246) );
  NAND2_X1 U5152 ( .A1(n5598), .A2(n8813), .ZN(n6449) );
  NAND2_X1 U5153 ( .A1(n5483), .A2(n5482), .ZN(n7848) );
  NAND2_X1 U5154 ( .A1(n5479), .A2(n5478), .ZN(n5483) );
  AND2_X1 U5155 ( .A1(n5443), .A2(n5430), .ZN(n5441) );
  NOR2_X1 U5156 ( .A1(n4920), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n4626) );
  AND2_X1 U5157 ( .A1(n5138), .A2(n5123), .ZN(n5136) );
  NOR2_X1 U5158 ( .A1(n5105), .A2(n4598), .ZN(n4597) );
  INV_X1 U5159 ( .A(n5084), .ZN(n4598) );
  NAND2_X1 U5160 ( .A1(n5066), .A2(n5065), .ZN(n5082) );
  INV_X1 U5161 ( .A(SI_8_), .ZN(n9496) );
  INV_X1 U5162 ( .A(SI_5_), .ZN(n9592) );
  NAND2_X1 U5163 ( .A1(n4734), .A2(n4733), .ZN(n7462) );
  AND2_X1 U5164 ( .A1(n5902), .A2(n5881), .ZN(n4733) );
  NAND2_X1 U5165 ( .A1(n5983), .A2(n4588), .ZN(n4587) );
  INV_X1 U5166 ( .A(n5984), .ZN(n4588) );
  NOR2_X1 U5167 ( .A1(n7808), .A2(n5972), .ZN(n4583) );
  NOR2_X1 U5168 ( .A1(n5848), .A2(n4601), .ZN(n4704) );
  INV_X1 U5169 ( .A(n5848), .ZN(n4602) );
  OAI21_X1 U5170 ( .B1(n4706), .B2(n4601), .A(n7163), .ZN(n4600) );
  INV_X1 U5171 ( .A(n6420), .ZN(n5726) );
  AND2_X1 U5172 ( .A1(n5814), .A2(n5797), .ZN(n4731) );
  OR2_X1 U5173 ( .A1(n5963), .A2(n9620), .ZN(n5974) );
  NAND2_X1 U5174 ( .A1(n5672), .A2(n5673), .ZN(n4730) );
  AND2_X1 U5175 ( .A1(n6663), .A2(n4322), .ZN(n4713) );
  OR2_X1 U5176 ( .A1(n6056), .A2(n6055), .ZN(n6073) );
  AOI21_X1 U5177 ( .B1(n7105), .B2(n7104), .A(n7103), .ZN(n7215) );
  NOR2_X1 U5178 ( .A1(n7994), .A2(n8052), .ZN(n8229) );
  NAND2_X1 U5179 ( .A1(n8288), .A2(n4861), .ZN(n4860) );
  NOR2_X1 U5180 ( .A1(n4862), .A2(n8225), .ZN(n4861) );
  INV_X1 U5181 ( .A(n4866), .ZN(n4862) );
  NAND2_X1 U5182 ( .A1(n8260), .A2(n4850), .ZN(n4848) );
  INV_X1 U5183 ( .A(n8224), .ZN(n8246) );
  NOR2_X1 U5184 ( .A1(n8260), .A2(n8261), .ZN(n8259) );
  INV_X1 U5185 ( .A(n4869), .ZN(n4868) );
  OAI21_X1 U5186 ( .B1(n4871), .B2(n8272), .A(n4870), .ZN(n4869) );
  NAND2_X1 U5187 ( .A1(n8198), .A2(n8262), .ZN(n4870) );
  NAND2_X1 U5188 ( .A1(n8222), .A2(n8269), .ZN(n4867) );
  INV_X1 U5189 ( .A(n4882), .ZN(n4880) );
  INV_X1 U5190 ( .A(n8359), .ZN(n8325) );
  AND2_X1 U5191 ( .A1(n8047), .A2(n7999), .ZN(n8343) );
  NAND3_X1 U5192 ( .A1(n8401), .A2(n8002), .A3(n8043), .ZN(n4820) );
  NAND2_X1 U5193 ( .A1(n4378), .A2(n8002), .ZN(n4821) );
  NAND2_X1 U5194 ( .A1(n8412), .A2(n8042), .ZN(n8401) );
  AND2_X1 U5195 ( .A1(n8042), .A2(n7952), .ZN(n8413) );
  AND2_X1 U5196 ( .A1(n7933), .A2(n7932), .ZN(n8022) );
  NAND2_X1 U5197 ( .A1(n7445), .A2(n8022), .ZN(n7444) );
  OR2_X1 U5198 ( .A1(n7340), .A2(n7416), .ZN(n7455) );
  NAND2_X1 U5199 ( .A1(n4853), .A2(n4852), .ZN(n7417) );
  AOI21_X1 U5200 ( .B1(n4854), .B2(n4857), .A(n4367), .ZN(n4852) );
  NAND2_X1 U5201 ( .A1(n7268), .A2(n4854), .ZN(n4853) );
  INV_X1 U5202 ( .A(n7187), .ZN(n4857) );
  OR2_X1 U5203 ( .A1(n7177), .A2(n7338), .ZN(n7340) );
  NAND2_X1 U5204 ( .A1(n7122), .A2(n4883), .ZN(n7186) );
  AND2_X1 U5205 ( .A1(n7123), .A2(n7121), .ZN(n4883) );
  AND2_X1 U5206 ( .A1(n7904), .A2(n7909), .ZN(n8016) );
  INV_X1 U5207 ( .A(n8014), .ZN(n7018) );
  OAI21_X1 U5208 ( .B1(n4826), .B2(n8011), .A(n4823), .ZN(n6632) );
  AOI21_X1 U5209 ( .B1(n4825), .B2(n7890), .A(n4824), .ZN(n4823) );
  NAND2_X1 U5210 ( .A1(n6632), .A2(n8013), .ZN(n6916) );
  AND2_X1 U5211 ( .A1(n7897), .A2(n7896), .ZN(n8013) );
  AND2_X1 U5212 ( .A1(n7869), .A2(n6568), .ZN(n7872) );
  NAND2_X1 U5213 ( .A1(n6505), .A2(n8009), .ZN(n6567) );
  NOR2_X1 U5214 ( .A1(n6758), .A2(n6512), .ZN(n6572) );
  NAND2_X1 U5215 ( .A1(n6753), .A2(n7879), .ZN(n6752) );
  INV_X1 U5216 ( .A(n8441), .ZN(n8326) );
  OR2_X1 U5217 ( .A1(n6222), .A2(n9992), .ZN(n7845) );
  AND2_X1 U5218 ( .A1(n6224), .A2(n6240), .ZN(n8440) );
  AND2_X1 U5219 ( .A1(n6224), .A2(n6150), .ZN(n8441) );
  NAND2_X1 U5220 ( .A1(n8581), .A2(n7981), .ZN(n4779) );
  NAND2_X1 U5221 ( .A1(n5923), .A2(n5922), .ZN(n8534) );
  AND2_X1 U5222 ( .A1(n8589), .A2(n6106), .ZN(n9991) );
  NAND2_X1 U5223 ( .A1(n6102), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6121) );
  OR2_X1 U5224 ( .A1(n5638), .A2(n8572), .ZN(n5634) );
  CLKBUF_X1 U5225 ( .A(n5746), .Z(n5766) );
  AOI21_X1 U5226 ( .B1(n4514), .B2(n4513), .A(n4348), .ZN(n4512) );
  INV_X1 U5227 ( .A(n8627), .ZN(n4513) );
  AND2_X1 U5228 ( .A1(n7702), .A2(n7701), .ZN(n7732) );
  NAND2_X1 U5229 ( .A1(n6862), .A2(n6861), .ZN(n6871) );
  XNOR2_X1 U5230 ( .A(n6868), .B(n7673), .ZN(n6872) );
  XNOR2_X1 U5231 ( .A(n6924), .B(n7736), .ZN(n6948) );
  AND2_X1 U5232 ( .A1(n7656), .A2(n4903), .ZN(n4900) );
  NAND2_X1 U5233 ( .A1(n4905), .A2(n4906), .ZN(n4517) );
  AOI21_X1 U5234 ( .B1(n7331), .B2(n7370), .A(n4907), .ZN(n4906) );
  INV_X1 U5235 ( .A(n7428), .ZN(n4907) );
  NAND2_X1 U5236 ( .A1(n5210), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n5234) );
  OR2_X1 U5237 ( .A1(n5234), .A2(n5233), .ZN(n5255) );
  INV_X1 U5238 ( .A(n5451), .ZN(n5486) );
  OR2_X1 U5239 ( .A1(n6474), .A2(n4384), .ZN(n4616) );
  INV_X1 U5240 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n4677) );
  NOR2_X1 U5241 ( .A1(n6347), .A2(n4393), .ZN(n6332) );
  AND2_X1 U5242 ( .A1(n9826), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6551) );
  NAND2_X1 U5243 ( .A1(n6767), .A2(n6766), .ZN(n6770) );
  OR2_X1 U5244 ( .A1(n7293), .A2(n7292), .ZN(n4614) );
  OR2_X1 U5245 ( .A1(n9026), .A2(n9025), .ZN(n4623) );
  NAND2_X1 U5246 ( .A1(n4623), .A2(n4622), .ZN(n4621) );
  NAND2_X1 U5247 ( .A1(n9039), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n4622) );
  AND2_X1 U5248 ( .A1(n4621), .A2(n4620), .ZN(n9861) );
  INV_X1 U5249 ( .A(n9862), .ZN(n4620) );
  OR2_X1 U5250 ( .A1(n9294), .A2(n4639), .ZN(n4638) );
  OR2_X1 U5251 ( .A1(n9060), .A2(n9299), .ZN(n4639) );
  AND2_X1 U5252 ( .A1(n4742), .A2(n9077), .ZN(n4741) );
  INV_X1 U5253 ( .A(n4925), .ZN(n4742) );
  AND2_X1 U5254 ( .A1(n8925), .A2(n4345), .ZN(n4743) );
  NAND2_X1 U5255 ( .A1(n5590), .A2(n8894), .ZN(n9071) );
  OR2_X1 U5256 ( .A1(n9110), .A2(n9887), .ZN(n4409) );
  AOI21_X1 U5257 ( .B1(n4772), .B2(n4770), .A(n4362), .ZN(n4769) );
  INV_X1 U5258 ( .A(n4339), .ZN(n4770) );
  NAND2_X1 U5259 ( .A1(n4687), .A2(n4686), .ZN(n9115) );
  NAND2_X1 U5260 ( .A1(n9161), .A2(n8758), .ZN(n9144) );
  NAND2_X1 U5261 ( .A1(n5586), .A2(n5585), .ZN(n9147) );
  NAND2_X1 U5262 ( .A1(n4440), .A2(n4439), .ZN(n9174) );
  AOI21_X1 U5263 ( .B1(n4323), .B2(n9205), .A(n4364), .ZN(n4439) );
  NAND2_X1 U5264 ( .A1(n9192), .A2(n8822), .ZN(n9176) );
  INV_X1 U5265 ( .A(n8827), .ZN(n4427) );
  AOI21_X1 U5266 ( .B1(n9209), .B2(n4443), .A(n4399), .ZN(n4442) );
  INV_X1 U5267 ( .A(n5582), .ZN(n4443) );
  NAND2_X1 U5268 ( .A1(n7506), .A2(n5573), .ZN(n5575) );
  NAND2_X1 U5269 ( .A1(n5569), .A2(n4398), .ZN(n9723) );
  AND2_X1 U5270 ( .A1(n8714), .A2(n9884), .ZN(n8909) );
  AND2_X1 U5271 ( .A1(n5071), .A2(n8706), .ZN(n4688) );
  INV_X1 U5272 ( .A(n8904), .ZN(n5561) );
  OR2_X1 U5273 ( .A1(n8810), .A2(n6898), .ZN(n9887) );
  INV_X1 U5274 ( .A(n9892), .ZN(n9732) );
  NAND2_X1 U5275 ( .A1(n8792), .A2(n8791), .ZN(n9053) );
  AND2_X1 U5276 ( .A1(n9946), .A2(n9945), .ZN(n9354) );
  OR2_X1 U5277 ( .A1(n5534), .A2(n5533), .ZN(n6207) );
  XNOR2_X1 U5278 ( .A(n7860), .B(n7859), .ZN(n8794) );
  NAND2_X1 U5279 ( .A1(n4947), .A2(n9411), .ZN(n4948) );
  NAND2_X1 U5280 ( .A1(n4484), .A2(n4483), .ZN(n4944) );
  INV_X1 U5281 ( .A(n4920), .ZN(n4625) );
  XNOR2_X1 U5282 ( .A(n5504), .B(P1_IR_REG_20__SCAN_IN), .ZN(n5591) );
  XNOR2_X1 U5283 ( .A(n5137), .B(n5136), .ZN(n6216) );
  NAND2_X1 U5284 ( .A1(n5013), .A2(SI_3_), .ZN(n5014) );
  NAND2_X1 U5285 ( .A1(n4716), .A2(n4720), .ZN(n7760) );
  NAND2_X1 U5286 ( .A1(n7795), .A2(n4723), .ZN(n4716) );
  NAND2_X1 U5287 ( .A1(n5683), .A2(n5682), .ZN(n6490) );
  NAND2_X1 U5288 ( .A1(n6297), .A2(n6093), .ZN(n5682) );
  NAND2_X1 U5289 ( .A1(n8524), .A2(n8086), .ZN(n5681) );
  INV_X1 U5290 ( .A(n8072), .ZN(n7469) );
  NAND2_X1 U5291 ( .A1(n4649), .A2(n4814), .ZN(n4813) );
  NAND2_X1 U5292 ( .A1(n6022), .A2(n6021), .ZN(n8304) );
  NAND2_X1 U5293 ( .A1(n6798), .A2(n6799), .ZN(n6802) );
  XNOR2_X1 U5294 ( .A(n4676), .B(n4675), .ZN(n9690) );
  INV_X1 U5295 ( .A(n9692), .ZN(n4675) );
  NOR2_X1 U5296 ( .A1(n8200), .A2(n8232), .ZN(n4676) );
  NAND2_X1 U5297 ( .A1(n5684), .A2(n4358), .ZN(n4710) );
  NAND2_X1 U5298 ( .A1(n5684), .A2(n4707), .ZN(n4709) );
  NAND2_X1 U5299 ( .A1(n5209), .A2(n5208), .ZN(n8719) );
  AOI21_X1 U5300 ( .B1(n4502), .B2(n4505), .A(n4377), .ZN(n4500) );
  NOR2_X1 U5301 ( .A1(n7633), .A2(n8678), .ZN(n4505) );
  NAND2_X1 U5302 ( .A1(n5167), .A2(n5166), .ZN(n7540) );
  OAI22_X2 U5303 ( .A1(n6974), .A2(n6975), .B1(n6884), .B2(n6883), .ZN(n6932)
         );
  NAND2_X1 U5304 ( .A1(n5115), .A2(n5114), .ZN(n9875) );
  NAND2_X1 U5305 ( .A1(n5359), .A2(n5358), .ZN(n9152) );
  XNOR2_X1 U5306 ( .A(n6882), .B(n6881), .ZN(n6975) );
  INV_X1 U5307 ( .A(n9117), .ZN(n9088) );
  AND2_X1 U5308 ( .A1(n5467), .A2(n5434), .ZN(n9093) );
  INV_X1 U5309 ( .A(n9722), .ZN(n8692) );
  AND2_X1 U5310 ( .A1(n6790), .A2(n9961), .ZN(n9717) );
  NAND2_X1 U5311 ( .A1(n5232), .A2(n5231), .ZN(n9712) );
  AOI21_X1 U5312 ( .B1(n8813), .B2(n8814), .A(n8816), .ZN(n4468) );
  NAND2_X1 U5313 ( .A1(n5401), .A2(n5400), .ZN(n8986) );
  NAND2_X1 U5314 ( .A1(n6621), .A2(n6622), .ZN(n6767) );
  NAND2_X1 U5315 ( .A1(n7061), .A2(n7060), .ZN(n7294) );
  OAI21_X1 U5316 ( .B1(n9041), .B2(n9847), .A(n4610), .ZN(n4609) );
  OR2_X1 U5317 ( .A1(n9042), .A2(n9797), .ZN(n4610) );
  OAI21_X1 U5318 ( .B1(n9045), .B2(n9044), .A(n9043), .ZN(n4604) );
  AOI21_X1 U5319 ( .B1(n4699), .B2(n9892), .A(n4696), .ZN(n9301) );
  NAND2_X1 U5320 ( .A1(n4698), .A2(n4697), .ZN(n4696) );
  NAND2_X1 U5321 ( .A1(n9080), .A2(n9730), .ZN(n4697) );
  NAND2_X1 U5322 ( .A1(n5142), .A2(n5141), .ZN(n9738) );
  INV_X1 U5323 ( .A(n9059), .ZN(n9881) );
  NAND2_X1 U5324 ( .A1(n4519), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5310) );
  OR2_X1 U5325 ( .A1(n5112), .A2(n4406), .ZN(n4984) );
  INV_X1 U5326 ( .A(n5591), .ZN(n9921) );
  OAI21_X1 U5327 ( .B1(n7892), .B2(n7872), .A(n4360), .ZN(n7873) );
  NAND2_X1 U5328 ( .A1(n4482), .A2(n4480), .ZN(n8700) );
  OAI21_X1 U5329 ( .B1(n6854), .B2(n8696), .A(n8799), .ZN(n4480) );
  NAND2_X1 U5330 ( .A1(n8697), .A2(n8805), .ZN(n4482) );
  NAND2_X1 U5331 ( .A1(n4651), .A2(n4650), .ZN(n7908) );
  NAND2_X1 U5332 ( .A1(n7907), .A2(n7893), .ZN(n4650) );
  OAI21_X1 U5333 ( .B1(n7914), .B2(n4652), .A(n4363), .ZN(n4651) );
  OAI21_X1 U5334 ( .B1(n4553), .B2(n7927), .A(n4549), .ZN(n4548) );
  NOR2_X1 U5335 ( .A1(n4550), .A2(n7893), .ZN(n4549) );
  INV_X1 U5336 ( .A(n7929), .ZN(n4550) );
  OAI21_X1 U5337 ( .B1(n4553), .B2(n7931), .A(n4552), .ZN(n4551) );
  AND2_X1 U5338 ( .A1(n7930), .A2(n7893), .ZN(n4552) );
  OAI21_X1 U5339 ( .B1(n4474), .B2(n8709), .A(n8799), .ZN(n4473) );
  OAI21_X1 U5340 ( .B1(n4476), .B2(n8717), .A(n8805), .ZN(n4475) );
  NOR2_X1 U5341 ( .A1(n7951), .A2(n8409), .ZN(n4655) );
  AOI21_X1 U5342 ( .B1(n4371), .B2(n4535), .A(n4533), .ZN(n4532) );
  OAI21_X1 U5343 ( .B1(n4542), .B2(n8003), .A(n7893), .ZN(n4533) );
  NOR2_X1 U5344 ( .A1(n8437), .A2(n7949), .ZN(n4656) );
  OR2_X1 U5345 ( .A1(n7943), .A2(n4658), .ZN(n4657) );
  AOI21_X1 U5346 ( .B1(n4375), .B2(n4536), .A(n7893), .ZN(n4530) );
  NAND2_X1 U5347 ( .A1(n4538), .A2(n8002), .ZN(n4537) );
  INV_X1 U5348 ( .A(n4653), .ZN(n4538) );
  AND2_X1 U5349 ( .A1(n4532), .A2(n4534), .ZN(n4529) );
  NAND2_X1 U5350 ( .A1(n4541), .A2(n4535), .ZN(n4534) );
  AND2_X1 U5351 ( .A1(n4655), .A2(n8043), .ZN(n4541) );
  OR2_X1 U5352 ( .A1(n7965), .A2(n7966), .ZN(n4560) );
  NAND2_X1 U5353 ( .A1(n4648), .A2(n4647), .ZN(n4646) );
  AND2_X1 U5354 ( .A1(n8047), .A2(n7966), .ZN(n4647) );
  OR2_X1 U5355 ( .A1(n7960), .A2(n7962), .ZN(n4648) );
  NOR2_X1 U5356 ( .A1(n4347), .A2(n7966), .ZN(n4645) );
  INV_X1 U5357 ( .A(n8867), .ZN(n4471) );
  NAND2_X1 U5358 ( .A1(n5997), .A2(n5998), .ZN(n4586) );
  AOI21_X1 U5359 ( .B1(n4557), .B2(n4556), .A(n4554), .ZN(n7976) );
  INV_X1 U5360 ( .A(n4583), .ZN(n4580) );
  INV_X1 U5361 ( .A(n4586), .ZN(n4584) );
  NOR2_X1 U5362 ( .A1(n8057), .A2(n4811), .ZN(n4810) );
  NAND2_X1 U5363 ( .A1(n7990), .A2(n4812), .ZN(n4811) );
  NAND2_X1 U5364 ( .A1(n7994), .A2(n7966), .ZN(n4812) );
  INV_X1 U5365 ( .A(n6931), .ZN(n4488) );
  INV_X1 U5366 ( .A(n6930), .ZN(n4487) );
  NAND2_X1 U5367 ( .A1(n6854), .A2(n8839), .ZN(n8697) );
  INV_X1 U5368 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n5304) );
  INV_X1 U5369 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n5244) );
  INV_X1 U5370 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n5157) );
  INV_X1 U5371 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n5156) );
  INV_X1 U5372 ( .A(n4595), .ZN(n4594) );
  OAI21_X1 U5373 ( .B1(n4597), .B2(n4596), .A(n5116), .ZN(n4595) );
  INV_X1 U5374 ( .A(n5106), .ZN(n4596) );
  INV_X1 U5375 ( .A(SI_10_), .ZN(n5120) );
  INV_X1 U5376 ( .A(SI_28_), .ZN(n9596) );
  OAI21_X1 U5377 ( .B1(n4849), .B2(n8051), .A(n4847), .ZN(n8228) );
  INV_X1 U5378 ( .A(n8050), .ZN(n4850) );
  OR2_X1 U5379 ( .A1(n8483), .A2(n8262), .ZN(n7973) );
  INV_X1 U5380 ( .A(n5988), .ZN(n5987) );
  INV_X1 U5381 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n9620) );
  OR2_X1 U5382 ( .A1(n8530), .A2(n8210), .ZN(n8042) );
  OR2_X1 U5383 ( .A1(n4667), .A2(n8539), .ZN(n4666) );
  NAND2_X1 U5384 ( .A1(n5890), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5913) );
  OR2_X1 U5385 ( .A1(n8544), .A2(n8550), .ZN(n4667) );
  NAND2_X1 U5386 ( .A1(n5868), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5891) );
  INV_X1 U5387 ( .A(n5870), .ZN(n5868) );
  AND2_X1 U5388 ( .A1(n8019), .A2(n4855), .ZN(n4854) );
  NAND2_X1 U5389 ( .A1(n4856), .A2(n7187), .ZN(n4855) );
  INV_X1 U5390 ( .A(n8017), .ZN(n4856) );
  INV_X1 U5391 ( .A(n5821), .ZN(n5820) );
  NOR2_X1 U5392 ( .A1(n7026), .A2(n4844), .ZN(n4843) );
  INV_X1 U5393 ( .A(n7871), .ZN(n4824) );
  INV_X1 U5394 ( .A(n4544), .ZN(n7890) );
  AND2_X1 U5395 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5733) );
  NAND2_X1 U5396 ( .A1(n8083), .A2(n6500), .ZN(n7887) );
  AOI21_X1 U5397 ( .B1(n9991), .B2(n9996), .A(n9997), .ZN(n6646) );
  NOR2_X1 U5398 ( .A1(n6701), .A2(n6731), .ZN(n6698) );
  NOR2_X1 U5399 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n5637) );
  INV_X1 U5400 ( .A(n7641), .ZN(n4890) );
  AND3_X1 U5401 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n5038) );
  OAI21_X1 U5402 ( .B1(n8802), .B2(n8788), .A(n4478), .ZN(n4477) );
  NOR2_X1 U5403 ( .A1(n8807), .A2(n4479), .ZN(n4478) );
  NAND2_X1 U5404 ( .A1(n8789), .A2(n4395), .ZN(n4479) );
  OR2_X1 U5405 ( .A1(n9053), .A2(n8793), .ZN(n8892) );
  OR2_X1 U5406 ( .A1(n9060), .A2(n7707), .ZN(n8817) );
  OAI21_X1 U5407 ( .B1(n4686), .B2(n4683), .A(n8820), .ZN(n4682) );
  INV_X1 U5408 ( .A(n8962), .ZN(n4683) );
  AND2_X1 U5409 ( .A1(n9116), .A2(n8866), .ZN(n4686) );
  OR2_X1 U5410 ( .A1(n9152), .A2(n9166), .ZN(n8896) );
  AND2_X1 U5411 ( .A1(n9207), .A2(n9206), .ZN(n8899) );
  OR2_X1 U5412 ( .A1(n4750), .A2(n4320), .ZN(n4749) );
  INV_X1 U5413 ( .A(n5574), .ZN(n4755) );
  NAND2_X1 U5414 ( .A1(n4637), .A2(n9747), .ZN(n4636) );
  AND2_X1 U5415 ( .A1(n5168), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5189) );
  NOR2_X1 U5416 ( .A1(n7561), .A2(n7540), .ZN(n4637) );
  OR2_X1 U5417 ( .A1(n7540), .A2(n7559), .ZN(n8729) );
  NOR2_X1 U5418 ( .A1(n5144), .A2(n5143), .ZN(n5168) );
  INV_X1 U5419 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5097) );
  NAND2_X1 U5420 ( .A1(n7190), .A2(n5566), .ZN(n9874) );
  NAND2_X1 U5421 ( .A1(n4633), .A2(n7203), .ZN(n7199) );
  INV_X1 U5422 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5053) );
  NOR2_X1 U5423 ( .A1(n7304), .A2(n7308), .ZN(n4633) );
  NAND2_X1 U5424 ( .A1(n6741), .A2(n6935), .ZN(n8841) );
  NAND2_X1 U5425 ( .A1(n9001), .A2(n7231), .ZN(n8838) );
  OAI211_X1 U5426 ( .C1(n5017), .C2(n4762), .A(n4761), .B(n4760), .ZN(n6864)
         );
  INV_X1 U5427 ( .A(n7726), .ZN(n4762) );
  NAND2_X1 U5428 ( .A1(n5017), .A2(n4759), .ZN(n4760) );
  NAND2_X1 U5429 ( .A1(n9231), .A2(n4629), .ZN(n9181) );
  NAND2_X1 U5430 ( .A1(n9231), .A2(n9400), .ZN(n9216) );
  NAND2_X1 U5431 ( .A1(n7852), .A2(n7851), .ZN(n7867) );
  NOR2_X1 U5432 ( .A1(n4940), .A2(n4373), .ZN(n4483) );
  NAND2_X1 U5433 ( .A1(n5461), .A2(n5460), .ZN(n5479) );
  NAND2_X1 U5434 ( .A1(n4783), .A2(n4781), .ZN(n5461) );
  AOI21_X1 U5435 ( .B1(n4784), .B2(n4787), .A(n4782), .ZN(n4781) );
  AND2_X1 U5436 ( .A1(n4327), .A2(n4459), .ZN(n4458) );
  AND2_X1 U5437 ( .A1(n5460), .A2(n5448), .ZN(n5458) );
  AOI21_X1 U5438 ( .B1(n4789), .B2(n4786), .A(n4785), .ZN(n4784) );
  INV_X1 U5439 ( .A(n5443), .ZN(n4785) );
  INV_X1 U5440 ( .A(n5423), .ZN(n4786) );
  INV_X1 U5441 ( .A(n4789), .ZN(n4787) );
  INV_X1 U5442 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5519) );
  NAND2_X1 U5443 ( .A1(n4941), .A2(n4933), .ZN(n4920) );
  OAI21_X1 U5444 ( .B1(n5369), .B2(n5368), .A(n5367), .ZN(n5388) );
  AND2_X1 U5445 ( .A1(n5389), .A2(n5374), .ZN(n5387) );
  NAND2_X1 U5446 ( .A1(n4491), .A2(n5501), .ZN(n4490) );
  NAND2_X1 U5447 ( .A1(n4492), .A2(P1_IR_REG_20__SCAN_IN), .ZN(n4491) );
  NOR2_X1 U5448 ( .A1(n9410), .A2(n4493), .ZN(n4492) );
  NOR2_X1 U5449 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n4493) );
  AND2_X1 U5450 ( .A1(n5339), .A2(n5328), .ZN(n5337) );
  AOI21_X1 U5451 ( .B1(n4324), .B2(n4797), .A(n4400), .ZN(n4791) );
  AOI21_X1 U5452 ( .B1(n4799), .B2(n4796), .A(n4795), .ZN(n4794) );
  INV_X1 U5453 ( .A(n5264), .ZN(n4795) );
  INV_X1 U5454 ( .A(n5240), .ZN(n4796) );
  INV_X1 U5455 ( .A(n4799), .ZN(n4797) );
  NOR2_X1 U5456 ( .A1(n5203), .A2(P1_IR_REG_13__SCAN_IN), .ZN(n5249) );
  OAI21_X1 U5457 ( .B1(n5177), .B2(n5178), .A(n5179), .ZN(n5200) );
  AND2_X1 U5458 ( .A1(n5201), .A2(n5184), .ZN(n5199) );
  NAND2_X1 U5459 ( .A1(n6170), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n4405) );
  INV_X1 U5460 ( .A(SI_14_), .ZN(n9533) );
  INV_X1 U5461 ( .A(SI_13_), .ZN(n9617) );
  INV_X1 U5462 ( .A(SI_21_), .ZN(n9589) );
  NAND2_X1 U5463 ( .A1(n4700), .A2(n4340), .ZN(n4734) );
  AND2_X1 U5464 ( .A1(n4726), .A2(n4725), .ZN(n4723) );
  NAND2_X1 U5465 ( .A1(n6157), .A2(n6066), .ZN(n4576) );
  OR2_X1 U5466 ( .A1(n5853), .A2(n9593), .ZN(n5870) );
  INV_X1 U5467 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n9593) );
  OR2_X1 U5468 ( .A1(n5913), .A2(n5912), .ZN(n5925) );
  XNOR2_X1 U5469 ( .A(n6010), .B(n6011), .ZN(n7815) );
  NAND2_X1 U5470 ( .A1(n7815), .A2(n7814), .ZN(n7813) );
  NAND2_X1 U5471 ( .A1(n5954), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5963) );
  OR2_X1 U5472 ( .A1(n5949), .A2(n5948), .ZN(n4726) );
  NAND2_X1 U5473 ( .A1(n5745), .A2(n4715), .ZN(n4714) );
  INV_X1 U5474 ( .A(n6428), .ZN(n4715) );
  NOR2_X1 U5475 ( .A1(n6148), .A2(n7844), .ZN(n7763) );
  OR2_X1 U5476 ( .A1(n7178), .A2(n8063), .ZN(n4816) );
  AND2_X1 U5477 ( .A1(n7993), .A2(n7893), .ZN(n4805) );
  INV_X1 U5478 ( .A(n8065), .ZN(n4814) );
  INV_X1 U5479 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n4416) );
  XNOR2_X1 U5480 ( .A(n8228), .B(n8229), .ZN(n4438) );
  AND2_X1 U5481 ( .A1(n6139), .A2(n6085), .ZN(n8242) );
  INV_X1 U5482 ( .A(n8199), .ZN(n8255) );
  NOR2_X1 U5483 ( .A1(n8253), .A2(n4867), .ZN(n4866) );
  NAND2_X1 U5484 ( .A1(n8294), .A2(n8198), .ZN(n8278) );
  NAND3_X1 U5485 ( .A1(n8289), .A2(n8272), .A3(n8273), .ZN(n8271) );
  OR2_X1 U5486 ( .A1(n8488), .A2(n8220), .ZN(n8273) );
  NAND2_X1 U5487 ( .A1(n8290), .A2(n8291), .ZN(n8289) );
  NOR2_X1 U5488 ( .A1(n8329), .A2(n4670), .ZN(n4668) );
  NAND2_X1 U5489 ( .A1(n4376), .A2(n8044), .ZN(n4818) );
  NAND2_X1 U5490 ( .A1(n8384), .A2(n4672), .ZN(n8351) );
  AND2_X1 U5491 ( .A1(n8000), .A2(n8045), .ZN(n8356) );
  NAND2_X1 U5492 ( .A1(n8384), .A2(n8371), .ZN(n8365) );
  AOI21_X1 U5493 ( .B1(n4319), .B2(n8436), .A(n4370), .ZN(n4884) );
  OR2_X1 U5494 ( .A1(n5940), .A2(n9500), .ZN(n5956) );
  NAND2_X1 U5495 ( .A1(n5924), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5940) );
  INV_X1 U5496 ( .A(n5925), .ZN(n5924) );
  NAND2_X1 U5497 ( .A1(n4665), .A2(n4664), .ZN(n8449) );
  NOR2_X1 U5498 ( .A1(n4666), .A2(n8534), .ZN(n4664) );
  INV_X1 U5499 ( .A(n7455), .ZN(n4665) );
  INV_X1 U5500 ( .A(n4829), .ZN(n4828) );
  OAI21_X1 U5501 ( .B1(n7936), .B2(n4830), .A(n7938), .ZN(n4829) );
  NOR2_X1 U5502 ( .A1(n7455), .A2(n4666), .ZN(n8448) );
  NOR2_X1 U5503 ( .A1(n7455), .A2(n4667), .ZN(n7492) );
  NOR2_X1 U5504 ( .A1(n7455), .A2(n8550), .ZN(n7454) );
  INV_X1 U5505 ( .A(n8073), .ZN(n7446) );
  NAND2_X1 U5506 ( .A1(n7268), .A2(n8017), .ZN(n7267) );
  OR2_X1 U5507 ( .A1(n5802), .A2(n5801), .ZN(n5821) );
  OR2_X1 U5508 ( .A1(n5788), .A2(n9590), .ZN(n5802) );
  OAI21_X1 U5509 ( .B1(n6916), .B2(n4838), .A(n4836), .ZN(n7174) );
  INV_X1 U5510 ( .A(n4837), .ZN(n4836) );
  NAND2_X1 U5511 ( .A1(n4840), .A2(n7900), .ZN(n7126) );
  NAND2_X1 U5512 ( .A1(n6916), .A2(n4843), .ZN(n4840) );
  NAND2_X1 U5513 ( .A1(n6636), .A2(n6664), .ZN(n6912) );
  OR2_X1 U5514 ( .A1(n8421), .A2(n8283), .ZN(n7450) );
  NAND2_X1 U5515 ( .A1(n4413), .A2(n4412), .ZN(n4411) );
  INV_X1 U5516 ( .A(n6174), .ZN(n4412) );
  NOR2_X1 U5517 ( .A1(n7712), .A2(n4708), .ZN(n4707) );
  OR2_X1 U5518 ( .A1(n8086), .A2(n6297), .ZN(n6443) );
  AND2_X1 U5519 ( .A1(n8467), .A2(n9693), .ZN(n8468) );
  NAND2_X1 U5520 ( .A1(n4886), .A2(n4319), .ZN(n8408) );
  AND2_X1 U5521 ( .A1(n4886), .A2(n4380), .ZN(n8410) );
  NAND3_X1 U5522 ( .A1(n5720), .A2(n4641), .A3(n4640), .ZN(n6512) );
  NAND2_X1 U5523 ( .A1(n4642), .A2(n4413), .ZN(n4641) );
  NAND2_X1 U5524 ( .A1(n4316), .A2(n8094), .ZN(n4640) );
  INV_X1 U5525 ( .A(n10031), .ZN(n9693) );
  INV_X1 U5526 ( .A(n10034), .ZN(n8549) );
  AND2_X1 U5527 ( .A1(n4334), .A2(n5655), .ZN(n4887) );
  NOR2_X1 U5528 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n5630) );
  OR3_X1 U5529 ( .A1(n5849), .A2(P2_IR_REG_10__SCAN_IN), .A3(
        P2_IR_REG_11__SCAN_IN), .ZN(n5865) );
  OR2_X1 U5530 ( .A1(n5781), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n5782) );
  NOR2_X1 U5531 ( .A1(n5782), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n5817) );
  INV_X1 U5532 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5624) );
  AND2_X1 U5533 ( .A1(n4368), .A2(n4503), .ZN(n4502) );
  OR2_X1 U5534 ( .A1(n7632), .A2(n4504), .ZN(n4503) );
  INV_X1 U5535 ( .A(n8678), .ZN(n4504) );
  NAND2_X1 U5536 ( .A1(n5413), .A2(n5412), .ZN(n5549) );
  NAND2_X1 U5537 ( .A1(n8603), .A2(n8605), .ZN(n4898) );
  NAND2_X1 U5538 ( .A1(n4494), .A2(n7670), .ZN(n8602) );
  NAND2_X1 U5539 ( .A1(n8675), .A2(n8678), .ZN(n7634) );
  NAND2_X1 U5540 ( .A1(n5360), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n5379) );
  INV_X1 U5541 ( .A(n5362), .ZN(n5360) );
  NAND2_X1 U5542 ( .A1(n7631), .A2(n7632), .ZN(n8675) );
  NAND2_X1 U5543 ( .A1(n4501), .A2(n7633), .ZN(n8676) );
  INV_X1 U5544 ( .A(n7631), .ZN(n4501) );
  NAND2_X1 U5545 ( .A1(n5275), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5316) );
  INV_X1 U5546 ( .A(n5291), .ZN(n5275) );
  INV_X1 U5547 ( .A(n9709), .ZN(n8669) );
  AND2_X1 U5548 ( .A1(n4894), .A2(n7607), .ZN(n4893) );
  OR2_X1 U5549 ( .A1(n4895), .A2(n4896), .ZN(n4894) );
  NAND2_X1 U5550 ( .A1(n4892), .A2(n7608), .ZN(n9713) );
  NAND2_X1 U5551 ( .A1(n8814), .A2(n8979), .ZN(n8810) );
  NAND2_X1 U5552 ( .A1(n5005), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n4953) );
  XNOR2_X1 U5553 ( .A(n7726), .B(n6320), .ZN(n7721) );
  OR2_X1 U5554 ( .A1(n6474), .A2(n6473), .ZN(n4618) );
  AOI21_X1 U5555 ( .B1(n6311), .B2(n6310), .A(n6341), .ZN(n6314) );
  NOR2_X1 U5556 ( .A1(n6538), .A2(n6539), .ZN(n9818) );
  NAND2_X1 U5557 ( .A1(n9832), .A2(n4392), .ZN(n9845) );
  NAND2_X1 U5558 ( .A1(n9845), .A2(n9844), .ZN(n9843) );
  NAND2_X1 U5559 ( .A1(n6611), .A2(n4421), .ZN(n6612) );
  OR2_X1 U5560 ( .A1(n6620), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n4421) );
  NAND2_X1 U5561 ( .A1(n6612), .A2(n6613), .ZN(n6775) );
  AND2_X1 U5562 ( .A1(n6770), .A2(n6769), .ZN(n7050) );
  AOI21_X1 U5563 ( .B1(P1_REG1_REG_17__SCAN_IN), .B2(n9039), .A(n9038), .ZN(
        n9865) );
  NOR2_X1 U5564 ( .A1(n9072), .A2(n9060), .ZN(n5607) );
  NOR2_X1 U5565 ( .A1(n9089), .A2(n4638), .ZN(n9054) );
  AOI21_X1 U5566 ( .B1(n9078), .B2(n9070), .A(n8883), .ZN(n5601) );
  OR2_X1 U5567 ( .A1(n9089), .A2(n9299), .ZN(n9072) );
  AOI21_X1 U5568 ( .B1(n9084), .B2(n8819), .A(n8879), .ZN(n9078) );
  NAND2_X1 U5569 ( .A1(n9079), .A2(n9925), .ZN(n4698) );
  NAND2_X1 U5570 ( .A1(n4448), .A2(n4447), .ZN(n9083) );
  AOI21_X1 U5571 ( .B1(n4450), .B2(n4765), .A(n4365), .ZN(n4447) );
  AOI21_X1 U5572 ( .B1(n4452), .B2(n4764), .A(n4451), .ZN(n4450) );
  INV_X1 U5573 ( .A(n4680), .ZN(n9084) );
  OAI21_X1 U5574 ( .B1(n9137), .B2(n4684), .A(n4681), .ZN(n4680) );
  NAND2_X1 U5575 ( .A1(n8962), .A2(n4685), .ZN(n4684) );
  INV_X1 U5576 ( .A(n4682), .ZN(n4681) );
  NOR2_X1 U5577 ( .A1(n9130), .A2(n9120), .ZN(n9123) );
  OR2_X1 U5578 ( .A1(n9149), .A2(n9319), .ZN(n9130) );
  AND2_X1 U5579 ( .A1(n9231), .A2(n4333), .ZN(n9167) );
  NAND2_X1 U5580 ( .A1(n4430), .A2(n4429), .ZN(n9161) );
  INV_X1 U5581 ( .A(n9164), .ZN(n4429) );
  AND2_X1 U5582 ( .A1(n8898), .A2(n8897), .ZN(n9175) );
  NAND2_X1 U5583 ( .A1(n4432), .A2(n4431), .ZN(n9192) );
  INV_X1 U5584 ( .A(n8989), .ZN(n9197) );
  NAND2_X1 U5585 ( .A1(n5253), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5289) );
  OR2_X1 U5586 ( .A1(n5289), .A2(n5288), .ZN(n5291) );
  INV_X1 U5587 ( .A(n8990), .ZN(n9230) );
  AND2_X1 U5588 ( .A1(n8858), .A2(n8857), .ZN(n4692) );
  INV_X1 U5589 ( .A(n8899), .ZN(n9227) );
  AND2_X1 U5590 ( .A1(n8857), .A2(n8862), .ZN(n9258) );
  NOR2_X1 U5591 ( .A1(n9740), .A2(n4635), .ZN(n7581) );
  INV_X1 U5592 ( .A(n4637), .ZN(n4635) );
  NAND2_X1 U5593 ( .A1(n5150), .A2(n8726), .ZN(n7477) );
  NOR2_X1 U5594 ( .A1(n9740), .A2(n7540), .ZN(n7516) );
  NAND2_X1 U5595 ( .A1(n9723), .A2(n5571), .ZN(n7480) );
  NAND2_X1 U5596 ( .A1(n7480), .A2(n8914), .ZN(n7479) );
  OR2_X1 U5597 ( .A1(n9739), .A2(n9738), .ZN(n9740) );
  OR2_X1 U5598 ( .A1(n5129), .A2(n7383), .ZN(n5144) );
  INV_X1 U5599 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5143) );
  NAND2_X1 U5600 ( .A1(n9876), .A2(n9683), .ZN(n9739) );
  NOR2_X1 U5601 ( .A1(n7199), .A2(n9875), .ZN(n9876) );
  INV_X1 U5602 ( .A(n4633), .ZN(n7305) );
  NAND2_X1 U5603 ( .A1(n6838), .A2(n4344), .ZN(n7080) );
  AND2_X1 U5604 ( .A1(n8701), .A2(n8835), .ZN(n8904) );
  CLKBUF_X1 U5605 ( .A(n6842), .Z(n7084) );
  NAND2_X1 U5606 ( .A1(n8841), .A2(n8839), .ZN(n8902) );
  NOR2_X1 U5607 ( .A1(n6853), .A2(n6935), .ZN(n6852) );
  INV_X1 U5608 ( .A(n9000), .ZN(n6741) );
  CLKBUF_X1 U5609 ( .A(n6604), .Z(n8941) );
  AND2_X1 U5610 ( .A1(n7092), .A2(n4738), .ZN(n6601) );
  NAND2_X1 U5611 ( .A1(n9941), .A2(n9926), .ZN(n4738) );
  NOR2_X1 U5612 ( .A1(n9941), .A2(n9930), .ZN(n7098) );
  AND2_X1 U5613 ( .A1(n6454), .A2(n9930), .ZN(n7093) );
  NAND2_X1 U5614 ( .A1(n5556), .A2(n7093), .ZN(n7092) );
  INV_X1 U5615 ( .A(n9887), .ZN(n9925) );
  NOR2_X1 U5616 ( .A1(n5308), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n4518) );
  AND2_X1 U5617 ( .A1(n5600), .A2(n5599), .ZN(n9946) );
  INV_X1 U5618 ( .A(n9961), .ZN(n9942) );
  AND3_X1 U5619 ( .A1(n6785), .A2(n5614), .A3(n5613), .ZN(n5619) );
  OAI22_X1 U5620 ( .A1(n6207), .A2(P1_D_REG_0__SCAN_IN), .B1(n9429), .B2(n5546), .ZN(n6784) );
  INV_X1 U5621 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n4918) );
  XNOR2_X1 U5622 ( .A(n7867), .B(n7866), .ZN(n8790) );
  XNOR2_X1 U5623 ( .A(n7848), .B(n7847), .ZN(n8578) );
  XNOR2_X1 U5624 ( .A(n5479), .B(n5478), .ZN(n8581) );
  XNOR2_X1 U5625 ( .A(n5459), .B(n5458), .ZN(n6067) );
  NAND2_X1 U5626 ( .A1(n4780), .A2(n4784), .ZN(n5459) );
  OR2_X1 U5627 ( .A1(n5425), .A2(n4787), .ZN(n4780) );
  NAND2_X1 U5628 ( .A1(n4788), .A2(n5423), .ZN(n5442) );
  OR2_X1 U5629 ( .A1(n5425), .A2(n5424), .ZN(n4788) );
  INV_X1 U5630 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5524) );
  NAND2_X1 U5631 ( .A1(n4798), .A2(n5240), .ZN(n5263) );
  NAND2_X1 U5632 ( .A1(n4593), .A2(n5106), .ZN(n5117) );
  NAND2_X1 U5633 ( .A1(n5085), .A2(n4597), .ZN(n4593) );
  NAND2_X1 U5634 ( .A1(n5085), .A2(n5084), .ZN(n5104) );
  INV_X1 U5635 ( .A(n5033), .ZN(n4566) );
  AOI21_X1 U5636 ( .B1(n10091), .B2(n9443), .A(n10089), .ZN(n9444) );
  AND2_X1 U5637 ( .A1(n4420), .A2(n5763), .ZN(n4711) );
  AND2_X1 U5638 ( .A1(n6157), .A2(n7836), .ZN(n4577) );
  OR2_X1 U5639 ( .A1(n6052), .A2(n4575), .ZN(n4574) );
  OR2_X1 U5640 ( .A1(n6051), .A2(n4575), .ZN(n4567) );
  AND2_X1 U5641 ( .A1(n4572), .A2(n4569), .ZN(n4568) );
  OR3_X1 U5642 ( .A1(n6157), .A2(n7836), .A3(n6066), .ZN(n4572) );
  NOR2_X1 U5643 ( .A1(n4571), .A2(n4570), .ZN(n4569) );
  INV_X1 U5644 ( .A(n4576), .ZN(n4571) );
  NAND2_X1 U5645 ( .A1(n4734), .A2(n5881), .ZN(n7464) );
  OR2_X1 U5646 ( .A1(n5695), .A2(n5694), .ZN(n5696) );
  INV_X1 U5647 ( .A(n4728), .ZN(n4727) );
  NAND2_X1 U5648 ( .A1(n7758), .A2(n4583), .ZN(n4589) );
  NAND2_X1 U5649 ( .A1(n4702), .A2(n4705), .ZN(n7257) );
  AND2_X1 U5650 ( .A1(n4700), .A2(n4701), .ZN(n7256) );
  NAND2_X1 U5651 ( .A1(n7011), .A2(n4704), .ZN(n4702) );
  NAND2_X1 U5652 ( .A1(n7763), .A2(n8441), .ZN(n7827) );
  OR2_X1 U5653 ( .A1(n5764), .A2(n6183), .ZN(n5730) );
  OR2_X1 U5654 ( .A1(n5933), .A2(n5932), .ZN(n5934) );
  NAND2_X1 U5655 ( .A1(n6436), .A2(n6437), .ZN(n4735) );
  INV_X1 U5656 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n9616) );
  NAND2_X1 U5657 ( .A1(n6218), .A2(n7981), .ZN(n4599) );
  XNOR2_X1 U5658 ( .A(n5695), .B(n5694), .ZN(n6483) );
  NAND2_X1 U5659 ( .A1(n7763), .A2(n8440), .ZN(n7826) );
  AND2_X1 U5660 ( .A1(n4714), .A2(n4322), .ZN(n6662) );
  AND2_X1 U5661 ( .A1(n6052), .A2(n6051), .ZN(n7833) );
  AND2_X1 U5662 ( .A1(n6057), .A2(n6073), .ZN(n8281) );
  NAND2_X1 U5663 ( .A1(n6442), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7825) );
  INV_X1 U5664 ( .A(n7843), .ZN(n7830) );
  INV_X2 U5665 ( .A(P2_U3966), .ZN(n8085) );
  NAND2_X1 U5666 ( .A1(n4402), .A2(n6592), .ZN(n6798) );
  NOR2_X1 U5667 ( .A1(n6824), .A2(n6823), .ZN(n6826) );
  NOR2_X1 U5668 ( .A1(n7218), .A2(n7217), .ZN(n7223) );
  AND2_X1 U5669 ( .A1(n6242), .A2(n6241), .ZN(n9980) );
  NAND2_X1 U5670 ( .A1(n4419), .A2(n4418), .ZN(n8169) );
  NAND2_X1 U5671 ( .A1(n8168), .A2(n8182), .ZN(n4418) );
  INV_X1 U5672 ( .A(n8187), .ZN(n4419) );
  NAND2_X1 U5673 ( .A1(n7863), .A2(n7862), .ZN(n9692) );
  NAND2_X1 U5674 ( .A1(n4860), .A2(n4858), .ZN(n8227) );
  AOI21_X1 U5675 ( .B1(n4863), .B2(n8244), .A(n4859), .ZN(n4858) );
  NAND2_X1 U5676 ( .A1(n4437), .A2(n4435), .ZN(n8465) );
  INV_X1 U5677 ( .A(n4436), .ZN(n4435) );
  NAND2_X1 U5678 ( .A1(n4438), .A2(n8411), .ZN(n4437) );
  OAI22_X1 U5679 ( .A1(n8263), .A2(n8326), .B1(n8231), .B2(n8230), .ZN(n4436)
         );
  NOR2_X1 U5680 ( .A1(n8259), .A2(n8050), .ZN(n8245) );
  NAND2_X1 U5681 ( .A1(n4864), .A2(n4868), .ZN(n8254) );
  INV_X1 U5682 ( .A(n4867), .ZN(n4865) );
  NOR2_X1 U5683 ( .A1(n4872), .A2(n4321), .ZN(n8310) );
  INV_X1 U5684 ( .A(n4874), .ZN(n4872) );
  AND2_X1 U5685 ( .A1(n4833), .A2(n4347), .ZN(n8303) );
  NAND2_X1 U5686 ( .A1(n4877), .A2(n4882), .ZN(n8334) );
  INV_X1 U5687 ( .A(n4881), .ZN(n4877) );
  NOR2_X1 U5688 ( .A1(n4881), .A2(n4878), .ZN(n8498) );
  INV_X1 U5689 ( .A(n4833), .ZN(n8319) );
  NAND2_X1 U5690 ( .A1(n4820), .A2(n4821), .ZN(n8372) );
  INV_X1 U5691 ( .A(n8283), .ZN(n8425) );
  NAND2_X1 U5692 ( .A1(n7444), .A2(n7932), .ZN(n7496) );
  NAND2_X1 U5693 ( .A1(n7122), .A2(n7121), .ZN(n7125) );
  NAND2_X1 U5694 ( .A1(n6916), .A2(n7897), .ZN(n7027) );
  NAND2_X1 U5695 ( .A1(n6567), .A2(n6566), .ZN(n6626) );
  NAND2_X1 U5696 ( .A1(n6752), .A2(n7872), .ZN(n6631) );
  INV_X1 U5697 ( .A(n6512), .ZN(n6686) );
  NAND2_X1 U5698 ( .A1(n8422), .A2(n6651), .ZN(n8455) );
  OR2_X1 U5699 ( .A1(n7845), .A2(n6649), .ZN(n8426) );
  INV_X1 U5700 ( .A(n8455), .ZN(n8430) );
  INV_X1 U5701 ( .A(n8332), .ZN(n8461) );
  NOR3_X1 U5702 ( .A1(n4674), .A2(n9691), .A3(n4673), .ZN(n9701) );
  AND2_X1 U5703 ( .A1(n9692), .A2(n9693), .ZN(n4673) );
  NOR2_X1 U5704 ( .A1(n9690), .A2(n8524), .ZN(n4674) );
  NAND2_X1 U5705 ( .A1(n6300), .A2(n6679), .ZN(n10036) );
  AND2_X1 U5706 ( .A1(n6187), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9998) );
  XNOR2_X1 U5707 ( .A(n6099), .B(P2_IR_REG_25__SCAN_IN), .ZN(n7504) );
  XNOR2_X1 U5708 ( .A(n6104), .B(P2_IR_REG_24__SCAN_IN), .ZN(n7475) );
  INV_X1 U5709 ( .A(n8054), .ZN(n7874) );
  AND2_X1 U5710 ( .A1(n5904), .A2(n5887), .ZN(n7108) );
  XNOR2_X1 U5711 ( .A(n5659), .B(P2_IR_REG_1__SCAN_IN), .ZN(n9662) );
  BUF_X1 U5712 ( .A(P2_IR_REG_0__SCAN_IN), .Z(n9990) );
  INV_X1 U5713 ( .A(n4512), .ZN(n4508) );
  NAND2_X1 U5714 ( .A1(n4514), .A2(n7704), .ZN(n4511) );
  NAND2_X1 U5715 ( .A1(n7599), .A2(n7600), .ZN(n8592) );
  AND2_X1 U5716 ( .A1(n8686), .A2(n4914), .ZN(n4916) );
  NOR2_X1 U5717 ( .A1(n7732), .A2(n4348), .ZN(n4914) );
  AND2_X1 U5718 ( .A1(n7740), .A2(n9717), .ZN(n7741) );
  NAND2_X1 U5719 ( .A1(n6874), .A2(n6873), .ZN(n6967) );
  INV_X1 U5720 ( .A(n6871), .ZN(n6874) );
  INV_X1 U5721 ( .A(n4909), .ZN(n4908) );
  NAND2_X1 U5722 ( .A1(n5286), .A2(n5285), .ZN(n9351) );
  NAND2_X1 U5723 ( .A1(n7657), .A2(n4900), .ZN(n8665) );
  NAND2_X1 U5724 ( .A1(n7657), .A2(n7656), .ZN(n4904) );
  XNOR2_X1 U5725 ( .A(n7661), .B(n7736), .ZN(n8668) );
  INV_X1 U5726 ( .A(n9729), .ZN(n9888) );
  NAND2_X1 U5727 ( .A1(n4517), .A2(n4361), .ZN(n7531) );
  INV_X1 U5728 ( .A(n9707), .ZN(n8689) );
  NAND2_X1 U5729 ( .A1(n4515), .A2(n4514), .ZN(n8686) );
  AND2_X1 U5730 ( .A1(n4515), .A2(n4350), .ZN(n8685) );
  AND2_X1 U5731 ( .A1(n6896), .A2(n6895), .ZN(n9722) );
  INV_X1 U5732 ( .A(n8982), .ZN(n4464) );
  NAND2_X1 U5733 ( .A1(n5457), .A2(n5456), .ZN(n8985) );
  NAND2_X1 U5734 ( .A1(n5440), .A2(n5439), .ZN(n9080) );
  NAND2_X1 U5735 ( .A1(n5422), .A2(n5421), .ZN(n9117) );
  OR2_X1 U5736 ( .A1(n9104), .A2(n5486), .ZN(n5422) );
  NAND2_X1 U5737 ( .A1(n5386), .A2(n5385), .ZN(n9118) );
  NAND4_X1 U5738 ( .A1(n4970), .A2(n4969), .A3(n4968), .A4(n4967), .ZN(n9002)
         );
  NOR2_X1 U5739 ( .A1(n9800), .A2(n9799), .ZN(n9798) );
  AOI21_X1 U5740 ( .B1(n6328), .B2(n6308), .A(n6468), .ZN(n9812) );
  NAND2_X1 U5741 ( .A1(n4616), .A2(n4326), .ZN(n9806) );
  AND2_X1 U5742 ( .A1(n4618), .A2(n4617), .ZN(n9807) );
  NOR2_X1 U5743 ( .A1(n4318), .A2(n6348), .ZN(n6347) );
  AND2_X1 U5744 ( .A1(n4931), .A2(n4677), .ZN(n4444) );
  AND2_X1 U5745 ( .A1(n6332), .A2(n6331), .ZN(n6538) );
  AND2_X1 U5746 ( .A1(n6619), .A2(n4394), .ZN(n6621) );
  NAND2_X1 U5747 ( .A1(n7057), .A2(n4422), .ZN(n7061) );
  OR2_X1 U5748 ( .A1(n7058), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n4422) );
  INV_X1 U5749 ( .A(n4614), .ZN(n9004) );
  NOR2_X1 U5750 ( .A1(n9011), .A2(n9010), .ZN(n9013) );
  OAI21_X1 U5751 ( .B1(n7293), .B2(n4612), .A(n4611), .ZN(n9024) );
  NAND2_X1 U5752 ( .A1(n4615), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n4612) );
  NAND2_X1 U5753 ( .A1(n9005), .A2(n4615), .ZN(n4611) );
  INV_X1 U5754 ( .A(n9007), .ZN(n4615) );
  INV_X1 U5755 ( .A(n9005), .ZN(n4613) );
  INV_X1 U5756 ( .A(n4623), .ZN(n9034) );
  INV_X1 U5757 ( .A(n4621), .ZN(n9863) );
  AND2_X1 U5758 ( .A1(n6304), .A2(n4317), .ZN(n9860) );
  NOR2_X1 U5759 ( .A1(n9873), .A2(n9047), .ZN(n4607) );
  INV_X1 U5760 ( .A(n9046), .ZN(n4606) );
  NOR2_X1 U5761 ( .A1(n9048), .A2(n9263), .ZN(n9286) );
  AND2_X1 U5762 ( .A1(n5517), .A2(n5516), .ZN(n9296) );
  XNOR2_X1 U5763 ( .A(n4745), .B(n8927), .ZN(n9297) );
  NAND2_X1 U5764 ( .A1(n4740), .A2(n4739), .ZN(n4745) );
  OR2_X1 U5765 ( .A1(n4743), .A2(n4925), .ZN(n4739) );
  OR2_X1 U5766 ( .A1(n5596), .A2(n5595), .ZN(n9069) );
  AND2_X1 U5767 ( .A1(n4744), .A2(n4743), .ZN(n5596) );
  AOI21_X1 U5768 ( .B1(n4744), .B2(n4345), .A(n8925), .ZN(n5595) );
  NAND2_X1 U5769 ( .A1(n9071), .A2(n9077), .ZN(n4744) );
  OAI21_X1 U5770 ( .B1(n4410), .B2(n9732), .A(n4401), .ZN(n9308) );
  XNOR2_X1 U5771 ( .A(n9109), .B(n9108), .ZN(n4410) );
  OR2_X1 U5772 ( .A1(n9138), .A2(n9889), .ZN(n4408) );
  NAND2_X1 U5773 ( .A1(n4449), .A2(n4764), .ZN(n9099) );
  NAND2_X1 U5774 ( .A1(n5586), .A2(n4453), .ZN(n4449) );
  NAND2_X1 U5775 ( .A1(n4763), .A2(n4769), .ZN(n9113) );
  NAND2_X1 U5776 ( .A1(n9147), .A2(n4772), .ZN(n4763) );
  NAND2_X1 U5777 ( .A1(n4774), .A2(n4776), .ZN(n9129) );
  NAND2_X1 U5778 ( .A1(n4775), .A2(n4339), .ZN(n4774) );
  INV_X1 U5779 ( .A(n9147), .ZN(n4775) );
  NAND2_X1 U5780 ( .A1(n5313), .A2(n5312), .ZN(n9341) );
  NAND2_X1 U5781 ( .A1(n4441), .A2(n4442), .ZN(n9191) );
  OR2_X1 U5782 ( .A1(n5583), .A2(n9205), .ZN(n4441) );
  INV_X1 U5783 ( .A(n4748), .ZN(n9240) );
  AOI21_X1 U5784 ( .B1(n4752), .B2(n4750), .A(n4320), .ZN(n4748) );
  NAND2_X1 U5785 ( .A1(n4693), .A2(n8857), .ZN(n9242) );
  NAND2_X1 U5786 ( .A1(n7510), .A2(n8720), .ZN(n7575) );
  NAND2_X1 U5787 ( .A1(n5575), .A2(n5574), .ZN(n7580) );
  NAND2_X1 U5788 ( .A1(n5569), .A2(n5568), .ZN(n9725) );
  NAND2_X1 U5789 ( .A1(n4691), .A2(n8911), .ZN(n7398) );
  NAND2_X1 U5790 ( .A1(n5128), .A2(n5127), .ZN(n7408) );
  NAND2_X1 U5791 ( .A1(n7303), .A2(n5564), .ZN(n7191) );
  NAND2_X1 U5792 ( .A1(n4689), .A2(n8706), .ZN(n7312) );
  INV_X1 U5793 ( .A(n9253), .ZN(n9277) );
  AND2_X2 U5794 ( .A1(n5619), .A2(n9409), .ZN(n9978) );
  AND2_X1 U5795 ( .A1(n9290), .A2(n9289), .ZN(n9371) );
  INV_X1 U5796 ( .A(n9092), .ZN(n9379) );
  AND2_X1 U5797 ( .A1(n9313), .A2(n4433), .ZN(n9381) );
  AOI21_X1 U5798 ( .B1(n9315), .B2(n9957), .A(n9314), .ZN(n4433) );
  INV_X1 U5799 ( .A(n7231), .ZN(n6901) );
  AND2_X2 U5800 ( .A1(n5619), .A2(n6784), .ZN(n9968) );
  AND2_X1 U5801 ( .A1(n6450), .A2(n5528), .ZN(n9408) );
  INV_X1 U5802 ( .A(n4948), .ZN(n9418) );
  INV_X1 U5803 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5522) );
  INV_X1 U5804 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7368) );
  INV_X1 U5805 ( .A(n8979), .ZN(n8813) );
  INV_X1 U5806 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7171) );
  INV_X1 U5807 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7118) );
  INV_X1 U5808 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6597) );
  AND2_X1 U5809 ( .A1(n5165), .A2(n5203), .ZN(n6776) );
  INV_X1 U5810 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6221) );
  INV_X1 U5811 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6186) );
  AND2_X1 U5812 ( .A1(n4982), .A2(n4999), .ZN(n9792) );
  XNOR2_X1 U5813 ( .A(n4624), .B(P1_IR_REG_1__SCAN_IN), .ZN(n7726) );
  NAND2_X1 U5814 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n4624) );
  NOR2_X1 U5815 ( .A1(n9454), .A2(n10077), .ZN(n10076) );
  AOI21_X1 U5816 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10074), .ZN(n10073) );
  NOR2_X1 U5817 ( .A1(n10073), .A2(n10072), .ZN(n10071) );
  AOI21_X1 U5818 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10071), .ZN(n10070) );
  OAI21_X1 U5819 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10068), .ZN(n10066) );
  OR2_X1 U5820 ( .A1(n8069), .A2(n8068), .ZN(n4414) );
  NAND2_X1 U5821 ( .A1(n8976), .A2(n4464), .ZN(n4463) );
  NOR2_X1 U5822 ( .A1(n4607), .A2(n4606), .ZN(n4605) );
  NAND2_X1 U5823 ( .A1(n4609), .A2(n9911), .ZN(n4608) );
  OAI21_X1 U5824 ( .B1(n9301), .B2(n9938), .A(n4695), .ZN(n4694) );
  AOI21_X1 U5825 ( .B1(n9298), .B2(n9881), .A(n9081), .ZN(n4695) );
  NAND2_X2 U5826 ( .A1(n7865), .A2(n7864), .ZN(n7893) );
  INV_X2 U5827 ( .A(n7178), .ZN(n10022) );
  NAND2_X1 U5828 ( .A1(n4616), .A2(n4387), .ZN(n4318) );
  AND2_X1 U5829 ( .A1(n8409), .A2(n4380), .ZN(n4319) );
  AND2_X1 U5830 ( .A1(n9712), .A2(n8991), .ZN(n4320) );
  OR2_X1 U5831 ( .A1(n4875), .A2(n8216), .ZN(n4321) );
  OR2_X1 U5832 ( .A1(n9319), .A2(n9146), .ZN(n8866) );
  NAND2_X1 U5833 ( .A1(n5744), .A2(n5743), .ZN(n4322) );
  AND2_X1 U5834 ( .A1(n4442), .A2(n4352), .ZN(n4323) );
  INV_X1 U5835 ( .A(n8263), .ZN(n4777) );
  AND2_X1 U5836 ( .A1(n4794), .A2(n5282), .ZN(n4324) );
  OR3_X1 U5837 ( .A1(n9089), .A2(n4638), .A3(n9053), .ZN(n4325) );
  AND2_X1 U5838 ( .A1(n8687), .A2(n4350), .ZN(n4514) );
  OR2_X1 U5839 ( .A1(n9808), .A2(n4617), .ZN(n4326) );
  AND2_X1 U5840 ( .A1(n4626), .A2(n4928), .ZN(n4327) );
  AND2_X1 U5841 ( .A1(n8911), .A2(n8714), .ZN(n4328) );
  INV_X1 U5842 ( .A(n4765), .ZN(n4764) );
  OAI21_X1 U5843 ( .B1(n5589), .B2(n4766), .A(n5588), .ZN(n4765) );
  OR2_X1 U5844 ( .A1(n8476), .A2(n8224), .ZN(n4329) );
  NAND2_X1 U5845 ( .A1(n6014), .A2(n6013), .ZN(n8329) );
  AND2_X1 U5846 ( .A1(n7992), .A2(n7893), .ZN(n4330) );
  NAND2_X1 U5847 ( .A1(n5830), .A2(n5829), .ZN(n5831) );
  INV_X1 U5848 ( .A(n5831), .ZN(n4601) );
  AND3_X1 U5849 ( .A1(n4627), .A2(n4921), .A3(n4626), .ZN(n4331) );
  AND2_X1 U5850 ( .A1(n8658), .A2(n4890), .ZN(n4332) );
  INV_X1 U5851 ( .A(n7901), .ZN(n4839) );
  AND2_X1 U5852 ( .A1(n4629), .A2(n4628), .ZN(n4333) );
  AND2_X1 U5853 ( .A1(n5654), .A2(n4888), .ZN(n4334) );
  AND2_X1 U5854 ( .A1(n5565), .A2(n5564), .ZN(n4335) );
  NAND2_X1 U5855 ( .A1(n8813), .A2(n9920), .ZN(n8805) );
  NAND2_X1 U5856 ( .A1(n7531), .A2(n7530), .ZN(n7532) );
  OR2_X1 U5857 ( .A1(n9740), .A2(n4636), .ZN(n4336) );
  OR2_X1 U5858 ( .A1(n7599), .A2(n7600), .ZN(n4337) );
  OAI21_X1 U5859 ( .B1(n6932), .B2(n6931), .A(n6930), .ZN(n6945) );
  OAI21_X1 U5860 ( .B1(n7011), .B2(n7010), .A(n5831), .ZN(n7162) );
  NAND2_X1 U5861 ( .A1(n4732), .A2(n5797), .ZN(n6984) );
  AND2_X1 U5862 ( .A1(n4730), .A2(n4729), .ZN(n6488) );
  NAND2_X1 U5863 ( .A1(n5575), .A2(n4753), .ZN(n4752) );
  AND2_X1 U5864 ( .A1(n4701), .A2(n5864), .ZN(n4338) );
  XNOR2_X1 U5865 ( .A(n8476), .B(n8246), .ZN(n8261) );
  OR2_X1 U5866 ( .A1(n9137), .A2(n9136), .ZN(n4687) );
  OR2_X1 U5867 ( .A1(n8514), .A2(n7957), .ZN(n8044) );
  NAND2_X1 U5868 ( .A1(n9152), .A2(n8987), .ZN(n4339) );
  AND2_X1 U5869 ( .A1(n4338), .A2(n5876), .ZN(n4340) );
  OR2_X1 U5870 ( .A1(n6225), .A2(n5687), .ZN(n4341) );
  OR2_X1 U5871 ( .A1(n6012), .A2(n6011), .ZN(n4342) );
  XOR2_X1 U5872 ( .A(n8329), .B(n6093), .Z(n4343) );
  INV_X1 U5873 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9410) );
  AND2_X1 U5874 ( .A1(n8906), .A2(n5562), .ZN(n4344) );
  NAND2_X1 U5875 ( .A1(n4778), .A2(n4777), .ZN(n7996) );
  INV_X1 U5876 ( .A(n4721), .ZN(n4720) );
  AOI21_X1 U5877 ( .B1(n4724), .B2(n7823), .A(n4722), .ZN(n4721) );
  INV_X1 U5878 ( .A(n6170), .ZN(n4708) );
  OR2_X1 U5879 ( .A1(n9299), .A2(n8985), .ZN(n4345) );
  OR2_X1 U5880 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n9805), .ZN(n4346) );
  NAND2_X1 U5881 ( .A1(n6568), .A2(n7889), .ZN(n8011) );
  NAND2_X1 U5882 ( .A1(n4752), .A2(n5576), .ZN(n9257) );
  NAND2_X1 U5883 ( .A1(n4889), .A2(n7641), .ZN(n8657) );
  INV_X1 U5884 ( .A(n9108), .ZN(n4451) );
  NAND4_X2 U5885 ( .A1(n5693), .A2(n5692), .A3(n5691), .A4(n5690), .ZN(n8083)
         );
  INV_X1 U5886 ( .A(n8083), .ZN(n4846) );
  OR2_X1 U5887 ( .A1(n8499), .A2(n8304), .ZN(n4347) );
  INV_X1 U5888 ( .A(n9194), .ZN(n4431) );
  INV_X1 U5889 ( .A(n9136), .ZN(n4685) );
  AND2_X1 U5890 ( .A1(n7693), .A2(n7692), .ZN(n4348) );
  NAND2_X1 U5891 ( .A1(n5125), .A2(n5124), .ZN(n5309) );
  NAND2_X1 U5892 ( .A1(n5684), .A2(n6170), .ZN(n5764) );
  INV_X1 U5893 ( .A(n5764), .ZN(n4413) );
  INV_X1 U5894 ( .A(n6701), .ZN(n6492) );
  OAI211_X1 U5895 ( .C1(n5660), .C2(n6225), .A(n4710), .B(n4709), .ZN(n6701)
         );
  OR3_X1 U5896 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .A3(
        n9990), .ZN(n4349) );
  NAND2_X1 U5897 ( .A1(n7686), .A2(n7685), .ZN(n4350) );
  NAND2_X1 U5898 ( .A1(n4898), .A2(n8602), .ZN(n8648) );
  AND3_X1 U5899 ( .A1(n7888), .A2(n7966), .A3(n7887), .ZN(n4351) );
  NAND2_X1 U5900 ( .A1(n7996), .A2(n7995), .ZN(n8244) );
  OR2_X1 U5901 ( .A1(n8504), .A2(n8325), .ZN(n8047) );
  NAND2_X1 U5902 ( .A1(n5685), .A2(n4851), .ZN(n5717) );
  NAND2_X1 U5903 ( .A1(n5187), .A2(n5186), .ZN(n7561) );
  AND2_X1 U5904 ( .A1(n7973), .A2(n8049), .ZN(n8272) );
  INV_X1 U5905 ( .A(n9183), .ZN(n5548) );
  NAND2_X1 U5906 ( .A1(n5330), .A2(n5329), .ZN(n9183) );
  NAND2_X1 U5907 ( .A1(n9341), .A2(n9212), .ZN(n4352) );
  AND2_X1 U5908 ( .A1(n4850), .A2(n8261), .ZN(n4353) );
  AND2_X1 U5909 ( .A1(n4685), .A2(n9107), .ZN(n4354) );
  AND2_X1 U5910 ( .A1(n7648), .A2(n7647), .ZN(n4355) );
  AND2_X1 U5911 ( .A1(n5217), .A2(n8720), .ZN(n4356) );
  AND2_X1 U5912 ( .A1(n4687), .A2(n8866), .ZN(n4357) );
  AND2_X1 U5913 ( .A1(n5462), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n4358) );
  AND2_X1 U5914 ( .A1(n4848), .A2(n4849), .ZN(n4359) );
  NOR2_X1 U5915 ( .A1(n7998), .A2(n7997), .ZN(n8302) );
  AND2_X1 U5916 ( .A1(n7897), .A2(n7871), .ZN(n4360) );
  INV_X1 U5917 ( .A(n9219), .ZN(n9400) );
  NAND2_X1 U5918 ( .A1(n5273), .A2(n5272), .ZN(n9219) );
  AND2_X1 U5919 ( .A1(n7437), .A2(n7430), .ZN(n4361) );
  AND2_X1 U5920 ( .A1(n9319), .A2(n9118), .ZN(n4362) );
  INV_X1 U5921 ( .A(n9053), .ZN(n9373) );
  INV_X1 U5922 ( .A(n4879), .ZN(n4878) );
  NOR2_X1 U5923 ( .A1(n8333), .A2(n4880), .ZN(n4879) );
  NOR2_X1 U5924 ( .A1(n7903), .A2(n7893), .ZN(n4363) );
  NOR2_X1 U5925 ( .A1(n9341), .A2(n9212), .ZN(n4364) );
  NOR2_X1 U5926 ( .A1(n9310), .A2(n9117), .ZN(n4365) );
  AND2_X1 U5927 ( .A1(n6948), .A2(n6947), .ZN(n4366) );
  AND2_X1 U5928 ( .A1(n7338), .A2(n8074), .ZN(n4367) );
  INV_X1 U5929 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n4954) );
  AND2_X1 U5930 ( .A1(n8658), .A2(n4891), .ZN(n4368) );
  AND2_X1 U5931 ( .A1(n8014), .A2(n7898), .ZN(n4369) );
  AND2_X1 U5932 ( .A1(n8211), .A2(n8210), .ZN(n4370) );
  AND2_X1 U5933 ( .A1(n4653), .A2(n8043), .ZN(n4371) );
  INV_X1 U5934 ( .A(n4670), .ZN(n4669) );
  NAND2_X1 U5935 ( .A1(n4671), .A2(n4672), .ZN(n4670) );
  OR2_X1 U5936 ( .A1(n5549), .A2(n9088), .ZN(n8820) );
  OR2_X1 U5937 ( .A1(n8469), .A2(n8468), .ZN(n4372) );
  INV_X1 U5938 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n5124) );
  OR2_X1 U5939 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .ZN(
        n4373) );
  AND2_X1 U5940 ( .A1(n8273), .A2(n7970), .ZN(n8291) );
  NAND2_X1 U5941 ( .A1(n8849), .A2(n8912), .ZN(n4374) );
  INV_X1 U5942 ( .A(n4585), .ZN(n4582) );
  NAND2_X1 U5943 ( .A1(n4586), .A2(n4587), .ZN(n4585) );
  INV_X1 U5944 ( .A(n7996), .ZN(n8051) );
  AND2_X1 U5945 ( .A1(n4537), .A2(n8044), .ZN(n4375) );
  NAND2_X1 U5946 ( .A1(n5911), .A2(n5910), .ZN(n5919) );
  NAND2_X1 U5947 ( .A1(n8044), .A2(n8001), .ZN(n4376) );
  INV_X1 U5948 ( .A(n8038), .ZN(n8025) );
  AND2_X1 U5949 ( .A1(n7945), .A2(n7944), .ZN(n8038) );
  OR2_X1 U5950 ( .A1(n4332), .A2(n4355), .ZN(n4377) );
  NAND2_X1 U5951 ( .A1(n8381), .A2(n4822), .ZN(n4378) );
  OR2_X1 U5952 ( .A1(n4868), .A2(n8253), .ZN(n4379) );
  NAND2_X1 U5953 ( .A1(n8534), .A2(n8415), .ZN(n4380) );
  AND2_X1 U5954 ( .A1(n6170), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4381) );
  AND2_X1 U5955 ( .A1(n7258), .A2(n4704), .ZN(n4382) );
  NAND2_X1 U5956 ( .A1(n5907), .A2(n5906), .ZN(n8539) );
  AND2_X1 U5957 ( .A1(n8920), .A2(n4749), .ZN(n4383) );
  OR2_X1 U5958 ( .A1(n9808), .A2(n6473), .ZN(n4384) );
  AND2_X1 U5959 ( .A1(n5047), .A2(SI_5_), .ZN(n4385) );
  AND2_X1 U5960 ( .A1(n4930), .A2(n6566), .ZN(n4386) );
  AND2_X1 U5961 ( .A1(n4326), .A2(n4346), .ZN(n4387) );
  INV_X1 U5962 ( .A(n8221), .ZN(n4871) );
  NOR2_X1 U5963 ( .A1(n8488), .A2(n8305), .ZN(n8221) );
  AND2_X1 U5964 ( .A1(n7996), .A2(n4850), .ZN(n4388) );
  AND2_X1 U5965 ( .A1(n4657), .A2(n4656), .ZN(n4389) );
  INV_X1 U5966 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n4888) );
  INV_X1 U5967 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n4459) );
  AND2_X1 U5968 ( .A1(n4445), .A2(n4444), .ZN(n4390) );
  NAND2_X1 U5969 ( .A1(n6000), .A2(n5999), .ZN(n8504) );
  INV_X1 U5970 ( .A(n8504), .ZN(n4671) );
  INV_X1 U5971 ( .A(n7662), .ZN(n4903) );
  AND2_X1 U5972 ( .A1(n8384), .A2(n4669), .ZN(n4391) );
  OR2_X1 U5973 ( .A1(n9831), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n4392) );
  AND2_X1 U5974 ( .A1(n6351), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n4393) );
  NAND2_X1 U5975 ( .A1(n7758), .A2(n5973), .ZN(n7807) );
  NAND2_X1 U5976 ( .A1(n7371), .A2(n7370), .ZN(n7429) );
  NAND2_X1 U5977 ( .A1(n5583), .A2(n5582), .ZN(n9204) );
  NAND2_X1 U5978 ( .A1(n4589), .A2(n4587), .ZN(n7768) );
  NAND2_X1 U5979 ( .A1(n4779), .A2(n6083), .ZN(n8471) );
  INV_X1 U5980 ( .A(n8471), .ZN(n4778) );
  NAND2_X1 U5981 ( .A1(n5096), .A2(n5095), .ZN(n7357) );
  OR2_X1 U5982 ( .A1(n7329), .A2(n7331), .ZN(n7371) );
  OR2_X1 U5983 ( .A1(n6620), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n4394) );
  NAND2_X1 U5984 ( .A1(n4517), .A2(n7430), .ZN(n7435) );
  OR2_X1 U5985 ( .A1(n8884), .A2(n8799), .ZN(n4395) );
  NAND2_X1 U5986 ( .A1(n8716), .A2(n8911), .ZN(n4396) );
  INV_X1 U5987 ( .A(n4772), .ZN(n4771) );
  NOR2_X1 U5988 ( .A1(n5587), .A2(n4773), .ZN(n4772) );
  NAND2_X1 U5989 ( .A1(n9231), .A2(n4631), .ZN(n4632) );
  INV_X1 U5990 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n4757) );
  AND2_X1 U5991 ( .A1(n4614), .A2(n4613), .ZN(n4397) );
  AND2_X1 U5992 ( .A1(n5570), .A2(n5568), .ZN(n4398) );
  AND2_X1 U5993 ( .A1(n9219), .A2(n8990), .ZN(n4399) );
  AND2_X1 U5994 ( .A1(n5266), .A2(SI_17_), .ZN(n4400) );
  INV_X1 U5995 ( .A(n4754), .ZN(n4753) );
  OR2_X1 U5996 ( .A1(n5577), .A2(n4755), .ZN(n4754) );
  AND2_X1 U5997 ( .A1(n4409), .A2(n4408), .ZN(n4401) );
  INV_X1 U5998 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n4406) );
  INV_X1 U5999 ( .A(n7835), .ZN(n4570) );
  NAND2_X1 U6000 ( .A1(n5342), .A2(n5341), .ZN(n9328) );
  INV_X1 U6001 ( .A(n9328), .ZN(n4628) );
  NAND2_X1 U6002 ( .A1(n4338), .A2(n4700), .ZN(n7281) );
  NAND2_X1 U6003 ( .A1(n4909), .A2(n4911), .ZN(n7067) );
  NAND2_X1 U6004 ( .A1(n7267), .A2(n7187), .ZN(n7337) );
  XNOR2_X1 U6005 ( .A(n5520), .B(n5519), .ZN(n5533) );
  NAND2_X1 U6006 ( .A1(n7080), .A2(n5563), .ZN(n7302) );
  NAND2_X1 U6007 ( .A1(n4908), .A2(n4911), .ZN(n6992) );
  NAND2_X1 U6008 ( .A1(n4714), .A2(n4713), .ZN(n6661) );
  NAND2_X1 U6009 ( .A1(n5653), .A2(n5766), .ZN(n6098) );
  AND2_X1 U6010 ( .A1(n6590), .A2(n6589), .ZN(n4402) );
  NAND2_X1 U6011 ( .A1(n4921), .A2(n4919), .ZN(n4403) );
  AND2_X1 U6012 ( .A1(n6838), .A2(n5562), .ZN(n4404) );
  INV_X1 U6013 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n4933) );
  NAND2_X1 U6014 ( .A1(n4728), .A2(n4730), .ZN(n6482) );
  OAI21_X1 U6015 ( .B1(n6482), .B2(n6483), .A(n5696), .ZN(n6436) );
  NAND2_X1 U6016 ( .A1(n4727), .A2(n4730), .ZN(n6489) );
  NAND2_X1 U6017 ( .A1(n4735), .A2(n5710), .ZN(n6417) );
  AND2_X1 U6018 ( .A1(n6294), .A2(n6293), .ZN(n8444) );
  INV_X1 U6019 ( .A(n4949), .ZN(n9415) );
  INV_X1 U6020 ( .A(n6251), .ZN(n4426) );
  OAI21_X1 U6021 ( .B1(n6170), .B2(n4406), .A(n4405), .ZN(n4995) );
  NAND2_X1 U6022 ( .A1(n5202), .A2(n5201), .ZN(n5222) );
  NAND2_X1 U6023 ( .A1(n4793), .A2(n4794), .ZN(n5283) );
  NAND2_X1 U6024 ( .A1(n4407), .A2(n8067), .ZN(n4415) );
  NAND3_X1 U6025 ( .A1(n8064), .A2(n4815), .A3(n4813), .ZN(n4407) );
  NAND2_X1 U6026 ( .A1(n4792), .A2(n4791), .ZN(n5300) );
  NAND2_X1 U6027 ( .A1(n5303), .A2(n5302), .ZN(n5322) );
  INV_X1 U6028 ( .A(n4649), .ZN(n8066) );
  NAND2_X1 U6029 ( .A1(n5388), .A2(n5387), .ZN(n5390) );
  AOI21_X1 U6030 ( .B1(n4806), .B2(n8059), .A(n4805), .ZN(n4561) );
  OAI21_X1 U6031 ( .B1(n7988), .B2(n7994), .A(n4810), .ZN(n4809) );
  AND2_X1 U6032 ( .A1(n5688), .A2(n4411), .ZN(n4845) );
  NAND2_X1 U6033 ( .A1(n4428), .A2(n4427), .ZN(n5297) );
  AOI21_X1 U6034 ( .B1(n8357), .B2(n8356), .A(n8046), .ZN(n8344) );
  NAND2_X1 U6035 ( .A1(n6753), .A2(n7890), .ZN(n4826) );
  AOI21_X1 U6036 ( .B1(n8438), .B2(n8041), .A(n8040), .ZN(n8414) );
  OAI21_X2 U6037 ( .B1(n7423), .B2(n7422), .A(n7929), .ZN(n7445) );
  INV_X1 U6038 ( .A(n6096), .ZN(n4736) );
  NAND2_X1 U6039 ( .A1(n7024), .A2(n7901), .ZN(n7122) );
  NAND2_X1 U6040 ( .A1(n4885), .A2(n4884), .ZN(n8394) );
  OAI22_X1 U6041 ( .A1(n7417), .A2(n8021), .B1(n7416), .B2(n8073), .ZN(n7448)
         );
  AOI21_X1 U6042 ( .B1(n6910), .B2(n6909), .A(n6908), .ZN(n7019) );
  NAND2_X1 U6043 ( .A1(n4415), .A2(n4414), .ZN(P2_U3244) );
  NAND2_X1 U6044 ( .A1(n5746), .A2(n4663), .ZN(n4662) );
  INV_X1 U6045 ( .A(n5045), .ZN(n4564) );
  NAND2_X1 U6046 ( .A1(n4602), .A2(n4600), .ZN(n4705) );
  XNOR2_X1 U6047 ( .A(n4417), .B(n4416), .ZN(n8192) );
  OR2_X1 U6048 ( .A1(n8186), .A2(n8187), .ZN(n4417) );
  INV_X1 U6049 ( .A(n6859), .ZN(n6860) );
  NAND2_X1 U6050 ( .A1(n6456), .A2(n6457), .ZN(n6859) );
  NAND2_X1 U6051 ( .A1(n6953), .A2(n6952), .ZN(n4911) );
  NAND2_X1 U6052 ( .A1(n5518), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5520) );
  NAND2_X1 U6053 ( .A1(n7609), .A2(n9713), .ZN(n8633) );
  NOR2_X1 U6054 ( .A1(n7588), .A2(n7587), .ZN(n7593) );
  NAND2_X1 U6055 ( .A1(n5920), .A2(n5630), .ZN(n5950) );
  NAND2_X1 U6056 ( .A1(n6816), .A2(n6817), .ZN(n4732) );
  NAND3_X1 U6057 ( .A1(n6427), .A2(n6663), .A3(n4322), .ZN(n4420) );
  NAND2_X1 U6058 ( .A1(n4604), .A2(n9920), .ZN(n4603) );
  INV_X1 U6059 ( .A(n6761), .ZN(n10008) );
  NAND2_X1 U6060 ( .A1(n4660), .A2(n5653), .ZN(n6096) );
  NAND2_X1 U6061 ( .A1(n6629), .A2(n6628), .ZN(n6910) );
  AND2_X2 U6062 ( .A1(n4424), .A2(n4423), .ZN(n8378) );
  NAND2_X1 U6063 ( .A1(n8525), .A2(n8416), .ZN(n4423) );
  OR2_X2 U6064 ( .A1(n8394), .A2(n4425), .ZN(n4424) );
  NAND2_X1 U6065 ( .A1(n8470), .A2(n4434), .ZN(n8555) );
  OR2_X1 U6066 ( .A1(n6225), .A2(n4426), .ZN(n5705) );
  NAND2_X1 U6067 ( .A1(n5062), .A2(n5061), .ZN(n5066) );
  AOI21_X2 U6068 ( .B1(n8039), .B2(n8038), .A(n8037), .ZN(n8438) );
  INV_X1 U6069 ( .A(n7897), .ZN(n4844) );
  NAND2_X1 U6070 ( .A1(n4819), .A2(n4818), .ZN(n8357) );
  INV_X1 U6071 ( .A(n4843), .ZN(n4842) );
  NAND2_X1 U6072 ( .A1(n4956), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4957) );
  NAND2_X4 U6073 ( .A1(n5508), .A2(n8977), .ZN(n5017) );
  INV_X1 U6074 ( .A(n9195), .ZN(n4432) );
  AND2_X1 U6075 ( .A1(n5002), .A2(n4679), .ZN(n4678) );
  INV_X1 U6076 ( .A(n9163), .ZN(n4430) );
  AND2_X2 U6077 ( .A1(n4921), .A2(n4327), .ZN(n4484) );
  NAND2_X1 U6078 ( .A1(n8834), .A2(n8903), .ZN(n4481) );
  NAND2_X1 U6079 ( .A1(n6604), .A2(n6599), .ZN(n4985) );
  NAND2_X1 U6080 ( .A1(n4736), .A2(n4887), .ZN(n5664) );
  NAND2_X1 U6081 ( .A1(n5583), .A2(n4323), .ZN(n4440) );
  NAND2_X1 U6082 ( .A1(n4978), .A2(n4922), .ZN(n5018) );
  AND4_X2 U6083 ( .A1(n4978), .A2(n4922), .A3(n4516), .A4(n4931), .ZN(n5067)
         );
  NOR2_X4 U6084 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n4978) );
  NAND3_X1 U6085 ( .A1(n4978), .A2(n4922), .A3(n4931), .ZN(n5020) );
  INV_X1 U6086 ( .A(n5018), .ZN(n4445) );
  NAND2_X1 U6087 ( .A1(n5586), .A2(n4450), .ZN(n4448) );
  OAI21_X1 U6088 ( .B1(n6838), .B2(n4457), .A(n4455), .ZN(n7303) );
  NAND2_X1 U6089 ( .A1(n4627), .A2(n4484), .ZN(n4956) );
  INV_X1 U6090 ( .A(n4940), .ZN(n4627) );
  NAND3_X1 U6091 ( .A1(n4627), .A2(n4458), .A3(n4921), .ZN(n4460) );
  INV_X1 U6092 ( .A(n8901), .ZN(n4461) );
  OAI21_X1 U6093 ( .B1(n4465), .B2(n4463), .A(n4462), .ZN(P1_U3240) );
  OR2_X1 U6094 ( .A1(n8981), .A2(n8980), .ZN(n4462) );
  NAND2_X1 U6095 ( .A1(n8816), .A2(n8815), .ZN(n4466) );
  NOR2_X1 U6096 ( .A1(n4468), .A2(n8929), .ZN(n4467) );
  OAI21_X1 U6097 ( .B1(n4472), .B2(n4470), .A(n4469), .ZN(n8780) );
  INV_X1 U6098 ( .A(n8768), .ZN(n4469) );
  AOI21_X1 U6099 ( .B1(n8763), .B2(n4354), .A(n4471), .ZN(n4470) );
  AOI21_X1 U6100 ( .B1(n8755), .B2(n8867), .A(n8805), .ZN(n4472) );
  NAND3_X1 U6101 ( .A1(n4475), .A2(n8718), .A3(n4473), .ZN(n8734) );
  INV_X2 U6102 ( .A(n5091), .ZN(n4921) );
  NAND2_X1 U6103 ( .A1(n4488), .A2(n6944), .ZN(n4485) );
  INV_X1 U6104 ( .A(n4489), .ZN(n5499) );
  NAND2_X1 U6105 ( .A1(n5498), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5504) );
  NAND3_X1 U6106 ( .A1(n4898), .A2(n8602), .A3(n7676), .ZN(n8649) );
  INV_X1 U6107 ( .A(n4495), .ZN(n4494) );
  NAND2_X1 U6108 ( .A1(n4495), .A2(n7669), .ZN(n8603) );
  OAI21_X2 U6109 ( .B1(n7657), .B2(n4899), .A(n4496), .ZN(n4495) );
  INV_X1 U6110 ( .A(n4901), .ZN(n4498) );
  NAND2_X1 U6111 ( .A1(n7631), .A2(n4502), .ZN(n4499) );
  NAND2_X1 U6112 ( .A1(n4499), .A2(n4500), .ZN(n8618) );
  NAND2_X1 U6113 ( .A1(n8626), .A2(n8627), .ZN(n4515) );
  OAI211_X1 U6114 ( .C1(n8626), .C2(n4511), .A(n4509), .B(n4506), .ZN(n7710)
         );
  NAND2_X1 U6115 ( .A1(n8626), .A2(n4507), .ZN(n4506) );
  NOR2_X1 U6116 ( .A1(n4508), .A2(n7704), .ZN(n4507) );
  OAI21_X1 U6117 ( .B1(n7704), .B2(n4512), .A(n4510), .ZN(n4509) );
  OAI21_X1 U6118 ( .B1(n7704), .B2(n4514), .A(n4512), .ZN(n4510) );
  NAND2_X1 U6119 ( .A1(n5125), .A2(n4518), .ZN(n4519) );
  INV_X1 U6120 ( .A(n4519), .ZN(n5497) );
  NAND3_X1 U6121 ( .A1(n6865), .A2(n6454), .A3(n6449), .ZN(n6453) );
  AND2_X4 U6122 ( .A1(n4522), .A2(n4521), .ZN(n6170) );
  NAND3_X1 U6123 ( .A1(n4522), .A2(n6278), .A3(n4521), .ZN(n4523) );
  NAND2_X1 U6124 ( .A1(n4389), .A2(n4526), .ZN(n4527) );
  NAND3_X1 U6125 ( .A1(n4551), .A2(n4548), .A3(n8022), .ZN(n4547) );
  NAND3_X1 U6126 ( .A1(n4646), .A2(n8333), .A3(n4560), .ZN(n4559) );
  NAND2_X1 U6127 ( .A1(n4563), .A2(n5919), .ZN(n7565) );
  AND3_X2 U6128 ( .A1(n4563), .A2(n5919), .A3(n4562), .ZN(n7564) );
  INV_X1 U6129 ( .A(n7566), .ZN(n4562) );
  NAND2_X1 U6130 ( .A1(n5909), .A2(n5908), .ZN(n4563) );
  NAND2_X1 U6131 ( .A1(n5034), .A2(n5033), .ZN(n5046) );
  NAND3_X1 U6132 ( .A1(n6052), .A2(n6051), .A3(n7836), .ZN(n7834) );
  NAND4_X1 U6133 ( .A1(n4573), .A2(n4574), .A3(n4568), .A4(n4567), .ZN(n6165)
         );
  NAND3_X1 U6134 ( .A1(n6052), .A2(n6051), .A3(n4577), .ZN(n4573) );
  OR2_X1 U6135 ( .A1(n6157), .A2(n6066), .ZN(n4575) );
  OAI21_X2 U6136 ( .B1(n7758), .B2(n4585), .A(n4578), .ZN(n6010) );
  NAND2_X1 U6137 ( .A1(n5085), .A2(n4594), .ZN(n4590) );
  NAND2_X1 U6138 ( .A1(n4590), .A2(n4591), .ZN(n5137) );
  MUX2_X1 U6139 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(P1_DATAO_REG_3__SCAN_IN), 
        .S(n6170), .Z(n5013) );
  NAND3_X1 U6140 ( .A1(n4608), .A2(n4605), .A3(n4603), .ZN(P1_U3260) );
  XNOR2_X1 U6141 ( .A(n9003), .B(n9009), .ZN(n7293) );
  INV_X1 U6142 ( .A(n4618), .ZN(n6472) );
  NAND2_X1 U6143 ( .A1(n6328), .A2(n6327), .ZN(n4617) );
  NAND3_X1 U6144 ( .A1(n4627), .A2(n4921), .A3(n4625), .ZN(n5521) );
  INV_X1 U6145 ( .A(n4632), .ZN(n9180) );
  INV_X1 U6146 ( .A(n4634), .ZN(n9262) );
  MUX2_X1 U6147 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(P1_DATAO_REG_1__SCAN_IN), 
        .S(n6170), .Z(n4971) );
  NAND2_X1 U6148 ( .A1(n4803), .A2(n5014), .ZN(n4643) );
  NOR2_X2 U6149 ( .A1(n8278), .A2(n8476), .ZN(n8199) );
  INV_X1 U6150 ( .A(n4662), .ZN(n4660) );
  NAND2_X1 U6151 ( .A1(n5653), .A2(n4888), .ZN(n4661) );
  OAI21_X1 U6152 ( .B1(n4661), .B2(n4662), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n4929) );
  MUX2_X1 U6153 ( .A(n9990), .B(n8591), .S(n5684), .Z(n6731) );
  NAND2_X2 U6154 ( .A1(n8202), .A2(n6149), .ZN(n5684) );
  OR2_X1 U6155 ( .A1(n6760), .A2(n6761), .ZN(n6758) );
  NAND2_X1 U6156 ( .A1(n8384), .A2(n4668), .ZN(n8327) );
  NAND2_X2 U6157 ( .A1(n8944), .A2(n8838), .ZN(n6739) );
  OR2_X2 U6158 ( .A1(n9001), .A2(n7231), .ZN(n8944) );
  AND2_X2 U6159 ( .A1(n5003), .A2(n4678), .ZN(n7231) );
  OR2_X1 U6160 ( .A1(n5060), .A2(n6176), .ZN(n4679) );
  NAND2_X2 U6161 ( .A1(n7507), .A2(n5198), .ZN(n7510) );
  NAND2_X2 U6162 ( .A1(n4689), .A2(n4688), .ZN(n7310) );
  NAND2_X1 U6163 ( .A1(n4691), .A2(n4690), .ZN(n7401) );
  NAND2_X1 U6164 ( .A1(n4693), .A2(n4692), .ZN(n5261) );
  INV_X1 U6165 ( .A(n4694), .ZN(n9082) );
  XNOR2_X1 U6166 ( .A(n9078), .B(n9077), .ZN(n4699) );
  NAND2_X1 U6167 ( .A1(n4809), .A2(n4807), .ZN(n4806) );
  NAND2_X1 U6168 ( .A1(n7011), .A2(n4382), .ZN(n4700) );
  INV_X1 U6169 ( .A(n7010), .ZN(n4706) );
  AND2_X2 U6170 ( .A1(n5684), .A2(n5462), .ZN(n5715) );
  NAND2_X1 U6172 ( .A1(n6428), .A2(n4713), .ZN(n4712) );
  NAND2_X1 U6173 ( .A1(n4712), .A2(n4711), .ZN(n6672) );
  OAI21_X1 U6174 ( .B1(n7795), .B2(n7794), .A(n4726), .ZN(n7824) );
  NAND2_X1 U6175 ( .A1(n5961), .A2(n5962), .ZN(n4725) );
  NAND2_X1 U6176 ( .A1(n5675), .A2(n5674), .ZN(n4729) );
  NAND2_X1 U6177 ( .A1(n4732), .A2(n4731), .ZN(n6985) );
  NAND3_X1 U6178 ( .A1(n4735), .A2(n5710), .A3(n5726), .ZN(n6418) );
  NAND2_X1 U6179 ( .A1(n4736), .A2(n4334), .ZN(n5657) );
  NAND2_X1 U6180 ( .A1(n4737), .A2(n5561), .ZN(n6838) );
  INV_X1 U6181 ( .A(n6839), .ZN(n4737) );
  XNOR2_X2 U6182 ( .A(n8939), .B(n6863), .ZN(n5556) );
  NAND2_X1 U6183 ( .A1(n9071), .A2(n4741), .ZN(n4740) );
  NAND2_X1 U6184 ( .A1(n4746), .A2(n4383), .ZN(n5580) );
  NAND2_X1 U6185 ( .A1(n5017), .A2(n4381), .ZN(n4761) );
  NAND2_X2 U6186 ( .A1(n4958), .A2(n4460), .ZN(n8977) );
  NAND2_X2 U6187 ( .A1(n5017), .A2(n5462), .ZN(n5060) );
  INV_X1 U6188 ( .A(n5017), .ZN(n5001) );
  NAND2_X1 U6189 ( .A1(n7303), .A2(n4335), .ZN(n7190) );
  NAND2_X1 U6190 ( .A1(n5425), .A2(n4784), .ZN(n4783) );
  OR2_X1 U6191 ( .A1(n5242), .A2(n4797), .ZN(n4793) );
  NAND2_X1 U6192 ( .A1(n5242), .A2(n4324), .ZN(n4792) );
  OR2_X1 U6193 ( .A1(n5242), .A2(n5241), .ZN(n4798) );
  NAND2_X1 U6194 ( .A1(n4997), .A2(n4996), .ZN(n5012) );
  OAI211_X1 U6195 ( .C1(n5011), .C2(n4804), .A(n4801), .B(n5031), .ZN(n5034)
         );
  NAND2_X1 U6196 ( .A1(n4997), .A2(n4802), .ZN(n4801) );
  AND2_X1 U6197 ( .A1(n5014), .A2(n4996), .ZN(n4802) );
  NAND2_X1 U6198 ( .A1(n5012), .A2(n5011), .ZN(n4803) );
  INV_X1 U6199 ( .A(n5014), .ZN(n4804) );
  OAI21_X2 U6200 ( .B1(n5351), .B2(n5350), .A(n5353), .ZN(n5369) );
  OAI21_X2 U6201 ( .B1(n5155), .B2(n5154), .A(n5153), .ZN(n5177) );
  NAND2_X1 U6202 ( .A1(n4817), .A2(n4816), .ZN(n4815) );
  XNOR2_X1 U6203 ( .A(n8062), .B(n8283), .ZN(n4817) );
  NOR2_X2 U6204 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n4851) );
  NAND3_X1 U6205 ( .A1(n4820), .A2(n8044), .A3(n4821), .ZN(n4819) );
  OAI21_X1 U6206 ( .B1(n8401), .B2(n8400), .A(n8043), .ZN(n8380) );
  NAND2_X1 U6207 ( .A1(n8400), .A2(n8043), .ZN(n4822) );
  INV_X1 U6208 ( .A(n7872), .ZN(n4825) );
  INV_X1 U6209 ( .A(n7936), .ZN(n4827) );
  NAND2_X1 U6210 ( .A1(n4827), .A2(n7932), .ZN(n4831) );
  NAND2_X1 U6211 ( .A1(n4313), .A2(n7932), .ZN(n4830) );
  OAI21_X2 U6212 ( .B1(n7445), .B2(n4831), .A(n4828), .ZN(n8039) );
  NAND2_X1 U6213 ( .A1(n8342), .A2(n8047), .ZN(n8320) );
  NOR2_X1 U6214 ( .A1(n8321), .A2(n4835), .ZN(n4834) );
  INV_X1 U6215 ( .A(n8047), .ZN(n4835) );
  OAI21_X1 U6216 ( .B1(n7901), .B2(n4841), .A(n7902), .ZN(n4837) );
  NAND2_X1 U6217 ( .A1(n4839), .A2(n7900), .ZN(n4838) );
  INV_X2 U6218 ( .A(n6724), .ZN(n6500) );
  NAND2_X1 U6219 ( .A1(n7887), .A2(n7884), .ZN(n6387) );
  NAND2_X1 U6220 ( .A1(n4846), .A2(n6724), .ZN(n7884) );
  NAND2_X1 U6221 ( .A1(n8260), .A2(n4388), .ZN(n4847) );
  NAND3_X1 U6222 ( .A1(n4851), .A2(n5685), .A3(n5624), .ZN(n5716) );
  NOR2_X4 U6223 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5685) );
  AOI21_X1 U6224 ( .B1(n8288), .B2(n4866), .A(n4863), .ZN(n8240) );
  NAND2_X1 U6225 ( .A1(n8288), .A2(n4865), .ZN(n4864) );
  AOI21_X1 U6226 ( .B1(n8288), .B2(n8222), .A(n8221), .ZN(n8270) );
  OR2_X1 U6227 ( .A1(n8504), .A2(n8359), .ZN(n4882) );
  NAND2_X1 U6228 ( .A1(n6567), .A2(n4386), .ZN(n6629) );
  NAND2_X1 U6229 ( .A1(n8435), .A2(n4319), .ZN(n4885) );
  INV_X1 U6230 ( .A(n4886), .ZN(n8434) );
  NAND3_X1 U6231 ( .A1(n7634), .A2(n8676), .A3(n4891), .ZN(n4889) );
  NAND2_X1 U6232 ( .A1(n7634), .A2(n8676), .ZN(n8611) );
  INV_X1 U6233 ( .A(n8612), .ZN(n4891) );
  AOI21_X1 U6234 ( .B1(n7599), .B2(n4896), .A(n4895), .ZN(n4892) );
  OAI21_X1 U6235 ( .B1(n7599), .B2(n4895), .A(n4893), .ZN(n9714) );
  NAND2_X1 U6236 ( .A1(n4904), .A2(n7662), .ZN(n8666) );
  NAND2_X1 U6237 ( .A1(n7329), .A2(n7370), .ZN(n4905) );
  NAND2_X1 U6238 ( .A1(n4910), .A2(n6957), .ZN(n4909) );
  AND2_X1 U6239 ( .A1(n4911), .A2(n4910), .ZN(n6956) );
  NAND2_X1 U6240 ( .A1(n7531), .A2(n4912), .ZN(n7549) );
  OAI211_X1 U6241 ( .C1(n4916), .C2(n7750), .A(n4915), .B(n7749), .ZN(P1_U3218) );
  NAND2_X1 U6242 ( .A1(n4916), .A2(n7741), .ZN(n4915) );
  NOR2_X2 U6243 ( .A1(n4956), .A2(n4917), .ZN(n4946) );
  NAND3_X1 U6244 ( .A1(n4954), .A2(n4459), .A3(n4918), .ZN(n4917) );
  OR2_X2 U6245 ( .A1(n4946), .A2(n9410), .ZN(n4943) );
  NAND2_X1 U6246 ( .A1(n4921), .A2(n4933), .ZN(n5093) );
  NOR2_X1 U6247 ( .A1(n4940), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n4919) );
  CLKBUF_X1 U6248 ( .A(n6149), .Z(n6240) );
  NAND2_X1 U6249 ( .A1(n5698), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5690) );
  NAND2_X1 U6250 ( .A1(n5698), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5670) );
  INV_X1 U6251 ( .A(n8576), .ZN(n5667) );
  INV_X1 U6252 ( .A(n5621), .ZN(n5623) );
  INV_X1 U6253 ( .A(n5615), .ZN(n5618) );
  CLKBUF_X1 U6254 ( .A(n6695), .Z(n6703) );
  NAND2_X1 U6255 ( .A1(n5664), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5665) );
  AND2_X2 U6256 ( .A1(n9415), .A2(n4948), .ZN(n4988) );
  NAND2_X1 U6257 ( .A1(n8084), .A2(n6492), .ZN(n7883) );
  OR2_X1 U6258 ( .A1(n9297), .A2(n9253), .ZN(n5593) );
  AND2_X1 U6259 ( .A1(n5746), .A2(n5652), .ZN(n5920) );
  XNOR2_X1 U6260 ( .A(n6035), .B(n6036), .ZN(n7800) );
  INV_X1 U6261 ( .A(n8530), .ZN(n8211) );
  INV_X1 U6262 ( .A(n8814), .ZN(n5503) );
  INV_X1 U6263 ( .A(n8492), .ZN(n8218) );
  AND2_X1 U6264 ( .A1(n6154), .A2(n6153), .ZN(n4923) );
  OR2_X1 U6265 ( .A1(n9296), .A2(n9938), .ZN(n4924) );
  AND2_X1 U6266 ( .A1(n9060), .A2(n9079), .ZN(n4925) );
  OR2_X1 U6267 ( .A1(n8934), .A2(n9921), .ZN(n4926) );
  NOR2_X1 U6268 ( .A1(n6794), .A2(n9896), .ZN(n8695) );
  AND2_X1 U6269 ( .A1(n7592), .A2(n7591), .ZN(n4927) );
  AND2_X1 U6270 ( .A1(n5524), .A2(n5519), .ZN(n4928) );
  INV_X1 U6271 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5661) );
  INV_X1 U6272 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n8572) );
  NAND2_X1 U6273 ( .A1(n6300), .A2(n6648), .ZN(n10046) );
  INV_X2 U6274 ( .A(n10046), .ZN(n10048) );
  INV_X1 U6275 ( .A(SI_17_), .ZN(n5265) );
  INV_X1 U6276 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5801) );
  INV_X1 U6277 ( .A(n8305), .ZN(n8220) );
  OR2_X1 U6278 ( .A1(n8080), .A2(n6627), .ZN(n4930) );
  INV_X1 U6279 ( .A(n8908), .ZN(n5071) );
  MUX2_X1 U6280 ( .A(n8778), .B(n8777), .S(n8805), .Z(n8779) );
  INV_X1 U6281 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5627) );
  INV_X1 U6282 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n4932) );
  XNOR2_X1 U6283 ( .A(n6093), .B(n6701), .ZN(n5674) );
  INV_X1 U6284 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5654) );
  NAND2_X1 U6285 ( .A1(n9294), .A2(n8799), .ZN(n8789) );
  INV_X1 U6286 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n4941) );
  INV_X1 U6287 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n5243) );
  INV_X1 U6288 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n4931) );
  INV_X1 U6289 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5912) );
  NAND2_X1 U6290 ( .A1(n8524), .A2(n8084), .ZN(n5673) );
  INV_X1 U6291 ( .A(n6002), .ZN(n6001) );
  INV_X1 U6292 ( .A(n5956), .ZN(n5954) );
  AND2_X1 U6293 ( .A1(n8467), .A2(n8247), .ZN(n8052) );
  AND2_X1 U6294 ( .A1(n7875), .A2(n7883), .ZN(n6388) );
  INV_X1 U6295 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5935) );
  INV_X1 U6296 ( .A(n6954), .ZN(n6952) );
  INV_X1 U6297 ( .A(n5255), .ZN(n5253) );
  INV_X1 U6298 ( .A(n9726), .ZN(n5570) );
  NOR2_X1 U6299 ( .A1(n6454), .A2(n8900), .ZN(n8901) );
  INV_X1 U6300 ( .A(SI_23_), .ZN(n9614) );
  INV_X1 U6301 ( .A(SI_20_), .ZN(n9595) );
  INV_X1 U6302 ( .A(SI_16_), .ZN(n9613) );
  INV_X1 U6303 ( .A(SI_12_), .ZN(n5158) );
  INV_X1 U6304 ( .A(SI_9_), .ZN(n9527) );
  INV_X1 U6305 ( .A(n7465), .ZN(n5902) );
  OR2_X1 U6306 ( .A1(n5779), .A2(n5778), .ZN(n5780) );
  INV_X1 U6307 ( .A(n6027), .ZN(n6026) );
  OR2_X1 U6308 ( .A1(n6015), .A2(n9502), .ZN(n6027) );
  NAND2_X1 U6309 ( .A1(n5987), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n6002) );
  NAND2_X1 U6310 ( .A1(n5820), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5839) );
  INV_X1 U6311 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5655) );
  INV_X1 U6312 ( .A(n8439), .ZN(n8210) );
  INV_X1 U6313 ( .A(n8016), .ZN(n7123) );
  INV_X1 U6314 ( .A(n8426), .ZN(n8452) );
  OR2_X1 U6315 ( .A1(n10022), .A2(n8425), .ZN(n6649) );
  INV_X1 U6316 ( .A(n6872), .ZN(n6873) );
  INV_X1 U6317 ( .A(n8651), .ZN(n7676) );
  AND2_X1 U6318 ( .A1(n5189), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n5210) );
  OR2_X1 U6319 ( .A1(n5395), .A2(n5394), .ZN(n5416) );
  OR2_X1 U6320 ( .A1(n5331), .A2(n8659), .ZN(n5343) );
  OR2_X1 U6321 ( .A1(n5098), .A2(n5097), .ZN(n5129) );
  AND2_X1 U6322 ( .A1(n8983), .A2(n9049), .ZN(n5515) );
  OR2_X1 U6323 ( .A1(n5267), .A2(P1_IR_REG_16__SCAN_IN), .ZN(n5268) );
  INV_X1 U6324 ( .A(SI_11_), .ZN(n9522) );
  NAND2_X1 U6325 ( .A1(n6026), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6056) );
  INV_X1 U6326 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n9500) );
  AND2_X1 U6327 ( .A1(n6084), .A2(n6074), .ZN(n8256) );
  OR2_X1 U6328 ( .A1(n5974), .A2(n9616), .ZN(n5988) );
  INV_X1 U6329 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n9590) );
  INV_X1 U6330 ( .A(n8413), .ZN(n8409) );
  INV_X1 U6331 ( .A(n8076), .ZN(n7266) );
  OR2_X1 U6332 ( .A1(n6681), .A2(n6648), .ZN(n6650) );
  INV_X1 U6333 ( .A(n8329), .ZN(n8499) );
  AND2_X1 U6334 ( .A1(n8034), .A2(n8425), .ZN(n6147) );
  INV_X1 U6335 ( .A(n8440), .ZN(n8324) );
  AND2_X1 U6336 ( .A1(n9991), .A2(n9993), .ZN(n6117) );
  INV_X1 U6337 ( .A(n5636), .ZN(n6124) );
  NAND2_X1 U6338 ( .A1(n7377), .A2(n7378), .ZN(n7428) );
  INV_X1 U6339 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n5233) );
  OR2_X1 U6340 ( .A1(n5343), .A2(n8620), .ZN(n5362) );
  INV_X1 U6341 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n7383) );
  OR2_X1 U6342 ( .A1(n9922), .A2(n9921), .ZN(n9908) );
  INV_X1 U6343 ( .A(n8985), .ZN(n9087) );
  INV_X1 U6344 ( .A(n9706), .ZN(n9256) );
  INV_X1 U6345 ( .A(n8913), .ZN(n5135) );
  NAND2_X1 U6346 ( .A1(n8797), .A2(n8796), .ZN(n8803) );
  AND2_X1 U6347 ( .A1(n9908), .A2(n5616), .ZN(n9961) );
  OR2_X1 U6348 ( .A1(n8810), .A2(n4317), .ZN(n9889) );
  OR2_X1 U6349 ( .A1(n9945), .A2(n8814), .ZN(n5613) );
  NAND2_X1 U6350 ( .A1(n5390), .A2(n5389), .ZN(n5402) );
  AND2_X1 U6351 ( .A1(n5264), .A2(n5247), .ZN(n5262) );
  OR2_X1 U6352 ( .A1(n5164), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n5203) );
  OAI21_X1 U6353 ( .B1(n8258), .B2(n7843), .A(n6162), .ZN(n6163) );
  INV_X1 U6354 ( .A(n7825), .ZN(n7840) );
  AND2_X1 U6355 ( .A1(n6146), .A2(n6125), .ZN(n7835) );
  AND2_X1 U6356 ( .A1(n6092), .A2(n6091), .ZN(n8263) );
  AND4_X1 U6357 ( .A1(n5918), .A2(n5917), .A3(n5916), .A4(n5915), .ZN(n7789)
         );
  INV_X1 U6358 ( .A(n9983), .ZN(n9979) );
  INV_X1 U6359 ( .A(n9981), .ZN(n9674) );
  AND2_X1 U6360 ( .A1(n8003), .A2(n8002), .ZN(n8381) );
  AND2_X1 U6361 ( .A1(n7930), .A2(n7929), .ZN(n8021) );
  INV_X1 U6362 ( .A(n8444), .ZN(n8411) );
  INV_X1 U6363 ( .A(n6679), .ZN(n6648) );
  AND2_X1 U6364 ( .A1(n8346), .A2(n8345), .ZN(n8507) );
  OR2_X1 U6365 ( .A1(n6147), .A2(n6123), .ZN(n10031) );
  OR2_X1 U6366 ( .A1(n9994), .A2(n6117), .ZN(n6679) );
  NAND2_X1 U6367 ( .A1(n7450), .A2(n10006), .ZN(n10034) );
  XNOR2_X1 U6368 ( .A(n6097), .B(P2_IR_REG_26__SCAN_IN), .ZN(n8589) );
  AND2_X1 U6369 ( .A1(n5785), .A2(n5784), .ZN(n8124) );
  OR2_X1 U6370 ( .A1(n7742), .A2(n5486), .ZN(n5476) );
  NAND2_X1 U6371 ( .A1(n6279), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5009) );
  INV_X1 U6372 ( .A(n9873), .ZN(n9854) );
  INV_X1 U6373 ( .A(n9797), .ZN(n9868) );
  INV_X1 U6374 ( .A(n9263), .ZN(n9877) );
  INV_X1 U6375 ( .A(n9077), .ZN(n9070) );
  INV_X1 U6376 ( .A(n9889), .ZN(n9730) );
  INV_X1 U6377 ( .A(n9896), .ZN(n9272) );
  AND2_X1 U6378 ( .A1(n9978), .A2(n9942), .ZN(n9284) );
  INV_X1 U6379 ( .A(n9354), .ZN(n9957) );
  AND2_X1 U6380 ( .A1(n5207), .A2(n5227), .ZN(n7295) );
  NOR2_X1 U6381 ( .A1(n9442), .A2(n9441), .ZN(n10090) );
  OAI21_X1 U6382 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10053), .ZN(n10084) );
  AND2_X1 U6383 ( .A1(n7475), .A2(n6119), .ZN(n6222) );
  INV_X1 U6384 ( .A(n8521), .ZN(n8390) );
  OR2_X1 U6385 ( .A1(n6491), .A2(n10031), .ZN(n7843) );
  NAND2_X1 U6386 ( .A1(n6080), .A2(n6079), .ZN(n8224) );
  NAND2_X1 U6387 ( .A1(n6034), .A2(n6033), .ZN(n8217) );
  OR2_X1 U6388 ( .A1(n5947), .A2(n5946), .ZN(n8439) );
  OR2_X1 U6389 ( .A1(n6229), .A2(n8585), .ZN(n9983) );
  INV_X1 U6390 ( .A(n9980), .ZN(n8191) );
  OR2_X1 U6391 ( .A1(n9992), .A2(n9991), .ZN(n9995) );
  INV_X1 U6392 ( .A(n9717), .ZN(n8683) );
  NAND2_X1 U6393 ( .A1(n5476), .A2(n5475), .ZN(n9079) );
  OR2_X1 U6394 ( .A1(P1_U3083), .A2(n6465), .ZN(n9873) );
  NAND2_X1 U6395 ( .A1(n9918), .A2(n6786), .ZN(n9899) );
  NAND2_X1 U6396 ( .A1(n9918), .A2(n9903), .ZN(n9253) );
  INV_X1 U6397 ( .A(n9284), .ZN(n9360) );
  INV_X1 U6398 ( .A(n9978), .ZN(n9975) );
  INV_X1 U6399 ( .A(n9152), .ZN(n9389) );
  INV_X1 U6400 ( .A(n9365), .ZN(n9405) );
  INV_X1 U6401 ( .A(n9968), .ZN(n9966) );
  NAND2_X1 U6402 ( .A1(n9408), .A2(n6207), .ZN(n9939) );
  INV_X1 U6403 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7543) );
  XNOR2_X1 U6404 ( .A(n5523), .B(n5522), .ZN(n7503) );
  INV_X1 U6405 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6206) );
  INV_X1 U6406 ( .A(n9428), .ZN(n7729) );
  INV_X1 U6407 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n10091) );
  NOR2_X1 U6408 ( .A1(n10076), .A2(n10075), .ZN(n10074) );
  OAI21_X1 U6409 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10065), .ZN(n10063) );
  AND2_X1 U6410 ( .A1(n6222), .A2(n9998), .ZN(P2_U3966) );
  INV_X1 U6411 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  NOR2_X1 U6412 ( .A1(n6450), .A2(n6166), .ZN(P1_U4006) );
  NAND2_X1 U6413 ( .A1(n5067), .A2(n4932), .ZN(n5091) );
  NOR2_X1 U6414 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n4936) );
  NOR2_X1 U6415 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n4935) );
  NOR2_X1 U6416 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n4934) );
  NAND4_X1 U6417 ( .A1(n4937), .A2(n4936), .A3(n4935), .A4(n4934), .ZN(n5308)
         );
  INV_X1 U6418 ( .A(n5308), .ZN(n4939) );
  NOR3_X1 U6419 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .A3(
        P1_IR_REG_22__SCAN_IN), .ZN(n4938) );
  NAND4_X1 U6420 ( .A1(n4939), .A2(n4938), .A3(n5496), .A4(n5501), .ZN(n4940)
         );
  XNOR2_X2 U6421 ( .A(n4943), .B(n4942), .ZN(n4949) );
  NAND2_X1 U6422 ( .A1(n4944), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4945) );
  MUX2_X1 U6423 ( .A(P1_IR_REG_31__SCAN_IN), .B(n4945), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n4947) );
  INV_X1 U6424 ( .A(n4946), .ZN(n9411) );
  NAND2_X1 U6425 ( .A1(n4988), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n4952) );
  NAND2_X1 U6426 ( .A1(n4987), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n4951) );
  NAND2_X1 U6427 ( .A1(n5004), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n4950) );
  NAND4_X1 U6428 ( .A1(n4953), .A2(n4952), .A3(n4951), .A4(n4950), .ZN(n6863)
         );
  MUX2_X1 U6429 ( .A(P1_IR_REG_31__SCAN_IN), .B(n4957), .S(
        P1_IR_REG_27__SCAN_IN), .Z(n4958) );
  XNOR2_X1 U6430 ( .A(n4973), .B(SI_1_), .ZN(n4972) );
  XNOR2_X1 U6431 ( .A(n4972), .B(n4971), .ZN(n7712) );
  NAND2_X1 U6432 ( .A1(n4988), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n4964) );
  NAND2_X1 U6433 ( .A1(n5005), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n4963) );
  NAND2_X1 U6434 ( .A1(n4987), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n4962) );
  NAND2_X1 U6435 ( .A1(n5004), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n4961) );
  NAND2_X1 U6436 ( .A1(n5462), .A2(SI_0_), .ZN(n4965) );
  XNOR2_X1 U6437 ( .A(n4965), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n6168) );
  INV_X1 U6438 ( .A(n9930), .ZN(n8900) );
  CLKBUF_X2 U6439 ( .A(n6863), .Z(n9926) );
  INV_X1 U6440 ( .A(n9926), .ZN(n6606) );
  NAND2_X1 U6441 ( .A1(n6606), .A2(n9941), .ZN(n4966) );
  NAND2_X1 U6442 ( .A1(n5005), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n4970) );
  NAND2_X1 U6443 ( .A1(n4988), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n4969) );
  NAND2_X1 U6444 ( .A1(n4987), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n4968) );
  NAND2_X1 U6445 ( .A1(n5004), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n4967) );
  NAND2_X1 U6446 ( .A1(n4972), .A2(n4971), .ZN(n4976) );
  INV_X1 U6447 ( .A(n4973), .ZN(n4974) );
  NAND2_X1 U6448 ( .A1(n4974), .A2(SI_1_), .ZN(n4975) );
  NAND2_X1 U6449 ( .A1(n4976), .A2(n4975), .ZN(n4994) );
  INV_X1 U6450 ( .A(SI_2_), .ZN(n4977) );
  XNOR2_X1 U6451 ( .A(n4995), .B(n4977), .ZN(n4993) );
  XNOR2_X1 U6452 ( .A(n4994), .B(n4993), .ZN(n6174) );
  NOR2_X1 U6453 ( .A1(n4978), .A2(n9410), .ZN(n4979) );
  NAND2_X1 U6454 ( .A1(n4979), .A2(P1_IR_REG_2__SCAN_IN), .ZN(n4982) );
  INV_X1 U6455 ( .A(n4979), .ZN(n4981) );
  INV_X1 U6456 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n4980) );
  NAND2_X1 U6457 ( .A1(n4981), .A2(n4980), .ZN(n4999) );
  NAND2_X1 U6458 ( .A1(n5001), .A2(n9792), .ZN(n4983) );
  OAI211_X2 U6459 ( .C1(n5060), .C2(n6174), .A(n4984), .B(n4983), .ZN(n6879)
         );
  XNOR2_X1 U6460 ( .A(n9002), .B(n6879), .ZN(n6599) );
  INV_X1 U6461 ( .A(n9002), .ZN(n8940) );
  NAND2_X1 U6462 ( .A1(n8940), .A2(n6879), .ZN(n8943) );
  NAND2_X1 U6463 ( .A1(n4985), .A2(n8943), .ZN(n8834) );
  INV_X1 U6464 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n4986) );
  NAND2_X1 U6465 ( .A1(n5005), .A2(n4986), .ZN(n4992) );
  NAND2_X1 U6466 ( .A1(n5509), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n4991) );
  NAND2_X1 U6467 ( .A1(n4988), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n4990) );
  NAND2_X1 U6468 ( .A1(n5510), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n4989) );
  NAND2_X1 U6469 ( .A1(n4994), .A2(n4993), .ZN(n4997) );
  NAND2_X1 U6470 ( .A1(n4995), .A2(SI_2_), .ZN(n4996) );
  INV_X1 U6471 ( .A(SI_3_), .ZN(n4998) );
  XNOR2_X1 U6472 ( .A(n5013), .B(n4998), .ZN(n5011) );
  XNOR2_X1 U6473 ( .A(n5012), .B(n5011), .ZN(n6176) );
  INV_X1 U6474 ( .A(n5112), .ZN(n5016) );
  NAND2_X1 U6475 ( .A1(n5016), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n5003) );
  NAND2_X1 U6476 ( .A1(n4999), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5000) );
  XNOR2_X1 U6477 ( .A(n5000), .B(P1_IR_REG_3__SCAN_IN), .ZN(n6324) );
  NAND2_X1 U6478 ( .A1(n5001), .A2(n6324), .ZN(n5002) );
  INV_X1 U6479 ( .A(n6739), .ZN(n8903) );
  NAND2_X1 U6480 ( .A1(n4308), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5010) );
  NAND2_X1 U6481 ( .A1(n6280), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5008) );
  INV_X1 U6482 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n5006) );
  XNOR2_X1 U6483 ( .A(n5006), .B(P1_REG3_REG_3__SCAN_IN), .ZN(n7247) );
  NAND2_X1 U6484 ( .A1(n5451), .A2(n7247), .ZN(n5007) );
  MUX2_X1 U6485 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n4708), .Z(n5032) );
  INV_X1 U6486 ( .A(SI_4_), .ZN(n5015) );
  XNOR2_X1 U6487 ( .A(n5032), .B(n5015), .ZN(n5031) );
  NAND2_X1 U6488 ( .A1(n5016), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n5023) );
  NAND2_X1 U6489 ( .A1(n5018), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5019) );
  MUX2_X1 U6490 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5019), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n5021) );
  AND2_X1 U6491 ( .A1(n5021), .A2(n5020), .ZN(n6478) );
  NAND2_X1 U6492 ( .A1(n5311), .A2(n6478), .ZN(n5022) );
  INV_X1 U6493 ( .A(n6935), .ZN(n7246) );
  NAND2_X1 U6494 ( .A1(n9000), .A2(n7246), .ZN(n8839) );
  NAND2_X1 U6495 ( .A1(n8697), .A2(n8841), .ZN(n6842) );
  NAND2_X1 U6496 ( .A1(n6280), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5030) );
  INV_X1 U6497 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n6329) );
  OR2_X1 U6498 ( .A1(n5489), .A2(n6329), .ZN(n5029) );
  NAND2_X1 U6499 ( .A1(n4308), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5028) );
  INV_X1 U6500 ( .A(n5038), .ZN(n5039) );
  INV_X1 U6501 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5025) );
  NAND2_X1 U6502 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n5024) );
  NAND2_X1 U6503 ( .A1(n5025), .A2(n5024), .ZN(n5026) );
  AND2_X1 U6504 ( .A1(n5039), .A2(n5026), .ZN(n9905) );
  NAND2_X1 U6505 ( .A1(n5451), .A2(n9905), .ZN(n5027) );
  NAND4_X1 U6506 ( .A1(n5030), .A2(n5029), .A3(n5028), .A4(n5027), .ZN(n8999)
         );
  INV_X1 U6507 ( .A(n8999), .ZN(n7087) );
  NAND2_X1 U6508 ( .A1(n5032), .A2(SI_4_), .ZN(n5033) );
  MUX2_X1 U6509 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n4708), .Z(n5047) );
  XNOR2_X1 U6510 ( .A(n5046), .B(n5045), .ZN(n6183) );
  INV_X2 U6511 ( .A(n5112), .ZN(n8795) );
  NAND2_X1 U6512 ( .A1(n8795), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n5037) );
  NAND2_X1 U6513 ( .A1(n5020), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5035) );
  XNOR2_X1 U6514 ( .A(n5035), .B(P1_IR_REG_5__SCAN_IN), .ZN(n9805) );
  NAND2_X1 U6515 ( .A1(n5311), .A2(n9805), .ZN(n5036) );
  OAI211_X1 U6516 ( .C1(n5060), .C2(n6183), .A(n5037), .B(n5036), .ZN(n6962)
         );
  NAND2_X1 U6517 ( .A1(n7087), .A2(n6962), .ZN(n8701) );
  INV_X1 U6518 ( .A(n8701), .ZN(n8842) );
  INV_X1 U6519 ( .A(n6962), .ZN(n9909) );
  NAND2_X1 U6520 ( .A1(n8999), .A2(n9909), .ZN(n8835) );
  OAI21_X1 U6521 ( .B1(n6842), .B2(n8842), .A(n8835), .ZN(n5052) );
  NAND2_X1 U6522 ( .A1(n6280), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5044) );
  NAND2_X1 U6523 ( .A1(n4308), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5043) );
  NAND2_X1 U6524 ( .A1(n5038), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5054) );
  INV_X1 U6525 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6344) );
  NAND2_X1 U6526 ( .A1(n5039), .A2(n6344), .ZN(n5040) );
  AND2_X1 U6527 ( .A1(n5054), .A2(n5040), .ZN(n7003) );
  NAND2_X1 U6528 ( .A1(n5451), .A2(n7003), .ZN(n5042) );
  CLKBUF_X3 U6529 ( .A(n4988), .Z(n6279) );
  NAND2_X1 U6530 ( .A1(n6279), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5041) );
  NAND4_X1 U6531 ( .A1(n5044), .A2(n5043), .A3(n5042), .A4(n5041), .ZN(n8998)
         );
  INV_X1 U6532 ( .A(n8998), .ZN(n7314) );
  INV_X1 U6533 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n5048) );
  MUX2_X1 U6534 ( .A(n5048), .B(n6186), .S(n5462), .Z(n5063) );
  XNOR2_X1 U6535 ( .A(n5063), .B(SI_6_), .ZN(n5061) );
  XNOR2_X1 U6536 ( .A(n5062), .B(n5061), .ZN(n6185) );
  NAND2_X1 U6537 ( .A1(n8795), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n5051) );
  OR2_X1 U6538 ( .A1(n4390), .A2(n9410), .ZN(n5049) );
  XNOR2_X1 U6539 ( .A(n5049), .B(P1_IR_REG_6__SCAN_IN), .ZN(n6351) );
  NAND2_X1 U6540 ( .A1(n5311), .A2(n6351), .ZN(n5050) );
  OAI211_X1 U6541 ( .C1(n5060), .C2(n6185), .A(n5051), .B(n5050), .ZN(n9276)
         );
  NAND2_X1 U6542 ( .A1(n7314), .A2(n9276), .ZN(n8949) );
  INV_X1 U6543 ( .A(n9276), .ZN(n7081) );
  NAND2_X1 U6544 ( .A1(n8998), .A2(n7081), .ZN(n8706) );
  NAND2_X1 U6545 ( .A1(n6280), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5059) );
  NAND2_X1 U6546 ( .A1(n4308), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5058) );
  NOR2_X1 U6547 ( .A1(n5054), .A2(n5053), .ZN(n5073) );
  INV_X1 U6548 ( .A(n5073), .ZN(n5074) );
  NAND2_X1 U6549 ( .A1(n5054), .A2(n5053), .ZN(n5055) );
  AND2_X1 U6550 ( .A1(n5074), .A2(n5055), .ZN(n7307) );
  NAND2_X1 U6551 ( .A1(n5451), .A2(n7307), .ZN(n5057) );
  NAND2_X1 U6552 ( .A1(n6279), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5056) );
  NAND4_X1 U6553 ( .A1(n5059), .A2(n5058), .A3(n5057), .A4(n5056), .ZN(n8997)
         );
  INV_X1 U6554 ( .A(n8997), .ZN(n7088) );
  INV_X1 U6555 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6201) );
  INV_X2 U6556 ( .A(n5060), .ZN(n5090) );
  INV_X1 U6557 ( .A(n5063), .ZN(n5064) );
  NAND2_X1 U6558 ( .A1(n5064), .A2(SI_6_), .ZN(n5065) );
  MUX2_X1 U6559 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n5462), .Z(n5083) );
  XNOR2_X1 U6560 ( .A(n5083), .B(SI_7_), .ZN(n5080) );
  XNOR2_X1 U6561 ( .A(n5082), .B(n5080), .ZN(n6193) );
  NAND2_X1 U6562 ( .A1(n5090), .A2(n6193), .ZN(n5070) );
  OR2_X1 U6563 ( .A1(n5067), .A2(n9410), .ZN(n5068) );
  XNOR2_X1 U6564 ( .A(n5068), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6548) );
  NAND2_X1 U6565 ( .A1(n5311), .A2(n6548), .ZN(n5069) );
  OAI211_X1 U6566 ( .C1(n5112), .C2(n6201), .A(n5070), .B(n5069), .ZN(n7308)
         );
  NAND2_X1 U6567 ( .A1(n7088), .A2(n7308), .ZN(n8710) );
  INV_X1 U6568 ( .A(n7308), .ZN(n9953) );
  NAND2_X1 U6569 ( .A1(n8997), .A2(n9953), .ZN(n8712) );
  NAND2_X1 U6570 ( .A1(n8710), .A2(n8712), .ZN(n8908) );
  NAND2_X1 U6571 ( .A1(n4308), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5079) );
  INV_X1 U6572 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n5072) );
  OR2_X1 U6573 ( .A1(n5489), .A2(n5072), .ZN(n5078) );
  NAND2_X1 U6574 ( .A1(n5073), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5098) );
  INV_X1 U6575 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n7153) );
  NAND2_X1 U6576 ( .A1(n5074), .A2(n7153), .ZN(n5075) );
  AND2_X1 U6577 ( .A1(n5098), .A2(n5075), .ZN(n7201) );
  NAND2_X1 U6578 ( .A1(n5451), .A2(n7201), .ZN(n5077) );
  NAND2_X1 U6579 ( .A1(n6280), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5076) );
  NAND4_X1 U6580 ( .A1(n5079), .A2(n5078), .A3(n5077), .A4(n5076), .ZN(n8996)
         );
  INV_X1 U6581 ( .A(n8996), .ZN(n9890) );
  INV_X1 U6582 ( .A(n5080), .ZN(n5081) );
  NAND2_X1 U6583 ( .A1(n5083), .A2(SI_7_), .ZN(n5084) );
  INV_X1 U6584 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n5086) );
  MUX2_X1 U6585 ( .A(n5086), .B(n6206), .S(n4708), .Z(n5087) );
  NAND2_X1 U6586 ( .A1(n5087), .A2(n9496), .ZN(n5106) );
  INV_X1 U6587 ( .A(n5087), .ZN(n5088) );
  NAND2_X1 U6588 ( .A1(n5088), .A2(SI_8_), .ZN(n5089) );
  NAND2_X1 U6589 ( .A1(n5106), .A2(n5089), .ZN(n5105) );
  XNOR2_X1 U6590 ( .A(n5104), .B(n5105), .ZN(n6203) );
  NAND2_X1 U6591 ( .A1(n6203), .A2(n5090), .ZN(n5096) );
  NAND2_X1 U6592 ( .A1(n5091), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5092) );
  MUX2_X1 U6593 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5092), .S(
        P1_IR_REG_8__SCAN_IN), .Z(n5094) );
  AND2_X1 U6594 ( .A1(n5094), .A2(n5093), .ZN(n9821) );
  AOI22_X1 U6595 ( .A1(n8795), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n5311), .B2(
        n9821), .ZN(n5095) );
  NAND2_X1 U6596 ( .A1(n9890), .A2(n7357), .ZN(n8714) );
  AND2_X1 U6597 ( .A1(n8710), .A2(n8714), .ZN(n8828) );
  NAND2_X1 U6598 ( .A1(n7310), .A2(n8828), .ZN(n9883) );
  NAND2_X1 U6599 ( .A1(n5098), .A2(n5097), .ZN(n5099) );
  AND2_X1 U6600 ( .A1(n5129), .A2(n5099), .ZN(n9897) );
  NAND2_X1 U6601 ( .A1(n5451), .A2(n9897), .ZN(n5103) );
  NAND2_X1 U6602 ( .A1(n4308), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5102) );
  NAND2_X1 U6603 ( .A1(n6279), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5101) );
  NAND2_X1 U6604 ( .A1(n6280), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5100) );
  NAND4_X1 U6605 ( .A1(n5103), .A2(n5102), .A3(n5101), .A4(n5100), .ZN(n8995)
         );
  INV_X1 U6606 ( .A(n8995), .ZN(n7399) );
  INV_X1 U6607 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n5108) );
  INV_X1 U6608 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n5107) );
  MUX2_X1 U6609 ( .A(n5108), .B(n5107), .S(n5462), .Z(n5109) );
  NAND2_X1 U6610 ( .A1(n5109), .A2(n9527), .ZN(n5118) );
  INV_X1 U6611 ( .A(n5109), .ZN(n5110) );
  NAND2_X1 U6612 ( .A1(n5110), .A2(SI_9_), .ZN(n5111) );
  XNOR2_X1 U6613 ( .A(n5117), .B(n5116), .ZN(n6212) );
  NAND2_X1 U6614 ( .A1(n6212), .A2(n5090), .ZN(n5115) );
  NAND2_X1 U6615 ( .A1(n5093), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5113) );
  XNOR2_X1 U6616 ( .A(n5113), .B(P1_IR_REG_9__SCAN_IN), .ZN(n9831) );
  AOI22_X1 U6617 ( .A1(n8795), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5311), .B2(
        n9831), .ZN(n5114) );
  OR2_X1 U6618 ( .A1(n7399), .A2(n9875), .ZN(n8912) );
  INV_X1 U6619 ( .A(n7357), .ZN(n7203) );
  NAND2_X1 U6620 ( .A1(n7203), .A2(n8996), .ZN(n9884) );
  AND2_X1 U6621 ( .A1(n8912), .A2(n9884), .ZN(n8848) );
  NAND2_X1 U6622 ( .A1(n7399), .A2(n9875), .ZN(n8911) );
  MUX2_X1 U6623 ( .A(n5119), .B(n6221), .S(n5462), .Z(n5121) );
  NAND2_X1 U6624 ( .A1(n5121), .A2(n5120), .ZN(n5138) );
  INV_X1 U6625 ( .A(n5121), .ZN(n5122) );
  NAND2_X1 U6626 ( .A1(n5122), .A2(SI_10_), .ZN(n5123) );
  NAND2_X1 U6627 ( .A1(n6216), .A2(n5090), .ZN(n5128) );
  INV_X1 U6628 ( .A(n5093), .ZN(n5125) );
  NAND2_X1 U6629 ( .A1(n5309), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5126) );
  XNOR2_X1 U6630 ( .A(n5126), .B(P1_IR_REG_10__SCAN_IN), .ZN(n9853) );
  AOI22_X1 U6631 ( .A1(n8795), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5311), .B2(
        n9853), .ZN(n5127) );
  NAND2_X1 U6632 ( .A1(n4308), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5134) );
  NAND2_X1 U6633 ( .A1(n5510), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5133) );
  NAND2_X1 U6634 ( .A1(n5129), .A2(n7383), .ZN(n5130) );
  AND2_X1 U6635 ( .A1(n5144), .A2(n5130), .ZN(n7382) );
  NAND2_X1 U6636 ( .A1(n5451), .A2(n7382), .ZN(n5132) );
  NAND2_X1 U6637 ( .A1(n6279), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5131) );
  NAND4_X1 U6638 ( .A1(n5134), .A2(n5133), .A3(n5132), .A4(n5131), .ZN(n9729)
         );
  NAND2_X1 U6639 ( .A1(n7408), .A2(n9888), .ZN(n8716) );
  NAND2_X1 U6640 ( .A1(n8849), .A2(n8716), .ZN(n8913) );
  NAND2_X1 U6641 ( .A1(n7401), .A2(n8849), .ZN(n9727) );
  NAND2_X1 U6642 ( .A1(n5137), .A2(n5136), .ZN(n5139) );
  MUX2_X1 U6643 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n5462), .Z(n5152) );
  XNOR2_X1 U6644 ( .A(n5152), .B(n9522), .ZN(n5151) );
  NAND2_X1 U6645 ( .A1(n6218), .A2(n5090), .ZN(n5142) );
  NOR2_X1 U6646 ( .A1(n5309), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n5162) );
  OR2_X1 U6647 ( .A1(n5162), .A2(n9410), .ZN(n5140) );
  XNOR2_X1 U6648 ( .A(n5140), .B(P1_IR_REG_11__SCAN_IN), .ZN(n6620) );
  AOI22_X1 U6649 ( .A1(n8795), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5311), .B2(
        n6620), .ZN(n5141) );
  NAND2_X1 U6650 ( .A1(n6280), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5149) );
  NAND2_X1 U6651 ( .A1(n4308), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5148) );
  INV_X1 U6652 ( .A(n5168), .ZN(n5170) );
  NAND2_X1 U6653 ( .A1(n5144), .A2(n5143), .ZN(n5145) );
  AND2_X1 U6654 ( .A1(n5170), .A2(n5145), .ZN(n9736) );
  NAND2_X1 U6655 ( .A1(n5451), .A2(n9736), .ZN(n5147) );
  NAND2_X1 U6656 ( .A1(n6279), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5146) );
  NAND4_X1 U6657 ( .A1(n5149), .A2(n5148), .A3(n5147), .A4(n5146), .ZN(n8994)
         );
  INV_X1 U6658 ( .A(n8994), .ZN(n7538) );
  NAND2_X1 U6659 ( .A1(n9738), .A2(n7538), .ZN(n8721) );
  NAND2_X1 U6660 ( .A1(n9727), .A2(n8721), .ZN(n5150) );
  OR2_X1 U6661 ( .A1(n9738), .A2(n7538), .ZN(n8726) );
  INV_X1 U6662 ( .A(n5151), .ZN(n5154) );
  NAND2_X1 U6663 ( .A1(n5152), .A2(SI_11_), .ZN(n5153) );
  MUX2_X1 U6664 ( .A(n5157), .B(n5156), .S(n5462), .Z(n5159) );
  NAND2_X1 U6665 ( .A1(n5159), .A2(n5158), .ZN(n5179) );
  INV_X1 U6666 ( .A(n5159), .ZN(n5160) );
  NAND2_X1 U6667 ( .A1(n5160), .A2(SI_12_), .ZN(n5161) );
  NAND2_X1 U6668 ( .A1(n5179), .A2(n5161), .ZN(n5178) );
  XNOR2_X1 U6669 ( .A(n5177), .B(n5178), .ZN(n6337) );
  NAND2_X1 U6670 ( .A1(n6337), .A2(n5090), .ZN(n5167) );
  NAND2_X1 U6671 ( .A1(n5162), .A2(n4757), .ZN(n5164) );
  NAND2_X1 U6672 ( .A1(n5164), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5163) );
  MUX2_X1 U6673 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5163), .S(
        P1_IR_REG_12__SCAN_IN), .Z(n5165) );
  AOI22_X1 U6674 ( .A1(n8795), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5311), .B2(
        n6776), .ZN(n5166) );
  NAND2_X1 U6675 ( .A1(n6280), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5175) );
  NAND2_X1 U6676 ( .A1(n4308), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5174) );
  INV_X1 U6677 ( .A(n5189), .ZN(n5191) );
  INV_X1 U6678 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5169) );
  NAND2_X1 U6679 ( .A1(n5170), .A2(n5169), .ZN(n5171) );
  AND2_X1 U6680 ( .A1(n5191), .A2(n5171), .ZN(n7535) );
  NAND2_X1 U6681 ( .A1(n5451), .A2(n7535), .ZN(n5173) );
  NAND2_X1 U6682 ( .A1(n6279), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5172) );
  NAND4_X1 U6683 ( .A1(n5175), .A2(n5174), .A3(n5173), .A4(n5172), .ZN(n9728)
         );
  INV_X1 U6684 ( .A(n9728), .ZN(n7559) );
  NAND2_X1 U6685 ( .A1(n7540), .A2(n7559), .ZN(n8728) );
  NAND2_X1 U6686 ( .A1(n8729), .A2(n8728), .ZN(n8914) );
  INV_X1 U6687 ( .A(n8914), .ZN(n5176) );
  NAND2_X1 U6688 ( .A1(n7477), .A2(n5176), .ZN(n7507) );
  MUX2_X1 U6689 ( .A(n5181), .B(n5180), .S(n5462), .Z(n5182) );
  NAND2_X1 U6690 ( .A1(n5182), .A2(n9617), .ZN(n5201) );
  INV_X1 U6691 ( .A(n5182), .ZN(n5183) );
  NAND2_X1 U6692 ( .A1(n5183), .A2(SI_13_), .ZN(n5184) );
  XNOR2_X1 U6693 ( .A(n5200), .B(n5199), .ZN(n6413) );
  NAND2_X1 U6694 ( .A1(n6413), .A2(n5090), .ZN(n5187) );
  NAND2_X1 U6695 ( .A1(n5203), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5185) );
  XNOR2_X1 U6696 ( .A(n5185), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7058) );
  AOI22_X1 U6697 ( .A1(n8795), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n5311), .B2(
        n7058), .ZN(n5186) );
  NAND2_X1 U6698 ( .A1(n6280), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5196) );
  INV_X1 U6699 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n5188) );
  OR2_X1 U6700 ( .A1(n5489), .A2(n5188), .ZN(n5195) );
  NAND2_X1 U6701 ( .A1(n4308), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5194) );
  INV_X1 U6702 ( .A(n5210), .ZN(n5211) );
  INV_X1 U6703 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5190) );
  NAND2_X1 U6704 ( .A1(n5191), .A2(n5190), .ZN(n5192) );
  AND2_X1 U6705 ( .A1(n5211), .A2(n5192), .ZN(n7555) );
  NAND2_X1 U6706 ( .A1(n5451), .A2(n7555), .ZN(n5193) );
  NAND4_X1 U6707 ( .A1(n5196), .A2(n5195), .A3(n5194), .A4(n5193), .ZN(n8993)
         );
  INV_X1 U6708 ( .A(n8993), .ZN(n7576) );
  OR2_X1 U6709 ( .A1(n7561), .A2(n7576), .ZN(n8723) );
  NAND2_X1 U6710 ( .A1(n7561), .A2(n7576), .ZN(n8720) );
  NAND2_X1 U6711 ( .A1(n8723), .A2(n8720), .ZN(n7508) );
  INV_X1 U6712 ( .A(n8729), .ZN(n5197) );
  NOR2_X1 U6713 ( .A1(n7508), .A2(n5197), .ZN(n5198) );
  NAND2_X1 U6714 ( .A1(n5200), .A2(n5199), .ZN(n5202) );
  MUX2_X1 U6715 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n5462), .Z(n5219) );
  XNOR2_X1 U6716 ( .A(n5219), .B(n9533), .ZN(n5218) );
  XNOR2_X1 U6717 ( .A(n5222), .B(n5218), .ZN(n6425) );
  NAND2_X1 U6718 ( .A1(n6425), .A2(n5090), .ZN(n5209) );
  NOR2_X1 U6719 ( .A1(n5249), .A2(n9410), .ZN(n5204) );
  NAND2_X1 U6720 ( .A1(n5204), .A2(P1_IR_REG_14__SCAN_IN), .ZN(n5207) );
  INV_X1 U6721 ( .A(n5204), .ZN(n5206) );
  INV_X1 U6722 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5205) );
  NAND2_X1 U6723 ( .A1(n5206), .A2(n5205), .ZN(n5227) );
  AOI22_X1 U6724 ( .A1(n8795), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5311), .B2(
        n7295), .ZN(n5208) );
  NAND2_X1 U6725 ( .A1(n6280), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5216) );
  NAND2_X1 U6726 ( .A1(n4308), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5215) );
  INV_X1 U6727 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n7053) );
  NAND2_X1 U6728 ( .A1(n5211), .A2(n7053), .ZN(n5212) );
  AND2_X1 U6729 ( .A1(n5234), .A2(n5212), .ZN(n8595) );
  NAND2_X1 U6730 ( .A1(n5451), .A2(n8595), .ZN(n5214) );
  NAND2_X1 U6731 ( .A1(n6279), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5213) );
  NAND4_X1 U6732 ( .A1(n5216), .A2(n5215), .A3(n5214), .A4(n5213), .ZN(n8992)
         );
  INV_X1 U6733 ( .A(n8992), .ZN(n9710) );
  XNOR2_X1 U6734 ( .A(n8719), .B(n9710), .ZN(n8918) );
  INV_X1 U6735 ( .A(n8918), .ZN(n5217) );
  OR2_X1 U6736 ( .A1(n8719), .A2(n9710), .ZN(n8732) );
  INV_X1 U6737 ( .A(n5218), .ZN(n5221) );
  NAND2_X1 U6738 ( .A1(n5219), .A2(SI_14_), .ZN(n5220) );
  MUX2_X1 U6739 ( .A(n5223), .B(n6597), .S(n5462), .Z(n5224) );
  NAND2_X1 U6740 ( .A1(n5224), .A2(n9619), .ZN(n5240) );
  INV_X1 U6741 ( .A(n5224), .ZN(n5225) );
  NAND2_X1 U6742 ( .A1(n5225), .A2(SI_15_), .ZN(n5226) );
  NAND2_X1 U6743 ( .A1(n5240), .A2(n5226), .ZN(n5241) );
  XNOR2_X1 U6744 ( .A(n5242), .B(n5241), .ZN(n6564) );
  NAND2_X1 U6745 ( .A1(n6564), .A2(n5090), .ZN(n5232) );
  NAND2_X1 U6746 ( .A1(n5227), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5229) );
  INV_X1 U6747 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5228) );
  XNOR2_X1 U6748 ( .A(n5229), .B(n5228), .ZN(n9009) );
  INV_X1 U6749 ( .A(n9009), .ZN(n5230) );
  AOI22_X1 U6750 ( .A1(n5230), .A2(n5311), .B1(n8795), .B2(
        P2_DATAO_REG_15__SCAN_IN), .ZN(n5231) );
  NAND2_X1 U6751 ( .A1(n4308), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5239) );
  NAND2_X1 U6752 ( .A1(n6279), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5238) );
  NAND2_X1 U6753 ( .A1(n6280), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5237) );
  NAND2_X1 U6754 ( .A1(n5234), .A2(n5233), .ZN(n5235) );
  NAND2_X1 U6755 ( .A1(n5255), .A2(n5235), .ZN(n9721) );
  INV_X1 U6756 ( .A(n9721), .ZN(n9264) );
  NAND2_X1 U6757 ( .A1(n5451), .A2(n9264), .ZN(n5236) );
  NAND4_X1 U6758 ( .A1(n5239), .A2(n5238), .A3(n5237), .A4(n5236), .ZN(n8991)
         );
  INV_X1 U6759 ( .A(n8991), .ZN(n9245) );
  NAND2_X1 U6760 ( .A1(n9712), .A2(n9245), .ZN(n8862) );
  OR2_X1 U6761 ( .A1(n9712), .A2(n9245), .ZN(n8857) );
  MUX2_X1 U6762 ( .A(n5244), .B(n5243), .S(n5462), .Z(n5245) );
  NAND2_X1 U6763 ( .A1(n5245), .A2(n9613), .ZN(n5264) );
  INV_X1 U6764 ( .A(n5245), .ZN(n5246) );
  NAND2_X1 U6765 ( .A1(n5246), .A2(SI_16_), .ZN(n5247) );
  XNOR2_X1 U6766 ( .A(n5263), .B(n5262), .ZN(n6691) );
  NAND2_X1 U6767 ( .A1(n6691), .A2(n5090), .ZN(n5252) );
  NOR2_X1 U6768 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n5248) );
  NAND2_X1 U6769 ( .A1(n5249), .A2(n5248), .ZN(n5267) );
  NAND2_X1 U6770 ( .A1(n5267), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5250) );
  XNOR2_X1 U6771 ( .A(n5250), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9028) );
  AOI22_X1 U6772 ( .A1(n8795), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n5311), .B2(
        n9028), .ZN(n5251) );
  NAND2_X1 U6773 ( .A1(n4308), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n5260) );
  NAND2_X1 U6774 ( .A1(n6279), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5259) );
  INV_X1 U6775 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n5254) );
  NAND2_X1 U6776 ( .A1(n5255), .A2(n5254), .ZN(n5256) );
  AND2_X1 U6777 ( .A1(n5289), .A2(n5256), .ZN(n9248) );
  NAND2_X1 U6778 ( .A1(n5451), .A2(n9248), .ZN(n5258) );
  NAND2_X1 U6779 ( .A1(n6280), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5257) );
  NAND4_X1 U6780 ( .A1(n5260), .A2(n5259), .A3(n5258), .A4(n5257), .ZN(n9706)
         );
  OR2_X1 U6781 ( .A1(n9247), .A2(n9256), .ZN(n8858) );
  NAND2_X1 U6782 ( .A1(n9247), .A2(n9256), .ZN(n8825) );
  NAND2_X1 U6783 ( .A1(n5261), .A2(n8825), .ZN(n9228) );
  MUX2_X1 U6784 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .S(n5462), .Z(n5266) );
  XNOR2_X1 U6785 ( .A(n5266), .B(n5265), .ZN(n5282) );
  MUX2_X1 U6786 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n5462), .Z(n5301) );
  XNOR2_X1 U6787 ( .A(n5301), .B(SI_18_), .ZN(n5298) );
  XNOR2_X1 U6788 ( .A(n5300), .B(n5298), .ZN(n6941) );
  NAND2_X1 U6789 ( .A1(n6941), .A2(n5090), .ZN(n5273) );
  NAND2_X1 U6790 ( .A1(n5268), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5284) );
  INV_X1 U6791 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5269) );
  NAND2_X1 U6792 ( .A1(n5284), .A2(n5269), .ZN(n5270) );
  NAND2_X1 U6793 ( .A1(n5270), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5271) );
  XNOR2_X1 U6794 ( .A(n5271), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9859) );
  AOI22_X1 U6795 ( .A1(n9859), .A2(n5311), .B1(n8795), .B2(
        P2_DATAO_REG_18__SCAN_IN), .ZN(n5272) );
  NAND2_X1 U6796 ( .A1(n4308), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n5281) );
  INV_X1 U6797 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n5274) );
  OR2_X1 U6798 ( .A1(n5489), .A2(n5274), .ZN(n5280) );
  INV_X1 U6799 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n5288) );
  INV_X1 U6800 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n5276) );
  NAND2_X1 U6801 ( .A1(n5291), .A2(n5276), .ZN(n5277) );
  AND2_X1 U6802 ( .A1(n5316), .A2(n5277), .ZN(n9220) );
  NAND2_X1 U6803 ( .A1(n5451), .A2(n9220), .ZN(n5279) );
  NAND2_X1 U6804 ( .A1(n6280), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n5278) );
  NAND4_X1 U6805 ( .A1(n5281), .A2(n5280), .A3(n5279), .A4(n5278), .ZN(n8990)
         );
  NAND2_X1 U6806 ( .A1(n9219), .A2(n9230), .ZN(n8747) );
  XNOR2_X1 U6807 ( .A(n5283), .B(n5282), .ZN(n6745) );
  NAND2_X1 U6808 ( .A1(n6745), .A2(n5090), .ZN(n5286) );
  XNOR2_X1 U6809 ( .A(n5284), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9039) );
  AOI22_X1 U6810 ( .A1(n8795), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n9039), .B2(
        n5311), .ZN(n5285) );
  NAND2_X1 U6811 ( .A1(n4308), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n5295) );
  INV_X1 U6812 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n5287) );
  OR2_X1 U6813 ( .A1(n5489), .A2(n5287), .ZN(n5294) );
  NAND2_X1 U6814 ( .A1(n5289), .A2(n5288), .ZN(n5290) );
  AND2_X1 U6815 ( .A1(n5291), .A2(n5290), .ZN(n9234) );
  NAND2_X1 U6816 ( .A1(n5451), .A2(n9234), .ZN(n5293) );
  NAND2_X1 U6817 ( .A1(n6280), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5292) );
  NAND4_X1 U6818 ( .A1(n5295), .A2(n5294), .A3(n5293), .A4(n5292), .ZN(n9213)
         );
  INV_X1 U6819 ( .A(n9213), .ZN(n9244) );
  NAND2_X1 U6820 ( .A1(n9351), .A2(n9244), .ZN(n9206) );
  NAND2_X1 U6821 ( .A1(n8747), .A2(n9206), .ZN(n8827) );
  OR2_X1 U6822 ( .A1(n9219), .A2(n9230), .ZN(n8745) );
  OR2_X1 U6823 ( .A1(n9351), .A2(n9244), .ZN(n9207) );
  NAND2_X1 U6824 ( .A1(n8745), .A2(n9207), .ZN(n8871) );
  NAND2_X1 U6825 ( .A1(n8871), .A2(n8747), .ZN(n5296) );
  NAND2_X1 U6826 ( .A1(n5297), .A2(n5296), .ZN(n9195) );
  INV_X1 U6827 ( .A(n5298), .ZN(n5299) );
  NAND2_X1 U6828 ( .A1(n5300), .A2(n5299), .ZN(n5303) );
  NAND2_X1 U6829 ( .A1(n5301), .A2(SI_18_), .ZN(n5302) );
  MUX2_X1 U6830 ( .A(n5304), .B(n7118), .S(n5462), .Z(n5305) );
  INV_X1 U6831 ( .A(SI_19_), .ZN(n9632) );
  NAND2_X1 U6832 ( .A1(n5305), .A2(n9632), .ZN(n5324) );
  INV_X1 U6833 ( .A(n5305), .ZN(n5306) );
  NAND2_X1 U6834 ( .A1(n5306), .A2(SI_19_), .ZN(n5307) );
  NAND2_X1 U6835 ( .A1(n5324), .A2(n5307), .ZN(n5323) );
  XNOR2_X1 U6836 ( .A(n5322), .B(n5323), .ZN(n7048) );
  NAND2_X1 U6837 ( .A1(n7048), .A2(n5090), .ZN(n5313) );
  XNOR2_X2 U6838 ( .A(n5310), .B(P1_IR_REG_19__SCAN_IN), .ZN(n9920) );
  AOI22_X1 U6839 ( .A1(n8795), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9920), .B2(
        n5311), .ZN(n5312) );
  NAND2_X1 U6840 ( .A1(n4308), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n5321) );
  NAND2_X1 U6841 ( .A1(n6279), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n5320) );
  INV_X1 U6842 ( .A(n5316), .ZN(n5314) );
  NAND2_X1 U6843 ( .A1(n5314), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5331) );
  INV_X1 U6844 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n5315) );
  NAND2_X1 U6845 ( .A1(n5316), .A2(n5315), .ZN(n5317) );
  AND2_X1 U6846 ( .A1(n5331), .A2(n5317), .ZN(n9198) );
  NAND2_X1 U6847 ( .A1(n5451), .A2(n9198), .ZN(n5319) );
  NAND2_X1 U6848 ( .A1(n6280), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5318) );
  NAND4_X1 U6849 ( .A1(n5321), .A2(n5320), .A3(n5319), .A4(n5318), .ZN(n9212)
         );
  INV_X1 U6850 ( .A(n9212), .ZN(n9179) );
  OR2_X1 U6851 ( .A1(n9341), .A2(n9179), .ZN(n8749) );
  NAND2_X1 U6852 ( .A1(n9341), .A2(n9179), .ZN(n8822) );
  NAND2_X1 U6853 ( .A1(n8749), .A2(n8822), .ZN(n9194) );
  INV_X1 U6854 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n5325) );
  MUX2_X1 U6855 ( .A(n5325), .B(n7171), .S(n5462), .Z(n5326) );
  NAND2_X1 U6856 ( .A1(n5326), .A2(n9595), .ZN(n5339) );
  INV_X1 U6857 ( .A(n5326), .ZN(n5327) );
  NAND2_X1 U6858 ( .A1(n5327), .A2(SI_20_), .ZN(n5328) );
  XNOR2_X1 U6859 ( .A(n5338), .B(n5337), .ZN(n7160) );
  NAND2_X1 U6860 ( .A1(n7160), .A2(n5090), .ZN(n5330) );
  NAND2_X1 U6861 ( .A1(n8795), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n5329) );
  INV_X1 U6862 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n8659) );
  NAND2_X1 U6863 ( .A1(n5331), .A2(n8659), .ZN(n5332) );
  NAND2_X1 U6864 ( .A1(n5343), .A2(n5332), .ZN(n9184) );
  OR2_X1 U6865 ( .A1(n5486), .A2(n9184), .ZN(n5336) );
  NAND2_X1 U6866 ( .A1(n4308), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n5335) );
  NAND2_X1 U6867 ( .A1(n6279), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n5334) );
  NAND2_X1 U6868 ( .A1(n5510), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n5333) );
  NAND4_X1 U6869 ( .A1(n5336), .A2(n5335), .A3(n5334), .A4(n5333), .ZN(n8989)
         );
  AND2_X1 U6870 ( .A1(n9183), .A2(n9197), .ZN(n8756) );
  NAND2_X1 U6871 ( .A1(n5338), .A2(n5337), .ZN(n5340) );
  NAND2_X1 U6872 ( .A1(n5340), .A2(n5339), .ZN(n5351) );
  MUX2_X1 U6873 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n5462), .Z(n5352) );
  XNOR2_X1 U6874 ( .A(n5352), .B(n9589), .ZN(n5349) );
  XNOR2_X1 U6875 ( .A(n5351), .B(n5349), .ZN(n7169) );
  NAND2_X1 U6876 ( .A1(n7169), .A2(n5090), .ZN(n5342) );
  NAND2_X1 U6877 ( .A1(n8795), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n5341) );
  INV_X1 U6878 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n8620) );
  NAND2_X1 U6879 ( .A1(n5343), .A2(n8620), .ZN(n5344) );
  NAND2_X1 U6880 ( .A1(n5362), .A2(n5344), .ZN(n9168) );
  NAND2_X1 U6881 ( .A1(n5510), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5346) );
  NAND2_X1 U6882 ( .A1(n4308), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n5345) );
  AND2_X1 U6883 ( .A1(n5346), .A2(n5345), .ZN(n5348) );
  NAND2_X1 U6884 ( .A1(n6279), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n5347) );
  OAI211_X1 U6885 ( .C1(n9168), .C2(n5486), .A(n5348), .B(n5347), .ZN(n8988)
         );
  INV_X1 U6886 ( .A(n8988), .ZN(n9178) );
  OR2_X1 U6887 ( .A1(n9328), .A2(n9178), .ZN(n8757) );
  NAND2_X1 U6888 ( .A1(n9328), .A2(n9178), .ZN(n8758) );
  NAND2_X1 U6889 ( .A1(n8757), .A2(n8758), .ZN(n9164) );
  INV_X1 U6890 ( .A(n5349), .ZN(n5350) );
  NAND2_X1 U6891 ( .A1(n5352), .A2(SI_21_), .ZN(n5353) );
  INV_X1 U6892 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n5354) );
  MUX2_X1 U6893 ( .A(n5354), .B(n7368), .S(n5462), .Z(n5355) );
  INV_X1 U6894 ( .A(SI_22_), .ZN(n9526) );
  NAND2_X1 U6895 ( .A1(n5355), .A2(n9526), .ZN(n5367) );
  INV_X1 U6896 ( .A(n5355), .ZN(n5356) );
  NAND2_X1 U6897 ( .A1(n5356), .A2(SI_22_), .ZN(n5357) );
  NAND2_X1 U6898 ( .A1(n5367), .A2(n5357), .ZN(n5368) );
  XNOR2_X1 U6899 ( .A(n5369), .B(n5368), .ZN(n7350) );
  NAND2_X1 U6900 ( .A1(n7350), .A2(n5090), .ZN(n5359) );
  NAND2_X1 U6901 ( .A1(n8795), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n5358) );
  INV_X1 U6902 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n9154) );
  INV_X1 U6903 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n5361) );
  NAND2_X1 U6904 ( .A1(n5362), .A2(n5361), .ZN(n5363) );
  NAND2_X1 U6905 ( .A1(n5379), .A2(n5363), .ZN(n9153) );
  OR2_X1 U6906 ( .A1(n9153), .A2(n5486), .ZN(n5365) );
  AOI22_X1 U6907 ( .A1(n5510), .A2(P1_REG0_REG_22__SCAN_IN), .B1(n4308), .B2(
        P1_REG1_REG_22__SCAN_IN), .ZN(n5364) );
  OAI211_X1 U6908 ( .C1(n5489), .C2(n9154), .A(n5365), .B(n5364), .ZN(n8987)
         );
  INV_X1 U6909 ( .A(n8987), .ZN(n9166) );
  NAND2_X1 U6910 ( .A1(n9144), .A2(n8896), .ZN(n5366) );
  NAND2_X1 U6911 ( .A1(n9152), .A2(n9166), .ZN(n8895) );
  NAND2_X1 U6912 ( .A1(n5366), .A2(n8895), .ZN(n9137) );
  INV_X1 U6913 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n5371) );
  INV_X1 U6914 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n5370) );
  MUX2_X1 U6915 ( .A(n5371), .B(n5370), .S(n5462), .Z(n5372) );
  NAND2_X1 U6916 ( .A1(n5372), .A2(n9614), .ZN(n5389) );
  INV_X1 U6917 ( .A(n5372), .ZN(n5373) );
  NAND2_X1 U6918 ( .A1(n5373), .A2(SI_23_), .ZN(n5374) );
  XNOR2_X1 U6919 ( .A(n5388), .B(n5387), .ZN(n7411) );
  NAND2_X1 U6920 ( .A1(n7411), .A2(n5090), .ZN(n5376) );
  NAND2_X1 U6921 ( .A1(n8795), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n5375) );
  INV_X1 U6922 ( .A(n5379), .ZN(n5377) );
  NAND2_X1 U6923 ( .A1(n5377), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5395) );
  INV_X1 U6924 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n5378) );
  NAND2_X1 U6925 ( .A1(n5379), .A2(n5378), .ZN(n5380) );
  NAND2_X1 U6926 ( .A1(n5395), .A2(n5380), .ZN(n9132) );
  OR2_X1 U6927 ( .A1(n9132), .A2(n5486), .ZN(n5386) );
  INV_X1 U6928 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n5383) );
  NAND2_X1 U6929 ( .A1(n5510), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5382) );
  NAND2_X1 U6930 ( .A1(n4308), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n5381) );
  OAI211_X1 U6931 ( .C1(n5383), .C2(n5489), .A(n5382), .B(n5381), .ZN(n5384)
         );
  INV_X1 U6932 ( .A(n5384), .ZN(n5385) );
  INV_X1 U6933 ( .A(n9118), .ZN(n9146) );
  NAND2_X1 U6934 ( .A1(n9319), .A2(n9146), .ZN(n8765) );
  NAND2_X1 U6935 ( .A1(n8866), .A2(n8765), .ZN(n9136) );
  MUX2_X1 U6936 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(P2_DATAO_REG_24__SCAN_IN), 
        .S(n5462), .Z(n5405) );
  INV_X1 U6937 ( .A(SI_24_), .ZN(n5391) );
  XNOR2_X1 U6938 ( .A(n5405), .B(n5391), .ZN(n5403) );
  XNOR2_X1 U6939 ( .A(n5402), .B(n5403), .ZN(n7474) );
  NAND2_X1 U6940 ( .A1(n7474), .A2(n5090), .ZN(n5393) );
  NAND2_X1 U6941 ( .A1(n8795), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n5392) );
  INV_X1 U6942 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n5394) );
  NAND2_X1 U6943 ( .A1(n5395), .A2(n5394), .ZN(n5396) );
  AND2_X1 U6944 ( .A1(n5416), .A2(n5396), .ZN(n9124) );
  NAND2_X1 U6945 ( .A1(n9124), .A2(n5451), .ZN(n5401) );
  INV_X1 U6946 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n9114) );
  NAND2_X1 U6947 ( .A1(n5510), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5398) );
  NAND2_X1 U6948 ( .A1(n4308), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n5397) );
  OAI211_X1 U6949 ( .C1(n9114), .C2(n5489), .A(n5398), .B(n5397), .ZN(n5399)
         );
  INV_X1 U6950 ( .A(n5399), .ZN(n5400) );
  XNOR2_X1 U6951 ( .A(n9120), .B(n8986), .ZN(n9116) );
  INV_X1 U6952 ( .A(n5402), .ZN(n5404) );
  NAND2_X1 U6953 ( .A1(n5404), .A2(n5403), .ZN(n5407) );
  NAND2_X1 U6954 ( .A1(n5405), .A2(SI_24_), .ZN(n5406) );
  NAND2_X1 U6955 ( .A1(n5407), .A2(n5406), .ZN(n5425) );
  INV_X1 U6956 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n5408) );
  MUX2_X1 U6957 ( .A(n5408), .B(n7543), .S(n5462), .Z(n5409) );
  INV_X1 U6958 ( .A(SI_25_), .ZN(n9498) );
  NAND2_X1 U6959 ( .A1(n5409), .A2(n9498), .ZN(n5423) );
  INV_X1 U6960 ( .A(n5409), .ZN(n5410) );
  NAND2_X1 U6961 ( .A1(n5410), .A2(SI_25_), .ZN(n5411) );
  NAND2_X1 U6962 ( .A1(n5423), .A2(n5411), .ZN(n5424) );
  XNOR2_X1 U6963 ( .A(n5425), .B(n5424), .ZN(n6039) );
  NAND2_X1 U6964 ( .A1(n6039), .A2(n5090), .ZN(n5413) );
  NAND2_X1 U6965 ( .A1(n8795), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n5412) );
  INV_X1 U6966 ( .A(n5416), .ZN(n5414) );
  NAND2_X1 U6967 ( .A1(n5414), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n5433) );
  INV_X1 U6968 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n5415) );
  NAND2_X1 U6969 ( .A1(n5416), .A2(n5415), .ZN(n5417) );
  NAND2_X1 U6970 ( .A1(n5433), .A2(n5417), .ZN(n9104) );
  INV_X1 U6971 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n9103) );
  NAND2_X1 U6972 ( .A1(n4308), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n5419) );
  NAND2_X1 U6973 ( .A1(n5510), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5418) );
  OAI211_X1 U6974 ( .C1(n9103), .C2(n5489), .A(n5419), .B(n5418), .ZN(n5420)
         );
  INV_X1 U6975 ( .A(n5420), .ZN(n5421) );
  NAND2_X1 U6976 ( .A1(n5549), .A2(n9088), .ZN(n8775) );
  INV_X1 U6977 ( .A(n8986), .ZN(n9138) );
  NAND2_X1 U6978 ( .A1(n9120), .A2(n9138), .ZN(n9107) );
  AND2_X1 U6979 ( .A1(n8775), .A2(n9107), .ZN(n8962) );
  INV_X1 U6980 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n5427) );
  INV_X1 U6981 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n5426) );
  MUX2_X1 U6982 ( .A(n5427), .B(n5426), .S(n5462), .Z(n5428) );
  INV_X1 U6983 ( .A(SI_26_), .ZN(n9520) );
  NAND2_X1 U6984 ( .A1(n5428), .A2(n9520), .ZN(n5443) );
  INV_X1 U6985 ( .A(n5428), .ZN(n5429) );
  NAND2_X1 U6986 ( .A1(n5429), .A2(SI_26_), .ZN(n5430) );
  NAND2_X1 U6987 ( .A1(n8587), .A2(n5090), .ZN(n5432) );
  NAND2_X1 U6988 ( .A1(n8795), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n5431) );
  INV_X1 U6989 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n8688) );
  NAND2_X1 U6990 ( .A1(n5433), .A2(n8688), .ZN(n5434) );
  NAND2_X1 U6991 ( .A1(n9093), .A2(n5451), .ZN(n5440) );
  INV_X1 U6992 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n5437) );
  NAND2_X1 U6993 ( .A1(n5510), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5436) );
  NAND2_X1 U6994 ( .A1(n4308), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n5435) );
  OAI211_X1 U6995 ( .C1(n5437), .C2(n5489), .A(n5436), .B(n5435), .ZN(n5438)
         );
  INV_X1 U6996 ( .A(n5438), .ZN(n5439) );
  INV_X1 U6997 ( .A(n9080), .ZN(n9110) );
  OR2_X1 U6998 ( .A1(n9092), .A2(n9110), .ZN(n8819) );
  AND2_X1 U6999 ( .A1(n9092), .A2(n9110), .ZN(n8879) );
  INV_X1 U7000 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n5445) );
  INV_X1 U7001 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n5444) );
  MUX2_X1 U7002 ( .A(n5445), .B(n5444), .S(n5462), .Z(n5446) );
  INV_X1 U7003 ( .A(SI_27_), .ZN(n9536) );
  NAND2_X1 U7004 ( .A1(n5446), .A2(n9536), .ZN(n5460) );
  INV_X1 U7005 ( .A(n5446), .ZN(n5447) );
  NAND2_X1 U7006 ( .A1(n5447), .A2(SI_27_), .ZN(n5448) );
  NAND2_X1 U7007 ( .A1(n6067), .A2(n5090), .ZN(n5450) );
  NAND2_X1 U7008 ( .A1(n8795), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n5449) );
  NAND2_X2 U7009 ( .A1(n5450), .A2(n5449), .ZN(n9299) );
  XNOR2_X1 U7010 ( .A(n5467), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n9074) );
  NAND2_X1 U7011 ( .A1(n9074), .A2(n5451), .ZN(n5457) );
  INV_X1 U7012 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n5454) );
  NAND2_X1 U7013 ( .A1(n4308), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n5453) );
  NAND2_X1 U7014 ( .A1(n5510), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5452) );
  OAI211_X1 U7015 ( .C1(n5454), .C2(n5489), .A(n5453), .B(n5452), .ZN(n5455)
         );
  INV_X1 U7016 ( .A(n5455), .ZN(n5456) );
  NAND2_X1 U7017 ( .A1(n9299), .A2(n9087), .ZN(n8880) );
  INV_X1 U7018 ( .A(n8821), .ZN(n8883) );
  MUX2_X1 U7019 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n5462), .Z(n5480) );
  XNOR2_X1 U7020 ( .A(n5480), .B(n9596), .ZN(n5478) );
  NAND2_X1 U7021 ( .A1(n8581), .A2(n5090), .ZN(n5464) );
  NAND2_X1 U7022 ( .A1(n8795), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n5463) );
  INV_X1 U7023 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n5466) );
  INV_X1 U7024 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n5465) );
  OAI21_X1 U7025 ( .B1(n5467), .B2(n5466), .A(n5465), .ZN(n5470) );
  INV_X1 U7026 ( .A(n5467), .ZN(n5469) );
  AND2_X1 U7027 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n5468) );
  NAND2_X1 U7028 ( .A1(n5469), .A2(n5468), .ZN(n5551) );
  NAND2_X1 U7029 ( .A1(n5470), .A2(n5551), .ZN(n7742) );
  INV_X1 U7030 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n5473) );
  NAND2_X1 U7031 ( .A1(n5510), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5472) );
  NAND2_X1 U7032 ( .A1(n4308), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n5471) );
  OAI211_X1 U7033 ( .C1(n5473), .C2(n5489), .A(n5472), .B(n5471), .ZN(n5474)
         );
  INV_X1 U7034 ( .A(n5474), .ZN(n5475) );
  INV_X1 U7035 ( .A(n9079), .ZN(n7707) );
  NAND2_X1 U7036 ( .A1(n9060), .A2(n7707), .ZN(n8881) );
  INV_X1 U7037 ( .A(n8881), .ZN(n5477) );
  AOI21_X1 U7038 ( .B1(n5601), .B2(n8817), .A(n5477), .ZN(n5495) );
  INV_X1 U7039 ( .A(n5480), .ZN(n5481) );
  NAND2_X1 U7040 ( .A1(n5481), .A2(n9596), .ZN(n5482) );
  MUX2_X1 U7041 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .S(n5462), .Z(n7849) );
  INV_X1 U7042 ( .A(SI_29_), .ZN(n9514) );
  XNOR2_X1 U7043 ( .A(n7849), .B(n9514), .ZN(n7847) );
  NAND2_X1 U7044 ( .A1(n8578), .A2(n5090), .ZN(n5485) );
  NAND2_X1 U7045 ( .A1(n8795), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n5484) );
  OR2_X1 U7046 ( .A1(n5551), .A2(n5486), .ZN(n5493) );
  INV_X1 U7047 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n5490) );
  NAND2_X1 U7048 ( .A1(n5510), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n5488) );
  NAND2_X1 U7049 ( .A1(n4308), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n5487) );
  OAI211_X1 U7050 ( .C1(n5490), .C2(n5489), .A(n5488), .B(n5487), .ZN(n5491)
         );
  INV_X1 U7051 ( .A(n5491), .ZN(n5492) );
  NAND2_X1 U7052 ( .A1(n5493), .A2(n5492), .ZN(n8984) );
  XNOR2_X1 U7053 ( .A(n9294), .B(n8984), .ZN(n8927) );
  INV_X1 U7054 ( .A(n8927), .ZN(n5494) );
  XNOR2_X1 U7055 ( .A(n5495), .B(n5494), .ZN(n5507) );
  NAND2_X1 U7056 ( .A1(n5497), .A2(n5496), .ZN(n5498) );
  OR2_X1 U7057 ( .A1(n8813), .A2(n9911), .ZN(n5506) );
  OR2_X1 U7058 ( .A1(n5503), .A2(n9921), .ZN(n5505) );
  NAND2_X1 U7059 ( .A1(n5507), .A2(n9892), .ZN(n5517) );
  NAND2_X1 U7060 ( .A1(n4308), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n5513) );
  NAND2_X1 U7061 ( .A1(n6279), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n5512) );
  NAND2_X1 U7062 ( .A1(n5510), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n5511) );
  NAND3_X1 U7063 ( .A1(n5513), .A2(n5512), .A3(n5511), .ZN(n8983) );
  INV_X1 U7064 ( .A(n4317), .ZN(n6898) );
  INV_X1 U7065 ( .A(P1_B_REG_SCAN_IN), .ZN(n5530) );
  NOR2_X1 U7066 ( .A1(n8977), .A2(n5530), .ZN(n5514) );
  NOR2_X1 U7067 ( .A1(n9887), .A2(n5514), .ZN(n9049) );
  AOI21_X1 U7068 ( .B1(n9079), .B2(n9730), .A(n5515), .ZN(n5516) );
  OR2_X1 U7069 ( .A1(n8805), .A2(n5591), .ZN(n9945) );
  NAND2_X1 U7070 ( .A1(n5525), .A2(n5524), .ZN(n5518) );
  NAND2_X1 U7071 ( .A1(n5521), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5523) );
  NAND2_X1 U7072 ( .A1(n4403), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5526) );
  MUX2_X1 U7073 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5526), .S(
        P1_IR_REG_23__SCAN_IN), .Z(n5527) );
  NAND2_X1 U7074 ( .A1(n5527), .A2(n5521), .ZN(n6890) );
  NAND2_X1 U7075 ( .A1(n6890), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6166) );
  INV_X1 U7076 ( .A(n6166), .ZN(n5528) );
  NAND2_X1 U7077 ( .A1(n9408), .A2(n5503), .ZN(n5529) );
  NOR2_X4 U7078 ( .A1(n9945), .A2(n5529), .ZN(n9896) );
  OR2_X1 U7079 ( .A1(n8810), .A2(n5598), .ZN(n6891) );
  AND2_X1 U7080 ( .A1(n6891), .A2(n9408), .ZN(n6785) );
  NAND3_X1 U7081 ( .A1(n7545), .A2(P1_B_REG_SCAN_IN), .A3(n7503), .ZN(n5532)
         );
  INV_X1 U7082 ( .A(n7503), .ZN(n5546) );
  NAND2_X1 U7083 ( .A1(n5546), .A2(n5530), .ZN(n5531) );
  NAND2_X1 U7084 ( .A1(n5532), .A2(n5531), .ZN(n5534) );
  NOR4_X1 U7085 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n5538) );
  NOR4_X1 U7086 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n5537) );
  NOR4_X1 U7087 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5536) );
  NOR4_X1 U7088 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n5535) );
  AND4_X1 U7089 ( .A1(n5538), .A2(n5537), .A3(n5536), .A4(n5535), .ZN(n5544)
         );
  NOR2_X1 U7090 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .ZN(
        n5542) );
  NOR4_X1 U7091 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n5541) );
  NOR4_X1 U7092 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n5540) );
  NOR4_X1 U7093 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n5539) );
  AND4_X1 U7094 ( .A1(n5542), .A2(n5541), .A3(n5540), .A4(n5539), .ZN(n5543)
         );
  NAND2_X1 U7095 ( .A1(n5544), .A2(n5543), .ZN(n5609) );
  INV_X1 U7096 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n6211) );
  NOR2_X1 U7097 ( .A1(n5609), .A2(n6211), .ZN(n5545) );
  NAND2_X1 U7098 ( .A1(n5533), .A2(n7545), .ZN(n6208) );
  OAI21_X1 U7099 ( .B1(n6207), .B2(n5545), .A(n6208), .ZN(n6783) );
  INV_X1 U7100 ( .A(n6783), .ZN(n5547) );
  INV_X1 U7101 ( .A(n5533), .ZN(n9429) );
  NAND3_X1 U7102 ( .A1(n6785), .A2(n5547), .A3(n6784), .ZN(n7200) );
  INV_X1 U7103 ( .A(n6879), .ZN(n7237) );
  NAND2_X1 U7104 ( .A1(n7098), .A2(n7237), .ZN(n6738) );
  OR2_X1 U7105 ( .A1(n6738), .A2(n6901), .ZN(n6853) );
  AND2_X1 U7106 ( .A1(n6852), .A2(n9909), .ZN(n7082) );
  NAND2_X1 U7107 ( .A1(n7082), .A2(n7081), .ZN(n7304) );
  INV_X1 U7108 ( .A(n7408), .ZN(n9683) );
  INV_X1 U7109 ( .A(n7561), .ZN(n9751) );
  INV_X1 U7110 ( .A(n8719), .ZN(n9747) );
  INV_X1 U7111 ( .A(n9351), .ZN(n9237) );
  NAND2_X1 U7112 ( .A1(n9167), .A2(n9389), .ZN(n9149) );
  INV_X1 U7113 ( .A(n9310), .ZN(n9102) );
  NAND2_X1 U7114 ( .A1(n9100), .A2(n9379), .ZN(n9089) );
  INV_X1 U7115 ( .A(n5607), .ZN(n5550) );
  NAND2_X1 U7116 ( .A1(n8813), .A2(n5503), .ZN(n9922) );
  INV_X1 U7117 ( .A(n9294), .ZN(n5554) );
  AND2_X1 U7118 ( .A1(n9918), .A2(n9911), .ZN(n9233) );
  INV_X1 U7119 ( .A(n9908), .ZN(n6786) );
  INV_X1 U7120 ( .A(n5551), .ZN(n5552) );
  AOI22_X1 U7121 ( .A1(n5552), .A2(n9896), .B1(P1_REG2_REG_29__SCAN_IN), .B2(
        n9938), .ZN(n5553) );
  OAI21_X1 U7122 ( .B1(n5554), .B2(n9899), .A(n5553), .ZN(n5555) );
  AOI21_X1 U7123 ( .B1(n9293), .B2(n9233), .A(n5555), .ZN(n5594) );
  INV_X1 U7124 ( .A(n6599), .ZN(n5557) );
  NAND2_X1 U7125 ( .A1(n6601), .A2(n5557), .ZN(n6600) );
  NAND2_X1 U7126 ( .A1(n8940), .A2(n7237), .ZN(n5558) );
  NAND2_X1 U7127 ( .A1(n6600), .A2(n5558), .ZN(n6736) );
  NAND2_X1 U7128 ( .A1(n6736), .A2(n6739), .ZN(n6735) );
  INV_X1 U7129 ( .A(n9001), .ZN(n6977) );
  NAND2_X1 U7130 ( .A1(n6977), .A2(n7231), .ZN(n5559) );
  NAND2_X1 U7131 ( .A1(n6735), .A2(n5559), .ZN(n6851) );
  NAND2_X1 U7132 ( .A1(n6851), .A2(n8902), .ZN(n6850) );
  NAND2_X1 U7133 ( .A1(n6741), .A2(n7246), .ZN(n5560) );
  NAND2_X1 U7134 ( .A1(n6850), .A2(n5560), .ZN(n6839) );
  NAND2_X1 U7135 ( .A1(n8999), .A2(n6962), .ZN(n5562) );
  NAND2_X1 U7136 ( .A1(n8949), .A2(n8706), .ZN(n8906) );
  NAND2_X1 U7137 ( .A1(n7314), .A2(n7081), .ZN(n5563) );
  NAND2_X1 U7138 ( .A1(n7088), .A2(n9953), .ZN(n5564) );
  INV_X1 U7139 ( .A(n8909), .ZN(n5565) );
  NAND2_X1 U7140 ( .A1(n8996), .A2(n7357), .ZN(n5566) );
  AND2_X1 U7141 ( .A1(n9875), .A2(n8995), .ZN(n5567) );
  OR2_X1 U7142 ( .A1(n7408), .A2(n9729), .ZN(n5568) );
  XNOR2_X1 U7143 ( .A(n9738), .B(n8994), .ZN(n9726) );
  NAND2_X1 U7144 ( .A1(n9738), .A2(n8994), .ZN(n5571) );
  NAND2_X1 U7145 ( .A1(n7540), .A2(n9728), .ZN(n5572) );
  OR2_X1 U7146 ( .A1(n7561), .A2(n8993), .ZN(n5573) );
  NAND2_X1 U7147 ( .A1(n7561), .A2(n8993), .ZN(n5574) );
  AND2_X1 U7148 ( .A1(n8719), .A2(n8992), .ZN(n5577) );
  OR2_X1 U7149 ( .A1(n8719), .A2(n8992), .ZN(n5576) );
  NOR2_X1 U7150 ( .A1(n9712), .A2(n8991), .ZN(n5578) );
  NAND2_X1 U7151 ( .A1(n8858), .A2(n8825), .ZN(n8920) );
  NAND2_X1 U7152 ( .A1(n9247), .A2(n9706), .ZN(n5579) );
  NAND2_X1 U7153 ( .A1(n5580), .A2(n5579), .ZN(n9226) );
  OR2_X1 U7154 ( .A1(n9351), .A2(n9213), .ZN(n5581) );
  NAND2_X1 U7155 ( .A1(n9226), .A2(n5581), .ZN(n5583) );
  NAND2_X1 U7156 ( .A1(n9351), .A2(n9213), .ZN(n5582) );
  NAND2_X1 U7157 ( .A1(n8745), .A2(n8747), .ZN(n9209) );
  NOR2_X1 U7158 ( .A1(n9183), .A2(n8989), .ZN(n5584) );
  NAND2_X1 U7159 ( .A1(n9160), .A2(n9164), .ZN(n5586) );
  NAND2_X1 U7160 ( .A1(n9328), .A2(n8988), .ZN(n5585) );
  NOR2_X1 U7161 ( .A1(n9319), .A2(n9118), .ZN(n5587) );
  AND2_X1 U7162 ( .A1(n9120), .A2(n8986), .ZN(n5589) );
  OR2_X1 U7163 ( .A1(n9120), .A2(n8986), .ZN(n5588) );
  NAND2_X1 U7164 ( .A1(n8820), .A2(n8775), .ZN(n9108) );
  NAND2_X1 U7165 ( .A1(n9092), .A2(n9080), .ZN(n8893) );
  NAND2_X1 U7166 ( .A1(n9083), .A2(n8893), .ZN(n5590) );
  NAND2_X1 U7167 ( .A1(n8817), .A2(n8881), .ZN(n8925) );
  INV_X1 U7168 ( .A(n5592), .ZN(n5597) );
  AND2_X1 U7169 ( .A1(n5597), .A2(n7193), .ZN(n9923) );
  NOR2_X1 U7170 ( .A1(n7673), .A2(n9923), .ZN(n9903) );
  NAND3_X1 U7171 ( .A1(n4924), .A2(n5594), .A3(n5593), .ZN(P1_U3355) );
  NAND2_X1 U7172 ( .A1(n5597), .A2(n6448), .ZN(n5600) );
  OR2_X1 U7173 ( .A1(n6449), .A2(n5503), .ZN(n5599) );
  INV_X1 U7174 ( .A(n8925), .ZN(n8784) );
  XNOR2_X1 U7175 ( .A(n5601), .B(n8784), .ZN(n5602) );
  NAND2_X1 U7176 ( .A1(n5602), .A2(n9892), .ZN(n5604) );
  AOI22_X1 U7177 ( .A1(n8985), .A2(n9730), .B1(n8984), .B2(n9925), .ZN(n5603)
         );
  NAND2_X1 U7178 ( .A1(n5604), .A2(n5603), .ZN(n9067) );
  NAND2_X1 U7179 ( .A1(n9072), .A2(n9060), .ZN(n5605) );
  NAND2_X1 U7180 ( .A1(n5605), .A2(n9877), .ZN(n5606) );
  NOR2_X1 U7181 ( .A1(n5607), .A2(n5606), .ZN(n9061) );
  OAI21_X1 U7182 ( .B1(n9069), .B2(n9354), .A(n5608), .ZN(n5620) );
  INV_X1 U7183 ( .A(n6207), .ZN(n5610) );
  NAND2_X1 U7184 ( .A1(n5610), .A2(n5609), .ZN(n5612) );
  OAI21_X1 U7185 ( .B1(n6207), .B2(P1_D_REG_1__SCAN_IN), .A(n6208), .ZN(n5611)
         );
  AND2_X1 U7186 ( .A1(n5612), .A2(n5611), .ZN(n5614) );
  INV_X1 U7187 ( .A(n6784), .ZN(n9409) );
  MUX2_X1 U7188 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n5620), .S(n9978), .Z(n5615)
         );
  OR2_X1 U7189 ( .A1(n9922), .A2(n9911), .ZN(n5616) );
  NAND2_X1 U7190 ( .A1(n9060), .A2(n9284), .ZN(n5617) );
  NAND2_X1 U7191 ( .A1(n5618), .A2(n5617), .ZN(P1_U3551) );
  MUX2_X1 U7192 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n5620), .S(n9968), .Z(n5621)
         );
  AND2_X1 U7193 ( .A1(n9968), .A2(n9942), .ZN(n9365) );
  NAND2_X1 U7194 ( .A1(n9060), .A2(n9365), .ZN(n5622) );
  NAND2_X1 U7195 ( .A1(n5623), .A2(n5622), .ZN(P1_U3519) );
  NOR2_X2 U7196 ( .A1(n5716), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n5746) );
  NOR2_X1 U7197 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n5626) );
  NAND4_X1 U7198 ( .A1(n5626), .A2(n5625), .A3(n5816), .A4(n5882), .ZN(n5629)
         );
  NAND4_X1 U7199 ( .A1(n5627), .A2(n5885), .A3(n5832), .A4(n5765), .ZN(n5628)
         );
  NAND2_X1 U7200 ( .A1(n5638), .A2(n5631), .ZN(n5632) );
  INV_X1 U7201 ( .A(n5634), .ZN(n5633) );
  NAND2_X1 U7202 ( .A1(n5633), .A2(P2_IR_REG_19__SCAN_IN), .ZN(n5635) );
  NAND2_X1 U7203 ( .A1(n5634), .A2(n5647), .ZN(n5641) );
  AND2_X2 U7204 ( .A1(n5635), .A2(n5641), .ZN(n8283) );
  NAND2_X1 U7205 ( .A1(n5638), .A2(n5637), .ZN(n5639) );
  NAND2_X1 U7206 ( .A1(n5639), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5640) );
  NAND2_X4 U7207 ( .A1(n5643), .A2(n6644), .ZN(n6093) );
  NOR2_X1 U7208 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n5645) );
  NAND4_X1 U7209 ( .A1(n5645), .A2(n5644), .A3(n5935), .A4(n6120), .ZN(n5650)
         );
  INV_X1 U7210 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5648) );
  INV_X1 U7211 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5646) );
  NAND4_X1 U7212 ( .A1(n5648), .A2(n5647), .A3(n6100), .A4(n5646), .ZN(n5649)
         );
  NOR2_X1 U7213 ( .A1(n5650), .A2(n5649), .ZN(n5651) );
  MUX2_X1 U7214 ( .A(P2_IR_REG_31__SCAN_IN), .B(n4929), .S(
        P2_IR_REG_27__SCAN_IN), .Z(n5658) );
  NAND2_X1 U7215 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n9990), .ZN(n5659) );
  INV_X1 U7216 ( .A(n9662), .ZN(n5660) );
  INV_X1 U7217 ( .A(n5674), .ZN(n5672) );
  INV_X1 U7218 ( .A(n5664), .ZN(n5662) );
  NAND2_X1 U7219 ( .A1(n5662), .A2(n5661), .ZN(n8573) );
  XNOR2_X2 U7220 ( .A(n5663), .B(P2_IR_REG_30__SCAN_IN), .ZN(n8576) );
  NAND2_X1 U7221 ( .A1(n5689), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n5671) );
  NAND2_X1 U7222 ( .A1(n5699), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5669) );
  NAND2_X1 U7223 ( .A1(n5697), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5668) );
  INV_X1 U7224 ( .A(n5673), .ZN(n5675) );
  NAND2_X1 U7225 ( .A1(n4312), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5679) );
  INV_X1 U7226 ( .A(n5942), .ZN(n5689) );
  NAND2_X1 U7227 ( .A1(n5689), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5678) );
  NAND2_X1 U7228 ( .A1(n5698), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5677) );
  NAND2_X1 U7229 ( .A1(n4309), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5676) );
  NAND4_X2 U7230 ( .A1(n5679), .A2(n5678), .A3(n5677), .A4(n5676), .ZN(n8086)
         );
  INV_X1 U7231 ( .A(SI_0_), .ZN(n9633) );
  OR2_X1 U7232 ( .A1(n5462), .A2(n9633), .ZN(n5680) );
  XNOR2_X1 U7233 ( .A(n5680), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n8591) );
  NAND2_X1 U7234 ( .A1(n5681), .A2(n6731), .ZN(n5683) );
  NAND2_X1 U7235 ( .A1(n5715), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n5688) );
  OR2_X1 U7236 ( .A1(n5685), .A2(n8572), .ZN(n5686) );
  XNOR2_X1 U7237 ( .A(n5686), .B(P2_IR_REG_2__SCAN_IN), .ZN(n9673) );
  INV_X1 U7238 ( .A(n9673), .ZN(n5687) );
  XNOR2_X1 U7239 ( .A(n6724), .B(n5732), .ZN(n5695) );
  NAND2_X1 U7240 ( .A1(n4310), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5693) );
  NAND2_X1 U7241 ( .A1(n4311), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5692) );
  NAND2_X1 U7242 ( .A1(n5689), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5691) );
  NAND2_X1 U7243 ( .A1(n8083), .A2(n8524), .ZN(n5694) );
  NAND2_X1 U7244 ( .A1(n4309), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5703) );
  INV_X2 U7245 ( .A(n5750), .ZN(n6140) );
  NAND2_X1 U7246 ( .A1(n6140), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5702) );
  INV_X1 U7247 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n9605) );
  NAND2_X1 U7248 ( .A1(n6145), .A2(n9605), .ZN(n5701) );
  NAND2_X1 U7249 ( .A1(n4312), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5700) );
  NAND2_X1 U7250 ( .A1(n8082), .A2(n8524), .ZN(n5707) );
  NAND2_X1 U7251 ( .A1(n5715), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n5706) );
  NAND2_X1 U7252 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n4349), .ZN(n5704) );
  XNOR2_X1 U7253 ( .A(n5704), .B(P2_IR_REG_3__SCAN_IN), .ZN(n6251) );
  OAI211_X1 U7254 ( .C1(n5764), .C2(n6176), .A(n5706), .B(n5705), .ZN(n6761)
         );
  XNOR2_X1 U7255 ( .A(n6761), .B(n6093), .ZN(n5708) );
  XNOR2_X1 U7256 ( .A(n5707), .B(n5708), .ZN(n6437) );
  INV_X1 U7257 ( .A(n5707), .ZN(n5709) );
  NAND2_X1 U7258 ( .A1(n5709), .A2(n5708), .ZN(n5710) );
  NAND2_X1 U7259 ( .A1(n4309), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5714) );
  NAND2_X1 U7260 ( .A1(n4312), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5713) );
  INV_X1 U7261 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n9629) );
  XNOR2_X1 U7262 ( .A(n9629), .B(P2_REG3_REG_3__SCAN_IN), .ZN(n6682) );
  NAND2_X1 U7263 ( .A1(n6145), .A2(n6682), .ZN(n5712) );
  NAND2_X1 U7264 ( .A1(n6140), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5711) );
  AND2_X1 U7265 ( .A1(n8081), .A2(n8524), .ZN(n5721) );
  NAND2_X1 U7266 ( .A1(n5715), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n5720) );
  NAND2_X1 U7267 ( .A1(n5717), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5718) );
  MUX2_X1 U7268 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5718), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n5719) );
  AND2_X1 U7269 ( .A1(n5716), .A2(n5719), .ZN(n8094) );
  XNOR2_X1 U7270 ( .A(n6512), .B(n6093), .ZN(n5722) );
  NAND2_X1 U7271 ( .A1(n5721), .A2(n5722), .ZN(n5725) );
  INV_X1 U7272 ( .A(n5721), .ZN(n5724) );
  INV_X1 U7273 ( .A(n5722), .ZN(n5723) );
  NAND2_X1 U7274 ( .A1(n5724), .A2(n5723), .ZN(n5727) );
  NAND2_X1 U7275 ( .A1(n5725), .A2(n5727), .ZN(n6420) );
  NAND2_X1 U7276 ( .A1(n6418), .A2(n5727), .ZN(n6428) );
  NAND2_X1 U7277 ( .A1(n5716), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5728) );
  XNOR2_X1 U7278 ( .A(n5728), .B(P2_IR_REG_5__SCAN_IN), .ZN(n8099) );
  INV_X1 U7279 ( .A(n8099), .ZN(n5731) );
  NAND2_X1 U7280 ( .A1(n5715), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n5729) );
  XNOR2_X1 U7281 ( .A(n6627), .B(n5732), .ZN(n5742) );
  NAND2_X1 U7282 ( .A1(n4310), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5740) );
  NAND2_X1 U7283 ( .A1(n6140), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5739) );
  NAND2_X1 U7284 ( .A1(n5733), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5752) );
  INV_X1 U7285 ( .A(n5733), .ZN(n5735) );
  INV_X1 U7286 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5734) );
  NAND2_X1 U7287 ( .A1(n5735), .A2(n5734), .ZN(n5736) );
  AND2_X1 U7288 ( .A1(n5752), .A2(n5736), .ZN(n6652) );
  NAND2_X1 U7289 ( .A1(n6145), .A2(n6652), .ZN(n5738) );
  NAND2_X1 U7290 ( .A1(n4312), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5737) );
  NAND4_X1 U7291 ( .A1(n5740), .A2(n5739), .A3(n5738), .A4(n5737), .ZN(n8080)
         );
  NAND2_X1 U7292 ( .A1(n8080), .A2(n8524), .ZN(n5741) );
  XNOR2_X1 U7293 ( .A(n5742), .B(n5741), .ZN(n6427) );
  INV_X1 U7294 ( .A(n6427), .ZN(n5745) );
  INV_X1 U7295 ( .A(n5741), .ZN(n5744) );
  INV_X1 U7296 ( .A(n5742), .ZN(n5743) );
  OR2_X1 U7297 ( .A1(n6185), .A2(n5764), .ZN(n5749) );
  OR2_X1 U7298 ( .A1(n5766), .A2(n8572), .ZN(n5747) );
  XNOR2_X1 U7299 ( .A(n5747), .B(P2_IR_REG_6__SCAN_IN), .ZN(n8111) );
  AOI22_X1 U7300 ( .A1(n7861), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n6188), .B2(
        n8111), .ZN(n5748) );
  NAND2_X1 U7301 ( .A1(n5749), .A2(n5748), .ZN(n6907) );
  XNOR2_X1 U7302 ( .A(n6907), .B(n6070), .ZN(n5758) );
  NAND2_X1 U7303 ( .A1(n4309), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5757) );
  INV_X2 U7304 ( .A(n5750), .ZN(n7868) );
  NAND2_X1 U7305 ( .A1(n7868), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5756) );
  INV_X1 U7306 ( .A(n5752), .ZN(n5751) );
  NAND2_X1 U7307 ( .A1(n5751), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5772) );
  INV_X1 U7308 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n9511) );
  NAND2_X1 U7309 ( .A1(n5752), .A2(n9511), .ZN(n5753) );
  AND2_X1 U7310 ( .A1(n5772), .A2(n5753), .ZN(n6713) );
  NAND2_X1 U7311 ( .A1(n6145), .A2(n6713), .ZN(n5755) );
  NAND2_X1 U7312 ( .A1(n4311), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5754) );
  NAND4_X1 U7313 ( .A1(n5757), .A2(n5756), .A3(n5755), .A4(n5754), .ZN(n8079)
         );
  NAND2_X1 U7314 ( .A1(n8079), .A2(n8524), .ZN(n5759) );
  NAND2_X1 U7315 ( .A1(n5758), .A2(n5759), .ZN(n5763) );
  INV_X1 U7316 ( .A(n5758), .ZN(n5761) );
  INV_X1 U7317 ( .A(n5759), .ZN(n5760) );
  NAND2_X1 U7318 ( .A1(n5761), .A2(n5760), .ZN(n5762) );
  AND2_X1 U7319 ( .A1(n5763), .A2(n5762), .ZN(n6663) );
  NAND2_X1 U7320 ( .A1(n6193), .A2(n4413), .ZN(n5769) );
  NAND2_X1 U7321 ( .A1(n5766), .A2(n5765), .ZN(n5781) );
  NAND2_X1 U7322 ( .A1(n5781), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5767) );
  XNOR2_X1 U7323 ( .A(n5767), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6369) );
  AOI22_X1 U7324 ( .A1(n7861), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6188), .B2(
        n6369), .ZN(n5768) );
  NAND2_X1 U7325 ( .A1(n5769), .A2(n5768), .ZN(n7020) );
  XNOR2_X1 U7326 ( .A(n7020), .B(n6070), .ZN(n5779) );
  NAND2_X1 U7327 ( .A1(n4309), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5777) );
  NAND2_X1 U7328 ( .A1(n4311), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5776) );
  INV_X1 U7329 ( .A(n5772), .ZN(n5770) );
  NAND2_X1 U7330 ( .A1(n5770), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5788) );
  INV_X1 U7331 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5771) );
  NAND2_X1 U7332 ( .A1(n5772), .A2(n5771), .ZN(n5773) );
  AND2_X1 U7333 ( .A1(n5788), .A2(n5773), .ZN(n6914) );
  NAND2_X1 U7334 ( .A1(n6145), .A2(n6914), .ZN(n5775) );
  NAND2_X1 U7335 ( .A1(n7868), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5774) );
  NAND4_X1 U7336 ( .A1(n5777), .A2(n5776), .A3(n5775), .A4(n5774), .ZN(n8078)
         );
  NAND2_X1 U7337 ( .A1(n8078), .A2(n10022), .ZN(n5778) );
  XNOR2_X1 U7338 ( .A(n5779), .B(n5778), .ZN(n6671) );
  NAND2_X1 U7339 ( .A1(n6203), .A2(n7981), .ZN(n5787) );
  INV_X1 U7340 ( .A(n5817), .ZN(n5785) );
  NAND2_X1 U7341 ( .A1(n5782), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5783) );
  MUX2_X1 U7342 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5783), .S(
        P2_IR_REG_8__SCAN_IN), .Z(n5784) );
  AOI22_X1 U7343 ( .A1(n7861), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6188), .B2(
        n8124), .ZN(n5786) );
  XNOR2_X1 U7344 ( .A(n7120), .B(n6093), .ZN(n5796) );
  NAND2_X1 U7345 ( .A1(n4310), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5793) );
  NAND2_X1 U7346 ( .A1(n7868), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5792) );
  NAND2_X1 U7347 ( .A1(n5788), .A2(n9590), .ZN(n5789) );
  AND2_X1 U7348 ( .A1(n5802), .A2(n5789), .ZN(n6818) );
  NAND2_X1 U7349 ( .A1(n6145), .A2(n6818), .ZN(n5791) );
  NAND2_X1 U7350 ( .A1(n4312), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5790) );
  NAND4_X1 U7351 ( .A1(n5793), .A2(n5792), .A3(n5791), .A4(n5790), .ZN(n8077)
         );
  NAND2_X1 U7352 ( .A1(n8077), .A2(n8524), .ZN(n5794) );
  XNOR2_X1 U7353 ( .A(n5796), .B(n5794), .ZN(n6817) );
  INV_X1 U7354 ( .A(n5794), .ZN(n5795) );
  NAND2_X1 U7355 ( .A1(n5796), .A2(n5795), .ZN(n5797) );
  NAND2_X1 U7356 ( .A1(n6212), .A2(n7981), .ZN(n5800) );
  OR2_X1 U7357 ( .A1(n5817), .A2(n8572), .ZN(n5798) );
  XNOR2_X1 U7358 ( .A(n5798), .B(P2_IR_REG_9__SCAN_IN), .ZN(n8136) );
  AOI22_X1 U7359 ( .A1(n7861), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6188), .B2(
        n8136), .ZN(n5799) );
  NAND2_X1 U7360 ( .A1(n5800), .A2(n5799), .ZN(n7184) );
  XNOR2_X1 U7361 ( .A(n7184), .B(n6070), .ZN(n5809) );
  NAND2_X1 U7362 ( .A1(n7868), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5808) );
  NAND2_X1 U7363 ( .A1(n4309), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5807) );
  NAND2_X1 U7364 ( .A1(n5802), .A2(n5801), .ZN(n5803) );
  NAND2_X1 U7365 ( .A1(n5821), .A2(n5803), .ZN(n7131) );
  INV_X1 U7366 ( .A(n7131), .ZN(n5804) );
  NAND2_X1 U7367 ( .A1(n6145), .A2(n5804), .ZN(n5806) );
  NAND2_X1 U7368 ( .A1(n4312), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5805) );
  NAND4_X1 U7369 ( .A1(n5808), .A2(n5807), .A3(n5806), .A4(n5805), .ZN(n8076)
         );
  NAND2_X1 U7370 ( .A1(n8076), .A2(n10022), .ZN(n5810) );
  NAND2_X1 U7371 ( .A1(n5809), .A2(n5810), .ZN(n5815) );
  INV_X1 U7372 ( .A(n5809), .ZN(n5812) );
  INV_X1 U7373 ( .A(n5810), .ZN(n5811) );
  NAND2_X1 U7374 ( .A1(n5812), .A2(n5811), .ZN(n5813) );
  NAND2_X1 U7375 ( .A1(n5815), .A2(n5813), .ZN(n6987) );
  INV_X1 U7376 ( .A(n6987), .ZN(n5814) );
  NAND2_X1 U7377 ( .A1(n6985), .A2(n5815), .ZN(n7011) );
  NAND2_X1 U7378 ( .A1(n6216), .A2(n7981), .ZN(n5819) );
  NAND2_X1 U7379 ( .A1(n5817), .A2(n5816), .ZN(n5849) );
  NAND2_X1 U7380 ( .A1(n5849), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5833) );
  XNOR2_X1 U7381 ( .A(n5833), .B(P2_IR_REG_10__SCAN_IN), .ZN(n6528) );
  AOI22_X1 U7382 ( .A1(n7861), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6188), .B2(
        n6528), .ZN(n5818) );
  NAND2_X1 U7383 ( .A1(n4309), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5826) );
  NAND2_X1 U7384 ( .A1(n7868), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5825) );
  INV_X1 U7385 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n7012) );
  NAND2_X1 U7386 ( .A1(n5821), .A2(n7012), .ZN(n5822) );
  AND2_X1 U7387 ( .A1(n5839), .A2(n5822), .ZN(n7275) );
  NAND2_X1 U7388 ( .A1(n6145), .A2(n7275), .ZN(n5824) );
  NAND2_X1 U7389 ( .A1(n4311), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5823) );
  NAND4_X1 U7390 ( .A1(n5826), .A2(n5825), .A3(n5824), .A4(n5823), .ZN(n8075)
         );
  NAND2_X1 U7391 ( .A1(n8075), .A2(n10022), .ZN(n5828) );
  XNOR2_X1 U7392 ( .A(n5827), .B(n5828), .ZN(n7010) );
  INV_X1 U7393 ( .A(n5827), .ZN(n5830) );
  INV_X1 U7394 ( .A(n5828), .ZN(n5829) );
  NAND2_X1 U7395 ( .A1(n5833), .A2(n5832), .ZN(n5834) );
  NAND2_X1 U7396 ( .A1(n5834), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5835) );
  XNOR2_X1 U7397 ( .A(n5835), .B(P2_IR_REG_11__SCAN_IN), .ZN(n6587) );
  AOI22_X1 U7398 ( .A1(n7861), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6188), .B2(
        n6587), .ZN(n5836) );
  XNOR2_X1 U7399 ( .A(n7338), .B(n6093), .ZN(n5847) );
  NAND2_X1 U7400 ( .A1(n4310), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n5844) );
  NAND2_X1 U7401 ( .A1(n7868), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5843) );
  INV_X1 U7402 ( .A(n5839), .ZN(n5837) );
  NAND2_X1 U7403 ( .A1(n5837), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5853) );
  INV_X1 U7404 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n5838) );
  NAND2_X1 U7405 ( .A1(n5839), .A2(n5838), .ZN(n5840) );
  AND2_X1 U7406 ( .A1(n5853), .A2(n5840), .ZN(n7179) );
  NAND2_X1 U7407 ( .A1(n6145), .A2(n7179), .ZN(n5842) );
  NAND2_X1 U7408 ( .A1(n4312), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5841) );
  NAND4_X1 U7409 ( .A1(n5844), .A2(n5843), .A3(n5842), .A4(n5841), .ZN(n8074)
         );
  NAND2_X1 U7410 ( .A1(n8074), .A2(n10022), .ZN(n5845) );
  XNOR2_X1 U7411 ( .A(n5847), .B(n5845), .ZN(n7163) );
  INV_X1 U7412 ( .A(n5845), .ZN(n5846) );
  AND2_X1 U7413 ( .A1(n5847), .A2(n5846), .ZN(n5848) );
  NAND2_X1 U7414 ( .A1(n6337), .A2(n7981), .ZN(n5852) );
  NAND2_X1 U7415 ( .A1(n5865), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5850) );
  XNOR2_X1 U7416 ( .A(n5850), .B(P2_IR_REG_12__SCAN_IN), .ZN(n6803) );
  AOI22_X1 U7417 ( .A1(n7861), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6188), .B2(
        n6803), .ZN(n5851) );
  XNOR2_X1 U7418 ( .A(n7416), .B(n6070), .ZN(n5859) );
  NAND2_X1 U7419 ( .A1(n4310), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5858) );
  NAND2_X1 U7420 ( .A1(n4312), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5857) );
  NAND2_X1 U7421 ( .A1(n5853), .A2(n9593), .ZN(n5854) );
  AND2_X1 U7422 ( .A1(n5870), .A2(n5854), .ZN(n7341) );
  NAND2_X1 U7423 ( .A1(n6145), .A2(n7341), .ZN(n5856) );
  NAND2_X1 U7424 ( .A1(n7868), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5855) );
  NAND4_X1 U7425 ( .A1(n5858), .A2(n5857), .A3(n5856), .A4(n5855), .ZN(n8073)
         );
  NAND2_X1 U7426 ( .A1(n8073), .A2(n10022), .ZN(n5860) );
  NAND2_X1 U7427 ( .A1(n5859), .A2(n5860), .ZN(n5864) );
  INV_X1 U7428 ( .A(n5859), .ZN(n5862) );
  INV_X1 U7429 ( .A(n5860), .ZN(n5861) );
  NAND2_X1 U7430 ( .A1(n5862), .A2(n5861), .ZN(n5863) );
  AND2_X1 U7431 ( .A1(n5864), .A2(n5863), .ZN(n7258) );
  NAND2_X1 U7432 ( .A1(n6413), .A2(n7981), .ZN(n5867) );
  OAI21_X1 U7433 ( .B1(n5865), .B2(P2_IR_REG_12__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5883) );
  XNOR2_X1 U7434 ( .A(n5883), .B(P2_IR_REG_13__SCAN_IN), .ZN(n6829) );
  AOI22_X1 U7435 ( .A1(n7861), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6188), .B2(
        n6829), .ZN(n5866) );
  XNOR2_X1 U7436 ( .A(n8550), .B(n6070), .ZN(n5877) );
  NAND2_X1 U7437 ( .A1(n4309), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5875) );
  NAND2_X1 U7438 ( .A1(n7868), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5874) );
  INV_X1 U7439 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5869) );
  NAND2_X1 U7440 ( .A1(n5870), .A2(n5869), .ZN(n5871) );
  AND2_X1 U7441 ( .A1(n5891), .A2(n5871), .ZN(n7456) );
  NAND2_X1 U7442 ( .A1(n6145), .A2(n7456), .ZN(n5873) );
  NAND2_X1 U7443 ( .A1(n4312), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n5872) );
  NAND4_X1 U7444 ( .A1(n5875), .A2(n5874), .A3(n5873), .A4(n5872), .ZN(n8072)
         );
  NAND2_X1 U7445 ( .A1(n8072), .A2(n10022), .ZN(n5878) );
  XNOR2_X1 U7446 ( .A(n5877), .B(n5878), .ZN(n7282) );
  INV_X1 U7447 ( .A(n7282), .ZN(n5876) );
  INV_X1 U7448 ( .A(n5877), .ZN(n5880) );
  INV_X1 U7449 ( .A(n5878), .ZN(n5879) );
  NAND2_X1 U7450 ( .A1(n5880), .A2(n5879), .ZN(n5881) );
  NAND2_X1 U7451 ( .A1(n6425), .A2(n7981), .ZN(n5889) );
  NAND2_X1 U7452 ( .A1(n5883), .A2(n5882), .ZN(n5884) );
  NAND2_X1 U7453 ( .A1(n5884), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5886) );
  NAND2_X1 U7454 ( .A1(n5886), .A2(n5885), .ZN(n5904) );
  OR2_X1 U7455 ( .A1(n5886), .A2(n5885), .ZN(n5887) );
  AOI22_X1 U7456 ( .A1(n7108), .A2(n6188), .B1(n5715), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n5888) );
  XNOR2_X1 U7457 ( .A(n8544), .B(n6070), .ZN(n5897) );
  NAND2_X1 U7458 ( .A1(n4309), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n5896) );
  NAND2_X1 U7459 ( .A1(n4311), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n5895) );
  INV_X1 U7460 ( .A(n5891), .ZN(n5890) );
  INV_X1 U7461 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n9537) );
  NAND2_X1 U7462 ( .A1(n5891), .A2(n9537), .ZN(n5892) );
  AND2_X1 U7463 ( .A1(n5913), .A2(n5892), .ZN(n7466) );
  NAND2_X1 U7464 ( .A1(n6145), .A2(n7466), .ZN(n5894) );
  NAND2_X1 U7465 ( .A1(n7868), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5893) );
  NAND4_X1 U7466 ( .A1(n5896), .A2(n5895), .A3(n5894), .A4(n5893), .ZN(n8071)
         );
  NAND2_X1 U7467 ( .A1(n8071), .A2(n10022), .ZN(n5898) );
  NAND2_X1 U7468 ( .A1(n5897), .A2(n5898), .ZN(n5903) );
  INV_X1 U7469 ( .A(n5897), .ZN(n5900) );
  INV_X1 U7470 ( .A(n5898), .ZN(n5899) );
  NAND2_X1 U7471 ( .A1(n5900), .A2(n5899), .ZN(n5901) );
  NAND2_X1 U7472 ( .A1(n5903), .A2(n5901), .ZN(n7465) );
  NAND2_X1 U7473 ( .A1(n7462), .A2(n5903), .ZN(n5911) );
  INV_X1 U7474 ( .A(n5911), .ZN(n5909) );
  NAND2_X1 U7475 ( .A1(n6564), .A2(n7981), .ZN(n5907) );
  NAND2_X1 U7476 ( .A1(n5904), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5905) );
  XNOR2_X1 U7477 ( .A(n5905), .B(P2_IR_REG_15__SCAN_IN), .ZN(n7216) );
  AOI22_X1 U7478 ( .A1(n7216), .A2(n6188), .B1(n5715), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n5906) );
  XNOR2_X1 U7479 ( .A(n8539), .B(n6070), .ZN(n5910) );
  INV_X1 U7480 ( .A(n5910), .ZN(n5908) );
  NAND2_X1 U7481 ( .A1(n4310), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n5918) );
  NAND2_X1 U7482 ( .A1(n4311), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n5917) );
  NAND2_X1 U7483 ( .A1(n5913), .A2(n5912), .ZN(n5914) );
  AND2_X1 U7484 ( .A1(n5925), .A2(n5914), .ZN(n7567) );
  NAND2_X1 U7485 ( .A1(n6145), .A2(n7567), .ZN(n5916) );
  NAND2_X1 U7486 ( .A1(n6140), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5915) );
  NOR2_X1 U7487 ( .A1(n7789), .A2(n7178), .ZN(n7566) );
  INV_X1 U7488 ( .A(n5919), .ZN(n7786) );
  NAND2_X1 U7489 ( .A1(n6691), .A2(n7981), .ZN(n5923) );
  OR2_X1 U7490 ( .A1(n5920), .A2(n8572), .ZN(n5921) );
  XNOR2_X1 U7491 ( .A(n5921), .B(P2_IR_REG_16__SCAN_IN), .ZN(n8153) );
  AOI22_X1 U7492 ( .A1(n7861), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n4316), .B2(
        n8153), .ZN(n5922) );
  XNOR2_X1 U7493 ( .A(n8534), .B(n6093), .ZN(n5933) );
  NAND2_X1 U7494 ( .A1(n4309), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n5930) );
  NAND2_X1 U7495 ( .A1(n6140), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5929) );
  INV_X1 U7496 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n9503) );
  NAND2_X1 U7497 ( .A1(n5925), .A2(n9503), .ZN(n5926) );
  AND2_X1 U7498 ( .A1(n5940), .A2(n5926), .ZN(n8453) );
  NAND2_X1 U7499 ( .A1(n6145), .A2(n8453), .ZN(n5928) );
  NAND2_X1 U7500 ( .A1(n4312), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n5927) );
  NAND4_X1 U7501 ( .A1(n5930), .A2(n5929), .A3(n5928), .A4(n5927), .ZN(n8415)
         );
  NAND2_X1 U7502 ( .A1(n8415), .A2(n10022), .ZN(n5931) );
  XNOR2_X1 U7503 ( .A(n5933), .B(n5931), .ZN(n7785) );
  INV_X1 U7504 ( .A(n5931), .ZN(n5932) );
  NAND2_X1 U7505 ( .A1(n6745), .A2(n7981), .ZN(n5939) );
  NAND2_X1 U7506 ( .A1(n5920), .A2(n5935), .ZN(n5936) );
  NAND2_X1 U7507 ( .A1(n5936), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5937) );
  XNOR2_X1 U7508 ( .A(n5937), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8171) );
  AOI22_X1 U7509 ( .A1(n7861), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6188), .B2(
        n8171), .ZN(n5938) );
  XNOR2_X1 U7510 ( .A(n8530), .B(n6070), .ZN(n5949) );
  NAND2_X1 U7511 ( .A1(n5940), .A2(n9500), .ZN(n5941) );
  NAND2_X1 U7512 ( .A1(n5956), .A2(n5941), .ZN(n8427) );
  INV_X1 U7513 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n5943) );
  OAI22_X1 U7514 ( .A1(n8427), .A2(n5942), .B1(n5750), .B2(n5943), .ZN(n5947)
         );
  NAND2_X1 U7515 ( .A1(n4309), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n5945) );
  NAND2_X1 U7516 ( .A1(n4312), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n5944) );
  NAND2_X1 U7517 ( .A1(n5945), .A2(n5944), .ZN(n5946) );
  NAND2_X1 U7518 ( .A1(n8439), .A2(n10022), .ZN(n5948) );
  XNOR2_X1 U7519 ( .A(n5949), .B(n5948), .ZN(n7794) );
  NAND2_X1 U7520 ( .A1(n6941), .A2(n7981), .ZN(n5953) );
  NAND2_X1 U7521 ( .A1(n5950), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5951) );
  XNOR2_X1 U7522 ( .A(n5951), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8182) );
  AOI22_X1 U7523 ( .A1(n7861), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6188), .B2(
        n8182), .ZN(n5952) );
  XNOR2_X1 U7524 ( .A(n8525), .B(n6093), .ZN(n5961) );
  INV_X1 U7525 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8172) );
  INV_X1 U7526 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n5955) );
  NAND2_X1 U7527 ( .A1(n5956), .A2(n5955), .ZN(n5957) );
  NAND2_X1 U7528 ( .A1(n5963), .A2(n5957), .ZN(n8396) );
  OR2_X1 U7529 ( .A1(n8396), .A2(n5942), .ZN(n5959) );
  AOI22_X1 U7530 ( .A1(n6140), .A2(P2_REG0_REG_18__SCAN_IN), .B1(n4309), .B2(
        P2_REG2_REG_18__SCAN_IN), .ZN(n5958) );
  OAI211_X1 U7531 ( .C1(n6088), .C2(n8172), .A(n5959), .B(n5958), .ZN(n8416)
         );
  NAND2_X1 U7532 ( .A1(n8416), .A2(n10022), .ZN(n5960) );
  XNOR2_X1 U7533 ( .A(n5961), .B(n5960), .ZN(n7823) );
  INV_X1 U7534 ( .A(n5960), .ZN(n5962) );
  INV_X1 U7535 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n5967) );
  NAND2_X1 U7536 ( .A1(n5963), .A2(n9620), .ZN(n5964) );
  NAND2_X1 U7537 ( .A1(n5974), .A2(n5964), .ZN(n7762) );
  OR2_X1 U7538 ( .A1(n7762), .A2(n5942), .ZN(n5966) );
  AOI22_X1 U7539 ( .A1(n7868), .A2(P2_REG0_REG_19__SCAN_IN), .B1(n4309), .B2(
        P2_REG2_REG_19__SCAN_IN), .ZN(n5965) );
  OAI211_X1 U7540 ( .C1(n6088), .C2(n5967), .A(n5966), .B(n5965), .ZN(n8402)
         );
  AND2_X1 U7541 ( .A1(n8402), .A2(n10022), .ZN(n5971) );
  NAND2_X1 U7542 ( .A1(n7048), .A2(n7981), .ZN(n5969) );
  AOI22_X1 U7543 ( .A1(n7861), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8283), .B2(
        n4316), .ZN(n5968) );
  XNOR2_X1 U7544 ( .A(n8521), .B(n6093), .ZN(n5970) );
  NOR2_X1 U7545 ( .A1(n5970), .A2(n5971), .ZN(n5972) );
  AOI21_X1 U7546 ( .B1(n5971), .B2(n5970), .A(n5972), .ZN(n7759) );
  INV_X1 U7547 ( .A(n5972), .ZN(n5973) );
  NAND2_X1 U7548 ( .A1(n5974), .A2(n9616), .ZN(n5975) );
  NAND2_X1 U7549 ( .A1(n5988), .A2(n5975), .ZN(n8368) );
  INV_X1 U7550 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n5978) );
  NAND2_X1 U7551 ( .A1(n4310), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n5977) );
  NAND2_X1 U7552 ( .A1(n6140), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n5976) );
  OAI211_X1 U7553 ( .C1(n6088), .C2(n5978), .A(n5977), .B(n5976), .ZN(n5979)
         );
  INV_X1 U7554 ( .A(n5979), .ZN(n5980) );
  OAI21_X1 U7555 ( .B1(n8368), .B2(n5942), .A(n5980), .ZN(n8358) );
  NAND2_X1 U7556 ( .A1(n8358), .A2(n10022), .ZN(n5984) );
  NAND2_X1 U7557 ( .A1(n7160), .A2(n7981), .ZN(n5982) );
  NAND2_X1 U7558 ( .A1(n5715), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n5981) );
  XNOR2_X1 U7559 ( .A(n8514), .B(n6093), .ZN(n5983) );
  XOR2_X1 U7560 ( .A(n5984), .B(n5983), .Z(n7808) );
  NAND2_X1 U7561 ( .A1(n7169), .A2(n7981), .ZN(n5986) );
  NAND2_X1 U7562 ( .A1(n5715), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n5985) );
  XNOR2_X1 U7563 ( .A(n8509), .B(n6093), .ZN(n5997) );
  INV_X1 U7564 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n9468) );
  NAND2_X1 U7565 ( .A1(n5988), .A2(n9468), .ZN(n5989) );
  AND2_X1 U7566 ( .A1(n6002), .A2(n5989), .ZN(n8353) );
  NAND2_X1 U7567 ( .A1(n8353), .A2(n6145), .ZN(n5995) );
  INV_X1 U7568 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n5992) );
  NAND2_X1 U7569 ( .A1(n4309), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n5991) );
  NAND2_X1 U7570 ( .A1(n6140), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n5990) );
  OAI211_X1 U7571 ( .C1(n5992), .C2(n6088), .A(n5991), .B(n5990), .ZN(n5993)
         );
  INV_X1 U7572 ( .A(n5993), .ZN(n5994) );
  NAND2_X1 U7573 ( .A1(n5995), .A2(n5994), .ZN(n8373) );
  NAND2_X1 U7574 ( .A1(n8373), .A2(n10022), .ZN(n5996) );
  XNOR2_X1 U7575 ( .A(n5997), .B(n5996), .ZN(n7769) );
  INV_X1 U7576 ( .A(n5996), .ZN(n5998) );
  NAND2_X1 U7577 ( .A1(n7350), .A2(n7981), .ZN(n6000) );
  NAND2_X1 U7578 ( .A1(n5715), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n5999) );
  XNOR2_X1 U7579 ( .A(n8504), .B(n6093), .ZN(n6011) );
  INV_X1 U7580 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n7819) );
  NAND2_X1 U7581 ( .A1(n6002), .A2(n7819), .ZN(n6003) );
  NAND2_X1 U7582 ( .A1(n6015), .A2(n6003), .ZN(n7817) );
  OR2_X1 U7583 ( .A1(n7817), .A2(n5942), .ZN(n6009) );
  INV_X1 U7584 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n6006) );
  NAND2_X1 U7585 ( .A1(n4309), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n6005) );
  NAND2_X1 U7586 ( .A1(n7868), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n6004) );
  OAI211_X1 U7587 ( .C1(n6006), .C2(n6088), .A(n6005), .B(n6004), .ZN(n6007)
         );
  INV_X1 U7588 ( .A(n6007), .ZN(n6008) );
  NAND2_X1 U7589 ( .A1(n6009), .A2(n6008), .ZN(n8359) );
  NAND2_X1 U7590 ( .A1(n8359), .A2(n10022), .ZN(n7814) );
  INV_X1 U7591 ( .A(n6010), .ZN(n6012) );
  NAND2_X2 U7592 ( .A1(n7813), .A2(n4342), .ZN(n6023) );
  NAND2_X1 U7593 ( .A1(n7411), .A2(n7981), .ZN(n6014) );
  NAND2_X1 U7594 ( .A1(n5715), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n6013) );
  XNOR2_X2 U7595 ( .A(n6023), .B(n4343), .ZN(n7751) );
  INV_X1 U7596 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n9502) );
  NAND2_X1 U7597 ( .A1(n6015), .A2(n9502), .ZN(n6016) );
  AND2_X1 U7598 ( .A1(n6027), .A2(n6016), .ZN(n8328) );
  NAND2_X1 U7599 ( .A1(n8328), .A2(n6145), .ZN(n6022) );
  INV_X1 U7600 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n6019) );
  NAND2_X1 U7601 ( .A1(n4309), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n6018) );
  NAND2_X1 U7602 ( .A1(n6140), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n6017) );
  OAI211_X1 U7603 ( .C1(n6019), .C2(n6088), .A(n6018), .B(n6017), .ZN(n6020)
         );
  INV_X1 U7604 ( .A(n6020), .ZN(n6021) );
  NAND2_X1 U7605 ( .A1(n8304), .A2(n10022), .ZN(n7752) );
  OAI22_X2 U7606 ( .A1(n7751), .A2(n7752), .B1(n4343), .B2(n6023), .ZN(n6035)
         );
  NAND2_X1 U7607 ( .A1(n7474), .A2(n7981), .ZN(n6025) );
  NAND2_X1 U7608 ( .A1(n5715), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n6024) );
  XNOR2_X1 U7609 ( .A(n8492), .B(n6093), .ZN(n6036) );
  INV_X1 U7610 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n7802) );
  NAND2_X1 U7611 ( .A1(n6027), .A2(n7802), .ZN(n6028) );
  NAND2_X1 U7612 ( .A1(n6056), .A2(n6028), .ZN(n8313) );
  OR2_X1 U7613 ( .A1(n8313), .A2(n5942), .ZN(n6034) );
  INV_X1 U7614 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n6031) );
  NAND2_X1 U7615 ( .A1(n7868), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n6030) );
  NAND2_X1 U7616 ( .A1(n4310), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n6029) );
  OAI211_X1 U7617 ( .C1(n6031), .C2(n6088), .A(n6030), .B(n6029), .ZN(n6032)
         );
  INV_X1 U7618 ( .A(n6032), .ZN(n6033) );
  NAND2_X1 U7619 ( .A1(n8217), .A2(n10022), .ZN(n7801) );
  INV_X1 U7620 ( .A(n6035), .ZN(n6038) );
  INV_X1 U7621 ( .A(n6036), .ZN(n6037) );
  OAI22_X2 U7622 ( .A1(n7800), .A2(n7801), .B1(n6038), .B2(n6037), .ZN(n7775)
         );
  NAND2_X1 U7623 ( .A1(n6039), .A2(n7981), .ZN(n6041) );
  NAND2_X1 U7624 ( .A1(n5715), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n6040) );
  XNOR2_X1 U7625 ( .A(n8488), .B(n6093), .ZN(n7777) );
  NAND2_X1 U7626 ( .A1(n7775), .A2(n7777), .ZN(n6048) );
  XNOR2_X1 U7627 ( .A(n6056), .B(P2_REG3_REG_25__SCAN_IN), .ZN(n8295) );
  NAND2_X1 U7628 ( .A1(n8295), .A2(n6145), .ZN(n6047) );
  INV_X1 U7629 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n6044) );
  NAND2_X1 U7630 ( .A1(n6140), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6043) );
  NAND2_X1 U7631 ( .A1(n4309), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n6042) );
  OAI211_X1 U7632 ( .C1(n6044), .C2(n6088), .A(n6043), .B(n6042), .ZN(n6045)
         );
  INV_X1 U7633 ( .A(n6045), .ZN(n6046) );
  NAND2_X1 U7634 ( .A1(n6047), .A2(n6046), .ZN(n8305) );
  NAND2_X1 U7635 ( .A1(n8305), .A2(n10022), .ZN(n7776) );
  INV_X1 U7636 ( .A(n7775), .ZN(n6050) );
  INV_X1 U7637 ( .A(n7777), .ZN(n6049) );
  NAND2_X1 U7638 ( .A1(n6050), .A2(n6049), .ZN(n6051) );
  NAND2_X1 U7639 ( .A1(n8587), .A2(n7981), .ZN(n6054) );
  NAND2_X1 U7640 ( .A1(n5715), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n6053) );
  XNOR2_X1 U7641 ( .A(n8483), .B(n6070), .ZN(n6065) );
  INV_X1 U7642 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n7779) );
  INV_X1 U7643 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n7837) );
  OAI21_X1 U7644 ( .B1(n6056), .B2(n7779), .A(n7837), .ZN(n6057) );
  NAND2_X1 U7645 ( .A1(P2_REG3_REG_25__SCAN_IN), .A2(P2_REG3_REG_26__SCAN_IN), 
        .ZN(n6055) );
  NAND2_X1 U7646 ( .A1(n8281), .A2(n6145), .ZN(n6063) );
  INV_X1 U7647 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n6060) );
  NAND2_X1 U7648 ( .A1(n7868), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6059) );
  NAND2_X1 U7649 ( .A1(n4310), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n6058) );
  OAI211_X1 U7650 ( .C1(n6060), .C2(n6088), .A(n6059), .B(n6058), .ZN(n6061)
         );
  INV_X1 U7651 ( .A(n6061), .ZN(n6062) );
  NAND2_X1 U7652 ( .A1(n6063), .A2(n6062), .ZN(n8223) );
  NAND2_X1 U7653 ( .A1(n8223), .A2(n10022), .ZN(n6064) );
  NOR2_X1 U7654 ( .A1(n6065), .A2(n6064), .ZN(n6066) );
  AOI21_X1 U7655 ( .B1(n6065), .B2(n6064), .A(n6066), .ZN(n7836) );
  NAND2_X1 U7656 ( .A1(n6067), .A2(n7981), .ZN(n6069) );
  NAND2_X1 U7657 ( .A1(n7861), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n6068) );
  XNOR2_X1 U7658 ( .A(n8476), .B(n6070), .ZN(n6082) );
  INV_X1 U7659 ( .A(n6073), .ZN(n6071) );
  NAND2_X1 U7660 ( .A1(n6071), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6084) );
  INV_X1 U7661 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n6072) );
  NAND2_X1 U7662 ( .A1(n6073), .A2(n6072), .ZN(n6074) );
  NAND2_X1 U7663 ( .A1(n8256), .A2(n6145), .ZN(n6080) );
  INV_X1 U7664 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n6077) );
  NAND2_X1 U7665 ( .A1(n6140), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6076) );
  NAND2_X1 U7666 ( .A1(n4310), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n6075) );
  OAI211_X1 U7667 ( .C1(n6077), .C2(n6088), .A(n6076), .B(n6075), .ZN(n6078)
         );
  INV_X1 U7668 ( .A(n6078), .ZN(n6079) );
  NAND2_X1 U7669 ( .A1(n8224), .A2(n8524), .ZN(n6081) );
  NOR2_X1 U7670 ( .A1(n6082), .A2(n6081), .ZN(n6131) );
  AOI21_X1 U7671 ( .B1(n6082), .B2(n6081), .A(n6131), .ZN(n6157) );
  INV_X1 U7672 ( .A(n6158), .ZN(n6127) );
  NAND2_X1 U7673 ( .A1(n5715), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n6083) );
  INV_X1 U7674 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n6137) );
  NAND2_X1 U7675 ( .A1(n6084), .A2(n6137), .ZN(n6085) );
  NAND2_X1 U7676 ( .A1(n8242), .A2(n6145), .ZN(n6092) );
  INV_X1 U7677 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n6089) );
  NAND2_X1 U7678 ( .A1(n6140), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6087) );
  NAND2_X1 U7679 ( .A1(n4309), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n6086) );
  OAI211_X1 U7680 ( .C1(n6089), .C2(n6088), .A(n6087), .B(n6086), .ZN(n6090)
         );
  INV_X1 U7681 ( .A(n6090), .ZN(n6091) );
  NOR2_X1 U7682 ( .A1(n8263), .A2(n7178), .ZN(n6094) );
  XNOR2_X1 U7683 ( .A(n6094), .B(n6093), .ZN(n6095) );
  XNOR2_X1 U7684 ( .A(n8471), .B(n6095), .ZN(n6130) );
  NAND2_X1 U7685 ( .A1(n6096), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6097) );
  NAND2_X1 U7686 ( .A1(n6098), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6099) );
  NAND2_X1 U7687 ( .A1(n6101), .A2(n6100), .ZN(n6102) );
  NAND2_X1 U7688 ( .A1(n6121), .A2(n6120), .ZN(n6103) );
  NAND2_X1 U7689 ( .A1(n6103), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6104) );
  XNOR2_X1 U7690 ( .A(n7475), .B(P2_B_REG_SCAN_IN), .ZN(n6105) );
  OR2_X1 U7691 ( .A1(n7504), .A2(n6105), .ZN(n6106) );
  INV_X1 U7692 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n9996) );
  NOR2_X1 U7693 ( .A1(n8589), .A2(n7504), .ZN(n9997) );
  NOR4_X1 U7694 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n6110) );
  NOR4_X1 U7695 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n6109) );
  NOR4_X1 U7696 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n6108) );
  NOR4_X1 U7697 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n6107) );
  NAND4_X1 U7698 ( .A1(n6110), .A2(n6109), .A3(n6108), .A4(n6107), .ZN(n6116)
         );
  NOR2_X1 U7699 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .ZN(
        n6114) );
  NOR4_X1 U7700 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n6113) );
  NOR4_X1 U7701 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n6112) );
  NOR4_X1 U7702 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n6111) );
  NAND4_X1 U7703 ( .A1(n6114), .A2(n6113), .A3(n6112), .A4(n6111), .ZN(n6115)
         );
  OAI21_X1 U7704 ( .B1(n6116), .B2(n6115), .A(n9991), .ZN(n6289) );
  NOR2_X1 U7705 ( .A1(n7475), .A2(n8589), .ZN(n9994) );
  INV_X1 U7706 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n9993) );
  AND2_X1 U7707 ( .A1(n6289), .A2(n6648), .ZN(n6118) );
  NAND2_X1 U7708 ( .A1(n6646), .A2(n6118), .ZN(n6132) );
  AND2_X1 U7709 ( .A1(n8589), .A2(n7504), .ZN(n6119) );
  XNOR2_X1 U7710 ( .A(n6121), .B(n6120), .ZN(n6187) );
  INV_X1 U7711 ( .A(n9998), .ZN(n9992) );
  NOR2_X1 U7712 ( .A1(n6132), .A2(n7845), .ZN(n6146) );
  NAND2_X1 U7713 ( .A1(n6124), .A2(n7874), .ZN(n6190) );
  AND2_X1 U7714 ( .A1(n10031), .A2(n6190), .ZN(n6125) );
  AND2_X1 U7715 ( .A1(n6130), .A2(n7835), .ZN(n6126) );
  NAND2_X1 U7716 ( .A1(n6127), .A2(n6126), .ZN(n6156) );
  INV_X1 U7717 ( .A(n6131), .ZN(n6129) );
  INV_X1 U7718 ( .A(n6130), .ZN(n6128) );
  NAND4_X1 U7719 ( .A1(n6158), .A2(n7835), .A3(n6129), .A4(n6128), .ZN(n6155)
         );
  NAND3_X1 U7720 ( .A1(n6131), .A2(n7835), .A3(n6130), .ZN(n6154) );
  NAND2_X1 U7721 ( .A1(n6132), .A2(n6649), .ZN(n6136) );
  INV_X1 U7722 ( .A(n7845), .ZN(n6133) );
  NAND2_X1 U7723 ( .A1(n6136), .A2(n6133), .ZN(n6491) );
  INV_X1 U7724 ( .A(n8242), .ZN(n6138) );
  OR2_X1 U7725 ( .A1(n6147), .A2(n6190), .ZN(n6286) );
  NAND2_X1 U7726 ( .A1(n6286), .A2(n6187), .ZN(n6134) );
  NOR2_X1 U7727 ( .A1(n6222), .A2(n6134), .ZN(n6135) );
  NAND2_X1 U7728 ( .A1(n6136), .A2(n6135), .ZN(n6442) );
  OAI22_X1 U7729 ( .A1(n6138), .A2(n7825), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6137), .ZN(n6152) );
  INV_X1 U7730 ( .A(n6139), .ZN(n8233) );
  NAND2_X1 U7731 ( .A1(n4311), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6143) );
  NAND2_X1 U7732 ( .A1(n6140), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6142) );
  NAND2_X1 U7733 ( .A1(n4310), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n6141) );
  NAND3_X1 U7734 ( .A1(n6143), .A2(n6142), .A3(n6141), .ZN(n6144) );
  AOI21_X1 U7735 ( .B1(n8233), .B2(n6145), .A(n6144), .ZN(n8247) );
  INV_X1 U7736 ( .A(n6146), .ZN(n6148) );
  INV_X1 U7737 ( .A(n6147), .ZN(n7844) );
  INV_X1 U7738 ( .A(n6190), .ZN(n6224) );
  INV_X1 U7739 ( .A(n6240), .ZN(n6150) );
  OAI22_X1 U7740 ( .A1(n8247), .A2(n7826), .B1(n8246), .B2(n7827), .ZN(n6151)
         );
  AOI211_X1 U7741 ( .C1(n8471), .C2(n7830), .A(n6152), .B(n6151), .ZN(n6153)
         );
  NAND3_X1 U7742 ( .A1(n6156), .A2(n6155), .A3(n4923), .ZN(P2_U3222) );
  INV_X1 U7743 ( .A(n8476), .ZN(n8258) );
  INV_X1 U7744 ( .A(n8256), .ZN(n6159) );
  NOR2_X1 U7745 ( .A1(n6159), .A2(n7825), .ZN(n6161) );
  INV_X1 U7746 ( .A(n8223), .ZN(n8262) );
  OAI22_X1 U7747 ( .A1(n8263), .A2(n7826), .B1(n8262), .B2(n7827), .ZN(n6160)
         );
  AOI211_X1 U7748 ( .C1(P2_REG3_REG_27__SCAN_IN), .C2(P2_U3152), .A(n6161), 
        .B(n6160), .ZN(n6162) );
  INV_X1 U7749 ( .A(n6163), .ZN(n6164) );
  NAND2_X1 U7750 ( .A1(n6165), .A2(n6164), .ZN(P2_U3216) );
  NAND2_X1 U7751 ( .A1(n8810), .A2(n6450), .ZN(n6167) );
  NAND2_X1 U7752 ( .A1(n6167), .A2(n6890), .ZN(n6316) );
  NAND2_X1 U7753 ( .A1(n6316), .A2(n5017), .ZN(n9778) );
  NAND2_X1 U7754 ( .A1(n9778), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  INV_X2 U7755 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  XNOR2_X1 U7756 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  INV_X1 U7757 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n7713) );
  NOR2_X1 U7758 ( .A1(n7713), .A2(P1_U3084), .ZN(n6462) );
  AOI21_X1 U7759 ( .B1(n6168), .B2(P1_U3084), .A(n6462), .ZN(n6169) );
  INV_X1 U7760 ( .A(n6169), .ZN(P1_U3353) );
  NOR2_X1 U7761 ( .A1(n6170), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8583) );
  AOI22_X1 U7762 ( .A1(n8583), .A2(P1_DATAO_REG_1__SCAN_IN), .B1(n9662), .B2(
        P2_STATE_REG_SCAN_IN), .ZN(n6171) );
  OAI21_X1 U7763 ( .B1(n7712), .B2(n6195), .A(n6171), .ZN(P2_U3357) );
  AOI22_X1 U7764 ( .A1(n8583), .A2(P1_DATAO_REG_2__SCAN_IN), .B1(n9673), .B2(
        P2_STATE_REG_SCAN_IN), .ZN(n6172) );
  OAI21_X1 U7765 ( .B1(n6174), .B2(n6195), .A(n6172), .ZN(P2_U3356) );
  NOR2_X2 U7766 ( .A1(n5462), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9428) );
  AOI22_X1 U7767 ( .A1(n9792), .A2(P1_STATE_REG_SCAN_IN), .B1(n9428), .B2(
        P2_DATAO_REG_2__SCAN_IN), .ZN(n6173) );
  OAI21_X1 U7768 ( .B1(n6174), .B2(n9420), .A(n6173), .ZN(P1_U3351) );
  AOI22_X1 U7769 ( .A1(n8583), .A2(P1_DATAO_REG_3__SCAN_IN), .B1(n6251), .B2(
        P2_STATE_REG_SCAN_IN), .ZN(n6175) );
  OAI21_X1 U7770 ( .B1(n6176), .B2(n6195), .A(n6175), .ZN(P2_U3355) );
  INV_X1 U7771 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6177) );
  INV_X1 U7772 ( .A(n6324), .ZN(n6404) );
  OAI222_X1 U7773 ( .A1(n7729), .A2(n6177), .B1(n9420), .B2(n6176), .C1(n6404), 
        .C2(P1_U3084), .ZN(P1_U3350) );
  CLKBUF_X1 U7774 ( .A(n8583), .Z(n8588) );
  AOI22_X1 U7775 ( .A1(n8094), .A2(P2_STATE_REG_SCAN_IN), .B1(n8588), .B2(
        P1_DATAO_REG_4__SCAN_IN), .ZN(n6178) );
  OAI21_X1 U7776 ( .B1(n6179), .B2(n6195), .A(n6178), .ZN(P2_U3354) );
  INV_X1 U7777 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6180) );
  INV_X1 U7778 ( .A(n6478), .ZN(n6328) );
  AOI22_X1 U7779 ( .A1(n9805), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n9428), .ZN(n6181) );
  OAI21_X1 U7780 ( .B1(n6183), .B2(n9420), .A(n6181), .ZN(P1_U3348) );
  AOI22_X1 U7781 ( .A1(n8099), .A2(P2_STATE_REG_SCAN_IN), .B1(n8588), .B2(
        P1_DATAO_REG_5__SCAN_IN), .ZN(n6182) );
  OAI21_X1 U7782 ( .B1(n6183), .B2(n6195), .A(n6182), .ZN(P2_U3353) );
  AOI22_X1 U7783 ( .A1(n8111), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_6__SCAN_IN), .B2(n8588), .ZN(n6184) );
  OAI21_X1 U7784 ( .B1(n6185), .B2(n6195), .A(n6184), .ZN(P2_U3352) );
  INV_X1 U7785 ( .A(n6351), .ZN(n6310) );
  OAI222_X1 U7786 ( .A1(n7729), .A2(n6186), .B1(n9420), .B2(n6185), .C1(n6310), 
        .C2(P1_U3084), .ZN(P1_U3347) );
  OR2_X1 U7787 ( .A1(n6187), .A2(P2_U3152), .ZN(n7846) );
  NAND2_X1 U7788 ( .A1(n7845), .A2(n7846), .ZN(n6189) );
  NAND2_X1 U7789 ( .A1(n6189), .A2(n6188), .ZN(n6192) );
  OR2_X1 U7790 ( .A1(n7845), .A2(n6190), .ZN(n6191) );
  NAND2_X1 U7791 ( .A1(n6192), .A2(n6191), .ZN(n9985) );
  NOR2_X1 U7792 ( .A1(n9985), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U7793 ( .A(n6193), .ZN(n6202) );
  AOI22_X1 U7794 ( .A1(n6369), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n8588), .ZN(n6194) );
  OAI21_X1 U7795 ( .B1(n6202), .B2(n6195), .A(n6194), .ZN(P2_U3351) );
  INV_X1 U7796 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n6200) );
  NAND2_X1 U7797 ( .A1(n4311), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n6198) );
  NAND2_X1 U7798 ( .A1(n4309), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n6197) );
  NAND2_X1 U7799 ( .A1(n7868), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n6196) );
  NAND3_X1 U7800 ( .A1(n6198), .A2(n6197), .A3(n6196), .ZN(n8055) );
  NAND2_X1 U7801 ( .A1(n8055), .A2(P2_U3966), .ZN(n6199) );
  OAI21_X1 U7802 ( .B1(n6200), .B2(P2_U3966), .A(n6199), .ZN(P2_U3583) );
  INV_X1 U7803 ( .A(n6548), .ZN(n6312) );
  OAI222_X1 U7804 ( .A1(n6312), .A2(P1_U3084), .B1(n9420), .B2(n6202), .C1(
        n6201), .C2(n7729), .ZN(P1_U3346) );
  INV_X1 U7805 ( .A(n6203), .ZN(n6205) );
  AOI22_X1 U7806 ( .A1(n8124), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_8__SCAN_IN), .B2(n8588), .ZN(n6204) );
  OAI21_X1 U7807 ( .B1(n6205), .B2(n6195), .A(n6204), .ZN(P2_U3350) );
  INV_X1 U7808 ( .A(n9821), .ZN(n9824) );
  OAI222_X1 U7809 ( .A1(n7729), .A2(n6206), .B1(n9420), .B2(n6205), .C1(n9824), 
        .C2(P1_U3084), .ZN(P1_U3345) );
  INV_X1 U7810 ( .A(n9939), .ZN(n6209) );
  OAI21_X1 U7811 ( .B1(n6209), .B2(P1_D_REG_1__SCAN_IN), .A(n6208), .ZN(n6210)
         );
  OAI21_X1 U7812 ( .B1(n6211), .B2(n9408), .A(n6210), .ZN(P1_U3441) );
  INV_X1 U7813 ( .A(n6212), .ZN(n6215) );
  AOI22_X1 U7814 ( .A1(n9831), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n9428), .ZN(n6213) );
  OAI21_X1 U7815 ( .B1(n6215), .B2(n9420), .A(n6213), .ZN(P1_U3344) );
  AOI22_X1 U7816 ( .A1(n8136), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n8588), .ZN(n6214) );
  OAI21_X1 U7817 ( .B1(n6215), .B2(n6195), .A(n6214), .ZN(P2_U3349) );
  INV_X1 U7818 ( .A(n6216), .ZN(n6220) );
  AOI22_X1 U7819 ( .A1(n6528), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_10__SCAN_IN), .B2(n8588), .ZN(n6217) );
  OAI21_X1 U7820 ( .B1(n6220), .B2(n6195), .A(n6217), .ZN(P2_U3348) );
  INV_X1 U7821 ( .A(n6218), .ZN(n6248) );
  AOI22_X1 U7822 ( .A1(n6587), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n8588), .ZN(n6219) );
  OAI21_X1 U7823 ( .B1(n6248), .B2(n6195), .A(n6219), .ZN(P2_U3347) );
  INV_X1 U7824 ( .A(n9853), .ZN(n6553) );
  OAI222_X1 U7825 ( .A1(n7729), .A2(n6221), .B1(n9420), .B2(n6220), .C1(
        P1_U3084), .C2(n6553), .ZN(P1_U3343) );
  NOR2_X1 U7826 ( .A1(n6240), .A2(P2_U3152), .ZN(n8582) );
  INV_X1 U7827 ( .A(n7846), .ZN(n8067) );
  AOI21_X1 U7828 ( .B1(n6222), .B2(n8582), .A(n8067), .ZN(n6223) );
  OAI21_X1 U7829 ( .B1(n7845), .B2(n6224), .A(n6223), .ZN(n6226) );
  NAND2_X1 U7830 ( .A1(n6226), .A2(n6225), .ZN(n6229) );
  NAND2_X1 U7831 ( .A1(n6229), .A2(n8085), .ZN(n6242) );
  NAND2_X1 U7832 ( .A1(n6242), .A2(n6240), .ZN(n9981) );
  NOR2_X1 U7833 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9605), .ZN(n6233) );
  INV_X1 U7834 ( .A(n9990), .ZN(n9988) );
  INV_X1 U7835 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n6303) );
  NAND2_X1 U7836 ( .A1(n9662), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6227) );
  OAI21_X1 U7837 ( .B1(n9662), .B2(P2_REG1_REG_1__SCAN_IN), .A(n6227), .ZN(
        n9658) );
  NOR3_X1 U7838 ( .A1(n9988), .A2(n6303), .A3(n9658), .ZN(n9657) );
  AOI21_X1 U7839 ( .B1(n9662), .B2(P2_REG1_REG_1__SCAN_IN), .A(n9657), .ZN(
        n9671) );
  NAND2_X1 U7840 ( .A1(n9673), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6228) );
  OAI21_X1 U7841 ( .B1(n9673), .B2(P2_REG1_REG_2__SCAN_IN), .A(n6228), .ZN(
        n9670) );
  NOR2_X1 U7842 ( .A1(n9671), .A2(n9670), .ZN(n9669) );
  AOI21_X1 U7843 ( .B1(n9673), .B2(P2_REG1_REG_2__SCAN_IN), .A(n9669), .ZN(
        n6231) );
  NAND2_X1 U7844 ( .A1(n6251), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6264) );
  OAI21_X1 U7845 ( .B1(n6251), .B2(P2_REG1_REG_3__SCAN_IN), .A(n6264), .ZN(
        n6230) );
  NOR2_X1 U7846 ( .A1(n6231), .A2(n6230), .ZN(n6262) );
  INV_X1 U7847 ( .A(n8202), .ZN(n8585) );
  AOI211_X1 U7848 ( .C1(n6231), .C2(n6230), .A(n6262), .B(n9983), .ZN(n6232)
         );
  AOI211_X1 U7849 ( .C1(P2_ADDR_REG_3__SCAN_IN), .C2(n9985), .A(n6233), .B(
        n6232), .ZN(n6246) );
  NAND2_X1 U7850 ( .A1(n9673), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6238) );
  INV_X1 U7851 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6234) );
  MUX2_X1 U7852 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n6234), .S(n9673), .Z(n9676)
         );
  NAND2_X1 U7853 ( .A1(n9662), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n6237) );
  INV_X1 U7854 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6235) );
  MUX2_X1 U7855 ( .A(n6235), .B(P2_REG2_REG_1__SCAN_IN), .S(n9662), .Z(n6236)
         );
  INV_X1 U7856 ( .A(n6236), .ZN(n9665) );
  NAND3_X1 U7857 ( .A1(n9990), .A2(P2_REG2_REG_0__SCAN_IN), .A3(n9665), .ZN(
        n9664) );
  NAND2_X1 U7858 ( .A1(n6237), .A2(n9664), .ZN(n9677) );
  NAND2_X1 U7859 ( .A1(n9676), .A2(n9677), .ZN(n9675) );
  NAND2_X1 U7860 ( .A1(n6238), .A2(n9675), .ZN(n6244) );
  INV_X1 U7861 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6239) );
  MUX2_X1 U7862 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n6239), .S(n6251), .Z(n6243)
         );
  NOR2_X1 U7863 ( .A1(n6240), .A2(n8202), .ZN(n6241) );
  NAND2_X1 U7864 ( .A1(n6243), .A2(n6244), .ZN(n6252) );
  OAI211_X1 U7865 ( .C1(n6244), .C2(n6243), .A(n9980), .B(n6252), .ZN(n6245)
         );
  OAI211_X1 U7866 ( .C1(n9981), .C2(n4426), .A(n6246), .B(n6245), .ZN(P2_U3248) );
  INV_X1 U7867 ( .A(n6620), .ZN(n6546) );
  INV_X1 U7868 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6247) );
  OAI222_X1 U7869 ( .A1(P1_U3084), .A2(n6546), .B1(n9420), .B2(n6248), .C1(
        n6247), .C2(n7729), .ZN(P1_U3342) );
  INV_X1 U7870 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6258) );
  INV_X1 U7871 ( .A(n8111), .ZN(n6257) );
  NAND2_X1 U7872 ( .A1(n8099), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6256) );
  INV_X1 U7873 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6249) );
  MUX2_X1 U7874 ( .A(n6249), .B(P2_REG2_REG_5__SCAN_IN), .S(n8099), .Z(n6250)
         );
  INV_X1 U7875 ( .A(n6250), .ZN(n8101) );
  INV_X1 U7876 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6255) );
  INV_X1 U7877 ( .A(n8094), .ZN(n6254) );
  NAND2_X1 U7878 ( .A1(n6251), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6253) );
  NAND2_X1 U7879 ( .A1(n6253), .A2(n6252), .ZN(n8093) );
  MUX2_X1 U7880 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n6255), .S(n8094), .Z(n8092)
         );
  NAND2_X1 U7881 ( .A1(n8093), .A2(n8092), .ZN(n8091) );
  OAI21_X1 U7882 ( .B1(n6255), .B2(n6254), .A(n8091), .ZN(n8102) );
  NAND2_X1 U7883 ( .A1(n8101), .A2(n8102), .ZN(n8100) );
  NAND2_X1 U7884 ( .A1(n6256), .A2(n8100), .ZN(n8114) );
  MUX2_X1 U7885 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n6258), .S(n8111), .Z(n8113)
         );
  NAND2_X1 U7886 ( .A1(n8114), .A2(n8113), .ZN(n8112) );
  OAI21_X1 U7887 ( .B1(n6258), .B2(n6257), .A(n8112), .ZN(n6372) );
  INV_X1 U7888 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6259) );
  MUX2_X1 U7889 ( .A(n6259), .B(P2_REG2_REG_7__SCAN_IN), .S(n6369), .Z(n6370)
         );
  XOR2_X1 U7890 ( .A(n6372), .B(n6370), .Z(n6276) );
  OR2_X1 U7891 ( .A1(n6369), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6260) );
  NAND2_X1 U7892 ( .A1(n6369), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6354) );
  AND2_X1 U7893 ( .A1(n6260), .A2(n6354), .ZN(n6270) );
  INV_X1 U7894 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6261) );
  XNOR2_X1 U7895 ( .A(n8094), .B(n6261), .ZN(n8089) );
  INV_X1 U7896 ( .A(n6262), .ZN(n6263) );
  NAND2_X1 U7897 ( .A1(n6264), .A2(n6263), .ZN(n8088) );
  NAND2_X1 U7898 ( .A1(n8089), .A2(n8088), .ZN(n8087) );
  NAND2_X1 U7899 ( .A1(n8094), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6265) );
  NAND2_X1 U7900 ( .A1(n8087), .A2(n6265), .ZN(n8105) );
  OR2_X1 U7901 ( .A1(n8099), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6266) );
  NAND2_X1 U7902 ( .A1(n8099), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6267) );
  AND2_X1 U7903 ( .A1(n6266), .A2(n6267), .ZN(n8106) );
  NAND2_X1 U7904 ( .A1(n8105), .A2(n8106), .ZN(n8104) );
  NAND2_X1 U7905 ( .A1(n8104), .A2(n6267), .ZN(n8118) );
  INV_X1 U7906 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6643) );
  MUX2_X1 U7907 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n6643), .S(n8111), .Z(n8119)
         );
  NAND2_X1 U7908 ( .A1(n8118), .A2(n8119), .ZN(n8117) );
  NAND2_X1 U7909 ( .A1(n8111), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6268) );
  NAND2_X1 U7910 ( .A1(n8117), .A2(n6268), .ZN(n6269) );
  NAND2_X1 U7911 ( .A1(n6269), .A2(n6270), .ZN(n6355) );
  OAI211_X1 U7912 ( .C1(n6270), .C2(n6269), .A(n9979), .B(n6355), .ZN(n6273)
         );
  NOR2_X1 U7913 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5771), .ZN(n6271) );
  AOI21_X1 U7914 ( .B1(n9985), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n6271), .ZN(
        n6272) );
  NAND2_X1 U7915 ( .A1(n6273), .A2(n6272), .ZN(n6274) );
  AOI21_X1 U7916 ( .B1(n6369), .B2(n9674), .A(n6274), .ZN(n6275) );
  OAI21_X1 U7917 ( .B1(n8191), .B2(n6276), .A(n6275), .ZN(P2_U3252) );
  INV_X1 U7918 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n6278) );
  NAND2_X1 U7919 ( .A1(n6454), .A2(n4315), .ZN(n6277) );
  OAI21_X1 U7920 ( .B1(n4315), .B2(n6278), .A(n6277), .ZN(P1_U3555) );
  INV_X1 U7921 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6285) );
  NAND2_X1 U7922 ( .A1(n4308), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6283) );
  NAND2_X1 U7923 ( .A1(n6279), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6282) );
  NAND2_X1 U7924 ( .A1(n6280), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6281) );
  NAND3_X1 U7925 ( .A1(n6283), .A2(n6282), .A3(n6281), .ZN(n9050) );
  NAND2_X1 U7926 ( .A1(n9050), .A2(n4315), .ZN(n6284) );
  OAI21_X1 U7927 ( .B1(n4315), .B2(n6285), .A(n6284), .ZN(P1_U3586) );
  INV_X1 U7928 ( .A(n6286), .ZN(n6287) );
  NOR2_X1 U7929 ( .A1(n7845), .A2(n6287), .ZN(n6288) );
  NAND2_X1 U7930 ( .A1(n6289), .A2(n6288), .ZN(n6645) );
  INV_X1 U7931 ( .A(n6649), .ZN(n6290) );
  NOR2_X1 U7932 ( .A1(n6645), .A2(n6290), .ZN(n6292) );
  INV_X1 U7933 ( .A(n6646), .ZN(n6291) );
  AND2_X1 U7934 ( .A1(n6292), .A2(n6291), .ZN(n6300) );
  INV_X1 U7935 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n6299) );
  INV_X1 U7936 ( .A(n6731), .ZN(n6297) );
  NAND2_X1 U7937 ( .A1(n8086), .A2(n6297), .ZN(n8005) );
  NAND2_X1 U7938 ( .A1(n6443), .A2(n8005), .ZN(n6728) );
  AND2_X1 U7939 ( .A1(n7874), .A2(n8006), .ZN(n8063) );
  INV_X1 U7940 ( .A(n8063), .ZN(n6294) );
  AND2_X1 U7941 ( .A1(n8084), .A2(n8440), .ZN(n6295) );
  AOI21_X1 U7942 ( .B1(n6728), .B2(n8411), .A(n6295), .ZN(n6729) );
  XNOR2_X1 U7943 ( .A(n7864), .B(n6644), .ZN(n8421) );
  NAND3_X1 U7944 ( .A1(n8034), .A2(n7864), .A3(n8283), .ZN(n10006) );
  NAND2_X1 U7945 ( .A1(n6728), .A2(n10034), .ZN(n6296) );
  OAI211_X1 U7946 ( .C1(n6297), .C2(n6123), .A(n6729), .B(n6296), .ZN(n6301)
         );
  NAND2_X1 U7947 ( .A1(n4314), .A2(n6301), .ZN(n6298) );
  OAI21_X1 U7948 ( .B1(n4314), .B2(n6299), .A(n6298), .ZN(P2_U3451) );
  NAND2_X1 U7949 ( .A1(n10048), .A2(n6301), .ZN(n6302) );
  OAI21_X1 U7950 ( .B1(n10048), .B2(n6303), .A(n6302), .ZN(P2_U3520) );
  INV_X1 U7951 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n6336) );
  INV_X1 U7952 ( .A(n6890), .ZN(n7413) );
  NOR2_X1 U7953 ( .A1(n6450), .A2(n7413), .ZN(n6465) );
  NOR2_X1 U7954 ( .A1(n8977), .A2(P1_U3084), .ZN(n9425) );
  NAND2_X1 U7955 ( .A1(n6316), .A2(n9425), .ZN(n9044) );
  INV_X1 U7956 ( .A(n9044), .ZN(n6304) );
  AND2_X1 U7957 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7073) );
  INV_X1 U7958 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6311) );
  NAND2_X1 U7959 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(n9805), .ZN(n6309) );
  INV_X1 U7960 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6305) );
  MUX2_X1 U7961 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n6305), .S(n9805), .Z(n9811)
         );
  INV_X1 U7962 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6308) );
  MUX2_X1 U7963 ( .A(n6308), .B(P1_REG1_REG_4__SCAN_IN), .S(n6478), .Z(n6469)
         );
  INV_X1 U7964 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6307) );
  INV_X1 U7965 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n9971) );
  MUX2_X1 U7966 ( .A(n9971), .B(P1_REG1_REG_1__SCAN_IN), .S(n7726), .Z(n7714)
         );
  INV_X1 U7967 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9969) );
  NOR3_X1 U7968 ( .A1(n7714), .A2(n9969), .A3(n7713), .ZN(n7715) );
  AOI21_X1 U7969 ( .B1(P1_REG1_REG_1__SCAN_IN), .B2(n7726), .A(n7715), .ZN(
        n9800) );
  INV_X1 U7970 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6306) );
  MUX2_X1 U7971 ( .A(n6306), .B(P1_REG1_REG_2__SCAN_IN), .S(n9792), .Z(n9799)
         );
  AND2_X1 U7972 ( .A1(n9792), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6398) );
  MUX2_X1 U7973 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n6307), .S(n6324), .Z(n6399)
         );
  OAI21_X1 U7974 ( .B1(n9798), .B2(n6398), .A(n6399), .ZN(n6401) );
  OAI21_X1 U7975 ( .B1(n6307), .B2(n6404), .A(n6401), .ZN(n6470) );
  NOR2_X1 U7976 ( .A1(n6469), .A2(n6470), .ZN(n6468) );
  NAND2_X1 U7977 ( .A1(n9811), .A2(n9812), .ZN(n9810) );
  NAND2_X1 U7978 ( .A1(n6309), .A2(n9810), .ZN(n6343) );
  MUX2_X1 U7979 ( .A(n6311), .B(P1_REG1_REG_6__SCAN_IN), .S(n6351), .Z(n6342)
         );
  NOR2_X1 U7980 ( .A1(n6343), .A2(n6342), .ZN(n6341) );
  INV_X1 U7981 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n9973) );
  AOI22_X1 U7982 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(n6312), .B1(n6548), .B2(
        n9973), .ZN(n6313) );
  NOR2_X1 U7983 ( .A1(n6314), .A2(n6313), .ZN(n6549) );
  AOI21_X1 U7984 ( .B1(n6314), .B2(n6313), .A(n6549), .ZN(n6317) );
  OR2_X1 U7985 ( .A1(n4317), .A2(P1_U3084), .ZN(n9422) );
  INV_X1 U7986 ( .A(n8977), .ZN(n6461) );
  NOR2_X1 U7987 ( .A1(n9422), .A2(n6461), .ZN(n6315) );
  NAND2_X1 U7988 ( .A1(n6316), .A2(n6315), .ZN(n9797) );
  NOR2_X1 U7989 ( .A1(n6317), .A2(n9797), .ZN(n6318) );
  AOI211_X1 U7990 ( .C1(n9860), .C2(n6548), .A(n7073), .B(n6318), .ZN(n6335)
         );
  INV_X1 U7991 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6327) );
  INV_X1 U7992 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6326) );
  INV_X1 U7993 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6319) );
  MUX2_X1 U7994 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n6319), .S(n9792), .Z(n6323)
         );
  INV_X1 U7995 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6320) );
  AND2_X1 U7996 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n6321) );
  NAND2_X1 U7997 ( .A1(n7721), .A2(n6321), .ZN(n7720) );
  NAND2_X1 U7998 ( .A1(n7726), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6322) );
  NAND2_X1 U7999 ( .A1(n7720), .A2(n6322), .ZN(n9787) );
  NAND2_X1 U8000 ( .A1(n6323), .A2(n9787), .ZN(n9791) );
  NAND2_X1 U8001 ( .A1(n9792), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6406) );
  MUX2_X1 U8002 ( .A(n6326), .B(P1_REG2_REG_3__SCAN_IN), .S(n6324), .Z(n6407)
         );
  AOI21_X1 U8003 ( .B1(n9791), .B2(n6406), .A(n6407), .ZN(n6325) );
  INV_X1 U8004 ( .A(n6325), .ZN(n6409) );
  OAI21_X1 U8005 ( .B1(n6326), .B2(n6404), .A(n6409), .ZN(n6474) );
  MUX2_X1 U8006 ( .A(n6327), .B(P1_REG2_REG_4__SCAN_IN), .S(n6478), .Z(n6473)
         );
  MUX2_X1 U8007 ( .A(n6329), .B(P1_REG2_REG_5__SCAN_IN), .S(n9805), .Z(n9808)
         );
  INV_X1 U8008 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n9274) );
  MUX2_X1 U8009 ( .A(n9274), .B(P1_REG2_REG_6__SCAN_IN), .S(n6351), .Z(n6348)
         );
  INV_X1 U8010 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n6330) );
  MUX2_X1 U8011 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n6330), .S(n6548), .Z(n6331)
         );
  NOR2_X1 U8012 ( .A1(n6332), .A2(n6331), .ZN(n6333) );
  OR2_X1 U8013 ( .A1(n9044), .A2(n4317), .ZN(n9847) );
  INV_X1 U8014 ( .A(n9847), .ZN(n9869) );
  OAI21_X1 U8015 ( .B1(n6538), .B2(n6333), .A(n9869), .ZN(n6334) );
  OAI211_X1 U8016 ( .C1(n6336), .C2(n9873), .A(n6335), .B(n6334), .ZN(P1_U3248) );
  INV_X1 U8017 ( .A(n6337), .ZN(n6340) );
  AOI22_X1 U8018 ( .A1(n6776), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n9428), .ZN(n6338) );
  OAI21_X1 U8019 ( .B1(n6340), .B2(n9420), .A(n6338), .ZN(P1_U3341) );
  AOI22_X1 U8020 ( .A1(n6803), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_12__SCAN_IN), .B2(n8588), .ZN(n6339) );
  OAI21_X1 U8021 ( .B1(n6340), .B2(n6195), .A(n6339), .ZN(P2_U3346) );
  INV_X1 U8022 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n6353) );
  AOI21_X1 U8023 ( .B1(n6343), .B2(n6342), .A(n6341), .ZN(n6346) );
  NOR2_X1 U8024 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6344), .ZN(n7004) );
  INV_X1 U8025 ( .A(n7004), .ZN(n6345) );
  OAI21_X1 U8026 ( .B1(n6346), .B2(n9797), .A(n6345), .ZN(n6350) );
  AOI211_X1 U8027 ( .C1(n4318), .C2(n6348), .A(n6347), .B(n9847), .ZN(n6349)
         );
  AOI211_X1 U8028 ( .C1(n9860), .C2(n6351), .A(n6350), .B(n6349), .ZN(n6352)
         );
  OAI21_X1 U8029 ( .B1(n9873), .B2(n6353), .A(n6352), .ZN(P1_U3247) );
  NAND2_X1 U8030 ( .A1(n6355), .A2(n6354), .ZN(n8130) );
  INV_X1 U8031 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n7044) );
  MUX2_X1 U8032 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n7044), .S(n8124), .Z(n8131)
         );
  NAND2_X1 U8033 ( .A1(n8130), .A2(n8131), .ZN(n8129) );
  NAND2_X1 U8034 ( .A1(n8124), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n6356) );
  NAND2_X1 U8035 ( .A1(n8129), .A2(n6356), .ZN(n8143) );
  INV_X1 U8036 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10044) );
  MUX2_X1 U8037 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n10044), .S(n8136), .Z(n8144)
         );
  NAND2_X1 U8038 ( .A1(n8143), .A2(n8144), .ZN(n8142) );
  NAND2_X1 U8039 ( .A1(n8136), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n6357) );
  AND2_X1 U8040 ( .A1(n8142), .A2(n6357), .ZN(n6360) );
  INV_X1 U8041 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n6358) );
  MUX2_X1 U8042 ( .A(n6358), .B(P2_REG1_REG_10__SCAN_IN), .S(n6528), .Z(n6359)
         );
  NAND2_X1 U8043 ( .A1(n6360), .A2(n6359), .ZN(n6362) );
  NOR2_X1 U8044 ( .A1(n6360), .A2(n6359), .ZN(n6520) );
  INV_X1 U8045 ( .A(n6520), .ZN(n6361) );
  NAND2_X1 U8046 ( .A1(n6362), .A2(n6361), .ZN(n6365) );
  NOR2_X1 U8047 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7012), .ZN(n6363) );
  AOI21_X1 U8048 ( .B1(n9985), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n6363), .ZN(
        n6364) );
  OAI21_X1 U8049 ( .B1(n9983), .B2(n6365), .A(n6364), .ZN(n6366) );
  AOI21_X1 U8050 ( .B1(n6528), .B2(n9674), .A(n6366), .ZN(n6382) );
  NAND2_X1 U8051 ( .A1(n8136), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6376) );
  INV_X1 U8052 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n6367) );
  MUX2_X1 U8053 ( .A(n6367), .B(P2_REG2_REG_9__SCAN_IN), .S(n8136), .Z(n6368)
         );
  INV_X1 U8054 ( .A(n6368), .ZN(n8138) );
  INV_X1 U8055 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7032) );
  INV_X1 U8056 ( .A(n8124), .ZN(n6375) );
  NAND2_X1 U8057 ( .A1(n6369), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6374) );
  INV_X1 U8058 ( .A(n6370), .ZN(n6371) );
  NAND2_X1 U8059 ( .A1(n6372), .A2(n6371), .ZN(n6373) );
  NAND2_X1 U8060 ( .A1(n6374), .A2(n6373), .ZN(n8127) );
  MUX2_X1 U8061 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n7032), .S(n8124), .Z(n8126)
         );
  NAND2_X1 U8062 ( .A1(n8127), .A2(n8126), .ZN(n8125) );
  OAI21_X1 U8063 ( .B1(n7032), .B2(n6375), .A(n8125), .ZN(n8139) );
  NAND2_X1 U8064 ( .A1(n8138), .A2(n8139), .ZN(n8137) );
  NAND2_X1 U8065 ( .A1(n6376), .A2(n8137), .ZN(n6380) );
  INV_X1 U8066 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n6377) );
  MUX2_X1 U8067 ( .A(n6377), .B(P2_REG2_REG_10__SCAN_IN), .S(n6528), .Z(n6378)
         );
  INV_X1 U8068 ( .A(n6378), .ZN(n6379) );
  NAND2_X1 U8069 ( .A1(n6379), .A2(n6380), .ZN(n6529) );
  OAI211_X1 U8070 ( .C1(n6380), .C2(n6379), .A(n9980), .B(n6529), .ZN(n6381)
         );
  NAND2_X1 U8071 ( .A1(n6382), .A2(n6381), .ZN(P2_U3255) );
  INV_X1 U8072 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n6394) );
  INV_X1 U8073 ( .A(n8084), .ZN(n6383) );
  NAND2_X1 U8074 ( .A1(n6383), .A2(n6701), .ZN(n7886) );
  NAND2_X1 U8075 ( .A1(n7886), .A2(n7883), .ZN(n6695) );
  NAND2_X1 U8076 ( .A1(n8086), .A2(n6731), .ZN(n6697) );
  NAND2_X1 U8077 ( .A1(n6695), .A2(n6697), .ZN(n6696) );
  NAND2_X1 U8078 ( .A1(n6383), .A2(n6492), .ZN(n6384) );
  NAND2_X1 U8079 ( .A1(n6696), .A2(n6384), .ZN(n6385) );
  NAND2_X1 U8080 ( .A1(n6385), .A2(n6387), .ZN(n6502) );
  OAI21_X1 U8081 ( .B1(n6385), .B2(n6387), .A(n6502), .ZN(n6725) );
  NAND2_X1 U8082 ( .A1(n6698), .A2(n6500), .ZN(n6760) );
  OR2_X1 U8083 ( .A1(n6698), .A2(n6500), .ZN(n6386) );
  NAND2_X1 U8084 ( .A1(n6760), .A2(n6386), .ZN(n6720) );
  OAI22_X1 U8085 ( .A1(n6720), .A2(n10022), .B1(n6500), .B2(n10031), .ZN(n6392) );
  INV_X1 U8086 ( .A(n6387), .ZN(n8008) );
  NAND2_X1 U8087 ( .A1(n6443), .A2(n7886), .ZN(n7875) );
  NAND2_X1 U8088 ( .A1(n6388), .A2(n8008), .ZN(n6506) );
  OAI21_X1 U8089 ( .B1(n8008), .B2(n6388), .A(n6506), .ZN(n6389) );
  NAND2_X1 U8090 ( .A1(n6389), .A2(n8411), .ZN(n6391) );
  AOI22_X1 U8091 ( .A1(n8441), .A2(n8084), .B1(n8082), .B2(n8440), .ZN(n6390)
         );
  NAND2_X1 U8092 ( .A1(n6391), .A2(n6390), .ZN(n6723) );
  AOI211_X1 U8093 ( .C1(n10034), .C2(n6725), .A(n6392), .B(n6723), .ZN(n6395)
         );
  OR2_X1 U8094 ( .A1(n6395), .A2(n10036), .ZN(n6393) );
  OAI21_X1 U8095 ( .B1(n4314), .B2(n6394), .A(n6393), .ZN(P2_U3457) );
  INV_X1 U8096 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6397) );
  OR2_X1 U8097 ( .A1(n6395), .A2(n10046), .ZN(n6396) );
  OAI21_X1 U8098 ( .B1(n10048), .B2(n6397), .A(n6396), .ZN(P2_U3522) );
  INV_X1 U8099 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n6412) );
  INV_X1 U8100 ( .A(n9860), .ZN(n9023) );
  NOR2_X1 U8101 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n4986), .ZN(n6900) );
  INV_X1 U8102 ( .A(n6900), .ZN(n6403) );
  OR3_X1 U8103 ( .A1(n6399), .A2(n9798), .A3(n6398), .ZN(n6400) );
  NAND3_X1 U8104 ( .A1(n9868), .A2(n6401), .A3(n6400), .ZN(n6402) );
  OAI211_X1 U8105 ( .C1(n9023), .C2(n6404), .A(n6403), .B(n6402), .ZN(n6405)
         );
  INV_X1 U8106 ( .A(n6405), .ZN(n6411) );
  NAND3_X1 U8107 ( .A1(n6407), .A2(n9791), .A3(n6406), .ZN(n6408) );
  NAND3_X1 U8108 ( .A1(n9869), .A2(n6409), .A3(n6408), .ZN(n6410) );
  OAI211_X1 U8109 ( .C1(n6412), .C2(n9873), .A(n6411), .B(n6410), .ZN(P1_U3244) );
  INV_X1 U8110 ( .A(n6413), .ZN(n6416) );
  AOI22_X1 U8111 ( .A1(n7058), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n9428), .ZN(n6414) );
  OAI21_X1 U8112 ( .B1(n6416), .B2(n9420), .A(n6414), .ZN(P1_U3340) );
  AOI22_X1 U8113 ( .A1(n6829), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(n8588), .ZN(n6415) );
  OAI21_X1 U8114 ( .B1(n6416), .B2(n6195), .A(n6415), .ZN(P2_U3345) );
  INV_X1 U8115 ( .A(n6418), .ZN(n6419) );
  AOI21_X1 U8116 ( .B1(n6417), .B2(n6420), .A(n6419), .ZN(n6424) );
  INV_X1 U8117 ( .A(n8082), .ZN(n6503) );
  INV_X1 U8118 ( .A(n8080), .ZN(n6666) );
  OAI22_X1 U8119 ( .A1(n6503), .A2(n8326), .B1(n6666), .B2(n8324), .ZN(n6508)
         );
  NOR2_X1 U8120 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9629), .ZN(n8090) );
  AOI21_X1 U8121 ( .B1(n7763), .B2(n6508), .A(n8090), .ZN(n6421) );
  OAI21_X1 U8122 ( .B1(n6686), .B2(n7843), .A(n6421), .ZN(n6422) );
  AOI21_X1 U8123 ( .B1(n6682), .B2(n7840), .A(n6422), .ZN(n6423) );
  OAI21_X1 U8124 ( .B1(n6424), .B2(n4570), .A(n6423), .ZN(P2_U3232) );
  INV_X1 U8125 ( .A(n6425), .ZN(n6499) );
  AOI22_X1 U8126 ( .A1(n7108), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_14__SCAN_IN), .B2(n8588), .ZN(n6426) );
  OAI21_X1 U8127 ( .B1(n6499), .B2(n6195), .A(n6426), .ZN(P2_U3344) );
  XNOR2_X1 U8128 ( .A(n6428), .B(n6427), .ZN(n6435) );
  INV_X1 U8129 ( .A(n6652), .ZN(n6432) );
  NAND2_X1 U8130 ( .A1(n8079), .A2(n8440), .ZN(n6430) );
  NAND2_X1 U8131 ( .A1(n8081), .A2(n8441), .ZN(n6429) );
  NAND2_X1 U8132 ( .A1(n6430), .A2(n6429), .ZN(n6570) );
  AOI22_X1 U8133 ( .A1(n7763), .A2(n6570), .B1(P2_REG3_REG_5__SCAN_IN), .B2(
        P2_U3152), .ZN(n6431) );
  OAI21_X1 U8134 ( .B1(n6432), .B2(n7825), .A(n6431), .ZN(n6433) );
  AOI21_X1 U8135 ( .B1(n7830), .B2(n6627), .A(n6433), .ZN(n6434) );
  OAI21_X1 U8136 ( .B1(n6435), .B2(n4570), .A(n6434), .ZN(P2_U3229) );
  XNOR2_X1 U8137 ( .A(n6436), .B(n6437), .ZN(n6441) );
  INV_X1 U8138 ( .A(n7827), .ZN(n6675) );
  INV_X1 U8139 ( .A(n8081), .ZN(n6754) );
  OAI22_X1 U8140 ( .A1(n7826), .A2(n6754), .B1(n10008), .B2(n7843), .ZN(n6438)
         );
  AOI21_X1 U8141 ( .B1(n6675), .B2(n8083), .A(n6438), .ZN(n6440) );
  MUX2_X1 U8142 ( .A(n7825), .B(P2_STATE_REG_SCAN_IN), .S(
        P2_REG3_REG_3__SCAN_IN), .Z(n6439) );
  OAI211_X1 U8143 ( .C1(n4570), .C2(n6441), .A(n6440), .B(n6439), .ZN(P2_U3220) );
  OR2_X1 U8144 ( .A1(n6442), .A2(P2_U3152), .ZN(n6484) );
  INV_X1 U8145 ( .A(n6484), .ZN(n6497) );
  INV_X1 U8146 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n9524) );
  INV_X1 U8147 ( .A(n7826), .ZN(n6673) );
  AOI22_X1 U8148 ( .A1(n6673), .A2(n8084), .B1(n7830), .B2(n6731), .ZN(n6447)
         );
  INV_X1 U8149 ( .A(n6443), .ZN(n6702) );
  INV_X1 U8150 ( .A(n8005), .ZN(n6444) );
  MUX2_X1 U8151 ( .A(n6731), .B(n6444), .S(n8524), .Z(n6445) );
  OAI21_X1 U8152 ( .B1(n6702), .B2(n6445), .A(n7835), .ZN(n6446) );
  OAI211_X1 U8153 ( .C1(n6497), .C2(n9524), .A(n6447), .B(n6446), .ZN(P2_U3234) );
  INV_X1 U8154 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n6481) );
  INV_X1 U8155 ( .A(n6450), .ZN(n6451) );
  AOI22_X1 U8156 ( .A1(n9930), .A2(n7146), .B1(n6451), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n6452) );
  AND2_X1 U8157 ( .A1(n6453), .A2(n6452), .ZN(n6458) );
  NAND2_X1 U8158 ( .A1(n6454), .A2(n7146), .ZN(n6457) );
  NOR2_X1 U8159 ( .A1(n6450), .A2(n9969), .ZN(n6455) );
  AOI21_X1 U8160 ( .B1(n9930), .B2(n6865), .A(n6455), .ZN(n6456) );
  NAND2_X1 U8161 ( .A1(n6458), .A2(n6859), .ZN(n6861) );
  OAI21_X1 U8162 ( .B1(n6458), .B2(n6859), .A(n6861), .ZN(n6791) );
  NAND2_X1 U8163 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n7719) );
  NAND2_X1 U8164 ( .A1(n6461), .A2(n7719), .ZN(n6459) );
  NAND2_X1 U8165 ( .A1(n6898), .A2(n6459), .ZN(n9777) );
  AOI21_X1 U8166 ( .B1(n6791), .B2(n8977), .A(n9777), .ZN(n6467) );
  INV_X1 U8167 ( .A(n9422), .ZN(n6464) );
  INV_X1 U8168 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n6460) );
  NAND2_X1 U8169 ( .A1(n6461), .A2(n6460), .ZN(n6463) );
  AOI21_X1 U8170 ( .B1(n6464), .B2(n6463), .A(n6462), .ZN(n9780) );
  INV_X1 U8171 ( .A(n6465), .ZN(n6466) );
  NOR3_X1 U8172 ( .A1(n6467), .A2(n9780), .A3(n6466), .ZN(n9795) );
  INV_X1 U8173 ( .A(n9795), .ZN(n6480) );
  AOI21_X1 U8174 ( .B1(n6470), .B2(n6469), .A(n6468), .ZN(n6471) );
  NAND2_X1 U8175 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n6933) );
  OAI21_X1 U8176 ( .B1(n9797), .B2(n6471), .A(n6933), .ZN(n6477) );
  AOI21_X1 U8177 ( .B1(n6474), .B2(n6473), .A(n6472), .ZN(n6475) );
  NOR2_X1 U8178 ( .A1(n9847), .A2(n6475), .ZN(n6476) );
  AOI211_X1 U8179 ( .C1(n9860), .C2(n6478), .A(n6477), .B(n6476), .ZN(n6479)
         );
  OAI211_X1 U8180 ( .C1(n9873), .C2(n6481), .A(n6480), .B(n6479), .ZN(P1_U3245) );
  XNOR2_X1 U8181 ( .A(n6482), .B(n6483), .ZN(n6487) );
  AOI22_X1 U8182 ( .A1(n6675), .A2(n8084), .B1(n6673), .B2(n8082), .ZN(n6486)
         );
  AOI22_X1 U8183 ( .A1(n7830), .A2(n6724), .B1(P2_REG3_REG_2__SCAN_IN), .B2(
        n6484), .ZN(n6485) );
  OAI211_X1 U8184 ( .C1(n6487), .C2(n4570), .A(n6486), .B(n6485), .ZN(P2_U3239) );
  INV_X1 U8185 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n9654) );
  AOI22_X1 U8186 ( .A1(n6675), .A2(n8086), .B1(n6673), .B2(n8083), .ZN(n6496)
         );
  OAI21_X1 U8187 ( .B1(n6488), .B2(n6490), .A(n6489), .ZN(n6494) );
  INV_X1 U8188 ( .A(n6491), .ZN(n6493) );
  NOR2_X1 U8189 ( .A1(n6492), .A2(n10031), .ZN(n9999) );
  AOI22_X1 U8190 ( .A1(n7835), .A2(n6494), .B1(n6493), .B2(n9999), .ZN(n6495)
         );
  OAI211_X1 U8191 ( .C1(n6497), .C2(n9654), .A(n6496), .B(n6495), .ZN(P2_U3224) );
  INV_X1 U8192 ( .A(n7295), .ZN(n7288) );
  INV_X1 U8193 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6498) );
  OAI222_X1 U8194 ( .A1(P1_U3084), .A2(n7288), .B1(n9420), .B2(n6499), .C1(
        n6498), .C2(n7729), .ZN(P1_U3339) );
  INV_X1 U8195 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n6516) );
  NAND2_X1 U8196 ( .A1(n4846), .A2(n6500), .ZN(n6501) );
  NAND2_X1 U8197 ( .A1(n6502), .A2(n6501), .ZN(n6750) );
  NAND2_X1 U8198 ( .A1(n8082), .A2(n10008), .ZN(n7889) );
  NAND2_X1 U8199 ( .A1(n6750), .A2(n8011), .ZN(n6749) );
  NAND2_X1 U8200 ( .A1(n6503), .A2(n10008), .ZN(n6504) );
  NAND2_X1 U8201 ( .A1(n6749), .A2(n6504), .ZN(n6505) );
  OR2_X1 U8202 ( .A1(n8081), .A2(n6686), .ZN(n7869) );
  NAND2_X1 U8203 ( .A1(n7869), .A2(n6630), .ZN(n8009) );
  OAI21_X1 U8204 ( .B1(n6505), .B2(n8009), .A(n6567), .ZN(n6688) );
  INV_X1 U8205 ( .A(n6688), .ZN(n6514) );
  NAND2_X1 U8206 ( .A1(n6506), .A2(n7884), .ZN(n6753) );
  INV_X1 U8207 ( .A(n8011), .ZN(n7879) );
  NAND2_X1 U8208 ( .A1(n6752), .A2(n6568), .ZN(n6507) );
  XOR2_X1 U8209 ( .A(n8009), .B(n6507), .Z(n6509) );
  AOI21_X1 U8210 ( .B1(n6509), .B2(n8411), .A(n6508), .ZN(n6690) );
  NAND2_X1 U8211 ( .A1(n6758), .A2(n6512), .ZN(n6510) );
  NAND2_X1 U8212 ( .A1(n6510), .A2(n7178), .ZN(n6511) );
  NOR2_X1 U8213 ( .A1(n6572), .A2(n6511), .ZN(n6683) );
  AOI21_X1 U8214 ( .B1(n9693), .B2(n6512), .A(n6683), .ZN(n6513) );
  OAI211_X1 U8215 ( .C1(n6514), .C2(n8549), .A(n6690), .B(n6513), .ZN(n6517)
         );
  NAND2_X1 U8216 ( .A1(n6517), .A2(n4314), .ZN(n6515) );
  OAI21_X1 U8217 ( .B1(n4314), .B2(n6516), .A(n6515), .ZN(P2_U3463) );
  NAND2_X1 U8218 ( .A1(n6517), .A2(n10048), .ZN(n6518) );
  OAI21_X1 U8219 ( .B1(n10048), .B2(n6261), .A(n6518), .ZN(P2_U3524) );
  INV_X1 U8220 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n6519) );
  MUX2_X1 U8221 ( .A(n6519), .B(P2_REG1_REG_11__SCAN_IN), .S(n6587), .Z(n6521)
         );
  AOI21_X1 U8222 ( .B1(n6528), .B2(P2_REG1_REG_10__SCAN_IN), .A(n6520), .ZN(
        n6522) );
  NAND2_X1 U8223 ( .A1(n6521), .A2(n6522), .ZN(n6524) );
  NOR2_X1 U8224 ( .A1(n6522), .A2(n6521), .ZN(n6580) );
  INV_X1 U8225 ( .A(n6580), .ZN(n6523) );
  NAND2_X1 U8226 ( .A1(n6524), .A2(n6523), .ZN(n6527) );
  NOR2_X1 U8227 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5838), .ZN(n6525) );
  AOI21_X1 U8228 ( .B1(n9985), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n6525), .ZN(
        n6526) );
  OAI21_X1 U8229 ( .B1(n9983), .B2(n6527), .A(n6526), .ZN(n6536) );
  NAND2_X1 U8230 ( .A1(n6528), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6530) );
  NAND2_X1 U8231 ( .A1(n6530), .A2(n6529), .ZN(n6533) );
  INV_X1 U8232 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n6531) );
  MUX2_X1 U8233 ( .A(n6531), .B(P2_REG2_REG_11__SCAN_IN), .S(n6587), .Z(n6532)
         );
  NOR2_X1 U8234 ( .A1(n6533), .A2(n6532), .ZN(n6588) );
  AOI21_X1 U8235 ( .B1(n6533), .B2(n6532), .A(n6588), .ZN(n6534) );
  NOR2_X1 U8236 ( .A1(n6534), .A2(n8191), .ZN(n6535) );
  AOI211_X1 U8237 ( .C1(n9674), .C2(n6587), .A(n6536), .B(n6535), .ZN(n6537)
         );
  INV_X1 U8238 ( .A(n6537), .ZN(P2_U3256) );
  NOR2_X1 U8239 ( .A1(P1_REG2_REG_7__SCAN_IN), .A2(n6548), .ZN(n6539) );
  INV_X1 U8240 ( .A(n9818), .ZN(n6540) );
  NOR2_X1 U8241 ( .A1(n6540), .A2(n5072), .ZN(n6541) );
  OAI22_X1 U8242 ( .A1(n6541), .A2(n9821), .B1(P1_REG2_REG_8__SCAN_IN), .B2(
        n9818), .ZN(n9836) );
  NAND2_X1 U8243 ( .A1(n9831), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6542) );
  OAI21_X1 U8244 ( .B1(n9831), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6542), .ZN(
        n9837) );
  NOR2_X1 U8245 ( .A1(n9836), .A2(n9837), .ZN(n9835) );
  AOI21_X1 U8246 ( .B1(P1_REG2_REG_9__SCAN_IN), .B2(n9831), .A(n9835), .ZN(
        n9849) );
  XNOR2_X1 U8247 ( .A(n9853), .B(P1_REG2_REG_10__SCAN_IN), .ZN(n9848) );
  NOR2_X1 U8248 ( .A1(n9849), .A2(n9848), .ZN(n9846) );
  AOI21_X1 U8249 ( .B1(n9853), .B2(P1_REG2_REG_10__SCAN_IN), .A(n9846), .ZN(
        n6545) );
  INV_X1 U8250 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n6543) );
  AOI22_X1 U8251 ( .A1(P1_REG2_REG_11__SCAN_IN), .A2(n6620), .B1(n6546), .B2(
        n6543), .ZN(n6544) );
  NAND2_X1 U8252 ( .A1(n6544), .A2(n6545), .ZN(n6619) );
  OAI21_X1 U8253 ( .B1(n6545), .B2(n6544), .A(n6619), .ZN(n6562) );
  INV_X1 U8254 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n6560) );
  INV_X1 U8255 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n9767) );
  AOI22_X1 U8256 ( .A1(P1_REG1_REG_11__SCAN_IN), .A2(n6620), .B1(n6546), .B2(
        n9767), .ZN(n6556) );
  INV_X1 U8257 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6552) );
  MUX2_X1 U8258 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n6552), .S(n9853), .Z(n9844)
         );
  NOR2_X1 U8259 ( .A1(n9831), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6547) );
  AOI21_X1 U8260 ( .B1(P1_REG1_REG_9__SCAN_IN), .B2(n9831), .A(n6547), .ZN(
        n9833) );
  NOR2_X1 U8261 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(n6548), .ZN(n6550) );
  NOR2_X1 U8262 ( .A1(n6550), .A2(n6549), .ZN(n9826) );
  INV_X1 U8263 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9823) );
  OAI22_X1 U8264 ( .A1(n6551), .A2(n9821), .B1(P1_REG1_REG_8__SCAN_IN), .B2(
        n9826), .ZN(n9834) );
  NAND2_X1 U8265 ( .A1(n9833), .A2(n9834), .ZN(n9832) );
  NAND2_X1 U8266 ( .A1(n6553), .A2(n6552), .ZN(n6554) );
  NAND2_X1 U8267 ( .A1(n9843), .A2(n6554), .ZN(n6555) );
  NAND2_X1 U8268 ( .A1(n6556), .A2(n6555), .ZN(n6611) );
  OAI21_X1 U8269 ( .B1(n6556), .B2(n6555), .A(n6611), .ZN(n6557) );
  AND2_X1 U8270 ( .A1(P1_U3084), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n7439) );
  AOI21_X1 U8271 ( .B1(n9868), .B2(n6557), .A(n7439), .ZN(n6559) );
  NAND2_X1 U8272 ( .A1(n9860), .A2(n6620), .ZN(n6558) );
  OAI211_X1 U8273 ( .C1(n9873), .C2(n6560), .A(n6559), .B(n6558), .ZN(n6561)
         );
  AOI21_X1 U8274 ( .B1(n6562), .B2(n9869), .A(n6561), .ZN(n6563) );
  INV_X1 U8275 ( .A(n6563), .ZN(P1_U3252) );
  INV_X1 U8276 ( .A(n6564), .ZN(n6596) );
  AOI22_X1 U8277 ( .A1(n7216), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_15__SCAN_IN), .B2(n8588), .ZN(n6565) );
  OAI21_X1 U8278 ( .B1(n6596), .B2(n6195), .A(n6565), .ZN(P2_U3343) );
  INV_X1 U8279 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n6576) );
  NAND2_X1 U8280 ( .A1(n6754), .A2(n6686), .ZN(n6566) );
  NAND2_X1 U8281 ( .A1(n6666), .A2(n6627), .ZN(n7871) );
  NAND2_X1 U8282 ( .A1(n7871), .A2(n7891), .ZN(n8010) );
  XOR2_X1 U8283 ( .A(n6626), .B(n8010), .Z(n6660) );
  NAND2_X1 U8284 ( .A1(n6631), .A2(n6630), .ZN(n6569) );
  XNOR2_X1 U8285 ( .A(n6569), .B(n8010), .ZN(n6571) );
  AOI21_X1 U8286 ( .B1(n6571), .B2(n8411), .A(n6570), .ZN(n6657) );
  OAI21_X1 U8287 ( .B1(n6572), .B2(n6655), .A(n7178), .ZN(n6573) );
  NOR2_X1 U8288 ( .A1(n6573), .A2(n6636), .ZN(n6653) );
  AOI21_X1 U8289 ( .B1(n9693), .B2(n6627), .A(n6653), .ZN(n6574) );
  OAI211_X1 U8290 ( .C1(n6660), .C2(n8549), .A(n6657), .B(n6574), .ZN(n6577)
         );
  NAND2_X1 U8291 ( .A1(n6577), .A2(n4314), .ZN(n6575) );
  OAI21_X1 U8292 ( .B1(n4314), .B2(n6576), .A(n6575), .ZN(P2_U3466) );
  INV_X1 U8293 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6579) );
  NAND2_X1 U8294 ( .A1(n6577), .A2(n10048), .ZN(n6578) );
  OAI21_X1 U8295 ( .B1(n10048), .B2(n6579), .A(n6578), .ZN(P2_U3525) );
  INV_X1 U8296 ( .A(n6803), .ZN(n6595) );
  AOI21_X1 U8297 ( .B1(n6587), .B2(P2_REG1_REG_11__SCAN_IN), .A(n6580), .ZN(
        n6583) );
  INV_X1 U8298 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n6581) );
  MUX2_X1 U8299 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n6581), .S(n6803), .Z(n6582)
         );
  NAND2_X1 U8300 ( .A1(n6582), .A2(n6583), .ZN(n6805) );
  OAI21_X1 U8301 ( .B1(n6583), .B2(n6582), .A(n6805), .ZN(n6586) );
  AND2_X1 U8302 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3152), .ZN(n7261) );
  INV_X1 U8303 ( .A(n9985), .ZN(n9656) );
  INV_X1 U8304 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n6584) );
  NOR2_X1 U8305 ( .A1(n9656), .A2(n6584), .ZN(n6585) );
  AOI211_X1 U8306 ( .C1(n9979), .C2(n6586), .A(n7261), .B(n6585), .ZN(n6594)
         );
  OR2_X1 U8307 ( .A1(n6587), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n6590) );
  INV_X1 U8308 ( .A(n6588), .ZN(n6589) );
  INV_X1 U8309 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n6591) );
  MUX2_X1 U8310 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n6591), .S(n6803), .Z(n6592)
         );
  OAI211_X1 U8311 ( .C1(n4402), .C2(n6592), .A(n9980), .B(n6798), .ZN(n6593)
         );
  OAI211_X1 U8312 ( .C1(n9981), .C2(n6595), .A(n6594), .B(n6593), .ZN(P2_U3257) );
  OAI222_X1 U8313 ( .A1(n7729), .A2(n6597), .B1(n9420), .B2(n6596), .C1(n9009), 
        .C2(P1_U3084), .ZN(P1_U3338) );
  NAND2_X1 U8314 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(n8085), .ZN(n6598) );
  OAI21_X1 U8315 ( .B1(n8247), .B2(n8085), .A(n6598), .ZN(P2_U3581) );
  OAI21_X1 U8316 ( .B1(n6601), .B2(n5557), .A(n6600), .ZN(n7241) );
  INV_X1 U8317 ( .A(n7098), .ZN(n6603) );
  INV_X1 U8318 ( .A(n6738), .ZN(n6602) );
  AOI211_X1 U8319 ( .C1(n6879), .C2(n6603), .A(n9263), .B(n6602), .ZN(n7240)
         );
  XNOR2_X1 U8320 ( .A(n8941), .B(n5557), .ZN(n6605) );
  OAI222_X1 U8321 ( .A1(n9887), .A2(n6977), .B1(n9889), .B2(n6606), .C1(n9732), 
        .C2(n6605), .ZN(n7236) );
  AOI211_X1 U8322 ( .C1(n9957), .C2(n7241), .A(n7240), .B(n7236), .ZN(n6609)
         );
  AOI22_X1 U8323 ( .A1(n9284), .A2(n6879), .B1(n9975), .B2(
        P1_REG1_REG_2__SCAN_IN), .ZN(n6607) );
  OAI21_X1 U8324 ( .B1(n6609), .B2(n9975), .A(n6607), .ZN(P1_U3525) );
  AOI22_X1 U8325 ( .A1(n9365), .A2(n6879), .B1(n9966), .B2(
        P1_REG0_REG_2__SCAN_IN), .ZN(n6608) );
  OAI21_X1 U8326 ( .B1(n6609), .B2(n9966), .A(n6608), .ZN(P1_U3460) );
  INV_X1 U8327 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n6625) );
  INV_X1 U8328 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n6610) );
  MUX2_X1 U8329 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n6610), .S(n6776), .Z(n6613)
         );
  OAI21_X1 U8330 ( .B1(n6613), .B2(n6612), .A(n6775), .ZN(n6614) );
  NAND2_X1 U8331 ( .A1(n9868), .A2(n6614), .ZN(n6616) );
  NAND2_X1 U8332 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3084), .ZN(n6615) );
  NAND2_X1 U8333 ( .A1(n6616), .A2(n6615), .ZN(n6617) );
  AOI21_X1 U8334 ( .B1(n6776), .B2(n9860), .A(n6617), .ZN(n6624) );
  INV_X1 U8335 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n6618) );
  XNOR2_X1 U8336 ( .A(n6776), .B(n6618), .ZN(n6622) );
  OAI211_X1 U8337 ( .C1(n6622), .C2(n6621), .A(n9869), .B(n6767), .ZN(n6623)
         );
  OAI211_X1 U8338 ( .C1(n6625), .C2(n9873), .A(n6624), .B(n6623), .ZN(P1_U3253) );
  INV_X1 U8339 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n6640) );
  OR2_X1 U8340 ( .A1(n8010), .A2(n6666), .ZN(n6628) );
  INV_X1 U8341 ( .A(n8079), .ZN(n6918) );
  NAND2_X1 U8342 ( .A1(n6918), .A2(n6907), .ZN(n7897) );
  INV_X1 U8343 ( .A(n6907), .ZN(n6664) );
  NAND2_X1 U8344 ( .A1(n6664), .A2(n8079), .ZN(n7896) );
  INV_X1 U8345 ( .A(n8013), .ZN(n6909) );
  XNOR2_X1 U8346 ( .A(n6910), .B(n6909), .ZN(n6719) );
  OAI21_X1 U8347 ( .B1(n8013), .B2(n6632), .A(n6916), .ZN(n6633) );
  NAND2_X1 U8348 ( .A1(n6633), .A2(n8411), .ZN(n6635) );
  AOI22_X1 U8349 ( .A1(n8441), .A2(n8080), .B1(n8078), .B2(n8440), .ZN(n6634)
         );
  AND2_X1 U8350 ( .A1(n6635), .A2(n6634), .ZN(n6711) );
  OR2_X1 U8351 ( .A1(n6636), .A2(n6664), .ZN(n6637) );
  AND2_X1 U8352 ( .A1(n6912), .A2(n6637), .ZN(n6712) );
  AOI22_X1 U8353 ( .A1(n6712), .A2(n7178), .B1(n9693), .B2(n6907), .ZN(n6638)
         );
  OAI211_X1 U8354 ( .C1(n6719), .C2(n8549), .A(n6711), .B(n6638), .ZN(n6641)
         );
  NAND2_X1 U8355 ( .A1(n6641), .A2(n4314), .ZN(n6639) );
  OAI21_X1 U8356 ( .B1(n4314), .B2(n6640), .A(n6639), .ZN(P2_U3469) );
  NAND2_X1 U8357 ( .A1(n6641), .A2(n10048), .ZN(n6642) );
  OAI21_X1 U8358 ( .B1(n10048), .B2(n6643), .A(n6642), .ZN(P2_U3526) );
  INV_X1 U8359 ( .A(n7450), .ZN(n8447) );
  NOR2_X1 U8360 ( .A1(n6644), .A2(n8425), .ZN(n6751) );
  INV_X1 U8361 ( .A(n6645), .ZN(n6647) );
  NAND2_X1 U8362 ( .A1(n6647), .A2(n6646), .ZN(n6681) );
  OAI21_X2 U8363 ( .B1(n8447), .B2(n6751), .A(n8422), .ZN(n8407) );
  NOR2_X1 U8364 ( .A1(n6123), .A2(n8034), .ZN(n6651) );
  AND2_X1 U8365 ( .A1(n8422), .A2(n8425), .ZN(n8386) );
  AOI22_X1 U8366 ( .A1(n8386), .A2(n6653), .B1(n6652), .B2(n8452), .ZN(n6654)
         );
  OAI21_X1 U8367 ( .B1(n6655), .B2(n8455), .A(n6654), .ZN(n6656) );
  INV_X1 U8368 ( .A(n6656), .ZN(n6659) );
  MUX2_X1 U8369 ( .A(n6249), .B(n6657), .S(n8422), .Z(n6658) );
  OAI211_X1 U8370 ( .C1(n6660), .C2(n8407), .A(n6659), .B(n6658), .ZN(P2_U3291) );
  OAI21_X1 U8371 ( .B1(n6663), .B2(n6662), .A(n6661), .ZN(n6669) );
  INV_X1 U8372 ( .A(n8078), .ZN(n6911) );
  OAI22_X1 U8373 ( .A1(n7826), .A2(n6911), .B1(n6664), .B2(n7843), .ZN(n6668)
         );
  NAND2_X1 U8374 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3152), .ZN(n8115) );
  NAND2_X1 U8375 ( .A1(n7840), .A2(n6713), .ZN(n6665) );
  OAI211_X1 U8376 ( .C1(n7827), .C2(n6666), .A(n8115), .B(n6665), .ZN(n6667)
         );
  AOI211_X1 U8377 ( .C1(n6669), .C2(n7835), .A(n6668), .B(n6667), .ZN(n6670)
         );
  INV_X1 U8378 ( .A(n6670), .ZN(P2_U3241) );
  XNOR2_X1 U8379 ( .A(n6672), .B(n6671), .ZN(n6678) );
  AOI22_X1 U8380 ( .A1(n6673), .A2(n8077), .B1(n7840), .B2(n6914), .ZN(n6677)
         );
  INV_X1 U8381 ( .A(n7020), .ZN(n10014) );
  OAI22_X1 U8382 ( .A1(n7843), .A2(n10014), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5771), .ZN(n6674) );
  AOI21_X1 U8383 ( .B1(n6675), .B2(n8079), .A(n6674), .ZN(n6676) );
  OAI211_X1 U8384 ( .C1(n6678), .C2(n4570), .A(n6677), .B(n6676), .ZN(P2_U3215) );
  INV_X1 U8385 ( .A(n8407), .ZN(n8379) );
  NAND2_X1 U8386 ( .A1(n6679), .A2(n8425), .ZN(n6680) );
  NOR2_X1 U8387 ( .A1(n6681), .A2(n6680), .ZN(n7182) );
  AOI22_X1 U8388 ( .A1(n7182), .A2(n6683), .B1(n6682), .B2(n8452), .ZN(n6685)
         );
  NAND2_X1 U8389 ( .A1(n8463), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6684) );
  OAI211_X1 U8390 ( .C1(n8455), .C2(n6686), .A(n6685), .B(n6684), .ZN(n6687)
         );
  AOI21_X1 U8391 ( .B1(n8379), .B2(n6688), .A(n6687), .ZN(n6689) );
  OAI21_X1 U8392 ( .B1(n8463), .B2(n6690), .A(n6689), .ZN(P2_U3292) );
  INV_X1 U8393 ( .A(n6691), .ZN(n6694) );
  AOI22_X1 U8394 ( .A1(n9028), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n9428), .ZN(n6692) );
  OAI21_X1 U8395 ( .B1(n6694), .B2(n9420), .A(n6692), .ZN(P1_U3337) );
  AOI22_X1 U8396 ( .A1(n8153), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n8583), .ZN(n6693) );
  OAI21_X1 U8397 ( .B1(n6694), .B2(n6195), .A(n6693), .ZN(P2_U3342) );
  OAI21_X1 U8398 ( .B1(n6703), .B2(n6697), .A(n6696), .ZN(n10004) );
  INV_X1 U8399 ( .A(n10004), .ZN(n6710) );
  NAND2_X1 U8400 ( .A1(n7182), .A2(n7178), .ZN(n8332) );
  AND2_X1 U8401 ( .A1(n6701), .A2(n6731), .ZN(n6699) );
  OR2_X1 U8402 ( .A1(n6699), .A2(n6698), .ZN(n10001) );
  OAI22_X1 U8403 ( .A1(n8332), .A2(n10001), .B1(n9654), .B2(n8426), .ZN(n6700)
         );
  AOI21_X1 U8404 ( .B1(n8430), .B2(n6701), .A(n6700), .ZN(n6709) );
  NOR2_X1 U8405 ( .A1(n6703), .A2(n6702), .ZN(n8007) );
  NAND2_X1 U8406 ( .A1(n6703), .A2(n6702), .ZN(n6704) );
  NAND2_X1 U8407 ( .A1(n6704), .A2(n8411), .ZN(n6706) );
  AOI22_X1 U8408 ( .A1(n8441), .A2(n8086), .B1(n8083), .B2(n8440), .ZN(n6705)
         );
  OAI21_X1 U8409 ( .B1(n8007), .B2(n6706), .A(n6705), .ZN(n10002) );
  MUX2_X1 U8410 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n10002), .S(n8422), .Z(n6707)
         );
  INV_X1 U8411 ( .A(n6707), .ZN(n6708) );
  OAI211_X1 U8412 ( .C1(n6710), .C2(n8407), .A(n6709), .B(n6708), .ZN(P2_U3295) );
  MUX2_X1 U8413 ( .A(n6258), .B(n6711), .S(n8422), .Z(n6718) );
  INV_X1 U8414 ( .A(n6712), .ZN(n6715) );
  INV_X1 U8415 ( .A(n6713), .ZN(n6714) );
  OAI22_X1 U8416 ( .A1(n8332), .A2(n6715), .B1(n6714), .B2(n8426), .ZN(n6716)
         );
  AOI21_X1 U8417 ( .B1(n8430), .B2(n6907), .A(n6716), .ZN(n6717) );
  OAI211_X1 U8418 ( .C1(n6719), .C2(n8407), .A(n6718), .B(n6717), .ZN(P2_U3290) );
  INV_X1 U8419 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n9512) );
  NOR2_X1 U8420 ( .A1(n8426), .A2(n9512), .ZN(n6722) );
  OAI22_X1 U8421 ( .A1(n8332), .A2(n6720), .B1(n6234), .B2(n8422), .ZN(n6721)
         );
  AOI211_X1 U8422 ( .C1(n8422), .C2(n6723), .A(n6722), .B(n6721), .ZN(n6727)
         );
  AOI22_X1 U8423 ( .A1(n8379), .A2(n6725), .B1(n8430), .B2(n6724), .ZN(n6726)
         );
  NAND2_X1 U8424 ( .A1(n6727), .A2(n6726), .ZN(P2_U3294) );
  INV_X1 U8425 ( .A(n6728), .ZN(n6734) );
  INV_X1 U8426 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n9663) );
  OAI22_X1 U8427 ( .A1(n8463), .A2(n6729), .B1(n9524), .B2(n8426), .ZN(n6730)
         );
  AOI21_X1 U8428 ( .B1(n8463), .B2(P2_REG2_REG_0__SCAN_IN), .A(n6730), .ZN(
        n6733) );
  OAI21_X1 U8429 ( .B1(n8461), .B2(n8430), .A(n6731), .ZN(n6732) );
  OAI211_X1 U8430 ( .C1(n6734), .C2(n8407), .A(n6733), .B(n6732), .ZN(P2_U3296) );
  OAI21_X1 U8431 ( .B1(n6736), .B2(n6739), .A(n6735), .ZN(n7233) );
  INV_X1 U8432 ( .A(n6853), .ZN(n6737) );
  AOI211_X1 U8433 ( .C1(n6901), .C2(n6738), .A(n9263), .B(n6737), .ZN(n7228)
         );
  XNOR2_X1 U8434 ( .A(n8834), .B(n6739), .ZN(n6740) );
  OAI222_X1 U8435 ( .A1(n9889), .A2(n8940), .B1(n9887), .B2(n6741), .C1(n6740), 
        .C2(n9732), .ZN(n7227) );
  AOI211_X1 U8436 ( .C1(n9957), .C2(n7233), .A(n7228), .B(n7227), .ZN(n6744)
         );
  AOI22_X1 U8437 ( .A1(n9365), .A2(n6901), .B1(n9966), .B2(
        P1_REG0_REG_3__SCAN_IN), .ZN(n6742) );
  OAI21_X1 U8438 ( .B1(n6744), .B2(n9966), .A(n6742), .ZN(P1_U3463) );
  AOI22_X1 U8439 ( .A1(n9284), .A2(n6901), .B1(n9975), .B2(
        P1_REG1_REG_3__SCAN_IN), .ZN(n6743) );
  OAI21_X1 U8440 ( .B1(n6744), .B2(n9975), .A(n6743), .ZN(P1_U3526) );
  INV_X1 U8441 ( .A(n6745), .ZN(n6748) );
  AOI22_X1 U8442 ( .A1(n9039), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n9428), .ZN(n6746) );
  OAI21_X1 U8443 ( .B1(n6748), .B2(n9420), .A(n6746), .ZN(P1_U3336) );
  AOI22_X1 U8444 ( .A1(n8171), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n8588), .ZN(n6747) );
  OAI21_X1 U8445 ( .B1(n6748), .B2(n6195), .A(n6747), .ZN(P2_U3341) );
  OAI21_X1 U8446 ( .B1(n6750), .B2(n8011), .A(n6749), .ZN(n10012) );
  INV_X1 U8447 ( .A(n10012), .ZN(n6765) );
  NAND2_X1 U8448 ( .A1(n8422), .A2(n6751), .ZN(n8458) );
  OAI21_X1 U8449 ( .B1(n7879), .B2(n6753), .A(n6752), .ZN(n6756) );
  OAI22_X1 U8450 ( .A1(n4846), .A2(n8326), .B1(n6754), .B2(n8324), .ZN(n6755)
         );
  AOI21_X1 U8451 ( .B1(n6756), .B2(n8411), .A(n6755), .ZN(n6757) );
  OAI21_X1 U8452 ( .B1(n6765), .B2(n7450), .A(n6757), .ZN(n10010) );
  AOI22_X1 U8453 ( .A1(n10010), .A2(n8422), .B1(n8430), .B2(n6761), .ZN(n6764)
         );
  INV_X1 U8454 ( .A(n6758), .ZN(n6759) );
  AOI21_X1 U8455 ( .B1(n6761), .B2(n6760), .A(n6759), .ZN(n10007) );
  OAI22_X1 U8456 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(n8426), .B1(n8422), .B2(
        n6239), .ZN(n6762) );
  AOI21_X1 U8457 ( .B1(n8461), .B2(n10007), .A(n6762), .ZN(n6763) );
  OAI211_X1 U8458 ( .C1(n6765), .C2(n8458), .A(n6764), .B(n6763), .ZN(P2_U3293) );
  INV_X1 U8459 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n6782) );
  NAND2_X1 U8460 ( .A1(n6776), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n6766) );
  INV_X1 U8461 ( .A(n6770), .ZN(n6772) );
  NAND2_X1 U8462 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n7058), .ZN(n6768) );
  OAI21_X1 U8463 ( .B1(n7058), .B2(P1_REG2_REG_13__SCAN_IN), .A(n6768), .ZN(
        n6771) );
  INV_X1 U8464 ( .A(n6771), .ZN(n6769) );
  AOI211_X1 U8465 ( .C1(n6772), .C2(n6771), .A(n7050), .B(n9847), .ZN(n6773)
         );
  AOI21_X1 U8466 ( .B1(n9860), .B2(n7058), .A(n6773), .ZN(n6781) );
  INV_X1 U8467 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n6774) );
  MUX2_X1 U8468 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n6774), .S(n7058), .Z(n6778)
         );
  OAI21_X1 U8469 ( .B1(n6776), .B2(P1_REG1_REG_12__SCAN_IN), .A(n6775), .ZN(
        n6777) );
  NAND2_X1 U8470 ( .A1(n6777), .A2(n6778), .ZN(n7057) );
  OAI21_X1 U8471 ( .B1(n6778), .B2(n6777), .A(n7057), .ZN(n6779) );
  AND2_X1 U8472 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n7556) );
  AOI21_X1 U8473 ( .B1(n6779), .B2(n9868), .A(n7556), .ZN(n6780) );
  OAI211_X1 U8474 ( .C1(n9873), .C2(n6782), .A(n6781), .B(n6780), .ZN(P1_U3254) );
  OR2_X1 U8475 ( .A1(n6784), .A2(n6783), .ZN(n6792) );
  NAND2_X1 U8476 ( .A1(n9961), .A2(n6792), .ZN(n6892) );
  AND2_X1 U8477 ( .A1(n6892), .A2(n6785), .ZN(n6788) );
  NAND2_X1 U8478 ( .A1(n6786), .A2(n9408), .ZN(n6793) );
  INV_X1 U8479 ( .A(n6793), .ZN(n6787) );
  NAND2_X1 U8480 ( .A1(n6787), .A2(n6792), .ZN(n6895) );
  NAND2_X1 U8481 ( .A1(n6788), .A2(n6895), .ZN(n6979) );
  INV_X1 U8482 ( .A(n6979), .ZN(n6797) );
  INV_X1 U8483 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n9786) );
  NAND2_X1 U8484 ( .A1(n9408), .A2(n8810), .ZN(n6789) );
  NOR2_X1 U8485 ( .A1(n6792), .A2(n6789), .ZN(n6790) );
  NAND2_X1 U8486 ( .A1(n6791), .A2(n9717), .ZN(n6796) );
  NAND2_X1 U8487 ( .A1(n9923), .A2(n9408), .ZN(n8978) );
  OR2_X1 U8488 ( .A1(n6792), .A2(n8978), .ZN(n6897) );
  NOR2_X2 U8489 ( .A1(n6897), .A2(n6898), .ZN(n9707) );
  NOR2_X1 U8490 ( .A1(n6793), .A2(n6792), .ZN(n6794) );
  INV_X2 U8491 ( .A(n8695), .ZN(n8638) );
  AOI22_X1 U8492 ( .A1(n9707), .A2(n9926), .B1(n8638), .B2(n9930), .ZN(n6795)
         );
  OAI211_X1 U8493 ( .C1(n6797), .C2(n9786), .A(n6796), .B(n6795), .ZN(P1_U3230) );
  NAND2_X1 U8494 ( .A1(n6803), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n6799) );
  INV_X1 U8495 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n6800) );
  INV_X1 U8496 ( .A(n6829), .ZN(n6806) );
  AOI22_X1 U8497 ( .A1(n6829), .A2(n6800), .B1(P2_REG2_REG_13__SCAN_IN), .B2(
        n6806), .ZN(n6801) );
  NOR2_X1 U8498 ( .A1(n6802), .A2(n6801), .ZN(n6823) );
  AOI21_X1 U8499 ( .B1(n6802), .B2(n6801), .A(n6823), .ZN(n6815) );
  OR2_X1 U8500 ( .A1(n6803), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n6804) );
  NAND2_X1 U8501 ( .A1(n6805), .A2(n6804), .ZN(n6809) );
  INV_X1 U8502 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n6807) );
  AOI22_X1 U8503 ( .A1(n6829), .A2(P2_REG1_REG_13__SCAN_IN), .B1(n6807), .B2(
        n6806), .ZN(n6808) );
  NAND2_X1 U8504 ( .A1(n6808), .A2(n6809), .ZN(n6828) );
  OAI21_X1 U8505 ( .B1(n6809), .B2(n6808), .A(n6828), .ZN(n6810) );
  INV_X1 U8506 ( .A(n6810), .ZN(n6812) );
  AOI22_X1 U8507 ( .A1(n9985), .A2(P2_ADDR_REG_13__SCAN_IN), .B1(
        P2_REG3_REG_13__SCAN_IN), .B2(P2_U3152), .ZN(n6811) );
  OAI21_X1 U8508 ( .B1(n9983), .B2(n6812), .A(n6811), .ZN(n6813) );
  AOI21_X1 U8509 ( .B1(n6829), .B2(n9674), .A(n6813), .ZN(n6814) );
  OAI21_X1 U8510 ( .B1(n6815), .B2(n8191), .A(n6814), .ZN(P2_U3258) );
  XNOR2_X1 U8511 ( .A(n6816), .B(n6817), .ZN(n6822) );
  INV_X1 U8512 ( .A(n6818), .ZN(n7034) );
  OAI22_X1 U8513 ( .A1(n7825), .A2(n7034), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9590), .ZN(n6820) );
  OAI22_X1 U8514 ( .A1(n6911), .A2(n7827), .B1(n7826), .B2(n7266), .ZN(n6819)
         );
  AOI211_X1 U8515 ( .C1(n7830), .C2(n7120), .A(n6820), .B(n6819), .ZN(n6821)
         );
  OAI21_X1 U8516 ( .B1(n6822), .B2(n4570), .A(n6821), .ZN(P2_U3223) );
  NOR2_X1 U8517 ( .A1(n6829), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n6824) );
  INV_X1 U8518 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n7104) );
  INV_X1 U8519 ( .A(n7108), .ZN(n7105) );
  AOI22_X1 U8520 ( .A1(n7108), .A2(n7104), .B1(P2_REG2_REG_14__SCAN_IN), .B2(
        n7105), .ZN(n6825) );
  NOR2_X1 U8521 ( .A1(n6826), .A2(n6825), .ZN(n7103) );
  AOI21_X1 U8522 ( .B1(n6826), .B2(n6825), .A(n7103), .ZN(n6837) );
  INV_X1 U8523 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n6827) );
  AOI22_X1 U8524 ( .A1(n7108), .A2(P2_REG1_REG_14__SCAN_IN), .B1(n6827), .B2(
        n7105), .ZN(n6831) );
  OAI21_X1 U8525 ( .B1(n6829), .B2(P2_REG1_REG_13__SCAN_IN), .A(n6828), .ZN(
        n6830) );
  NAND2_X1 U8526 ( .A1(n6831), .A2(n6830), .ZN(n7107) );
  OAI21_X1 U8527 ( .B1(n6831), .B2(n6830), .A(n7107), .ZN(n6835) );
  NAND2_X1 U8528 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3152), .ZN(n7467) );
  INV_X1 U8529 ( .A(n7467), .ZN(n6832) );
  AOI21_X1 U8530 ( .B1(n9985), .B2(P2_ADDR_REG_14__SCAN_IN), .A(n6832), .ZN(
        n6833) );
  OAI21_X1 U8531 ( .B1(n9981), .B2(n7105), .A(n6833), .ZN(n6834) );
  AOI21_X1 U8532 ( .B1(n6835), .B2(n9979), .A(n6834), .ZN(n6836) );
  OAI21_X1 U8533 ( .B1(n6837), .B2(n8191), .A(n6836), .ZN(P2_U3259) );
  NAND2_X1 U8534 ( .A1(n6839), .A2(n8904), .ZN(n6840) );
  NAND2_X1 U8535 ( .A1(n6838), .A2(n6840), .ZN(n9915) );
  OAI21_X1 U8536 ( .B1(n6852), .B2(n9909), .A(n9877), .ZN(n6841) );
  OR2_X1 U8537 ( .A1(n6841), .A2(n7082), .ZN(n9904) );
  NAND2_X1 U8538 ( .A1(n8998), .A2(n9925), .ZN(n9907) );
  OAI211_X1 U8539 ( .C1(n9915), .C2(n9354), .A(n9904), .B(n9907), .ZN(n6846)
         );
  XNOR2_X1 U8540 ( .A(n7084), .B(n8904), .ZN(n6843) );
  NAND2_X1 U8541 ( .A1(n6843), .A2(n9892), .ZN(n6845) );
  NAND2_X1 U8542 ( .A1(n9000), .A2(n9730), .ZN(n6844) );
  NAND2_X1 U8543 ( .A1(n6845), .A2(n6844), .ZN(n9916) );
  NOR2_X1 U8544 ( .A1(n6846), .A2(n9916), .ZN(n6849) );
  AOI22_X1 U8545 ( .A1(n9284), .A2(n6962), .B1(n9975), .B2(
        P1_REG1_REG_5__SCAN_IN), .ZN(n6847) );
  OAI21_X1 U8546 ( .B1(n6849), .B2(n9975), .A(n6847), .ZN(P1_U3528) );
  AOI22_X1 U8547 ( .A1(n9365), .A2(n6962), .B1(n9966), .B2(
        P1_REG0_REG_5__SCAN_IN), .ZN(n6848) );
  OAI21_X1 U8548 ( .B1(n6849), .B2(n9966), .A(n6848), .ZN(P1_U3469) );
  OAI21_X1 U8549 ( .B1(n6851), .B2(n8902), .A(n6850), .ZN(n7252) );
  AOI211_X1 U8550 ( .C1(n6935), .C2(n6853), .A(n9263), .B(n6852), .ZN(n7251)
         );
  XNOR2_X1 U8551 ( .A(n6854), .B(n8902), .ZN(n6855) );
  OAI222_X1 U8552 ( .A1(n9887), .A2(n7087), .B1(n9889), .B2(n6977), .C1(n6855), 
        .C2(n9732), .ZN(n7245) );
  AOI211_X1 U8553 ( .C1(n9957), .C2(n7252), .A(n7251), .B(n7245), .ZN(n6858)
         );
  AOI22_X1 U8554 ( .A1(n9365), .A2(n6935), .B1(n9966), .B2(
        P1_REG0_REG_4__SCAN_IN), .ZN(n6856) );
  OAI21_X1 U8555 ( .B1(n6858), .B2(n9966), .A(n6856), .ZN(P1_U3466) );
  AOI22_X1 U8556 ( .A1(n9284), .A2(n6935), .B1(n9975), .B2(
        P1_REG1_REG_4__SCAN_IN), .ZN(n6857) );
  OAI21_X1 U8557 ( .B1(n6858), .B2(n9975), .A(n6857), .ZN(P1_U3527) );
  NAND2_X1 U8558 ( .A1(n6860), .A2(n7736), .ZN(n6862) );
  NAND2_X1 U8559 ( .A1(n6863), .A2(n7146), .ZN(n6867) );
  NAND2_X1 U8560 ( .A1(n6864), .A2(n6865), .ZN(n6866) );
  NAND2_X1 U8561 ( .A1(n6867), .A2(n6866), .ZN(n6868) );
  NAND2_X1 U8562 ( .A1(n6871), .A2(n6872), .ZN(n6966) );
  NAND2_X1 U8563 ( .A1(n9926), .A2(n7733), .ZN(n6870) );
  NAND2_X1 U8564 ( .A1(n9941), .A2(n7146), .ZN(n6869) );
  NAND2_X1 U8565 ( .A1(n6870), .A2(n6869), .ZN(n6969) );
  NAND2_X1 U8566 ( .A1(n6966), .A2(n6969), .ZN(n6875) );
  NAND2_X1 U8567 ( .A1(n6875), .A2(n6967), .ZN(n6974) );
  NAND2_X1 U8568 ( .A1(n9002), .A2(n7146), .ZN(n6877) );
  NAND2_X1 U8569 ( .A1(n6879), .A2(n6865), .ZN(n6876) );
  NAND2_X1 U8570 ( .A1(n6877), .A2(n6876), .ZN(n6878) );
  AND2_X1 U8571 ( .A1(n6879), .A2(n7146), .ZN(n6880) );
  AOI21_X1 U8572 ( .B1(n9002), .B2(n7733), .A(n6880), .ZN(n6881) );
  INV_X1 U8573 ( .A(n6881), .ZN(n6884) );
  INV_X1 U8574 ( .A(n6882), .ZN(n6883) );
  NAND2_X1 U8575 ( .A1(n9001), .A2(n7146), .ZN(n6886) );
  NAND2_X1 U8576 ( .A1(n6901), .A2(n6865), .ZN(n6885) );
  NAND2_X1 U8577 ( .A1(n6886), .A2(n6885), .ZN(n6887) );
  XNOR2_X1 U8578 ( .A(n6887), .B(n7673), .ZN(n6927) );
  AND2_X1 U8579 ( .A1(n6901), .A2(n7146), .ZN(n6888) );
  AOI21_X1 U8580 ( .B1(n9001), .B2(n7733), .A(n6888), .ZN(n6926) );
  INV_X1 U8581 ( .A(n6926), .ZN(n6928) );
  XNOR2_X1 U8582 ( .A(n6927), .B(n6928), .ZN(n6889) );
  XNOR2_X1 U8583 ( .A(n6932), .B(n6889), .ZN(n6905) );
  AND3_X1 U8584 ( .A1(n6891), .A2(n6450), .A3(n6890), .ZN(n6893) );
  NAND2_X1 U8585 ( .A1(n6893), .A2(n6892), .ZN(n6894) );
  NAND2_X1 U8586 ( .A1(n6894), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6896) );
  INV_X1 U8587 ( .A(n6897), .ZN(n6899) );
  NAND2_X1 U8588 ( .A1(n6899), .A2(n6898), .ZN(n9709) );
  AOI22_X1 U8589 ( .A1(n8669), .A2(n9002), .B1(n9707), .B2(n9000), .ZN(n6903)
         );
  AOI21_X1 U8590 ( .B1(n8638), .B2(n6901), .A(n6900), .ZN(n6902) );
  OAI211_X1 U8591 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n9722), .A(n6903), .B(
        n6902), .ZN(n6904) );
  AOI21_X1 U8592 ( .B1(n6905), .B2(n9717), .A(n6904), .ZN(n6906) );
  INV_X1 U8593 ( .A(n6906), .ZN(P1_U3216) );
  AND2_X1 U8594 ( .A1(n6907), .A2(n8079), .ZN(n6908) );
  OR2_X1 U8595 ( .A1(n7020), .A2(n6911), .ZN(n7900) );
  AND2_X1 U8596 ( .A1(n7020), .A2(n6911), .ZN(n7026) );
  INV_X1 U8597 ( .A(n7026), .ZN(n7915) );
  XNOR2_X1 U8598 ( .A(n7019), .B(n7018), .ZN(n10018) );
  OR2_X1 U8599 ( .A1(n6912), .A2(n7020), .ZN(n7033) );
  NAND2_X1 U8600 ( .A1(n6912), .A2(n7020), .ZN(n6913) );
  NAND2_X1 U8601 ( .A1(n7033), .A2(n6913), .ZN(n10015) );
  AOI22_X1 U8602 ( .A1(n8430), .A2(n7020), .B1(n8452), .B2(n6914), .ZN(n6915)
         );
  OAI21_X1 U8603 ( .B1(n8332), .B2(n10015), .A(n6915), .ZN(n6920) );
  INV_X1 U8604 ( .A(n8077), .ZN(n7127) );
  XNOR2_X1 U8605 ( .A(n7027), .B(n7018), .ZN(n6917) );
  OAI222_X1 U8606 ( .A1(n8324), .A2(n7127), .B1(n8326), .B2(n6918), .C1(n6917), 
        .C2(n8444), .ZN(n10016) );
  MUX2_X1 U8607 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n10016), .S(n8422), .Z(n6919)
         );
  AOI211_X1 U8608 ( .C1(n8379), .C2(n10018), .A(n6920), .B(n6919), .ZN(n6921)
         );
  INV_X1 U8609 ( .A(n6921), .ZN(P2_U3289) );
  NAND2_X1 U8610 ( .A1(n9000), .A2(n7146), .ZN(n6923) );
  NAND2_X1 U8611 ( .A1(n6935), .A2(n6865), .ZN(n6922) );
  NAND2_X1 U8612 ( .A1(n6923), .A2(n6922), .ZN(n6924) );
  AND2_X1 U8613 ( .A1(n6935), .A2(n7146), .ZN(n6925) );
  AOI21_X1 U8614 ( .B1(n9000), .B2(n7733), .A(n6925), .ZN(n6946) );
  XNOR2_X1 U8615 ( .A(n6948), .B(n6946), .ZN(n6944) );
  AND2_X1 U8616 ( .A1(n6927), .A2(n6926), .ZN(n6931) );
  INV_X1 U8617 ( .A(n6927), .ZN(n6929) );
  NAND2_X1 U8618 ( .A1(n6929), .A2(n6928), .ZN(n6930) );
  XNOR2_X1 U8619 ( .A(n6944), .B(n6945), .ZN(n6940) );
  INV_X1 U8620 ( .A(n6933), .ZN(n6934) );
  AOI21_X1 U8621 ( .B1(n8638), .B2(n6935), .A(n6934), .ZN(n6937) );
  NAND2_X1 U8622 ( .A1(n9707), .A2(n8999), .ZN(n6936) );
  OAI211_X1 U8623 ( .C1(n6977), .C2(n9709), .A(n6937), .B(n6936), .ZN(n6938)
         );
  AOI21_X1 U8624 ( .B1(n8692), .B2(n7247), .A(n6938), .ZN(n6939) );
  OAI21_X1 U8625 ( .B1(n6940), .B2(n8683), .A(n6939), .ZN(P1_U3228) );
  INV_X1 U8626 ( .A(n6941), .ZN(n6983) );
  AOI22_X1 U8627 ( .A1(n8182), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n8588), .ZN(n6942) );
  OAI21_X1 U8628 ( .B1(n6983), .B2(n6195), .A(n6942), .ZN(P2_U3340) );
  INV_X1 U8629 ( .A(n9905), .ZN(n6965) );
  AND2_X1 U8630 ( .A1(n6962), .A2(n7146), .ZN(n6943) );
  AOI21_X1 U8631 ( .B1(n8999), .B2(n7733), .A(n6943), .ZN(n6957) );
  INV_X1 U8632 ( .A(n6946), .ZN(n6947) );
  INV_X1 U8633 ( .A(n6955), .ZN(n6953) );
  NAND2_X1 U8634 ( .A1(n8999), .A2(n7666), .ZN(n6950) );
  NAND2_X1 U8635 ( .A1(n6962), .A2(n6865), .ZN(n6949) );
  NAND2_X1 U8636 ( .A1(n6950), .A2(n6949), .ZN(n6951) );
  XNOR2_X1 U8637 ( .A(n6951), .B(n7736), .ZN(n6954) );
  OAI21_X1 U8638 ( .B1(n6957), .B2(n6956), .A(n6992), .ZN(n6958) );
  NAND2_X1 U8639 ( .A1(n6958), .A2(n9717), .ZN(n6964) );
  NAND2_X1 U8640 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n9815) );
  INV_X1 U8641 ( .A(n9815), .ZN(n6959) );
  AOI21_X1 U8642 ( .B1(n8669), .B2(n9000), .A(n6959), .ZN(n6960) );
  OAI21_X1 U8643 ( .B1(n7314), .B2(n8689), .A(n6960), .ZN(n6961) );
  AOI21_X1 U8644 ( .B1(n6962), .B2(n8638), .A(n6961), .ZN(n6963) );
  OAI211_X1 U8645 ( .C1(n9722), .C2(n6965), .A(n6964), .B(n6963), .ZN(P1_U3225) );
  NAND2_X1 U8646 ( .A1(n6967), .A2(n6966), .ZN(n6968) );
  XOR2_X1 U8647 ( .A(n6969), .B(n6968), .Z(n6973) );
  INV_X1 U8648 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n7724) );
  AOI22_X1 U8649 ( .A1(n8669), .A2(n6454), .B1(n9941), .B2(n8638), .ZN(n6970)
         );
  OAI21_X1 U8650 ( .B1(n8940), .B2(n8689), .A(n6970), .ZN(n6971) );
  AOI21_X1 U8651 ( .B1(n6979), .B2(P1_REG3_REG_1__SCAN_IN), .A(n6971), .ZN(
        n6972) );
  OAI21_X1 U8652 ( .B1(n6973), .B2(n8683), .A(n6972), .ZN(P1_U3220) );
  XOR2_X1 U8653 ( .A(n6974), .B(n6975), .Z(n6981) );
  AOI22_X1 U8654 ( .A1(n8669), .A2(n9926), .B1(n6879), .B2(n8638), .ZN(n6976)
         );
  OAI21_X1 U8655 ( .B1(n6977), .B2(n8689), .A(n6976), .ZN(n6978) );
  AOI21_X1 U8656 ( .B1(P1_REG3_REG_2__SCAN_IN), .B2(n6979), .A(n6978), .ZN(
        n6980) );
  OAI21_X1 U8657 ( .B1(n6981), .B2(n8683), .A(n6980), .ZN(P1_U3235) );
  INV_X1 U8658 ( .A(n9859), .ZN(n9037) );
  INV_X1 U8659 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n6982) );
  OAI222_X1 U8660 ( .A1(n9037), .A2(P1_U3084), .B1(n9420), .B2(n6983), .C1(
        n6982), .C2(n7729), .ZN(P1_U3335) );
  INV_X1 U8661 ( .A(n6985), .ZN(n6986) );
  AOI21_X1 U8662 ( .B1(n6984), .B2(n6987), .A(n6986), .ZN(n6991) );
  NAND2_X1 U8663 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3152), .ZN(n8140) );
  OAI21_X1 U8664 ( .B1(n7825), .B2(n7131), .A(n8140), .ZN(n6989) );
  INV_X1 U8665 ( .A(n8075), .ZN(n7175) );
  OAI22_X1 U8666 ( .A1(n7127), .A2(n7827), .B1(n7826), .B2(n7175), .ZN(n6988)
         );
  AOI211_X1 U8667 ( .C1(n7830), .C2(n7184), .A(n6989), .B(n6988), .ZN(n6990)
         );
  OAI21_X1 U8668 ( .B1(n6991), .B2(n4570), .A(n6990), .ZN(P2_U3233) );
  NAND2_X1 U8669 ( .A1(n8998), .A2(n7146), .ZN(n6994) );
  NAND2_X1 U8670 ( .A1(n9276), .A2(n6865), .ZN(n6993) );
  NAND2_X1 U8671 ( .A1(n6994), .A2(n6993), .ZN(n6995) );
  XNOR2_X1 U8672 ( .A(n6995), .B(n7673), .ZN(n6997) );
  AND2_X1 U8673 ( .A1(n9276), .A2(n7146), .ZN(n6996) );
  AOI21_X1 U8674 ( .B1(n8998), .B2(n7733), .A(n6996), .ZN(n6998) );
  AND2_X1 U8675 ( .A1(n6997), .A2(n6998), .ZN(n7065) );
  INV_X1 U8676 ( .A(n7065), .ZN(n7001) );
  INV_X1 U8677 ( .A(n6997), .ZN(n7000) );
  INV_X1 U8678 ( .A(n6998), .ZN(n6999) );
  NAND2_X1 U8679 ( .A1(n7000), .A2(n6999), .ZN(n7066) );
  NAND2_X1 U8680 ( .A1(n7001), .A2(n7066), .ZN(n7002) );
  XNOR2_X1 U8681 ( .A(n7067), .B(n7002), .ZN(n7009) );
  INV_X1 U8682 ( .A(n7003), .ZN(n9273) );
  AOI21_X1 U8683 ( .B1(n8669), .B2(n8999), .A(n7004), .ZN(n7006) );
  NAND2_X1 U8684 ( .A1(n9707), .A2(n8997), .ZN(n7005) );
  OAI211_X1 U8685 ( .C1(n9722), .C2(n9273), .A(n7006), .B(n7005), .ZN(n7007)
         );
  AOI21_X1 U8686 ( .B1(n9276), .B2(n8638), .A(n7007), .ZN(n7008) );
  OAI21_X1 U8687 ( .B1(n7009), .B2(n8683), .A(n7008), .ZN(P1_U3237) );
  XNOR2_X1 U8688 ( .A(n7011), .B(n7010), .ZN(n7017) );
  INV_X1 U8689 ( .A(n7275), .ZN(n7013) );
  OAI22_X1 U8690 ( .A1(n7825), .A2(n7013), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7012), .ZN(n7015) );
  INV_X1 U8691 ( .A(n8074), .ZN(n7265) );
  OAI22_X1 U8692 ( .A1(n7266), .A2(n7827), .B1(n7826), .B2(n7265), .ZN(n7014)
         );
  AOI211_X1 U8693 ( .C1(n7830), .C2(n7389), .A(n7015), .B(n7014), .ZN(n7016)
         );
  OAI21_X1 U8694 ( .B1(n7017), .B2(n4570), .A(n7016), .ZN(P2_U3219) );
  OR2_X1 U8695 ( .A1(n7120), .A2(n7127), .ZN(n7905) );
  NAND2_X1 U8696 ( .A1(n7120), .A2(n7127), .ZN(n7902) );
  NAND2_X1 U8697 ( .A1(n7905), .A2(n7902), .ZN(n7901) );
  NAND2_X1 U8698 ( .A1(n7019), .A2(n7018), .ZN(n7022) );
  OR2_X1 U8699 ( .A1(n7020), .A2(n8078), .ZN(n7021) );
  NAND2_X1 U8700 ( .A1(n7022), .A2(n7021), .ZN(n7023) );
  INV_X1 U8701 ( .A(n7023), .ZN(n7024) );
  INV_X1 U8702 ( .A(n7122), .ZN(n7025) );
  AOI21_X1 U8703 ( .B1(n4839), .B2(n7023), .A(n7025), .ZN(n7031) );
  INV_X1 U8704 ( .A(n7031), .ZN(n7042) );
  XNOR2_X1 U8705 ( .A(n7126), .B(n4839), .ZN(n7029) );
  AOI22_X1 U8706 ( .A1(n8441), .A2(n8078), .B1(n8076), .B2(n8440), .ZN(n7028)
         );
  OAI21_X1 U8707 ( .B1(n7029), .B2(n8444), .A(n7028), .ZN(n7030) );
  AOI21_X1 U8708 ( .B1(n7031), .B2(n8447), .A(n7030), .ZN(n7041) );
  MUX2_X1 U8709 ( .A(n7032), .B(n7041), .S(n8422), .Z(n7038) );
  AOI21_X1 U8710 ( .B1(n7120), .B2(n7033), .A(n7132), .ZN(n7039) );
  INV_X1 U8711 ( .A(n7120), .ZN(n7035) );
  OAI22_X1 U8712 ( .A1(n8455), .A2(n7035), .B1(n8426), .B2(n7034), .ZN(n7036)
         );
  AOI21_X1 U8713 ( .B1(n7039), .B2(n8461), .A(n7036), .ZN(n7037) );
  OAI211_X1 U8714 ( .C1(n7042), .C2(n8458), .A(n7038), .B(n7037), .ZN(P2_U3288) );
  AOI22_X1 U8715 ( .A1(n7039), .A2(n7178), .B1(n9693), .B2(n7120), .ZN(n7040)
         );
  OAI211_X1 U8716 ( .C1(n10006), .C2(n7042), .A(n7041), .B(n7040), .ZN(n7045)
         );
  NAND2_X1 U8717 ( .A1(n7045), .A2(n10048), .ZN(n7043) );
  OAI21_X1 U8718 ( .B1(n10048), .B2(n7044), .A(n7043), .ZN(P2_U3528) );
  INV_X1 U8719 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n7047) );
  NAND2_X1 U8720 ( .A1(n7045), .A2(n4314), .ZN(n7046) );
  OAI21_X1 U8721 ( .B1(n4314), .B2(n7047), .A(n7046), .ZN(P2_U3475) );
  INV_X1 U8722 ( .A(n7048), .ZN(n7119) );
  AOI22_X1 U8723 ( .A1(n8283), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_19__SCAN_IN), .B2(n8588), .ZN(n7049) );
  OAI21_X1 U8724 ( .B1(n7119), .B2(n6195), .A(n7049), .ZN(P2_U3339) );
  AOI21_X1 U8725 ( .B1(n7058), .B2(P1_REG2_REG_13__SCAN_IN), .A(n7050), .ZN(
        n7289) );
  XNOR2_X1 U8726 ( .A(n7288), .B(n7289), .ZN(n7052) );
  INV_X1 U8727 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7051) );
  NOR2_X1 U8728 ( .A1(n7051), .A2(n7052), .ZN(n7290) );
  AOI211_X1 U8729 ( .C1(n7052), .C2(n7051), .A(n7290), .B(n9847), .ZN(n7056)
         );
  NOR2_X1 U8730 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7053), .ZN(n8596) );
  INV_X1 U8731 ( .A(n8596), .ZN(n7054) );
  OAI21_X1 U8732 ( .B1(n9023), .B2(n7288), .A(n7054), .ZN(n7055) );
  NOR2_X1 U8733 ( .A1(n7056), .A2(n7055), .ZN(n7064) );
  INV_X1 U8734 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n7059) );
  MUX2_X1 U8735 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n7059), .S(n7295), .Z(n7060)
         );
  OAI21_X1 U8736 ( .B1(n7061), .B2(n7060), .A(n7294), .ZN(n7062) );
  AOI22_X1 U8737 ( .A1(n9854), .A2(P1_ADDR_REG_14__SCAN_IN), .B1(n7062), .B2(
        n9868), .ZN(n7063) );
  NAND2_X1 U8738 ( .A1(n7064), .A2(n7063), .ZN(P1_U3255) );
  AOI21_X1 U8739 ( .B1(n7067), .B2(n7066), .A(n7065), .ZN(n7140) );
  NAND2_X1 U8740 ( .A1(n8997), .A2(n7146), .ZN(n7069) );
  NAND2_X1 U8741 ( .A1(n7308), .A2(n6865), .ZN(n7068) );
  NAND2_X1 U8742 ( .A1(n7069), .A2(n7068), .ZN(n7070) );
  XNOR2_X1 U8743 ( .A(n7070), .B(n7673), .ZN(n7141) );
  AND2_X1 U8744 ( .A1(n7308), .A2(n7146), .ZN(n7071) );
  AOI21_X1 U8745 ( .B1(n8997), .B2(n7733), .A(n7071), .ZN(n7138) );
  INV_X1 U8746 ( .A(n7138), .ZN(n7142) );
  XNOR2_X1 U8747 ( .A(n7141), .B(n7142), .ZN(n7072) );
  XNOR2_X1 U8748 ( .A(n7140), .B(n7072), .ZN(n7079) );
  INV_X1 U8749 ( .A(n7307), .ZN(n7076) );
  AOI21_X1 U8750 ( .B1(n8669), .B2(n8998), .A(n7073), .ZN(n7075) );
  NAND2_X1 U8751 ( .A1(n9707), .A2(n8996), .ZN(n7074) );
  OAI211_X1 U8752 ( .C1(n9722), .C2(n7076), .A(n7075), .B(n7074), .ZN(n7077)
         );
  AOI21_X1 U8753 ( .B1(n7308), .B2(n8638), .A(n7077), .ZN(n7078) );
  OAI21_X1 U8754 ( .B1(n7079), .B2(n8683), .A(n7078), .ZN(P1_U3211) );
  OAI21_X1 U8755 ( .B1(n4404), .B2(n8906), .A(n7080), .ZN(n9278) );
  OR2_X1 U8756 ( .A1(n7082), .A2(n7081), .ZN(n7083) );
  AND3_X1 U8757 ( .A1(n7304), .A2(n7083), .A3(n9877), .ZN(n9279) );
  AOI21_X1 U8758 ( .B1(n7084), .B2(n8835), .A(n8842), .ZN(n7085) );
  INV_X1 U8759 ( .A(n8906), .ZN(n8702) );
  XNOR2_X1 U8760 ( .A(n7085), .B(n8702), .ZN(n7086) );
  OAI222_X1 U8761 ( .A1(n9887), .A2(n7088), .B1(n9889), .B2(n7087), .C1(n7086), 
        .C2(n9732), .ZN(n9271) );
  AOI211_X1 U8762 ( .C1(n9957), .C2(n9278), .A(n9279), .B(n9271), .ZN(n7091)
         );
  AOI22_X1 U8763 ( .A1(n9365), .A2(n9276), .B1(n9966), .B2(
        P1_REG0_REG_6__SCAN_IN), .ZN(n7089) );
  OAI21_X1 U8764 ( .B1(n7091), .B2(n9966), .A(n7089), .ZN(P1_U3472) );
  AOI22_X1 U8765 ( .A1(n9284), .A2(n9276), .B1(n9975), .B2(
        P1_REG1_REG_6__SCAN_IN), .ZN(n7090) );
  OAI21_X1 U8766 ( .B1(n7091), .B2(n9975), .A(n7090), .ZN(P1_U3529) );
  OAI21_X1 U8767 ( .B1(n5556), .B2(n7093), .A(n7092), .ZN(n9947) );
  XNOR2_X1 U8768 ( .A(n5556), .B(n4461), .ZN(n7094) );
  NAND2_X1 U8769 ( .A1(n7094), .A2(n9892), .ZN(n7096) );
  AOI22_X1 U8770 ( .A1(n9730), .A2(n6454), .B1(n9002), .B2(n9925), .ZN(n7095)
         );
  NAND2_X1 U8771 ( .A1(n7096), .A2(n7095), .ZN(n9950) );
  NAND2_X1 U8772 ( .A1(n9941), .A2(n9930), .ZN(n7097) );
  NAND2_X1 U8773 ( .A1(n7097), .A2(n9877), .ZN(n7099) );
  OR2_X1 U8774 ( .A1(n7099), .A2(n7098), .ZN(n9944) );
  OAI22_X1 U8775 ( .A1(n9944), .A2(n9920), .B1(n7724), .B2(n9272), .ZN(n7100)
         );
  OAI21_X1 U8776 ( .B1(n9950), .B2(n7100), .A(n9918), .ZN(n7102) );
  INV_X1 U8777 ( .A(n9899), .ZN(n9737) );
  AOI22_X1 U8778 ( .A1(n9737), .A2(n9941), .B1(n9938), .B2(
        P1_REG2_REG_1__SCAN_IN), .ZN(n7101) );
  OAI211_X1 U8779 ( .C1(n9253), .C2(n9947), .A(n7102), .B(n7101), .ZN(P1_U3290) );
  XNOR2_X1 U8780 ( .A(n7215), .B(n7216), .ZN(n7106) );
  NOR2_X1 U8781 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n7106), .ZN(n7217) );
  AOI21_X1 U8782 ( .B1(n7106), .B2(P2_REG2_REG_15__SCAN_IN), .A(n7217), .ZN(
        n7117) );
  OAI21_X1 U8783 ( .B1(n7108), .B2(P2_REG1_REG_14__SCAN_IN), .A(n7107), .ZN(
        n7207) );
  INV_X1 U8784 ( .A(n7216), .ZN(n7208) );
  XNOR2_X1 U8785 ( .A(n7207), .B(n7208), .ZN(n7109) );
  INV_X1 U8786 ( .A(n7109), .ZN(n7112) );
  INV_X1 U8787 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n7110) );
  NOR2_X1 U8788 ( .A1(n7110), .A2(n7109), .ZN(n7209) );
  INV_X1 U8789 ( .A(n7209), .ZN(n7111) );
  OAI211_X1 U8790 ( .C1(n7112), .C2(P2_REG1_REG_15__SCAN_IN), .A(n9979), .B(
        n7111), .ZN(n7116) );
  NAND2_X1 U8791 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(P2_U3152), .ZN(n7568) );
  INV_X1 U8792 ( .A(n7568), .ZN(n7114) );
  NOR2_X1 U8793 ( .A1(n9981), .A2(n7208), .ZN(n7113) );
  AOI211_X1 U8794 ( .C1(P2_ADDR_REG_15__SCAN_IN), .C2(n9985), .A(n7114), .B(
        n7113), .ZN(n7115) );
  OAI211_X1 U8795 ( .C1(n7117), .C2(n8191), .A(n7116), .B(n7115), .ZN(P2_U3260) );
  OAI222_X1 U8796 ( .A1(P1_U3084), .A2(n9911), .B1(n9420), .B2(n7119), .C1(
        n7118), .C2(n7729), .ZN(P1_U3334) );
  OR2_X1 U8797 ( .A1(n7184), .A2(n7266), .ZN(n7904) );
  NAND2_X1 U8798 ( .A1(n7184), .A2(n7266), .ZN(n7909) );
  NAND2_X1 U8799 ( .A1(n7120), .A2(n8077), .ZN(n7121) );
  INV_X1 U8800 ( .A(n7186), .ZN(n7124) );
  AOI21_X1 U8801 ( .B1(n8016), .B2(n7125), .A(n7124), .ZN(n10020) );
  XNOR2_X1 U8802 ( .A(n7174), .B(n8016), .ZN(n7129) );
  OAI22_X1 U8803 ( .A1(n7127), .A2(n8326), .B1(n7175), .B2(n8324), .ZN(n7128)
         );
  AOI21_X1 U8804 ( .B1(n7129), .B2(n8411), .A(n7128), .ZN(n7130) );
  OAI21_X1 U8805 ( .B1(n10020), .B2(n7450), .A(n7130), .ZN(n10024) );
  NAND2_X1 U8806 ( .A1(n10024), .A2(n8422), .ZN(n7137) );
  OAI22_X1 U8807 ( .A1(n8422), .A2(n6367), .B1(n7131), .B2(n8426), .ZN(n7135)
         );
  INV_X1 U8808 ( .A(n7184), .ZN(n10021) );
  AND2_X1 U8809 ( .A1(n7132), .A2(n10021), .ZN(n7272) );
  NOR2_X1 U8810 ( .A1(n7132), .A2(n10021), .ZN(n7133) );
  OR2_X1 U8811 ( .A1(n7272), .A2(n7133), .ZN(n10023) );
  NOR2_X1 U8812 ( .A1(n10023), .A2(n8332), .ZN(n7134) );
  AOI211_X1 U8813 ( .C1(n8430), .C2(n7184), .A(n7135), .B(n7134), .ZN(n7136)
         );
  OAI211_X1 U8814 ( .C1(n10020), .C2(n8458), .A(n7137), .B(n7136), .ZN(
        P2_U3287) );
  NAND2_X1 U8815 ( .A1(n7141), .A2(n7138), .ZN(n7139) );
  NAND2_X1 U8816 ( .A1(n7140), .A2(n7139), .ZN(n7145) );
  INV_X1 U8817 ( .A(n7141), .ZN(n7143) );
  NAND2_X1 U8818 ( .A1(n7143), .A2(n7142), .ZN(n7144) );
  NAND2_X1 U8819 ( .A1(n7145), .A2(n7144), .ZN(n7326) );
  NAND2_X1 U8820 ( .A1(n8996), .A2(n7733), .ZN(n7148) );
  NAND2_X1 U8821 ( .A1(n7357), .A2(n7666), .ZN(n7147) );
  NAND2_X1 U8822 ( .A1(n7148), .A2(n7147), .ZN(n7325) );
  NAND2_X1 U8823 ( .A1(n8996), .A2(n7146), .ZN(n7150) );
  NAND2_X1 U8824 ( .A1(n7357), .A2(n6865), .ZN(n7149) );
  NAND2_X1 U8825 ( .A1(n7150), .A2(n7149), .ZN(n7151) );
  XNOR2_X1 U8826 ( .A(n7151), .B(n7736), .ZN(n7324) );
  XOR2_X1 U8827 ( .A(n7325), .B(n7324), .Z(n7152) );
  XNOR2_X1 U8828 ( .A(n7326), .B(n7152), .ZN(n7159) );
  INV_X1 U8829 ( .A(n7201), .ZN(n7156) );
  NOR2_X1 U8830 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7153), .ZN(n9820) );
  AOI21_X1 U8831 ( .B1(n8669), .B2(n8997), .A(n9820), .ZN(n7155) );
  NAND2_X1 U8832 ( .A1(n9707), .A2(n8995), .ZN(n7154) );
  OAI211_X1 U8833 ( .C1(n9722), .C2(n7156), .A(n7155), .B(n7154), .ZN(n7157)
         );
  AOI21_X1 U8834 ( .B1(n7357), .B2(n8638), .A(n7157), .ZN(n7158) );
  OAI21_X1 U8835 ( .B1(n7159), .B2(n8683), .A(n7158), .ZN(P1_U3219) );
  INV_X1 U8836 ( .A(n7160), .ZN(n7172) );
  AOI22_X1 U8837 ( .A1(n8006), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_20__SCAN_IN), .B2(n8583), .ZN(n7161) );
  OAI21_X1 U8838 ( .B1(n7172), .B2(n6195), .A(n7161), .ZN(P2_U3338) );
  XNOR2_X1 U8839 ( .A(n7162), .B(n7163), .ZN(n7168) );
  INV_X1 U8840 ( .A(n7179), .ZN(n7164) );
  OAI22_X1 U8841 ( .A1(n7825), .A2(n7164), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5838), .ZN(n7166) );
  OAI22_X1 U8842 ( .A1(n7175), .A2(n7827), .B1(n7826), .B2(n7446), .ZN(n7165)
         );
  AOI211_X1 U8843 ( .C1(n7830), .C2(n7338), .A(n7166), .B(n7165), .ZN(n7167)
         );
  OAI21_X1 U8844 ( .B1(n7168), .B2(n4570), .A(n7167), .ZN(P2_U3238) );
  INV_X1 U8845 ( .A(n7169), .ZN(n7731) );
  AOI22_X1 U8846 ( .A1(n7874), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_21__SCAN_IN), .B2(n8583), .ZN(n7170) );
  OAI21_X1 U8847 ( .B1(n7731), .B2(n6195), .A(n7170), .ZN(P2_U3337) );
  OAI222_X1 U8848 ( .A1(n9921), .A2(P1_U3084), .B1(n9420), .B2(n7172), .C1(
        n7171), .C2(n7729), .ZN(P1_U3333) );
  OR2_X1 U8849 ( .A1(n7338), .A2(n7265), .ZN(n7926) );
  AND2_X1 U8850 ( .A1(n7338), .A2(n7265), .ZN(n7344) );
  INV_X1 U8851 ( .A(n7344), .ZN(n7928) );
  NAND2_X1 U8852 ( .A1(n7926), .A2(n7928), .ZN(n8019) );
  INV_X1 U8853 ( .A(n7909), .ZN(n7173) );
  NOR2_X1 U8854 ( .A1(n7389), .A2(n7175), .ZN(n7912) );
  NAND2_X1 U8855 ( .A1(n7389), .A2(n7175), .ZN(n7920) );
  XOR2_X1 U8856 ( .A(n8019), .B(n7345), .Z(n7176) );
  AOI222_X1 U8857 ( .A1(n8411), .A2(n7176), .B1(n8073), .B2(n8440), .C1(n8075), 
        .C2(n8441), .ZN(n10030) );
  INV_X1 U8858 ( .A(n7389), .ZN(n7277) );
  NAND2_X1 U8859 ( .A1(n7272), .A2(n7277), .ZN(n7177) );
  INV_X1 U8860 ( .A(n7177), .ZN(n7273) );
  INV_X1 U8861 ( .A(n7338), .ZN(n10032) );
  OAI211_X1 U8862 ( .C1(n7273), .C2(n10032), .A(n7178), .B(n7340), .ZN(n10029)
         );
  INV_X1 U8863 ( .A(n10029), .ZN(n7183) );
  AOI22_X1 U8864 ( .A1(n8463), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n7179), .B2(
        n8452), .ZN(n7180) );
  OAI21_X1 U8865 ( .B1(n10032), .B2(n8455), .A(n7180), .ZN(n7181) );
  AOI21_X1 U8866 ( .B1(n7183), .B2(n7182), .A(n7181), .ZN(n7189) );
  OR2_X1 U8867 ( .A1(n7184), .A2(n8076), .ZN(n7185) );
  AND2_X2 U8868 ( .A1(n7186), .A2(n7185), .ZN(n7268) );
  INV_X1 U8869 ( .A(n7912), .ZN(n7917) );
  NAND2_X1 U8870 ( .A1(n7917), .A2(n7920), .ZN(n8017) );
  NAND2_X1 U8871 ( .A1(n7389), .A2(n8075), .ZN(n7187) );
  XOR2_X1 U8872 ( .A(n7337), .B(n8019), .Z(n10035) );
  NAND2_X1 U8873 ( .A1(n10035), .A2(n8379), .ZN(n7188) );
  OAI211_X1 U8874 ( .C1(n10030), .C2(n8463), .A(n7189), .B(n7188), .ZN(
        P2_U3285) );
  NAND2_X1 U8875 ( .A1(n7191), .A2(n8909), .ZN(n7192) );
  NAND2_X1 U8876 ( .A1(n7190), .A2(n7192), .ZN(n7352) );
  AND2_X1 U8877 ( .A1(n7193), .A2(n9920), .ZN(n7194) );
  NAND2_X1 U8878 ( .A1(n9918), .A2(n7194), .ZN(n9267) );
  AOI22_X1 U8879 ( .A1(n9730), .A2(n8997), .B1(n8995), .B2(n9925), .ZN(n7198)
         );
  AND2_X1 U8880 ( .A1(n7310), .A2(n8710), .ZN(n7196) );
  NAND3_X1 U8881 ( .A1(n7310), .A2(n8828), .A3(n9884), .ZN(n7195) );
  OAI211_X1 U8882 ( .C1(n7196), .C2(n8909), .A(n7195), .B(n9892), .ZN(n7197)
         );
  OAI211_X1 U8883 ( .C1(n7352), .C2(n9946), .A(n7198), .B(n7197), .ZN(n7353)
         );
  NAND2_X1 U8884 ( .A1(n7353), .A2(n9918), .ZN(n7206) );
  INV_X1 U8885 ( .A(n7199), .ZN(n9879) );
  AOI211_X1 U8886 ( .C1(n7357), .C2(n7305), .A(n9263), .B(n9879), .ZN(n7354)
         );
  OR2_X1 U8887 ( .A1(n7200), .A2(n9920), .ZN(n9059) );
  AOI22_X1 U8888 ( .A1(n9938), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n7201), .B2(
        n9896), .ZN(n7202) );
  OAI21_X1 U8889 ( .B1(n7203), .B2(n9899), .A(n7202), .ZN(n7204) );
  AOI21_X1 U8890 ( .B1(n7354), .B2(n9881), .A(n7204), .ZN(n7205) );
  OAI211_X1 U8891 ( .C1(n7352), .C2(n9267), .A(n7206), .B(n7205), .ZN(P1_U3283) );
  NOR2_X1 U8892 ( .A1(n7208), .A2(n7207), .ZN(n7210) );
  NOR2_X1 U8893 ( .A1(n7210), .A2(n7209), .ZN(n7212) );
  XOR2_X1 U8894 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8153), .Z(n7211) );
  NAND2_X1 U8895 ( .A1(n7211), .A2(n7212), .ZN(n8154) );
  OAI21_X1 U8896 ( .B1(n7212), .B2(n7211), .A(n8154), .ZN(n7213) );
  INV_X1 U8897 ( .A(n7213), .ZN(n7226) );
  NOR2_X1 U8898 ( .A1(n9503), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7791) );
  INV_X1 U8899 ( .A(n8153), .ZN(n7220) );
  NOR2_X1 U8900 ( .A1(n9981), .A2(n7220), .ZN(n7214) );
  AOI211_X1 U8901 ( .C1(P2_ADDR_REG_16__SCAN_IN), .C2(n9985), .A(n7791), .B(
        n7214), .ZN(n7225) );
  NOR2_X1 U8902 ( .A1(n7216), .A2(n7215), .ZN(n7218) );
  INV_X1 U8903 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n7221) );
  NAND2_X1 U8904 ( .A1(n8153), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n8150) );
  INV_X1 U8905 ( .A(n8150), .ZN(n7219) );
  AOI21_X1 U8906 ( .B1(n7221), .B2(n7220), .A(n7219), .ZN(n7222) );
  NAND2_X1 U8907 ( .A1(n7222), .A2(n7223), .ZN(n8149) );
  OAI211_X1 U8908 ( .C1(n7223), .C2(n7222), .A(n9980), .B(n8149), .ZN(n7224)
         );
  OAI211_X1 U8909 ( .C1(n7226), .C2(n9983), .A(n7225), .B(n7224), .ZN(P2_U3261) );
  INV_X1 U8910 ( .A(n7227), .ZN(n7235) );
  NAND2_X1 U8911 ( .A1(n7228), .A2(n9881), .ZN(n7230) );
  AOI22_X1 U8912 ( .A1(n9938), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n9896), .B2(
        n4986), .ZN(n7229) );
  OAI211_X1 U8913 ( .C1(n7231), .C2(n9899), .A(n7230), .B(n7229), .ZN(n7232)
         );
  AOI21_X1 U8914 ( .B1(n9277), .B2(n7233), .A(n7232), .ZN(n7234) );
  OAI21_X1 U8915 ( .B1(n7235), .B2(n9938), .A(n7234), .ZN(P1_U3288) );
  INV_X1 U8916 ( .A(n7236), .ZN(n7244) );
  NOR2_X1 U8917 ( .A1(n9899), .A2(n7237), .ZN(n7239) );
  INV_X1 U8918 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n9804) );
  OAI22_X1 U8919 ( .A1(n9918), .A2(n6319), .B1(n9804), .B2(n9272), .ZN(n7238)
         );
  AOI211_X1 U8920 ( .C1(n7240), .C2(n9881), .A(n7239), .B(n7238), .ZN(n7243)
         );
  NAND2_X1 U8921 ( .A1(n7241), .A2(n9277), .ZN(n7242) );
  OAI211_X1 U8922 ( .C1(n7244), .C2(n9938), .A(n7243), .B(n7242), .ZN(P1_U3289) );
  INV_X1 U8923 ( .A(n7245), .ZN(n7255) );
  NOR2_X1 U8924 ( .A1(n9899), .A2(n7246), .ZN(n7250) );
  INV_X1 U8925 ( .A(n7247), .ZN(n7248) );
  OAI22_X1 U8926 ( .A1(n9918), .A2(n6327), .B1(n7248), .B2(n9272), .ZN(n7249)
         );
  AOI211_X1 U8927 ( .C1(n7251), .C2(n9881), .A(n7250), .B(n7249), .ZN(n7254)
         );
  NAND2_X1 U8928 ( .A1(n7252), .A2(n9277), .ZN(n7253) );
  OAI211_X1 U8929 ( .C1(n7255), .C2(n9938), .A(n7254), .B(n7253), .ZN(P1_U3287) );
  INV_X1 U8930 ( .A(n7416), .ZN(n7343) );
  OAI21_X1 U8931 ( .B1(n7258), .B2(n7257), .A(n7256), .ZN(n7259) );
  NAND2_X1 U8932 ( .A1(n7259), .A2(n7835), .ZN(n7263) );
  OAI22_X1 U8933 ( .A1(n7265), .A2(n7827), .B1(n7826), .B2(n7469), .ZN(n7260)
         );
  AOI211_X1 U8934 ( .C1(n7341), .C2(n7840), .A(n7261), .B(n7260), .ZN(n7262)
         );
  OAI211_X1 U8935 ( .C1(n7343), .C2(n7843), .A(n7263), .B(n7262), .ZN(P2_U3226) );
  XNOR2_X1 U8936 ( .A(n7264), .B(n8017), .ZN(n7271) );
  OAI22_X1 U8937 ( .A1(n7266), .A2(n8326), .B1(n7265), .B2(n8324), .ZN(n7270)
         );
  OAI21_X1 U8938 ( .B1(n7268), .B2(n8017), .A(n7267), .ZN(n7393) );
  NOR2_X1 U8939 ( .A1(n7393), .A2(n7450), .ZN(n7269) );
  AOI211_X1 U8940 ( .C1(n7271), .C2(n8411), .A(n7270), .B(n7269), .ZN(n7392)
         );
  INV_X1 U8941 ( .A(n7272), .ZN(n7274) );
  AOI21_X1 U8942 ( .B1(n7389), .B2(n7274), .A(n7273), .ZN(n7390) );
  AOI22_X1 U8943 ( .A1(n8463), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n7275), .B2(
        n8452), .ZN(n7276) );
  OAI21_X1 U8944 ( .B1(n7277), .B2(n8455), .A(n7276), .ZN(n7279) );
  NOR2_X1 U8945 ( .A1(n7393), .A2(n8458), .ZN(n7278) );
  AOI211_X1 U8946 ( .C1(n7390), .C2(n8461), .A(n7279), .B(n7278), .ZN(n7280)
         );
  OAI21_X1 U8947 ( .B1(n7392), .B2(n8463), .A(n7280), .ZN(P2_U3286) );
  XNOR2_X1 U8948 ( .A(n7281), .B(n7282), .ZN(n7287) );
  INV_X1 U8949 ( .A(n7456), .ZN(n7283) );
  OAI22_X1 U8950 ( .A1(n7825), .A2(n7283), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5869), .ZN(n7285) );
  INV_X1 U8951 ( .A(n8071), .ZN(n7570) );
  OAI22_X1 U8952 ( .A1(n7446), .A2(n7827), .B1(n7826), .B2(n7570), .ZN(n7284)
         );
  AOI211_X1 U8953 ( .C1(n7830), .C2(n8550), .A(n7285), .B(n7284), .ZN(n7286)
         );
  OAI21_X1 U8954 ( .B1(n7287), .B2(n4570), .A(n7286), .ZN(P2_U3236) );
  NOR2_X1 U8955 ( .A1(n7289), .A2(n7288), .ZN(n7291) );
  NOR2_X1 U8956 ( .A1(n7291), .A2(n7290), .ZN(n9003) );
  INV_X1 U8957 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n7292) );
  AOI211_X1 U8958 ( .C1(n7293), .C2(n7292), .A(n9004), .B(n9847), .ZN(n7301)
         );
  OAI21_X1 U8959 ( .B1(n7295), .B2(P1_REG1_REG_14__SCAN_IN), .A(n7294), .ZN(
        n9008) );
  XNOR2_X1 U8960 ( .A(n9009), .B(n9008), .ZN(n7297) );
  INV_X1 U8961 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n7296) );
  NOR2_X1 U8962 ( .A1(n7296), .A2(n7297), .ZN(n9010) );
  AOI211_X1 U8963 ( .C1(n7297), .C2(n7296), .A(n9010), .B(n9797), .ZN(n7300)
         );
  NAND2_X1 U8964 ( .A1(n9854), .A2(P1_ADDR_REG_15__SCAN_IN), .ZN(n7298) );
  NAND2_X1 U8965 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9704) );
  OAI211_X1 U8966 ( .C1(n9023), .C2(n9009), .A(n7298), .B(n9704), .ZN(n7299)
         );
  OR3_X1 U8967 ( .A1(n7301), .A2(n7300), .A3(n7299), .ZN(P1_U3256) );
  OAI21_X1 U8968 ( .B1(n7302), .B2(n8908), .A(n7303), .ZN(n9956) );
  INV_X1 U8969 ( .A(n7304), .ZN(n7306) );
  OAI211_X1 U8970 ( .C1(n7306), .C2(n9953), .A(n9877), .B(n7305), .ZN(n9952)
         );
  AOI22_X1 U8971 ( .A1(n9737), .A2(n7308), .B1(n9896), .B2(n7307), .ZN(n7309)
         );
  OAI21_X1 U8972 ( .B1(n9952), .B2(n9059), .A(n7309), .ZN(n7316) );
  INV_X1 U8973 ( .A(n7310), .ZN(n7311) );
  AOI21_X1 U8974 ( .B1(n8908), .B2(n7312), .A(n7311), .ZN(n7313) );
  OAI222_X1 U8975 ( .A1(n9889), .A2(n7314), .B1(n9887), .B2(n9890), .C1(n9732), 
        .C2(n7313), .ZN(n9954) );
  MUX2_X1 U8976 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n9954), .S(n9918), .Z(n7315)
         );
  AOI211_X1 U8977 ( .C1(n9277), .C2(n9956), .A(n7316), .B(n7315), .ZN(n7317)
         );
  INV_X1 U8978 ( .A(n7317), .ZN(P1_U3284) );
  NAND2_X1 U8979 ( .A1(n9875), .A2(n6865), .ZN(n7319) );
  NAND2_X1 U8980 ( .A1(n8995), .A2(n7146), .ZN(n7318) );
  NAND2_X1 U8981 ( .A1(n7319), .A2(n7318), .ZN(n7320) );
  XNOR2_X1 U8982 ( .A(n7320), .B(n7673), .ZN(n7322) );
  AOI22_X1 U8983 ( .A1(n9875), .A2(n7666), .B1(n8995), .B2(n7733), .ZN(n7321)
         );
  NAND2_X1 U8984 ( .A1(n7322), .A2(n7321), .ZN(n7370) );
  OR2_X1 U8985 ( .A1(n7322), .A2(n7321), .ZN(n7323) );
  NAND2_X1 U8986 ( .A1(n7370), .A2(n7323), .ZN(n7331) );
  OAI21_X1 U8987 ( .B1(n7326), .B2(n7325), .A(n7324), .ZN(n7328) );
  NAND2_X1 U8988 ( .A1(n7326), .A2(n7325), .ZN(n7327) );
  NAND2_X1 U8989 ( .A1(n7328), .A2(n7327), .ZN(n7329) );
  INV_X1 U8990 ( .A(n7371), .ZN(n7330) );
  AOI21_X1 U8991 ( .B1(n7331), .B2(n7329), .A(n7330), .ZN(n7336) );
  NAND2_X1 U8992 ( .A1(n8692), .A2(n9897), .ZN(n7333) );
  AND2_X1 U8993 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n9839) );
  AOI21_X1 U8994 ( .B1(n8996), .B2(n8669), .A(n9839), .ZN(n7332) );
  OAI211_X1 U8995 ( .C1(n9888), .C2(n8689), .A(n7333), .B(n7332), .ZN(n7334)
         );
  AOI21_X1 U8996 ( .B1(n9875), .B2(n8638), .A(n7334), .ZN(n7335) );
  OAI21_X1 U8997 ( .B1(n7336), .B2(n8683), .A(n7335), .ZN(P1_U3229) );
  NOR2_X1 U8998 ( .A1(n7416), .A2(n7446), .ZN(n7422) );
  INV_X1 U8999 ( .A(n7422), .ZN(n7930) );
  NAND2_X1 U9000 ( .A1(n7416), .A2(n7446), .ZN(n7929) );
  XOR2_X1 U9001 ( .A(n7417), .B(n8021), .Z(n7363) );
  INV_X1 U9002 ( .A(n7455), .ZN(n7339) );
  AOI21_X1 U9003 ( .B1(n7416), .B2(n7340), .A(n7339), .ZN(n7360) );
  AOI22_X1 U9004 ( .A1(n8463), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n7341), .B2(
        n8452), .ZN(n7342) );
  OAI21_X1 U9005 ( .B1(n7343), .B2(n8455), .A(n7342), .ZN(n7348) );
  OAI21_X2 U9006 ( .B1(n7345), .B2(n7344), .A(n7926), .ZN(n7423) );
  XOR2_X1 U9007 ( .A(n8021), .B(n7423), .Z(n7346) );
  AOI222_X1 U9008 ( .A1(n8411), .A2(n7346), .B1(n8072), .B2(n8440), .C1(n8074), 
        .C2(n8441), .ZN(n7362) );
  NOR2_X1 U9009 ( .A1(n7362), .A2(n8463), .ZN(n7347) );
  AOI211_X1 U9010 ( .C1(n7360), .C2(n8461), .A(n7348), .B(n7347), .ZN(n7349)
         );
  OAI21_X1 U9011 ( .B1(n8407), .B2(n7363), .A(n7349), .ZN(P2_U3284) );
  INV_X1 U9012 ( .A(n7350), .ZN(n7369) );
  AOI22_X1 U9013 ( .A1(n6124), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_22__SCAN_IN), .B2(n8583), .ZN(n7351) );
  OAI21_X1 U9014 ( .B1(n7369), .B2(n6195), .A(n7351), .ZN(P2_U3336) );
  INV_X1 U9015 ( .A(n7352), .ZN(n7355) );
  INV_X1 U9016 ( .A(n9945), .ZN(n9965) );
  AOI211_X1 U9017 ( .C1(n7355), .C2(n9965), .A(n7354), .B(n7353), .ZN(n7359)
         );
  AOI22_X1 U9018 ( .A1(n9284), .A2(n7357), .B1(n9975), .B2(
        P1_REG1_REG_8__SCAN_IN), .ZN(n7356) );
  OAI21_X1 U9019 ( .B1(n7359), .B2(n9975), .A(n7356), .ZN(P1_U3531) );
  AOI22_X1 U9020 ( .A1(n9365), .A2(n7357), .B1(n9966), .B2(
        P1_REG0_REG_8__SCAN_IN), .ZN(n7358) );
  OAI21_X1 U9021 ( .B1(n7359), .B2(n9966), .A(n7358), .ZN(P1_U3478) );
  AOI22_X1 U9022 ( .A1(n7360), .A2(n7178), .B1(n9693), .B2(n7416), .ZN(n7361)
         );
  OAI211_X1 U9023 ( .C1(n8549), .C2(n7363), .A(n7362), .B(n7361), .ZN(n7365)
         );
  NAND2_X1 U9024 ( .A1(n7365), .A2(n10048), .ZN(n7364) );
  OAI21_X1 U9025 ( .B1(n10048), .B2(n6581), .A(n7364), .ZN(P2_U3532) );
  INV_X1 U9026 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n7367) );
  NAND2_X1 U9027 ( .A1(n7365), .A2(n4314), .ZN(n7366) );
  OAI21_X1 U9028 ( .B1(n4314), .B2(n7367), .A(n7366), .ZN(P2_U3487) );
  OAI222_X1 U9029 ( .A1(P1_U3084), .A2(n8813), .B1(n9420), .B2(n7369), .C1(
        n7368), .C2(n7729), .ZN(P1_U3331) );
  NAND2_X1 U9030 ( .A1(n7408), .A2(n6865), .ZN(n7373) );
  NAND2_X1 U9031 ( .A1(n9729), .A2(n7666), .ZN(n7372) );
  NAND2_X1 U9032 ( .A1(n7373), .A2(n7372), .ZN(n7374) );
  XNOR2_X1 U9033 ( .A(n7374), .B(n7736), .ZN(n7377) );
  NAND2_X1 U9034 ( .A1(n7408), .A2(n7146), .ZN(n7376) );
  NAND2_X1 U9035 ( .A1(n9729), .A2(n7733), .ZN(n7375) );
  NAND2_X1 U9036 ( .A1(n7376), .A2(n7375), .ZN(n7378) );
  INV_X1 U9037 ( .A(n7377), .ZN(n7380) );
  INV_X1 U9038 ( .A(n7378), .ZN(n7379) );
  NAND2_X1 U9039 ( .A1(n7380), .A2(n7379), .ZN(n7430) );
  NAND2_X1 U9040 ( .A1(n7428), .A2(n7430), .ZN(n7381) );
  XNOR2_X1 U9041 ( .A(n7429), .B(n7381), .ZN(n7388) );
  INV_X1 U9042 ( .A(n7382), .ZN(n7404) );
  NOR2_X1 U9043 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7383), .ZN(n9851) );
  AOI21_X1 U9044 ( .B1(n8669), .B2(n8995), .A(n9851), .ZN(n7385) );
  NAND2_X1 U9045 ( .A1(n9707), .A2(n8994), .ZN(n7384) );
  OAI211_X1 U9046 ( .C1(n9722), .C2(n7404), .A(n7385), .B(n7384), .ZN(n7386)
         );
  AOI21_X1 U9047 ( .B1(n7408), .B2(n8638), .A(n7386), .ZN(n7387) );
  OAI21_X1 U9048 ( .B1(n7388), .B2(n8683), .A(n7387), .ZN(P1_U3215) );
  AOI22_X1 U9049 ( .A1(n7390), .A2(n7178), .B1(n9693), .B2(n7389), .ZN(n7391)
         );
  OAI211_X1 U9050 ( .C1(n10006), .C2(n7393), .A(n7392), .B(n7391), .ZN(n7395)
         );
  NAND2_X1 U9051 ( .A1(n7395), .A2(n10048), .ZN(n7394) );
  OAI21_X1 U9052 ( .B1(n10048), .B2(n6358), .A(n7394), .ZN(P2_U3530) );
  INV_X1 U9053 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n7397) );
  NAND2_X1 U9054 ( .A1(n7395), .A2(n4314), .ZN(n7396) );
  OAI21_X1 U9055 ( .B1(n4314), .B2(n7397), .A(n7396), .ZN(P2_U3481) );
  AOI21_X1 U9056 ( .B1(n7398), .B2(n8913), .A(n9732), .ZN(n7402) );
  OAI22_X1 U9057 ( .A1(n7399), .A2(n9889), .B1(n7538), .B2(n9887), .ZN(n7400)
         );
  AOI21_X1 U9058 ( .B1(n7402), .B2(n7401), .A(n7400), .ZN(n9682) );
  XOR2_X1 U9059 ( .A(n8913), .B(n7403), .Z(n9684) );
  INV_X1 U9060 ( .A(n9684), .ZN(n9687) );
  NAND2_X1 U9061 ( .A1(n9687), .A2(n9277), .ZN(n7410) );
  INV_X1 U9062 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7405) );
  OAI22_X1 U9063 ( .A1(n9918), .A2(n7405), .B1(n7404), .B2(n9272), .ZN(n7407)
         );
  OAI211_X1 U9064 ( .C1(n9876), .C2(n9683), .A(n9739), .B(n9877), .ZN(n9681)
         );
  NOR2_X1 U9065 ( .A1(n9681), .A2(n9059), .ZN(n7406) );
  AOI211_X1 U9066 ( .C1(n9737), .C2(n7408), .A(n7407), .B(n7406), .ZN(n7409)
         );
  OAI211_X1 U9067 ( .C1(n9938), .C2(n9682), .A(n7410), .B(n7409), .ZN(P1_U3281) );
  INV_X1 U9068 ( .A(n7411), .ZN(n7415) );
  AOI21_X1 U9069 ( .B1(P1_DATAO_REG_23__SCAN_IN), .B2(n8588), .A(n8067), .ZN(
        n7412) );
  OAI21_X1 U9070 ( .B1(n7415), .B2(n6195), .A(n7412), .ZN(P2_U3335) );
  NAND2_X1 U9071 ( .A1(n7413), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8982) );
  NAND2_X1 U9072 ( .A1(n9428), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n7414) );
  OAI211_X1 U9073 ( .C1(n7415), .C2(n9420), .A(n8982), .B(n7414), .ZN(P1_U3330) );
  INV_X1 U9074 ( .A(n8550), .ZN(n7458) );
  INV_X1 U9075 ( .A(n7448), .ZN(n7418) );
  OR2_X1 U9076 ( .A1(n8550), .A2(n7469), .ZN(n7933) );
  NAND2_X1 U9077 ( .A1(n8550), .A2(n7469), .ZN(n7932) );
  NAND2_X1 U9078 ( .A1(n7418), .A2(n4313), .ZN(n7447) );
  OAI21_X1 U9079 ( .B1(n7458), .B2(n7469), .A(n7447), .ZN(n7489) );
  OR2_X1 U9080 ( .A1(n8544), .A2(n7570), .ZN(n7938) );
  NAND2_X1 U9081 ( .A1(n8544), .A2(n7570), .ZN(n7939) );
  NAND2_X1 U9082 ( .A1(n7938), .A2(n7939), .ZN(n7936) );
  XNOR2_X1 U9083 ( .A(n7489), .B(n7936), .ZN(n8548) );
  INV_X1 U9084 ( .A(n7454), .ZN(n7419) );
  INV_X1 U9085 ( .A(n8544), .ZN(n7421) );
  AOI21_X1 U9086 ( .B1(n8544), .B2(n7419), .A(n7492), .ZN(n8545) );
  AOI22_X1 U9087 ( .A1(n8463), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n7466), .B2(
        n8452), .ZN(n7420) );
  OAI21_X1 U9088 ( .B1(n7421), .B2(n8455), .A(n7420), .ZN(n7426) );
  INV_X1 U9089 ( .A(n7936), .ZN(n8023) );
  XNOR2_X1 U9090 ( .A(n7496), .B(n8023), .ZN(n7424) );
  INV_X1 U9091 ( .A(n7789), .ZN(n8442) );
  AOI222_X1 U9092 ( .A1(n8411), .A2(n7424), .B1(n8072), .B2(n8441), .C1(n8442), 
        .C2(n8440), .ZN(n8547) );
  NOR2_X1 U9093 ( .A1(n8547), .A2(n8463), .ZN(n7425) );
  AOI211_X1 U9094 ( .C1(n8545), .C2(n8461), .A(n7426), .B(n7425), .ZN(n7427)
         );
  OAI21_X1 U9095 ( .B1(n8407), .B2(n8548), .A(n7427), .ZN(P2_U3282) );
  INV_X1 U9096 ( .A(n9738), .ZN(n9762) );
  NAND2_X1 U9097 ( .A1(n9738), .A2(n6865), .ZN(n7432) );
  NAND2_X1 U9098 ( .A1(n8994), .A2(n7146), .ZN(n7431) );
  NAND2_X1 U9099 ( .A1(n7432), .A2(n7431), .ZN(n7433) );
  XNOR2_X1 U9100 ( .A(n7433), .B(n7673), .ZN(n7526) );
  AND2_X1 U9101 ( .A1(n8994), .A2(n7733), .ZN(n7434) );
  AOI21_X1 U9102 ( .B1(n9738), .B2(n7666), .A(n7434), .ZN(n7527) );
  XNOR2_X1 U9103 ( .A(n7526), .B(n7527), .ZN(n7436) );
  AOI21_X1 U9104 ( .B1(n7435), .B2(n7436), .A(n8683), .ZN(n7438) );
  INV_X1 U9105 ( .A(n7436), .ZN(n7437) );
  NAND2_X1 U9106 ( .A1(n7438), .A2(n7531), .ZN(n7443) );
  AOI21_X1 U9107 ( .B1(n9707), .B2(n9728), .A(n7439), .ZN(n7440) );
  OAI21_X1 U9108 ( .B1(n9888), .B2(n9709), .A(n7440), .ZN(n7441) );
  AOI21_X1 U9109 ( .B1(n9736), .B2(n8692), .A(n7441), .ZN(n7442) );
  OAI211_X1 U9110 ( .C1(n9762), .C2(n8695), .A(n7443), .B(n7442), .ZN(P1_U3234) );
  OAI21_X1 U9111 ( .B1(n8022), .B2(n7445), .A(n7444), .ZN(n7453) );
  OAI22_X1 U9112 ( .A1(n7446), .A2(n8326), .B1(n7570), .B2(n8324), .ZN(n7452)
         );
  NAND2_X1 U9113 ( .A1(n7448), .A2(n8022), .ZN(n7449) );
  NAND2_X1 U9114 ( .A1(n7447), .A2(n7449), .ZN(n8554) );
  NOR2_X1 U9115 ( .A1(n8554), .A2(n7450), .ZN(n7451) );
  AOI211_X1 U9116 ( .C1(n8411), .C2(n7453), .A(n7452), .B(n7451), .ZN(n8553)
         );
  AOI21_X1 U9117 ( .B1(n8550), .B2(n7455), .A(n7454), .ZN(n8551) );
  AOI22_X1 U9118 ( .A1(n8463), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n7456), .B2(
        n8452), .ZN(n7457) );
  OAI21_X1 U9119 ( .B1(n7458), .B2(n8455), .A(n7457), .ZN(n7460) );
  NOR2_X1 U9120 ( .A1(n8554), .A2(n8458), .ZN(n7459) );
  AOI211_X1 U9121 ( .C1(n8551), .C2(n8461), .A(n7460), .B(n7459), .ZN(n7461)
         );
  OAI21_X1 U9122 ( .B1(n8553), .B2(n8463), .A(n7461), .ZN(P2_U3283) );
  INV_X1 U9123 ( .A(n7462), .ZN(n7463) );
  AOI21_X1 U9124 ( .B1(n7465), .B2(n7464), .A(n7463), .ZN(n7473) );
  INV_X1 U9125 ( .A(n7466), .ZN(n7468) );
  OAI21_X1 U9126 ( .B1(n7825), .B2(n7468), .A(n7467), .ZN(n7471) );
  OAI22_X1 U9127 ( .A1(n7789), .A2(n7826), .B1(n7827), .B2(n7469), .ZN(n7470)
         );
  AOI211_X1 U9128 ( .C1(n7830), .C2(n8544), .A(n7471), .B(n7470), .ZN(n7472)
         );
  OAI21_X1 U9129 ( .B1(n7473), .B2(n4570), .A(n7472), .ZN(P2_U3217) );
  INV_X1 U9130 ( .A(n7474), .ZN(n7502) );
  AOI22_X1 U9131 ( .A1(n7475), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_24__SCAN_IN), .B2(n8583), .ZN(n7476) );
  OAI21_X1 U9132 ( .B1(n7502), .B2(n6195), .A(n7476), .ZN(P2_U3334) );
  XNOR2_X1 U9133 ( .A(n7477), .B(n8914), .ZN(n7478) );
  AOI222_X1 U9134 ( .A1(n9892), .A2(n7478), .B1(n8993), .B2(n9925), .C1(n8994), 
        .C2(n9730), .ZN(n9757) );
  OAI21_X1 U9135 ( .B1(n7480), .B2(n8914), .A(n7479), .ZN(n7481) );
  INV_X1 U9136 ( .A(n7481), .ZN(n9760) );
  NAND2_X1 U9137 ( .A1(n9760), .A2(n9277), .ZN(n7488) );
  INV_X1 U9138 ( .A(n7540), .ZN(n9758) );
  INV_X1 U9139 ( .A(n9740), .ZN(n7483) );
  INV_X1 U9140 ( .A(n7516), .ZN(n7482) );
  OAI211_X1 U9141 ( .C1(n9758), .C2(n7483), .A(n7482), .B(n9877), .ZN(n9756)
         );
  INV_X1 U9142 ( .A(n9756), .ZN(n7486) );
  AOI22_X1 U9143 ( .A1(n9938), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n7535), .B2(
        n9896), .ZN(n7484) );
  OAI21_X1 U9144 ( .B1(n9758), .B2(n9899), .A(n7484), .ZN(n7485) );
  AOI21_X1 U9145 ( .B1(n7486), .B2(n9881), .A(n7485), .ZN(n7487) );
  OAI211_X1 U9146 ( .C1(n9938), .C2(n9757), .A(n7488), .B(n7487), .ZN(P1_U3279) );
  OR2_X1 U9147 ( .A1(n8539), .A2(n7789), .ZN(n7945) );
  NAND2_X1 U9148 ( .A1(n8539), .A2(n7789), .ZN(n7944) );
  NAND2_X1 U9149 ( .A1(n7490), .A2(n8025), .ZN(n8209) );
  OAI21_X1 U9150 ( .B1(n7490), .B2(n8025), .A(n8209), .ZN(n7491) );
  INV_X1 U9151 ( .A(n7491), .ZN(n8543) );
  INV_X1 U9152 ( .A(n7492), .ZN(n7493) );
  INV_X1 U9153 ( .A(n8539), .ZN(n7495) );
  AOI21_X1 U9154 ( .B1(n8539), .B2(n7493), .A(n8448), .ZN(n8540) );
  AOI22_X1 U9155 ( .A1(n8463), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n7567), .B2(
        n8452), .ZN(n7494) );
  OAI21_X1 U9156 ( .B1(n7495), .B2(n8455), .A(n7494), .ZN(n7499) );
  XNOR2_X1 U9157 ( .A(n8039), .B(n8025), .ZN(n7497) );
  AOI222_X1 U9158 ( .A1(n8411), .A2(n7497), .B1(n8071), .B2(n8441), .C1(n8415), 
        .C2(n8440), .ZN(n8542) );
  NOR2_X1 U9159 ( .A1(n8542), .A2(n8463), .ZN(n7498) );
  AOI211_X1 U9160 ( .C1(n8540), .C2(n8461), .A(n7499), .B(n7498), .ZN(n7500)
         );
  OAI21_X1 U9161 ( .B1(n8543), .B2(n8407), .A(n7500), .ZN(P2_U3281) );
  INV_X1 U9162 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7501) );
  OAI222_X1 U9163 ( .A1(n7503), .A2(P1_U3084), .B1(n9420), .B2(n7502), .C1(
        n7501), .C2(n7729), .ZN(P1_U3329) );
  INV_X1 U9164 ( .A(n6039), .ZN(n7544) );
  AOI22_X1 U9165 ( .A1(n7504), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_25__SCAN_IN), .B2(n8583), .ZN(n7505) );
  OAI21_X1 U9166 ( .B1(n7544), .B2(n6195), .A(n7505), .ZN(P2_U3333) );
  INV_X1 U9167 ( .A(n7508), .ZN(n8917) );
  XNOR2_X1 U9168 ( .A(n7506), .B(n8917), .ZN(n9753) );
  INV_X1 U9169 ( .A(n9946), .ZN(n9735) );
  NAND2_X1 U9170 ( .A1(n7507), .A2(n8729), .ZN(n7509) );
  NAND2_X1 U9171 ( .A1(n7509), .A2(n7508), .ZN(n7511) );
  NAND2_X1 U9172 ( .A1(n7511), .A2(n7510), .ZN(n7512) );
  NAND2_X1 U9173 ( .A1(n7512), .A2(n9892), .ZN(n7514) );
  AOI22_X1 U9174 ( .A1(n9730), .A2(n9728), .B1(n8992), .B2(n9925), .ZN(n7513)
         );
  NAND2_X1 U9175 ( .A1(n7514), .A2(n7513), .ZN(n7515) );
  AOI21_X1 U9176 ( .B1(n9753), .B2(n9735), .A(n7515), .ZN(n9755) );
  INV_X1 U9177 ( .A(n9267), .ZN(n9882) );
  OAI21_X1 U9178 ( .B1(n7516), .B2(n9751), .A(n9877), .ZN(n7517) );
  OR2_X1 U9179 ( .A1(n7517), .A2(n7581), .ZN(n9750) );
  AOI22_X1 U9180 ( .A1(n9938), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n7555), .B2(
        n9896), .ZN(n7519) );
  NAND2_X1 U9181 ( .A1(n7561), .A2(n9737), .ZN(n7518) );
  OAI211_X1 U9182 ( .C1(n9750), .C2(n9059), .A(n7519), .B(n7518), .ZN(n7520)
         );
  AOI21_X1 U9183 ( .B1(n9753), .B2(n9882), .A(n7520), .ZN(n7521) );
  OAI21_X1 U9184 ( .B1(n9755), .B2(n9938), .A(n7521), .ZN(P1_U3278) );
  NAND2_X1 U9185 ( .A1(n7540), .A2(n6865), .ZN(n7523) );
  NAND2_X1 U9186 ( .A1(n9728), .A2(n7666), .ZN(n7522) );
  NAND2_X1 U9187 ( .A1(n7523), .A2(n7522), .ZN(n7524) );
  XNOR2_X1 U9188 ( .A(n7524), .B(n7673), .ZN(n7547) );
  AND2_X1 U9189 ( .A1(n9728), .A2(n7733), .ZN(n7525) );
  AOI21_X1 U9190 ( .B1(n7540), .B2(n7666), .A(n7525), .ZN(n7546) );
  XNOR2_X1 U9191 ( .A(n7547), .B(n7546), .ZN(n7534) );
  INV_X1 U9192 ( .A(n7526), .ZN(n7529) );
  INV_X1 U9193 ( .A(n7527), .ZN(n7528) );
  NAND2_X1 U9194 ( .A1(n7529), .A2(n7528), .ZN(n7530) );
  INV_X1 U9195 ( .A(n7549), .ZN(n7533) );
  AOI21_X1 U9196 ( .B1(n7534), .B2(n7532), .A(n7533), .ZN(n7542) );
  NAND2_X1 U9197 ( .A1(n8692), .A2(n7535), .ZN(n7537) );
  AOI22_X1 U9198 ( .A1(n9707), .A2(n8993), .B1(P1_REG3_REG_12__SCAN_IN), .B2(
        P1_U3084), .ZN(n7536) );
  OAI211_X1 U9199 ( .C1(n7538), .C2(n9709), .A(n7537), .B(n7536), .ZN(n7539)
         );
  AOI21_X1 U9200 ( .B1(n7540), .B2(n8638), .A(n7539), .ZN(n7541) );
  OAI21_X1 U9201 ( .B1(n7542), .B2(n8683), .A(n7541), .ZN(P1_U3222) );
  OAI222_X1 U9202 ( .A1(P1_U3084), .A2(n7545), .B1(n9420), .B2(n7544), .C1(
        n7543), .C2(n7729), .ZN(P1_U3328) );
  NAND2_X1 U9203 ( .A1(n7547), .A2(n7546), .ZN(n7548) );
  NAND2_X1 U9204 ( .A1(n7549), .A2(n7548), .ZN(n7588) );
  NAND2_X1 U9205 ( .A1(n7561), .A2(n6865), .ZN(n7551) );
  NAND2_X1 U9206 ( .A1(n8993), .A2(n7146), .ZN(n7550) );
  NAND2_X1 U9207 ( .A1(n7551), .A2(n7550), .ZN(n7552) );
  XNOR2_X1 U9208 ( .A(n7552), .B(n7673), .ZN(n7589) );
  AND2_X1 U9209 ( .A1(n8993), .A2(n7733), .ZN(n7553) );
  AOI21_X1 U9210 ( .B1(n7561), .B2(n7666), .A(n7553), .ZN(n7590) );
  XNOR2_X1 U9211 ( .A(n7589), .B(n7590), .ZN(n7554) );
  XNOR2_X1 U9212 ( .A(n7588), .B(n7554), .ZN(n7563) );
  NAND2_X1 U9213 ( .A1(n8692), .A2(n7555), .ZN(n7558) );
  AOI21_X1 U9214 ( .B1(n9707), .B2(n8992), .A(n7556), .ZN(n7557) );
  OAI211_X1 U9215 ( .C1(n7559), .C2(n9709), .A(n7558), .B(n7557), .ZN(n7560)
         );
  AOI21_X1 U9216 ( .B1(n7561), .B2(n8638), .A(n7560), .ZN(n7562) );
  OAI21_X1 U9217 ( .B1(n7563), .B2(n8683), .A(n7562), .ZN(P1_U3232) );
  AOI21_X1 U9218 ( .B1(n7566), .B2(n7565), .A(n7564), .ZN(n7574) );
  INV_X1 U9219 ( .A(n7567), .ZN(n7569) );
  OAI21_X1 U9220 ( .B1(n7825), .B2(n7569), .A(n7568), .ZN(n7572) );
  INV_X1 U9221 ( .A(n8415), .ZN(n7947) );
  OAI22_X1 U9222 ( .A1(n7947), .A2(n7826), .B1(n7827), .B2(n7570), .ZN(n7571)
         );
  AOI211_X1 U9223 ( .C1(n8539), .C2(n7830), .A(n7572), .B(n7571), .ZN(n7573)
         );
  OAI21_X1 U9224 ( .B1(n7574), .B2(n4570), .A(n7573), .ZN(P2_U3243) );
  AOI21_X1 U9225 ( .B1(n7575), .B2(n8918), .A(n9732), .ZN(n7579) );
  OAI22_X1 U9226 ( .A1(n9245), .A2(n9887), .B1(n7576), .B2(n9889), .ZN(n7577)
         );
  AOI21_X1 U9227 ( .B1(n7579), .B2(n7578), .A(n7577), .ZN(n9746) );
  XOR2_X1 U9228 ( .A(n8918), .B(n7580), .Z(n9749) );
  NAND2_X1 U9229 ( .A1(n9749), .A2(n9277), .ZN(n7586) );
  OAI211_X1 U9230 ( .C1(n7581), .C2(n9747), .A(n9877), .B(n4336), .ZN(n9745)
         );
  INV_X1 U9231 ( .A(n9745), .ZN(n7584) );
  AOI22_X1 U9232 ( .A1(n9938), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n8595), .B2(
        n9896), .ZN(n7582) );
  OAI21_X1 U9233 ( .B1(n9747), .B2(n9899), .A(n7582), .ZN(n7583) );
  AOI21_X1 U9234 ( .B1(n7584), .B2(n9881), .A(n7583), .ZN(n7585) );
  OAI211_X1 U9235 ( .C1(n9938), .C2(n9746), .A(n7586), .B(n7585), .ZN(P1_U3277) );
  AND2_X1 U9236 ( .A1(n7589), .A2(n7590), .ZN(n7587) );
  INV_X1 U9237 ( .A(n7589), .ZN(n7592) );
  INV_X1 U9238 ( .A(n7590), .ZN(n7591) );
  NOR2_X2 U9239 ( .A1(n7593), .A2(n4927), .ZN(n7599) );
  NAND2_X1 U9240 ( .A1(n8719), .A2(n6865), .ZN(n7595) );
  NAND2_X1 U9241 ( .A1(n8992), .A2(n7666), .ZN(n7594) );
  NAND2_X1 U9242 ( .A1(n7595), .A2(n7594), .ZN(n7596) );
  XNOR2_X1 U9243 ( .A(n7596), .B(n7673), .ZN(n7600) );
  NAND2_X1 U9244 ( .A1(n8719), .A2(n7146), .ZN(n7598) );
  NAND2_X1 U9245 ( .A1(n8992), .A2(n7733), .ZN(n7597) );
  NAND2_X1 U9246 ( .A1(n7598), .A2(n7597), .ZN(n8594) );
  INV_X1 U9247 ( .A(n7600), .ZN(n7601) );
  NAND2_X1 U9248 ( .A1(n9712), .A2(n6865), .ZN(n7603) );
  NAND2_X1 U9249 ( .A1(n8991), .A2(n7666), .ZN(n7602) );
  NAND2_X1 U9250 ( .A1(n7603), .A2(n7602), .ZN(n7604) );
  XNOR2_X1 U9251 ( .A(n7604), .B(n7673), .ZN(n7607) );
  NAND2_X1 U9252 ( .A1(n9712), .A2(n7666), .ZN(n7606) );
  NAND2_X1 U9253 ( .A1(n8991), .A2(n7733), .ZN(n7605) );
  NAND2_X1 U9254 ( .A1(n7606), .A2(n7605), .ZN(n9715) );
  NAND2_X1 U9255 ( .A1(n9714), .A2(n9715), .ZN(n7609) );
  INV_X1 U9256 ( .A(n7607), .ZN(n7608) );
  NAND2_X1 U9257 ( .A1(n9247), .A2(n6865), .ZN(n7611) );
  NAND2_X1 U9258 ( .A1(n9706), .A2(n7146), .ZN(n7610) );
  NAND2_X1 U9259 ( .A1(n7611), .A2(n7610), .ZN(n7612) );
  XNOR2_X1 U9260 ( .A(n7612), .B(n7673), .ZN(n7615) );
  AND2_X1 U9261 ( .A1(n9706), .A2(n7733), .ZN(n7613) );
  AOI21_X1 U9262 ( .B1(n9247), .B2(n7666), .A(n7613), .ZN(n7614) );
  XNOR2_X1 U9263 ( .A(n7615), .B(n7614), .ZN(n8634) );
  NAND2_X1 U9264 ( .A1(n7615), .A2(n7614), .ZN(n7616) );
  OAI21_X1 U9265 ( .B1(n8633), .B2(n8634), .A(n7616), .ZN(n8641) );
  NAND2_X1 U9266 ( .A1(n9351), .A2(n6865), .ZN(n7618) );
  NAND2_X1 U9267 ( .A1(n9213), .A2(n7666), .ZN(n7617) );
  NAND2_X1 U9268 ( .A1(n7618), .A2(n7617), .ZN(n7619) );
  XNOR2_X1 U9269 ( .A(n7619), .B(n7736), .ZN(n7621) );
  AND2_X1 U9270 ( .A1(n9213), .A2(n7733), .ZN(n7620) );
  AOI21_X1 U9271 ( .B1(n9351), .B2(n7666), .A(n7620), .ZN(n7622) );
  XNOR2_X1 U9272 ( .A(n7621), .B(n7622), .ZN(n8642) );
  NAND2_X1 U9273 ( .A1(n8641), .A2(n8642), .ZN(n7625) );
  INV_X1 U9274 ( .A(n7621), .ZN(n7623) );
  NAND2_X1 U9275 ( .A1(n7623), .A2(n7622), .ZN(n7624) );
  NAND2_X1 U9276 ( .A1(n9219), .A2(n6865), .ZN(n7627) );
  NAND2_X1 U9277 ( .A1(n8990), .A2(n7666), .ZN(n7626) );
  NAND2_X1 U9278 ( .A1(n7627), .A2(n7626), .ZN(n7628) );
  XNOR2_X1 U9279 ( .A(n7628), .B(n7673), .ZN(n7632) );
  NAND2_X1 U9280 ( .A1(n9219), .A2(n7666), .ZN(n7630) );
  NAND2_X1 U9281 ( .A1(n8990), .A2(n7733), .ZN(n7629) );
  NAND2_X1 U9282 ( .A1(n7630), .A2(n7629), .ZN(n8678) );
  INV_X1 U9283 ( .A(n7632), .ZN(n7633) );
  NAND2_X1 U9284 ( .A1(n9341), .A2(n6865), .ZN(n7636) );
  NAND2_X1 U9285 ( .A1(n9212), .A2(n7146), .ZN(n7635) );
  NAND2_X1 U9286 ( .A1(n7636), .A2(n7635), .ZN(n7637) );
  XNOR2_X1 U9287 ( .A(n7637), .B(n7673), .ZN(n7640) );
  AND2_X1 U9288 ( .A1(n9212), .A2(n7733), .ZN(n7638) );
  AOI21_X1 U9289 ( .B1(n9341), .B2(n7666), .A(n7638), .ZN(n7639) );
  XNOR2_X1 U9290 ( .A(n7640), .B(n7639), .ZN(n8612) );
  NAND2_X1 U9291 ( .A1(n7640), .A2(n7639), .ZN(n7641) );
  NAND2_X1 U9292 ( .A1(n9183), .A2(n6865), .ZN(n7643) );
  NAND2_X1 U9293 ( .A1(n8989), .A2(n7146), .ZN(n7642) );
  NAND2_X1 U9294 ( .A1(n7643), .A2(n7642), .ZN(n7644) );
  XNOR2_X1 U9295 ( .A(n7644), .B(n7736), .ZN(n7646) );
  AND2_X1 U9296 ( .A1(n8989), .A2(n7733), .ZN(n7645) );
  AOI21_X1 U9297 ( .B1(n9183), .B2(n7666), .A(n7645), .ZN(n7647) );
  XNOR2_X1 U9298 ( .A(n7646), .B(n7647), .ZN(n8658) );
  INV_X1 U9299 ( .A(n7646), .ZN(n7648) );
  NAND2_X1 U9300 ( .A1(n9328), .A2(n6865), .ZN(n7650) );
  NAND2_X1 U9301 ( .A1(n8988), .A2(n7666), .ZN(n7649) );
  NAND2_X1 U9302 ( .A1(n7650), .A2(n7649), .ZN(n7651) );
  XNOR2_X1 U9303 ( .A(n7651), .B(n7736), .ZN(n7653) );
  AND2_X1 U9304 ( .A1(n8988), .A2(n7733), .ZN(n7652) );
  AOI21_X1 U9305 ( .B1(n9328), .B2(n7666), .A(n7652), .ZN(n7654) );
  XNOR2_X1 U9306 ( .A(n7653), .B(n7654), .ZN(n8619) );
  NAND2_X1 U9307 ( .A1(n8618), .A2(n8619), .ZN(n7657) );
  INV_X1 U9308 ( .A(n7653), .ZN(n7655) );
  NAND2_X1 U9309 ( .A1(n7655), .A2(n7654), .ZN(n7656) );
  AND2_X1 U9310 ( .A1(n8987), .A2(n7733), .ZN(n7658) );
  AOI21_X1 U9311 ( .B1(n9152), .B2(n7666), .A(n7658), .ZN(n7662) );
  NAND2_X1 U9312 ( .A1(n9152), .A2(n6865), .ZN(n7660) );
  NAND2_X1 U9313 ( .A1(n8987), .A2(n7146), .ZN(n7659) );
  NAND2_X1 U9314 ( .A1(n7660), .A2(n7659), .ZN(n7661) );
  NAND2_X1 U9315 ( .A1(n9319), .A2(n6865), .ZN(n7664) );
  NAND2_X1 U9316 ( .A1(n9118), .A2(n7666), .ZN(n7663) );
  NAND2_X1 U9317 ( .A1(n7664), .A2(n7663), .ZN(n7665) );
  XNOR2_X1 U9318 ( .A(n7665), .B(n7673), .ZN(n7669) );
  NAND2_X1 U9319 ( .A1(n9319), .A2(n7666), .ZN(n7668) );
  NAND2_X1 U9320 ( .A1(n9118), .A2(n7733), .ZN(n7667) );
  NAND2_X1 U9321 ( .A1(n7668), .A2(n7667), .ZN(n8605) );
  INV_X1 U9322 ( .A(n7669), .ZN(n7670) );
  NAND2_X1 U9323 ( .A1(n9120), .A2(n6865), .ZN(n7672) );
  NAND2_X1 U9324 ( .A1(n8986), .A2(n7146), .ZN(n7671) );
  NAND2_X1 U9325 ( .A1(n7672), .A2(n7671), .ZN(n7674) );
  XNOR2_X1 U9326 ( .A(n7674), .B(n7673), .ZN(n7678) );
  AND2_X1 U9327 ( .A1(n8986), .A2(n7733), .ZN(n7675) );
  AOI21_X1 U9328 ( .B1(n9120), .B2(n7146), .A(n7675), .ZN(n7677) );
  XNOR2_X1 U9329 ( .A(n7678), .B(n7677), .ZN(n8651) );
  NAND2_X1 U9330 ( .A1(n7678), .A2(n7677), .ZN(n7679) );
  NAND2_X1 U9331 ( .A1(n8649), .A2(n7679), .ZN(n8626) );
  NAND2_X1 U9332 ( .A1(n9310), .A2(n6865), .ZN(n7681) );
  NAND2_X1 U9333 ( .A1(n9117), .A2(n7146), .ZN(n7680) );
  NAND2_X1 U9334 ( .A1(n7681), .A2(n7680), .ZN(n7682) );
  XNOR2_X1 U9335 ( .A(n7682), .B(n7736), .ZN(n7684) );
  AND2_X1 U9336 ( .A1(n9117), .A2(n7733), .ZN(n7683) );
  AOI21_X1 U9337 ( .B1(n9310), .B2(n7146), .A(n7683), .ZN(n7685) );
  XNOR2_X1 U9338 ( .A(n7684), .B(n7685), .ZN(n8627) );
  INV_X1 U9339 ( .A(n7684), .ZN(n7686) );
  NAND2_X1 U9340 ( .A1(n9092), .A2(n6865), .ZN(n7688) );
  NAND2_X1 U9341 ( .A1(n9080), .A2(n7666), .ZN(n7687) );
  NAND2_X1 U9342 ( .A1(n7688), .A2(n7687), .ZN(n7689) );
  XNOR2_X1 U9343 ( .A(n7689), .B(n7736), .ZN(n7693) );
  AND2_X1 U9344 ( .A1(n9080), .A2(n7733), .ZN(n7690) );
  AOI21_X1 U9345 ( .B1(n9092), .B2(n7146), .A(n7690), .ZN(n7691) );
  XNOR2_X1 U9346 ( .A(n7693), .B(n7691), .ZN(n8687) );
  INV_X1 U9347 ( .A(n7691), .ZN(n7692) );
  NAND2_X1 U9348 ( .A1(n9299), .A2(n6865), .ZN(n7695) );
  NAND2_X1 U9349 ( .A1(n8985), .A2(n7666), .ZN(n7694) );
  NAND2_X1 U9350 ( .A1(n7695), .A2(n7694), .ZN(n7696) );
  XNOR2_X1 U9351 ( .A(n7696), .B(n7736), .ZN(n7702) );
  INV_X1 U9352 ( .A(n7702), .ZN(n7700) );
  NAND2_X1 U9353 ( .A1(n9299), .A2(n7666), .ZN(n7698) );
  NAND2_X1 U9354 ( .A1(n8985), .A2(n7733), .ZN(n7697) );
  NAND2_X1 U9355 ( .A1(n7698), .A2(n7697), .ZN(n7701) );
  INV_X1 U9356 ( .A(n7701), .ZN(n7699) );
  NAND2_X1 U9357 ( .A1(n7700), .A2(n7699), .ZN(n7745) );
  INV_X1 U9358 ( .A(n7745), .ZN(n7703) );
  NOR2_X1 U9359 ( .A1(n7703), .A2(n7732), .ZN(n7704) );
  AOI22_X1 U9360 ( .A1(n9080), .A2(n8669), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3084), .ZN(n7706) );
  NAND2_X1 U9361 ( .A1(n9074), .A2(n8692), .ZN(n7705) );
  OAI211_X1 U9362 ( .C1(n7707), .C2(n8689), .A(n7706), .B(n7705), .ZN(n7708)
         );
  AOI21_X1 U9363 ( .B1(n9299), .B2(n8638), .A(n7708), .ZN(n7709) );
  OAI21_X1 U9364 ( .B1(n7710), .B2(n8683), .A(n7709), .ZN(P1_U3212) );
  AOI22_X1 U9365 ( .A1(n9428), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        P1_STATE_REG_SCAN_IN), .B2(n7726), .ZN(n7711) );
  OAI21_X1 U9366 ( .B1(n7712), .B2(n9420), .A(n7711), .ZN(P1_U3352) );
  INV_X1 U9367 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n7728) );
  NOR2_X1 U9368 ( .A1(n7713), .A2(n9969), .ZN(n7718) );
  INV_X1 U9369 ( .A(n7714), .ZN(n7717) );
  INV_X1 U9370 ( .A(n7715), .ZN(n7716) );
  OAI211_X1 U9371 ( .C1(n7718), .C2(n7717), .A(n9868), .B(n7716), .ZN(n7723)
         );
  OAI211_X1 U9372 ( .C1(n7721), .C2(n6321), .A(n9869), .B(n7720), .ZN(n7722)
         );
  OAI211_X1 U9373 ( .C1(P1_STATE_REG_SCAN_IN), .C2(n7724), .A(n7723), .B(n7722), .ZN(n7725) );
  AOI21_X1 U9374 ( .B1(n9860), .B2(n7726), .A(n7725), .ZN(n7727) );
  OAI21_X1 U9375 ( .B1(n9873), .B2(n7728), .A(n7727), .ZN(P1_U3242) );
  INV_X1 U9376 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7730) );
  OAI222_X1 U9377 ( .A1(n5503), .A2(P1_U3084), .B1(n9420), .B2(n7731), .C1(
        n7730), .C2(n7729), .ZN(P1_U3332) );
  NAND2_X1 U9378 ( .A1(n9060), .A2(n7666), .ZN(n7735) );
  NAND2_X1 U9379 ( .A1(n9079), .A2(n7733), .ZN(n7734) );
  NAND2_X1 U9380 ( .A1(n7735), .A2(n7734), .ZN(n7737) );
  XNOR2_X1 U9381 ( .A(n7737), .B(n7736), .ZN(n7739) );
  AOI22_X1 U9382 ( .A1(n9060), .A2(n6865), .B1(n7146), .B2(n9079), .ZN(n7738)
         );
  XNOR2_X1 U9383 ( .A(n7739), .B(n7738), .ZN(n7740) );
  INV_X1 U9384 ( .A(n7740), .ZN(n7746) );
  NAND3_X1 U9385 ( .A1(n7746), .A2(n9717), .A3(n7745), .ZN(n7750) );
  INV_X1 U9386 ( .A(n7742), .ZN(n9062) );
  AOI22_X1 U9387 ( .A1(n9062), .A2(n8692), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n7744) );
  NAND2_X1 U9388 ( .A1(n8984), .A2(n9707), .ZN(n7743) );
  OAI211_X1 U9389 ( .C1(n9087), .C2(n9709), .A(n7744), .B(n7743), .ZN(n7748)
         );
  NOR3_X1 U9390 ( .A1(n7746), .A2(n8683), .A3(n7745), .ZN(n7747) );
  AOI211_X1 U9391 ( .C1(n8638), .C2(n9060), .A(n7748), .B(n7747), .ZN(n7749)
         );
  XNOR2_X1 U9392 ( .A(n7751), .B(n7752), .ZN(n7757) );
  INV_X1 U9393 ( .A(n8328), .ZN(n7753) );
  OAI22_X1 U9394 ( .A1(n7825), .A2(n7753), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9502), .ZN(n7755) );
  INV_X1 U9395 ( .A(n8217), .ZN(n8323) );
  OAI22_X1 U9396 ( .A1(n8323), .A2(n7826), .B1(n7827), .B2(n8325), .ZN(n7754)
         );
  AOI211_X1 U9397 ( .C1(n8329), .C2(n7830), .A(n7755), .B(n7754), .ZN(n7756)
         );
  OAI21_X1 U9398 ( .B1(n7757), .B2(n4570), .A(n7756), .ZN(P2_U3218) );
  OAI21_X1 U9399 ( .B1(n7760), .B2(n7759), .A(n7758), .ZN(n7761) );
  NAND2_X1 U9400 ( .A1(n7761), .A2(n7835), .ZN(n7767) );
  INV_X1 U9401 ( .A(n7762), .ZN(n8387) );
  INV_X1 U9402 ( .A(n7763), .ZN(n7838) );
  AND2_X1 U9403 ( .A1(n8416), .A2(n8441), .ZN(n7764) );
  AOI21_X1 U9404 ( .B1(n8358), .B2(n8440), .A(n7764), .ZN(n8382) );
  NAND2_X1 U9405 ( .A1(P2_U3152), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8179) );
  OAI21_X1 U9406 ( .B1(n7838), .B2(n8382), .A(n8179), .ZN(n7765) );
  AOI21_X1 U9407 ( .B1(n8387), .B2(n7840), .A(n7765), .ZN(n7766) );
  OAI211_X1 U9408 ( .C1(n8390), .C2(n7843), .A(n7767), .B(n7766), .ZN(P2_U3221) );
  XNOR2_X1 U9409 ( .A(n7768), .B(n7769), .ZN(n7774) );
  INV_X1 U9410 ( .A(n8353), .ZN(n7770) );
  OAI22_X1 U9411 ( .A1(n7825), .A2(n7770), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9468), .ZN(n7772) );
  INV_X1 U9412 ( .A(n8358), .ZN(n7957) );
  OAI22_X1 U9413 ( .A1(n7957), .A2(n7827), .B1(n7826), .B2(n8325), .ZN(n7771)
         );
  AOI211_X1 U9414 ( .C1(n8509), .C2(n7830), .A(n7772), .B(n7771), .ZN(n7773)
         );
  OAI21_X1 U9415 ( .B1(n7774), .B2(n4570), .A(n7773), .ZN(P2_U3225) );
  XNOR2_X1 U9416 ( .A(n7777), .B(n7776), .ZN(n7778) );
  XNOR2_X1 U9417 ( .A(n7775), .B(n7778), .ZN(n7783) );
  AOI22_X1 U9418 ( .A1(n8223), .A2(n8440), .B1(n8441), .B2(n8217), .ZN(n8292)
         );
  OAI22_X1 U9419 ( .A1(n8292), .A2(n7838), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7779), .ZN(n7780) );
  AOI21_X1 U9420 ( .B1(n8295), .B2(n7840), .A(n7780), .ZN(n7782) );
  NAND2_X1 U9421 ( .A1(n8488), .A2(n7830), .ZN(n7781) );
  OAI211_X1 U9422 ( .C1(n7783), .C2(n4570), .A(n7782), .B(n7781), .ZN(P2_U3227) );
  INV_X1 U9423 ( .A(n8534), .ZN(n8456) );
  INV_X1 U9424 ( .A(n7784), .ZN(n7788) );
  NOR3_X1 U9425 ( .A1(n7564), .A2(n7786), .A3(n7785), .ZN(n7787) );
  OAI21_X1 U9426 ( .B1(n7788), .B2(n7787), .A(n7835), .ZN(n7793) );
  OAI22_X1 U9427 ( .A1(n7789), .A2(n7827), .B1(n7826), .B2(n8210), .ZN(n7790)
         );
  AOI211_X1 U9428 ( .C1(n7840), .C2(n8453), .A(n7791), .B(n7790), .ZN(n7792)
         );
  OAI211_X1 U9429 ( .C1(n8456), .C2(n7843), .A(n7793), .B(n7792), .ZN(P2_U3228) );
  XNOR2_X1 U9430 ( .A(n7795), .B(n7794), .ZN(n7799) );
  OAI22_X1 U9431 ( .A1(n7825), .A2(n8427), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9500), .ZN(n7797) );
  INV_X1 U9432 ( .A(n8416), .ZN(n8212) );
  OAI22_X1 U9433 ( .A1(n7947), .A2(n7827), .B1(n7826), .B2(n8212), .ZN(n7796)
         );
  AOI211_X1 U9434 ( .C1(n8530), .C2(n7830), .A(n7797), .B(n7796), .ZN(n7798)
         );
  OAI21_X1 U9435 ( .B1(n7799), .B2(n4570), .A(n7798), .ZN(P2_U3230) );
  XNOR2_X1 U9436 ( .A(n7800), .B(n7801), .ZN(n7806) );
  OAI22_X1 U9437 ( .A1(n7825), .A2(n8313), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7802), .ZN(n7804) );
  INV_X1 U9438 ( .A(n8304), .ZN(n7967) );
  OAI22_X1 U9439 ( .A1(n8220), .A2(n7826), .B1(n7827), .B2(n7967), .ZN(n7803)
         );
  AOI211_X1 U9440 ( .C1(n8492), .C2(n7830), .A(n7804), .B(n7803), .ZN(n7805)
         );
  OAI21_X1 U9441 ( .B1(n7806), .B2(n4570), .A(n7805), .ZN(P2_U3231) );
  XNOR2_X1 U9442 ( .A(n7807), .B(n7808), .ZN(n7812) );
  OAI22_X1 U9443 ( .A1(n7825), .A2(n8368), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9616), .ZN(n7810) );
  INV_X1 U9444 ( .A(n8402), .ZN(n8213) );
  INV_X1 U9445 ( .A(n8373), .ZN(n8214) );
  OAI22_X1 U9446 ( .A1(n8213), .A2(n7827), .B1(n7826), .B2(n8214), .ZN(n7809)
         );
  AOI211_X1 U9447 ( .C1(n8514), .C2(n7830), .A(n7810), .B(n7809), .ZN(n7811)
         );
  OAI21_X1 U9448 ( .B1(n7812), .B2(n4570), .A(n7811), .ZN(P2_U3235) );
  OAI21_X1 U9449 ( .B1(n7815), .B2(n7814), .A(n7813), .ZN(n7816) );
  NAND2_X1 U9450 ( .A1(n7816), .A2(n7835), .ZN(n7822) );
  INV_X1 U9451 ( .A(n7817), .ZN(n8340) );
  AND2_X1 U9452 ( .A1(n8373), .A2(n8441), .ZN(n7818) );
  AOI21_X1 U9453 ( .B1(n8304), .B2(n8440), .A(n7818), .ZN(n8345) );
  OAI22_X1 U9454 ( .A1(n7838), .A2(n8345), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7819), .ZN(n7820) );
  AOI21_X1 U9455 ( .B1(n8340), .B2(n7840), .A(n7820), .ZN(n7821) );
  OAI211_X1 U9456 ( .C1(n4671), .C2(n7843), .A(n7822), .B(n7821), .ZN(P2_U3237) );
  XNOR2_X1 U9457 ( .A(n7824), .B(n7823), .ZN(n7832) );
  NAND2_X1 U9458 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8174) );
  OAI21_X1 U9459 ( .B1(n7825), .B2(n8396), .A(n8174), .ZN(n7829) );
  OAI22_X1 U9460 ( .A1(n8210), .A2(n7827), .B1(n7826), .B2(n8213), .ZN(n7828)
         );
  AOI211_X1 U9461 ( .C1(n8525), .C2(n7830), .A(n7829), .B(n7828), .ZN(n7831)
         );
  OAI21_X1 U9462 ( .B1(n7832), .B2(n4570), .A(n7831), .ZN(P2_U3240) );
  INV_X1 U9463 ( .A(n8483), .ZN(n8198) );
  OAI211_X1 U9464 ( .C1(n7833), .C2(n7836), .A(n7834), .B(n7835), .ZN(n7842)
         );
  AOI22_X1 U9465 ( .A1(n8224), .A2(n8440), .B1(n8441), .B2(n8305), .ZN(n8276)
         );
  OAI22_X1 U9466 ( .A1(n8276), .A2(n7838), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7837), .ZN(n7839) );
  AOI21_X1 U9467 ( .B1(n8281), .B2(n7840), .A(n7839), .ZN(n7841) );
  OAI211_X1 U9468 ( .C1(n8198), .C2(n7843), .A(n7842), .B(n7841), .ZN(P2_U3242) );
  NOR4_X1 U9469 ( .A1(n7845), .A2(n8326), .A3(n8202), .A4(n7844), .ZN(n8069)
         );
  OAI21_X1 U9470 ( .B1(n7846), .B2(n6124), .A(P2_B_REG_SCAN_IN), .ZN(n8068) );
  NAND2_X1 U9471 ( .A1(n7848), .A2(n7847), .ZN(n7852) );
  INV_X1 U9472 ( .A(n7849), .ZN(n7850) );
  NAND2_X1 U9473 ( .A1(n7850), .A2(n9514), .ZN(n7851) );
  MUX2_X1 U9474 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .S(n5462), .Z(n7853) );
  INV_X1 U9475 ( .A(SI_30_), .ZN(n9604) );
  XNOR2_X1 U9476 ( .A(n7853), .B(n9604), .ZN(n7866) );
  NAND2_X1 U9477 ( .A1(n7867), .A2(n7866), .ZN(n7856) );
  INV_X1 U9478 ( .A(n7853), .ZN(n7854) );
  NAND2_X1 U9479 ( .A1(n7854), .A2(n9604), .ZN(n7855) );
  NAND2_X1 U9480 ( .A1(n7856), .A2(n7855), .ZN(n7860) );
  MUX2_X1 U9481 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n5462), .Z(n7858) );
  INV_X1 U9482 ( .A(SI_31_), .ZN(n7857) );
  XNOR2_X1 U9483 ( .A(n7858), .B(n7857), .ZN(n7859) );
  NAND2_X1 U9484 ( .A1(n8794), .A2(n7981), .ZN(n7863) );
  NAND2_X1 U9485 ( .A1(n7861), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n7862) );
  INV_X1 U9486 ( .A(n8055), .ZN(n8203) );
  NOR2_X1 U9487 ( .A1(n9692), .A2(n8203), .ZN(n7992) );
  NOR2_X1 U9488 ( .A1(n8425), .A2(n8054), .ZN(n7865) );
  AOI222_X1 U9489 ( .A1(n4312), .A2(P2_REG1_REG_30__SCAN_IN), .B1(n7868), .B2(
        P2_REG0_REG_30__SCAN_IN), .C1(n4309), .C2(P2_REG2_REG_30__SCAN_IN), 
        .ZN(n8230) );
  INV_X1 U9490 ( .A(n8230), .ZN(n8070) );
  NOR2_X1 U9491 ( .A1(n9696), .A2(n8070), .ZN(n7989) );
  NOR2_X1 U9492 ( .A1(n7992), .A2(n7989), .ZN(n8056) );
  NOR2_X1 U9493 ( .A1(n8217), .A2(n7893), .ZN(n7969) );
  NAND2_X1 U9494 ( .A1(n8488), .A2(n8220), .ZN(n7970) );
  INV_X1 U9495 ( .A(n8291), .ZN(n8222) );
  NAND2_X1 U9496 ( .A1(n7871), .A2(n7869), .ZN(n7870) );
  NAND2_X1 U9497 ( .A1(n7873), .A2(n7893), .ZN(n7882) );
  INV_X1 U9498 ( .A(n7892), .ZN(n7880) );
  AND2_X1 U9499 ( .A1(n8005), .A2(n7874), .ZN(n7876) );
  OAI211_X1 U9500 ( .C1(n7876), .C2(n7875), .A(n7883), .B(n7887), .ZN(n7877)
         );
  NAND3_X1 U9501 ( .A1(n7877), .A2(n7893), .A3(n7884), .ZN(n7878) );
  NAND3_X1 U9502 ( .A1(n7880), .A2(n7879), .A3(n7878), .ZN(n7881) );
  NAND2_X1 U9503 ( .A1(n7883), .A2(n8005), .ZN(n7885) );
  NAND3_X1 U9504 ( .A1(n7886), .A2(n7885), .A3(n7884), .ZN(n7888) );
  AOI22_X1 U9505 ( .A1(n7892), .A2(n7891), .B1(n7890), .B2(n7889), .ZN(n7895)
         );
  INV_X1 U9506 ( .A(n7896), .ZN(n7894) );
  OAI21_X1 U9507 ( .B1(n7895), .B2(n7894), .A(n7966), .ZN(n7899) );
  MUX2_X1 U9508 ( .A(n7897), .B(n7896), .S(n7893), .Z(n7898) );
  INV_X1 U9509 ( .A(n7902), .ZN(n7903) );
  INV_X1 U9510 ( .A(n7904), .ZN(n7911) );
  INV_X1 U9511 ( .A(n7905), .ZN(n7906) );
  NOR2_X1 U9512 ( .A1(n7911), .A2(n7906), .ZN(n7907) );
  NAND2_X1 U9513 ( .A1(n7908), .A2(n7909), .ZN(n7925) );
  NAND2_X1 U9514 ( .A1(n7920), .A2(n7909), .ZN(n7910) );
  MUX2_X1 U9515 ( .A(n7911), .B(n7910), .S(n7893), .Z(n7913) );
  OR2_X1 U9516 ( .A1(n7913), .A2(n7912), .ZN(n7918) );
  INV_X1 U9517 ( .A(n7918), .ZN(n7924) );
  NAND3_X1 U9518 ( .A1(n7916), .A2(n4839), .A3(n7915), .ZN(n7919) );
  OAI211_X1 U9519 ( .C1(n7919), .C2(n7918), .A(n7917), .B(n7926), .ZN(n7922)
         );
  NAND2_X1 U9520 ( .A1(n7928), .A2(n7920), .ZN(n7921) );
  MUX2_X1 U9521 ( .A(n7922), .B(n7921), .S(n7966), .Z(n7923) );
  NAND2_X1 U9522 ( .A1(n7930), .A2(n7926), .ZN(n7927) );
  NAND2_X1 U9523 ( .A1(n7929), .A2(n7928), .ZN(n7931) );
  INV_X1 U9524 ( .A(n7932), .ZN(n7935) );
  INV_X1 U9525 ( .A(n7933), .ZN(n7934) );
  MUX2_X1 U9526 ( .A(n7935), .B(n7934), .S(n7893), .Z(n7937) );
  INV_X1 U9527 ( .A(n7938), .ZN(n7941) );
  INV_X1 U9528 ( .A(n7939), .ZN(n7940) );
  MUX2_X1 U9529 ( .A(n7941), .B(n7940), .S(n7893), .Z(n7942) );
  INV_X1 U9530 ( .A(n7944), .ZN(n7946) );
  INV_X1 U9531 ( .A(n7945), .ZN(n8037) );
  MUX2_X1 U9532 ( .A(n7946), .B(n8037), .S(n7893), .Z(n7949) );
  OR2_X1 U9533 ( .A1(n8534), .A2(n7947), .ZN(n8041) );
  AND2_X1 U9534 ( .A1(n8534), .A2(n7947), .ZN(n8040) );
  INV_X1 U9535 ( .A(n8040), .ZN(n7948) );
  NAND2_X1 U9536 ( .A1(n8041), .A2(n7948), .ZN(n8437) );
  INV_X1 U9537 ( .A(n8041), .ZN(n7950) );
  MUX2_X1 U9538 ( .A(n7950), .B(n8040), .S(n7893), .Z(n7951) );
  NAND2_X1 U9539 ( .A1(n8530), .A2(n8210), .ZN(n7952) );
  OR2_X1 U9540 ( .A1(n8525), .A2(n8212), .ZN(n8004) );
  INV_X1 U9541 ( .A(n8004), .ZN(n7956) );
  NAND2_X1 U9542 ( .A1(n8043), .A2(n7952), .ZN(n7954) );
  INV_X1 U9543 ( .A(n8042), .ZN(n7953) );
  MUX2_X1 U9544 ( .A(n7954), .B(n7953), .S(n7893), .Z(n7955) );
  OR2_X1 U9545 ( .A1(n8521), .A2(n8213), .ZN(n8003) );
  INV_X1 U9546 ( .A(n8003), .ZN(n7958) );
  NAND2_X1 U9547 ( .A1(n8521), .A2(n8213), .ZN(n8002) );
  NAND2_X1 U9548 ( .A1(n8514), .A2(n7957), .ZN(n8001) );
  OR2_X1 U9549 ( .A1(n8509), .A2(n8214), .ZN(n8000) );
  INV_X1 U9550 ( .A(n8000), .ZN(n7959) );
  AOI21_X1 U9551 ( .B1(n7961), .B2(n8001), .A(n7959), .ZN(n7960) );
  NAND2_X1 U9552 ( .A1(n8504), .A2(n8325), .ZN(n7999) );
  NAND2_X1 U9553 ( .A1(n8509), .A2(n8214), .ZN(n8045) );
  NAND2_X1 U9554 ( .A1(n7999), .A2(n8045), .ZN(n7962) );
  NAND3_X1 U9555 ( .A1(n7961), .A2(n8044), .A3(n8000), .ZN(n7964) );
  INV_X1 U9556 ( .A(n7962), .ZN(n7963) );
  AOI21_X1 U9557 ( .B1(n7964), .B2(n7963), .A(n4835), .ZN(n7965) );
  XOR2_X1 U9558 ( .A(n8304), .B(n8329), .Z(n8321) );
  INV_X1 U9559 ( .A(n8321), .ZN(n8333) );
  NOR2_X1 U9560 ( .A1(n8218), .A2(n8217), .ZN(n7998) );
  NOR2_X1 U9561 ( .A1(n8492), .A2(n8323), .ZN(n7997) );
  INV_X1 U9562 ( .A(n7997), .ZN(n8048) );
  OAI21_X1 U9563 ( .B1(n7967), .B2(n8329), .A(n8048), .ZN(n7968) );
  NAND2_X1 U9564 ( .A1(n7973), .A2(n8273), .ZN(n7972) );
  NAND2_X1 U9565 ( .A1(n8483), .A2(n8262), .ZN(n8049) );
  NAND2_X1 U9566 ( .A1(n8272), .A2(n7970), .ZN(n7971) );
  MUX2_X1 U9567 ( .A(n7972), .B(n7971), .S(n7893), .Z(n7975) );
  MUX2_X1 U9568 ( .A(n8049), .B(n7973), .S(n7893), .Z(n7974) );
  INV_X1 U9569 ( .A(n8261), .ZN(n8253) );
  OAI211_X1 U9570 ( .C1(n7976), .C2(n7975), .A(n7974), .B(n8253), .ZN(n7980)
         );
  NAND2_X1 U9571 ( .A1(n8471), .A2(n8263), .ZN(n7995) );
  NOR2_X1 U9572 ( .A1(n8476), .A2(n8246), .ZN(n8050) );
  NOR2_X1 U9573 ( .A1(n8051), .A2(n8050), .ZN(n7978) );
  NAND2_X1 U9574 ( .A1(n8476), .A2(n8246), .ZN(n7977) );
  MUX2_X1 U9575 ( .A(n7978), .B(n7977), .S(n7893), .Z(n7979) );
  NAND3_X1 U9576 ( .A1(n7980), .A2(n7995), .A3(n7979), .ZN(n7987) );
  NAND2_X1 U9577 ( .A1(n8578), .A2(n7981), .ZN(n7983) );
  NAND2_X1 U9578 ( .A1(n5715), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n7982) );
  NAND2_X1 U9579 ( .A1(n7983), .A2(n7982), .ZN(n8467) );
  INV_X1 U9580 ( .A(n8052), .ZN(n7984) );
  OAI211_X1 U9581 ( .C1(n7966), .C2(n8471), .A(n7984), .B(n7995), .ZN(n7985)
         );
  OAI21_X1 U9582 ( .B1(n7966), .B2(n4777), .A(n7985), .ZN(n7986) );
  AOI22_X1 U9583 ( .A1(n7987), .A2(n7986), .B1(n8052), .B2(n7893), .ZN(n7988)
         );
  OR2_X1 U9584 ( .A1(n8467), .A2(n8247), .ZN(n8053) );
  INV_X1 U9585 ( .A(n9696), .ZN(n8200) );
  NOR2_X1 U9586 ( .A1(n8200), .A2(n8230), .ZN(n8057) );
  INV_X1 U9587 ( .A(n8057), .ZN(n7991) );
  INV_X1 U9588 ( .A(n7989), .ZN(n7990) );
  NAND2_X1 U9589 ( .A1(n9692), .A2(n8203), .ZN(n8059) );
  NAND2_X1 U9590 ( .A1(n8059), .A2(n7991), .ZN(n7993) );
  INV_X1 U9591 ( .A(n7993), .ZN(n8032) );
  INV_X1 U9592 ( .A(n8272), .ZN(n8269) );
  INV_X1 U9593 ( .A(n8343), .ZN(n8338) );
  INV_X1 U9594 ( .A(n8356), .ZN(n8028) );
  NAND2_X1 U9595 ( .A1(n8004), .A2(n8043), .ZN(n8400) );
  INV_X1 U9596 ( .A(n8400), .ZN(n8393) );
  NAND4_X1 U9597 ( .A1(n8008), .A2(n8007), .A3(n8006), .A4(n8005), .ZN(n8012)
         );
  NOR4_X1 U9598 ( .A1(n8012), .A2(n8011), .A3(n8010), .A4(n8009), .ZN(n8015)
         );
  NAND4_X1 U9599 ( .A1(n8015), .A2(n8014), .A3(n4839), .A4(n8013), .ZN(n8018)
         );
  NOR4_X1 U9600 ( .A1(n8019), .A2(n8018), .A3(n8017), .A4(n7123), .ZN(n8020)
         );
  NAND4_X1 U9601 ( .A1(n8023), .A2(n8022), .A3(n8021), .A4(n8020), .ZN(n8024)
         );
  NOR4_X1 U9602 ( .A1(n8409), .A2(n8437), .A3(n8025), .A4(n8024), .ZN(n8026)
         );
  NAND3_X1 U9603 ( .A1(n8381), .A2(n8393), .A3(n8026), .ZN(n8027) );
  NOR4_X1 U9604 ( .A1(n8338), .A2(n8028), .A3(n4376), .A4(n8027), .ZN(n8029)
         );
  NAND4_X1 U9605 ( .A1(n8291), .A2(n8302), .A3(n8029), .A4(n8333), .ZN(n8030)
         );
  NOR4_X1 U9606 ( .A1(n8244), .A2(n8261), .A3(n8269), .A4(n8030), .ZN(n8031)
         );
  NAND4_X1 U9607 ( .A1(n8056), .A2(n8032), .A3(n8229), .A4(n8031), .ZN(n8033)
         );
  XNOR2_X1 U9608 ( .A(n8033), .B(n8283), .ZN(n8036) );
  INV_X1 U9609 ( .A(n6293), .ZN(n8035) );
  AOI22_X1 U9610 ( .A1(n8036), .A2(n8054), .B1(n8035), .B2(n8034), .ZN(n8065)
         );
  NAND2_X1 U9611 ( .A1(n8414), .A2(n8413), .ZN(n8412) );
  INV_X1 U9612 ( .A(n8045), .ZN(n8046) );
  NAND2_X1 U9613 ( .A1(n8301), .A2(n8048), .ZN(n8290) );
  AOI211_X1 U9614 ( .C1(n8058), .C2(n9696), .A(n8055), .B(n8054), .ZN(n8061)
         );
  OAI21_X1 U9615 ( .B1(n8058), .B2(n8057), .A(n8056), .ZN(n8060) );
  OAI21_X1 U9616 ( .B1(n8061), .B2(n8060), .A(n8059), .ZN(n8062) );
  NAND3_X1 U9617 ( .A1(n8066), .A2(n6293), .A3(n6123), .ZN(n8064) );
  MUX2_X1 U9618 ( .A(n8070), .B(P2_DATAO_REG_30__SCAN_IN), .S(n8085), .Z(
        P2_U3582) );
  MUX2_X1 U9619 ( .A(n4777), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8085), .Z(
        P2_U3580) );
  MUX2_X1 U9620 ( .A(n8224), .B(P2_DATAO_REG_27__SCAN_IN), .S(n8085), .Z(
        P2_U3579) );
  MUX2_X1 U9621 ( .A(n8223), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8085), .Z(
        P2_U3578) );
  MUX2_X1 U9622 ( .A(n8305), .B(P2_DATAO_REG_25__SCAN_IN), .S(n8085), .Z(
        P2_U3577) );
  MUX2_X1 U9623 ( .A(n8217), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8085), .Z(
        P2_U3576) );
  MUX2_X1 U9624 ( .A(n8304), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8085), .Z(
        P2_U3575) );
  MUX2_X1 U9625 ( .A(n8359), .B(P2_DATAO_REG_22__SCAN_IN), .S(n8085), .Z(
        P2_U3574) );
  MUX2_X1 U9626 ( .A(n8373), .B(P2_DATAO_REG_21__SCAN_IN), .S(n8085), .Z(
        P2_U3573) );
  MUX2_X1 U9627 ( .A(n8358), .B(P2_DATAO_REG_20__SCAN_IN), .S(n8085), .Z(
        P2_U3572) );
  MUX2_X1 U9628 ( .A(n8402), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8085), .Z(
        P2_U3571) );
  MUX2_X1 U9629 ( .A(n8416), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8085), .Z(
        P2_U3570) );
  MUX2_X1 U9630 ( .A(n8439), .B(P2_DATAO_REG_17__SCAN_IN), .S(n8085), .Z(
        P2_U3569) );
  MUX2_X1 U9631 ( .A(n8415), .B(P2_DATAO_REG_16__SCAN_IN), .S(n8085), .Z(
        P2_U3568) );
  MUX2_X1 U9632 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8442), .S(P2_U3966), .Z(
        P2_U3567) );
  MUX2_X1 U9633 ( .A(n8071), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8085), .Z(
        P2_U3566) );
  MUX2_X1 U9634 ( .A(n8072), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8085), .Z(
        P2_U3565) );
  MUX2_X1 U9635 ( .A(n8073), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8085), .Z(
        P2_U3564) );
  MUX2_X1 U9636 ( .A(n8074), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8085), .Z(
        P2_U3563) );
  MUX2_X1 U9637 ( .A(n8075), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8085), .Z(
        P2_U3562) );
  MUX2_X1 U9638 ( .A(n8076), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8085), .Z(
        P2_U3561) );
  MUX2_X1 U9639 ( .A(n8077), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8085), .Z(
        P2_U3560) );
  MUX2_X1 U9640 ( .A(n8078), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8085), .Z(
        P2_U3559) );
  MUX2_X1 U9641 ( .A(n8079), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8085), .Z(
        P2_U3558) );
  MUX2_X1 U9642 ( .A(n8080), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8085), .Z(
        P2_U3557) );
  MUX2_X1 U9643 ( .A(n8081), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8085), .Z(
        P2_U3556) );
  MUX2_X1 U9644 ( .A(n8082), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8085), .Z(
        P2_U3555) );
  MUX2_X1 U9645 ( .A(n8083), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8085), .Z(
        P2_U3554) );
  MUX2_X1 U9646 ( .A(n8084), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8085), .Z(
        P2_U3553) );
  MUX2_X1 U9647 ( .A(n8086), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8085), .Z(
        P2_U3552) );
  OAI211_X1 U9648 ( .C1(n8089), .C2(n8088), .A(n9979), .B(n8087), .ZN(n8098)
         );
  AOI21_X1 U9649 ( .B1(n9985), .B2(P2_ADDR_REG_4__SCAN_IN), .A(n8090), .ZN(
        n8097) );
  OAI211_X1 U9650 ( .C1(n8093), .C2(n8092), .A(n9980), .B(n8091), .ZN(n8096)
         );
  NAND2_X1 U9651 ( .A1(n9674), .A2(n8094), .ZN(n8095) );
  NAND4_X1 U9652 ( .A1(n8098), .A2(n8097), .A3(n8096), .A4(n8095), .ZN(
        P2_U3249) );
  NAND2_X1 U9653 ( .A1(n9674), .A2(n8099), .ZN(n8110) );
  OAI211_X1 U9654 ( .C1(n8102), .C2(n8101), .A(n9980), .B(n8100), .ZN(n8109)
         );
  AND2_X1 U9655 ( .A1(P2_U3152), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n8103) );
  AOI21_X1 U9656 ( .B1(n9985), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n8103), .ZN(
        n8108) );
  OAI211_X1 U9657 ( .C1(n8106), .C2(n8105), .A(n9979), .B(n8104), .ZN(n8107)
         );
  NAND4_X1 U9658 ( .A1(n8110), .A2(n8109), .A3(n8108), .A4(n8107), .ZN(
        P2_U3250) );
  NAND2_X1 U9659 ( .A1(n9674), .A2(n8111), .ZN(n8123) );
  OAI211_X1 U9660 ( .C1(n8114), .C2(n8113), .A(n9980), .B(n8112), .ZN(n8122)
         );
  INV_X1 U9661 ( .A(n8115), .ZN(n8116) );
  AOI21_X1 U9662 ( .B1(n9985), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n8116), .ZN(
        n8121) );
  OAI211_X1 U9663 ( .C1(n8119), .C2(n8118), .A(n9979), .B(n8117), .ZN(n8120)
         );
  NAND4_X1 U9664 ( .A1(n8123), .A2(n8122), .A3(n8121), .A4(n8120), .ZN(
        P2_U3251) );
  NAND2_X1 U9665 ( .A1(n9674), .A2(n8124), .ZN(n8135) );
  OAI211_X1 U9666 ( .C1(n8127), .C2(n8126), .A(n9980), .B(n8125), .ZN(n8134)
         );
  NOR2_X1 U9667 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9590), .ZN(n8128) );
  AOI21_X1 U9668 ( .B1(n9985), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n8128), .ZN(
        n8133) );
  OAI211_X1 U9669 ( .C1(n8131), .C2(n8130), .A(n9979), .B(n8129), .ZN(n8132)
         );
  NAND4_X1 U9670 ( .A1(n8135), .A2(n8134), .A3(n8133), .A4(n8132), .ZN(
        P2_U3253) );
  NAND2_X1 U9671 ( .A1(n9674), .A2(n8136), .ZN(n8148) );
  OAI211_X1 U9672 ( .C1(n8139), .C2(n8138), .A(n9980), .B(n8137), .ZN(n8147)
         );
  INV_X1 U9673 ( .A(n8140), .ZN(n8141) );
  AOI21_X1 U9674 ( .B1(n9985), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n8141), .ZN(
        n8146) );
  OAI211_X1 U9675 ( .C1(n8144), .C2(n8143), .A(n9979), .B(n8142), .ZN(n8145)
         );
  NAND4_X1 U9676 ( .A1(n8148), .A2(n8147), .A3(n8146), .A4(n8145), .ZN(
        P2_U3254) );
  NAND2_X1 U9677 ( .A1(n8150), .A2(n8149), .ZN(n8152) );
  INV_X1 U9678 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8428) );
  XNOR2_X1 U9679 ( .A(n8171), .B(n8428), .ZN(n8151) );
  NAND2_X1 U9680 ( .A1(n8151), .A2(n8152), .ZN(n8166) );
  OAI211_X1 U9681 ( .C1(n8152), .C2(n8151), .A(n9980), .B(n8166), .ZN(n8165)
         );
  XNOR2_X1 U9682 ( .A(n8171), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n8157) );
  OR2_X1 U9683 ( .A1(n8153), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n8155) );
  NAND2_X1 U9684 ( .A1(n8155), .A2(n8154), .ZN(n8156) );
  NAND2_X1 U9685 ( .A1(n8157), .A2(n8156), .ZN(n8159) );
  NOR2_X1 U9686 ( .A1(n8157), .A2(n8156), .ZN(n8170) );
  INV_X1 U9687 ( .A(n8170), .ZN(n8158) );
  NAND2_X1 U9688 ( .A1(n8159), .A2(n8158), .ZN(n8162) );
  NOR2_X1 U9689 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9500), .ZN(n8160) );
  AOI21_X1 U9690 ( .B1(n9985), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n8160), .ZN(
        n8161) );
  OAI21_X1 U9691 ( .B1(n9983), .B2(n8162), .A(n8161), .ZN(n8163) );
  AOI21_X1 U9692 ( .B1(n8171), .B2(n9674), .A(n8163), .ZN(n8164) );
  NAND2_X1 U9693 ( .A1(n8165), .A2(n8164), .ZN(P2_U3262) );
  NAND2_X1 U9694 ( .A1(n8171), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8167) );
  NAND2_X1 U9695 ( .A1(n8167), .A2(n8166), .ZN(n8168) );
  NOR2_X1 U9696 ( .A1(n8168), .A2(n8182), .ZN(n8187) );
  NOR2_X1 U9697 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n8169), .ZN(n8186) );
  AOI21_X1 U9698 ( .B1(n8169), .B2(P2_REG2_REG_18__SCAN_IN), .A(n8186), .ZN(
        n8178) );
  AOI21_X1 U9699 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n8171), .A(n8170), .ZN(
        n8180) );
  XNOR2_X1 U9700 ( .A(n8182), .B(n8172), .ZN(n8181) );
  XOR2_X1 U9701 ( .A(n8180), .B(n8181), .Z(n8175) );
  NAND2_X1 U9702 ( .A1(n9985), .A2(P2_ADDR_REG_18__SCAN_IN), .ZN(n8173) );
  OAI211_X1 U9703 ( .C1(n9983), .C2(n8175), .A(n8174), .B(n8173), .ZN(n8176)
         );
  AOI21_X1 U9704 ( .B1(n8182), .B2(n9674), .A(n8176), .ZN(n8177) );
  OAI21_X1 U9705 ( .B1(n8178), .B2(n8191), .A(n8177), .ZN(P2_U3263) );
  INV_X1 U9706 ( .A(n8179), .ZN(n8196) );
  NAND2_X1 U9707 ( .A1(n8181), .A2(n8180), .ZN(n8184) );
  OR2_X1 U9708 ( .A1(n8182), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8183) );
  NAND2_X1 U9709 ( .A1(n8184), .A2(n8183), .ZN(n8185) );
  XNOR2_X1 U9710 ( .A(n8185), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8189) );
  NAND2_X1 U9711 ( .A1(n8192), .A2(n9980), .ZN(n8188) );
  OAI211_X1 U9712 ( .C1(n8189), .C2(n9983), .A(n8188), .B(n9981), .ZN(n8194)
         );
  INV_X1 U9713 ( .A(n8189), .ZN(n8190) );
  OAI22_X1 U9714 ( .A1(n8192), .A2(n8191), .B1(n8190), .B2(n9983), .ZN(n8193)
         );
  AOI211_X1 U9715 ( .C1(P2_ADDR_REG_19__SCAN_IN), .C2(n9985), .A(n8196), .B(
        n8195), .ZN(n8197) );
  INV_X1 U9716 ( .A(n8197), .ZN(P2_U3264) );
  INV_X1 U9717 ( .A(n8467), .ZN(n8235) );
  OR2_X1 U9718 ( .A1(n8449), .A2(n8530), .ZN(n8419) );
  NOR2_X2 U9719 ( .A1(n8419), .A2(n8525), .ZN(n8395) );
  AND2_X2 U9720 ( .A1(n8395), .A2(n8390), .ZN(n8384) );
  INV_X1 U9721 ( .A(n8514), .ZN(n8371) );
  NOR2_X2 U9722 ( .A1(n8255), .A2(n8471), .ZN(n8241) );
  NAND2_X1 U9723 ( .A1(n8235), .A2(n8241), .ZN(n8232) );
  INV_X1 U9724 ( .A(P2_B_REG_SCAN_IN), .ZN(n8201) );
  OAI21_X1 U9725 ( .B1(n8202), .B2(n8201), .A(n8440), .ZN(n8231) );
  NOR2_X1 U9726 ( .A1(n8203), .A2(n8231), .ZN(n9691) );
  INV_X1 U9727 ( .A(n9691), .ZN(n9695) );
  NOR2_X1 U9728 ( .A1(n8463), .A2(n9695), .ZN(n8206) );
  AOI21_X1 U9729 ( .B1(n8463), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8206), .ZN(
        n8205) );
  NAND2_X1 U9730 ( .A1(n9692), .A2(n8430), .ZN(n8204) );
  OAI211_X1 U9731 ( .C1(n9690), .C2(n8332), .A(n8205), .B(n8204), .ZN(P2_U3265) );
  XNOR2_X1 U9732 ( .A(n9696), .B(n8232), .ZN(n9698) );
  NAND2_X1 U9733 ( .A1(n9698), .A2(n8461), .ZN(n8208) );
  AOI21_X1 U9734 ( .B1(n8463), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8206), .ZN(
        n8207) );
  OAI211_X1 U9735 ( .C1(n9696), .C2(n8455), .A(n8208), .B(n8207), .ZN(P2_U3266) );
  INV_X1 U9736 ( .A(n8525), .ZN(n8399) );
  OAI21_X1 U9737 ( .B1(n8442), .B2(n8539), .A(n8209), .ZN(n8435) );
  INV_X1 U9738 ( .A(n8437), .ZN(n8436) );
  NAND2_X1 U9739 ( .A1(n8509), .A2(n8373), .ZN(n8215) );
  INV_X1 U9740 ( .A(n8509), .ZN(n8355) );
  INV_X1 U9741 ( .A(n8302), .ZN(n8309) );
  NAND2_X1 U9742 ( .A1(n8218), .A2(n8323), .ZN(n8219) );
  NAND2_X2 U9743 ( .A1(n8308), .A2(n8219), .ZN(n8288) );
  INV_X1 U9744 ( .A(n8488), .ZN(n8298) );
  INV_X1 U9745 ( .A(n8244), .ZN(n8225) );
  INV_X1 U9746 ( .A(n8229), .ZN(n8226) );
  XNOR2_X1 U9747 ( .A(n8227), .B(n8226), .ZN(n8464) );
  INV_X1 U9748 ( .A(n8464), .ZN(n8239) );
  OAI21_X1 U9749 ( .B1(n8235), .B2(n8241), .A(n8232), .ZN(n8466) );
  NOR2_X1 U9750 ( .A1(n8466), .A2(n8332), .ZN(n8237) );
  AOI22_X1 U9751 ( .A1(n8233), .A2(n8452), .B1(P2_REG2_REG_29__SCAN_IN), .B2(
        n8463), .ZN(n8234) );
  OAI21_X1 U9752 ( .B1(n8235), .B2(n8455), .A(n8234), .ZN(n8236) );
  AOI211_X1 U9753 ( .C1(n8465), .C2(n8422), .A(n8237), .B(n8236), .ZN(n8238)
         );
  OAI21_X1 U9754 ( .B1(n8239), .B2(n8407), .A(n8238), .ZN(P2_U3267) );
  XNOR2_X1 U9755 ( .A(n8240), .B(n8244), .ZN(n8475) );
  AOI21_X1 U9756 ( .B1(n8471), .B2(n8255), .A(n8241), .ZN(n8472) );
  AOI22_X1 U9757 ( .A1(n8242), .A2(n8452), .B1(P2_REG2_REG_28__SCAN_IN), .B2(
        n8463), .ZN(n8243) );
  OAI21_X1 U9758 ( .B1(n4778), .B2(n8455), .A(n8243), .ZN(n8251) );
  AOI211_X1 U9759 ( .C1(n8245), .C2(n8244), .A(n8444), .B(n4359), .ZN(n8249)
         );
  OAI22_X1 U9760 ( .A1(n8247), .A2(n8324), .B1(n8246), .B2(n8326), .ZN(n8248)
         );
  NOR2_X1 U9761 ( .A1(n8249), .A2(n8248), .ZN(n8474) );
  NOR2_X1 U9762 ( .A1(n8474), .A2(n8463), .ZN(n8250) );
  AOI211_X1 U9763 ( .C1(n8461), .C2(n8472), .A(n8251), .B(n8250), .ZN(n8252)
         );
  OAI21_X1 U9764 ( .B1(n8475), .B2(n8407), .A(n8252), .ZN(P2_U3268) );
  XNOR2_X1 U9765 ( .A(n8254), .B(n8253), .ZN(n8480) );
  AOI21_X1 U9766 ( .B1(n8476), .B2(n8278), .A(n8199), .ZN(n8477) );
  AOI22_X1 U9767 ( .A1(n8256), .A2(n8452), .B1(P2_REG2_REG_27__SCAN_IN), .B2(
        n8463), .ZN(n8257) );
  OAI21_X1 U9768 ( .B1(n8258), .B2(n8455), .A(n8257), .ZN(n8267) );
  AOI211_X1 U9769 ( .C1(n8261), .C2(n8260), .A(n8444), .B(n8259), .ZN(n8265)
         );
  OAI22_X1 U9770 ( .A1(n8263), .A2(n8324), .B1(n8262), .B2(n8326), .ZN(n8264)
         );
  NOR2_X1 U9771 ( .A1(n8265), .A2(n8264), .ZN(n8479) );
  NOR2_X1 U9772 ( .A1(n8479), .A2(n8463), .ZN(n8266) );
  AOI211_X1 U9773 ( .C1(n8461), .C2(n8477), .A(n8267), .B(n8266), .ZN(n8268)
         );
  OAI21_X1 U9774 ( .B1(n8480), .B2(n8407), .A(n8268), .ZN(P2_U3269) );
  XNOR2_X1 U9775 ( .A(n8270), .B(n8269), .ZN(n8485) );
  AOI22_X1 U9776 ( .A1(n8483), .A2(n8430), .B1(n8463), .B2(
        P2_REG2_REG_26__SCAN_IN), .ZN(n8287) );
  INV_X1 U9777 ( .A(n8271), .ZN(n8275) );
  AOI21_X1 U9778 ( .B1(n8289), .B2(n8273), .A(n8272), .ZN(n8274) );
  NOR2_X1 U9779 ( .A1(n8275), .A2(n8274), .ZN(n8277) );
  OAI21_X1 U9780 ( .B1(n8277), .B2(n8444), .A(n8276), .ZN(n8481) );
  INV_X1 U9781 ( .A(n8294), .ZN(n8280) );
  INV_X1 U9782 ( .A(n8278), .ZN(n8279) );
  AOI211_X1 U9783 ( .C1(n8483), .C2(n8280), .A(n10022), .B(n8279), .ZN(n8482)
         );
  INV_X1 U9784 ( .A(n8482), .ZN(n8284) );
  INV_X1 U9785 ( .A(n8281), .ZN(n8282) );
  OAI22_X1 U9786 ( .A1(n8284), .A2(n8283), .B1(n8426), .B2(n8282), .ZN(n8285)
         );
  OAI21_X1 U9787 ( .B1(n8481), .B2(n8285), .A(n8422), .ZN(n8286) );
  OAI211_X1 U9788 ( .C1(n8485), .C2(n8407), .A(n8287), .B(n8286), .ZN(P2_U3270) );
  XNOR2_X1 U9789 ( .A(n8288), .B(n8291), .ZN(n8490) );
  OAI211_X1 U9790 ( .C1(n8291), .C2(n8290), .A(n8289), .B(n8411), .ZN(n8293)
         );
  NAND2_X1 U9791 ( .A1(n8293), .A2(n8292), .ZN(n8486) );
  AOI211_X1 U9792 ( .C1(n8488), .C2(n8311), .A(n10022), .B(n8294), .ZN(n8487)
         );
  NAND2_X1 U9793 ( .A1(n8487), .A2(n8386), .ZN(n8297) );
  AOI22_X1 U9794 ( .A1(n8463), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n8295), .B2(
        n8452), .ZN(n8296) );
  OAI211_X1 U9795 ( .C1(n8298), .C2(n8455), .A(n8297), .B(n8296), .ZN(n8299)
         );
  AOI21_X1 U9796 ( .B1(n8486), .B2(n8422), .A(n8299), .ZN(n8300) );
  OAI21_X1 U9797 ( .B1(n8490), .B2(n8407), .A(n8300), .ZN(P2_U3271) );
  OAI211_X1 U9798 ( .C1(n8303), .C2(n8302), .A(n8301), .B(n8411), .ZN(n8307)
         );
  AOI22_X1 U9799 ( .A1(n8305), .A2(n8440), .B1(n8441), .B2(n8304), .ZN(n8306)
         );
  AND2_X1 U9800 ( .A1(n8307), .A2(n8306), .ZN(n8495) );
  OAI21_X1 U9801 ( .B1(n8310), .B2(n8309), .A(n8308), .ZN(n8491) );
  NAND2_X1 U9802 ( .A1(n8491), .A2(n8379), .ZN(n8318) );
  INV_X1 U9803 ( .A(n8311), .ZN(n8312) );
  AOI21_X1 U9804 ( .B1(n8492), .B2(n8327), .A(n8312), .ZN(n8493) );
  INV_X1 U9805 ( .A(n8313), .ZN(n8314) );
  AOI22_X1 U9806 ( .A1(n8463), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n8314), .B2(
        n8452), .ZN(n8315) );
  OAI21_X1 U9807 ( .B1(n8218), .B2(n8455), .A(n8315), .ZN(n8316) );
  AOI21_X1 U9808 ( .B1(n8493), .B2(n8461), .A(n8316), .ZN(n8317) );
  OAI211_X1 U9809 ( .C1(n8463), .C2(n8495), .A(n8318), .B(n8317), .ZN(P2_U3272) );
  AOI21_X1 U9810 ( .B1(n8321), .B2(n8320), .A(n8319), .ZN(n8322) );
  OAI222_X1 U9811 ( .A1(n8326), .A2(n8325), .B1(n8324), .B2(n8323), .C1(n8444), 
        .C2(n8322), .ZN(n8502) );
  OAI21_X1 U9812 ( .B1(n8499), .B2(n4391), .A(n8327), .ZN(n8500) );
  AOI22_X1 U9813 ( .A1(n8463), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n8328), .B2(
        n8452), .ZN(n8331) );
  NAND2_X1 U9814 ( .A1(n8329), .A2(n8430), .ZN(n8330) );
  OAI211_X1 U9815 ( .C1(n8500), .C2(n8332), .A(n8331), .B(n8330), .ZN(n8336)
         );
  AND2_X1 U9816 ( .A1(n8334), .A2(n8333), .ZN(n8497) );
  NOR3_X1 U9817 ( .A1(n8498), .A2(n8497), .A3(n8407), .ZN(n8335) );
  AOI211_X1 U9818 ( .C1(n8422), .C2(n8502), .A(n8336), .B(n8335), .ZN(n8337)
         );
  INV_X1 U9819 ( .A(n8337), .ZN(P2_U3273) );
  XNOR2_X1 U9820 ( .A(n8339), .B(n8338), .ZN(n8508) );
  AOI21_X1 U9821 ( .B1(n8504), .B2(n8351), .A(n4391), .ZN(n8505) );
  AOI22_X1 U9822 ( .A1(n8463), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8340), .B2(
        n8452), .ZN(n8341) );
  OAI21_X1 U9823 ( .B1(n4671), .B2(n8455), .A(n8341), .ZN(n8348) );
  OAI211_X1 U9824 ( .C1(n8344), .C2(n8343), .A(n8342), .B(n8411), .ZN(n8346)
         );
  NOR2_X1 U9825 ( .A1(n8507), .A2(n8463), .ZN(n8347) );
  AOI211_X1 U9826 ( .C1(n8505), .C2(n8461), .A(n8348), .B(n8347), .ZN(n8349)
         );
  OAI21_X1 U9827 ( .B1(n8508), .B2(n8407), .A(n8349), .ZN(P2_U3274) );
  XNOR2_X1 U9828 ( .A(n8350), .B(n8356), .ZN(n8513) );
  INV_X1 U9829 ( .A(n8351), .ZN(n8352) );
  AOI21_X1 U9830 ( .B1(n8509), .B2(n8365), .A(n8352), .ZN(n8510) );
  AOI22_X1 U9831 ( .A1(n8463), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8353), .B2(
        n8452), .ZN(n8354) );
  OAI21_X1 U9832 ( .B1(n8355), .B2(n8455), .A(n8354), .ZN(n8362) );
  XNOR2_X1 U9833 ( .A(n8357), .B(n8356), .ZN(n8360) );
  AOI222_X1 U9834 ( .A1(n8411), .A2(n8360), .B1(n8359), .B2(n8440), .C1(n8358), 
        .C2(n8441), .ZN(n8512) );
  NOR2_X1 U9835 ( .A1(n8512), .A2(n8463), .ZN(n8361) );
  AOI211_X1 U9836 ( .C1(n8510), .C2(n8461), .A(n8362), .B(n8361), .ZN(n8363)
         );
  OAI21_X1 U9837 ( .B1(n8407), .B2(n8513), .A(n8363), .ZN(P2_U3275) );
  XNOR2_X1 U9838 ( .A(n8364), .B(n4376), .ZN(n8518) );
  INV_X1 U9839 ( .A(n8384), .ZN(n8367) );
  INV_X1 U9840 ( .A(n8365), .ZN(n8366) );
  AOI21_X1 U9841 ( .B1(n8514), .B2(n8367), .A(n8366), .ZN(n8515) );
  INV_X1 U9842 ( .A(n8368), .ZN(n8369) );
  AOI22_X1 U9843 ( .A1(n8463), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8369), .B2(
        n8452), .ZN(n8370) );
  OAI21_X1 U9844 ( .B1(n8371), .B2(n8455), .A(n8370), .ZN(n8376) );
  XNOR2_X1 U9845 ( .A(n8372), .B(n4376), .ZN(n8374) );
  AOI222_X1 U9846 ( .A1(n8411), .A2(n8374), .B1(n8373), .B2(n8440), .C1(n8402), 
        .C2(n8441), .ZN(n8517) );
  NOR2_X1 U9847 ( .A1(n8517), .A2(n8463), .ZN(n8375) );
  AOI211_X1 U9848 ( .C1(n8515), .C2(n8461), .A(n8376), .B(n8375), .ZN(n8377)
         );
  OAI21_X1 U9849 ( .B1(n8407), .B2(n8518), .A(n8377), .ZN(P2_U3276) );
  XNOR2_X1 U9850 ( .A(n8378), .B(n8381), .ZN(n8523) );
  XOR2_X1 U9851 ( .A(n8381), .B(n8380), .Z(n8383) );
  OAI21_X1 U9852 ( .B1(n8383), .B2(n8444), .A(n8382), .ZN(n8519) );
  INV_X1 U9853 ( .A(n8395), .ZN(n8385) );
  AOI211_X1 U9854 ( .C1(n8521), .C2(n8385), .A(n10022), .B(n8384), .ZN(n8520)
         );
  NAND2_X1 U9855 ( .A1(n8520), .A2(n8386), .ZN(n8389) );
  AOI22_X1 U9856 ( .A1(n8463), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n8387), .B2(
        n8452), .ZN(n8388) );
  OAI211_X1 U9857 ( .C1(n8390), .C2(n8455), .A(n8389), .B(n8388), .ZN(n8391)
         );
  AOI21_X1 U9858 ( .B1(n8519), .B2(n8422), .A(n8391), .ZN(n8392) );
  OAI21_X1 U9859 ( .B1(n8523), .B2(n8407), .A(n8392), .ZN(P2_U3277) );
  XNOR2_X1 U9860 ( .A(n8394), .B(n8393), .ZN(n8529) );
  AOI21_X1 U9861 ( .B1(n8525), .B2(n8419), .A(n8395), .ZN(n8526) );
  INV_X1 U9862 ( .A(n8396), .ZN(n8397) );
  AOI22_X1 U9863 ( .A1(n8463), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8397), .B2(
        n8452), .ZN(n8398) );
  OAI21_X1 U9864 ( .B1(n8399), .B2(n8455), .A(n8398), .ZN(n8405) );
  XNOR2_X1 U9865 ( .A(n8401), .B(n8400), .ZN(n8403) );
  AOI222_X1 U9866 ( .A1(n8411), .A2(n8403), .B1(n8402), .B2(n8440), .C1(n8439), 
        .C2(n8441), .ZN(n8528) );
  NOR2_X1 U9867 ( .A1(n8528), .A2(n8463), .ZN(n8404) );
  AOI211_X1 U9868 ( .C1(n8526), .C2(n8461), .A(n8405), .B(n8404), .ZN(n8406)
         );
  OAI21_X1 U9869 ( .B1(n8529), .B2(n8407), .A(n8406), .ZN(P2_U3278) );
  OAI21_X1 U9870 ( .B1(n8410), .B2(n8409), .A(n8408), .ZN(n8531) );
  INV_X1 U9871 ( .A(n8531), .ZN(n8433) );
  OAI211_X1 U9872 ( .C1(n8414), .C2(n8413), .A(n8412), .B(n8411), .ZN(n8418)
         );
  AOI22_X1 U9873 ( .A1(n8416), .A2(n8440), .B1(n8441), .B2(n8415), .ZN(n8417)
         );
  NAND2_X1 U9874 ( .A1(n8418), .A2(n8417), .ZN(n8424) );
  AOI21_X1 U9875 ( .B1(n8449), .B2(n8530), .A(n10022), .ZN(n8420) );
  AOI21_X1 U9876 ( .B1(n8420), .B2(n8419), .A(n8424), .ZN(n8532) );
  OAI21_X1 U9877 ( .B1(n8433), .B2(n8421), .A(n8532), .ZN(n8423) );
  OAI211_X1 U9878 ( .C1(n8425), .C2(n8424), .A(n8423), .B(n8422), .ZN(n8432)
         );
  OAI22_X1 U9879 ( .A1(n8422), .A2(n8428), .B1(n8427), .B2(n8426), .ZN(n8429)
         );
  AOI21_X1 U9880 ( .B1(n8530), .B2(n8430), .A(n8429), .ZN(n8431) );
  OAI211_X1 U9881 ( .C1(n8433), .C2(n8458), .A(n8432), .B(n8431), .ZN(P2_U3279) );
  AOI21_X1 U9882 ( .B1(n8436), .B2(n8435), .A(n8434), .ZN(n8457) );
  XNOR2_X1 U9883 ( .A(n8438), .B(n8437), .ZN(n8445) );
  AOI22_X1 U9884 ( .A1(n8442), .A2(n8441), .B1(n8440), .B2(n8439), .ZN(n8443)
         );
  OAI21_X1 U9885 ( .B1(n8445), .B2(n8444), .A(n8443), .ZN(n8446) );
  AOI21_X1 U9886 ( .B1(n8457), .B2(n8447), .A(n8446), .ZN(n8537) );
  INV_X1 U9887 ( .A(n8448), .ZN(n8451) );
  INV_X1 U9888 ( .A(n8449), .ZN(n8450) );
  AOI21_X1 U9889 ( .B1(n8534), .B2(n8451), .A(n8450), .ZN(n8535) );
  AOI22_X1 U9890 ( .A1(n8463), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n8453), .B2(
        n8452), .ZN(n8454) );
  OAI21_X1 U9891 ( .B1(n8456), .B2(n8455), .A(n8454), .ZN(n8460) );
  INV_X1 U9892 ( .A(n8457), .ZN(n8538) );
  NOR2_X1 U9893 ( .A1(n8538), .A2(n8458), .ZN(n8459) );
  AOI211_X1 U9894 ( .C1(n8535), .C2(n8461), .A(n8460), .B(n8459), .ZN(n8462)
         );
  OAI21_X1 U9895 ( .B1(n8463), .B2(n8537), .A(n8462), .ZN(P2_U3280) );
  NOR2_X1 U9896 ( .A1(n8466), .A2(n10022), .ZN(n8469) );
  MUX2_X1 U9897 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n8555), .S(n10048), .Z(
        P2_U3549) );
  AOI22_X1 U9898 ( .A1(n8472), .A2(n7178), .B1(n9693), .B2(n8471), .ZN(n8473)
         );
  OAI211_X1 U9899 ( .C1(n8475), .C2(n8549), .A(n8474), .B(n8473), .ZN(n8556)
         );
  MUX2_X1 U9900 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n8556), .S(n10048), .Z(
        P2_U3548) );
  AOI22_X1 U9901 ( .A1(n8477), .A2(n7178), .B1(n9693), .B2(n8476), .ZN(n8478)
         );
  OAI211_X1 U9902 ( .C1(n8480), .C2(n8549), .A(n8479), .B(n8478), .ZN(n8557)
         );
  MUX2_X1 U9903 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8557), .S(n10048), .Z(
        P2_U3547) );
  AOI211_X1 U9904 ( .C1(n9693), .C2(n8483), .A(n8482), .B(n8481), .ZN(n8484)
         );
  OAI21_X1 U9905 ( .B1(n8485), .B2(n8549), .A(n8484), .ZN(n8558) );
  MUX2_X1 U9906 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n8558), .S(n10048), .Z(
        P2_U3546) );
  AOI211_X1 U9907 ( .C1(n9693), .C2(n8488), .A(n8487), .B(n8486), .ZN(n8489)
         );
  OAI21_X1 U9908 ( .B1(n8490), .B2(n8549), .A(n8489), .ZN(n8559) );
  MUX2_X1 U9909 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8559), .S(n10048), .Z(
        P2_U3545) );
  INV_X1 U9910 ( .A(n8491), .ZN(n8496) );
  AOI22_X1 U9911 ( .A1(n8493), .A2(n7178), .B1(n9693), .B2(n8492), .ZN(n8494)
         );
  OAI211_X1 U9912 ( .C1(n8496), .C2(n8549), .A(n8495), .B(n8494), .ZN(n8560)
         );
  MUX2_X1 U9913 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8560), .S(n10048), .Z(
        P2_U3544) );
  NOR3_X1 U9914 ( .A1(n8498), .A2(n8497), .A3(n8549), .ZN(n8503) );
  OAI22_X1 U9915 ( .A1(n8500), .A2(n10022), .B1(n8499), .B2(n10031), .ZN(n8501) );
  MUX2_X1 U9916 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8561), .S(n10048), .Z(
        P2_U3543) );
  AOI22_X1 U9917 ( .A1(n8505), .A2(n7178), .B1(n9693), .B2(n8504), .ZN(n8506)
         );
  OAI211_X1 U9918 ( .C1(n8508), .C2(n8549), .A(n8507), .B(n8506), .ZN(n8562)
         );
  MUX2_X1 U9919 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n8562), .S(n10048), .Z(
        P2_U3542) );
  AOI22_X1 U9920 ( .A1(n8510), .A2(n7178), .B1(n9693), .B2(n8509), .ZN(n8511)
         );
  OAI211_X1 U9921 ( .C1(n8513), .C2(n8549), .A(n8512), .B(n8511), .ZN(n8563)
         );
  MUX2_X1 U9922 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n8563), .S(n10048), .Z(
        P2_U3541) );
  AOI22_X1 U9923 ( .A1(n8515), .A2(n7178), .B1(n9693), .B2(n8514), .ZN(n8516)
         );
  OAI211_X1 U9924 ( .C1(n8518), .C2(n8549), .A(n8517), .B(n8516), .ZN(n8564)
         );
  MUX2_X1 U9925 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n8564), .S(n10048), .Z(
        P2_U3540) );
  AOI211_X1 U9926 ( .C1(n9693), .C2(n8521), .A(n8520), .B(n8519), .ZN(n8522)
         );
  OAI21_X1 U9927 ( .B1(n8523), .B2(n8549), .A(n8522), .ZN(n8565) );
  MUX2_X1 U9928 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8565), .S(n10048), .Z(
        P2_U3539) );
  AOI22_X1 U9929 ( .A1(n8526), .A2(n7178), .B1(n9693), .B2(n8525), .ZN(n8527)
         );
  OAI211_X1 U9930 ( .C1(n8529), .C2(n8549), .A(n8528), .B(n8527), .ZN(n8566)
         );
  MUX2_X1 U9931 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n8566), .S(n10048), .Z(
        P2_U3538) );
  NAND2_X1 U9932 ( .A1(n8531), .A2(n10034), .ZN(n8533) );
  OAI211_X1 U9933 ( .C1(n8211), .C2(n10031), .A(n8533), .B(n8532), .ZN(n8567)
         );
  MUX2_X1 U9934 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8567), .S(n10048), .Z(
        P2_U3537) );
  AOI22_X1 U9935 ( .A1(n8535), .A2(n7178), .B1(n9693), .B2(n8534), .ZN(n8536)
         );
  OAI211_X1 U9936 ( .C1(n8538), .C2(n10006), .A(n8537), .B(n8536), .ZN(n8568)
         );
  MUX2_X1 U9937 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8568), .S(n10048), .Z(
        P2_U3536) );
  AOI22_X1 U9938 ( .A1(n8540), .A2(n7178), .B1(n9693), .B2(n8539), .ZN(n8541)
         );
  OAI211_X1 U9939 ( .C1(n8549), .C2(n8543), .A(n8542), .B(n8541), .ZN(n8569)
         );
  MUX2_X1 U9940 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n8569), .S(n10048), .Z(
        P2_U3535) );
  AOI22_X1 U9941 ( .A1(n8545), .A2(n7178), .B1(n9693), .B2(n8544), .ZN(n8546)
         );
  OAI211_X1 U9942 ( .C1(n8549), .C2(n8548), .A(n8547), .B(n8546), .ZN(n8570)
         );
  MUX2_X1 U9943 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n8570), .S(n10048), .Z(
        P2_U3534) );
  AOI22_X1 U9944 ( .A1(n8551), .A2(n7178), .B1(n9693), .B2(n8550), .ZN(n8552)
         );
  OAI211_X1 U9945 ( .C1(n10006), .C2(n8554), .A(n8553), .B(n8552), .ZN(n8571)
         );
  MUX2_X1 U9946 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n8571), .S(n10048), .Z(
        P2_U3533) );
  MUX2_X1 U9947 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n8555), .S(n4314), .Z(
        P2_U3517) );
  MUX2_X1 U9948 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n8556), .S(n4314), .Z(
        P2_U3516) );
  MUX2_X1 U9949 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8557), .S(n4314), .Z(
        P2_U3515) );
  MUX2_X1 U9950 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n8558), .S(n4314), .Z(
        P2_U3514) );
  MUX2_X1 U9951 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n8559), .S(n4314), .Z(
        P2_U3513) );
  MUX2_X1 U9952 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n8560), .S(n4314), .Z(
        P2_U3512) );
  MUX2_X1 U9953 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n8561), .S(n4314), .Z(
        P2_U3511) );
  MUX2_X1 U9954 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n8562), .S(n4314), .Z(
        P2_U3510) );
  MUX2_X1 U9955 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n8563), .S(n4314), .Z(
        P2_U3509) );
  MUX2_X1 U9956 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n8564), .S(n4314), .Z(
        P2_U3508) );
  MUX2_X1 U9957 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n8565), .S(n4314), .Z(
        P2_U3507) );
  MUX2_X1 U9958 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n8566), .S(n4314), .Z(
        P2_U3505) );
  MUX2_X1 U9959 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n8567), .S(n4314), .Z(
        P2_U3502) );
  MUX2_X1 U9960 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n8568), .S(n4314), .Z(
        P2_U3499) );
  MUX2_X1 U9961 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n8569), .S(n4314), .Z(
        P2_U3496) );
  MUX2_X1 U9962 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n8570), .S(n4314), .Z(
        P2_U3493) );
  MUX2_X1 U9963 ( .A(P2_REG0_REG_13__SCAN_IN), .B(n8571), .S(n4314), .Z(
        P2_U3490) );
  INV_X1 U9964 ( .A(n8794), .ZN(n9414) );
  NOR4_X1 U9965 ( .A1(n8573), .A2(P2_IR_REG_30__SCAN_IN), .A3(n8572), .A4(
        P2_U3152), .ZN(n8574) );
  AOI21_X1 U9966 ( .B1(n8583), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n8574), .ZN(
        n8575) );
  OAI21_X1 U9967 ( .B1(n9414), .B2(n6195), .A(n8575), .ZN(P2_U3327) );
  INV_X1 U9968 ( .A(n8790), .ZN(n9417) );
  AOI22_X1 U9969 ( .A1(n8576), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n8588), .ZN(n8577) );
  OAI21_X1 U9970 ( .B1(n9417), .B2(n6195), .A(n8577), .ZN(P2_U3328) );
  INV_X1 U9971 ( .A(n8578), .ZN(n9421) );
  AOI22_X1 U9972 ( .A1(n8579), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n8588), .ZN(n8580) );
  OAI21_X1 U9973 ( .B1(n9421), .B2(n6195), .A(n8580), .ZN(P2_U3329) );
  INV_X1 U9974 ( .A(n8581), .ZN(n9424) );
  AOI21_X1 U9975 ( .B1(n8583), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n8582), .ZN(
        n8584) );
  OAI21_X1 U9976 ( .B1(n9424), .B2(n6195), .A(n8584), .ZN(P2_U3330) );
  INV_X1 U9977 ( .A(n6067), .ZN(n9427) );
  AOI22_X1 U9978 ( .A1(n8585), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_27__SCAN_IN), .B2(n8588), .ZN(n8586) );
  OAI21_X1 U9979 ( .B1(n9427), .B2(n6195), .A(n8586), .ZN(P2_U3331) );
  INV_X1 U9980 ( .A(n8587), .ZN(n9431) );
  AOI22_X1 U9981 ( .A1(n8589), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n8588), .ZN(n8590) );
  OAI21_X1 U9982 ( .B1(n9431), .B2(n6195), .A(n8590), .ZN(P2_U3332) );
  MUX2_X1 U9983 ( .A(n8591), .B(n9990), .S(P2_STATE_REG_SCAN_IN), .Z(P2_U3358)
         );
  NAND2_X1 U9984 ( .A1(n8592), .A2(n4337), .ZN(n8593) );
  XOR2_X1 U9985 ( .A(n8594), .B(n8593), .Z(n8601) );
  NAND2_X1 U9986 ( .A1(n8692), .A2(n8595), .ZN(n8598) );
  AOI21_X1 U9987 ( .B1(n8669), .B2(n8993), .A(n8596), .ZN(n8597) );
  OAI211_X1 U9988 ( .C1(n9245), .C2(n8689), .A(n8598), .B(n8597), .ZN(n8599)
         );
  AOI21_X1 U9989 ( .B1(n8719), .B2(n8638), .A(n8599), .ZN(n8600) );
  OAI21_X1 U9990 ( .B1(n8601), .B2(n8683), .A(n8600), .ZN(P1_U3213) );
  NAND2_X1 U9991 ( .A1(n8603), .A2(n8602), .ZN(n8604) );
  XOR2_X1 U9992 ( .A(n8605), .B(n8604), .Z(n8610) );
  NAND2_X1 U9993 ( .A1(n8986), .A2(n9707), .ZN(n8607) );
  AOI22_X1 U9994 ( .A1(n8987), .A2(n8669), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3084), .ZN(n8606) );
  OAI211_X1 U9995 ( .C1(n9722), .C2(n9132), .A(n8607), .B(n8606), .ZN(n8608)
         );
  AOI21_X1 U9996 ( .B1(n9319), .B2(n8638), .A(n8608), .ZN(n8609) );
  OAI21_X1 U9997 ( .B1(n8610), .B2(n8683), .A(n8609), .ZN(P1_U3214) );
  XOR2_X1 U9998 ( .A(n8611), .B(n8612), .Z(n8617) );
  NAND2_X1 U9999 ( .A1(n9707), .A2(n8989), .ZN(n8613) );
  NAND2_X1 U10000 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9046) );
  OAI211_X1 U10001 ( .C1(n9230), .C2(n9709), .A(n8613), .B(n9046), .ZN(n8614)
         );
  AOI21_X1 U10002 ( .B1(n8692), .B2(n9198), .A(n8614), .ZN(n8616) );
  NAND2_X1 U10003 ( .A1(n9341), .A2(n8638), .ZN(n8615) );
  OAI211_X1 U10004 ( .C1(n8617), .C2(n8683), .A(n8616), .B(n8615), .ZN(
        P1_U3217) );
  XOR2_X1 U10005 ( .A(n8619), .B(n8618), .Z(n8625) );
  OAI22_X1 U10006 ( .A1(n9166), .A2(n8689), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8620), .ZN(n8621) );
  AOI21_X1 U10007 ( .B1(n8669), .B2(n8989), .A(n8621), .ZN(n8622) );
  OAI21_X1 U10008 ( .B1(n9722), .B2(n9168), .A(n8622), .ZN(n8623) );
  AOI21_X1 U10009 ( .B1(n9328), .B2(n8638), .A(n8623), .ZN(n8624) );
  OAI21_X1 U10010 ( .B1(n8625), .B2(n8683), .A(n8624), .ZN(P1_U3221) );
  XOR2_X1 U10011 ( .A(n8627), .B(n8626), .Z(n8632) );
  NAND2_X1 U10012 ( .A1(n9080), .A2(n9707), .ZN(n8629) );
  AOI22_X1 U10013 ( .A1(n8986), .A2(n8669), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3084), .ZN(n8628) );
  OAI211_X1 U10014 ( .C1(n9722), .C2(n9104), .A(n8629), .B(n8628), .ZN(n8630)
         );
  AOI21_X1 U10015 ( .B1(n9310), .B2(n8638), .A(n8630), .ZN(n8631) );
  OAI21_X1 U10016 ( .B1(n8632), .B2(n8683), .A(n8631), .ZN(P1_U3223) );
  XOR2_X1 U10017 ( .A(n8633), .B(n8634), .Z(n8640) );
  NAND2_X1 U10018 ( .A1(n8692), .A2(n9248), .ZN(n8636) );
  AOI22_X1 U10019 ( .A1(n8669), .A2(n8991), .B1(P1_REG3_REG_16__SCAN_IN), .B2(
        P1_U3084), .ZN(n8635) );
  OAI211_X1 U10020 ( .C1(n9244), .C2(n8689), .A(n8636), .B(n8635), .ZN(n8637)
         );
  AOI21_X1 U10021 ( .B1(n9247), .B2(n8638), .A(n8637), .ZN(n8639) );
  OAI21_X1 U10022 ( .B1(n8640), .B2(n8683), .A(n8639), .ZN(P1_U3224) );
  XOR2_X1 U10023 ( .A(n8641), .B(n8642), .Z(n8647) );
  NAND2_X1 U10024 ( .A1(n8692), .A2(n9234), .ZN(n8644) );
  AOI22_X1 U10025 ( .A1(n9707), .A2(n8990), .B1(P1_REG3_REG_17__SCAN_IN), .B2(
        P1_U3084), .ZN(n8643) );
  OAI211_X1 U10026 ( .C1(n9256), .C2(n9709), .A(n8644), .B(n8643), .ZN(n8645)
         );
  AOI21_X1 U10027 ( .B1(n9351), .B2(n8638), .A(n8645), .ZN(n8646) );
  OAI21_X1 U10028 ( .B1(n8647), .B2(n8683), .A(n8646), .ZN(P1_U3226) );
  INV_X1 U10029 ( .A(n8649), .ZN(n8650) );
  AOI21_X1 U10030 ( .B1(n8651), .B2(n8648), .A(n8650), .ZN(n8656) );
  AOI22_X1 U10031 ( .A1(n9118), .A2(n8669), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3084), .ZN(n8653) );
  NAND2_X1 U10032 ( .A1(n8692), .A2(n9124), .ZN(n8652) );
  OAI211_X1 U10033 ( .C1(n9088), .C2(n8689), .A(n8653), .B(n8652), .ZN(n8654)
         );
  AOI21_X1 U10034 ( .B1(n9120), .B2(n8638), .A(n8654), .ZN(n8655) );
  OAI21_X1 U10035 ( .B1(n8656), .B2(n8683), .A(n8655), .ZN(P1_U3227) );
  XOR2_X1 U10036 ( .A(n8657), .B(n8658), .Z(n8664) );
  OAI22_X1 U10037 ( .A1(n9178), .A2(n8689), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8659), .ZN(n8660) );
  AOI21_X1 U10038 ( .B1(n8669), .B2(n9212), .A(n8660), .ZN(n8661) );
  OAI21_X1 U10039 ( .B1(n9722), .B2(n9184), .A(n8661), .ZN(n8662) );
  AOI21_X1 U10040 ( .B1(n9183), .B2(n8638), .A(n8662), .ZN(n8663) );
  OAI21_X1 U10041 ( .B1(n8664), .B2(n8683), .A(n8663), .ZN(P1_U3231) );
  NAND2_X1 U10042 ( .A1(n8665), .A2(n8666), .ZN(n8667) );
  XOR2_X1 U10043 ( .A(n8668), .B(n8667), .Z(n8674) );
  NAND2_X1 U10044 ( .A1(n9118), .A2(n9707), .ZN(n8671) );
  AOI22_X1 U10045 ( .A1(n8669), .A2(n8988), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3084), .ZN(n8670) );
  OAI211_X1 U10046 ( .C1(n9722), .C2(n9153), .A(n8671), .B(n8670), .ZN(n8672)
         );
  AOI21_X1 U10047 ( .B1(n9152), .B2(n8638), .A(n8672), .ZN(n8673) );
  OAI21_X1 U10048 ( .B1(n8674), .B2(n8683), .A(n8673), .ZN(P1_U3233) );
  NAND2_X1 U10049 ( .A1(n8676), .A2(n8675), .ZN(n8677) );
  XOR2_X1 U10050 ( .A(n8678), .B(n8677), .Z(n8684) );
  NAND2_X1 U10051 ( .A1(n9707), .A2(n9212), .ZN(n8679) );
  NAND2_X1 U10052 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9857) );
  OAI211_X1 U10053 ( .C1(n9244), .C2(n9709), .A(n8679), .B(n9857), .ZN(n8681)
         );
  NOR2_X1 U10054 ( .A1(n9400), .A2(n8695), .ZN(n8680) );
  AOI211_X1 U10055 ( .C1(n9220), .C2(n8692), .A(n8681), .B(n8680), .ZN(n8682)
         );
  OAI21_X1 U10056 ( .B1(n8684), .B2(n8683), .A(n8682), .ZN(P1_U3236) );
  OAI211_X1 U10057 ( .C1(n8685), .C2(n8687), .A(n8686), .B(n9717), .ZN(n8694)
         );
  OAI22_X1 U10058 ( .A1(n9088), .A2(n9709), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8688), .ZN(n8691) );
  NOR2_X1 U10059 ( .A1(n9087), .A2(n8689), .ZN(n8690) );
  AOI211_X1 U10060 ( .C1(n9093), .C2(n8692), .A(n8691), .B(n8690), .ZN(n8693)
         );
  OAI211_X1 U10061 ( .C1(n9379), .C2(n8695), .A(n8694), .B(n8693), .ZN(
        P1_U3238) );
  INV_X1 U10062 ( .A(n8984), .ZN(n8884) );
  INV_X1 U10063 ( .A(n8841), .ZN(n8696) );
  NAND2_X1 U10064 ( .A1(n8701), .A2(n8841), .ZN(n8946) );
  NAND2_X1 U10065 ( .A1(n8835), .A2(n8839), .ZN(n8840) );
  INV_X1 U10066 ( .A(n8805), .ZN(n8799) );
  MUX2_X1 U10067 ( .A(n8946), .B(n8840), .S(n8799), .Z(n8698) );
  INV_X1 U10068 ( .A(n8698), .ZN(n8699) );
  NAND2_X1 U10069 ( .A1(n8700), .A2(n8699), .ZN(n8705) );
  MUX2_X1 U10070 ( .A(n8701), .B(n8835), .S(n8805), .Z(n8703) );
  AND2_X1 U10071 ( .A1(n8703), .A2(n8702), .ZN(n8704) );
  NAND2_X1 U10072 ( .A1(n8705), .A2(n8704), .ZN(n8711) );
  AND2_X1 U10073 ( .A1(n8712), .A2(n8706), .ZN(n8836) );
  NAND2_X1 U10074 ( .A1(n8711), .A2(n8836), .ZN(n8707) );
  NAND2_X1 U10075 ( .A1(n8707), .A2(n8828), .ZN(n8708) );
  INV_X1 U10076 ( .A(n8849), .ZN(n8709) );
  NAND3_X1 U10077 ( .A1(n8711), .A2(n8710), .A3(n8949), .ZN(n8713) );
  NAND3_X1 U10078 ( .A1(n8713), .A2(n9884), .A3(n8712), .ZN(n8715) );
  NAND2_X1 U10079 ( .A1(n8728), .A2(n8716), .ZN(n8717) );
  AND2_X1 U10080 ( .A1(n8729), .A2(n9726), .ZN(n8718) );
  NAND2_X1 U10081 ( .A1(n8719), .A2(n9710), .ZN(n8724) );
  NAND2_X1 U10082 ( .A1(n8724), .A2(n8720), .ZN(n8855) );
  NAND2_X1 U10083 ( .A1(n8728), .A2(n8721), .ZN(n8829) );
  AND2_X1 U10084 ( .A1(n8829), .A2(n8729), .ZN(n8722) );
  NOR2_X1 U10085 ( .A1(n8855), .A2(n8722), .ZN(n8725) );
  NAND2_X1 U10086 ( .A1(n8732), .A2(n8723), .ZN(n8731) );
  AND2_X1 U10087 ( .A1(n8731), .A2(n8724), .ZN(n8853) );
  AOI21_X1 U10088 ( .B1(n8734), .B2(n8725), .A(n8853), .ZN(n8736) );
  INV_X1 U10089 ( .A(n8726), .ZN(n8727) );
  NAND2_X1 U10090 ( .A1(n8728), .A2(n8727), .ZN(n8730) );
  NAND2_X1 U10091 ( .A1(n8730), .A2(n8729), .ZN(n8850) );
  NOR2_X1 U10092 ( .A1(n8731), .A2(n8850), .ZN(n8733) );
  AOI22_X1 U10093 ( .A1(n8734), .A2(n8733), .B1(n8732), .B2(n8855), .ZN(n8735)
         );
  MUX2_X1 U10094 ( .A(n8736), .B(n8735), .S(n8805), .Z(n8739) );
  INV_X1 U10095 ( .A(n8920), .ZN(n9241) );
  MUX2_X1 U10096 ( .A(n8857), .B(n8862), .S(n8799), .Z(n8737) );
  NAND2_X1 U10097 ( .A1(n9241), .A2(n8737), .ZN(n8738) );
  AOI21_X1 U10098 ( .B1(n8739), .B2(n9258), .A(n8738), .ZN(n8744) );
  MUX2_X1 U10099 ( .A(n8858), .B(n8825), .S(n8805), .Z(n8740) );
  NAND2_X1 U10100 ( .A1(n8899), .A2(n8740), .ZN(n8743) );
  MUX2_X1 U10101 ( .A(n8827), .B(n8871), .S(n8805), .Z(n8741) );
  INV_X1 U10102 ( .A(n8741), .ZN(n8742) );
  OAI21_X1 U10103 ( .B1(n8744), .B2(n8743), .A(n8742), .ZN(n8748) );
  NAND3_X1 U10104 ( .A1(n8748), .A2(n8745), .A3(n8749), .ZN(n8746) );
  INV_X1 U10105 ( .A(n8756), .ZN(n8898) );
  NAND3_X1 U10106 ( .A1(n8746), .A2(n8898), .A3(n8822), .ZN(n8752) );
  AND2_X1 U10107 ( .A1(n8822), .A2(n8747), .ZN(n8872) );
  NAND2_X1 U10108 ( .A1(n8748), .A2(n8872), .ZN(n8750) );
  AND2_X1 U10109 ( .A1(n8897), .A2(n8749), .ZN(n8868) );
  NAND2_X1 U10110 ( .A1(n8750), .A2(n8868), .ZN(n8751) );
  MUX2_X1 U10111 ( .A(n8752), .B(n8751), .S(n8805), .Z(n8761) );
  INV_X1 U10112 ( .A(n8758), .ZN(n8753) );
  AOI21_X1 U10113 ( .B1(n8761), .B2(n8897), .A(n8753), .ZN(n8754) );
  NAND2_X1 U10114 ( .A1(n8896), .A2(n8757), .ZN(n8869) );
  OAI21_X1 U10115 ( .B1(n8754), .B2(n8869), .A(n8895), .ZN(n8755) );
  OR2_X1 U10116 ( .A1(n9120), .A2(n9138), .ZN(n8867) );
  NAND2_X1 U10117 ( .A1(n8757), .A2(n8756), .ZN(n8759) );
  AND2_X1 U10118 ( .A1(n8759), .A2(n8758), .ZN(n8760) );
  NAND2_X1 U10119 ( .A1(n8760), .A2(n8895), .ZN(n8824) );
  NAND2_X1 U10120 ( .A1(n8824), .A2(n8896), .ZN(n8873) );
  OAI21_X1 U10121 ( .B1(n8761), .B2(n8869), .A(n8873), .ZN(n8762) );
  NAND2_X1 U10122 ( .A1(n8762), .A2(n8805), .ZN(n8763) );
  INV_X1 U10123 ( .A(n9107), .ZN(n8764) );
  OAI21_X1 U10124 ( .B1(n8764), .B2(n8866), .A(n8820), .ZN(n8767) );
  INV_X1 U10125 ( .A(n8765), .ZN(n8959) );
  NAND2_X1 U10126 ( .A1(n8867), .A2(n8959), .ZN(n8766) );
  NAND2_X1 U10127 ( .A1(n8962), .A2(n8766), .ZN(n8877) );
  MUX2_X1 U10128 ( .A(n8767), .B(n8877), .S(n8799), .Z(n8768) );
  AND2_X1 U10129 ( .A1(n8820), .A2(n9110), .ZN(n8769) );
  OR2_X1 U10130 ( .A1(n8879), .A2(n8769), .ZN(n8772) );
  NOR2_X1 U10131 ( .A1(n8775), .A2(n9080), .ZN(n8770) );
  NOR2_X1 U10132 ( .A1(n8770), .A2(n9092), .ZN(n8771) );
  MUX2_X1 U10133 ( .A(n8772), .B(n8771), .S(n8805), .Z(n8773) );
  OAI21_X1 U10134 ( .B1(n8780), .B2(n8894), .A(n8773), .ZN(n8782) );
  NAND2_X1 U10135 ( .A1(n9092), .A2(n8820), .ZN(n8774) );
  NAND2_X1 U10136 ( .A1(n8880), .A2(n8774), .ZN(n8778) );
  NAND2_X1 U10137 ( .A1(n8775), .A2(n9080), .ZN(n8776) );
  NAND2_X1 U10138 ( .A1(n8821), .A2(n8776), .ZN(n8777) );
  NAND2_X1 U10139 ( .A1(n8782), .A2(n8781), .ZN(n8785) );
  MUX2_X1 U10140 ( .A(n8821), .B(n8880), .S(n8805), .Z(n8783) );
  NAND3_X1 U10141 ( .A1(n8785), .A2(n8784), .A3(n8783), .ZN(n8787) );
  MUX2_X1 U10142 ( .A(n8881), .B(n8817), .S(n8805), .Z(n8786) );
  INV_X1 U10143 ( .A(n8802), .ZN(n8800) );
  NAND2_X1 U10144 ( .A1(n5554), .A2(n8884), .ZN(n8788) );
  NAND2_X1 U10145 ( .A1(n8790), .A2(n5090), .ZN(n8792) );
  NAND2_X1 U10146 ( .A1(n8795), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n8791) );
  INV_X1 U10147 ( .A(n8983), .ZN(n8793) );
  NAND2_X1 U10148 ( .A1(n8892), .A2(n9050), .ZN(n8798) );
  NAND2_X1 U10149 ( .A1(n8794), .A2(n5090), .ZN(n8797) );
  NAND2_X1 U10150 ( .A1(n8795), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n8796) );
  NAND2_X1 U10151 ( .A1(n8983), .A2(n9050), .ZN(n8801) );
  NAND2_X1 U10152 ( .A1(n9053), .A2(n8801), .ZN(n8887) );
  INV_X1 U10153 ( .A(n8807), .ZN(n8890) );
  NAND3_X1 U10154 ( .A1(n8890), .A2(n8802), .A3(n9294), .ZN(n8804) );
  INV_X1 U10155 ( .A(n9050), .ZN(n8812) );
  AND2_X1 U10156 ( .A1(n8803), .A2(n8812), .ZN(n8926) );
  AOI21_X1 U10157 ( .B1(n8804), .B2(n8887), .A(n8926), .ZN(n8806) );
  MUX2_X1 U10158 ( .A(n8807), .B(n8806), .S(n8805), .Z(n8808) );
  INV_X1 U10159 ( .A(n8810), .ZN(n8811) );
  NAND2_X1 U10160 ( .A1(n8811), .A2(n9920), .ZN(n8815) );
  NOR2_X1 U10161 ( .A1(n8803), .A2(n8812), .ZN(n8929) );
  OR2_X1 U10162 ( .A1(n9294), .A2(n8884), .ZN(n8818) );
  AND2_X1 U10163 ( .A1(n8818), .A2(n8817), .ZN(n8886) );
  NAND4_X1 U10164 ( .A1(n8886), .A2(n8821), .A3(n8820), .A4(n8819), .ZN(n8935)
         );
  INV_X1 U10165 ( .A(n8822), .ZN(n8823) );
  NOR2_X1 U10166 ( .A1(n8824), .A2(n8823), .ZN(n8955) );
  INV_X1 U10167 ( .A(n8825), .ZN(n8826) );
  OR2_X1 U10168 ( .A1(n8827), .A2(n8826), .ZN(n8864) );
  INV_X1 U10169 ( .A(n8864), .ZN(n8833) );
  INV_X1 U10170 ( .A(n8828), .ZN(n8831) );
  AOI21_X1 U10171 ( .B1(n8849), .B2(n4396), .A(n8829), .ZN(n8852) );
  INV_X1 U10172 ( .A(n8852), .ZN(n8830) );
  NOR3_X1 U10173 ( .A1(n8855), .A2(n8831), .A3(n8830), .ZN(n8832) );
  NAND3_X1 U10174 ( .A1(n8833), .A2(n8832), .A3(n8862), .ZN(n8951) );
  INV_X1 U10175 ( .A(n8834), .ZN(n8847) );
  INV_X1 U10176 ( .A(n8835), .ZN(n8837) );
  INV_X1 U10177 ( .A(n8836), .ZN(n8845) );
  AOI21_X1 U10178 ( .B1(n8837), .B2(n8949), .A(n8845), .ZN(n8947) );
  NAND3_X1 U10179 ( .A1(n8947), .A2(n8839), .A3(n8838), .ZN(n8937) );
  AOI21_X1 U10180 ( .B1(n8841), .B2(n8944), .A(n8840), .ZN(n8844) );
  INV_X1 U10181 ( .A(n8949), .ZN(n8843) );
  NOR3_X1 U10182 ( .A1(n8844), .A2(n8843), .A3(n8842), .ZN(n8846) );
  OAI22_X1 U10183 ( .A1(n8847), .A2(n8937), .B1(n8846), .B2(n8845), .ZN(n8865)
         );
  NAND2_X1 U10184 ( .A1(n8849), .A2(n8848), .ZN(n8851) );
  AOI21_X1 U10185 ( .B1(n8852), .B2(n8851), .A(n8850), .ZN(n8856) );
  INV_X1 U10186 ( .A(n8853), .ZN(n8854) );
  OAI21_X1 U10187 ( .B1(n8856), .B2(n8855), .A(n8854), .ZN(n8861) );
  INV_X1 U10188 ( .A(n8857), .ZN(n8860) );
  INV_X1 U10189 ( .A(n8858), .ZN(n8859) );
  AOI211_X1 U10190 ( .C1(n8862), .C2(n8861), .A(n8860), .B(n8859), .ZN(n8863)
         );
  OR2_X1 U10191 ( .A1(n8864), .A2(n8863), .ZN(n8936) );
  OAI21_X1 U10192 ( .B1(n8951), .B2(n8865), .A(n8936), .ZN(n8876) );
  NAND2_X1 U10193 ( .A1(n8867), .A2(n8866), .ZN(n8963) );
  INV_X1 U10194 ( .A(n8868), .ZN(n8870) );
  AOI211_X1 U10195 ( .C1(n8872), .C2(n8871), .A(n8870), .B(n8869), .ZN(n8875)
         );
  INV_X1 U10196 ( .A(n8873), .ZN(n8874) );
  NOR2_X1 U10197 ( .A1(n8875), .A2(n8874), .ZN(n8958) );
  AOI211_X1 U10198 ( .C1(n8955), .C2(n8876), .A(n8963), .B(n8958), .ZN(n8878)
         );
  NOR2_X1 U10199 ( .A1(n8878), .A2(n8877), .ZN(n8888) );
  INV_X1 U10200 ( .A(n8879), .ZN(n8882) );
  OAI211_X1 U10201 ( .C1(n8883), .C2(n8882), .A(n8881), .B(n8880), .ZN(n8885)
         );
  AOI22_X1 U10202 ( .A1(n8886), .A2(n8885), .B1(n8884), .B2(n9294), .ZN(n8965)
         );
  OAI211_X1 U10203 ( .C1(n8935), .C2(n8888), .A(n8965), .B(n8887), .ZN(n8889)
         );
  AOI211_X1 U10204 ( .C1(n8890), .C2(n8889), .A(n5503), .B(n8929), .ZN(n8891)
         );
  NOR2_X1 U10205 ( .A1(n8891), .A2(n9920), .ZN(n8933) );
  INV_X1 U10206 ( .A(n8892), .ZN(n8969) );
  NAND2_X1 U10207 ( .A1(n8894), .A2(n8893), .ZN(n9085) );
  NAND2_X1 U10208 ( .A1(n8896), .A2(n8895), .ZN(n9148) );
  INV_X1 U10209 ( .A(n9209), .ZN(n9205) );
  AND2_X1 U10210 ( .A1(n6454), .A2(n8900), .ZN(n8938) );
  NOR2_X1 U10211 ( .A1(n8901), .A2(n8938), .ZN(n9924) );
  INV_X1 U10212 ( .A(n8902), .ZN(n8905) );
  NAND4_X1 U10213 ( .A1(n9924), .A2(n8905), .A3(n8904), .A4(n8903), .ZN(n8907)
         );
  NOR4_X1 U10214 ( .A1(n8907), .A2(n5557), .A3(n8906), .A4(n5556), .ZN(n8910)
         );
  NAND3_X1 U10215 ( .A1(n8910), .A2(n8909), .A3(n5071), .ZN(n8915) );
  NAND2_X1 U10216 ( .A1(n8912), .A2(n8911), .ZN(n9885) );
  NOR4_X1 U10217 ( .A1(n8915), .A2(n8914), .A3(n8913), .A4(n9885), .ZN(n8916)
         );
  NAND4_X1 U10218 ( .A1(n9258), .A2(n8917), .A3(n8916), .A4(n9726), .ZN(n8919)
         );
  NOR4_X1 U10219 ( .A1(n9227), .A2(n8920), .A3(n8919), .A4(n8918), .ZN(n8921)
         );
  NAND4_X1 U10220 ( .A1(n9175), .A2(n9205), .A3(n4431), .A4(n8921), .ZN(n8922)
         );
  NOR4_X1 U10221 ( .A1(n9136), .A2(n9164), .A3(n9148), .A4(n8922), .ZN(n8923)
         );
  NAND4_X1 U10222 ( .A1(n9085), .A2(n4451), .A3(n8923), .A4(n9116), .ZN(n8924)
         );
  NOR4_X1 U10223 ( .A1(n8969), .A2(n9077), .A3(n8925), .A4(n8924), .ZN(n8928)
         );
  INV_X1 U10224 ( .A(n8926), .ZN(n8971) );
  NAND3_X1 U10225 ( .A1(n8928), .A2(n8927), .A3(n8971), .ZN(n8931) );
  INV_X1 U10226 ( .A(n8929), .ZN(n8930) );
  OAI21_X1 U10227 ( .B1(n9373), .B2(n8983), .A(n8930), .ZN(n8972) );
  OAI21_X1 U10228 ( .B1(n8931), .B2(n8972), .A(n5503), .ZN(n8932) );
  MUX2_X1 U10229 ( .A(n9920), .B(n8933), .S(n8932), .Z(n8934) );
  INV_X1 U10230 ( .A(n8935), .ZN(n8968) );
  INV_X1 U10231 ( .A(n8936), .ZN(n8957) );
  INV_X1 U10232 ( .A(n8937), .ZN(n8954) );
  AOI211_X1 U10233 ( .C1(n8939), .C2(n9926), .A(n5503), .B(n8938), .ZN(n8942)
         );
  OAI22_X1 U10234 ( .A1(n8942), .A2(n8941), .B1(n8940), .B2(n6879), .ZN(n8945)
         );
  NAND3_X1 U10235 ( .A1(n8945), .A2(n8944), .A3(n8943), .ZN(n8953) );
  INV_X1 U10236 ( .A(n8946), .ZN(n8950) );
  INV_X1 U10237 ( .A(n8947), .ZN(n8948) );
  AOI21_X1 U10238 ( .B1(n8950), .B2(n8949), .A(n8948), .ZN(n8952) );
  AOI211_X1 U10239 ( .C1(n8954), .C2(n8953), .A(n8952), .B(n8951), .ZN(n8956)
         );
  OAI21_X1 U10240 ( .B1(n8957), .B2(n8956), .A(n8955), .ZN(n8961) );
  INV_X1 U10241 ( .A(n8958), .ZN(n8960) );
  AOI21_X1 U10242 ( .B1(n8961), .B2(n8960), .A(n8959), .ZN(n8964) );
  OAI21_X1 U10243 ( .B1(n8964), .B2(n8963), .A(n8962), .ZN(n8967) );
  INV_X1 U10244 ( .A(n8965), .ZN(n8966) );
  AOI21_X1 U10245 ( .B1(n8968), .B2(n8967), .A(n8966), .ZN(n8970) );
  NOR2_X1 U10246 ( .A1(n8970), .A2(n8969), .ZN(n8973) );
  OAI21_X1 U10247 ( .B1(n8973), .B2(n8972), .A(n8971), .ZN(n8974) );
  XNOR2_X1 U10248 ( .A(n8974), .B(n9911), .ZN(n8975) );
  NAND2_X1 U10249 ( .A1(n8975), .A2(n9921), .ZN(n8976) );
  NOR3_X1 U10250 ( .A1(n8978), .A2(n4317), .A3(n8977), .ZN(n8981) );
  OAI21_X1 U10251 ( .B1(n8979), .B2(n8982), .A(P1_B_REG_SCAN_IN), .ZN(n8980)
         );
  MUX2_X1 U10252 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n8983), .S(n4315), .Z(
        P1_U3585) );
  MUX2_X1 U10253 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n8984), .S(n4315), .Z(
        P1_U3584) );
  MUX2_X1 U10254 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9079), .S(n4315), .Z(
        P1_U3583) );
  MUX2_X1 U10255 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n8985), .S(n4315), .Z(
        P1_U3582) );
  MUX2_X1 U10256 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9080), .S(n4315), .Z(
        P1_U3581) );
  MUX2_X1 U10257 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9117), .S(P1_U4006), .Z(
        P1_U3580) );
  MUX2_X1 U10258 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n8986), .S(P1_U4006), .Z(
        P1_U3579) );
  MUX2_X1 U10259 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9118), .S(P1_U4006), .Z(
        P1_U3578) );
  MUX2_X1 U10260 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n8987), .S(P1_U4006), .Z(
        P1_U3577) );
  MUX2_X1 U10261 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n8988), .S(n4315), .Z(
        P1_U3576) );
  MUX2_X1 U10262 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n8989), .S(n4315), .Z(
        P1_U3575) );
  MUX2_X1 U10263 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9212), .S(n4315), .Z(
        P1_U3574) );
  MUX2_X1 U10264 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n8990), .S(n4315), .Z(
        P1_U3573) );
  MUX2_X1 U10265 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9213), .S(n4315), .Z(
        P1_U3572) );
  MUX2_X1 U10266 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9706), .S(n4315), .Z(
        P1_U3571) );
  MUX2_X1 U10267 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n8991), .S(n4315), .Z(
        P1_U3570) );
  MUX2_X1 U10268 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n8992), .S(n4315), .Z(
        P1_U3569) );
  MUX2_X1 U10269 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n8993), .S(n4315), .Z(
        P1_U3568) );
  MUX2_X1 U10270 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9728), .S(n4315), .Z(
        P1_U3567) );
  MUX2_X1 U10271 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n8994), .S(n4315), .Z(
        P1_U3566) );
  MUX2_X1 U10272 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9729), .S(n4315), .Z(
        P1_U3565) );
  MUX2_X1 U10273 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n8995), .S(n4315), .Z(
        P1_U3564) );
  MUX2_X1 U10274 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n8996), .S(n4315), .Z(
        P1_U3563) );
  MUX2_X1 U10275 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n8997), .S(n4315), .Z(
        P1_U3562) );
  MUX2_X1 U10276 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n8998), .S(n4315), .Z(
        P1_U3561) );
  MUX2_X1 U10277 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n8999), .S(n4315), .Z(
        P1_U3560) );
  MUX2_X1 U10278 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9000), .S(n4315), .Z(
        P1_U3559) );
  MUX2_X1 U10279 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9001), .S(n4315), .Z(
        P1_U3558) );
  MUX2_X1 U10280 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n9002), .S(n4315), .Z(
        P1_U3557) );
  MUX2_X1 U10281 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n9926), .S(n4315), .Z(
        P1_U3556) );
  NOR2_X1 U10282 ( .A1(n9003), .A2(n9009), .ZN(n9005) );
  NAND2_X1 U10283 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n9028), .ZN(n9006) );
  OAI21_X1 U10284 ( .B1(n9028), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9006), .ZN(
        n9007) );
  AOI211_X1 U10285 ( .C1(n4397), .C2(n9007), .A(n9024), .B(n9847), .ZN(n9019)
         );
  NOR2_X1 U10286 ( .A1(n9009), .A2(n9008), .ZN(n9011) );
  XNOR2_X1 U10287 ( .A(n9028), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n9012) );
  NOR2_X1 U10288 ( .A1(n9013), .A2(n9012), .ZN(n9027) );
  AOI211_X1 U10289 ( .C1(n9013), .C2(n9012), .A(n9027), .B(n9797), .ZN(n9018)
         );
  INV_X1 U10290 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n9016) );
  NAND2_X1 U10291 ( .A1(P1_REG3_REG_16__SCAN_IN), .A2(P1_U3084), .ZN(n9015) );
  NAND2_X1 U10292 ( .A1(n9860), .A2(n9028), .ZN(n9014) );
  OAI211_X1 U10293 ( .C1(n9873), .C2(n9016), .A(n9015), .B(n9014), .ZN(n9017)
         );
  OR3_X1 U10294 ( .A1(n9019), .A2(n9018), .A3(n9017), .ZN(P1_U3257) );
  INV_X1 U10295 ( .A(n9039), .ZN(n9022) );
  NAND2_X1 U10296 ( .A1(n9854), .A2(P1_ADDR_REG_17__SCAN_IN), .ZN(n9021) );
  NAND2_X1 U10297 ( .A1(P1_REG3_REG_17__SCAN_IN), .A2(P1_U3084), .ZN(n9020) );
  OAI211_X1 U10298 ( .C1(n9023), .C2(n9022), .A(n9021), .B(n9020), .ZN(n9033)
         );
  AOI21_X1 U10299 ( .B1(n9028), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9024), .ZN(
        n9026) );
  XNOR2_X1 U10300 ( .A(n9039), .B(P1_REG2_REG_17__SCAN_IN), .ZN(n9025) );
  AOI211_X1 U10301 ( .C1(n9026), .C2(n9025), .A(n9034), .B(n9847), .ZN(n9032)
         );
  XNOR2_X1 U10302 ( .A(n9039), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9030) );
  AOI21_X1 U10303 ( .B1(n9028), .B2(P1_REG1_REG_16__SCAN_IN), .A(n9027), .ZN(
        n9029) );
  NOR2_X1 U10304 ( .A1(n9029), .A2(n9030), .ZN(n9038) );
  AOI211_X1 U10305 ( .C1(n9030), .C2(n9029), .A(n9038), .B(n9797), .ZN(n9031)
         );
  OR3_X1 U10306 ( .A1(n9033), .A2(n9032), .A3(n9031), .ZN(P1_U3258) );
  INV_X1 U10307 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n9047) );
  NAND2_X1 U10308 ( .A1(n9859), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9035) );
  OAI21_X1 U10309 ( .B1(n9859), .B2(P1_REG2_REG_18__SCAN_IN), .A(n9035), .ZN(
        n9862) );
  XNOR2_X1 U10310 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n9036), .ZN(n9045) );
  INV_X1 U10311 ( .A(n9045), .ZN(n9041) );
  INV_X1 U10312 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9347) );
  AOI22_X1 U10313 ( .A1(n9859), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n9347), .B2(
        n9037), .ZN(n9866) );
  NAND2_X1 U10314 ( .A1(n9866), .A2(n9865), .ZN(n9864) );
  OAI21_X1 U10315 ( .B1(n9859), .B2(P1_REG1_REG_18__SCAN_IN), .A(n9864), .ZN(
        n9040) );
  XOR2_X1 U10316 ( .A(n9040), .B(P1_REG1_REG_19__SCAN_IN), .Z(n9042) );
  AOI21_X1 U10317 ( .B1(n9042), .B2(n9868), .A(n9860), .ZN(n9043) );
  INV_X1 U10318 ( .A(n8803), .ZN(n9369) );
  XNOR2_X1 U10319 ( .A(n4325), .B(n8803), .ZN(n9048) );
  NAND2_X1 U10320 ( .A1(n9286), .A2(n9881), .ZN(n9052) );
  AND2_X1 U10321 ( .A1(n9050), .A2(n9049), .ZN(n9285) );
  INV_X1 U10322 ( .A(n9285), .ZN(n9289) );
  NOR2_X1 U10323 ( .A1(n9289), .A2(n9938), .ZN(n9057) );
  AOI21_X1 U10324 ( .B1(n9938), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9057), .ZN(
        n9051) );
  OAI211_X1 U10325 ( .C1(n9369), .C2(n9899), .A(n9052), .B(n9051), .ZN(
        P1_U3261) );
  XNOR2_X1 U10326 ( .A(n9054), .B(n9053), .ZN(n9055) );
  NAND2_X1 U10327 ( .A1(n9055), .A2(n9877), .ZN(n9290) );
  NOR2_X1 U10328 ( .A1(n9373), .A2(n9899), .ZN(n9056) );
  AOI211_X1 U10329 ( .C1(n9938), .C2(P1_REG2_REG_30__SCAN_IN), .A(n9057), .B(
        n9056), .ZN(n9058) );
  OAI21_X1 U10330 ( .B1(n9059), .B2(n9290), .A(n9058), .ZN(P1_U3262) );
  INV_X1 U10331 ( .A(n9060), .ZN(n9065) );
  NAND2_X1 U10332 ( .A1(n9061), .A2(n9233), .ZN(n9064) );
  AOI22_X1 U10333 ( .A1(n9062), .A2(n9896), .B1(P1_REG2_REG_28__SCAN_IN), .B2(
        n9938), .ZN(n9063) );
  OAI211_X1 U10334 ( .C1(n9065), .C2(n9899), .A(n9064), .B(n9063), .ZN(n9066)
         );
  AOI21_X1 U10335 ( .B1(n9067), .B2(n9918), .A(n9066), .ZN(n9068) );
  OAI21_X1 U10336 ( .B1(n9069), .B2(n9253), .A(n9068), .ZN(P1_U3263) );
  XNOR2_X1 U10337 ( .A(n9071), .B(n9070), .ZN(n9302) );
  INV_X1 U10338 ( .A(n9072), .ZN(n9073) );
  AOI211_X1 U10339 ( .C1(n9299), .C2(n9089), .A(n9263), .B(n9073), .ZN(n9298)
         );
  INV_X1 U10340 ( .A(n9299), .ZN(n9076) );
  AOI22_X1 U10341 ( .A1(n9074), .A2(n9896), .B1(P1_REG2_REG_27__SCAN_IN), .B2(
        n9938), .ZN(n9075) );
  OAI21_X1 U10342 ( .B1(n9076), .B2(n9899), .A(n9075), .ZN(n9081) );
  OAI21_X1 U10343 ( .B1(n9302), .B2(n9253), .A(n9082), .ZN(P1_U3264) );
  XOR2_X1 U10344 ( .A(n9085), .B(n9083), .Z(n9305) );
  INV_X1 U10345 ( .A(n9305), .ZN(n9098) );
  XOR2_X1 U10346 ( .A(n9085), .B(n9084), .Z(n9086) );
  OAI222_X1 U10347 ( .A1(n9889), .A2(n9088), .B1(n9887), .B2(n9087), .C1(n9086), .C2(n9732), .ZN(n9303) );
  INV_X1 U10348 ( .A(n9100), .ZN(n9091) );
  INV_X1 U10349 ( .A(n9089), .ZN(n9090) );
  AOI211_X1 U10350 ( .C1(n9092), .C2(n9091), .A(n9263), .B(n9090), .ZN(n9304)
         );
  NAND2_X1 U10351 ( .A1(n9304), .A2(n9881), .ZN(n9095) );
  AOI22_X1 U10352 ( .A1(n9093), .A2(n9896), .B1(P1_REG2_REG_26__SCAN_IN), .B2(
        n9938), .ZN(n9094) );
  OAI211_X1 U10353 ( .C1(n9379), .C2(n9899), .A(n9095), .B(n9094), .ZN(n9096)
         );
  AOI21_X1 U10354 ( .B1(n9303), .B2(n9918), .A(n9096), .ZN(n9097) );
  OAI21_X1 U10355 ( .B1(n9098), .B2(n9253), .A(n9097), .ZN(P1_U3265) );
  XOR2_X1 U10356 ( .A(n9099), .B(n9108), .Z(n9312) );
  INV_X1 U10357 ( .A(n9123), .ZN(n9101) );
  AOI211_X1 U10358 ( .C1(n9310), .C2(n9101), .A(n9263), .B(n9100), .ZN(n9309)
         );
  NOR2_X1 U10359 ( .A1(n9102), .A2(n9899), .ZN(n9106) );
  OAI22_X1 U10360 ( .A1(n9104), .A2(n9272), .B1(n9103), .B2(n9918), .ZN(n9105)
         );
  AOI211_X1 U10361 ( .C1(n9309), .C2(n9233), .A(n9106), .B(n9105), .ZN(n9112)
         );
  NAND2_X1 U10362 ( .A1(n9115), .A2(n9107), .ZN(n9109) );
  NAND2_X1 U10363 ( .A1(n9308), .A2(n9918), .ZN(n9111) );
  OAI211_X1 U10364 ( .C1(n9312), .C2(n9253), .A(n9112), .B(n9111), .ZN(
        P1_U3266) );
  XNOR2_X1 U10365 ( .A(n9113), .B(n9116), .ZN(n9315) );
  INV_X1 U10366 ( .A(n9120), .ZN(n9384) );
  OAI22_X1 U10367 ( .A1(n9384), .A2(n9899), .B1(n9114), .B2(n9918), .ZN(n9127)
         );
  OAI21_X1 U10368 ( .B1(n4357), .B2(n9116), .A(n9115), .ZN(n9119) );
  AOI222_X1 U10369 ( .A1(n9892), .A2(n9119), .B1(n9118), .B2(n9730), .C1(n9117), .C2(n9925), .ZN(n9313) );
  NAND2_X1 U10370 ( .A1(n9130), .A2(n9120), .ZN(n9121) );
  NAND2_X1 U10371 ( .A1(n9121), .A2(n9877), .ZN(n9122) );
  NOR2_X1 U10372 ( .A1(n9123), .A2(n9122), .ZN(n9314) );
  AOI22_X1 U10373 ( .A1(n9314), .A2(n9911), .B1(n9896), .B2(n9124), .ZN(n9125)
         );
  AOI21_X1 U10374 ( .B1(n9313), .B2(n9125), .A(n9938), .ZN(n9126) );
  AOI211_X1 U10375 ( .C1(n9277), .C2(n9315), .A(n9127), .B(n9126), .ZN(n9128)
         );
  INV_X1 U10376 ( .A(n9128), .ZN(P1_U3267) );
  XNOR2_X1 U10377 ( .A(n9129), .B(n4685), .ZN(n9322) );
  INV_X1 U10378 ( .A(n9130), .ZN(n9131) );
  AOI211_X1 U10379 ( .C1(n9319), .C2(n9149), .A(n9263), .B(n9131), .ZN(n9318)
         );
  INV_X1 U10380 ( .A(n9319), .ZN(n9135) );
  INV_X1 U10381 ( .A(n9132), .ZN(n9133) );
  AOI22_X1 U10382 ( .A1(n9133), .A2(n9896), .B1(n9938), .B2(
        P1_REG2_REG_23__SCAN_IN), .ZN(n9134) );
  OAI21_X1 U10383 ( .B1(n9135), .B2(n9899), .A(n9134), .ZN(n9142) );
  AOI21_X1 U10384 ( .B1(n9137), .B2(n9136), .A(n9732), .ZN(n9140) );
  OAI22_X1 U10385 ( .A1(n9138), .A2(n9887), .B1(n9166), .B2(n9889), .ZN(n9139)
         );
  AOI21_X1 U10386 ( .B1(n9140), .B2(n4687), .A(n9139), .ZN(n9321) );
  NOR2_X1 U10387 ( .A1(n9321), .A2(n9938), .ZN(n9141) );
  AOI211_X1 U10388 ( .C1(n9318), .C2(n9233), .A(n9142), .B(n9141), .ZN(n9143)
         );
  OAI21_X1 U10389 ( .B1(n9322), .B2(n9253), .A(n9143), .ZN(P1_U3268) );
  XNOR2_X1 U10390 ( .A(n9144), .B(n9148), .ZN(n9145) );
  OAI222_X1 U10391 ( .A1(n9887), .A2(n9146), .B1(n9889), .B2(n9178), .C1(n9145), .C2(n9732), .ZN(n9323) );
  INV_X1 U10392 ( .A(n9323), .ZN(n9159) );
  XOR2_X1 U10393 ( .A(n9148), .B(n9147), .Z(n9325) );
  NAND2_X1 U10394 ( .A1(n9325), .A2(n9277), .ZN(n9158) );
  INV_X1 U10395 ( .A(n9167), .ZN(n9151) );
  INV_X1 U10396 ( .A(n9149), .ZN(n9150) );
  AOI211_X1 U10397 ( .C1(n9152), .C2(n9151), .A(n9263), .B(n9150), .ZN(n9324)
         );
  NOR2_X1 U10398 ( .A1(n9389), .A2(n9899), .ZN(n9156) );
  OAI22_X1 U10399 ( .A1(n9154), .A2(n9918), .B1(n9153), .B2(n9272), .ZN(n9155)
         );
  AOI211_X1 U10400 ( .C1(n9324), .C2(n9881), .A(n9156), .B(n9155), .ZN(n9157)
         );
  OAI211_X1 U10401 ( .C1(n9938), .C2(n9159), .A(n9158), .B(n9157), .ZN(
        P1_U3269) );
  XOR2_X1 U10402 ( .A(n9160), .B(n9164), .Z(n9331) );
  INV_X1 U10403 ( .A(n9331), .ZN(n9173) );
  AOI22_X1 U10404 ( .A1(n9328), .A2(n9737), .B1(P1_REG2_REG_21__SCAN_IN), .B2(
        n9938), .ZN(n9172) );
  INV_X1 U10405 ( .A(n9161), .ZN(n9162) );
  AOI21_X1 U10406 ( .B1(n9164), .B2(n9163), .A(n9162), .ZN(n9165) );
  OAI222_X1 U10407 ( .A1(n9889), .A2(n9197), .B1(n9887), .B2(n9166), .C1(n9732), .C2(n9165), .ZN(n9329) );
  AOI211_X1 U10408 ( .C1(n9328), .C2(n9181), .A(n9263), .B(n9167), .ZN(n9330)
         );
  INV_X1 U10409 ( .A(n9330), .ZN(n9169) );
  OAI22_X1 U10410 ( .A1(n9169), .A2(n9920), .B1(n9272), .B2(n9168), .ZN(n9170)
         );
  OAI21_X1 U10411 ( .B1(n9329), .B2(n9170), .A(n9918), .ZN(n9171) );
  OAI211_X1 U10412 ( .C1(n9173), .C2(n9253), .A(n9172), .B(n9171), .ZN(
        P1_U3270) );
  XOR2_X1 U10413 ( .A(n9174), .B(n9175), .Z(n9336) );
  INV_X1 U10414 ( .A(n9336), .ZN(n9190) );
  XOR2_X1 U10415 ( .A(n9176), .B(n9175), .Z(n9177) );
  OAI222_X1 U10416 ( .A1(n9889), .A2(n9179), .B1(n9887), .B2(n9178), .C1(n9177), .C2(n9732), .ZN(n9334) );
  INV_X1 U10417 ( .A(n9181), .ZN(n9182) );
  AOI211_X1 U10418 ( .C1(n9183), .C2(n4632), .A(n9263), .B(n9182), .ZN(n9335)
         );
  NAND2_X1 U10419 ( .A1(n9335), .A2(n9233), .ZN(n9187) );
  INV_X1 U10420 ( .A(n9184), .ZN(n9185) );
  AOI22_X1 U10421 ( .A1(n9938), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9185), .B2(
        n9896), .ZN(n9186) );
  OAI211_X1 U10422 ( .C1(n5548), .C2(n9899), .A(n9187), .B(n9186), .ZN(n9188)
         );
  AOI21_X1 U10423 ( .B1(n9334), .B2(n9918), .A(n9188), .ZN(n9189) );
  OAI21_X1 U10424 ( .B1(n9190), .B2(n9253), .A(n9189), .ZN(P1_U3271) );
  XNOR2_X1 U10425 ( .A(n9191), .B(n9194), .ZN(n9343) );
  INV_X1 U10426 ( .A(n9192), .ZN(n9193) );
  AOI21_X1 U10427 ( .B1(n9195), .B2(n9194), .A(n9193), .ZN(n9196) );
  OAI222_X1 U10428 ( .A1(n9889), .A2(n9230), .B1(n9887), .B2(n9197), .C1(n9732), .C2(n9196), .ZN(n9339) );
  INV_X1 U10429 ( .A(n9341), .ZN(n9201) );
  AOI211_X1 U10430 ( .C1(n9341), .C2(n9216), .A(n9263), .B(n9180), .ZN(n9340)
         );
  NAND2_X1 U10431 ( .A1(n9340), .A2(n9233), .ZN(n9200) );
  AOI22_X1 U10432 ( .A1(n9938), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9198), .B2(
        n9896), .ZN(n9199) );
  OAI211_X1 U10433 ( .C1(n9201), .C2(n9899), .A(n9200), .B(n9199), .ZN(n9202)
         );
  AOI21_X1 U10434 ( .B1(n9339), .B2(n9918), .A(n9202), .ZN(n9203) );
  OAI21_X1 U10435 ( .B1(n9253), .B2(n9343), .A(n9203), .ZN(P1_U3272) );
  XNOR2_X1 U10436 ( .A(n9204), .B(n9205), .ZN(n9346) );
  INV_X1 U10437 ( .A(n9346), .ZN(n9225) );
  INV_X1 U10438 ( .A(n9206), .ZN(n9208) );
  OAI21_X1 U10439 ( .B1(n9228), .B2(n9208), .A(n9207), .ZN(n9210) );
  XNOR2_X1 U10440 ( .A(n9210), .B(n9209), .ZN(n9211) );
  NAND2_X1 U10441 ( .A1(n9211), .A2(n9892), .ZN(n9215) );
  AOI22_X1 U10442 ( .A1(n9730), .A2(n9213), .B1(n9212), .B2(n9925), .ZN(n9214)
         );
  NAND2_X1 U10443 ( .A1(n9215), .A2(n9214), .ZN(n9344) );
  INV_X1 U10444 ( .A(n9231), .ZN(n9218) );
  INV_X1 U10445 ( .A(n9216), .ZN(n9217) );
  AOI211_X1 U10446 ( .C1(n9219), .C2(n9218), .A(n9263), .B(n9217), .ZN(n9345)
         );
  NAND2_X1 U10447 ( .A1(n9345), .A2(n9881), .ZN(n9222) );
  AOI22_X1 U10448 ( .A1(n9938), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9220), .B2(
        n9896), .ZN(n9221) );
  OAI211_X1 U10449 ( .C1(n9400), .C2(n9899), .A(n9222), .B(n9221), .ZN(n9223)
         );
  AOI21_X1 U10450 ( .B1(n9344), .B2(n9918), .A(n9223), .ZN(n9224) );
  OAI21_X1 U10451 ( .B1(n9225), .B2(n9253), .A(n9224), .ZN(P1_U3273) );
  XNOR2_X1 U10452 ( .A(n9226), .B(n9227), .ZN(n9353) );
  XNOR2_X1 U10453 ( .A(n9228), .B(n9227), .ZN(n9229) );
  OAI222_X1 U10454 ( .A1(n9887), .A2(n9230), .B1(n9889), .B2(n9256), .C1(n9229), .C2(n9732), .ZN(n9349) );
  INV_X1 U10455 ( .A(n9246), .ZN(n9232) );
  AOI211_X1 U10456 ( .C1(n9351), .C2(n9232), .A(n9263), .B(n9231), .ZN(n9350)
         );
  NAND2_X1 U10457 ( .A1(n9350), .A2(n9233), .ZN(n9236) );
  AOI22_X1 U10458 ( .A1(n9938), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9234), .B2(
        n9896), .ZN(n9235) );
  OAI211_X1 U10459 ( .C1(n9237), .C2(n9899), .A(n9236), .B(n9235), .ZN(n9238)
         );
  AOI21_X1 U10460 ( .B1(n9349), .B2(n9918), .A(n9238), .ZN(n9239) );
  OAI21_X1 U10461 ( .B1(n9353), .B2(n9253), .A(n9239), .ZN(P1_U3274) );
  XNOR2_X1 U10462 ( .A(n9240), .B(n9241), .ZN(n9357) );
  INV_X1 U10463 ( .A(n9357), .ZN(n9254) );
  XNOR2_X1 U10464 ( .A(n9242), .B(n9241), .ZN(n9243) );
  OAI222_X1 U10465 ( .A1(n9889), .A2(n9245), .B1(n9887), .B2(n9244), .C1(n9732), .C2(n9243), .ZN(n9355) );
  INV_X1 U10466 ( .A(n9247), .ZN(n9406) );
  AOI211_X1 U10467 ( .C1(n9247), .C2(n9262), .A(n9263), .B(n9246), .ZN(n9356)
         );
  NAND2_X1 U10468 ( .A1(n9356), .A2(n9881), .ZN(n9250) );
  AOI22_X1 U10469 ( .A1(n9938), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9248), .B2(
        n9896), .ZN(n9249) );
  OAI211_X1 U10470 ( .C1(n9406), .C2(n9899), .A(n9250), .B(n9249), .ZN(n9251)
         );
  AOI21_X1 U10471 ( .B1(n9355), .B2(n9918), .A(n9251), .ZN(n9252) );
  OAI21_X1 U10472 ( .B1(n9254), .B2(n9253), .A(n9252), .ZN(P1_U3275) );
  XOR2_X1 U10473 ( .A(n9255), .B(n9258), .Z(n9261) );
  OAI22_X1 U10474 ( .A1(n9710), .A2(n9889), .B1(n9256), .B2(n9887), .ZN(n9260)
         );
  XNOR2_X1 U10475 ( .A(n9257), .B(n9258), .ZN(n9364) );
  NOR2_X1 U10476 ( .A1(n9364), .A2(n9946), .ZN(n9259) );
  AOI211_X1 U10477 ( .C1(n9892), .C2(n9261), .A(n9260), .B(n9259), .ZN(n9363)
         );
  AOI211_X1 U10478 ( .C1(n9712), .C2(n4336), .A(n9263), .B(n4634), .ZN(n9361)
         );
  INV_X1 U10479 ( .A(n9712), .ZN(n9266) );
  AOI22_X1 U10480 ( .A1(n9938), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n9264), .B2(
        n9896), .ZN(n9265) );
  OAI21_X1 U10481 ( .B1(n9266), .B2(n9899), .A(n9265), .ZN(n9269) );
  NOR2_X1 U10482 ( .A1(n9364), .A2(n9267), .ZN(n9268) );
  AOI211_X1 U10483 ( .C1(n9361), .C2(n9881), .A(n9269), .B(n9268), .ZN(n9270)
         );
  OAI21_X1 U10484 ( .B1(n9363), .B2(n9938), .A(n9270), .ZN(P1_U3276) );
  NAND2_X1 U10485 ( .A1(n9271), .A2(n9918), .ZN(n9283) );
  OAI22_X1 U10486 ( .A1(n9918), .A2(n9274), .B1(n9273), .B2(n9272), .ZN(n9275)
         );
  AOI21_X1 U10487 ( .B1(n9737), .B2(n9276), .A(n9275), .ZN(n9282) );
  NAND2_X1 U10488 ( .A1(n9278), .A2(n9277), .ZN(n9281) );
  NAND2_X1 U10489 ( .A1(n9279), .A2(n9881), .ZN(n9280) );
  NAND4_X1 U10490 ( .A1(n9283), .A2(n9282), .A3(n9281), .A4(n9280), .ZN(
        P1_U3285) );
  INV_X1 U10491 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9287) );
  NOR2_X1 U10492 ( .A1(n9286), .A2(n9285), .ZN(n9366) );
  MUX2_X1 U10493 ( .A(n9287), .B(n9366), .S(n9978), .Z(n9288) );
  OAI21_X1 U10494 ( .B1(n9369), .B2(n9360), .A(n9288), .ZN(P1_U3554) );
  INV_X1 U10495 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9291) );
  MUX2_X1 U10496 ( .A(n9291), .B(n9371), .S(n9978), .Z(n9292) );
  OAI21_X1 U10497 ( .B1(n9373), .B2(n9360), .A(n9292), .ZN(P1_U3553) );
  AOI21_X1 U10498 ( .B1(n9942), .B2(n9294), .A(n9293), .ZN(n9295) );
  OAI211_X1 U10499 ( .C1(n9297), .C2(n9354), .A(n9296), .B(n9295), .ZN(n9374)
         );
  MUX2_X1 U10500 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9374), .S(n9978), .Z(
        P1_U3552) );
  AOI21_X1 U10501 ( .B1(n9942), .B2(n9299), .A(n9298), .ZN(n9300) );
  OAI211_X1 U10502 ( .C1(n9302), .C2(n9354), .A(n9301), .B(n9300), .ZN(n9375)
         );
  MUX2_X1 U10503 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9375), .S(n9978), .Z(
        P1_U3550) );
  INV_X1 U10504 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n9306) );
  AOI211_X1 U10505 ( .C1(n9305), .C2(n9957), .A(n9304), .B(n9303), .ZN(n9376)
         );
  MUX2_X1 U10506 ( .A(n9306), .B(n9376), .S(n9978), .Z(n9307) );
  OAI21_X1 U10507 ( .B1(n9379), .B2(n9360), .A(n9307), .ZN(P1_U3549) );
  AOI211_X1 U10508 ( .C1(n9942), .C2(n9310), .A(n9309), .B(n9308), .ZN(n9311)
         );
  OAI21_X1 U10509 ( .B1(n9312), .B2(n9354), .A(n9311), .ZN(n9380) );
  MUX2_X1 U10510 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9380), .S(n9978), .Z(
        P1_U3548) );
  INV_X1 U10511 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n9316) );
  MUX2_X1 U10512 ( .A(n9316), .B(n9381), .S(n9978), .Z(n9317) );
  OAI21_X1 U10513 ( .B1(n9384), .B2(n9360), .A(n9317), .ZN(P1_U3547) );
  AOI21_X1 U10514 ( .B1(n9942), .B2(n9319), .A(n9318), .ZN(n9320) );
  OAI211_X1 U10515 ( .C1(n9322), .C2(n9354), .A(n9321), .B(n9320), .ZN(n9385)
         );
  MUX2_X1 U10516 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9385), .S(n9978), .Z(
        P1_U3546) );
  INV_X1 U10517 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n9326) );
  AOI211_X1 U10518 ( .C1(n9325), .C2(n9957), .A(n9324), .B(n9323), .ZN(n9386)
         );
  MUX2_X1 U10519 ( .A(n9326), .B(n9386), .S(n9978), .Z(n9327) );
  OAI21_X1 U10520 ( .B1(n9389), .B2(n9360), .A(n9327), .ZN(P1_U3545) );
  INV_X1 U10521 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n9332) );
  AOI211_X1 U10522 ( .C1(n9331), .C2(n9957), .A(n9330), .B(n9329), .ZN(n9390)
         );
  MUX2_X1 U10523 ( .A(n9332), .B(n9390), .S(n9978), .Z(n9333) );
  OAI21_X1 U10524 ( .B1(n4628), .B2(n9360), .A(n9333), .ZN(P1_U3544) );
  INV_X1 U10525 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n9337) );
  AOI211_X1 U10526 ( .C1(n9336), .C2(n9957), .A(n9335), .B(n9334), .ZN(n9393)
         );
  MUX2_X1 U10527 ( .A(n9337), .B(n9393), .S(n9978), .Z(n9338) );
  OAI21_X1 U10528 ( .B1(n5548), .B2(n9360), .A(n9338), .ZN(P1_U3543) );
  AOI211_X1 U10529 ( .C1(n9942), .C2(n9341), .A(n9340), .B(n9339), .ZN(n9342)
         );
  OAI21_X1 U10530 ( .B1(n9354), .B2(n9343), .A(n9342), .ZN(n9396) );
  MUX2_X1 U10531 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9396), .S(n9978), .Z(
        P1_U3542) );
  AOI211_X1 U10532 ( .C1(n9346), .C2(n9957), .A(n9345), .B(n9344), .ZN(n9397)
         );
  MUX2_X1 U10533 ( .A(n9347), .B(n9397), .S(n9978), .Z(n9348) );
  OAI21_X1 U10534 ( .B1(n9400), .B2(n9360), .A(n9348), .ZN(P1_U3541) );
  AOI211_X1 U10535 ( .C1(n9942), .C2(n9351), .A(n9350), .B(n9349), .ZN(n9352)
         );
  OAI21_X1 U10536 ( .B1(n9354), .B2(n9353), .A(n9352), .ZN(n9401) );
  MUX2_X1 U10537 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9401), .S(n9978), .Z(
        P1_U3540) );
  INV_X1 U10538 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9358) );
  AOI211_X1 U10539 ( .C1(n9357), .C2(n9957), .A(n9356), .B(n9355), .ZN(n9402)
         );
  MUX2_X1 U10540 ( .A(n9358), .B(n9402), .S(n9978), .Z(n9359) );
  OAI21_X1 U10541 ( .B1(n9406), .B2(n9360), .A(n9359), .ZN(P1_U3539) );
  AOI21_X1 U10542 ( .B1(n9942), .B2(n9712), .A(n9361), .ZN(n9362) );
  OAI211_X1 U10543 ( .C1(n9364), .C2(n9945), .A(n9363), .B(n9362), .ZN(n9407)
         );
  MUX2_X1 U10544 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9407), .S(n9978), .Z(
        P1_U3538) );
  INV_X1 U10545 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n9367) );
  MUX2_X1 U10546 ( .A(n9367), .B(n9366), .S(n9968), .Z(n9368) );
  OAI21_X1 U10547 ( .B1(n9369), .B2(n9405), .A(n9368), .ZN(P1_U3522) );
  INV_X1 U10548 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9370) );
  MUX2_X1 U10549 ( .A(n9371), .B(n9370), .S(n9966), .Z(n9372) );
  OAI21_X1 U10550 ( .B1(n9373), .B2(n9405), .A(n9372), .ZN(P1_U3521) );
  MUX2_X1 U10551 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9374), .S(n9968), .Z(
        P1_U3520) );
  MUX2_X1 U10552 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9375), .S(n9968), .Z(
        P1_U3518) );
  INV_X1 U10553 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n9377) );
  MUX2_X1 U10554 ( .A(n9377), .B(n9376), .S(n9968), .Z(n9378) );
  OAI21_X1 U10555 ( .B1(n9379), .B2(n9405), .A(n9378), .ZN(P1_U3517) );
  MUX2_X1 U10556 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9380), .S(n9968), .Z(
        P1_U3516) );
  INV_X1 U10557 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n9382) );
  MUX2_X1 U10558 ( .A(n9382), .B(n9381), .S(n9968), .Z(n9383) );
  OAI21_X1 U10559 ( .B1(n9384), .B2(n9405), .A(n9383), .ZN(P1_U3515) );
  MUX2_X1 U10560 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9385), .S(n9968), .Z(
        P1_U3514) );
  INV_X1 U10561 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n9387) );
  MUX2_X1 U10562 ( .A(n9387), .B(n9386), .S(n9968), .Z(n9388) );
  OAI21_X1 U10563 ( .B1(n9389), .B2(n9405), .A(n9388), .ZN(P1_U3513) );
  INV_X1 U10564 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n9391) );
  MUX2_X1 U10565 ( .A(n9391), .B(n9390), .S(n9968), .Z(n9392) );
  OAI21_X1 U10566 ( .B1(n4628), .B2(n9405), .A(n9392), .ZN(P1_U3512) );
  INV_X1 U10567 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n9394) );
  MUX2_X1 U10568 ( .A(n9394), .B(n9393), .S(n9968), .Z(n9395) );
  OAI21_X1 U10569 ( .B1(n5548), .B2(n9405), .A(n9395), .ZN(P1_U3511) );
  MUX2_X1 U10570 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9396), .S(n9968), .Z(
        P1_U3510) );
  INV_X1 U10571 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n9398) );
  MUX2_X1 U10572 ( .A(n9398), .B(n9397), .S(n9968), .Z(n9399) );
  OAI21_X1 U10573 ( .B1(n9400), .B2(n9405), .A(n9399), .ZN(P1_U3508) );
  MUX2_X1 U10574 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9401), .S(n9968), .Z(
        P1_U3505) );
  INV_X1 U10575 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n9403) );
  MUX2_X1 U10576 ( .A(n9403), .B(n9402), .S(n9968), .Z(n9404) );
  OAI21_X1 U10577 ( .B1(n9406), .B2(n9405), .A(n9404), .ZN(P1_U3502) );
  MUX2_X1 U10578 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n9407), .S(n9968), .Z(
        P1_U3499) );
  MUX2_X1 U10579 ( .A(P1_D_REG_0__SCAN_IN), .B(n9409), .S(n9408), .Z(P1_U3440)
         );
  NOR4_X1 U10580 ( .A1(n9411), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3084), .A4(
        n9410), .ZN(n9412) );
  AOI21_X1 U10581 ( .B1(n9428), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9412), .ZN(
        n9413) );
  OAI21_X1 U10582 ( .B1(n9414), .B2(n9420), .A(n9413), .ZN(P1_U3322) );
  AOI22_X1 U10583 ( .A1(n9415), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n9428), .ZN(n9416) );
  OAI21_X1 U10584 ( .B1(n9417), .B2(n9420), .A(n9416), .ZN(P1_U3323) );
  AOI22_X1 U10585 ( .A1(n9418), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n9428), .ZN(n9419) );
  OAI21_X1 U10586 ( .B1(n9421), .B2(n9420), .A(n9419), .ZN(P1_U3324) );
  NAND2_X1 U10587 ( .A1(n9428), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n9423) );
  OAI211_X1 U10588 ( .C1(n9424), .C2(n9420), .A(n9423), .B(n9422), .ZN(
        P1_U3325) );
  AOI21_X1 U10589 ( .B1(n9428), .B2(P2_DATAO_REG_27__SCAN_IN), .A(n9425), .ZN(
        n9426) );
  OAI21_X1 U10590 ( .B1(n9427), .B2(n9420), .A(n9426), .ZN(P1_U3326) );
  AOI22_X1 U10591 ( .A1(n9429), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n9428), .ZN(n9430) );
  OAI21_X1 U10592 ( .B1(n9431), .B2(n9420), .A(n9430), .ZN(P1_U3327) );
  INV_X1 U10593 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10085) );
  NOR2_X1 U10594 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n9432) );
  AOI21_X1 U10595 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n9432), .ZN(n10055) );
  NOR2_X1 U10596 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n9433) );
  AOI21_X1 U10597 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n9433), .ZN(n10058) );
  NOR2_X1 U10598 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n9434) );
  AOI21_X1 U10599 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n9434), .ZN(n10061) );
  NOR2_X1 U10600 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n9435) );
  AOI21_X1 U10601 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n9435), .ZN(n10064) );
  NOR2_X1 U10602 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n9436) );
  AOI21_X1 U10603 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n9436), .ZN(n10067) );
  NOR2_X1 U10604 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n9442) );
  XNOR2_X1 U10605 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10096) );
  NAND2_X1 U10606 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n9440) );
  XOR2_X1 U10607 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10094) );
  NAND2_X1 U10608 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n9438) );
  XOR2_X1 U10609 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(P1_ADDR_REG_2__SCAN_IN), .Z(
        n10081) );
  AOI21_X1 U10610 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10049) );
  INV_X1 U10611 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n9655) );
  NAND3_X1 U10612 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n10051) );
  OAI21_X1 U10613 ( .B1(n10049), .B2(n9655), .A(n10051), .ZN(n10080) );
  NAND2_X1 U10614 ( .A1(n10081), .A2(n10080), .ZN(n9437) );
  NAND2_X1 U10615 ( .A1(n9438), .A2(n9437), .ZN(n10093) );
  NAND2_X1 U10616 ( .A1(n10094), .A2(n10093), .ZN(n9439) );
  NAND2_X1 U10617 ( .A1(n9440), .A2(n9439), .ZN(n10095) );
  NOR2_X1 U10618 ( .A1(n10096), .A2(n10095), .ZN(n9441) );
  NAND2_X1 U10619 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n10090), .ZN(n9443) );
  NOR2_X1 U10620 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n10090), .ZN(n10089) );
  NAND2_X1 U10621 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(n9444), .ZN(n9446) );
  XOR2_X1 U10622 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(n9444), .Z(n10088) );
  NAND2_X1 U10623 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(n10088), .ZN(n9445) );
  NAND2_X1 U10624 ( .A1(n9446), .A2(n9445), .ZN(n9447) );
  NAND2_X1 U10625 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n9447), .ZN(n9449) );
  XOR2_X1 U10626 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n9447), .Z(n10087) );
  NAND2_X1 U10627 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n10087), .ZN(n9448) );
  NAND2_X1 U10628 ( .A1(n9449), .A2(n9448), .ZN(n9450) );
  NAND2_X1 U10629 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n9450), .ZN(n9452) );
  XOR2_X1 U10630 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n9450), .Z(n10082) );
  NAND2_X1 U10631 ( .A1(n10082), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n9451) );
  NAND2_X1 U10632 ( .A1(n9452), .A2(n9451), .ZN(n9453) );
  AND2_X1 U10633 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n9453), .ZN(n9454) );
  XNOR2_X1 U10634 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n9453), .ZN(n10079) );
  INV_X1 U10635 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10078) );
  NOR2_X1 U10636 ( .A1(n10079), .A2(n10078), .ZN(n10077) );
  NAND2_X1 U10637 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n9455) );
  OAI21_X1 U10638 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n9455), .ZN(n10075) );
  NAND2_X1 U10639 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n9456) );
  OAI21_X1 U10640 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n9456), .ZN(n10072) );
  NOR2_X1 U10641 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n9457) );
  AOI21_X1 U10642 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n9457), .ZN(n10069) );
  NAND2_X1 U10643 ( .A1(n10070), .A2(n10069), .ZN(n10068) );
  NAND2_X1 U10644 ( .A1(n10067), .A2(n10066), .ZN(n10065) );
  NAND2_X1 U10645 ( .A1(n10064), .A2(n10063), .ZN(n10062) );
  OAI21_X1 U10646 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10062), .ZN(n10060) );
  NAND2_X1 U10647 ( .A1(n10061), .A2(n10060), .ZN(n10059) );
  OAI21_X1 U10648 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10059), .ZN(n10057) );
  NAND2_X1 U10649 ( .A1(n10058), .A2(n10057), .ZN(n10056) );
  OAI21_X1 U10650 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10056), .ZN(n10054) );
  NAND2_X1 U10651 ( .A1(n10055), .A2(n10054), .ZN(n10053) );
  NOR2_X1 U10652 ( .A1(n10085), .A2(n10084), .ZN(n9458) );
  NAND2_X1 U10653 ( .A1(n10085), .A2(n10084), .ZN(n10083) );
  OAI21_X1 U10654 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n9458), .A(n10083), .ZN(
        n9649) );
  AOI22_X1 U10655 ( .A1(P2_REG3_REG_1__SCAN_IN), .A2(keyinput_f44), .B1(SI_10_), .B2(keyinput_f22), .ZN(n9459) );
  OAI221_X1 U10656 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(keyinput_f44), .C1(
        SI_10_), .C2(keyinput_f22), .A(n9459), .ZN(n9466) );
  AOI22_X1 U10657 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(keyinput_f43), .B1(SI_13_), .B2(keyinput_f19), .ZN(n9460) );
  OAI221_X1 U10658 ( .B1(P2_REG3_REG_8__SCAN_IN), .B2(keyinput_f43), .C1(
        SI_13_), .C2(keyinput_f19), .A(n9460), .ZN(n9465) );
  AOI22_X1 U10659 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(keyinput_f49), .B1(SI_19_), .B2(keyinput_f13), .ZN(n9461) );
  OAI221_X1 U10660 ( .B1(P2_REG3_REG_5__SCAN_IN), .B2(keyinput_f49), .C1(
        SI_19_), .C2(keyinput_f13), .A(n9461), .ZN(n9464) );
  AOI22_X1 U10661 ( .A1(P2_REG3_REG_25__SCAN_IN), .A2(keyinput_f47), .B1(SI_7_), .B2(keyinput_f25), .ZN(n9462) );
  OAI221_X1 U10662 ( .B1(P2_REG3_REG_25__SCAN_IN), .B2(keyinput_f47), .C1(
        SI_7_), .C2(keyinput_f25), .A(n9462), .ZN(n9463) );
  NOR4_X1 U10663 ( .A1(n9466), .A2(n9465), .A3(n9464), .A4(n9463), .ZN(n9494)
         );
  XNOR2_X1 U10664 ( .A(P2_RD_REG_SCAN_IN), .B(keyinput_f33), .ZN(n9474) );
  AOI22_X1 U10665 ( .A1(SI_17_), .A2(keyinput_f15), .B1(n9468), .B2(
        keyinput_f45), .ZN(n9467) );
  OAI221_X1 U10666 ( .B1(SI_17_), .B2(keyinput_f15), .C1(n9468), .C2(
        keyinput_f45), .A(n9467), .ZN(n9473) );
  AOI22_X1 U10667 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(keyinput_f60), .B1(SI_0_), .B2(keyinput_f32), .ZN(n9469) );
  OAI221_X1 U10668 ( .B1(P2_REG3_REG_18__SCAN_IN), .B2(keyinput_f60), .C1(
        SI_0_), .C2(keyinput_f32), .A(n9469), .ZN(n9472) );
  AOI22_X1 U10669 ( .A1(SI_12_), .A2(keyinput_f20), .B1(SI_20_), .B2(
        keyinput_f12), .ZN(n9470) );
  OAI221_X1 U10670 ( .B1(SI_12_), .B2(keyinput_f20), .C1(SI_20_), .C2(
        keyinput_f12), .A(n9470), .ZN(n9471) );
  NOR4_X1 U10671 ( .A1(n9474), .A2(n9473), .A3(n9472), .A4(n9471), .ZN(n9493)
         );
  AOI22_X1 U10672 ( .A1(SI_5_), .A2(keyinput_f27), .B1(SI_23_), .B2(
        keyinput_f9), .ZN(n9475) );
  OAI221_X1 U10673 ( .B1(SI_5_), .B2(keyinput_f27), .C1(SI_23_), .C2(
        keyinput_f9), .A(n9475), .ZN(n9482) );
  AOI22_X1 U10674 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(keyinput_f51), .B1(
        SI_18_), .B2(keyinput_f14), .ZN(n9476) );
  OAI221_X1 U10675 ( .B1(P2_REG3_REG_24__SCAN_IN), .B2(keyinput_f51), .C1(
        SI_18_), .C2(keyinput_f14), .A(n9476), .ZN(n9481) );
  AOI22_X1 U10676 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(keyinput_f41), .B1(SI_3_), .B2(keyinput_f29), .ZN(n9477) );
  OAI221_X1 U10677 ( .B1(P2_REG3_REG_19__SCAN_IN), .B2(keyinput_f41), .C1(
        SI_3_), .C2(keyinput_f29), .A(n9477), .ZN(n9480) );
  AOI22_X1 U10678 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(keyinput_f39), .B1(
        P2_REG3_REG_20__SCAN_IN), .B2(keyinput_f55), .ZN(n9478) );
  OAI221_X1 U10679 ( .B1(P2_REG3_REG_10__SCAN_IN), .B2(keyinput_f39), .C1(
        P2_REG3_REG_20__SCAN_IN), .C2(keyinput_f55), .A(n9478), .ZN(n9479) );
  NOR4_X1 U10680 ( .A1(n9482), .A2(n9481), .A3(n9480), .A4(n9479), .ZN(n9492)
         );
  AOI22_X1 U10681 ( .A1(SI_30_), .A2(keyinput_f2), .B1(P2_REG3_REG_26__SCAN_IN), .B2(keyinput_f62), .ZN(n9483) );
  OAI221_X1 U10682 ( .B1(SI_30_), .B2(keyinput_f2), .C1(
        P2_REG3_REG_26__SCAN_IN), .C2(keyinput_f62), .A(n9483), .ZN(n9490) );
  AOI22_X1 U10683 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(keyinput_f36), .B1(
        SI_16_), .B2(keyinput_f16), .ZN(n9484) );
  OAI221_X1 U10684 ( .B1(P2_REG3_REG_27__SCAN_IN), .B2(keyinput_f36), .C1(
        SI_16_), .C2(keyinput_f16), .A(n9484), .ZN(n9489) );
  AOI22_X1 U10685 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(keyinput_f53), .B1(
        P2_REG3_REG_11__SCAN_IN), .B2(keyinput_f58), .ZN(n9485) );
  OAI221_X1 U10686 ( .B1(P2_REG3_REG_9__SCAN_IN), .B2(keyinput_f53), .C1(
        P2_REG3_REG_11__SCAN_IN), .C2(keyinput_f58), .A(n9485), .ZN(n9488) );
  AOI22_X1 U10687 ( .A1(SI_4_), .A2(keyinput_f28), .B1(SI_21_), .B2(
        keyinput_f11), .ZN(n9486) );
  OAI221_X1 U10688 ( .B1(SI_4_), .B2(keyinput_f28), .C1(SI_21_), .C2(
        keyinput_f11), .A(n9486), .ZN(n9487) );
  NOR4_X1 U10689 ( .A1(n9490), .A2(n9489), .A3(n9488), .A4(n9487), .ZN(n9491)
         );
  NAND4_X1 U10690 ( .A1(n9494), .A2(n9493), .A3(n9492), .A4(n9491), .ZN(n9549)
         );
  INV_X1 U10691 ( .A(P2_WR_REG_SCAN_IN), .ZN(n9587) );
  AOI22_X1 U10692 ( .A1(n9496), .A2(keyinput_f24), .B1(keyinput_f0), .B2(n9587), .ZN(n9495) );
  OAI221_X1 U10693 ( .B1(n9496), .B2(keyinput_f24), .C1(n9587), .C2(
        keyinput_f0), .A(n9495), .ZN(n9507) );
  AOI22_X1 U10694 ( .A1(n5771), .A2(keyinput_f35), .B1(n9498), .B2(keyinput_f7), .ZN(n9497) );
  OAI221_X1 U10695 ( .B1(n5771), .B2(keyinput_f35), .C1(n9498), .C2(
        keyinput_f7), .A(n9497), .ZN(n9506) );
  AOI22_X1 U10696 ( .A1(n9500), .A2(keyinput_f50), .B1(keyinput_f46), .B2(
        n9593), .ZN(n9499) );
  OAI221_X1 U10697 ( .B1(n9500), .B2(keyinput_f50), .C1(n9593), .C2(
        keyinput_f46), .A(n9499), .ZN(n9505) );
  AOI22_X1 U10698 ( .A1(n9503), .A2(keyinput_f48), .B1(n9502), .B2(
        keyinput_f38), .ZN(n9501) );
  OAI221_X1 U10699 ( .B1(n9503), .B2(keyinput_f48), .C1(n9502), .C2(
        keyinput_f38), .A(n9501), .ZN(n9504) );
  NOR4_X1 U10700 ( .A1(n9507), .A2(n9506), .A3(n9505), .A4(n9504), .ZN(n9547)
         );
  AOI22_X1 U10701 ( .A1(P2_REG3_REG_28__SCAN_IN), .A2(keyinput_f42), .B1(
        SI_28_), .B2(keyinput_f4), .ZN(n9508) );
  OAI221_X1 U10702 ( .B1(P2_REG3_REG_28__SCAN_IN), .B2(keyinput_f42), .C1(
        SI_28_), .C2(keyinput_f4), .A(n9508), .ZN(n9518) );
  AOI22_X1 U10703 ( .A1(P2_REG3_REG_22__SCAN_IN), .A2(keyinput_f57), .B1(
        SI_15_), .B2(keyinput_f17), .ZN(n9509) );
  OAI221_X1 U10704 ( .B1(P2_REG3_REG_22__SCAN_IN), .B2(keyinput_f57), .C1(
        SI_15_), .C2(keyinput_f17), .A(n9509), .ZN(n9517) );
  AOI22_X1 U10705 ( .A1(n9512), .A2(keyinput_f59), .B1(n9511), .B2(
        keyinput_f61), .ZN(n9510) );
  OAI221_X1 U10706 ( .B1(n9512), .B2(keyinput_f59), .C1(n9511), .C2(
        keyinput_f61), .A(n9510), .ZN(n9516) );
  AOI22_X1 U10707 ( .A1(P2_STATE_REG_SCAN_IN), .A2(keyinput_f34), .B1(n9514), 
        .B2(keyinput_f3), .ZN(n9513) );
  OAI221_X1 U10708 ( .B1(P2_STATE_REG_SCAN_IN), .B2(keyinput_f34), .C1(n9514), 
        .C2(keyinput_f3), .A(n9513), .ZN(n9515) );
  NOR4_X1 U10709 ( .A1(n9518), .A2(n9517), .A3(n9516), .A4(n9515), .ZN(n9546)
         );
  AOI22_X1 U10710 ( .A1(n5869), .A2(keyinput_f56), .B1(n9520), .B2(keyinput_f6), .ZN(n9519) );
  OAI221_X1 U10711 ( .B1(n5869), .B2(keyinput_f56), .C1(n9520), .C2(
        keyinput_f6), .A(n9519), .ZN(n9531) );
  AOI22_X1 U10712 ( .A1(n9522), .A2(keyinput_f21), .B1(keyinput_f1), .B2(n7857), .ZN(n9521) );
  OAI221_X1 U10713 ( .B1(n9522), .B2(keyinput_f21), .C1(n7857), .C2(
        keyinput_f1), .A(n9521), .ZN(n9530) );
  AOI22_X1 U10714 ( .A1(n9524), .A2(keyinput_f54), .B1(n5912), .B2(
        keyinput_f63), .ZN(n9523) );
  OAI221_X1 U10715 ( .B1(n9524), .B2(keyinput_f54), .C1(n5912), .C2(
        keyinput_f63), .A(n9523), .ZN(n9529) );
  AOI22_X1 U10716 ( .A1(n9527), .A2(keyinput_f23), .B1(n9526), .B2(
        keyinput_f10), .ZN(n9525) );
  OAI221_X1 U10717 ( .B1(n9527), .B2(keyinput_f23), .C1(n9526), .C2(
        keyinput_f10), .A(n9525), .ZN(n9528) );
  NOR4_X1 U10718 ( .A1(n9531), .A2(n9530), .A3(n9529), .A4(n9528), .ZN(n9545)
         );
  INV_X1 U10719 ( .A(SI_6_), .ZN(n9630) );
  AOI22_X1 U10720 ( .A1(n9533), .A2(keyinput_f18), .B1(keyinput_f26), .B2(
        n9630), .ZN(n9532) );
  OAI221_X1 U10721 ( .B1(n9533), .B2(keyinput_f18), .C1(n9630), .C2(
        keyinput_f26), .A(n9532), .ZN(n9543) );
  AOI22_X1 U10722 ( .A1(n9605), .A2(keyinput_f40), .B1(keyinput_f52), .B2(
        n9629), .ZN(n9534) );
  OAI221_X1 U10723 ( .B1(n9605), .B2(keyinput_f40), .C1(n9629), .C2(
        keyinput_f52), .A(n9534), .ZN(n9542) );
  AOI22_X1 U10724 ( .A1(n9537), .A2(keyinput_f37), .B1(n9536), .B2(keyinput_f5), .ZN(n9535) );
  OAI221_X1 U10725 ( .B1(n9537), .B2(keyinput_f37), .C1(n9536), .C2(
        keyinput_f5), .A(n9535), .ZN(n9541) );
  XOR2_X1 U10726 ( .A(n5391), .B(keyinput_f8), .Z(n9539) );
  XNOR2_X1 U10727 ( .A(SI_1_), .B(keyinput_f31), .ZN(n9538) );
  NAND2_X1 U10728 ( .A1(n9539), .A2(n9538), .ZN(n9540) );
  NOR4_X1 U10729 ( .A1(n9543), .A2(n9542), .A3(n9541), .A4(n9540), .ZN(n9544)
         );
  NAND4_X1 U10730 ( .A1(n9547), .A2(n9546), .A3(n9545), .A4(n9544), .ZN(n9548)
         );
  OAI22_X1 U10731 ( .A1(n9549), .A2(n9548), .B1(keyinput_f30), .B2(SI_2_), 
        .ZN(n9550) );
  AOI21_X1 U10732 ( .B1(keyinput_f30), .B2(SI_2_), .A(n9550), .ZN(n9647) );
  AOI22_X1 U10733 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(keyinput_g49), .B1(SI_7_), 
        .B2(keyinput_g25), .ZN(n9551) );
  OAI221_X1 U10734 ( .B1(P2_REG3_REG_5__SCAN_IN), .B2(keyinput_g49), .C1(SI_7_), .C2(keyinput_g25), .A(n9551), .ZN(n9558) );
  AOI22_X1 U10735 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(keyinput_g56), .B1(
        SI_26_), .B2(keyinput_g6), .ZN(n9552) );
  OAI221_X1 U10736 ( .B1(P2_REG3_REG_13__SCAN_IN), .B2(keyinput_g56), .C1(
        SI_26_), .C2(keyinput_g6), .A(n9552), .ZN(n9557) );
  AOI22_X1 U10737 ( .A1(P2_REG3_REG_22__SCAN_IN), .A2(keyinput_g57), .B1(
        P2_REG3_REG_23__SCAN_IN), .B2(keyinput_g38), .ZN(n9553) );
  OAI221_X1 U10738 ( .B1(P2_REG3_REG_22__SCAN_IN), .B2(keyinput_g57), .C1(
        P2_REG3_REG_23__SCAN_IN), .C2(keyinput_g38), .A(n9553), .ZN(n9556) );
  AOI22_X1 U10739 ( .A1(P2_STATE_REG_SCAN_IN), .A2(keyinput_g34), .B1(SI_11_), 
        .B2(keyinput_g21), .ZN(n9554) );
  OAI221_X1 U10740 ( .B1(P2_STATE_REG_SCAN_IN), .B2(keyinput_g34), .C1(SI_11_), 
        .C2(keyinput_g21), .A(n9554), .ZN(n9555) );
  NOR4_X1 U10741 ( .A1(n9558), .A2(n9557), .A3(n9556), .A4(n9555), .ZN(n9585)
         );
  XOR2_X1 U10742 ( .A(SI_14_), .B(keyinput_g18), .Z(n9565) );
  AOI22_X1 U10743 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(keyinput_g51), .B1(
        SI_22_), .B2(keyinput_g10), .ZN(n9559) );
  OAI221_X1 U10744 ( .B1(P2_REG3_REG_24__SCAN_IN), .B2(keyinput_g51), .C1(
        SI_22_), .C2(keyinput_g10), .A(n9559), .ZN(n9564) );
  AOI22_X1 U10745 ( .A1(P2_REG3_REG_0__SCAN_IN), .A2(keyinput_g54), .B1(SI_12_), .B2(keyinput_g20), .ZN(n9560) );
  OAI221_X1 U10746 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(keyinput_g54), .C1(
        SI_12_), .C2(keyinput_g20), .A(n9560), .ZN(n9563) );
  AOI22_X1 U10747 ( .A1(P2_REG3_REG_1__SCAN_IN), .A2(keyinput_g44), .B1(
        P2_REG3_REG_7__SCAN_IN), .B2(keyinput_g35), .ZN(n9561) );
  OAI221_X1 U10748 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(keyinput_g44), .C1(
        P2_REG3_REG_7__SCAN_IN), .C2(keyinput_g35), .A(n9561), .ZN(n9562) );
  NOR4_X1 U10749 ( .A1(n9565), .A2(n9564), .A3(n9563), .A4(n9562), .ZN(n9584)
         );
  AOI22_X1 U10750 ( .A1(P2_REG3_REG_26__SCAN_IN), .A2(keyinput_g62), .B1(
        SI_27_), .B2(keyinput_g5), .ZN(n9566) );
  OAI221_X1 U10751 ( .B1(P2_REG3_REG_26__SCAN_IN), .B2(keyinput_g62), .C1(
        SI_27_), .C2(keyinput_g5), .A(n9566), .ZN(n9573) );
  AOI22_X1 U10752 ( .A1(SI_29_), .A2(keyinput_g3), .B1(P2_REG3_REG_25__SCAN_IN), .B2(keyinput_g47), .ZN(n9567) );
  OAI221_X1 U10753 ( .B1(SI_29_), .B2(keyinput_g3), .C1(
        P2_REG3_REG_25__SCAN_IN), .C2(keyinput_g47), .A(n9567), .ZN(n9572) );
  AOI22_X1 U10754 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(keyinput_g63), .B1(SI_8_), .B2(keyinput_g24), .ZN(n9568) );
  OAI221_X1 U10755 ( .B1(P2_REG3_REG_15__SCAN_IN), .B2(keyinput_g63), .C1(
        SI_8_), .C2(keyinput_g24), .A(n9568), .ZN(n9571) );
  AOI22_X1 U10756 ( .A1(SI_3_), .A2(keyinput_g29), .B1(SI_10_), .B2(
        keyinput_g22), .ZN(n9569) );
  OAI221_X1 U10757 ( .B1(SI_3_), .B2(keyinput_g29), .C1(SI_10_), .C2(
        keyinput_g22), .A(n9569), .ZN(n9570) );
  NOR4_X1 U10758 ( .A1(n9573), .A2(n9572), .A3(n9571), .A4(n9570), .ZN(n9583)
         );
  AOI22_X1 U10759 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(keyinput_g61), .B1(SI_4_), 
        .B2(keyinput_g28), .ZN(n9574) );
  OAI221_X1 U10760 ( .B1(P2_REG3_REG_6__SCAN_IN), .B2(keyinput_g61), .C1(SI_4_), .C2(keyinput_g28), .A(n9574), .ZN(n9581) );
  AOI22_X1 U10761 ( .A1(SI_31_), .A2(keyinput_g1), .B1(P2_REG3_REG_10__SCAN_IN), .B2(keyinput_g39), .ZN(n9575) );
  OAI221_X1 U10762 ( .B1(SI_31_), .B2(keyinput_g1), .C1(
        P2_REG3_REG_10__SCAN_IN), .C2(keyinput_g39), .A(n9575), .ZN(n9580) );
  AOI22_X1 U10763 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(keyinput_g48), .B1(SI_9_), .B2(keyinput_g23), .ZN(n9576) );
  OAI221_X1 U10764 ( .B1(P2_REG3_REG_16__SCAN_IN), .B2(keyinput_g48), .C1(
        SI_9_), .C2(keyinput_g23), .A(n9576), .ZN(n9579) );
  AOI22_X1 U10765 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(keyinput_g50), .B1(
        P2_REG3_REG_18__SCAN_IN), .B2(keyinput_g60), .ZN(n9577) );
  OAI221_X1 U10766 ( .B1(P2_REG3_REG_17__SCAN_IN), .B2(keyinput_g50), .C1(
        P2_REG3_REG_18__SCAN_IN), .C2(keyinput_g60), .A(n9577), .ZN(n9578) );
  NOR4_X1 U10767 ( .A1(n9581), .A2(n9580), .A3(n9579), .A4(n9578), .ZN(n9582)
         );
  NAND4_X1 U10768 ( .A1(n9585), .A2(n9584), .A3(n9583), .A4(n9582), .ZN(n9645)
         );
  AOI22_X1 U10769 ( .A1(n9587), .A2(keyinput_g0), .B1(n5391), .B2(keyinput_g8), 
        .ZN(n9586) );
  OAI221_X1 U10770 ( .B1(n9587), .B2(keyinput_g0), .C1(n5391), .C2(keyinput_g8), .A(n9586), .ZN(n9600) );
  AOI22_X1 U10771 ( .A1(n9590), .A2(keyinput_g43), .B1(n9589), .B2(
        keyinput_g11), .ZN(n9588) );
  OAI221_X1 U10772 ( .B1(n9590), .B2(keyinput_g43), .C1(n9589), .C2(
        keyinput_g11), .A(n9588), .ZN(n9599) );
  AOI22_X1 U10773 ( .A1(n9593), .A2(keyinput_g46), .B1(n9592), .B2(
        keyinput_g27), .ZN(n9591) );
  OAI221_X1 U10774 ( .B1(n9593), .B2(keyinput_g46), .C1(n9592), .C2(
        keyinput_g27), .A(n9591), .ZN(n9598) );
  AOI22_X1 U10775 ( .A1(n9596), .A2(keyinput_g4), .B1(n9595), .B2(keyinput_g12), .ZN(n9594) );
  OAI221_X1 U10776 ( .B1(n9596), .B2(keyinput_g4), .C1(n9595), .C2(
        keyinput_g12), .A(n9594), .ZN(n9597) );
  NOR4_X1 U10777 ( .A1(n9600), .A2(n9599), .A3(n9598), .A4(n9597), .ZN(n9643)
         );
  AOI22_X1 U10778 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(keyinput_g58), .B1(
        P2_REG3_REG_14__SCAN_IN), .B2(keyinput_g37), .ZN(n9601) );
  OAI221_X1 U10779 ( .B1(P2_REG3_REG_11__SCAN_IN), .B2(keyinput_g58), .C1(
        P2_REG3_REG_14__SCAN_IN), .C2(keyinput_g37), .A(n9601), .ZN(n9611) );
  AOI22_X1 U10780 ( .A1(P2_REG3_REG_2__SCAN_IN), .A2(keyinput_g59), .B1(SI_25_), .B2(keyinput_g7), .ZN(n9602) );
  OAI221_X1 U10781 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(keyinput_g59), .C1(
        SI_25_), .C2(keyinput_g7), .A(n9602), .ZN(n9610) );
  AOI22_X1 U10782 ( .A1(n9605), .A2(keyinput_g40), .B1(keyinput_g2), .B2(n9604), .ZN(n9603) );
  OAI221_X1 U10783 ( .B1(n9605), .B2(keyinput_g40), .C1(n9604), .C2(
        keyinput_g2), .A(n9603), .ZN(n9609) );
  INV_X1 U10784 ( .A(SI_18_), .ZN(n9607) );
  AOI22_X1 U10785 ( .A1(n5801), .A2(keyinput_g53), .B1(n9607), .B2(
        keyinput_g14), .ZN(n9606) );
  OAI221_X1 U10786 ( .B1(n5801), .B2(keyinput_g53), .C1(n9607), .C2(
        keyinput_g14), .A(n9606), .ZN(n9608) );
  NOR4_X1 U10787 ( .A1(n9611), .A2(n9610), .A3(n9609), .A4(n9608), .ZN(n9642)
         );
  AOI22_X1 U10788 ( .A1(n9614), .A2(keyinput_g9), .B1(keyinput_g16), .B2(n9613), .ZN(n9612) );
  OAI221_X1 U10789 ( .B1(n9614), .B2(keyinput_g9), .C1(n9613), .C2(
        keyinput_g16), .A(n9612), .ZN(n9626) );
  AOI22_X1 U10790 ( .A1(n9617), .A2(keyinput_g19), .B1(keyinput_g55), .B2(
        n9616), .ZN(n9615) );
  OAI221_X1 U10791 ( .B1(n9617), .B2(keyinput_g19), .C1(n9616), .C2(
        keyinput_g55), .A(n9615), .ZN(n9625) );
  AOI22_X1 U10792 ( .A1(n9620), .A2(keyinput_g41), .B1(n9619), .B2(
        keyinput_g17), .ZN(n9618) );
  OAI221_X1 U10793 ( .B1(n9620), .B2(keyinput_g41), .C1(n9619), .C2(
        keyinput_g17), .A(n9618), .ZN(n9624) );
  XNOR2_X1 U10794 ( .A(P2_REG3_REG_21__SCAN_IN), .B(keyinput_g45), .ZN(n9622)
         );
  XNOR2_X1 U10795 ( .A(SI_1_), .B(keyinput_g31), .ZN(n9621) );
  NAND2_X1 U10796 ( .A1(n9622), .A2(n9621), .ZN(n9623) );
  NOR4_X1 U10797 ( .A1(n9626), .A2(n9625), .A3(n9624), .A4(n9623), .ZN(n9641)
         );
  AOI22_X1 U10798 ( .A1(n5265), .A2(keyinput_g15), .B1(keyinput_g42), .B2(
        n6137), .ZN(n9627) );
  OAI221_X1 U10799 ( .B1(n5265), .B2(keyinput_g15), .C1(n6137), .C2(
        keyinput_g42), .A(n9627), .ZN(n9639) );
  AOI22_X1 U10800 ( .A1(n9630), .A2(keyinput_g26), .B1(keyinput_g52), .B2(
        n9629), .ZN(n9628) );
  OAI221_X1 U10801 ( .B1(n9630), .B2(keyinput_g26), .C1(n9629), .C2(
        keyinput_g52), .A(n9628), .ZN(n9638) );
  AOI22_X1 U10802 ( .A1(n9633), .A2(keyinput_g32), .B1(n9632), .B2(
        keyinput_g13), .ZN(n9631) );
  OAI221_X1 U10803 ( .B1(n9633), .B2(keyinput_g32), .C1(n9632), .C2(
        keyinput_g13), .A(n9631), .ZN(n9637) );
  XNOR2_X1 U10804 ( .A(P2_REG3_REG_27__SCAN_IN), .B(keyinput_g36), .ZN(n9635)
         );
  XNOR2_X1 U10805 ( .A(P2_RD_REG_SCAN_IN), .B(keyinput_g33), .ZN(n9634) );
  NAND2_X1 U10806 ( .A1(n9635), .A2(n9634), .ZN(n9636) );
  NOR4_X1 U10807 ( .A1(n9639), .A2(n9638), .A3(n9637), .A4(n9636), .ZN(n9640)
         );
  NAND4_X1 U10808 ( .A1(n9643), .A2(n9642), .A3(n9641), .A4(n9640), .ZN(n9644)
         );
  OAI22_X1 U10809 ( .A1(SI_2_), .A2(keyinput_g30), .B1(n9645), .B2(n9644), 
        .ZN(n9646) );
  AOI211_X1 U10810 ( .C1(SI_2_), .C2(keyinput_g30), .A(n9647), .B(n9646), .ZN(
        n9648) );
  XNOR2_X1 U10811 ( .A(n9649), .B(n9648), .ZN(n9653) );
  NOR2_X1 U10812 ( .A1(n9651), .A2(n9650), .ZN(n9652) );
  XOR2_X1 U10813 ( .A(n9653), .B(n9652), .Z(ADD_1071_U4) );
  OAI22_X1 U10814 ( .A1(n9656), .A2(n9655), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9654), .ZN(n9661) );
  NAND2_X1 U10815 ( .A1(n9990), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n9659) );
  AOI211_X1 U10816 ( .C1(n9659), .C2(n9658), .A(n9657), .B(n9983), .ZN(n9660)
         );
  AOI211_X1 U10817 ( .C1(n9674), .C2(n9662), .A(n9661), .B(n9660), .ZN(n9668)
         );
  NOR2_X1 U10818 ( .A1(n9988), .A2(n9663), .ZN(n9666) );
  OAI211_X1 U10819 ( .C1(n9666), .C2(n9665), .A(n9980), .B(n9664), .ZN(n9667)
         );
  NAND2_X1 U10820 ( .A1(n9668), .A2(n9667), .ZN(P2_U3246) );
  AOI22_X1 U10821 ( .A1(n9985), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n9680) );
  AOI211_X1 U10822 ( .C1(n9671), .C2(n9670), .A(n9669), .B(n9983), .ZN(n9672)
         );
  AOI21_X1 U10823 ( .B1(n9674), .B2(n9673), .A(n9672), .ZN(n9679) );
  OAI211_X1 U10824 ( .C1(n9677), .C2(n9676), .A(n9980), .B(n9675), .ZN(n9678)
         );
  NAND3_X1 U10825 ( .A1(n9680), .A2(n9679), .A3(n9678), .ZN(P2_U3247) );
  OAI211_X1 U10826 ( .C1(n9961), .C2(n9683), .A(n9682), .B(n9681), .ZN(n9686)
         );
  NOR2_X1 U10827 ( .A1(n9684), .A2(n9946), .ZN(n9685) );
  AOI211_X1 U10828 ( .C1(n9965), .C2(n9687), .A(n9686), .B(n9685), .ZN(n9689)
         );
  INV_X1 U10829 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n9688) );
  AOI22_X1 U10830 ( .A1(n9968), .A2(n9689), .B1(n9688), .B2(n9966), .ZN(
        P1_U3484) );
  AOI22_X1 U10831 ( .A1(n9978), .A2(n9689), .B1(n6552), .B2(n9975), .ZN(
        P1_U3533) );
  INV_X1 U10832 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n9694) );
  AOI22_X1 U10833 ( .A1(n10048), .A2(n9701), .B1(n9694), .B2(n10046), .ZN(
        P2_U3551) );
  OAI21_X1 U10834 ( .B1(n9696), .B2(n10031), .A(n9695), .ZN(n9697) );
  AOI21_X1 U10835 ( .B1(n9698), .B2(n7178), .A(n9697), .ZN(n9703) );
  INV_X1 U10836 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n9699) );
  AOI22_X1 U10837 ( .A1(n10048), .A2(n9703), .B1(n9699), .B2(n10046), .ZN(
        P2_U3550) );
  INV_X1 U10838 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n9700) );
  AOI22_X1 U10839 ( .A1(n4314), .A2(n9701), .B1(n9700), .B2(n10036), .ZN(
        P2_U3519) );
  INV_X1 U10840 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n9702) );
  AOI22_X1 U10841 ( .A1(n4314), .A2(n9703), .B1(n9702), .B2(n10036), .ZN(
        P2_U3518) );
  INV_X1 U10842 ( .A(n9704), .ZN(n9705) );
  AOI21_X1 U10843 ( .B1(n9707), .B2(n9706), .A(n9705), .ZN(n9708) );
  OAI21_X1 U10844 ( .B1(n9710), .B2(n9709), .A(n9708), .ZN(n9711) );
  AOI21_X1 U10845 ( .B1(n9712), .B2(n8638), .A(n9711), .ZN(n9720) );
  NAND2_X1 U10846 ( .A1(n9714), .A2(n9713), .ZN(n9716) );
  XNOR2_X1 U10847 ( .A(n9716), .B(n9715), .ZN(n9718) );
  NAND2_X1 U10848 ( .A1(n9718), .A2(n9717), .ZN(n9719) );
  OAI211_X1 U10849 ( .C1(n9722), .C2(n9721), .A(n9720), .B(n9719), .ZN(
        P1_U3239) );
  INV_X1 U10850 ( .A(n9723), .ZN(n9724) );
  AOI21_X1 U10851 ( .B1(n9726), .B2(n9725), .A(n9724), .ZN(n9766) );
  XNOR2_X1 U10852 ( .A(n9727), .B(n9726), .ZN(n9733) );
  AOI22_X1 U10853 ( .A1(n9730), .A2(n9729), .B1(n9728), .B2(n9925), .ZN(n9731)
         );
  OAI21_X1 U10854 ( .B1(n9733), .B2(n9732), .A(n9731), .ZN(n9734) );
  AOI21_X1 U10855 ( .B1(n9766), .B2(n9735), .A(n9734), .ZN(n9763) );
  AOI222_X1 U10856 ( .A1(n9738), .A2(n9737), .B1(P1_REG2_REG_11__SCAN_IN), 
        .B2(n9938), .C1(n9896), .C2(n9736), .ZN(n9744) );
  INV_X1 U10857 ( .A(n9739), .ZN(n9741) );
  OAI211_X1 U10858 ( .C1(n9741), .C2(n9762), .A(n9877), .B(n9740), .ZN(n9761)
         );
  INV_X1 U10859 ( .A(n9761), .ZN(n9742) );
  AOI22_X1 U10860 ( .A1(n9766), .A2(n9882), .B1(n9881), .B2(n9742), .ZN(n9743)
         );
  OAI211_X1 U10861 ( .C1(n9938), .C2(n9763), .A(n9744), .B(n9743), .ZN(
        P1_U3280) );
  OAI211_X1 U10862 ( .C1(n9961), .C2(n9747), .A(n9746), .B(n9745), .ZN(n9748)
         );
  AOI21_X1 U10863 ( .B1(n9749), .B2(n9957), .A(n9748), .ZN(n9769) );
  AOI22_X1 U10864 ( .A1(n9978), .A2(n9769), .B1(n7059), .B2(n9975), .ZN(
        P1_U3537) );
  OAI21_X1 U10865 ( .B1(n9961), .B2(n9751), .A(n9750), .ZN(n9752) );
  AOI21_X1 U10866 ( .B1(n9753), .B2(n9965), .A(n9752), .ZN(n9754) );
  AND2_X1 U10867 ( .A1(n9755), .A2(n9754), .ZN(n9771) );
  AOI22_X1 U10868 ( .A1(n9978), .A2(n9771), .B1(n6774), .B2(n9975), .ZN(
        P1_U3536) );
  OAI211_X1 U10869 ( .C1(n9961), .C2(n9758), .A(n9757), .B(n9756), .ZN(n9759)
         );
  AOI21_X1 U10870 ( .B1(n9760), .B2(n9957), .A(n9759), .ZN(n9773) );
  AOI22_X1 U10871 ( .A1(n9978), .A2(n9773), .B1(n6610), .B2(n9975), .ZN(
        P1_U3535) );
  OAI21_X1 U10872 ( .B1(n9961), .B2(n9762), .A(n9761), .ZN(n9765) );
  INV_X1 U10873 ( .A(n9763), .ZN(n9764) );
  AOI211_X1 U10874 ( .C1(n9965), .C2(n9766), .A(n9765), .B(n9764), .ZN(n9775)
         );
  AOI22_X1 U10875 ( .A1(n9978), .A2(n9775), .B1(n9767), .B2(n9975), .ZN(
        P1_U3534) );
  INV_X1 U10876 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n9768) );
  AOI22_X1 U10877 ( .A1(n9968), .A2(n9769), .B1(n9768), .B2(n9966), .ZN(
        P1_U3496) );
  INV_X1 U10878 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n9770) );
  AOI22_X1 U10879 ( .A1(n9968), .A2(n9771), .B1(n9770), .B2(n9966), .ZN(
        P1_U3493) );
  INV_X1 U10880 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n9772) );
  AOI22_X1 U10881 ( .A1(n9968), .A2(n9773), .B1(n9772), .B2(n9966), .ZN(
        P1_U3490) );
  INV_X1 U10882 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n9774) );
  AOI22_X1 U10883 ( .A1(n9968), .A2(n9775), .B1(n9774), .B2(n9966), .ZN(
        P1_U3487) );
  XNOR2_X1 U10884 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  INV_X1 U10885 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n9782) );
  NOR2_X1 U10886 ( .A1(n9969), .A2(P1_IR_REG_0__SCAN_IN), .ZN(n9776) );
  NOR2_X1 U10887 ( .A1(n9777), .A2(n9776), .ZN(n9779) );
  OR3_X1 U10888 ( .A1(n9780), .A2(n9779), .A3(n9778), .ZN(n9781) );
  OAI21_X1 U10889 ( .B1(n9873), .B2(n9782), .A(n9781), .ZN(n9783) );
  INV_X1 U10890 ( .A(n9783), .ZN(n9785) );
  OR3_X1 U10891 ( .A1(n9797), .A2(P1_REG1_REG_0__SCAN_IN), .A3(n7713), .ZN(
        n9784) );
  OAI211_X1 U10892 ( .C1(P1_STATE_REG_SCAN_IN), .C2(n9786), .A(n9785), .B(
        n9784), .ZN(P1_U3241) );
  MUX2_X1 U10893 ( .A(n6319), .B(P1_REG2_REG_2__SCAN_IN), .S(n9792), .Z(n9789)
         );
  INV_X1 U10894 ( .A(n9787), .ZN(n9788) );
  NAND2_X1 U10895 ( .A1(n9789), .A2(n9788), .ZN(n9790) );
  NAND3_X1 U10896 ( .A1(n9869), .A2(n9791), .A3(n9790), .ZN(n9794) );
  NAND2_X1 U10897 ( .A1(n9860), .A2(n9792), .ZN(n9793) );
  NAND2_X1 U10898 ( .A1(n9794), .A2(n9793), .ZN(n9796) );
  AOI211_X1 U10899 ( .C1(n9854), .C2(P1_ADDR_REG_2__SCAN_IN), .A(n9796), .B(
        n9795), .ZN(n9803) );
  AOI211_X1 U10900 ( .C1(n9800), .C2(n9799), .A(n9798), .B(n9797), .ZN(n9801)
         );
  INV_X1 U10901 ( .A(n9801), .ZN(n9802) );
  OAI211_X1 U10902 ( .C1(P1_STATE_REG_SCAN_IN), .C2(n9804), .A(n9803), .B(
        n9802), .ZN(P1_U3243) );
  AOI22_X1 U10903 ( .A1(n9854), .A2(P1_ADDR_REG_5__SCAN_IN), .B1(n9805), .B2(
        n9860), .ZN(n9816) );
  AOI21_X1 U10904 ( .B1(n9808), .B2(n9807), .A(n9806), .ZN(n9809) );
  OR2_X1 U10905 ( .A1(n9847), .A2(n9809), .ZN(n9814) );
  OAI211_X1 U10906 ( .C1(n9812), .C2(n9811), .A(n9868), .B(n9810), .ZN(n9813)
         );
  NAND4_X1 U10907 ( .A1(n9816), .A2(n9815), .A3(n9814), .A4(n9813), .ZN(
        P1_U3246) );
  XOR2_X1 U10908 ( .A(n5072), .B(n9821), .Z(n9817) );
  XNOR2_X1 U10909 ( .A(n9818), .B(n9817), .ZN(n9819) );
  AOI22_X1 U10910 ( .A1(n9819), .A2(n9869), .B1(n9854), .B2(
        P1_ADDR_REG_8__SCAN_IN), .ZN(n9830) );
  INV_X1 U10911 ( .A(n9820), .ZN(n9829) );
  AND3_X1 U10912 ( .A1(n9826), .A2(P1_REG1_REG_8__SCAN_IN), .A3(n9868), .ZN(
        n9822) );
  OAI21_X1 U10913 ( .B1(n9822), .B2(n9860), .A(n9821), .ZN(n9828) );
  NAND2_X1 U10914 ( .A1(n9824), .A2(n9823), .ZN(n9825) );
  OAI211_X1 U10915 ( .C1(n9826), .C2(n9825), .A(n9834), .B(n9868), .ZN(n9827)
         );
  NAND4_X1 U10916 ( .A1(n9830), .A2(n9829), .A3(n9828), .A4(n9827), .ZN(
        P1_U3249) );
  AOI22_X1 U10917 ( .A1(n9854), .A2(P1_ADDR_REG_9__SCAN_IN), .B1(n9831), .B2(
        n9860), .ZN(n9842) );
  OAI21_X1 U10918 ( .B1(n9834), .B2(n9833), .A(n9832), .ZN(n9840) );
  AOI211_X1 U10919 ( .C1(n9837), .C2(n9836), .A(n9847), .B(n9835), .ZN(n9838)
         );
  AOI211_X1 U10920 ( .C1(n9868), .C2(n9840), .A(n9839), .B(n9838), .ZN(n9841)
         );
  NAND2_X1 U10921 ( .A1(n9842), .A2(n9841), .ZN(P1_U3250) );
  OAI21_X1 U10922 ( .B1(n9845), .B2(n9844), .A(n9843), .ZN(n9852) );
  AOI211_X1 U10923 ( .C1(n9849), .C2(n9848), .A(n9847), .B(n9846), .ZN(n9850)
         );
  AOI211_X1 U10924 ( .C1(n9868), .C2(n9852), .A(n9851), .B(n9850), .ZN(n9856)
         );
  AOI22_X1 U10925 ( .A1(n9854), .A2(P1_ADDR_REG_10__SCAN_IN), .B1(n9853), .B2(
        n9860), .ZN(n9855) );
  NAND2_X1 U10926 ( .A1(n9856), .A2(n9855), .ZN(P1_U3251) );
  INV_X1 U10927 ( .A(n9857), .ZN(n9858) );
  AOI21_X1 U10928 ( .B1(n9860), .B2(n9859), .A(n9858), .ZN(n9872) );
  AOI21_X1 U10929 ( .B1(n9863), .B2(n9862), .A(n9861), .ZN(n9870) );
  OAI21_X1 U10930 ( .B1(n9866), .B2(n9865), .A(n9864), .ZN(n9867) );
  AOI22_X1 U10931 ( .A1(n9870), .A2(n9869), .B1(n9868), .B2(n9867), .ZN(n9871)
         );
  OAI211_X1 U10932 ( .C1(n9873), .C2(n10085), .A(n9872), .B(n9871), .ZN(
        P1_U3259) );
  XNOR2_X1 U10933 ( .A(n9874), .B(n9885), .ZN(n9895) );
  INV_X1 U10934 ( .A(n9895), .ZN(n9964) );
  INV_X1 U10935 ( .A(n9875), .ZN(n9960) );
  INV_X1 U10936 ( .A(n9876), .ZN(n9878) );
  OAI211_X1 U10937 ( .C1(n9960), .C2(n9879), .A(n9878), .B(n9877), .ZN(n9959)
         );
  INV_X1 U10938 ( .A(n9959), .ZN(n9880) );
  AOI22_X1 U10939 ( .A1(n9964), .A2(n9882), .B1(n9881), .B2(n9880), .ZN(n9902)
         );
  NAND2_X1 U10940 ( .A1(n9883), .A2(n9884), .ZN(n9886) );
  XNOR2_X1 U10941 ( .A(n9886), .B(n9885), .ZN(n9893) );
  OAI22_X1 U10942 ( .A1(n9890), .A2(n9889), .B1(n9888), .B2(n9887), .ZN(n9891)
         );
  AOI21_X1 U10943 ( .B1(n9893), .B2(n9892), .A(n9891), .ZN(n9894) );
  OAI21_X1 U10944 ( .B1(n9895), .B2(n9946), .A(n9894), .ZN(n9962) );
  AOI22_X1 U10945 ( .A1(n9938), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n9897), .B2(
        n9896), .ZN(n9898) );
  OAI21_X1 U10946 ( .B1(n9960), .B2(n9899), .A(n9898), .ZN(n9900) );
  AOI21_X1 U10947 ( .B1(n9962), .B2(n9918), .A(n9900), .ZN(n9901) );
  NAND2_X1 U10948 ( .A1(n9902), .A2(n9901), .ZN(P1_U3282) );
  INV_X1 U10949 ( .A(n9903), .ZN(n9914) );
  INV_X1 U10950 ( .A(n9904), .ZN(n9912) );
  NAND2_X1 U10951 ( .A1(n9896), .A2(n9905), .ZN(n9906) );
  OAI211_X1 U10952 ( .C1(n9909), .C2(n9908), .A(n9907), .B(n9906), .ZN(n9910)
         );
  AOI21_X1 U10953 ( .B1(n9912), .B2(n9911), .A(n9910), .ZN(n9913) );
  OAI21_X1 U10954 ( .B1(n9915), .B2(n9914), .A(n9913), .ZN(n9917) );
  NOR2_X1 U10955 ( .A1(n9917), .A2(n9916), .ZN(n9919) );
  AOI22_X1 U10956 ( .A1(n9938), .A2(n6329), .B1(n9919), .B2(n9918), .ZN(
        P1_U3286) );
  NAND2_X1 U10957 ( .A1(n9921), .A2(n9920), .ZN(n9935) );
  INV_X1 U10958 ( .A(n9922), .ZN(n9929) );
  OR3_X1 U10959 ( .A1(n9924), .A2(n9929), .A3(n9923), .ZN(n9928) );
  NAND2_X1 U10960 ( .A1(n9926), .A2(n9925), .ZN(n9927) );
  AND2_X1 U10961 ( .A1(n9928), .A2(n9927), .ZN(n9932) );
  INV_X1 U10962 ( .A(n9932), .ZN(n9934) );
  NAND2_X1 U10963 ( .A1(n9930), .A2(n9929), .ZN(n9931) );
  AND2_X1 U10964 ( .A1(n9932), .A2(n9931), .ZN(n9970) );
  INV_X1 U10965 ( .A(n9970), .ZN(n9933) );
  OAI21_X1 U10966 ( .B1(n9935), .B2(n9934), .A(n9933), .ZN(n9937) );
  AOI22_X1 U10967 ( .A1(n9896), .A2(P1_REG3_REG_0__SCAN_IN), .B1(
        P1_REG2_REG_0__SCAN_IN), .B2(n9938), .ZN(n9936) );
  OAI21_X1 U10968 ( .B1(n9938), .B2(n9937), .A(n9936), .ZN(P1_U3291) );
  AND2_X1 U10969 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9939), .ZN(P1_U3292) );
  AND2_X1 U10970 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9939), .ZN(P1_U3293) );
  AND2_X1 U10971 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9939), .ZN(P1_U3294) );
  AND2_X1 U10972 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9939), .ZN(P1_U3295) );
  AND2_X1 U10973 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9939), .ZN(P1_U3296) );
  AND2_X1 U10974 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9939), .ZN(P1_U3297) );
  AND2_X1 U10975 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9939), .ZN(P1_U3298) );
  AND2_X1 U10976 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9939), .ZN(P1_U3299) );
  AND2_X1 U10977 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9939), .ZN(P1_U3300) );
  AND2_X1 U10978 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9939), .ZN(P1_U3301) );
  AND2_X1 U10979 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9939), .ZN(P1_U3302) );
  AND2_X1 U10980 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9939), .ZN(P1_U3303) );
  AND2_X1 U10981 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9939), .ZN(P1_U3304) );
  AND2_X1 U10982 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9939), .ZN(P1_U3305) );
  AND2_X1 U10983 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9939), .ZN(P1_U3306) );
  AND2_X1 U10984 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9939), .ZN(P1_U3307) );
  AND2_X1 U10985 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9939), .ZN(P1_U3308) );
  AND2_X1 U10986 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9939), .ZN(P1_U3309) );
  AND2_X1 U10987 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9939), .ZN(P1_U3310) );
  AND2_X1 U10988 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9939), .ZN(P1_U3311) );
  AND2_X1 U10989 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9939), .ZN(P1_U3312) );
  AND2_X1 U10990 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9939), .ZN(P1_U3313) );
  AND2_X1 U10991 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9939), .ZN(P1_U3314) );
  AND2_X1 U10992 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9939), .ZN(P1_U3315) );
  AND2_X1 U10993 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9939), .ZN(P1_U3316) );
  AND2_X1 U10994 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9939), .ZN(P1_U3317) );
  AND2_X1 U10995 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9939), .ZN(P1_U3318) );
  AND2_X1 U10996 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9939), .ZN(P1_U3319) );
  AND2_X1 U10997 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9939), .ZN(P1_U3320) );
  AND2_X1 U10998 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9939), .ZN(P1_U3321) );
  INV_X1 U10999 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n9940) );
  AOI22_X1 U11000 ( .A1(n9968), .A2(n9970), .B1(n9940), .B2(n9966), .ZN(
        P1_U3454) );
  NAND2_X1 U11001 ( .A1(n9942), .A2(n9941), .ZN(n9943) );
  OAI211_X1 U11002 ( .C1(n9947), .C2(n9945), .A(n9944), .B(n9943), .ZN(n9949)
         );
  NOR2_X1 U11003 ( .A1(n9947), .A2(n9946), .ZN(n9948) );
  NOR3_X1 U11004 ( .A1(n9950), .A2(n9949), .A3(n9948), .ZN(n9972) );
  INV_X1 U11005 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9951) );
  AOI22_X1 U11006 ( .A1(n9968), .A2(n9972), .B1(n9951), .B2(n9966), .ZN(
        P1_U3457) );
  OAI21_X1 U11007 ( .B1(n9961), .B2(n9953), .A(n9952), .ZN(n9955) );
  AOI211_X1 U11008 ( .C1(n9957), .C2(n9956), .A(n9955), .B(n9954), .ZN(n9974)
         );
  INV_X1 U11009 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9958) );
  AOI22_X1 U11010 ( .A1(n9968), .A2(n9974), .B1(n9958), .B2(n9966), .ZN(
        P1_U3475) );
  OAI21_X1 U11011 ( .B1(n9961), .B2(n9960), .A(n9959), .ZN(n9963) );
  AOI211_X1 U11012 ( .C1(n9965), .C2(n9964), .A(n9963), .B(n9962), .ZN(n9977)
         );
  INV_X1 U11013 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9967) );
  AOI22_X1 U11014 ( .A1(n9968), .A2(n9977), .B1(n9967), .B2(n9966), .ZN(
        P1_U3481) );
  AOI22_X1 U11015 ( .A1(n9978), .A2(n9970), .B1(n9969), .B2(n9975), .ZN(
        P1_U3523) );
  AOI22_X1 U11016 ( .A1(n9978), .A2(n9972), .B1(n9971), .B2(n9975), .ZN(
        P1_U3524) );
  AOI22_X1 U11017 ( .A1(n9978), .A2(n9974), .B1(n9973), .B2(n9975), .ZN(
        P1_U3530) );
  INV_X1 U11018 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n9976) );
  AOI22_X1 U11019 ( .A1(n9978), .A2(n9977), .B1(n9976), .B2(n9975), .ZN(
        P1_U3532) );
  AOI22_X1 U11020 ( .A1(n9980), .A2(P2_REG2_REG_0__SCAN_IN), .B1(n9979), .B2(
        P2_REG1_REG_0__SCAN_IN), .ZN(n9989) );
  NAND2_X1 U11021 ( .A1(n9980), .A2(n9663), .ZN(n9982) );
  OAI211_X1 U11022 ( .C1(P2_REG1_REG_0__SCAN_IN), .C2(n9983), .A(n9982), .B(
        n9981), .ZN(n9984) );
  INV_X1 U11023 ( .A(n9984), .ZN(n9987) );
  AOI22_X1 U11024 ( .A1(n9985), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n9986) );
  OAI221_X1 U11025 ( .B1(n9990), .B2(n9989), .C1(n9988), .C2(n9987), .A(n9986), 
        .ZN(P2_U3245) );
  AND2_X1 U11026 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n9995), .ZN(P2_U3297) );
  AND2_X1 U11027 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n9995), .ZN(P2_U3298) );
  AND2_X1 U11028 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n9995), .ZN(P2_U3299) );
  AND2_X1 U11029 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n9995), .ZN(P2_U3300) );
  AND2_X1 U11030 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n9995), .ZN(P2_U3301) );
  AND2_X1 U11031 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n9995), .ZN(P2_U3302) );
  AND2_X1 U11032 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n9995), .ZN(P2_U3303) );
  AND2_X1 U11033 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n9995), .ZN(P2_U3304) );
  AND2_X1 U11034 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n9995), .ZN(P2_U3305) );
  AND2_X1 U11035 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n9995), .ZN(P2_U3306) );
  AND2_X1 U11036 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n9995), .ZN(P2_U3307) );
  AND2_X1 U11037 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n9995), .ZN(P2_U3308) );
  AND2_X1 U11038 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n9995), .ZN(P2_U3309) );
  AND2_X1 U11039 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n9995), .ZN(P2_U3310) );
  AND2_X1 U11040 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n9995), .ZN(P2_U3311) );
  AND2_X1 U11041 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n9995), .ZN(P2_U3312) );
  AND2_X1 U11042 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n9995), .ZN(P2_U3313) );
  AND2_X1 U11043 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n9995), .ZN(P2_U3314) );
  AND2_X1 U11044 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n9995), .ZN(P2_U3315) );
  AND2_X1 U11045 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n9995), .ZN(P2_U3316) );
  AND2_X1 U11046 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n9995), .ZN(P2_U3317) );
  AND2_X1 U11047 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n9995), .ZN(P2_U3318) );
  AND2_X1 U11048 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n9995), .ZN(P2_U3319) );
  AND2_X1 U11049 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n9995), .ZN(P2_U3320) );
  AND2_X1 U11050 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n9995), .ZN(P2_U3321) );
  AND2_X1 U11051 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n9995), .ZN(P2_U3322) );
  AND2_X1 U11052 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n9995), .ZN(P2_U3323) );
  AND2_X1 U11053 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n9995), .ZN(P2_U3324) );
  AND2_X1 U11054 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n9995), .ZN(P2_U3325) );
  AND2_X1 U11055 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n9995), .ZN(P2_U3326) );
  AOI22_X1 U11056 ( .A1(n9998), .A2(n9994), .B1(n9993), .B2(n9995), .ZN(
        P2_U3437) );
  AOI22_X1 U11057 ( .A1(n9998), .A2(n9997), .B1(n9996), .B2(n9995), .ZN(
        P2_U3438) );
  INV_X1 U11058 ( .A(n9999), .ZN(n10000) );
  OAI21_X1 U11059 ( .B1(n10001), .B2(n10022), .A(n10000), .ZN(n10003) );
  AOI211_X1 U11060 ( .C1(n10034), .C2(n10004), .A(n10003), .B(n10002), .ZN(
        n10039) );
  INV_X1 U11061 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10005) );
  AOI22_X1 U11062 ( .A1(n4314), .A2(n10039), .B1(n10005), .B2(n10036), .ZN(
        P2_U3454) );
  INV_X1 U11063 ( .A(n10006), .ZN(n10027) );
  INV_X1 U11064 ( .A(n10007), .ZN(n10009) );
  OAI22_X1 U11065 ( .A1(n10009), .A2(n10022), .B1(n10008), .B2(n10031), .ZN(
        n10011) );
  AOI211_X1 U11066 ( .C1(n10027), .C2(n10012), .A(n10011), .B(n10010), .ZN(
        n10041) );
  INV_X1 U11067 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10013) );
  AOI22_X1 U11068 ( .A1(n4314), .A2(n10041), .B1(n10013), .B2(n10036), .ZN(
        P2_U3460) );
  OAI22_X1 U11069 ( .A1(n10015), .A2(n10022), .B1(n10014), .B2(n10031), .ZN(
        n10017) );
  AOI211_X1 U11070 ( .C1(n10018), .C2(n10034), .A(n10017), .B(n10016), .ZN(
        n10043) );
  INV_X1 U11071 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10019) );
  AOI22_X1 U11072 ( .A1(n4314), .A2(n10043), .B1(n10019), .B2(n10036), .ZN(
        P2_U3472) );
  INV_X1 U11073 ( .A(n10020), .ZN(n10026) );
  OAI22_X1 U11074 ( .A1(n10023), .A2(n10022), .B1(n10021), .B2(n10031), .ZN(
        n10025) );
  AOI211_X1 U11075 ( .C1(n10027), .C2(n10026), .A(n10025), .B(n10024), .ZN(
        n10045) );
  INV_X1 U11076 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10028) );
  AOI22_X1 U11077 ( .A1(n4314), .A2(n10045), .B1(n10028), .B2(n10036), .ZN(
        P2_U3478) );
  OAI211_X1 U11078 ( .C1(n10032), .C2(n10031), .A(n10030), .B(n10029), .ZN(
        n10033) );
  AOI21_X1 U11079 ( .B1(n10035), .B2(n10034), .A(n10033), .ZN(n10047) );
  INV_X1 U11080 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10037) );
  AOI22_X1 U11081 ( .A1(n4314), .A2(n10047), .B1(n10037), .B2(n10036), .ZN(
        P2_U3484) );
  INV_X1 U11082 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10038) );
  AOI22_X1 U11083 ( .A1(n10048), .A2(n10039), .B1(n10038), .B2(n10046), .ZN(
        P2_U3521) );
  INV_X1 U11084 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10040) );
  AOI22_X1 U11085 ( .A1(n10048), .A2(n10041), .B1(n10040), .B2(n10046), .ZN(
        P2_U3523) );
  INV_X1 U11086 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n10042) );
  AOI22_X1 U11087 ( .A1(n10048), .A2(n10043), .B1(n10042), .B2(n10046), .ZN(
        P2_U3527) );
  AOI22_X1 U11088 ( .A1(n10048), .A2(n10045), .B1(n10044), .B2(n10046), .ZN(
        P2_U3529) );
  AOI22_X1 U11089 ( .A1(n10048), .A2(n10047), .B1(n6519), .B2(n10046), .ZN(
        P2_U3531) );
  INV_X1 U11090 ( .A(n10049), .ZN(n10050) );
  NAND2_X1 U11091 ( .A1(n10051), .A2(n10050), .ZN(n10052) );
  XNOR2_X1 U11092 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n10052), .ZN(ADD_1071_U5)
         );
  XOR2_X1 U11093 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  OAI21_X1 U11094 ( .B1(n10055), .B2(n10054), .A(n10053), .ZN(ADD_1071_U56) );
  OAI21_X1 U11095 ( .B1(n10058), .B2(n10057), .A(n10056), .ZN(ADD_1071_U57) );
  OAI21_X1 U11096 ( .B1(n10061), .B2(n10060), .A(n10059), .ZN(ADD_1071_U58) );
  OAI21_X1 U11097 ( .B1(n10064), .B2(n10063), .A(n10062), .ZN(ADD_1071_U59) );
  OAI21_X1 U11098 ( .B1(n10067), .B2(n10066), .A(n10065), .ZN(ADD_1071_U60) );
  OAI21_X1 U11099 ( .B1(n10070), .B2(n10069), .A(n10068), .ZN(ADD_1071_U61) );
  AOI21_X1 U11100 ( .B1(n10073), .B2(n10072), .A(n10071), .ZN(ADD_1071_U62) );
  AOI21_X1 U11101 ( .B1(n10076), .B2(n10075), .A(n10074), .ZN(ADD_1071_U63) );
  AOI21_X1 U11102 ( .B1(n10079), .B2(n10078), .A(n10077), .ZN(ADD_1071_U47) );
  XOR2_X1 U11103 ( .A(n10081), .B(n10080), .Z(ADD_1071_U54) );
  XOR2_X1 U11104 ( .A(n10082), .B(P2_ADDR_REG_8__SCAN_IN), .Z(ADD_1071_U48) );
  OAI21_X1 U11105 ( .B1(n10085), .B2(n10084), .A(n10083), .ZN(n10086) );
  XNOR2_X1 U11106 ( .A(n10086), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  XOR2_X1 U11107 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(n10087), .Z(ADD_1071_U49) );
  XOR2_X1 U11108 ( .A(P2_ADDR_REG_6__SCAN_IN), .B(n10088), .Z(ADD_1071_U50) );
  AOI21_X1 U11109 ( .B1(n10090), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n10089), .ZN(
        n10092) );
  XNOR2_X1 U11110 ( .A(n10092), .B(n10091), .ZN(ADD_1071_U51) );
  XOR2_X1 U11111 ( .A(n10094), .B(n10093), .Z(ADD_1071_U53) );
  XNOR2_X1 U11112 ( .A(n10096), .B(n10095), .ZN(ADD_1071_U52) );
  INV_X2 U4814 ( .A(n7736), .ZN(n7673) );
  XNOR2_X1 U4845 ( .A(n5656), .B(n5655), .ZN(n6149) );
  CLKBUF_X1 U6171 ( .A(n5508), .Z(n4317) );
endmodule

