

module b21_C_SARLock_k_64_1 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3, 
        keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, 
        keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, 
        keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, 
        keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, 
        keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, 
        keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, 
        keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, 
        keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, 
        keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, 
        keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, 
        ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58, 
        ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63, 
        ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51, 
        ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46, 
        U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, 
        P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, 
        P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, 
        P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, 
        P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440, P1_U3441, 
        P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, 
        P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, 
        P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, 
        P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, 
        P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463, P1_U3466, 
        P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484, P1_U3487, 
        P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505, P1_U3508, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289, P1_U3288, 
        P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, 
        P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, 
        P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, 
        P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262, P1_U3261, 
        P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, 
        P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, 
        P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238, P1_U3237, 
        P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, 
        P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, 
        P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, 
        P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084, P1_U3083, 
        P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354, P2_U3353, 
        P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347, P2_U3346, 
        P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340, P2_U3339, 
        P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333, P2_U3332, 
        P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437, P2_U3438, 
        P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, 
        P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, 
        P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, 
        P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, 
        P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, 
        P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, 
        P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502, P2_U3505, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, 
        P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533, P2_U3534, 
        P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, 
        P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, 
        P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294, P2_U3293, 
        P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, 
        P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, 
        P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, 
        P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, 
        P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, 
        P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, 
        P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3552, 
        P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, 
        P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565, P2_U3566, 
        P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572, P2_U3573, 
        P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579, P2_U3580, 
        P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152, P2_U3151, 
        P2_U3966 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4273, n4274, n4275, n4276, n4277, n4278, n4280, n4281, n4282, n4283,
         n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293,
         n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303,
         n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
         n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
         n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333,
         n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
         n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353,
         n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
         n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373,
         n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383,
         n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
         n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403,
         n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413,
         n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423,
         n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433,
         n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443,
         n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453,
         n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
         n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473,
         n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
         n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
         n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
         n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
         n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
         n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
         n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
         n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
         n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
         n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
         n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693,
         n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703,
         n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713,
         n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723,
         n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733,
         n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743,
         n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753,
         n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763,
         n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773,
         n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783,
         n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793,
         n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803,
         n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813,
         n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823,
         n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833,
         n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843,
         n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853,
         n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863,
         n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873,
         n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883,
         n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893,
         n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903,
         n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913,
         n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923,
         n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933,
         n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943,
         n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953,
         n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963,
         n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973,
         n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983,
         n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993,
         n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003,
         n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013,
         n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023,
         n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033,
         n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043,
         n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053,
         n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063,
         n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073,
         n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083,
         n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093,
         n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103,
         n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113,
         n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123,
         n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133,
         n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143,
         n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153,
         n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163,
         n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173,
         n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183,
         n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193,
         n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203,
         n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213,
         n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223,
         n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233,
         n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243,
         n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253,
         n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263,
         n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273,
         n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283,
         n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293,
         n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303,
         n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313,
         n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323,
         n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333,
         n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343,
         n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353,
         n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363,
         n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373,
         n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383,
         n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393,
         n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403,
         n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413,
         n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423,
         n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433,
         n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443,
         n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453,
         n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463,
         n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473,
         n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483,
         n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493,
         n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503,
         n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513,
         n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523,
         n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533,
         n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543,
         n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553,
         n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563,
         n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573,
         n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583,
         n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593,
         n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603,
         n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613,
         n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623,
         n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633,
         n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643,
         n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653,
         n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663,
         n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673,
         n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683,
         n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693,
         n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703,
         n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713,
         n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723,
         n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733,
         n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743,
         n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753,
         n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763,
         n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773,
         n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783,
         n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793,
         n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803,
         n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813,
         n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823,
         n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833,
         n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843,
         n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853,
         n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863,
         n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873,
         n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883,
         n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893,
         n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903,
         n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913,
         n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923,
         n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933,
         n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943,
         n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953,
         n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963,
         n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973,
         n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983,
         n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993,
         n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003,
         n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013,
         n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023,
         n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033,
         n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043,
         n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053,
         n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063,
         n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073,
         n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083,
         n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093,
         n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103,
         n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113,
         n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123,
         n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133,
         n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143,
         n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153,
         n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163,
         n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173,
         n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183,
         n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193,
         n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203,
         n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213,
         n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223,
         n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233,
         n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243,
         n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253,
         n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263,
         n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273,
         n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283,
         n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293,
         n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303,
         n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313,
         n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323,
         n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333,
         n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343,
         n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353,
         n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363,
         n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373,
         n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383,
         n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393,
         n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403,
         n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413,
         n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423,
         n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433,
         n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443,
         n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453,
         n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463,
         n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473,
         n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483,
         n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493,
         n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503,
         n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513,
         n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523,
         n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533,
         n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543,
         n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553,
         n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6563, n6564,
         n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
         n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
         n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
         n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
         n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
         n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624,
         n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634,
         n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644,
         n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654,
         n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664,
         n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674,
         n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684,
         n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694,
         n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704,
         n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714,
         n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724,
         n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734,
         n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744,
         n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754,
         n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764,
         n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774,
         n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784,
         n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794,
         n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804,
         n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814,
         n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824,
         n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834,
         n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844,
         n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854,
         n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864,
         n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874,
         n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884,
         n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894,
         n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904,
         n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914,
         n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924,
         n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934,
         n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944,
         n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954,
         n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964,
         n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974,
         n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984,
         n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994,
         n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004,
         n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014,
         n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024,
         n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034,
         n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044,
         n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054,
         n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064,
         n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074,
         n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084,
         n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094,
         n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104,
         n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114,
         n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124,
         n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134,
         n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144,
         n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154,
         n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164,
         n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174,
         n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184,
         n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194,
         n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204,
         n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214,
         n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224,
         n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234,
         n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244,
         n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254,
         n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264,
         n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274,
         n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284,
         n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294,
         n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304,
         n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314,
         n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324,
         n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334,
         n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344,
         n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354,
         n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364,
         n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374,
         n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384,
         n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394,
         n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404,
         n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414,
         n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424,
         n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434,
         n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444,
         n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454,
         n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464,
         n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474,
         n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484,
         n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494,
         n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504,
         n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514,
         n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524,
         n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534,
         n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544,
         n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554,
         n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564,
         n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574,
         n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584,
         n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594,
         n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604,
         n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614,
         n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624,
         n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634,
         n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644,
         n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654,
         n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664,
         n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674,
         n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684,
         n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694,
         n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704,
         n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714,
         n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724,
         n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734,
         n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744,
         n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754,
         n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764,
         n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774,
         n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784,
         n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794,
         n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804,
         n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814,
         n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824,
         n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834,
         n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844,
         n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854,
         n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864,
         n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874,
         n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884,
         n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894,
         n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904,
         n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914,
         n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924,
         n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934,
         n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944,
         n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954,
         n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964,
         n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974,
         n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984,
         n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994,
         n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004,
         n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014,
         n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024,
         n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034,
         n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044,
         n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054,
         n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064,
         n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074,
         n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084,
         n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094,
         n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104,
         n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114,
         n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124,
         n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134,
         n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144,
         n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154,
         n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164,
         n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174,
         n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184,
         n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194,
         n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204,
         n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214,
         n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224,
         n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234,
         n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244,
         n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254,
         n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264,
         n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274,
         n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284,
         n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294,
         n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304,
         n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314,
         n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324,
         n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334,
         n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344,
         n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354,
         n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364,
         n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374,
         n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384,
         n8385, n8386, n8387, n8388, n8389, n8391, n8392, n8393, n8394, n8395,
         n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405,
         n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415,
         n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425,
         n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435,
         n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445,
         n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455,
         n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465,
         n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475,
         n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485,
         n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495,
         n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505,
         n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515,
         n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525,
         n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535,
         n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545,
         n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555,
         n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565,
         n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575,
         n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585,
         n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595,
         n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605,
         n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615,
         n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625,
         n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635,
         n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645,
         n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655,
         n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665,
         n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675,
         n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685,
         n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695,
         n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705,
         n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715,
         n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725,
         n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735,
         n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745,
         n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755,
         n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765,
         n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775,
         n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785,
         n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795,
         n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805,
         n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815,
         n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825,
         n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835,
         n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845,
         n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855,
         n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865,
         n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875,
         n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885,
         n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895,
         n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905,
         n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915,
         n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925,
         n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935,
         n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945,
         n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955,
         n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965,
         n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975,
         n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985,
         n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995,
         n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005,
         n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015,
         n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025,
         n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035,
         n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045,
         n9046, n9047, n9048, n9049, n9050, n9052, n9053, n9054, n9055, n9056,
         n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066,
         n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076,
         n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086,
         n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096,
         n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106,
         n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116,
         n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126,
         n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136,
         n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146,
         n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156,
         n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166,
         n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176,
         n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186,
         n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196,
         n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206,
         n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216,
         n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226,
         n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236,
         n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246,
         n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256,
         n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266,
         n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276,
         n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286,
         n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296,
         n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306,
         n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316,
         n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326,
         n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336,
         n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346,
         n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356,
         n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366,
         n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376,
         n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386,
         n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396,
         n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406,
         n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416,
         n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426,
         n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436,
         n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446,
         n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456,
         n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466,
         n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476,
         n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486,
         n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496,
         n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506,
         n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516,
         n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526,
         n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536,
         n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546,
         n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556,
         n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566,
         n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576,
         n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586,
         n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596,
         n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606,
         n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616,
         n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626,
         n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636,
         n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646,
         n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656,
         n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666,
         n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676,
         n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686,
         n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696,
         n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706,
         n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716,
         n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726,
         n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736,
         n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746,
         n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756,
         n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766,
         n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776,
         n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786,
         n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796,
         n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806,
         n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816,
         n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826,
         n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836,
         n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846,
         n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856,
         n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866,
         n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876,
         n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886,
         n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896,
         n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906,
         n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916,
         n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926,
         n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936,
         n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946,
         n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956,
         n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966,
         n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976,
         n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986,
         n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996,
         n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005,
         n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013,
         n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021,
         n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029,
         n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037,
         n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045,
         n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053,
         n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061,
         n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069,
         n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077,
         n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085,
         n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093,
         n10096;

  INV_X2 U4779 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  CLKBUF_X2 U4780 ( .A(n5247), .Z(n4286) );
  AND3_X1 U4781 ( .A1(n5150), .A2(n5149), .A3(n5148), .ZN(n9829) );
  CLKBUF_X2 U4782 ( .A(n5792), .Z(n6722) );
  AND2_X1 U4783 ( .A1(n8059), .A2(n9050), .ZN(n5792) );
  NAND2_X2 U4784 ( .A1(n5035), .A2(n5038), .ZN(n5166) );
  INV_X1 U4785 ( .A(n9829), .ZN(n7116) );
  INV_X1 U4786 ( .A(n5797), .ZN(n8084) );
  NAND2_X1 U4787 ( .A1(n5700), .A2(n5051), .ZN(n5171) );
  INV_X1 U4788 ( .A(n5700), .ZN(n5570) );
  OR2_X1 U4789 ( .A1(n9246), .A2(n9401), .ZN(n9221) );
  INV_X1 U4790 ( .A(n6108), .ZN(n6152) );
  INV_X1 U4791 ( .A(n9815), .ZN(n7255) );
  NAND2_X1 U4792 ( .A1(n9258), .A2(n9406), .ZN(n9246) );
  AND2_X1 U4793 ( .A1(n4997), .A2(n4996), .ZN(n9307) );
  AND2_X1 U4794 ( .A1(n7829), .A2(n4363), .ZN(n8043) );
  AND3_X1 U4795 ( .A1(n5197), .A2(n5196), .A3(n5195), .ZN(n9836) );
  INV_X1 U4796 ( .A(n6305), .ZN(n4568) );
  AND2_X2 U4797 ( .A1(n4863), .A2(n4862), .ZN(n4873) );
  INV_X1 U4798 ( .A(n5108), .ZN(n6416) );
  OR2_X1 U4799 ( .A1(n9050), .A2(n5736), .ZN(n4273) );
  NAND2_X2 U4800 ( .A1(n7279), .A2(n5208), .ZN(n8308) );
  NAND2_X2 U4801 ( .A1(n6886), .A2(n5203), .ZN(n7279) );
  NAND2_X2 U4802 ( .A1(n4396), .A2(n4394), .ZN(n8487) );
  NAND2_X1 U4803 ( .A1(n5671), .A2(n4280), .ZN(n4274) );
  NAND2_X1 U4804 ( .A1(n5671), .A2(n4280), .ZN(n5110) );
  INV_X4 U4805 ( .A(n5110), .ZN(n6579) );
  INV_X2 U4806 ( .A(n4273), .ZN(n4275) );
  INV_X1 U4807 ( .A(n5093), .ZN(n4276) );
  OR2_X4 U4808 ( .A1(n5064), .A2(n5013), .ZN(n5093) );
  INV_X1 U4809 ( .A(n4873), .ZN(n4277) );
  INV_X2 U4810 ( .A(n4873), .ZN(n4278) );
  INV_X1 U4812 ( .A(n10096), .ZN(n4280) );
  NOR2_X2 U4813 ( .A1(n5344), .A2(n5008), .ZN(n5650) );
  AND2_X1 U4814 ( .A1(n6382), .A2(n6381), .ZN(n6426) );
  NAND2_X1 U4815 ( .A1(n4418), .A2(n4333), .ZN(n8755) );
  NAND2_X1 U4816 ( .A1(n8074), .A2(n4611), .ZN(n8798) );
  NOR2_X1 U4817 ( .A1(n8436), .A2(n4824), .ZN(n4823) );
  INV_X1 U4818 ( .A(n9307), .ZN(n9429) );
  OR2_X1 U4819 ( .A1(n7208), .A2(n9470), .ZN(n9570) );
  AND2_X1 U4820 ( .A1(n5125), .A2(n5086), .ZN(n6753) );
  NAND2_X1 U4821 ( .A1(n8143), .A2(n7590), .ZN(n7081) );
  NAND2_X1 U4822 ( .A1(n7071), .A2(n7070), .ZN(n8146) );
  INV_X4 U4823 ( .A(n5760), .ZN(n7043) );
  CLKBUF_X2 U4824 ( .A(P1_U4006), .Z(n4281) );
  NAND2_X2 U4825 ( .A1(n9953), .A2(n8265), .ZN(n5760) );
  INV_X2 U4826 ( .A(n7072), .ZN(n7071) );
  BUF_X2 U4827 ( .A(n5806), .Z(n6093) );
  BUF_X2 U4828 ( .A(n4275), .Z(n6068) );
  CLKBUF_X1 U4829 ( .A(n8088), .Z(n4284) );
  INV_X2 U4830 ( .A(n5166), .ZN(n5087) );
  NAND2_X1 U4831 ( .A1(n8389), .A2(n5038), .ZN(n5237) );
  INV_X1 U4832 ( .A(n5241), .ZN(n4290) );
  AND2_X1 U4833 ( .A1(n5739), .A2(n5738), .ZN(n5744) );
  INV_X4 U4834 ( .A(n4873), .ZN(n4283) );
  NAND2_X1 U4835 ( .A1(n5757), .A2(n4386), .ZN(n5798) );
  AND2_X1 U4836 ( .A1(n9135), .A2(n4858), .ZN(n5717) );
  OAI21_X1 U4837 ( .B1(n9239), .B2(n4795), .A(n4794), .ZN(n9184) );
  NOR2_X1 U4838 ( .A1(n8446), .A2(n8447), .ZN(n8445) );
  AOI21_X1 U4839 ( .B1(n9233), .B2(n9786), .A(n9232), .ZN(n9404) );
  NAND2_X1 U4840 ( .A1(n9240), .A2(n9199), .ZN(n9226) );
  OAI21_X1 U4841 ( .B1(n9098), .B2(n4618), .A(n4616), .ZN(n5525) );
  NAND2_X1 U4842 ( .A1(n9242), .A2(n9241), .ZN(n9240) );
  INV_X1 U4843 ( .A(n4796), .ZN(n4795) );
  AOI21_X1 U4844 ( .B1(n4796), .B2(n9241), .A(n4368), .ZN(n4794) );
  OAI22_X1 U4845 ( .A1(n8735), .A2(n8741), .B1(n8607), .B2(n8970), .ZN(n8723)
         );
  NOR2_X1 U4846 ( .A1(n9246), .A2(n4584), .ZN(n9212) );
  NAND2_X1 U4847 ( .A1(n4664), .A2(n4662), .ZN(n9282) );
  AOI21_X1 U4848 ( .B1(n4666), .B2(n4668), .A(n4663), .ZN(n4662) );
  OR2_X1 U4849 ( .A1(n7871), .A2(n5404), .ZN(n4445) );
  NAND2_X1 U4850 ( .A1(n8826), .A2(n8072), .ZN(n8827) );
  NAND2_X1 U4851 ( .A1(n4631), .A2(n5361), .ZN(n7871) );
  NAND2_X1 U4852 ( .A1(n9358), .A2(n9359), .ZN(n9365) );
  NAND2_X1 U4853 ( .A1(n5533), .A2(n5532), .ZN(n9423) );
  AOI21_X1 U4854 ( .B1(n4681), .B2(n4676), .A(n4675), .ZN(n7981) );
  NAND2_X1 U4855 ( .A1(n7640), .A2(n5316), .ZN(n7652) );
  NAND2_X1 U4856 ( .A1(n6084), .A2(n6083), .ZN(n8970) );
  OAI21_X1 U4857 ( .B1(n7851), .B2(n4836), .A(n4833), .ZN(n7992) );
  NAND2_X1 U4858 ( .A1(n6063), .A2(n6062), .ZN(n8983) );
  NAND2_X1 U4859 ( .A1(n7262), .A2(n5294), .ZN(n4621) );
  NAND2_X1 U4860 ( .A1(n5495), .A2(n5494), .ZN(n9438) );
  AND2_X1 U4861 ( .A1(n7557), .A2(n7556), .ZN(n7827) );
  NAND2_X1 U4862 ( .A1(n7784), .A2(n4832), .ZN(n10008) );
  NAND2_X1 U4863 ( .A1(n6037), .A2(n6036), .ZN(n8993) );
  OAI21_X1 U4864 ( .B1(n5493), .B2(n4966), .A(n4965), .ZN(n5511) );
  OAI21_X1 U4865 ( .B1(n7552), .B2(n7551), .A(n7550), .ZN(n9558) );
  NAND2_X1 U4866 ( .A1(n5473), .A2(n5472), .ZN(n9442) );
  NAND2_X1 U4867 ( .A1(n5455), .A2(n5454), .ZN(n9447) );
  NAND2_X1 U4868 ( .A1(n6011), .A2(n6010), .ZN(n9005) );
  NAND2_X1 U4869 ( .A1(n6025), .A2(n6024), .ZN(n9002) );
  OR2_X1 U4870 ( .A1(n9458), .A2(n8037), .ZN(n8032) );
  OAI21_X1 U4871 ( .B1(n4949), .B2(n5435), .A(n4731), .ZN(n5453) );
  NAND2_X1 U4872 ( .A1(n5391), .A2(n5390), .ZN(n7912) );
  NAND2_X1 U4873 ( .A1(n5412), .A2(n5411), .ZN(n9465) );
  NAND2_X1 U4874 ( .A1(n5995), .A2(n5994), .ZN(n9012) );
  AOI21_X1 U4875 ( .B1(n8481), .B2(n4690), .A(n4305), .ZN(n8402) );
  NOR2_X1 U4876 ( .A1(n7858), .A2(n7887), .ZN(n7859) );
  NAND2_X1 U4877 ( .A1(n6201), .A2(n6198), .ZN(n8593) );
  NAND2_X1 U4878 ( .A1(n8372), .A2(n8482), .ZN(n8481) );
  OR2_X1 U4879 ( .A1(n5364), .A2(n4925), .ZN(n4295) );
  AND2_X1 U4880 ( .A1(n6503), .A2(n7165), .ZN(n7194) );
  NAND2_X1 U4881 ( .A1(n5879), .A2(n5878), .ZN(n7887) );
  NOR2_X1 U4882 ( .A1(n9772), .A2(n7116), .ZN(n9773) );
  INV_X1 U4883 ( .A(n7106), .ZN(n9849) );
  OR2_X1 U4884 ( .A1(n7295), .A2(n7294), .ZN(n9772) );
  NAND2_X1 U4885 ( .A1(n4430), .A2(n4429), .ZN(n5318) );
  AND2_X1 U4886 ( .A1(n8137), .A2(n8128), .ZN(n9919) );
  XNOR2_X1 U4887 ( .A(n4552), .B(n5232), .ZN(n6655) );
  INV_X1 U4888 ( .A(n9161), .ZN(n6307) );
  INV_X1 U4889 ( .A(n9158), .ZN(n5181) );
  AND2_X1 U4890 ( .A1(n5139), .A2(n5138), .ZN(n9783) );
  AND3_X2 U4891 ( .A1(n5134), .A2(n5133), .A3(n5132), .ZN(n9823) );
  INV_X1 U4892 ( .A(n7779), .ZN(n8613) );
  AND2_X2 U4893 ( .A1(n5752), .A2(n8089), .ZN(n6108) );
  NAND2_X1 U4894 ( .A1(n8123), .A2(n8122), .ZN(n8257) );
  NAND4_X1 U4895 ( .A1(n5796), .A2(n5795), .A3(n5794), .A4(n5793), .ZN(n8619)
         );
  NAND2_X1 U4896 ( .A1(n4623), .A2(n4624), .ZN(n5254) );
  NAND3_X1 U4897 ( .A1(n5073), .A2(n5072), .A3(n5071), .ZN(n9815) );
  INV_X1 U4898 ( .A(n9932), .ZN(n9966) );
  NAND4_X1 U4899 ( .A1(n5170), .A2(n5169), .A3(n5168), .A4(n5167), .ZN(n9158)
         );
  AND4_X1 U4900 ( .A1(n5859), .A2(n5858), .A3(n5857), .A4(n5856), .ZN(n7726)
         );
  OAI21_X1 U4901 ( .B1(n5110), .B2(n6864), .A(n4649), .ZN(n4648) );
  AND4_X1 U4902 ( .A1(n6918), .A2(n6916), .A3(n6917), .A4(n6915), .ZN(n8413)
         );
  OAI211_X1 U4903 ( .C1(n6286), .C2(n7006), .A(n5785), .B(n5784), .ZN(n9932)
         );
  AND4_X1 U4904 ( .A1(n6923), .A2(n6925), .A3(n6924), .A4(n6922), .ZN(n8425)
         );
  AND4_X1 U4905 ( .A1(n5769), .A2(n5768), .A3(n5767), .A4(n5766), .ZN(n7072)
         );
  CLKBUF_X1 U4906 ( .A(n5631), .Z(n7648) );
  OAI21_X1 U4907 ( .B1(n4409), .B2(n4408), .A(n4406), .ZN(n5172) );
  XNOR2_X1 U4908 ( .A(n5048), .B(n5047), .ZN(n5631) );
  NAND2_X1 U4909 ( .A1(n5012), .A2(n5637), .ZN(n6568) );
  NAND2_X1 U4910 ( .A1(n5046), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5048) );
  NOR2_X1 U4911 ( .A1(n7941), .A2(n7896), .ZN(n5012) );
  NAND2_X1 U4912 ( .A1(n5632), .A2(n5658), .ZN(n5064) );
  INV_X2 U4913 ( .A(n5241), .ZN(n5446) );
  NAND2_X1 U4914 ( .A1(n4478), .A2(n4476), .ZN(n8414) );
  OR2_X1 U4915 ( .A1(n4879), .A2(n5129), .ZN(n4880) );
  MUX2_X1 U4916 ( .A(P2_IR_REG_0__SCAN_IN), .B(n9052), .S(n6286), .Z(n9952) );
  NAND2_X1 U4917 ( .A1(n6286), .A2(n4873), .ZN(n5797) );
  AND2_X1 U4918 ( .A1(n5658), .A2(n9298), .ZN(n5663) );
  NAND2_X2 U4919 ( .A1(n5035), .A2(n9499), .ZN(n5111) );
  NAND2_X4 U4920 ( .A1(n6286), .A2(n4283), .ZN(n6082) );
  XNOR2_X1 U4921 ( .A(n5037), .B(n5036), .ZN(n8389) );
  XNOR2_X1 U4922 ( .A(n5034), .B(n5033), .ZN(n9499) );
  MUX2_X1 U4923 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5729), .S(
        P2_IR_REG_29__SCAN_IN), .Z(n5732) );
  NAND2_X1 U4925 ( .A1(n4998), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5045) );
  OR2_X1 U4926 ( .A1(n9492), .A2(n9493), .ZN(n5037) );
  XNOR2_X1 U4927 ( .A(n5050), .B(P1_IR_REG_19__SCAN_IN), .ZN(n9757) );
  OR2_X1 U4928 ( .A1(n5753), .A2(n5728), .ZN(n4387) );
  XNOR2_X1 U4929 ( .A(n5756), .B(n5755), .ZN(n8264) );
  CLKBUF_X1 U4930 ( .A(n5737), .Z(n6008) );
  INV_X2 U4931 ( .A(n8053), .ZN(n4282) );
  AND2_X1 U4932 ( .A1(n5721), .A2(n5991), .ZN(n5722) );
  AND2_X1 U4933 ( .A1(n4984), .A2(n4981), .ZN(n4684) );
  AND2_X1 U4934 ( .A1(n4805), .A2(n4721), .ZN(n4720) );
  NOR2_X1 U4935 ( .A1(n4983), .A2(P1_IR_REG_13__SCAN_IN), .ZN(n4984) );
  NOR2_X1 U4936 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(n5975), .ZN(n5991) );
  AND3_X1 U4937 ( .A1(n4717), .A2(n4716), .A3(n4715), .ZN(n5718) );
  AND2_X1 U4938 ( .A1(n5719), .A2(n4723), .ZN(n4721) );
  AND3_X1 U4939 ( .A1(n5746), .A2(n5738), .A3(n5748), .ZN(n5726) );
  AND4_X1 U4940 ( .A1(n5007), .A2(n5006), .A3(n5437), .A4(n5047), .ZN(n4301)
         );
  INV_X1 U4941 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5211) );
  INV_X1 U4942 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n8307) );
  INV_X1 U4943 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5946) );
  INV_X1 U4944 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5437) );
  INV_X1 U4945 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n4981) );
  INV_X1 U4946 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5029) );
  NOR2_X2 U4947 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n5068) );
  INV_X1 U4948 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5047) );
  INV_X1 U4949 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5003) );
  NOR2_X1 U4950 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n4975) );
  INV_X1 U4951 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5386) );
  NOR2_X1 U4952 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n4386) );
  INV_X1 U4953 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5738) );
  INV_X1 U4954 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5748) );
  INV_X1 U4955 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5746) );
  AND2_X1 U4956 ( .A1(n7176), .A2(n7011), .ZN(n7013) );
  OAI222_X1 U4957 ( .A1(n9502), .A2(n6642), .B1(n4282), .B2(n6641), .C1(
        P1_U3084), .C2(n9635), .ZN(P1_U3347) );
  OAI222_X1 U4958 ( .A1(n9041), .A2(n6639), .B1(n9049), .B2(n6641), .C1(
        P2_U3152), .C2(n6946), .ZN(P2_U3352) );
  XNOR2_X1 U4959 ( .A(n5750), .B(P2_IR_REG_19__SCAN_IN), .ZN(n8088) );
  NAND2_X1 U4960 ( .A1(n5700), .A2(n5051), .ZN(n4285) );
  INV_X2 U4961 ( .A(n6414), .ZN(n4287) );
  INV_X1 U4962 ( .A(n6414), .ZN(n5213) );
  OAI21_X2 U4963 ( .B1(n9101), .B2(n9100), .A(n9099), .ZN(n9098) );
  NAND2_X4 U4964 ( .A1(n6206), .A2(n8264), .ZN(n6286) );
  OAI222_X1 U4965 ( .A1(n9047), .A2(n8461), .B1(P2_U3152), .B2(n6206), .C1(
        n9049), .C2(n8460), .ZN(P2_U3330) );
  XNOR2_X2 U4966 ( .A(n4387), .B(n5754), .ZN(n6206) );
  AOI21_X2 U4967 ( .B1(n9092), .B2(n5574), .A(n4319), .ZN(n9134) );
  NOR2_X2 U4968 ( .A1(n4434), .A2(n9054), .ZN(n9092) );
  INV_X1 U4969 ( .A(n5237), .ZN(n4288) );
  INV_X2 U4970 ( .A(n5237), .ZN(n4289) );
  NAND2_X1 U4971 ( .A1(n8389), .A2(n9499), .ZN(n5241) );
  XNOR2_X2 U4972 ( .A(n4994), .B(P1_IR_REG_28__SCAN_IN), .ZN(n5671) );
  AOI21_X1 U4973 ( .B1(n8582), .B2(n4708), .A(n4705), .ZN(n4704) );
  INV_X1 U4974 ( .A(n8462), .ZN(n4705) );
  AND2_X1 U4975 ( .A1(n5735), .A2(n5736), .ZN(n5806) );
  NAND2_X1 U4976 ( .A1(n9109), .A2(n9112), .ZN(n4435) );
  NAND2_X1 U4977 ( .A1(n4742), .A2(n4741), .ZN(n6396) );
  AOI21_X1 U4978 ( .B1(n4744), .B2(n4746), .A(n4372), .ZN(n4741) );
  NAND2_X1 U4979 ( .A1(n5691), .A2(n4744), .ZN(n4742) );
  NOR2_X1 U4981 ( .A1(n4540), .A2(n4539), .ZN(n4538) );
  OAI22_X1 U4982 ( .A1(n6376), .A2(n9412), .B1(n6418), .B2(n6368), .ZN(n6369)
         );
  AND2_X1 U4983 ( .A1(n8238), .A2(n8237), .ZN(n4533) );
  NOR2_X1 U4984 ( .A1(n8911), .A2(n8877), .ZN(n8191) );
  AND2_X1 U4985 ( .A1(n4731), .A2(n4730), .ZN(n4729) );
  INV_X1 U4986 ( .A(n4935), .ZN(n4749) );
  INV_X1 U4987 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n4937) );
  INV_X1 U4988 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n4936) );
  INV_X1 U4989 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n4929) );
  AND2_X1 U4990 ( .A1(n5851), .A2(n5832), .ZN(n4714) );
  NOR2_X1 U4991 ( .A1(n7883), .A2(n4412), .ZN(n5893) );
  INV_X1 U4992 ( .A(n7758), .ZN(n4412) );
  OR2_X1 U4993 ( .A1(n8966), .A2(n8745), .ZN(n8228) );
  AND2_X1 U4994 ( .A1(n8228), .A2(n8229), .ZN(n8437) );
  NAND2_X1 U4995 ( .A1(n8798), .A2(n8075), .ZN(n4418) );
  NOR2_X1 U4996 ( .A1(n9012), .A2(n8850), .ZN(n4824) );
  AND2_X1 U4997 ( .A1(n8875), .A2(n4422), .ZN(n4421) );
  AOI21_X1 U4998 ( .B1(n9938), .B2(n9949), .A(n9951), .ZN(n7515) );
  AND2_X1 U4999 ( .A1(n6189), .A2(n6188), .ZN(n6209) );
  OR2_X1 U5000 ( .A1(n6237), .A2(n6238), .ZN(n6189) );
  AND2_X1 U5001 ( .A1(n5740), .A2(n5742), .ZN(n4724) );
  INV_X1 U5002 ( .A(n7652), .ZN(n5338) );
  INV_X1 U5003 ( .A(n9499), .ZN(n5038) );
  OR2_X1 U5004 ( .A1(n9401), .A2(n9245), .ZN(n9200) );
  OR2_X1 U5005 ( .A1(n9248), .A2(n9267), .ZN(n9199) );
  AND2_X1 U5006 ( .A1(n4293), .A2(n4325), .ZN(n4773) );
  NOR2_X1 U5007 ( .A1(n9180), .A2(n4778), .ZN(n4777) );
  INV_X1 U5008 ( .A(n4842), .ZN(n4778) );
  NAND2_X1 U5009 ( .A1(n7294), .A2(n9783), .ZN(n6441) );
  INV_X1 U5010 ( .A(n9823), .ZN(n7294) );
  INV_X1 U5011 ( .A(n5528), .ZN(n4755) );
  NAND2_X1 U5012 ( .A1(n4295), .A2(n4315), .ZN(n5385) );
  OAI21_X1 U5013 ( .B1(n5318), .B2(n5317), .A(n4917), .ZN(n5343) );
  INV_X1 U5014 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n4977) );
  NAND2_X1 U5015 ( .A1(n4410), .A2(n6079), .ZN(n6101) );
  INV_X1 U5016 ( .A(n4701), .ZN(n4698) );
  AOI21_X1 U5017 ( .B1(n4701), .B2(n4703), .A(n6200), .ZN(n4700) );
  NOR2_X1 U5018 ( .A1(n6208), .A2(n9939), .ZN(n6201) );
  NOR2_X1 U5019 ( .A1(n4302), .A2(n8082), .ZN(n4602) );
  INV_X1 U5020 ( .A(n4526), .ZN(n4525) );
  NAND2_X1 U5021 ( .A1(n4504), .A2(n4503), .ZN(n4502) );
  INV_X1 U5022 ( .A(n6986), .ZN(n4503) );
  NAND2_X1 U5023 ( .A1(n4808), .A2(n4807), .ZN(n8671) );
  AOI21_X1 U5024 ( .B1(n4809), .B2(n4811), .A(n4348), .ZN(n4807) );
  AND3_X1 U5025 ( .A1(n6151), .A2(n6150), .A3(n6149), .ZN(n8694) );
  XNOR2_X1 U5026 ( .A(n8957), .B(n8586), .ZN(n8690) );
  AND4_X1 U5027 ( .A1(n6089), .A2(n6088), .A3(n6087), .A4(n6086), .ZN(n8756)
         );
  NAND2_X1 U5028 ( .A1(n4817), .A2(n4304), .ZN(n4816) );
  NAND2_X1 U5029 ( .A1(n4820), .A2(n4821), .ZN(n4814) );
  NOR2_X1 U5030 ( .A1(n8778), .A2(n4823), .ZN(n4820) );
  OR2_X1 U5031 ( .A1(n8927), .A2(n8904), .ZN(n8900) );
  INV_X1 U5032 ( .A(n6082), .ZN(n6023) );
  NAND2_X1 U5033 ( .A1(n9990), .A2(n7703), .ZN(n7706) );
  NAND2_X1 U5034 ( .A1(n4355), .A2(n4298), .ZN(n4828) );
  AND2_X1 U5035 ( .A1(n6185), .A2(n9938), .ZN(n7519) );
  NAND2_X1 U5036 ( .A1(n6143), .A2(n6142), .ZN(n8950) );
  AND2_X1 U5037 ( .A1(n8122), .A2(n8133), .ZN(n9953) );
  NAND2_X1 U5038 ( .A1(n5733), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5734) );
  AND2_X1 U5039 ( .A1(n5929), .A2(n4837), .ZN(n5731) );
  NOR2_X1 U5040 ( .A1(n4838), .A2(n4299), .ZN(n4837) );
  NAND2_X1 U5041 ( .A1(n5722), .A2(n5754), .ZN(n4838) );
  NAND4_X1 U5042 ( .A1(n4720), .A2(n5722), .A3(n4803), .A4(n4486), .ZN(n6171)
         );
  INV_X1 U5043 ( .A(n5727), .ZN(n4486) );
  INV_X1 U5044 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4725) );
  INV_X1 U5045 ( .A(n9153), .ZN(n9561) );
  INV_X1 U5046 ( .A(n5341), .ZN(n4635) );
  AND2_X1 U5047 ( .A1(n4433), .A2(n4432), .ZN(n9054) );
  OR2_X1 U5048 ( .A1(n9412), .A2(n9284), .ZN(n9181) );
  OR2_X1 U5049 ( .A1(n9432), .A2(n9346), .ZN(n9178) );
  NOR2_X1 U5050 ( .A1(n9084), .A2(n8037), .ZN(n8038) );
  AND4_X1 U5051 ( .A1(n5421), .A2(n5420), .A3(n5419), .A4(n5418), .ZN(n7982)
         );
  NAND2_X1 U5052 ( .A1(n4274), .A2(n4873), .ZN(n6414) );
  INV_X1 U5053 ( .A(n9781), .ZN(n9736) );
  NAND2_X1 U5054 ( .A1(n7020), .A2(n7019), .ZN(n9786) );
  NAND2_X1 U5055 ( .A1(n5604), .A2(n5603), .ZN(n5691) );
  NAND2_X1 U5056 ( .A1(n6081), .A2(n6080), .ZN(n8975) );
  NAND2_X1 U5057 ( .A1(n4444), .A2(n4443), .ZN(n4442) );
  NOR2_X1 U5058 ( .A1(n5703), .A2(n9131), .ZN(n4443) );
  INV_X1 U5059 ( .A(n5704), .ZN(n4444) );
  NAND2_X1 U5060 ( .A1(n4381), .A2(n4844), .ZN(n8162) );
  NOR2_X1 U5061 ( .A1(n4549), .A2(n8257), .ZN(n4548) );
  INV_X1 U5062 ( .A(n8178), .ZN(n4549) );
  NAND2_X1 U5063 ( .A1(n4392), .A2(n4543), .ZN(n4391) );
  NOR2_X1 U5064 ( .A1(n8879), .A2(n8192), .ZN(n4543) );
  NAND2_X1 U5065 ( .A1(n4393), .A2(n4544), .ZN(n4392) );
  NAND2_X1 U5066 ( .A1(n8892), .A2(n4542), .ZN(n4541) );
  NOR2_X1 U5067 ( .A1(n8127), .A2(n8906), .ZN(n4542) );
  AOI21_X1 U5068 ( .B1(n4308), .B2(n4291), .A(n4536), .ZN(n4535) );
  INV_X1 U5069 ( .A(n8221), .ZN(n8222) );
  OAI21_X1 U5070 ( .B1(n8217), .B2(n4378), .A(n8076), .ZN(n4377) );
  NAND2_X1 U5071 ( .A1(n8214), .A2(n4379), .ZN(n4378) );
  NOR2_X1 U5072 ( .A1(n8216), .A2(n8257), .ZN(n4379) );
  MUX2_X1 U5073 ( .A(n6374), .B(n6373), .S(n6430), .Z(n6375) );
  INV_X1 U5074 ( .A(n4660), .ZN(n4659) );
  OAI21_X1 U5075 ( .B1(n8041), .B2(n4661), .A(n9378), .ZN(n4660) );
  NAND2_X1 U5076 ( .A1(n6524), .A2(n6522), .ZN(n7109) );
  INV_X1 U5077 ( .A(SI_16_), .ZN(n4938) );
  AOI21_X1 U5078 ( .B1(n4904), .B2(n4903), .A(n4419), .ZN(n4740) );
  NAND2_X1 U5079 ( .A1(n4906), .A2(n4905), .ZN(n4909) );
  INV_X1 U5080 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n4976) );
  NAND2_X1 U5081 ( .A1(n4397), .A2(n4400), .ZN(n4395) );
  NAND2_X1 U5082 ( .A1(n5895), .A2(n4335), .ZN(n4416) );
  NAND2_X1 U5083 ( .A1(n7934), .A2(n5960), .ZN(n5965) );
  OAI21_X1 U5084 ( .B1(n4529), .B2(n4297), .A(n4527), .ZN(n8254) );
  INV_X1 U5085 ( .A(n4528), .ZN(n4527) );
  OAI21_X1 U5086 ( .B1(n4322), .B2(n4297), .A(n8253), .ZN(n4528) );
  NAND2_X1 U5087 ( .A1(n4481), .A2(n4480), .ZN(n4479) );
  NOR2_X1 U5088 ( .A1(n4596), .A2(n4595), .ZN(n4594) );
  OR2_X1 U5089 ( .A1(n4597), .A2(n4595), .ZN(n4592) );
  NOR2_X1 U5090 ( .A1(n7852), .A2(n4598), .ZN(n4597) );
  INV_X1 U5091 ( .A(n8173), .ZN(n4598) );
  NAND2_X1 U5092 ( .A1(n7727), .A2(n9972), .ZN(n4831) );
  AND2_X1 U5093 ( .A1(n4298), .A2(n8091), .ZN(n4830) );
  OAI211_X1 U5094 ( .C1(n4431), .C2(n4606), .A(n4604), .B(n8070), .ZN(n8826)
         );
  INV_X1 U5095 ( .A(n4314), .ZN(n4431) );
  NAND2_X1 U5096 ( .A1(n6163), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6187) );
  INV_X1 U5097 ( .A(n8310), .ZN(n4447) );
  NAND2_X1 U5098 ( .A1(n6421), .A2(n4852), .ZN(n6422) );
  NOR2_X1 U5099 ( .A1(n9653), .A2(n8277), .ZN(n8278) );
  OR2_X1 U5100 ( .A1(n9412), .A2(n6472), .ZN(n9198) );
  AND2_X1 U5101 ( .A1(n9280), .A2(n9293), .ZN(n9194) );
  AND2_X1 U5102 ( .A1(n4325), .A2(n4776), .ZN(n4772) );
  NOR2_X1 U5103 ( .A1(n9175), .A2(n4790), .ZN(n4789) );
  INV_X1 U5104 ( .A(n4792), .ZN(n4790) );
  INV_X1 U5105 ( .A(n7978), .ZN(n4678) );
  AND2_X1 U5106 ( .A1(n7914), .A2(n4801), .ZN(n4799) );
  AND2_X1 U5107 ( .A1(n7837), .A2(n7825), .ZN(n4682) );
  INV_X1 U5108 ( .A(n7827), .ZN(n4681) );
  INV_X1 U5109 ( .A(n7200), .ZN(n4783) );
  OR2_X1 U5110 ( .A1(n6314), .A2(n8315), .ZN(n6503) );
  NOR2_X1 U5111 ( .A1(n7284), .A2(n7106), .ZN(n4575) );
  NAND2_X1 U5112 ( .A1(n7315), .A2(n7106), .ZN(n7163) );
  OAI21_X1 U5113 ( .B1(n6396), .B2(n6395), .A(n6394), .ZN(n6409) );
  NAND2_X1 U5114 ( .A1(n4764), .A2(n4762), .ZN(n5602) );
  AOI21_X1 U5115 ( .B1(n4765), .B2(n4767), .A(n4763), .ZN(n4762) );
  INV_X1 U5116 ( .A(n5575), .ZN(n4763) );
  AND3_X1 U5117 ( .A1(n5652), .A2(n4985), .A3(n5029), .ZN(n4989) );
  NOR2_X1 U5118 ( .A1(n4757), .A2(n4752), .ZN(n4751) );
  INV_X1 U5119 ( .A(n4961), .ZN(n4752) );
  INV_X1 U5120 ( .A(n4758), .ZN(n4757) );
  INV_X1 U5121 ( .A(n4760), .ZN(n4756) );
  NAND2_X1 U5122 ( .A1(n4728), .A2(n4726), .ZN(n5471) );
  AND2_X1 U5123 ( .A1(n4727), .A2(n4957), .ZN(n4726) );
  AND2_X1 U5124 ( .A1(n4961), .A2(n4960), .ZN(n5470) );
  INV_X1 U5125 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n4952) );
  INV_X1 U5126 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n4982) );
  INV_X1 U5127 ( .A(SI_15_), .ZN(n4930) );
  NAND2_X1 U5128 ( .A1(n4976), .A2(n4786), .ZN(n4785) );
  INV_X1 U5129 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n4786) );
  AND2_X1 U5130 ( .A1(n4735), .A2(n4912), .ZN(n4429) );
  NAND2_X1 U5131 ( .A1(n4347), .A2(n5254), .ZN(n4430) );
  AOI21_X1 U5132 ( .B1(n4740), .B2(n4738), .A(n4737), .ZN(n4736) );
  INV_X1 U5133 ( .A(n4909), .ZN(n4737) );
  INV_X1 U5134 ( .A(n4903), .ZN(n4738) );
  INV_X1 U5135 ( .A(n4740), .ZN(n4739) );
  OR2_X1 U5136 ( .A1(n5252), .A2(n4902), .ZN(n4904) );
  NAND2_X1 U5137 ( .A1(n5881), .A2(n5880), .ZN(n5900) );
  NAND2_X1 U5138 ( .A1(n5806), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n6924) );
  NOR2_X1 U5139 ( .A1(n8553), .A2(n4713), .ZN(n4712) );
  INV_X1 U5140 ( .A(n6035), .ZN(n4713) );
  AOI21_X1 U5141 ( .B1(n4416), .B2(n4415), .A(n4375), .ZN(n4688) );
  NAND2_X1 U5142 ( .A1(n5895), .A2(n7600), .ZN(n4415) );
  INV_X1 U5143 ( .A(n4416), .ZN(n4689) );
  OR2_X1 U5144 ( .A1(n8523), .A2(n8524), .ZN(n8521) );
  AND2_X1 U5145 ( .A1(n7344), .A2(n5803), .ZN(n4691) );
  NAND2_X1 U5146 ( .A1(n5965), .A2(n5964), .ZN(n5966) );
  OR2_X1 U5147 ( .A1(n5965), .A2(n5964), .ZN(n5974) );
  AND3_X1 U5148 ( .A1(n6138), .A2(n6137), .A3(n6136), .ZN(n8586) );
  AND4_X1 U5149 ( .A1(n5875), .A2(n5874), .A3(n5873), .A4(n5872), .ZN(n7779)
         );
  NAND2_X1 U5150 ( .A1(n6217), .A2(n4489), .ZN(n4488) );
  INV_X1 U5151 ( .A(n9507), .ZN(n4489) );
  AOI21_X1 U5152 ( .B1(n6248), .B2(P2_REG2_REG_7__SCAN_IN), .A(n6961), .ZN(
        n6837) );
  NAND2_X1 U5153 ( .A1(n6659), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n4495) );
  NAND2_X1 U5154 ( .A1(n4310), .A2(n4518), .ZN(n4514) );
  NAND2_X1 U5155 ( .A1(n4310), .A2(n4516), .ZN(n4515) );
  INV_X1 U5156 ( .A(n7232), .ZN(n4516) );
  NAND2_X1 U5157 ( .A1(n4513), .A2(n4511), .ZN(n7744) );
  AOI21_X1 U5158 ( .B1(n4515), .B2(n4514), .A(n4512), .ZN(n4511) );
  NAND2_X1 U5159 ( .A1(n6227), .A2(n4514), .ZN(n4513) );
  INV_X1 U5160 ( .A(n7745), .ZN(n4512) );
  XNOR2_X1 U5161 ( .A(n4490), .B(n6235), .ZN(n6284) );
  NAND2_X1 U5162 ( .A1(n8650), .A2(n6234), .ZN(n4490) );
  NAND2_X1 U5163 ( .A1(n8244), .A2(n8251), .ZN(n8447) );
  INV_X1 U5164 ( .A(n8447), .ZN(n8441) );
  AND3_X1 U5165 ( .A1(n6129), .A2(n6128), .A3(n6127), .ZN(n8693) );
  OR2_X1 U5166 ( .A1(n8961), .A2(n8606), .ZN(n8439) );
  INV_X1 U5167 ( .A(n4810), .ZN(n4809) );
  OAI21_X1 U5168 ( .B1(n8705), .B2(n4811), .A(n8690), .ZN(n4810) );
  INV_X1 U5169 ( .A(n8439), .ZN(n4811) );
  AND2_X1 U5170 ( .A1(n8437), .A2(n4609), .ZN(n4608) );
  AND2_X1 U5171 ( .A1(n8078), .A2(n8437), .ZN(n4610) );
  INV_X1 U5172 ( .A(n8710), .ZN(n8705) );
  NAND2_X1 U5173 ( .A1(n8706), .A2(n8705), .ZN(n8704) );
  NOR2_X1 U5174 ( .A1(n8763), .A2(n4479), .ZN(n8725) );
  INV_X1 U5175 ( .A(n8437), .ZN(n8728) );
  NAND2_X1 U5176 ( .A1(n8755), .A2(n8078), .ZN(n8740) );
  NOR2_X1 U5177 ( .A1(n8763), .A2(n8970), .ZN(n8451) );
  AOI21_X1 U5178 ( .B1(n4823), .B2(n8858), .A(n4341), .ZN(n4821) );
  OR2_X1 U5179 ( .A1(n8993), .A2(n8833), .ZN(n8212) );
  INV_X1 U5180 ( .A(n8090), .ZN(n8817) );
  INV_X1 U5181 ( .A(n4824), .ZN(n4822) );
  NAND2_X1 U5182 ( .A1(n4817), .A2(n4826), .ZN(n4825) );
  AND4_X1 U5183 ( .A1(n5973), .A2(n5972), .A3(n5971), .A4(n5970), .ZN(n8877)
         );
  NAND2_X1 U5184 ( .A1(n6749), .A2(n8084), .ZN(n4417) );
  AOI21_X1 U5185 ( .B1(n4835), .B2(n4834), .A(n4307), .ZN(n4833) );
  NAND2_X1 U5186 ( .A1(n7851), .A2(n8102), .ZN(n7990) );
  NAND2_X1 U5187 ( .A1(n7704), .A2(n4596), .ZN(n7784) );
  AND2_X1 U5188 ( .A1(n8120), .A2(n8089), .ZN(n8920) );
  OR2_X1 U5189 ( .A1(n6912), .A2(n6206), .ZN(n8905) );
  INV_X1 U5190 ( .A(n7519), .ZN(n7517) );
  INV_X1 U5191 ( .A(n8862), .ZN(n8907) );
  INV_X1 U5192 ( .A(n8920), .ZN(n9922) );
  NOR2_X1 U5193 ( .A1(n8948), .A2(n4365), .ZN(n4484) );
  INV_X1 U5194 ( .A(n9913), .ZN(n10004) );
  AND2_X1 U5195 ( .A1(n6909), .A2(n6908), .ZN(n6933) );
  NAND2_X1 U5196 ( .A1(n6209), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9939) );
  AND2_X1 U5197 ( .A1(n6173), .A2(n6186), .ZN(n9938) );
  OR2_X1 U5198 ( .A1(n7943), .A2(n6168), .ZN(n6173) );
  INV_X1 U5199 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n6158) );
  NOR2_X1 U5200 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n5740) );
  NAND2_X1 U5201 ( .A1(n5745), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5750) );
  NOR2_X2 U5202 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5757) );
  NAND2_X1 U5203 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n4498) );
  NAND2_X1 U5204 ( .A1(n4436), .A2(n4435), .ZN(n9053) );
  CLKBUF_X1 U5205 ( .A(n5171), .Z(n5451) );
  INV_X1 U5206 ( .A(n9121), .ZN(n4639) );
  OR2_X1 U5207 ( .A1(n5535), .A2(n5534), .ZN(n5562) );
  NAND2_X1 U5208 ( .A1(n5018), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5349) );
  INV_X1 U5209 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5348) );
  OR2_X1 U5210 ( .A1(n5349), .A2(n5348), .ZN(n5370) );
  OR2_X1 U5211 ( .A1(n5497), .A2(n5496), .ZN(n5514) );
  NAND2_X1 U5212 ( .A1(n5136), .A2(n5135), .ZN(n5137) );
  NAND2_X1 U5213 ( .A1(n4294), .A2(n4338), .ZN(n4642) );
  NOR2_X1 U5214 ( .A1(n4294), .A2(n4338), .ZN(n4641) );
  NAND2_X1 U5215 ( .A1(n4645), .A2(n4646), .ZN(n4647) );
  NAND2_X1 U5216 ( .A1(n4629), .A2(n4627), .ZN(n7960) );
  NAND2_X1 U5217 ( .A1(n4628), .A2(n4346), .ZN(n4627) );
  NOR2_X1 U5218 ( .A1(n7960), .A2(n7959), .ZN(n8020) );
  NAND2_X1 U5219 ( .A1(n5655), .A2(n6705), .ZN(n6708) );
  OAI21_X1 U5220 ( .B1(n6855), .B2(n5074), .A(n4455), .ZN(n6851) );
  NAND2_X1 U5221 ( .A1(n6855), .A2(n5074), .ZN(n4455) );
  NAND2_X1 U5222 ( .A1(n6850), .A2(n6851), .ZN(n6849) );
  NAND2_X1 U5223 ( .A1(n9622), .A2(n9623), .ZN(n9621) );
  NAND2_X1 U5224 ( .A1(n4454), .A2(n4453), .ZN(n8356) );
  INV_X1 U5225 ( .A(n8359), .ZN(n4453) );
  INV_X1 U5226 ( .A(n8358), .ZN(n4454) );
  NOR2_X1 U5227 ( .A1(n8349), .A2(n4466), .ZN(n8333) );
  AND2_X1 U5228 ( .A1(n6776), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4466) );
  NAND2_X1 U5229 ( .A1(n8333), .A2(n8332), .ZN(n8331) );
  OR2_X1 U5230 ( .A1(n6779), .A2(n6780), .ZN(n8273) );
  XNOR2_X1 U5231 ( .A(n8278), .B(n4465), .ZN(n9671) );
  INV_X1 U5232 ( .A(n9674), .ZN(n4465) );
  OR2_X1 U5233 ( .A1(n9671), .A2(n7843), .ZN(n4464) );
  NAND2_X1 U5234 ( .A1(n4586), .A2(n4585), .ZN(n4584) );
  INV_X1 U5235 ( .A(n9398), .ZN(n4586) );
  NAND2_X1 U5236 ( .A1(n9226), .A2(n4652), .ZN(n9205) );
  AND2_X1 U5237 ( .A1(n9204), .A2(n9203), .ZN(n4652) );
  NAND2_X1 U5238 ( .A1(n9269), .A2(n9198), .ZN(n9242) );
  OR2_X1 U5239 ( .A1(n4672), .A2(n9192), .ZN(n4669) );
  AND2_X1 U5240 ( .A1(n9312), .A2(n4674), .ZN(n4672) );
  NAND2_X1 U5241 ( .A1(n9327), .A2(n4670), .ZN(n4665) );
  AOI21_X1 U5242 ( .B1(n4669), .B2(n4671), .A(n4667), .ZN(n4666) );
  INV_X1 U5243 ( .A(n9291), .ZN(n4667) );
  INV_X1 U5244 ( .A(n4669), .ZN(n4668) );
  INV_X1 U5245 ( .A(n4777), .ZN(n4776) );
  NAND2_X1 U5246 ( .A1(n9307), .A2(n9179), .ZN(n4780) );
  NAND2_X1 U5247 ( .A1(n4777), .A2(n4775), .ZN(n4774) );
  INV_X1 U5248 ( .A(n9178), .ZN(n4775) );
  AND2_X1 U5249 ( .A1(n6494), .A2(n9193), .ZN(n9291) );
  NOR2_X1 U5250 ( .A1(n9352), .A2(n4791), .ZN(n9176) );
  AND2_X1 U5251 ( .A1(n9442), .A2(n9381), .ZN(n4791) );
  AND2_X1 U5252 ( .A1(n9453), .A2(n9380), .ZN(n4792) );
  OR2_X1 U5253 ( .A1(n5416), .A2(n5057), .ZN(n5444) );
  NOR2_X1 U5254 ( .A1(n8040), .A2(n8041), .ZN(n9173) );
  NAND2_X1 U5255 ( .A1(n8035), .A2(n8041), .ZN(n9186) );
  NAND2_X1 U5256 ( .A1(n7972), .A2(n7971), .ZN(n8039) );
  NAND2_X1 U5257 ( .A1(n9465), .A2(n9150), .ZN(n7971) );
  INV_X1 U5258 ( .A(n7836), .ZN(n4679) );
  NAND2_X1 U5259 ( .A1(n4681), .A2(n4682), .ZN(n4680) );
  NAND2_X1 U5260 ( .A1(n4680), .A2(n4296), .ZN(n7979) );
  NAND2_X1 U5261 ( .A1(n9588), .A2(n7963), .ZN(n4801) );
  AND2_X1 U5262 ( .A1(n7877), .A2(n9152), .ZN(n4802) );
  OR2_X1 U5263 ( .A1(n9592), .A2(n9561), .ZN(n4841) );
  OR2_X1 U5264 ( .A1(n7823), .A2(n9153), .ZN(n7821) );
  AND2_X1 U5265 ( .A1(n6500), .A2(n7825), .ZN(n7556) );
  NAND2_X1 U5266 ( .A1(n4783), .A2(n7156), .ZN(n7198) );
  NAND2_X1 U5267 ( .A1(n4656), .A2(n4655), .ZN(n4654) );
  AND2_X1 U5268 ( .A1(n6440), .A2(n6530), .ZN(n9738) );
  INV_X1 U5269 ( .A(n9786), .ZN(n9766) );
  NAND2_X1 U5270 ( .A1(n7289), .A2(n7288), .ZN(n4567) );
  OAI21_X2 U5271 ( .B1(n6414), .B2(n6621), .A(n4648), .ZN(n6305) );
  NAND2_X1 U5272 ( .A1(n4274), .A2(n4650), .ZN(n4649) );
  NAND2_X1 U5273 ( .A1(n4651), .A2(n4278), .ZN(n4650) );
  OR2_X1 U5274 ( .A1(n6708), .A2(n7024), .ZN(n9781) );
  INV_X1 U5275 ( .A(n9280), .ZN(n9417) );
  NOR3_X1 U5276 ( .A1(n6716), .A2(n6704), .A3(n6703), .ZN(n7015) );
  XNOR2_X1 U5277 ( .A(n6409), .B(n6408), .ZN(n6407) );
  NAND2_X1 U5278 ( .A1(n4324), .A2(n4301), .ZN(n5008) );
  XNOR2_X1 U5279 ( .A(n6396), .B(n6387), .ZN(n9046) );
  AND2_X1 U5280 ( .A1(n5692), .A2(n5608), .ZN(n5690) );
  XNOR2_X1 U5281 ( .A(n5011), .B(P1_IR_REG_26__SCAN_IN), .ZN(n5637) );
  XNOR2_X1 U5282 ( .A(n5577), .B(n5576), .ZN(n7940) );
  NOR2_X1 U5283 ( .A1(n5510), .A2(n4761), .ZN(n4760) );
  INV_X1 U5284 ( .A(n4965), .ZN(n4761) );
  AND2_X1 U5285 ( .A1(n5530), .A2(n4974), .ZN(n5528) );
  AOI21_X1 U5286 ( .B1(n4760), .B2(n4966), .A(n4759), .ZN(n4758) );
  INV_X1 U5287 ( .A(n4971), .ZN(n4759) );
  AND2_X1 U5288 ( .A1(n5209), .A2(n5173), .ZN(n4555) );
  NOR2_X1 U5289 ( .A1(n5252), .A2(n4625), .ZN(n4622) );
  OR2_X1 U5290 ( .A1(n5069), .A2(P1_IR_REG_2__SCAN_IN), .ZN(n5130) );
  NAND2_X1 U5291 ( .A1(n6133), .A2(n6132), .ZN(n8957) );
  NAND2_X1 U5292 ( .A1(n5950), .A2(n5949), .ZN(n8927) );
  AND4_X1 U5293 ( .A1(n5908), .A2(n5907), .A3(n5906), .A4(n5905), .ZN(n7904)
         );
  AOI21_X1 U5294 ( .B1(n4700), .B2(n4698), .A(n4696), .ZN(n4695) );
  OAI21_X1 U5295 ( .B1(n4698), .B2(n4697), .A(n6199), .ZN(n4696) );
  NAND2_X1 U5296 ( .A1(n4703), .A2(n6197), .ZN(n4697) );
  INV_X1 U5297 ( .A(n4700), .ZN(n4699) );
  AND4_X1 U5298 ( .A1(n5890), .A2(n5889), .A3(n5888), .A4(n5887), .ZN(n7889)
         );
  NAND2_X1 U5299 ( .A1(n6286), .A2(n4477), .ZN(n4476) );
  OAI21_X1 U5300 ( .B1(n6634), .B2(n4278), .A(n4309), .ZN(n4477) );
  INV_X1 U5301 ( .A(n10020), .ZN(n8002) );
  NAND2_X1 U5302 ( .A1(n6105), .A2(n6104), .ZN(n8518) );
  INV_X1 U5303 ( .A(n8519), .ZN(n4404) );
  AND2_X1 U5304 ( .A1(n8966), .A2(n8589), .ZN(n4402) );
  NAND2_X1 U5305 ( .A1(n5974), .A2(n4719), .ZN(n8523) );
  OR2_X1 U5306 ( .A1(n8593), .A2(n7043), .ZN(n8592) );
  NAND2_X1 U5307 ( .A1(n5828), .A2(n8392), .ZN(n8405) );
  AND4_X1 U5308 ( .A1(n5813), .A2(n5812), .A3(n5811), .A4(n5810), .ZN(n7079)
         );
  AND4_X1 U5309 ( .A1(n5841), .A2(n5840), .A3(n5839), .A4(n5838), .ZN(n8396)
         );
  NAND2_X1 U5310 ( .A1(n8418), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8585) );
  AND2_X1 U5311 ( .A1(n7496), .A2(n5751), .ZN(n8265) );
  INV_X1 U5312 ( .A(n8905), .ZN(n8861) );
  NAND2_X1 U5313 ( .A1(n4526), .A2(n8262), .ZN(n4428) );
  NAND2_X1 U5314 ( .A1(n4525), .A2(n8261), .ZN(n4524) );
  NAND2_X1 U5315 ( .A1(n4599), .A2(n8263), .ZN(n4427) );
  INV_X1 U5316 ( .A(n8122), .ZN(n8268) );
  NOR2_X1 U5317 ( .A1(n6949), .A2(n4493), .ZN(n6975) );
  NOR2_X1 U5318 ( .A1(n6958), .A2(n6215), .ZN(n4493) );
  NAND2_X1 U5319 ( .A1(n6264), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n4501) );
  NAND2_X1 U5320 ( .A1(n7061), .A2(n4494), .ZN(n7231) );
  OR2_X1 U5321 ( .A1(n6265), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n4494) );
  INV_X1 U5322 ( .A(n4722), .ZN(n5912) );
  NAND2_X1 U5323 ( .A1(n8086), .A2(n8085), .ZN(n8938) );
  AND2_X1 U5324 ( .A1(n5892), .A2(n4354), .ZN(n4550) );
  OR2_X1 U5325 ( .A1(n6655), .A2(n5797), .ZN(n4551) );
  AND3_X1 U5326 ( .A1(n5802), .A2(n5801), .A3(n5800), .ZN(n7531) );
  INV_X1 U5327 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5730) );
  NAND2_X1 U5328 ( .A1(n6171), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5756) );
  XNOR2_X1 U5329 ( .A(n6162), .B(n6161), .ZN(n8122) );
  AND2_X1 U5330 ( .A1(n4858), .A2(n5716), .ZN(n4440) );
  OAI21_X1 U5331 ( .B1(n4442), .B2(n4858), .A(n4345), .ZN(n4438) );
  AND3_X1 U5332 ( .A1(n5449), .A2(n5448), .A3(n5447), .ZN(n9083) );
  OR2_X1 U5333 ( .A1(n6655), .A2(n5108), .ZN(n5236) );
  NAND2_X1 U5334 ( .A1(n5513), .A2(n5512), .ZN(n9432) );
  INV_X1 U5335 ( .A(n9148), .ZN(n9129) );
  INV_X1 U5336 ( .A(n9083), .ZN(n9380) );
  OAI21_X1 U5337 ( .B1(n8306), .B2(n8305), .A(n8304), .ZN(n4457) );
  OAI21_X1 U5338 ( .B1(n8302), .B2(n9681), .A(n4462), .ZN(n4461) );
  OR2_X1 U5339 ( .A1(n8303), .A2(n9724), .ZN(n4462) );
  OAI21_X1 U5340 ( .B1(n9727), .B2(n8307), .A(n9065), .ZN(n4459) );
  NAND2_X1 U5341 ( .A1(n9231), .A2(n9230), .ZN(n9232) );
  NAND2_X1 U5342 ( .A1(n9237), .A2(n4796), .ZN(n9219) );
  AND2_X1 U5343 ( .A1(n9237), .A2(n9182), .ZN(n9220) );
  NAND2_X1 U5344 ( .A1(n9797), .A2(n9769), .ZN(n9387) );
  INV_X1 U5345 ( .A(n9569), .ZN(n9791) );
  OR2_X1 U5346 ( .A1(n9818), .A2(n5661), .ZN(n9792) );
  AND2_X1 U5347 ( .A1(n9797), .A2(n9753), .ZN(n9569) );
  NAND2_X1 U5348 ( .A1(n4384), .A2(n4382), .ZN(n8140) );
  NAND2_X1 U5349 ( .A1(n4385), .A2(n8257), .ZN(n4384) );
  NAND2_X1 U5350 ( .A1(n8142), .A2(n4860), .ZN(n4383) );
  AOI21_X1 U5351 ( .B1(n4380), .B2(n8156), .A(n8174), .ZN(n8160) );
  NAND2_X1 U5352 ( .A1(n8162), .A2(n4329), .ZN(n4380) );
  AND2_X1 U5353 ( .A1(n6320), .A2(n6499), .ZN(n4557) );
  INV_X1 U5354 ( .A(n4559), .ZN(n4558) );
  OAI21_X1 U5355 ( .B1(n7920), .B2(n6430), .A(n6322), .ZN(n4559) );
  NAND2_X1 U5356 ( .A1(n8181), .A2(n4546), .ZN(n4545) );
  AOI21_X1 U5357 ( .B1(n8176), .B2(n4548), .A(n4349), .ZN(n4547) );
  AND2_X1 U5358 ( .A1(n8180), .A2(n8257), .ZN(n4546) );
  NOR2_X1 U5359 ( .A1(n8189), .A2(n8902), .ZN(n4544) );
  NAND2_X1 U5360 ( .A1(n4391), .A2(n4541), .ZN(n8198) );
  NAND2_X1 U5361 ( .A1(n4538), .A2(n8208), .ZN(n4537) );
  AND2_X1 U5362 ( .A1(n8215), .A2(n8212), .ZN(n8205) );
  NOR2_X1 U5363 ( .A1(n6365), .A2(n6418), .ZN(n4570) );
  OAI21_X1 U5364 ( .B1(n6366), .B2(n6430), .A(n6469), .ZN(n4569) );
  NAND2_X1 U5365 ( .A1(n4376), .A2(n4856), .ZN(n8227) );
  OAI21_X1 U5366 ( .B1(n8223), .B2(n4377), .A(n8222), .ZN(n4376) );
  INV_X1 U5367 ( .A(n8250), .ZN(n4532) );
  NAND2_X1 U5368 ( .A1(n4533), .A2(n8239), .ZN(n4530) );
  NAND2_X1 U5369 ( .A1(n4351), .A2(n4633), .ZN(n4632) );
  NAND2_X1 U5370 ( .A1(n5405), .A2(n4634), .ZN(n4633) );
  INV_X1 U5371 ( .A(n5361), .ZN(n4634) );
  AND2_X1 U5372 ( .A1(n9163), .A2(n6428), .ZN(n6517) );
  INV_X1 U5373 ( .A(n5692), .ZN(n4746) );
  INV_X1 U5374 ( .A(n4745), .ZN(n4744) );
  OAI21_X1 U5375 ( .B1(n5690), .B2(n4746), .A(n6383), .ZN(n4745) );
  NOR2_X1 U5376 ( .A1(n5576), .A2(n4766), .ZN(n4765) );
  INV_X1 U5377 ( .A(n5553), .ZN(n4766) );
  INV_X1 U5378 ( .A(n5452), .ZN(n4730) );
  INV_X1 U5379 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n4944) );
  OAI21_X1 U5380 ( .B1(n4873), .B2(P2_DATAO_REG_10__SCAN_IN), .A(n4420), .ZN(
        n4906) );
  NAND2_X1 U5381 ( .A1(n4873), .A2(n6660), .ZN(n4420) );
  AOI21_X1 U5382 ( .B1(n4704), .B2(n4702), .A(n4353), .ZN(n4701) );
  INV_X1 U5383 ( .A(n4708), .ZN(n4702) );
  INV_X1 U5384 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n4521) );
  AOI21_X1 U5385 ( .B1(P2_REG2_REG_17__SCAN_IN), .B2(n6246), .A(n8637), .ZN(
        n6233) );
  OR2_X1 U5386 ( .A1(n8950), .A2(n8694), .ZN(n8242) );
  AND2_X1 U5387 ( .A1(n8242), .A2(n8241), .ZN(n8238) );
  INV_X1 U5388 ( .A(n8224), .ZN(n4609) );
  NOR2_X1 U5389 ( .A1(n9002), .A2(n8993), .ZN(n4474) );
  NAND2_X1 U5390 ( .A1(n8106), .A2(n8900), .ZN(n4423) );
  NOR2_X1 U5391 ( .A1(n8911), .A2(n4469), .ZN(n4468) );
  INV_X1 U5392 ( .A(n4470), .ZN(n4469) );
  NOR2_X1 U5393 ( .A1(n8927), .A2(n8426), .ZN(n4470) );
  NOR2_X1 U5394 ( .A1(n9911), .A2(n8002), .ZN(n8004) );
  OR2_X1 U5395 ( .A1(n5884), .A2(n5883), .ZN(n5886) );
  INV_X1 U5396 ( .A(n8126), .ZN(n8131) );
  NAND2_X1 U5397 ( .A1(n7567), .A2(n8618), .ZN(n8126) );
  NAND2_X1 U5398 ( .A1(n8413), .A2(n8414), .ZN(n8143) );
  NOR3_X1 U5399 ( .A1(n8763), .A2(n8961), .A3(n4479), .ZN(n8714) );
  NAND2_X1 U5400 ( .A1(n7859), .A2(n10013), .ZN(n9911) );
  OR2_X1 U5401 ( .A1(n8414), .A2(n9952), .ZN(n7615) );
  INV_X1 U5402 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5943) );
  INV_X1 U5403 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n4804) );
  NOR2_X1 U5404 ( .A1(n5798), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n5814) );
  INV_X1 U5405 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4614) );
  AOI21_X1 U5406 ( .B1(n9073), .B2(n4617), .A(n4339), .ZN(n4616) );
  INV_X1 U5407 ( .A(n9073), .ZN(n4618) );
  INV_X1 U5408 ( .A(n5491), .ZN(n4617) );
  NOR2_X1 U5409 ( .A1(n4632), .A2(n7653), .ZN(n4630) );
  INV_X1 U5410 ( .A(n4632), .ZN(n4628) );
  AND2_X1 U5411 ( .A1(n9417), .A2(n9266), .ZN(n9196) );
  NAND2_X1 U5412 ( .A1(n4580), .A2(n9325), .ZN(n4579) );
  NOR2_X1 U5413 ( .A1(n9438), .A2(n9442), .ZN(n4580) );
  NAND2_X1 U5414 ( .A1(n9187), .A2(n9185), .ZN(n4658) );
  OR2_X1 U5415 ( .A1(n4659), .A2(n9188), .ZN(n4657) );
  NOR2_X1 U5416 ( .A1(n7912), .A2(n7877), .ZN(n4572) );
  NAND2_X1 U5417 ( .A1(n5017), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5326) );
  INV_X1 U5418 ( .A(n5304), .ZN(n5017) );
  INV_X1 U5419 ( .A(n7109), .ZN(n7248) );
  NAND2_X1 U5420 ( .A1(n7110), .A2(n7109), .ZN(n7245) );
  INV_X1 U5421 ( .A(n6634), .ZN(n4651) );
  INV_X1 U5422 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5006) );
  AND2_X1 U5423 ( .A1(n5603), .A2(n5581), .ZN(n5601) );
  INV_X1 U5424 ( .A(n5550), .ZN(n4767) );
  XNOR2_X1 U5425 ( .A(n5045), .B(P1_IR_REG_21__SCAN_IN), .ZN(n5632) );
  INV_X1 U5426 ( .A(SI_19_), .ZN(n4953) );
  INV_X1 U5427 ( .A(n4748), .ZN(n4747) );
  OAI21_X1 U5428 ( .B1(n4315), .B2(n4749), .A(n5408), .ZN(n4748) );
  INV_X1 U5429 ( .A(n4884), .ZN(n4407) );
  INV_X1 U5430 ( .A(n5144), .ZN(n4784) );
  OAI21_X1 U5431 ( .B1(n4278), .B2(P1_DATAO_REG_3__SCAN_IN), .A(n4874), .ZN(
        n4878) );
  OR2_X1 U5432 ( .A1(n6131), .A2(n6130), .ZN(n4708) );
  INV_X1 U5433 ( .A(n4704), .ZN(n4703) );
  NOR2_X1 U5434 ( .A1(n8530), .A2(n4710), .ZN(n4709) );
  INV_X1 U5435 ( .A(n5990), .ZN(n4710) );
  OR2_X1 U5436 ( .A1(n6092), .A2(n8546), .ZN(n6111) );
  AND2_X1 U5437 ( .A1(n6031), .A2(n4395), .ZN(n4394) );
  NAND2_X1 U5438 ( .A1(n8521), .A2(n4397), .ZN(n4396) );
  OR2_X1 U5439 ( .A1(n5919), .A2(n5918), .ZN(n5933) );
  INV_X1 U5440 ( .A(n6007), .ZN(n4400) );
  AND2_X1 U5441 ( .A1(n8572), .A2(n4398), .ZN(n4397) );
  NAND2_X1 U5442 ( .A1(n4399), .A2(n6007), .ZN(n4398) );
  INV_X1 U5443 ( .A(n4709), .ZN(n4399) );
  NAND2_X1 U5444 ( .A1(n5966), .A2(n4364), .ZN(n4719) );
  OR3_X1 U5445 ( .A1(n5968), .A2(n7952), .A3(n5967), .ZN(n5982) );
  INV_X1 U5446 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n7952) );
  NAND2_X1 U5447 ( .A1(n4388), .A2(n7496), .ZN(n4526) );
  NAND2_X1 U5448 ( .A1(n4389), .A2(n8260), .ZN(n4388) );
  NAND2_X1 U5449 ( .A1(n4390), .A2(n8255), .ZN(n4389) );
  AND4_X1 U5450 ( .A1(n6061), .A2(n6060), .A3(n6059), .A4(n6058), .ZN(n8431)
         );
  NAND2_X1 U5451 ( .A1(n5792), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n6918) );
  NAND2_X1 U5452 ( .A1(n5806), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n6916) );
  NAND2_X1 U5453 ( .A1(n9509), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n4487) );
  NOR2_X1 U5454 ( .A1(n9519), .A2(n4321), .ZN(n9518) );
  OR2_X1 U5455 ( .A1(n6975), .A2(n6974), .ZN(n4492) );
  NAND2_X1 U5456 ( .A1(n6838), .A2(n4505), .ZN(n4504) );
  NAND2_X1 U5457 ( .A1(n6224), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n4505) );
  NAND2_X1 U5458 ( .A1(n4323), .A2(n7062), .ZN(n7061) );
  NAND2_X1 U5459 ( .A1(n6676), .A2(n4523), .ZN(n4522) );
  INV_X1 U5460 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n4523) );
  OR2_X1 U5461 ( .A1(n6227), .A2(n7232), .ZN(n4520) );
  XNOR2_X1 U5462 ( .A(n6233), .B(n6245), .ZN(n8652) );
  NAND2_X1 U5463 ( .A1(n8652), .A2(n8651), .ZN(n8650) );
  NAND2_X1 U5464 ( .A1(n8063), .A2(n8062), .ZN(n8666) );
  NAND2_X1 U5465 ( .A1(n8065), .A2(n8064), .ZN(n8947) );
  OR2_X1 U5466 ( .A1(n8695), .A2(n8950), .ZN(n8674) );
  AND2_X1 U5467 ( .A1(n8234), .A2(n8231), .ZN(n8710) );
  AND4_X1 U5468 ( .A1(n6097), .A2(n6096), .A3(n6095), .A4(n6094), .ZN(n8746)
         );
  AND4_X1 U5469 ( .A1(n6116), .A2(n6115), .A3(n6114), .A4(n6113), .ZN(n8745)
         );
  NAND2_X1 U5470 ( .A1(n4418), .A2(n8214), .ZN(n8753) );
  NOR2_X1 U5471 ( .A1(n8076), .A2(n4819), .ZN(n4815) );
  NOR2_X1 U5472 ( .A1(n8792), .A2(n8983), .ZN(n8773) );
  NOR2_X1 U5473 ( .A1(n8797), .A2(n4612), .ZN(n4611) );
  INV_X1 U5474 ( .A(n8212), .ZN(n4612) );
  NAND2_X1 U5475 ( .A1(n8843), .A2(n4472), .ZN(n8792) );
  NOR2_X1 U5476 ( .A1(n8988), .A2(n4473), .ZN(n4472) );
  INV_X1 U5477 ( .A(n4474), .ZN(n4473) );
  NAND2_X1 U5478 ( .A1(n8843), .A2(n8450), .ZN(n8834) );
  NAND2_X1 U5479 ( .A1(n8268), .A2(n5751), .ZN(n4685) );
  OR2_X1 U5480 ( .A1(n8887), .A2(n9012), .ZN(n8866) );
  NOR2_X1 U5481 ( .A1(n8866), .A2(n9005), .ZN(n8843) );
  NAND2_X1 U5482 ( .A1(n4603), .A2(n4314), .ZN(n8859) );
  OR2_X1 U5483 ( .A1(n8899), .A2(n4605), .ZN(n4603) );
  NAND2_X1 U5484 ( .A1(n8004), .A2(n4467), .ZN(n8887) );
  AND2_X1 U5485 ( .A1(n4468), .A2(n8892), .ZN(n4467) );
  NAND2_X1 U5486 ( .A1(n8069), .A2(n8430), .ZN(n8875) );
  AND2_X1 U5487 ( .A1(n4607), .A2(n4422), .ZN(n8876) );
  OR2_X1 U5488 ( .A1(n8899), .A2(n4357), .ZN(n4607) );
  AND2_X1 U5489 ( .A1(n8004), .A2(n4468), .ZN(n8909) );
  NAND2_X1 U5490 ( .A1(n8900), .A2(n8184), .ZN(n8926) );
  NOR2_X1 U5491 ( .A1(n7992), .A2(n8182), .ZN(n8427) );
  NAND2_X1 U5492 ( .A1(n8004), .A2(n8003), .ZN(n8928) );
  AND2_X1 U5493 ( .A1(n4592), .A2(n8177), .ZN(n4591) );
  INV_X1 U5494 ( .A(n4597), .ZN(n4590) );
  AOI21_X1 U5495 ( .B1(n4597), .B2(n4596), .A(n4595), .ZN(n4589) );
  NAND2_X1 U5496 ( .A1(n7733), .A2(n4303), .ZN(n7858) );
  NAND2_X1 U5497 ( .A1(n7733), .A2(n7694), .ZN(n7716) );
  AND2_X1 U5498 ( .A1(n7574), .A2(n9972), .ZN(n7733) );
  NAND2_X1 U5499 ( .A1(n7681), .A2(n8154), .ZN(n7724) );
  OR2_X1 U5500 ( .A1(n9928), .A2(n7140), .ZN(n7138) );
  NOR2_X1 U5501 ( .A1(n7615), .A2(n8373), .ZN(n9927) );
  AND2_X1 U5502 ( .A1(n5759), .A2(n9952), .ZN(n7067) );
  NAND2_X1 U5503 ( .A1(n8425), .A2(n9952), .ZN(n7590) );
  AND2_X1 U5504 ( .A1(n6236), .A2(n6206), .ZN(n8862) );
  AND2_X1 U5505 ( .A1(n9953), .A2(n7496), .ZN(n9913) );
  AND2_X1 U5506 ( .A1(n7852), .A2(n7783), .ZN(n4832) );
  NOR2_X1 U5507 ( .A1(n7682), .A2(n4813), .ZN(n4812) );
  INV_X1 U5508 ( .A(n7687), .ZN(n4813) );
  AND2_X1 U5509 ( .A1(n6172), .A2(n6171), .ZN(n6186) );
  XNOR2_X1 U5510 ( .A(n6167), .B(n6166), .ZN(n6237) );
  NAND2_X1 U5511 ( .A1(n6165), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6167) );
  XNOR2_X1 U5512 ( .A(n6187), .B(P2_IR_REG_23__SCAN_IN), .ZN(n9945) );
  NAND2_X1 U5513 ( .A1(n6155), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6162) );
  INV_X1 U5514 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n6161) );
  INV_X1 U5515 ( .A(n5929), .ZN(n5976) );
  INV_X1 U5516 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n4717) );
  INV_X1 U5517 ( .A(n5798), .ZN(n4805) );
  AOI21_X1 U5518 ( .B1(n5625), .B2(n5624), .A(n5703), .ZN(n5629) );
  NAND2_X1 U5519 ( .A1(n4450), .A2(n7481), .ZN(n7262) );
  INV_X1 U5520 ( .A(n5250), .ZN(n4448) );
  AOI21_X1 U5521 ( .B1(n5250), .B2(n4447), .A(n4318), .ZN(n4446) );
  AND2_X1 U5522 ( .A1(n5623), .A2(n5622), .ZN(n5703) );
  OR2_X1 U5523 ( .A1(n5474), .A2(n9104), .ZN(n5497) );
  INV_X1 U5524 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n9104) );
  NAND2_X1 U5525 ( .A1(n4621), .A2(n4619), .ZN(n7640) );
  NOR2_X1 U5526 ( .A1(n7643), .A2(n4620), .ZN(n4619) );
  INV_X1 U5527 ( .A(n7263), .ZN(n4620) );
  INV_X1 U5528 ( .A(n6432), .ZN(n4565) );
  AND2_X1 U5529 ( .A1(n5591), .A2(n5590), .ZN(n6472) );
  NAND2_X1 U5530 ( .A1(n8356), .A2(n6591), .ZN(n6736) );
  OR2_X1 U5531 ( .A1(n5233), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n5255) );
  AND2_X1 U5532 ( .A1(n9640), .A2(n9639), .ZN(n9642) );
  AND2_X1 U5533 ( .A1(n4464), .A2(n4463), .ZN(n9684) );
  NAND2_X1 U5534 ( .A1(n8279), .A2(n9674), .ZN(n4463) );
  AND2_X1 U5535 ( .A1(n9200), .A2(n9203), .ZN(n9227) );
  NAND2_X1 U5536 ( .A1(n9228), .A2(n9734), .ZN(n9231) );
  OR2_X1 U5537 ( .A1(n9248), .A2(n9228), .ZN(n9182) );
  AND2_X1 U5538 ( .A1(n9183), .A2(n9182), .ZN(n4796) );
  AND2_X1 U5539 ( .A1(n5682), .A2(n5681), .ZN(n9245) );
  AND2_X1 U5540 ( .A1(n5616), .A2(n5615), .ZN(n9267) );
  NOR2_X1 U5541 ( .A1(n9194), .A2(n9196), .ZN(n9281) );
  INV_X1 U5542 ( .A(n9193), .ZN(n4663) );
  AOI21_X1 U5543 ( .B1(n4293), .B2(n4772), .A(n4771), .ZN(n4770) );
  NOR2_X1 U5544 ( .A1(n9301), .A2(n9316), .ZN(n4771) );
  NAND2_X1 U5545 ( .A1(n5024), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5535) );
  OR2_X1 U5546 ( .A1(n9442), .A2(n9177), .ZN(n9342) );
  NOR2_X1 U5547 ( .A1(n9371), .A2(n4578), .ZN(n9337) );
  INV_X1 U5548 ( .A(n4580), .ZN(n4578) );
  AND2_X1 U5549 ( .A1(n5504), .A2(n5503), .ZN(n9363) );
  NOR2_X1 U5550 ( .A1(n9371), .A2(n9442), .ZN(n9353) );
  OAI21_X1 U5551 ( .B1(n8040), .B2(n4317), .A(n4787), .ZN(n9352) );
  NOR2_X1 U5552 ( .A1(n4789), .A2(n4788), .ZN(n4787) );
  NOR2_X1 U5553 ( .A1(n9377), .A2(n9362), .ZN(n4788) );
  AND2_X1 U5554 ( .A1(n9342), .A2(n6496), .ZN(n9359) );
  NAND2_X1 U5555 ( .A1(n5021), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5456) );
  INV_X1 U5556 ( .A(n5444), .ZN(n5021) );
  NOR2_X1 U5557 ( .A1(n4678), .A2(n4677), .ZN(n4676) );
  OAI21_X1 U5558 ( .B1(n4296), .B2(n4678), .A(n6457), .ZN(n4675) );
  INV_X1 U5559 ( .A(n4682), .ZN(n4677) );
  NAND2_X1 U5560 ( .A1(n5020), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5416) );
  INV_X1 U5561 ( .A(n5414), .ZN(n5020) );
  AND3_X1 U5562 ( .A1(n5063), .A2(n5062), .A3(n5061), .ZN(n8037) );
  NAND2_X1 U5563 ( .A1(n7829), .A2(n4572), .ZN(n7916) );
  AOI21_X1 U5564 ( .B1(n4799), .B2(n4802), .A(n4340), .ZN(n4798) );
  NAND2_X1 U5565 ( .A1(n5019), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n5393) );
  INV_X1 U5566 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n5392) );
  NAND2_X1 U5567 ( .A1(n7829), .A2(n9588), .ZN(n7844) );
  AOI21_X1 U5568 ( .B1(n4783), .B2(n4332), .A(n4781), .ZN(n9555) );
  OAI21_X1 U5569 ( .B1(n7157), .B2(n6319), .A(n4782), .ZN(n4781) );
  INV_X1 U5570 ( .A(n7546), .ZN(n4782) );
  AND4_X1 U5571 ( .A1(n5246), .A2(n5245), .A3(n5244), .A4(n5243), .ZN(n7207)
         );
  NOR2_X1 U5572 ( .A1(n4576), .A2(n7334), .ZN(n7331) );
  INV_X1 U5573 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5239) );
  OR2_X1 U5574 ( .A1(n5263), .A2(n5239), .ZN(n5281) );
  AND4_X1 U5575 ( .A1(n5268), .A2(n5267), .A3(n5266), .A4(n5265), .ZN(n8315)
         );
  NAND2_X1 U5576 ( .A1(n7148), .A2(n7147), .ZN(n7193) );
  AND2_X1 U5577 ( .A1(n7099), .A2(n7148), .ZN(n4653) );
  NAND2_X1 U5578 ( .A1(n9750), .A2(n9841), .ZN(n9731) );
  NAND2_X1 U5579 ( .A1(n9750), .A2(n4575), .ZN(n7185) );
  OAI21_X1 U5580 ( .B1(n9779), .B2(n9758), .A(n6308), .ZN(n4566) );
  INV_X1 U5581 ( .A(n9159), .ZN(n9767) );
  INV_X1 U5582 ( .A(n7023), .ZN(n7012) );
  NAND2_X1 U5583 ( .A1(n5409), .A2(n4451), .ZN(n5049) );
  NOR2_X1 U5584 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(n4350), .ZN(n4451) );
  NAND2_X1 U5585 ( .A1(n7022), .A2(n7023), .ZN(n7021) );
  NAND2_X1 U5586 ( .A1(n5583), .A2(n5582), .ZN(n9412) );
  NOR2_X1 U5587 ( .A1(n7827), .A2(n7826), .ZN(n7838) );
  OR2_X1 U5588 ( .A1(n7029), .A2(n5660), .ZN(n9865) );
  INV_X1 U5589 ( .A(n9865), .ZN(n9857) );
  NAND2_X1 U5590 ( .A1(n5636), .A2(n5637), .ZN(n6701) );
  XNOR2_X1 U5591 ( .A(n6407), .B(SI_30_), .ZN(n8060) );
  NOR2_X1 U5592 ( .A1(n4306), .A2(P1_IR_REG_23__SCAN_IN), .ZN(n4793) );
  INV_X1 U5593 ( .A(n5671), .ZN(n7024) );
  XNOR2_X1 U5594 ( .A(n5691), .B(n5690), .ZN(n8029) );
  INV_X1 U5595 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5001) );
  AND2_X1 U5596 ( .A1(n4326), .A2(n4684), .ZN(n4683) );
  NAND2_X1 U5597 ( .A1(n4750), .A2(n4754), .ZN(n5531) );
  AOI21_X1 U5598 ( .B1(n4758), .B2(n4756), .A(n4755), .ZN(n4754) );
  INV_X1 U5599 ( .A(n6558), .ZN(n6577) );
  AOI21_X1 U5600 ( .B1(n4950), .B2(n4732), .A(n4369), .ZN(n4731) );
  INV_X1 U5601 ( .A(n4948), .ZN(n4732) );
  NAND2_X1 U5602 ( .A1(n4949), .A2(n4948), .ZN(n5436) );
  NAND2_X1 U5603 ( .A1(n5409), .A2(n5007), .ZN(n5054) );
  NAND2_X1 U5604 ( .A1(n5385), .A2(n4935), .ZN(n5407) );
  NAND2_X1 U5605 ( .A1(n5384), .A2(n5385), .ZN(n6749) );
  NAND2_X1 U5606 ( .A1(n4295), .A2(n4928), .ZN(n5383) );
  NAND2_X1 U5607 ( .A1(n4561), .A2(n4980), .ZN(n5344) );
  AND4_X1 U5608 ( .A1(n4560), .A2(n4981), .A3(n4975), .A4(n5068), .ZN(n4561)
         );
  NAND2_X1 U5609 ( .A1(n4734), .A2(n4736), .ZN(n5297) );
  OR2_X1 U5610 ( .A1(n5254), .A2(n4739), .ZN(n4734) );
  XNOR2_X1 U5611 ( .A(n4414), .B(n4848), .ZN(n6657) );
  OAI21_X1 U5612 ( .B1(n5254), .B2(n4904), .A(n4903), .ZN(n4414) );
  NOR2_X1 U5613 ( .A1(n5068), .A2(n9493), .ZN(n5069) );
  AND4_X1 U5614 ( .A1(n5823), .A2(n5822), .A3(n5821), .A4(n5820), .ZN(n7727)
         );
  NAND2_X1 U5615 ( .A1(n8405), .A2(n5832), .ZN(n6571) );
  NAND2_X1 U5616 ( .A1(n4413), .A2(n5900), .ZN(n7883) );
  NAND2_X1 U5617 ( .A1(n7760), .A2(n5882), .ZN(n4413) );
  NAND2_X1 U5618 ( .A1(n4687), .A2(n4686), .ZN(n7900) );
  AOI21_X1 U5619 ( .B1(n4688), .B2(n4689), .A(n4343), .ZN(n4686) );
  AND4_X1 U5620 ( .A1(n6017), .A2(n6016), .A3(n6015), .A4(n6014), .ZN(n8832)
         );
  NAND2_X1 U5621 ( .A1(n8521), .A2(n5990), .ZN(n4711) );
  NAND2_X1 U5622 ( .A1(n4692), .A2(n8481), .ZN(n7343) );
  NAND2_X1 U5623 ( .A1(n8487), .A2(n6035), .ZN(n8552) );
  NAND2_X1 U5624 ( .A1(n7772), .A2(n7773), .ZN(n7925) );
  AND4_X1 U5625 ( .A1(n6072), .A2(n6071), .A3(n6070), .A4(n6069), .ZN(n8757)
         );
  INV_X1 U5626 ( .A(n7988), .ZN(n10013) );
  OAI21_X1 U5627 ( .B1(n7534), .B2(n4689), .A(n4688), .ZN(n7761) );
  INV_X1 U5628 ( .A(n8592), .ZN(n8514) );
  INV_X1 U5629 ( .A(n8593), .ZN(n8488) );
  AND4_X1 U5630 ( .A1(n6029), .A2(n6028), .A3(n6027), .A4(n6026), .ZN(n8578)
         );
  OAI21_X1 U5631 ( .B1(n8521), .B2(n4400), .A(n4397), .ZN(n8486) );
  AND2_X1 U5632 ( .A1(n4691), .A2(n7044), .ZN(n4690) );
  NAND2_X1 U5633 ( .A1(n6191), .A2(n8718), .ZN(n8589) );
  AND4_X1 U5634 ( .A1(n5954), .A2(n5953), .A3(n5952), .A4(n5951), .ZN(n8904)
         );
  NAND2_X1 U5635 ( .A1(n8509), .A2(n8861), .ZN(n8598) );
  INV_X1 U5636 ( .A(n8589), .ZN(n8604) );
  NAND2_X1 U5637 ( .A1(n5974), .A2(n5966), .ZN(n8594) );
  NAND2_X1 U5638 ( .A1(n4718), .A2(n5974), .ZN(n8595) );
  INV_X1 U5639 ( .A(n4719), .ZN(n4718) );
  INV_X1 U5640 ( .A(n8270), .ZN(n4425) );
  AND3_X1 U5641 ( .A1(n6672), .A2(n6671), .A3(n6670), .ZN(n8449) );
  AND3_X1 U5642 ( .A1(n6205), .A2(n6204), .A3(n6203), .ZN(n8081) );
  OR2_X1 U5643 ( .A1(n6241), .A2(n9945), .ZN(n6760) );
  INV_X1 U5644 ( .A(n8578), .ZN(n8851) );
  INV_X1 U5645 ( .A(n7726), .ZN(n8615) );
  INV_X1 U5646 ( .A(n6217), .ZN(n9506) );
  INV_X1 U5647 ( .A(n4488), .ZN(n9505) );
  AOI21_X1 U5648 ( .B1(n9521), .B2(P2_REG2_REG_2__SCAN_IN), .A(n9518), .ZN(
        n6999) );
  AOI21_X1 U5649 ( .B1(n6254), .B2(P2_REG2_REG_3__SCAN_IN), .A(n6997), .ZN(
        n6951) );
  INV_X1 U5650 ( .A(n4492), .ZN(n6973) );
  NOR2_X1 U5651 ( .A1(n6939), .A2(n6938), .ZN(n6937) );
  AND2_X1 U5652 ( .A1(n4492), .A2(n4491), .ZN(n6939) );
  NAND2_X1 U5653 ( .A1(n6252), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n4491) );
  AOI21_X1 U5654 ( .B1(n6250), .B2(P2_REG2_REG_6__SCAN_IN), .A(n6937), .ZN(
        n6963) );
  OR2_X1 U5655 ( .A1(n6837), .A2(n6836), .ZN(n6838) );
  AND2_X1 U5656 ( .A1(n6279), .A2(n6278), .ZN(n9888) );
  INV_X1 U5657 ( .A(n4502), .ZN(n6985) );
  INV_X1 U5658 ( .A(n4504), .ZN(n6987) );
  OR2_X1 U5659 ( .A1(n6899), .A2(n6898), .ZN(n6900) );
  NAND2_X1 U5660 ( .A1(n4510), .A2(n4514), .ZN(n7746) );
  OR2_X1 U5661 ( .A1(n6227), .A2(n4515), .ZN(n4510) );
  AND2_X1 U5662 ( .A1(n5961), .A2(n5948), .ZN(n7751) );
  NAND2_X1 U5663 ( .A1(n7947), .A2(n4320), .ZN(n4507) );
  INV_X1 U5664 ( .A(n9895), .ZN(n9889) );
  INV_X1 U5665 ( .A(n8666), .ZN(n8945) );
  OR2_X1 U5666 ( .A1(n8950), .A2(n8605), .ZN(n8440) );
  AND2_X1 U5667 ( .A1(n6146), .A2(n6135), .ZN(n8698) );
  OAI21_X1 U5668 ( .B1(n8706), .B2(n4811), .A(n4809), .ZN(n8687) );
  NAND2_X1 U5669 ( .A1(n8704), .A2(n8439), .ZN(n8688) );
  NAND2_X1 U5670 ( .A1(n8740), .A2(n8224), .ZN(n8729) );
  INV_X1 U5671 ( .A(n8451), .ZN(n8737) );
  NAND2_X1 U5672 ( .A1(n8856), .A2(n4823), .ZN(n4818) );
  AND2_X1 U5673 ( .A1(n8788), .A2(n8787), .ZN(n8996) );
  AND2_X1 U5674 ( .A1(n5915), .A2(n5914), .ZN(n10020) );
  NAND2_X1 U5675 ( .A1(n7990), .A2(n4835), .ZN(n9909) );
  AND2_X1 U5676 ( .A1(n7990), .A2(n7989), .ZN(n9910) );
  NAND2_X1 U5677 ( .A1(n7784), .A2(n7783), .ZN(n7785) );
  NAND2_X1 U5678 ( .A1(n7778), .A2(n8173), .ZN(n7853) );
  NAND2_X1 U5679 ( .A1(n7688), .A2(n7687), .ZN(n7690) );
  NAND2_X1 U5680 ( .A1(n7569), .A2(n7568), .ZN(n7686) );
  OR2_X1 U5681 ( .A1(n9937), .A2(n7529), .ZN(n8918) );
  OR2_X1 U5682 ( .A1(n6082), .A2(n6629), .ZN(n5785) );
  AND2_X1 U5683 ( .A1(n7521), .A2(n7520), .ZN(n9933) );
  NAND2_X1 U5684 ( .A1(n7518), .A2(n8718), .ZN(n8916) );
  OR2_X1 U5685 ( .A1(n9939), .A2(n6905), .ZN(n8718) );
  INV_X1 U5686 ( .A(n9906), .ZN(n9931) );
  AND2_X1 U5687 ( .A1(n9933), .A2(n9913), .ZN(n8896) );
  AND2_X2 U5688 ( .A1(n6933), .A2(n7514), .ZN(n10045) );
  NAND2_X1 U5689 ( .A1(n4485), .A2(n4482), .ZN(n9023) );
  INV_X1 U5690 ( .A(n8946), .ZN(n4485) );
  INV_X1 U5691 ( .A(n4483), .ZN(n4482) );
  OAI21_X1 U5692 ( .B1(n8949), .B2(n10001), .A(n4484), .ZN(n4483) );
  AND2_X2 U5693 ( .A1(n6933), .A2(n6910), .ZN(n10028) );
  INV_X1 U5694 ( .A(n9944), .ZN(n9948) );
  NAND2_X1 U5695 ( .A1(n5732), .A2(n5733), .ZN(n9050) );
  OR2_X1 U5696 ( .A1(n5731), .A2(n5728), .ZN(n5729) );
  AND2_X1 U5697 ( .A1(n6160), .A2(n6169), .ZN(n7943) );
  INV_X1 U5698 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7867) );
  INV_X1 U5699 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7771) );
  INV_X1 U5700 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n8058) );
  INV_X1 U5701 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7511) );
  XNOR2_X1 U5702 ( .A(n5743), .B(n5742), .ZN(n8133) );
  INV_X1 U5703 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7497) );
  INV_X1 U5704 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6809) );
  INV_X1 U5705 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6687) );
  INV_X1 U5706 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n7440) );
  INV_X1 U5707 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6678) );
  INV_X1 U5708 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6660) );
  INV_X1 U5709 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6653) );
  INV_X1 U5710 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6646) );
  XNOR2_X1 U5711 ( .A(n5771), .B(n5770), .ZN(n6638) );
  NAND2_X1 U5712 ( .A1(n4499), .A2(n4496), .ZN(n6635) );
  NAND2_X1 U5713 ( .A1(n4498), .A2(n4497), .ZN(n4496) );
  INV_X1 U5714 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n4497) );
  OR2_X1 U5715 ( .A1(n6568), .A2(n6577), .ZN(n6613) );
  NAND2_X1 U5716 ( .A1(n7650), .A2(n4316), .ZN(n4631) );
  NOR2_X1 U5717 ( .A1(n4638), .A2(n4641), .ZN(n4637) );
  AOI22_X1 U5718 ( .A1(n4638), .A2(n4644), .B1(n4641), .B2(n9080), .ZN(n4636)
         );
  AND2_X1 U5719 ( .A1(n4642), .A2(n4639), .ZN(n4638) );
  AOI22_X1 U5720 ( .A1(n4287), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6579), .B2(
        n6745), .ZN(n5259) );
  OR2_X1 U5721 ( .A1(n5863), .A2(n5108), .ZN(n5260) );
  XNOR2_X1 U5722 ( .A(n4452), .B(n5247), .ZN(n6730) );
  OAI21_X1 U5723 ( .B1(n5093), .B2(n6693), .A(n5117), .ZN(n4452) );
  NAND2_X1 U5724 ( .A1(n9072), .A2(n9073), .ZN(n9071) );
  NAND2_X1 U5725 ( .A1(n9098), .A2(n5491), .ZN(n9072) );
  NOR2_X1 U5726 ( .A1(n8019), .A2(n4336), .ZN(n8023) );
  NAND2_X1 U5727 ( .A1(n5669), .A2(n6692), .ZN(n9140) );
  INV_X1 U5728 ( .A(n9114), .ZN(n9139) );
  NAND2_X1 U5729 ( .A1(n7650), .A2(n5341), .ZN(n7673) );
  NAND2_X1 U5730 ( .A1(n4621), .A2(n7263), .ZN(n7642) );
  AND4_X1 U5731 ( .A1(n5332), .A2(n5331), .A3(n5330), .A4(n5329), .ZN(n7674)
         );
  NOR2_X1 U5732 ( .A1(n4839), .A2(n5137), .ZN(n5138) );
  NAND2_X1 U5733 ( .A1(n4647), .A2(n4641), .ZN(n9120) );
  NAND2_X1 U5734 ( .A1(n4645), .A2(n4643), .ZN(n4640) );
  INV_X1 U5735 ( .A(n9140), .ZN(n9127) );
  INV_X1 U5736 ( .A(n9735), .ZN(n7315) );
  OR2_X1 U5737 ( .A1(n5683), .A2(n7024), .ZN(n9123) );
  INV_X1 U5738 ( .A(n7912), .ZN(n9580) );
  AND2_X1 U5739 ( .A1(n5662), .A2(n9792), .ZN(n9148) );
  OR2_X1 U5740 ( .A1(n5683), .A2(n5671), .ZN(n9114) );
  AND2_X1 U5741 ( .A1(n9863), .A2(n5656), .ZN(n9136) );
  INV_X1 U5742 ( .A(n9123), .ZN(n9145) );
  OAI21_X1 U5743 ( .B1(n6553), .B2(n4563), .A(n4562), .ZN(n6561) );
  NAND2_X1 U5744 ( .A1(n6491), .A2(n4564), .ZN(n4563) );
  NOR2_X1 U5745 ( .A1(n6552), .A2(n6551), .ZN(n4562) );
  NOR2_X1 U5746 ( .A1(n7019), .A2(n5655), .ZN(n4564) );
  INV_X1 U5747 ( .A(n9267), .ZN(n9228) );
  INV_X1 U5748 ( .A(n6472), .ZN(n9284) );
  INV_X1 U5749 ( .A(n8037), .ZN(n9149) );
  INV_X1 U5750 ( .A(n9783), .ZN(n9160) );
  NAND2_X1 U5751 ( .A1(n5586), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5089) );
  NAND2_X1 U5752 ( .A1(n6849), .A2(n6584), .ZN(n6826) );
  NAND2_X1 U5753 ( .A1(n6827), .A2(n6826), .ZN(n6825) );
  NAND2_X1 U5754 ( .A1(n9621), .A2(n6590), .ZN(n8358) );
  NAND2_X1 U5755 ( .A1(n8331), .A2(n6777), .ZN(n6779) );
  INV_X1 U5756 ( .A(n4464), .ZN(n9670) );
  OR2_X1 U5757 ( .A1(n8305), .A2(n7024), .ZN(n9717) );
  INV_X1 U5758 ( .A(n9724), .ZN(n9704) );
  NAND2_X1 U5759 ( .A1(n9258), .A2(n4582), .ZN(n9391) );
  NOR2_X1 U5760 ( .A1(n9169), .A2(n4583), .ZN(n4582) );
  OR2_X1 U5761 ( .A1(n4584), .A2(n9248), .ZN(n4583) );
  NAND2_X1 U5762 ( .A1(n6389), .A2(n6388), .ZN(n9398) );
  INV_X1 U5763 ( .A(n9412), .ZN(n9262) );
  AND2_X1 U5764 ( .A1(n5559), .A2(n5558), .ZN(n9280) );
  OAI21_X1 U5765 ( .B1(n9327), .B2(n4668), .A(n4666), .ZN(n9290) );
  NAND2_X1 U5766 ( .A1(n4665), .A2(n4669), .ZN(n9292) );
  NAND2_X1 U5767 ( .A1(n4769), .A2(n4293), .ZN(n9289) );
  OR2_X1 U5768 ( .A1(n9319), .A2(n4776), .ZN(n4769) );
  AND2_X1 U5769 ( .A1(n4673), .A2(n4674), .ZN(n9313) );
  NAND2_X1 U5770 ( .A1(n9327), .A2(n9191), .ZN(n4673) );
  NAND2_X1 U5771 ( .A1(n4779), .A2(n4842), .ZN(n9305) );
  NAND2_X1 U5772 ( .A1(n9319), .A2(n9178), .ZN(n4779) );
  INV_X1 U5773 ( .A(n9432), .ZN(n9325) );
  NAND2_X1 U5774 ( .A1(n9186), .A2(n9185), .ZN(n9379) );
  NOR2_X1 U5775 ( .A1(n9173), .A2(n4792), .ZN(n9370) );
  AND2_X1 U5776 ( .A1(n4680), .A2(n4679), .ZN(n7839) );
  AND2_X1 U5777 ( .A1(n4800), .A2(n4801), .ZN(n7915) );
  OR2_X1 U5778 ( .A1(n7841), .A2(n4802), .ZN(n4800) );
  NAND2_X1 U5779 ( .A1(n5347), .A2(n5346), .ZN(n7823) );
  NAND2_X1 U5780 ( .A1(n7198), .A2(n7157), .ZN(n7548) );
  OR2_X1 U5781 ( .A1(n6648), .A2(n5108), .ZN(n5215) );
  AND2_X1 U5782 ( .A1(n7125), .A2(n7124), .ZN(n9769) );
  OR2_X1 U5783 ( .A1(n5108), .A2(n6630), .ZN(n5133) );
  OR2_X1 U5784 ( .A1(n6414), .A2(n4870), .ZN(n5073) );
  OAI21_X1 U5785 ( .B1(n7012), .B2(n7013), .A(n7108), .ZN(n9810) );
  AND2_X2 U5786 ( .A1(n6718), .A2(n6717), .ZN(n9887) );
  AND2_X2 U5787 ( .A1(n7015), .A2(n6718), .ZN(n9872) );
  AND2_X1 U5788 ( .A1(n6568), .A2(n5654), .ZN(n6688) );
  OAI21_X1 U5789 ( .B1(n6407), .B2(n6406), .A(n6410), .ZN(n4733) );
  XNOR2_X1 U5790 ( .A(n6384), .B(n6383), .ZN(n8459) );
  NAND2_X1 U5791 ( .A1(n4743), .A2(n5692), .ZN(n6384) );
  INV_X1 U5792 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7942) );
  INV_X1 U5793 ( .A(n5634), .ZN(n7896) );
  NAND2_X1 U5794 ( .A1(n4753), .A2(n4758), .ZN(n5529) );
  NAND2_X1 U5795 ( .A1(n5493), .A2(n4760), .ZN(n4753) );
  INV_X1 U5796 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7757) );
  INV_X1 U5797 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7500) );
  INV_X1 U5798 ( .A(n6705), .ZN(n7499) );
  INV_X1 U5799 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n8386) );
  INV_X1 U5800 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7230) );
  INV_X1 U5801 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6675) );
  NAND2_X1 U5802 ( .A1(n5229), .A2(n5228), .ZN(n4552) );
  NAND2_X1 U5803 ( .A1(n4409), .A2(n4884), .ZN(n5192) );
  NOR2_X1 U5804 ( .A1(n4278), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9496) );
  NOR2_X1 U5805 ( .A1(n7814), .A2(n10084), .ZN(n10073) );
  AOI21_X1 U5806 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10071), .ZN(n10070) );
  NOR2_X1 U5807 ( .A1(n10070), .A2(n10069), .ZN(n10068) );
  AOI21_X1 U5808 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10068), .ZN(n10067) );
  OAI21_X1 U5809 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10065), .ZN(n10063) );
  AND2_X1 U5810 ( .A1(n6213), .A2(n6212), .ZN(n4706) );
  NAND2_X1 U5811 ( .A1(n4695), .A2(n4699), .ZN(n4694) );
  NAND2_X1 U5812 ( .A1(n4403), .A2(n4401), .ZN(P2_U3227) );
  NOR2_X1 U5813 ( .A1(n8520), .A2(n4402), .ZN(n4401) );
  NAND2_X1 U5814 ( .A1(n4424), .A2(n8269), .ZN(P2_U3244) );
  NAND2_X1 U5815 ( .A1(n4426), .A2(n4425), .ZN(n4424) );
  AOI21_X1 U5816 ( .B1(n6292), .B2(n5751), .A(n6291), .ZN(n6293) );
  INV_X1 U5817 ( .A(n4438), .ZN(n4437) );
  INV_X1 U5818 ( .A(n4459), .ZN(n4458) );
  NAND2_X1 U5819 ( .A1(n4461), .A2(n9298), .ZN(n4460) );
  NAND2_X1 U5820 ( .A1(n4457), .A2(n9757), .ZN(n4456) );
  NOR2_X1 U5821 ( .A1(n9404), .A2(n9568), .ZN(n9234) );
  AND2_X1 U5822 ( .A1(n8204), .A2(n8777), .ZN(n4291) );
  AND2_X1 U5823 ( .A1(n4572), .A2(n4571), .ZN(n4292) );
  INV_X2 U5824 ( .A(n5247), .ZN(n7124) );
  AND2_X1 U5825 ( .A1(n4774), .A2(n4780), .ZN(n4293) );
  XOR2_X1 U5826 ( .A(n5450), .B(n7124), .Z(n4294) );
  AND2_X1 U5827 ( .A1(n8173), .A2(n8164), .ZN(n8100) );
  INV_X1 U5828 ( .A(n8100), .ZN(n4596) );
  AND2_X1 U5829 ( .A1(n7842), .A2(n4679), .ZN(n4296) );
  OR2_X1 U5830 ( .A1(n4532), .A2(n4531), .ZN(n4297) );
  NAND2_X1 U5831 ( .A1(n4784), .A2(n4976), .ZN(n5146) );
  INV_X1 U5832 ( .A(n8858), .ZN(n4826) );
  OR2_X1 U5833 ( .A1(n7727), .A2(n9972), .ZN(n4298) );
  OR2_X1 U5834 ( .A1(n5727), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n4299) );
  INV_X1 U5835 ( .A(n8806), .ZN(n4539) );
  NAND2_X1 U5836 ( .A1(n4805), .A2(n4362), .ZN(n4300) );
  OR2_X1 U5837 ( .A1(n8666), .A2(n8449), .ZN(n4302) );
  AND2_X1 U5838 ( .A1(n7694), .A2(n9994), .ZN(n4303) );
  AND2_X1 U5839 ( .A1(n4821), .A2(n8772), .ZN(n4304) );
  INV_X1 U5840 ( .A(n9080), .ZN(n4646) );
  AND2_X1 U5841 ( .A1(n4344), .A2(n7344), .ZN(n4305) );
  NAND3_X1 U5842 ( .A1(n5031), .A2(n5030), .A3(n5029), .ZN(n4306) );
  NOR2_X1 U5843 ( .A1(n8002), .A2(n8611), .ZN(n4307) );
  NAND2_X1 U5844 ( .A1(n8205), .A2(n4537), .ZN(n4308) );
  NAND2_X1 U5845 ( .A1(n4278), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n4309) );
  AND2_X1 U5846 ( .A1(n5056), .A2(n5055), .ZN(n9084) );
  INV_X1 U5847 ( .A(n9084), .ZN(n9458) );
  INV_X1 U5848 ( .A(n8970), .ZN(n4480) );
  NAND2_X1 U5849 ( .A1(n8843), .A2(n4474), .ZN(n4475) );
  OR2_X1 U5850 ( .A1(n6681), .A2(n4521), .ZN(n4310) );
  NAND2_X1 U5851 ( .A1(n8628), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n4311) );
  INV_X1 U5852 ( .A(n7098), .ZN(n4655) );
  OR2_X1 U5853 ( .A1(n4311), .A2(n8638), .ZN(n4312) );
  INV_X1 U5854 ( .A(n8373), .ZN(n7070) );
  OAI211_X1 U5855 ( .C1(n6286), .C2(n6638), .A(n5773), .B(n5772), .ZN(n8373)
         );
  NAND2_X1 U5856 ( .A1(n4825), .A2(n4822), .ZN(n8785) );
  NAND2_X1 U5857 ( .A1(n4274), .A2(n4278), .ZN(n5108) );
  AND2_X1 U5858 ( .A1(n5190), .A2(n5189), .ZN(n4313) );
  INV_X1 U5859 ( .A(n8088), .ZN(n5751) );
  OAI21_X1 U5860 ( .B1(n5049), .B2(P1_IR_REG_19__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n4999) );
  OR2_X1 U5861 ( .A1(n8193), .A2(n4421), .ZN(n4314) );
  NAND2_X1 U5862 ( .A1(n4411), .A2(n8499), .ZN(n8502) );
  NAND2_X1 U5863 ( .A1(n6121), .A2(n6120), .ZN(n8961) );
  AND2_X1 U5864 ( .A1(n4934), .A2(n4928), .ZN(n4315) );
  NOR2_X1 U5865 ( .A1(n5362), .A2(n4635), .ZN(n4316) );
  AND2_X1 U5866 ( .A1(n5236), .A2(n5235), .ZN(n9864) );
  AND4_X1 U5867 ( .A1(n5781), .A2(n5780), .A3(n5779), .A4(n5778), .ZN(n7074)
         );
  OR2_X1 U5868 ( .A1(n9175), .A2(n8041), .ZN(n4317) );
  NOR2_X1 U5869 ( .A1(n5144), .A2(n4785), .ZN(n5174) );
  NOR2_X1 U5870 ( .A1(n5293), .A2(n7305), .ZN(n4318) );
  NOR2_X1 U5871 ( .A1(n5573), .A2(n8320), .ZN(n4319) );
  NAND2_X1 U5872 ( .A1(n4990), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5000) );
  AND2_X1 U5873 ( .A1(n6231), .A2(n4508), .ZN(n4320) );
  AND2_X1 U5874 ( .A1(n4488), .A2(n4487), .ZN(n4321) );
  NAND2_X1 U5875 ( .A1(n4818), .A2(n4821), .ZN(n8771) );
  AND2_X1 U5876 ( .A1(n4843), .A2(n4530), .ZN(n4322) );
  AND2_X1 U5877 ( .A1(n6900), .A2(n4495), .ZN(n4323) );
  INV_X1 U5878 ( .A(n8166), .ZN(n4595) );
  AND4_X1 U5879 ( .A1(n5005), .A2(n5004), .A3(n5003), .A4(n5386), .ZN(n4324)
         );
  OR2_X1 U5880 ( .A1(n9423), .A2(n9283), .ZN(n4325) );
  AND4_X1 U5881 ( .A1(n4989), .A2(n4988), .A3(n4987), .A4(n4986), .ZN(n4326)
         );
  OR2_X1 U5882 ( .A1(n5204), .A2(n7217), .ZN(n4327) );
  INV_X1 U5883 ( .A(n9190), .ZN(n4674) );
  AND2_X1 U5884 ( .A1(n5586), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n4328) );
  AND2_X1 U5885 ( .A1(n7682), .A2(n8155), .ZN(n4329) );
  AND2_X1 U5886 ( .A1(n8256), .A2(n8250), .ZN(n4330) );
  AND2_X1 U5887 ( .A1(n4806), .A2(n4804), .ZN(n4331) );
  AND2_X1 U5888 ( .A1(n7156), .A2(n7547), .ZN(n4332) );
  INV_X1 U5889 ( .A(n9185), .ZN(n4661) );
  NAND2_X1 U5890 ( .A1(n4417), .A2(n5963), .ZN(n8911) );
  INV_X1 U5891 ( .A(n7877), .ZN(n9588) );
  NAND2_X1 U5892 ( .A1(n5369), .A2(n5368), .ZN(n7877) );
  NAND2_X1 U5893 ( .A1(n6054), .A2(n6053), .ZN(n8988) );
  AND2_X1 U5894 ( .A1(n8076), .A2(n8214), .ZN(n4333) );
  INV_X1 U5895 ( .A(n9438), .ZN(n9341) );
  AND2_X1 U5896 ( .A1(n8074), .A2(n8212), .ZN(n4334) );
  NAND2_X1 U5897 ( .A1(n6398), .A2(n6397), .ZN(n9169) );
  INV_X1 U5898 ( .A(n4671), .ZN(n4670) );
  NAND2_X1 U5899 ( .A1(n6295), .A2(n9191), .ZN(n4671) );
  NAND2_X1 U5900 ( .A1(n7535), .A2(n5900), .ZN(n4335) );
  INV_X1 U5901 ( .A(n4644), .ZN(n4643) );
  NAND2_X1 U5902 ( .A1(n4294), .A2(n4646), .ZN(n4644) );
  OR2_X1 U5903 ( .A1(n8020), .A2(n8018), .ZN(n4336) );
  INV_X1 U5904 ( .A(n8210), .ZN(n4540) );
  INV_X1 U5905 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5033) );
  OR2_X1 U5906 ( .A1(n4698), .A2(n4707), .ZN(n4337) );
  INV_X1 U5907 ( .A(n6197), .ZN(n4707) );
  AND2_X1 U5908 ( .A1(n5433), .A2(n5434), .ZN(n4338) );
  INV_X1 U5909 ( .A(n4625), .ZN(n4624) );
  OAI21_X1 U5910 ( .B1(n4889), .B2(n4626), .A(n4893), .ZN(n4625) );
  NOR2_X1 U5911 ( .A1(n5509), .A2(n5508), .ZN(n4339) );
  NOR2_X1 U5912 ( .A1(n9580), .A2(n7913), .ZN(n4340) );
  NOR2_X1 U5913 ( .A1(n4859), .A2(n8435), .ZN(n4341) );
  AND2_X1 U5914 ( .A1(n4886), .A2(SI_5_), .ZN(n4342) );
  AND2_X1 U5915 ( .A1(n5911), .A2(n5910), .ZN(n4343) );
  AND2_X1 U5916 ( .A1(n5805), .A2(n5804), .ZN(n4344) );
  AND2_X1 U5917 ( .A1(n5715), .A2(n5714), .ZN(n4345) );
  NAND2_X1 U5918 ( .A1(n4316), .A2(n5405), .ZN(n4346) );
  AND2_X1 U5919 ( .A1(n4736), .A2(n5298), .ZN(n4347) );
  NOR2_X1 U5920 ( .A1(n8957), .A2(n8712), .ZN(n4348) );
  NAND2_X1 U5921 ( .A1(n5068), .A2(n4975), .ZN(n5144) );
  OR2_X1 U5922 ( .A1(n8926), .A2(n8183), .ZN(n4349) );
  INV_X1 U5923 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5755) );
  OR2_X1 U5924 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n4350) );
  INV_X1 U5925 ( .A(n4836), .ZN(n4835) );
  NAND2_X1 U5926 ( .A1(n7991), .A2(n7989), .ZN(n4836) );
  NOR2_X1 U5927 ( .A1(n5406), .A2(n5404), .ZN(n4351) );
  INV_X1 U5928 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6658) );
  OR2_X1 U5929 ( .A1(n8983), .A2(n8757), .ZN(n8214) );
  INV_X1 U5930 ( .A(n8214), .ZN(n4536) );
  AND2_X1 U5931 ( .A1(n4449), .A2(n7307), .ZN(n4352) );
  INV_X1 U5932 ( .A(n4419), .ZN(n4848) );
  NAND2_X1 U5933 ( .A1(n4908), .A2(n4909), .ZN(n4419) );
  INV_X1 U5934 ( .A(n4606), .ZN(n4605) );
  NOR2_X1 U5935 ( .A1(n4357), .A2(n8193), .ZN(n4606) );
  AND2_X1 U5936 ( .A1(n6141), .A2(n6140), .ZN(n4353) );
  OR2_X1 U5937 ( .A1(n6286), .A2(n6994), .ZN(n4354) );
  NAND2_X1 U5938 ( .A1(n7568), .A2(n4831), .ZN(n4355) );
  AND2_X1 U5939 ( .A1(n5406), .A2(n5405), .ZN(n4356) );
  OR2_X1 U5940 ( .A1(n8926), .A2(n8190), .ZN(n4357) );
  AND2_X1 U5941 ( .A1(n8129), .A2(n8128), .ZN(n4358) );
  INV_X1 U5942 ( .A(n5209), .ZN(n4626) );
  AND3_X1 U5943 ( .A1(n6345), .A2(n6343), .A3(n4558), .ZN(n4359) );
  AND2_X1 U5944 ( .A1(n4695), .A2(n4337), .ZN(n4360) );
  AND2_X1 U5945 ( .A1(n4793), .A2(n5033), .ZN(n4361) );
  AND2_X1 U5946 ( .A1(n5718), .A2(n4331), .ZN(n4362) );
  AND2_X1 U5947 ( .A1(n4292), .A2(n9084), .ZN(n4363) );
  INV_X1 U5948 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5719) );
  INV_X1 U5949 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n4723) );
  INV_X1 U5950 ( .A(n9081), .ZN(n4645) );
  INV_X1 U5951 ( .A(n6434), .ZN(n9163) );
  AOI21_X1 U5952 ( .B1(n9039), .B2(n6416), .A(n6415), .ZN(n6434) );
  INV_X1 U5953 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n4715) );
  NOR2_X1 U5954 ( .A1(n4722), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n5929) );
  NAND2_X1 U5955 ( .A1(n8521), .A2(n4709), .ZN(n8531) );
  NOR2_X1 U5956 ( .A1(n7043), .A2(n8877), .ZN(n4364) );
  NAND2_X1 U5957 ( .A1(n5694), .A2(n5693), .ZN(n9401) );
  INV_X1 U5958 ( .A(n9401), .ZN(n4585) );
  INV_X1 U5959 ( .A(n5344), .ZN(n5321) );
  INV_X1 U5960 ( .A(n8102), .ZN(n4834) );
  INV_X1 U5961 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n4806) );
  AND2_X1 U5962 ( .A1(n8947), .A2(n9016), .ZN(n4365) );
  OR3_X1 U5963 ( .A1(n8513), .A2(n8512), .A3(n8593), .ZN(n4366) );
  NAND2_X1 U5964 ( .A1(n5980), .A2(n5979), .ZN(n9015) );
  NAND2_X1 U5965 ( .A1(n6107), .A2(n6106), .ZN(n8966) );
  INV_X1 U5966 ( .A(n8966), .ZN(n4481) );
  INV_X1 U5967 ( .A(n8251), .ZN(n4531) );
  AND2_X1 U5968 ( .A1(n4980), .A2(n5174), .ZN(n5319) );
  NOR3_X1 U5969 ( .A1(n9371), .A2(n4579), .A3(n9429), .ZN(n4581) );
  NAND2_X1 U5970 ( .A1(n4803), .A2(n4805), .ZN(n5901) );
  NAND2_X1 U5971 ( .A1(n4551), .A2(n4550), .ZN(n7721) );
  XNOR2_X1 U5972 ( .A(n4733), .B(n6412), .ZN(n9039) );
  INV_X1 U5973 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n4716) );
  NAND2_X1 U5974 ( .A1(n7829), .A2(n4292), .ZN(n4573) );
  AND2_X1 U5975 ( .A1(n4507), .A2(n4311), .ZN(n4367) );
  NOR2_X1 U5976 ( .A1(n9245), .A2(n4585), .ZN(n4368) );
  INV_X1 U5977 ( .A(n4577), .ZN(n9320) );
  NOR2_X1 U5978 ( .A1(n9371), .A2(n4579), .ZN(n4577) );
  AND2_X1 U5979 ( .A1(n4951), .A2(SI_18_), .ZN(n4369) );
  AND2_X1 U5980 ( .A1(n4640), .A2(n4642), .ZN(n4370) );
  INV_X1 U5981 ( .A(n9248), .ZN(n9406) );
  NAND2_X1 U5982 ( .A1(n5610), .A2(n5609), .ZN(n9248) );
  INV_X1 U5983 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5742) );
  INV_X1 U5984 ( .A(n4827), .ZN(n4819) );
  INV_X1 U5985 ( .A(n9465), .ZN(n4571) );
  INV_X1 U5986 ( .A(n5631), .ZN(n5655) );
  XNOR2_X1 U5987 ( .A(n4999), .B(n5003), .ZN(n5658) );
  NAND2_X1 U5988 ( .A1(n7246), .A2(n6522), .ZN(n7289) );
  NAND2_X1 U5989 ( .A1(n5338), .A2(n5337), .ZN(n7650) );
  INV_X1 U5990 ( .A(n4518), .ZN(n4517) );
  OR2_X1 U5991 ( .A1(n7626), .A2(n4519), .ZN(n4518) );
  AND2_X1 U5992 ( .A1(n4520), .A2(n4517), .ZN(n4371) );
  NAND2_X1 U5993 ( .A1(n8004), .A2(n4470), .ZN(n4471) );
  AND2_X1 U5994 ( .A1(n6386), .A2(n6385), .ZN(n4372) );
  NAND2_X1 U5995 ( .A1(n7279), .A2(n7278), .ZN(n4373) );
  NAND2_X1 U5996 ( .A1(n7711), .A2(n8100), .ZN(n7778) );
  INV_X1 U5997 ( .A(n4500), .ZN(n6899) );
  NAND2_X1 U5998 ( .A1(n4502), .A2(n4501), .ZN(n4500) );
  AND2_X1 U5999 ( .A1(n4654), .A2(n7099), .ZN(n4374) );
  NAND2_X1 U6000 ( .A1(n4423), .A2(n8105), .ZN(n4422) );
  CLKBUF_X1 U6001 ( .A(n6305), .Z(n7034) );
  XOR2_X1 U6002 ( .A(n5910), .B(n5909), .Z(n4375) );
  NAND2_X1 U6003 ( .A1(n5260), .A2(n5259), .ZN(n6314) );
  INV_X1 U6004 ( .A(n6314), .ZN(n4574) );
  INV_X1 U6005 ( .A(n8638), .ZN(n4509) );
  INV_X1 U6006 ( .A(n9757), .ZN(n9298) );
  INV_X1 U6007 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5652) );
  XNOR2_X1 U6008 ( .A(n5749), .B(n5748), .ZN(n7496) );
  AND2_X1 U6009 ( .A1(n5650), .A2(n4361), .ZN(n9492) );
  INV_X1 U6010 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4615) );
  INV_X1 U6011 ( .A(n7661), .ZN(n7567) );
  NOR2_X1 U6012 ( .A1(n7138), .A2(n7661), .ZN(n7574) );
  OAI21_X1 U6013 ( .B1(n8153), .B2(n8257), .A(n8152), .ZN(n4381) );
  NOR2_X1 U6014 ( .A1(n8140), .A2(n4358), .ZN(n8132) );
  NAND2_X1 U6015 ( .A1(n4383), .A2(n8127), .ZN(n4382) );
  NAND2_X1 U6016 ( .A1(n8126), .A2(n8129), .ZN(n4385) );
  NAND2_X1 U6017 ( .A1(n8249), .A2(n8127), .ZN(n4390) );
  NAND2_X1 U6018 ( .A1(n4547), .A2(n4545), .ZN(n4393) );
  MUX2_X1 U6019 ( .A(n4366), .B(n4404), .S(n8518), .Z(n4403) );
  NAND2_X1 U6020 ( .A1(n5107), .A2(n4405), .ZN(n4869) );
  XNOR2_X1 U6021 ( .A(n5107), .B(n4405), .ZN(n6634) );
  XNOR2_X1 U6022 ( .A(n4867), .B(n4866), .ZN(n4405) );
  AOI21_X1 U6023 ( .B1(n5193), .B2(n4407), .A(n4342), .ZN(n4406) );
  INV_X1 U6024 ( .A(n5193), .ZN(n4408) );
  NAND3_X1 U6025 ( .A1(n4881), .A2(n4880), .A3(n5143), .ZN(n4409) );
  NAND2_X1 U6026 ( .A1(n8502), .A2(n6076), .ZN(n4410) );
  NAND2_X1 U6027 ( .A1(n8498), .A2(n6052), .ZN(n4411) );
  NAND3_X1 U6028 ( .A1(n4524), .A2(n4428), .A3(n4427), .ZN(n4426) );
  INV_X1 U6029 ( .A(n5527), .ZN(n4432) );
  NAND2_X1 U6030 ( .A1(n4435), .A2(n9110), .ZN(n4433) );
  AND2_X2 U6031 ( .A1(n9053), .A2(n9056), .ZN(n4434) );
  NAND2_X1 U6032 ( .A1(n5525), .A2(n5526), .ZN(n9109) );
  AND2_X2 U6033 ( .A1(n9110), .A2(n5527), .ZN(n4436) );
  OR2_X2 U6034 ( .A1(n5525), .A2(n5526), .ZN(n9110) );
  NAND3_X1 U6035 ( .A1(n4441), .A2(n4439), .A3(n4437), .ZN(P1_U3218) );
  NAND2_X1 U6036 ( .A1(n9135), .A2(n4440), .ZN(n4439) );
  OR2_X1 U6037 ( .A1(n9135), .A2(n4442), .ZN(n4441) );
  NAND2_X2 U6038 ( .A1(n9134), .A2(n5600), .ZN(n9135) );
  AND2_X2 U6039 ( .A1(n4445), .A2(n4356), .ZN(n8019) );
  AOI21_X2 U6040 ( .B1(n8308), .B2(n5274), .A(n4352), .ZN(n7481) );
  NAND2_X1 U6041 ( .A1(n8308), .A2(n8310), .ZN(n8309) );
  OAI21_X1 U6042 ( .B1(n8308), .B2(n4448), .A(n4446), .ZN(n4450) );
  OR2_X1 U6043 ( .A1(n5275), .A2(n7305), .ZN(n4449) );
  NOR2_X2 U6044 ( .A1(n9064), .A2(n9063), .ZN(n9101) );
  OAI21_X2 U6045 ( .B1(n4645), .B2(n4637), .A(n4636), .ZN(n9064) );
  NAND2_X1 U6046 ( .A1(n6728), .A2(n6730), .ZN(n5120) );
  AND2_X2 U6047 ( .A1(n7017), .A2(n5064), .ZN(n5247) );
  NAND3_X1 U6048 ( .A1(n4460), .A2(n4458), .A3(n4456), .ZN(P1_U3260) );
  INV_X1 U6049 ( .A(n4471), .ZN(n8929) );
  INV_X1 U6050 ( .A(n4475), .ZN(n8791) );
  OR2_X1 U6051 ( .A1(n6286), .A2(n6635), .ZN(n4478) );
  NAND3_X1 U6052 ( .A1(n4720), .A2(n5722), .A3(n4803), .ZN(n5737) );
  NAND3_X1 U6053 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_IR_REG_0__SCAN_IN), .ZN(n4499) );
  NAND3_X1 U6054 ( .A1(n7947), .A2(n4509), .A3(n4320), .ZN(n4506) );
  NAND2_X1 U6055 ( .A1(n4506), .A2(n4312), .ZN(n8637) );
  NAND2_X1 U6056 ( .A1(n7947), .A2(n6231), .ZN(n8634) );
  INV_X1 U6057 ( .A(n4507), .ZN(n8632) );
  INV_X1 U6058 ( .A(n8633), .ZN(n4508) );
  NAND2_X1 U6059 ( .A1(n4520), .A2(n4522), .ZN(n7625) );
  INV_X1 U6060 ( .A(n4522), .ZN(n4519) );
  NAND2_X1 U6061 ( .A1(n8240), .A2(n4533), .ZN(n4529) );
  NAND2_X1 U6062 ( .A1(n4529), .A2(n4322), .ZN(n8252) );
  NAND2_X1 U6063 ( .A1(n4534), .A2(n4535), .ZN(n8206) );
  NAND3_X1 U6064 ( .A1(n8203), .A2(n4538), .A3(n4291), .ZN(n4534) );
  NAND2_X1 U6065 ( .A1(n4881), .A2(n4880), .ZN(n4554) );
  XNOR2_X1 U6066 ( .A(n4554), .B(n4553), .ZN(n6632) );
  INV_X1 U6067 ( .A(n5143), .ZN(n4553) );
  NAND2_X1 U6068 ( .A1(n5172), .A2(n5173), .ZN(n4890) );
  NAND2_X1 U6069 ( .A1(n5172), .A2(n4555), .ZN(n4623) );
  NAND3_X1 U6070 ( .A1(n6344), .A2(n4359), .A3(n4556), .ZN(n6346) );
  NAND3_X1 U6071 ( .A1(n6321), .A2(n6342), .A3(n4557), .ZN(n4556) );
  INV_X1 U6072 ( .A(n4785), .ZN(n4560) );
  AOI21_X2 U6073 ( .B1(n6433), .B2(n6483), .A(n4565), .ZN(n6553) );
  AND2_X1 U6074 ( .A1(n4566), .A2(n7118), .ZN(n9737) );
  NAND2_X1 U6075 ( .A1(n4567), .A2(n6441), .ZN(n9779) );
  XNOR2_X2 U6076 ( .A(n6693), .B(n4568), .ZN(n7023) );
  AND4_X2 U6077 ( .A1(n5115), .A2(n5116), .A3(n5113), .A4(n5114), .ZN(n6693)
         );
  OAI21_X1 U6078 ( .B1(n4570), .B2(n4569), .A(n6367), .ZN(n6376) );
  INV_X1 U6079 ( .A(n4573), .ZN(n7975) );
  NAND3_X1 U6080 ( .A1(n9750), .A2(n4575), .A3(n4574), .ZN(n4576) );
  INV_X1 U6081 ( .A(n4576), .ZN(n7329) );
  INV_X1 U6082 ( .A(n4581), .ZN(n9306) );
  NAND2_X1 U6083 ( .A1(n5792), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n6923) );
  INV_X1 U6084 ( .A(n7731), .ZN(n4588) );
  NAND2_X1 U6085 ( .A1(n4587), .A2(n8155), .ZN(n7684) );
  NAND3_X1 U6086 ( .A1(n7681), .A2(n4588), .A3(n8154), .ZN(n4587) );
  NAND2_X1 U6087 ( .A1(n7571), .A2(n8092), .ZN(n7681) );
  OAI21_X2 U6088 ( .B1(n7570), .B2(n8131), .A(n8142), .ZN(n7571) );
  AND2_X1 U6089 ( .A1(n8149), .A2(n8154), .ZN(n8092) );
  OAI21_X1 U6090 ( .B1(n7711), .B2(n4590), .A(n4589), .ZN(n7995) );
  NAND2_X1 U6091 ( .A1(n4593), .A2(n4591), .ZN(n7996) );
  NAND2_X1 U6092 ( .A1(n7711), .A2(n4594), .ZN(n4593) );
  XNOR2_X1 U6093 ( .A(n4600), .B(n4284), .ZN(n4599) );
  NAND2_X1 U6094 ( .A1(n4601), .A2(n8246), .ZN(n4600) );
  OAI21_X1 U6095 ( .B1(n8083), .B2(n4602), .A(n4330), .ZN(n4601) );
  NAND2_X1 U6096 ( .A1(n8899), .A2(n4314), .ZN(n4604) );
  AOI211_X2 U6097 ( .C1(n8755), .C2(n4610), .A(n4608), .B(n8079), .ZN(n8709)
         );
  NAND2_X1 U6098 ( .A1(n4803), .A2(n4613), .ZN(n4722) );
  NOR2_X1 U6099 ( .A1(n5798), .A2(P2_IR_REG_11__SCAN_IN), .ZN(n4613) );
  OR2_X1 U6100 ( .A1(n5797), .A2(n6637), .ZN(n5772) );
  OR2_X1 U6101 ( .A1(n6082), .A2(n6636), .ZN(n5773) );
  NAND2_X1 U6102 ( .A1(n7133), .A2(n8129), .ZN(n7570) );
  NAND2_X1 U6103 ( .A1(n7072), .A2(n8373), .ZN(n9918) );
  NAND3_X1 U6104 ( .A1(n8307), .A2(n4615), .A3(n4614), .ZN(n4863) );
  NAND2_X1 U6105 ( .A1(n4623), .A2(n4622), .ZN(n5229) );
  NAND2_X1 U6106 ( .A1(n4890), .A2(n4889), .ZN(n5210) );
  NAND2_X1 U6107 ( .A1(n5338), .A2(n4630), .ZN(n4629) );
  INV_X1 U6108 ( .A(n4647), .ZN(n9079) );
  MUX2_X1 U6109 ( .A(n6631), .B(n6624), .S(n4278), .Z(n4882) );
  MUX2_X1 U6110 ( .A(n6628), .B(n6626), .S(n4283), .Z(n4885) );
  MUX2_X1 U6111 ( .A(n6639), .B(n6642), .S(n4283), .Z(n4887) );
  MUX2_X1 U6112 ( .A(n6652), .B(n6651), .S(n4283), .Z(n4895) );
  MUX2_X1 U6113 ( .A(n6653), .B(n6656), .S(n4278), .Z(n4900) );
  NAND2_X1 U6114 ( .A1(n4654), .A2(n4653), .ZN(n7164) );
  INV_X1 U6115 ( .A(n7289), .ZN(n4656) );
  OAI21_X1 U6116 ( .B1(n8035), .B2(n4658), .A(n4657), .ZN(n9358) );
  NAND2_X1 U6117 ( .A1(n9327), .A2(n4666), .ZN(n4664) );
  AND2_X1 U6118 ( .A1(n5319), .A2(n4684), .ZN(n5409) );
  NAND2_X1 U6119 ( .A1(n4683), .A2(n5319), .ZN(n4990) );
  NAND2_X1 U6120 ( .A1(n4685), .A2(n8133), .ZN(n5752) );
  NAND2_X1 U6121 ( .A1(n6911), .A2(n4685), .ZN(n6914) );
  NAND2_X1 U6122 ( .A1(n7534), .A2(n4688), .ZN(n4687) );
  AND2_X1 U6123 ( .A1(n7044), .A2(n5803), .ZN(n4692) );
  NAND2_X1 U6124 ( .A1(n8583), .A2(n4360), .ZN(n4693) );
  OAI211_X1 U6125 ( .C1(n8583), .C2(n4694), .A(n4706), .B(n4693), .ZN(P2_U3222) );
  OAI21_X1 U6126 ( .B1(n8583), .B2(n8582), .A(n4708), .ZN(n8463) );
  AOI21_X1 U6127 ( .B1(n4711), .B2(n8530), .A(n8593), .ZN(n8532) );
  NAND2_X1 U6128 ( .A1(n8487), .A2(n4712), .ZN(n8498) );
  NAND2_X1 U6129 ( .A1(n8405), .A2(n4714), .ZN(n6569) );
  NAND2_X1 U6130 ( .A1(n5744), .A2(n4724), .ZN(n6155) );
  NAND2_X1 U6131 ( .A1(n5744), .A2(n5740), .ZN(n5741) );
  NAND3_X1 U6132 ( .A1(n4725), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n4862) );
  NAND2_X1 U6133 ( .A1(n4949), .A2(n4729), .ZN(n4728) );
  NAND3_X1 U6134 ( .A1(n4731), .A2(n5435), .A3(n4730), .ZN(n4727) );
  NAND3_X1 U6135 ( .A1(n4736), .A2(n4739), .A3(n5298), .ZN(n4735) );
  NAND2_X1 U6136 ( .A1(n5691), .A2(n5690), .ZN(n4743) );
  OAI21_X1 U6137 ( .B1(n4295), .B2(n4749), .A(n4747), .ZN(n4943) );
  NAND2_X1 U6138 ( .A1(n4962), .A2(n4961), .ZN(n5493) );
  NAND2_X1 U6139 ( .A1(n4962), .A2(n4751), .ZN(n4750) );
  OAI21_X1 U6140 ( .B1(n5549), .B2(n4767), .A(n5553), .ZN(n5577) );
  NAND2_X1 U6141 ( .A1(n5549), .A2(n4765), .ZN(n4764) );
  NAND2_X1 U6142 ( .A1(n9319), .A2(n4773), .ZN(n4768) );
  NAND2_X1 U6143 ( .A1(n4768), .A2(n4770), .ZN(n9275) );
  NAND2_X1 U6144 ( .A1(n5650), .A2(n4793), .ZN(n5032) );
  NAND2_X1 U6145 ( .A1(n5650), .A2(n5652), .ZN(n5027) );
  NAND2_X1 U6146 ( .A1(n9239), .A2(n9238), .ZN(n9237) );
  NAND2_X1 U6147 ( .A1(n7841), .A2(n4799), .ZN(n4797) );
  NAND2_X1 U6148 ( .A1(n4797), .A2(n4798), .ZN(n7970) );
  AND3_X2 U6149 ( .A1(n5718), .A2(n4331), .A3(n4851), .ZN(n4803) );
  NAND3_X1 U6150 ( .A1(n4805), .A2(n5718), .A3(n4806), .ZN(n5860) );
  NAND2_X1 U6151 ( .A1(n8706), .A2(n4809), .ZN(n4808) );
  NAND2_X1 U6152 ( .A1(n7688), .A2(n4812), .ZN(n9990) );
  INV_X1 U6153 ( .A(n8856), .ZN(n4817) );
  NAND3_X1 U6154 ( .A1(n4816), .A2(n4814), .A3(n4827), .ZN(n8760) );
  NAND3_X1 U6155 ( .A1(n4816), .A2(n4815), .A3(n4814), .ZN(n8762) );
  OR2_X1 U6156 ( .A1(n8983), .A2(n8801), .ZN(n4827) );
  NAND2_X1 U6157 ( .A1(n7080), .A2(n8091), .ZN(n7569) );
  NAND2_X1 U6158 ( .A1(n4829), .A2(n4828), .ZN(n7732) );
  NAND2_X1 U6159 ( .A1(n7080), .A2(n4830), .ZN(n4829) );
  NOR2_X1 U6160 ( .A1(n5737), .A2(n4299), .ZN(n5753) );
  NAND2_X1 U6161 ( .A1(n5096), .A2(n4865), .ZN(n4867) );
  OAI22_X1 U6162 ( .A1(n9782), .A2(n5093), .B1(n9836), .B2(n5570), .ZN(n5198)
         );
  NAND2_X1 U6163 ( .A1(n6417), .A2(n9163), .ZN(n6487) );
  AND2_X2 U6164 ( .A1(n9773), .A2(n9836), .ZN(n9750) );
  INV_X1 U6165 ( .A(n9169), .ZN(n9394) );
  NOR2_X1 U6166 ( .A1(n6305), .A2(n7176), .ZN(n7254) );
  NAND2_X1 U6167 ( .A1(n5201), .A2(n4327), .ZN(n5206) );
  XNOR2_X1 U6168 ( .A(n5210), .B(n5209), .ZN(n6648) );
  NOR2_X1 U6169 ( .A1(n4328), .A2(n4847), .ZN(n5189) );
  OAI21_X1 U6170 ( .B1(n5717), .B2(n5657), .A(n9136), .ZN(n5689) );
  CLKBUF_X1 U6171 ( .A(n5632), .Z(n6705) );
  INV_X1 U6172 ( .A(n9733), .ZN(n9782) );
  NOR4_X1 U6173 ( .A1(n6547), .A2(n6517), .A3(n6543), .A4(n6516), .ZN(n6518)
         );
  NAND2_X1 U6174 ( .A1(n8137), .A2(n7075), .ZN(n7085) );
  NOR2_X1 U6175 ( .A1(n6155), .A2(n6154), .ZN(n6159) );
  AOI21_X1 U6176 ( .B1(n8470), .B2(n6099), .A(n6098), .ZN(n6105) );
  NAND2_X1 U6177 ( .A1(n8268), .A2(n8118), .ZN(n6912) );
  NAND2_X1 U6178 ( .A1(n5602), .A2(n5601), .ZN(n5604) );
  NAND2_X1 U6179 ( .A1(n6162), .A2(n6161), .ZN(n6163) );
  INV_X1 U6180 ( .A(n8039), .ZN(n7974) );
  INV_X1 U6181 ( .A(n6286), .ZN(n6022) );
  NAND2_X1 U6182 ( .A1(n7897), .A2(n7898), .ZN(n7772) );
  NAND2_X1 U6183 ( .A1(n7190), .A2(n7151), .ZN(n7319) );
  AND2_X1 U6184 ( .A1(n4288), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n4839) );
  OR2_X1 U6185 ( .A1(n9341), .A2(n9363), .ZN(n4840) );
  OR2_X1 U6186 ( .A1(n9325), .A2(n9315), .ZN(n4842) );
  AND2_X1 U6187 ( .A1(n8441), .A2(n8243), .ZN(n4843) );
  AND2_X1 U6188 ( .A1(n4588), .A2(n4850), .ZN(n4844) );
  AND2_X1 U6189 ( .A1(n7334), .A2(n9156), .ZN(n4845) );
  AND2_X1 U6190 ( .A1(n6274), .A2(n6273), .ZN(n4846) );
  AND2_X1 U6191 ( .A1(n4290), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n4847) );
  NAND2_X1 U6192 ( .A1(n7648), .A2(n9757), .ZN(n6430) );
  NAND2_X2 U6193 ( .A1(n7103), .A2(n9792), .ZN(n9797) );
  INV_X1 U6194 ( .A(n5658), .ZN(n5660) );
  AND2_X1 U6195 ( .A1(n8180), .A2(n8178), .ZN(n9908) );
  INV_X1 U6196 ( .A(n9908), .ZN(n7991) );
  INV_X1 U6197 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n5036) );
  AND2_X1 U6198 ( .A1(n7682), .A2(n8161), .ZN(n4849) );
  OR2_X1 U6199 ( .A1(n8154), .A2(n8257), .ZN(n4850) );
  NOR2_X1 U6200 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n4851) );
  AND2_X1 U6201 ( .A1(n6487), .A2(n6420), .ZN(n4852) );
  NAND2_X1 U6202 ( .A1(n9002), .A2(n8851), .ZN(n4853) );
  NOR2_X1 U6203 ( .A1(n9002), .A2(n8851), .ZN(n4854) );
  NAND2_X1 U6204 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), 
        .ZN(n4855) );
  AND2_X1 U6205 ( .A1(n8437), .A2(n8226), .ZN(n4856) );
  OR2_X1 U6206 ( .A1(n6568), .A2(n5098), .ZN(n4857) );
  AND2_X1 U6207 ( .A1(n5629), .A2(n5630), .ZN(n4858) );
  XNOR2_X1 U6208 ( .A(n5198), .B(n5247), .ZN(n5204) );
  NOR2_X1 U6209 ( .A1(n8988), .A2(n8808), .ZN(n4859) );
  OR2_X1 U6210 ( .A1(n8619), .A2(n7531), .ZN(n4860) );
  NAND2_X1 U6211 ( .A1(n6810), .A2(n5161), .ZN(n6886) );
  AND2_X1 U6212 ( .A1(n8426), .A2(n8610), .ZN(n4861) );
  NOR2_X1 U6213 ( .A1(n8427), .A2(n4861), .ZN(n8924) );
  NAND2_X1 U6214 ( .A1(n5931), .A2(n5930), .ZN(n8426) );
  INV_X1 U6215 ( .A(n8426), .ZN(n8003) );
  INV_X1 U6216 ( .A(n8257), .ZN(n8127) );
  AOI21_X1 U6217 ( .B1(n8198), .B2(n8858), .A(n8197), .ZN(n8209) );
  NOR2_X1 U6218 ( .A1(n6480), .A2(n6418), .ZN(n6419) );
  AOI21_X1 U6219 ( .B1(n9398), .B2(n6418), .A(n6419), .ZN(n6420) );
  AND2_X1 U6220 ( .A1(n4302), .A2(n8244), .ZN(n8245) );
  INV_X1 U6221 ( .A(n7689), .ZN(n7682) );
  INV_X1 U6222 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5721) );
  INV_X1 U6223 ( .A(n9151), .ZN(n7913) );
  INV_X1 U6224 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n4991) );
  INV_X1 U6225 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5883) );
  INV_X1 U6226 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5720) );
  NAND2_X1 U6227 ( .A1(n9815), .A2(n6307), .ZN(n6522) );
  AND4_X1 U6228 ( .A1(n4979), .A2(n4978), .A3(n5211), .A4(n4977), .ZN(n4980)
         );
  NOR2_X1 U6229 ( .A1(n6100), .A2(n8544), .ZN(n6098) );
  NAND2_X1 U6230 ( .A1(n8254), .A2(n8257), .ZN(n8255) );
  INV_X1 U6231 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6164) );
  INV_X1 U6232 ( .A(n5514), .ZN(n5023) );
  INV_X1 U6233 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n7268) );
  OR2_X1 U6234 ( .A1(n5584), .A2(n9143), .ZN(n5673) );
  INV_X1 U6235 ( .A(n5370), .ZN(n5019) );
  INV_X1 U6236 ( .A(SI_23_), .ZN(n7462) );
  INV_X1 U6237 ( .A(SI_20_), .ZN(n7387) );
  INV_X1 U6238 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5007) );
  INV_X1 U6239 ( .A(SI_13_), .ZN(n4919) );
  INV_X1 U6240 ( .A(n6570), .ZN(n5851) );
  OR2_X1 U6241 ( .A1(n6134), .A2(n8464), .ZN(n6146) );
  OR2_X1 U6242 ( .A1(n8413), .A2(n7043), .ZN(n5764) );
  OR2_X1 U6243 ( .A1(n6090), .A2(n8473), .ZN(n6092) );
  INV_X1 U6244 ( .A(n9050), .ZN(n5735) );
  OR2_X1 U6245 ( .A1(n8966), .A2(n8711), .ZN(n8438) );
  INV_X1 U6246 ( .A(n8752), .ZN(n8076) );
  INV_X1 U6247 ( .A(n7997), .ZN(n8180) );
  INV_X1 U6248 ( .A(n7131), .ZN(n7135) );
  INV_X1 U6249 ( .A(n8004), .ZN(n9912) );
  OR2_X1 U6250 ( .A1(n9939), .A2(n6906), .ZN(n6907) );
  INV_X1 U6251 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5754) );
  INV_X1 U6252 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n5057) );
  NAND2_X1 U6253 ( .A1(n5023), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n5516) );
  NAND2_X1 U6254 ( .A1(n5022), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5474) );
  OR2_X1 U6255 ( .A1(n5281), .A2(n7268), .ZN(n5304) );
  AND2_X1 U6256 ( .A1(n5673), .A2(n5585), .ZN(n9260) );
  OR2_X1 U6257 ( .A1(n5393), .A2(n5392), .ZN(n5414) );
  INV_X1 U6258 ( .A(n7204), .ZN(n7156) );
  INV_X1 U6259 ( .A(n5663), .ZN(n5633) );
  OR2_X1 U6260 ( .A1(n4902), .A2(n4901), .ZN(n4903) );
  NAND2_X1 U6261 ( .A1(n4283), .A2(n6623), .ZN(n4874) );
  OR2_X1 U6262 ( .A1(n6082), .A2(n8052), .ZN(n6132) );
  OR2_X1 U6263 ( .A1(n6196), .A2(n6195), .ZN(n6197) );
  OR2_X1 U6264 ( .A1(n6056), .A2(n6055), .ZN(n6066) );
  OR2_X1 U6265 ( .A1(n6012), .A2(n8577), .ZN(n6042) );
  OR2_X1 U6266 ( .A1(n7496), .A2(n8133), .ZN(n8089) );
  OR2_X1 U6267 ( .A1(n7749), .A2(n4615), .ZN(n6290) );
  INV_X1 U6268 ( .A(n8238), .ZN(n8680) );
  OR2_X1 U6269 ( .A1(n6082), .A2(n8015), .ZN(n6120) );
  INV_X1 U6270 ( .A(n8975), .ZN(n8767) );
  INV_X1 U6271 ( .A(n6912), .ZN(n6236) );
  INV_X1 U6272 ( .A(n8133), .ZN(n8118) );
  NAND2_X1 U6273 ( .A1(n8161), .A2(n8155), .ZN(n7731) );
  AND2_X1 U6274 ( .A1(n9953), .A2(n6911), .ZN(n9016) );
  NOR2_X1 U6275 ( .A1(n7519), .A2(n6907), .ZN(n6908) );
  INV_X1 U6276 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6166) );
  INV_X1 U6277 ( .A(n9293), .ZN(n9266) );
  AND2_X1 U6278 ( .A1(n9137), .A2(n9133), .ZN(n5600) );
  OR2_X1 U6279 ( .A1(n5166), .A2(n7032), .ZN(n5116) );
  INV_X1 U6280 ( .A(n9346), .ZN(n9315) );
  AND2_X1 U6281 ( .A1(n6497), .A2(n9185), .ZN(n8041) );
  AOI21_X1 U6282 ( .B1(n7319), .B2(n7152), .A(n4845), .ZN(n7153) );
  NAND2_X1 U6283 ( .A1(n7150), .A2(n7149), .ZN(n7190) );
  AND2_X1 U6284 ( .A1(n6499), .A2(n7920), .ZN(n7842) );
  AND2_X1 U6285 ( .A1(n6710), .A2(n5633), .ZN(n9856) );
  INV_X1 U6286 ( .A(n9734), .ZN(n9784) );
  OR2_X1 U6287 ( .A1(n6430), .A2(n5660), .ZN(n9818) );
  NAND2_X1 U6288 ( .A1(n6689), .A2(n6688), .ZN(n6716) );
  XNOR2_X1 U6289 ( .A(n5653), .B(n5652), .ZN(n6558) );
  AND2_X1 U6290 ( .A1(n4942), .A2(n4941), .ZN(n5408) );
  AND2_X1 U6291 ( .A1(n4923), .A2(n4922), .ZN(n5342) );
  AND2_X1 U6292 ( .A1(n6201), .A2(n8265), .ZN(n8509) );
  NAND2_X1 U6293 ( .A1(n8378), .A2(n8376), .ZN(n8372) );
  INV_X1 U6294 ( .A(n8585), .ZN(n8601) );
  OR2_X1 U6295 ( .A1(n7865), .A2(n6238), .ZN(n6241) );
  AND4_X1 U6296 ( .A1(n6047), .A2(n6046), .A3(n6045), .A4(n6044), .ZN(n8833)
         );
  NAND2_X1 U6297 ( .A1(n6290), .A2(n6289), .ZN(n6291) );
  INV_X1 U6298 ( .A(n8427), .ZN(n7994) );
  INV_X1 U6299 ( .A(n8918), .ZN(n9934) );
  AND2_X1 U6300 ( .A1(n6175), .A2(n6174), .ZN(n7514) );
  INV_X1 U6301 ( .A(n9016), .ZN(n10019) );
  AND2_X1 U6302 ( .A1(n8883), .A2(n9541), .ZN(n10001) );
  INV_X1 U6303 ( .A(n10001), .ZN(n10025) );
  INV_X1 U6304 ( .A(n7514), .ZN(n6910) );
  OAI21_X1 U6305 ( .B1(n9406), .B2(n9148), .A(n5686), .ZN(n5687) );
  AND2_X1 U6306 ( .A1(n5043), .A2(n5042), .ZN(n9179) );
  OR2_X1 U6307 ( .A1(n6597), .A2(n8031), .ZN(n8305) );
  INV_X1 U6308 ( .A(n9681), .ZN(n9714) );
  INV_X1 U6309 ( .A(n9717), .ZN(n9688) );
  AND2_X1 U6310 ( .A1(n4674), .A2(n9191), .ZN(n9326) );
  AND2_X1 U6311 ( .A1(n6498), .A2(n9187), .ZN(n9378) );
  NAND2_X1 U6312 ( .A1(n6457), .A2(n6460), .ZN(n7969) );
  AND2_X1 U6313 ( .A1(n9797), .A2(n9298), .ZN(n9350) );
  INV_X1 U6314 ( .A(n9864), .ZN(n7334) );
  AND2_X1 U6315 ( .A1(n7025), .A2(n7024), .ZN(n9734) );
  AND2_X1 U6316 ( .A1(n9350), .A2(n9857), .ZN(n9777) );
  INV_X1 U6317 ( .A(n9856), .ZN(n9863) );
  INV_X1 U6318 ( .A(n9853), .ZN(n9472) );
  NAND2_X1 U6319 ( .A1(n9789), .A2(n9818), .ZN(n9853) );
  AND2_X1 U6320 ( .A1(n6707), .A2(n6706), .ZN(n6718) );
  AND2_X1 U6321 ( .A1(n6558), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5654) );
  AND2_X1 U6322 ( .A1(n5258), .A2(n5257), .ZN(n6745) );
  AND2_X1 U6323 ( .A1(n4283), .A2(P1_U3084), .ZN(n8053) );
  INV_X1 U6324 ( .A(n7749), .ZN(n9892) );
  OR2_X1 U6325 ( .A1(n8676), .A2(n8585), .ZN(n6212) );
  NAND2_X1 U6326 ( .A1(n8509), .A2(n8862), .ZN(n8597) );
  INV_X1 U6327 ( .A(n8911), .ZN(n9529) );
  INV_X1 U6328 ( .A(n8431), .ZN(n8808) );
  INV_X1 U6329 ( .A(n8832), .ZN(n8863) );
  INV_X1 U6330 ( .A(n7074), .ZN(n8620) );
  NAND2_X1 U6331 ( .A1(n6244), .A2(n6243), .ZN(n9895) );
  INV_X1 U6332 ( .A(n9888), .ZN(n9894) );
  OR2_X1 U6333 ( .A1(n9937), .A2(n7527), .ZN(n9906) );
  INV_X1 U6334 ( .A(n8916), .ZN(n8932) );
  OR2_X1 U6335 ( .A1(n9937), .A2(n7707), .ZN(n8893) );
  INV_X2 U6336 ( .A(n8916), .ZN(n9937) );
  INV_X1 U6337 ( .A(n10045), .ZN(n10042) );
  INV_X1 U6338 ( .A(n10028), .ZN(n10026) );
  NOR2_X1 U6339 ( .A1(n9939), .A2(n9938), .ZN(n9944) );
  AND2_X1 U6340 ( .A1(n8017), .A2(n6237), .ZN(n9947) );
  INV_X1 U6341 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7946) );
  INV_X1 U6342 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7038) );
  INV_X1 U6343 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6669) );
  INV_X1 U6344 ( .A(n9136), .ZN(n9131) );
  INV_X1 U6345 ( .A(n9245), .ZN(n9208) );
  INV_X1 U6346 ( .A(n9179), .ZN(n9329) );
  INV_X1 U6347 ( .A(n7982), .ZN(n9150) );
  OR2_X1 U6348 ( .A1(n8305), .A2(n5671), .ZN(n9681) );
  OR3_X1 U6349 ( .A1(n6597), .A2(n5671), .A3(n6596), .ZN(n9724) );
  OR2_X1 U6350 ( .A1(P1_U3083), .A2(n6790), .ZN(n9727) );
  INV_X1 U6351 ( .A(n9797), .ZN(n9383) );
  INV_X1 U6352 ( .A(n9797), .ZN(n9568) );
  INV_X1 U6353 ( .A(n9887), .ZN(n9885) );
  INV_X1 U6354 ( .A(n9872), .ZN(n9871) );
  INV_X1 U6355 ( .A(n9809), .ZN(n9808) );
  NAND2_X1 U6356 ( .A1(n6688), .A2(n6701), .ZN(n9809) );
  INV_X1 U6357 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n8013) );
  INV_X1 U6358 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7649) );
  INV_X1 U6359 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6684) );
  INV_X1 U6360 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6667) );
  NOR2_X1 U6361 ( .A1(n10073), .A2(n10072), .ZN(n10071) );
  OAI21_X1 U6362 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10062), .ZN(n10060) );
  INV_X2 U6363 ( .A(n6760), .ZN(P2_U3966) );
  NAND2_X1 U6364 ( .A1(n6294), .A2(n6293), .ZN(P2_U3264) );
  NOR2_X1 U6365 ( .A1(n6613), .A2(P1_U3084), .ZN(P1_U4006) );
  AND2_X1 U6366 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n4864) );
  NAND2_X1 U6367 ( .A1(n4277), .A2(n4864), .ZN(n5096) );
  NAND3_X1 U6368 ( .A1(n4873), .A2(SI_0_), .A3(P1_DATAO_REG_0__SCAN_IN), .ZN(
        n4865) );
  INV_X1 U6369 ( .A(SI_1_), .ZN(n4866) );
  MUX2_X1 U6370 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(P1_DATAO_REG_1__SCAN_IN), 
        .S(n4873), .Z(n5107) );
  NAND2_X1 U6371 ( .A1(n4867), .A2(SI_1_), .ZN(n4868) );
  NAND2_X1 U6372 ( .A1(n4869), .A2(n4868), .ZN(n5067) );
  INV_X1 U6373 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6636) );
  INV_X1 U6374 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n4870) );
  MUX2_X1 U6375 ( .A(n6636), .B(n4870), .S(n4277), .Z(n4871) );
  XNOR2_X1 U6376 ( .A(n4871), .B(SI_2_), .ZN(n5066) );
  NAND2_X1 U6377 ( .A1(n5067), .A2(n5066), .ZN(n5127) );
  INV_X1 U6378 ( .A(n4871), .ZN(n4872) );
  NAND2_X1 U6379 ( .A1(n4872), .A2(SI_2_), .ZN(n5126) );
  INV_X1 U6380 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6629) );
  INV_X1 U6381 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6623) );
  INV_X1 U6382 ( .A(n4878), .ZN(n4875) );
  NAND2_X1 U6383 ( .A1(n4875), .A2(SI_3_), .ZN(n4877) );
  AND2_X1 U6384 ( .A1(n5126), .A2(n4877), .ZN(n4876) );
  NAND2_X1 U6385 ( .A1(n5127), .A2(n4876), .ZN(n4881) );
  INV_X1 U6386 ( .A(n4877), .ZN(n4879) );
  XNOR2_X1 U6387 ( .A(n4878), .B(SI_3_), .ZN(n5129) );
  INV_X1 U6388 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6631) );
  INV_X1 U6389 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6624) );
  XNOR2_X1 U6390 ( .A(n4882), .B(SI_4_), .ZN(n5143) );
  INV_X1 U6391 ( .A(n4882), .ZN(n4883) );
  NAND2_X1 U6392 ( .A1(n4883), .A2(SI_4_), .ZN(n4884) );
  INV_X1 U6393 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6628) );
  INV_X1 U6394 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6626) );
  XNOR2_X1 U6395 ( .A(n4885), .B(SI_5_), .ZN(n5193) );
  INV_X1 U6396 ( .A(n4885), .ZN(n4886) );
  INV_X1 U6397 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6639) );
  INV_X1 U6398 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6642) );
  XNOR2_X1 U6399 ( .A(n4887), .B(SI_6_), .ZN(n5173) );
  INV_X1 U6400 ( .A(n4887), .ZN(n4888) );
  NAND2_X1 U6401 ( .A1(n4888), .A2(SI_6_), .ZN(n4889) );
  INV_X1 U6402 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6649) );
  MUX2_X1 U6403 ( .A(n6646), .B(n6649), .S(n4278), .Z(n4891) );
  XNOR2_X1 U6404 ( .A(n4891), .B(SI_7_), .ZN(n5209) );
  INV_X1 U6405 ( .A(n4891), .ZN(n4892) );
  NAND2_X1 U6406 ( .A1(n4892), .A2(SI_7_), .ZN(n4893) );
  INV_X1 U6407 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6652) );
  INV_X1 U6408 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6651) );
  INV_X1 U6409 ( .A(SI_8_), .ZN(n4894) );
  NAND2_X1 U6410 ( .A1(n4895), .A2(n4894), .ZN(n5228) );
  INV_X1 U6411 ( .A(n4895), .ZN(n4896) );
  NAND2_X1 U6412 ( .A1(n4896), .A2(SI_8_), .ZN(n4897) );
  NAND2_X1 U6413 ( .A1(n5228), .A2(n4897), .ZN(n5252) );
  INV_X1 U6414 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6656) );
  INV_X1 U6415 ( .A(n4900), .ZN(n4898) );
  NAND2_X1 U6416 ( .A1(n4898), .A2(SI_9_), .ZN(n5230) );
  INV_X1 U6417 ( .A(n5230), .ZN(n4902) );
  INV_X1 U6418 ( .A(SI_9_), .ZN(n4899) );
  NAND2_X1 U6419 ( .A1(n4900), .A2(n4899), .ZN(n5231) );
  AND2_X1 U6420 ( .A1(n5228), .A2(n5231), .ZN(n4901) );
  INV_X1 U6421 ( .A(SI_10_), .ZN(n4905) );
  INV_X1 U6422 ( .A(n4906), .ZN(n4907) );
  NAND2_X1 U6423 ( .A1(n4907), .A2(SI_10_), .ZN(n4908) );
  MUX2_X1 U6424 ( .A(n6669), .B(n6667), .S(n4283), .Z(n4910) );
  XNOR2_X1 U6425 ( .A(n4910), .B(SI_11_), .ZN(n5298) );
  INV_X1 U6426 ( .A(n4910), .ZN(n4911) );
  NAND2_X1 U6427 ( .A1(n4911), .A2(SI_11_), .ZN(n4912) );
  MUX2_X1 U6428 ( .A(n6678), .B(n6675), .S(n4283), .Z(n4914) );
  INV_X1 U6429 ( .A(SI_12_), .ZN(n4913) );
  NAND2_X1 U6430 ( .A1(n4914), .A2(n4913), .ZN(n4917) );
  INV_X1 U6431 ( .A(n4914), .ZN(n4915) );
  NAND2_X1 U6432 ( .A1(n4915), .A2(SI_12_), .ZN(n4916) );
  NAND2_X1 U6433 ( .A1(n4917), .A2(n4916), .ZN(n5317) );
  INV_X1 U6434 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n4918) );
  MUX2_X1 U6435 ( .A(n7440), .B(n4918), .S(n4283), .Z(n4920) );
  NAND2_X1 U6436 ( .A1(n4920), .A2(n4919), .ZN(n4923) );
  INV_X1 U6437 ( .A(n4920), .ZN(n4921) );
  NAND2_X1 U6438 ( .A1(n4921), .A2(SI_13_), .ZN(n4922) );
  NAND2_X1 U6439 ( .A1(n5343), .A2(n5342), .ZN(n4924) );
  NAND2_X1 U6440 ( .A1(n4924), .A2(n4923), .ZN(n5364) );
  MUX2_X1 U6441 ( .A(n6687), .B(n6684), .S(n4283), .Z(n4926) );
  XNOR2_X1 U6442 ( .A(n4926), .B(SI_14_), .ZN(n5363) );
  INV_X1 U6443 ( .A(n5363), .ZN(n4925) );
  INV_X1 U6444 ( .A(n4926), .ZN(n4927) );
  NAND2_X1 U6445 ( .A1(n4927), .A2(SI_14_), .ZN(n4928) );
  MUX2_X1 U6446 ( .A(n6809), .B(n4929), .S(n4278), .Z(n4931) );
  NAND2_X1 U6447 ( .A1(n4931), .A2(n4930), .ZN(n4935) );
  INV_X1 U6448 ( .A(n4931), .ZN(n4932) );
  NAND2_X1 U6449 ( .A1(n4932), .A2(SI_15_), .ZN(n4933) );
  NAND2_X1 U6450 ( .A1(n4935), .A2(n4933), .ZN(n5382) );
  INV_X1 U6451 ( .A(n5382), .ZN(n4934) );
  MUX2_X1 U6452 ( .A(n4937), .B(n4936), .S(n4283), .Z(n4939) );
  NAND2_X1 U6453 ( .A1(n4939), .A2(n4938), .ZN(n4942) );
  INV_X1 U6454 ( .A(n4939), .ZN(n4940) );
  NAND2_X1 U6455 ( .A1(n4940), .A2(SI_16_), .ZN(n4941) );
  NAND2_X1 U6456 ( .A1(n4943), .A2(n4942), .ZN(n5053) );
  INV_X1 U6457 ( .A(n5053), .ZN(n4945) );
  MUX2_X1 U6458 ( .A(n7038), .B(n4944), .S(n4278), .Z(n4946) );
  XNOR2_X1 U6459 ( .A(n4946), .B(SI_17_), .ZN(n5052) );
  NAND2_X1 U6460 ( .A1(n4945), .A2(n5052), .ZN(n4949) );
  INV_X1 U6461 ( .A(n4946), .ZN(n4947) );
  NAND2_X1 U6462 ( .A1(n4947), .A2(SI_17_), .ZN(n4948) );
  MUX2_X1 U6463 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n4283), .Z(n4951) );
  XNOR2_X1 U6464 ( .A(n4951), .B(SI_18_), .ZN(n5435) );
  INV_X1 U6465 ( .A(n5435), .ZN(n4950) );
  MUX2_X1 U6466 ( .A(n4952), .B(n7230), .S(n4283), .Z(n4954) );
  NAND2_X1 U6467 ( .A1(n4954), .A2(n4953), .ZN(n4957) );
  INV_X1 U6468 ( .A(n4954), .ZN(n4955) );
  NAND2_X1 U6469 ( .A1(n4955), .A2(SI_19_), .ZN(n4956) );
  NAND2_X1 U6470 ( .A1(n4957), .A2(n4956), .ZN(n5452) );
  MUX2_X1 U6471 ( .A(n7497), .B(n8386), .S(n4283), .Z(n4958) );
  NAND2_X1 U6472 ( .A1(n4958), .A2(n7387), .ZN(n4961) );
  INV_X1 U6473 ( .A(n4958), .ZN(n4959) );
  NAND2_X1 U6474 ( .A1(n4959), .A2(SI_20_), .ZN(n4960) );
  NAND2_X1 U6475 ( .A1(n5471), .A2(n5470), .ZN(n4962) );
  MUX2_X1 U6476 ( .A(n7511), .B(n7500), .S(n4278), .Z(n4963) );
  XNOR2_X1 U6477 ( .A(n4963), .B(SI_21_), .ZN(n5492) );
  INV_X1 U6478 ( .A(n5492), .ZN(n4966) );
  INV_X1 U6479 ( .A(n4963), .ZN(n4964) );
  NAND2_X1 U6480 ( .A1(n4964), .A2(SI_21_), .ZN(n4965) );
  MUX2_X1 U6481 ( .A(n8058), .B(n7649), .S(n4283), .Z(n4968) );
  INV_X1 U6482 ( .A(SI_22_), .ZN(n4967) );
  NAND2_X1 U6483 ( .A1(n4968), .A2(n4967), .ZN(n4971) );
  INV_X1 U6484 ( .A(n4968), .ZN(n4969) );
  NAND2_X1 U6485 ( .A1(n4969), .A2(SI_22_), .ZN(n4970) );
  NAND2_X1 U6486 ( .A1(n4971), .A2(n4970), .ZN(n5510) );
  MUX2_X1 U6487 ( .A(n7771), .B(n7757), .S(n4278), .Z(n4972) );
  NAND2_X1 U6488 ( .A1(n4972), .A2(n7462), .ZN(n5530) );
  INV_X1 U6489 ( .A(n4972), .ZN(n4973) );
  NAND2_X1 U6490 ( .A1(n4973), .A2(SI_23_), .ZN(n4974) );
  XNOR2_X1 U6491 ( .A(n5529), .B(n5528), .ZN(n7769) );
  NOR2_X1 U6492 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n4979) );
  NOR2_X1 U6493 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n4978) );
  NAND2_X1 U6494 ( .A1(n5386), .A2(n4982), .ZN(n4983) );
  INV_X1 U6495 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n4985) );
  NOR2_X1 U6496 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n4988) );
  NOR2_X1 U6497 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n4987) );
  NOR2_X1 U6498 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n4986) );
  NAND2_X1 U6499 ( .A1(n5001), .A2(n4991), .ZN(n5028) );
  NAND2_X1 U6500 ( .A1(n5028), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4992) );
  NAND2_X1 U6501 ( .A1(n5000), .A2(n4992), .ZN(n4995) );
  INV_X1 U6502 ( .A(n4995), .ZN(n4993) );
  NAND2_X1 U6503 ( .A1(n4993), .A2(n4855), .ZN(n4994) );
  NAND2_X1 U6504 ( .A1(n7769), .A2(n6416), .ZN(n4997) );
  NAND2_X1 U6505 ( .A1(n4287), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n4996) );
  NAND2_X1 U6506 ( .A1(n4999), .A2(n5003), .ZN(n4998) );
  NAND2_X1 U6507 ( .A1(n5000), .A2(n5001), .ZN(n5010) );
  OR2_X1 U6508 ( .A1(n5000), .A2(n5001), .ZN(n5002) );
  NAND2_X1 U6509 ( .A1(n5010), .A2(n5002), .ZN(n7941) );
  NOR2_X1 U6510 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n5005) );
  NOR2_X1 U6511 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n5004) );
  NAND2_X1 U6512 ( .A1(n5027), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5009) );
  XNOR2_X1 U6513 ( .A(n5009), .B(P1_IR_REG_24__SCAN_IN), .ZN(n5634) );
  NAND2_X1 U6514 ( .A1(n5010), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5011) );
  INV_X1 U6515 ( .A(n6568), .ZN(n5013) );
  NAND3_X1 U6516 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n5188) );
  INV_X1 U6517 ( .A(n5188), .ZN(n5014) );
  NAND2_X1 U6518 ( .A1(n5014), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5217) );
  INV_X1 U6519 ( .A(n5217), .ZN(n5015) );
  NAND2_X1 U6520 ( .A1(n5015), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5261) );
  INV_X1 U6521 ( .A(n5261), .ZN(n5016) );
  NAND2_X1 U6522 ( .A1(n5016), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5263) );
  INV_X1 U6523 ( .A(n5326), .ZN(n5018) );
  INV_X1 U6524 ( .A(n5456), .ZN(n5022) );
  INV_X1 U6525 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n5496) );
  INV_X1 U6526 ( .A(n5516), .ZN(n5024) );
  INV_X1 U6527 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n5025) );
  NAND2_X1 U6528 ( .A1(n5516), .A2(n5025), .ZN(n5026) );
  NAND2_X1 U6529 ( .A1(n5535), .A2(n5026), .ZN(n9308) );
  INV_X1 U6530 ( .A(n5028), .ZN(n5031) );
  NOR2_X1 U6531 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), .ZN(
        n5030) );
  NAND2_X1 U6533 ( .A1(n5032), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5034) );
  OR2_X1 U6534 ( .A1(n9308), .A2(n5166), .ZN(n5043) );
  INV_X1 U6535 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n9309) );
  NAND2_X1 U6536 ( .A1(n4289), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n5040) );
  NAND2_X1 U6537 ( .A1(n4290), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5039) );
  OAI211_X1 U6538 ( .C1(n5111), .C2(n9309), .A(n5040), .B(n5039), .ZN(n5041)
         );
  INV_X1 U6539 ( .A(n5041), .ZN(n5042) );
  AND2_X4 U6540 ( .A1(n5064), .A2(n6568), .ZN(n5700) );
  INV_X1 U6541 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5044) );
  NAND2_X1 U6542 ( .A1(n5045), .A2(n5044), .ZN(n5046) );
  NAND2_X1 U6543 ( .A1(n5049), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5050) );
  NAND2_X1 U6544 ( .A1(n5631), .A2(n5663), .ZN(n5051) );
  OAI22_X1 U6545 ( .A1(n9307), .A2(n5093), .B1(n9179), .B2(n5451), .ZN(n9056)
         );
  XNOR2_X1 U6546 ( .A(n5053), .B(n5052), .ZN(n7009) );
  NAND2_X1 U6547 ( .A1(n7009), .A2(n6416), .ZN(n5056) );
  NAND2_X1 U6548 ( .A1(n5054), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5438) );
  XNOR2_X1 U6549 ( .A(n5438), .B(P1_IR_REG_17__SCAN_IN), .ZN(n8288) );
  AOI22_X1 U6550 ( .A1(n4287), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n6579), .B2(
        n8288), .ZN(n5055) );
  NAND2_X1 U6551 ( .A1(n5416), .A2(n5057), .ZN(n5058) );
  AND2_X1 U6552 ( .A1(n5444), .A2(n5058), .ZN(n9087) );
  NAND2_X1 U6553 ( .A1(n9087), .A2(n5087), .ZN(n5063) );
  NAND2_X1 U6554 ( .A1(n4289), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n5060) );
  NAND2_X1 U6555 ( .A1(n4290), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5059) );
  AND2_X1 U6556 ( .A1(n5060), .A2(n5059), .ZN(n5062) );
  INV_X4 U6557 ( .A(n5111), .ZN(n5586) );
  NAND2_X1 U6558 ( .A1(n5586), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5061) );
  OAI22_X1 U6559 ( .A1(n9084), .A2(n5093), .B1(n8037), .B2(n5451), .ZN(n5431)
         );
  INV_X1 U6560 ( .A(n5431), .ZN(n5434) );
  OAI22_X1 U6561 ( .A1(n9084), .A2(n5570), .B1(n8037), .B2(n5093), .ZN(n5065)
         );
  NAND2_X1 U6562 ( .A1(n5655), .A2(n9298), .ZN(n7017) );
  XNOR2_X1 U6563 ( .A(n5065), .B(n7124), .ZN(n5432) );
  INV_X1 U6564 ( .A(n5432), .ZN(n5433) );
  XNOR2_X1 U6565 ( .A(n5067), .B(n5066), .ZN(n6637) );
  OR2_X1 U6566 ( .A1(n5108), .A2(n6637), .ZN(n5072) );
  NAND2_X1 U6567 ( .A1(n5069), .A2(P1_IR_REG_2__SCAN_IN), .ZN(n5070) );
  AND2_X1 U6568 ( .A1(n5070), .A2(n5130), .ZN(n6855) );
  NAND2_X1 U6569 ( .A1(n6579), .A2(n6855), .ZN(n5071) );
  NAND2_X1 U6570 ( .A1(n5087), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5078) );
  NAND2_X1 U6571 ( .A1(n4288), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5077) );
  INV_X1 U6572 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n5074) );
  OR2_X1 U6573 ( .A1(n5111), .A2(n5074), .ZN(n5076) );
  NAND2_X1 U6574 ( .A1(n5446), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5075) );
  NAND4_X1 U6575 ( .A1(n5078), .A2(n5077), .A3(n5076), .A4(n5075), .ZN(n9161)
         );
  OAI22_X1 U6576 ( .A1(n7255), .A2(n5570), .B1(n5093), .B2(n6307), .ZN(n5079)
         );
  XNOR2_X1 U6577 ( .A(n5079), .B(n5247), .ZN(n5082) );
  OR2_X1 U6578 ( .A1(n4285), .A2(n6307), .ZN(n5081) );
  NAND2_X1 U6579 ( .A1(n9815), .A2(n5695), .ZN(n5080) );
  AND2_X1 U6580 ( .A1(n5081), .A2(n5080), .ZN(n5083) );
  NAND2_X1 U6581 ( .A1(n5082), .A2(n5083), .ZN(n5125) );
  INV_X1 U6582 ( .A(n5082), .ZN(n5085) );
  INV_X1 U6583 ( .A(n5083), .ZN(n5084) );
  NAND2_X1 U6584 ( .A1(n5085), .A2(n5084), .ZN(n5086) );
  NAND2_X1 U6585 ( .A1(n5446), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5091) );
  NAND2_X1 U6586 ( .A1(n5087), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5090) );
  NAND2_X1 U6587 ( .A1(n4288), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5088) );
  NAND4_X2 U6588 ( .A1(n5091), .A2(n5090), .A3(n5089), .A4(n5088), .ZN(n7011)
         );
  INV_X1 U6589 ( .A(n7011), .ZN(n5092) );
  NAND2_X1 U6590 ( .A1(n4278), .A2(SI_0_), .ZN(n5095) );
  INV_X1 U6591 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5094) );
  NAND2_X1 U6592 ( .A1(n5095), .A2(n5094), .ZN(n5097) );
  AND2_X1 U6593 ( .A1(n5097), .A2(n5096), .ZN(n6617) );
  MUX2_X1 U6594 ( .A(P1_IR_REG_0__SCAN_IN), .B(n6617), .S(n5110), .Z(n7176) );
  NAND2_X1 U6595 ( .A1(n5700), .A2(n7176), .ZN(n5099) );
  INV_X1 U6596 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n5098) );
  OAI211_X1 U6597 ( .C1(n5092), .C2(n5093), .A(n5099), .B(n4857), .ZN(n6695)
         );
  INV_X1 U6598 ( .A(n6695), .ZN(n5100) );
  NAND2_X1 U6599 ( .A1(n5100), .A2(n7124), .ZN(n5106) );
  INV_X1 U6600 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n5101) );
  NOR2_X1 U6601 ( .A1(n6568), .A2(n5101), .ZN(n5102) );
  AOI21_X1 U6602 ( .B1(n4276), .B2(n7176), .A(n5102), .ZN(n5105) );
  INV_X1 U6603 ( .A(n5171), .ZN(n5103) );
  NAND2_X1 U6604 ( .A1(n5103), .A2(n7011), .ZN(n5104) );
  AND2_X1 U6605 ( .A1(n5105), .A2(n5104), .ZN(n6696) );
  NAND2_X1 U6606 ( .A1(n6696), .A2(n6695), .ZN(n6694) );
  NAND2_X1 U6607 ( .A1(n5106), .A2(n6694), .ZN(n6728) );
  INV_X1 U6608 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6621) );
  NAND2_X1 U6609 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5109) );
  XNOR2_X1 U6610 ( .A(n5109), .B(P1_IR_REG_1__SCAN_IN), .ZN(n6864) );
  NAND2_X1 U6611 ( .A1(n5700), .A2(n6305), .ZN(n5117) );
  INV_X1 U6612 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n7032) );
  NAND2_X1 U6613 ( .A1(n4289), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5115) );
  NAND2_X1 U6614 ( .A1(n5586), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5114) );
  INV_X1 U6615 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n5112) );
  OR2_X1 U6616 ( .A1(n5241), .A2(n5112), .ZN(n5113) );
  OR2_X1 U6617 ( .A1(n5171), .A2(n6693), .ZN(n5119) );
  INV_X2 U6618 ( .A(n5093), .ZN(n5621) );
  NAND2_X1 U6619 ( .A1(n5621), .A2(n7034), .ZN(n5118) );
  NAND2_X1 U6620 ( .A1(n5119), .A2(n5118), .ZN(n6727) );
  NAND2_X1 U6621 ( .A1(n5120), .A2(n6727), .ZN(n5124) );
  INV_X1 U6622 ( .A(n6728), .ZN(n5122) );
  INV_X1 U6623 ( .A(n6730), .ZN(n5121) );
  NAND2_X1 U6624 ( .A1(n5122), .A2(n5121), .ZN(n5123) );
  AND2_X2 U6625 ( .A1(n5124), .A2(n5123), .ZN(n6752) );
  NAND2_X1 U6626 ( .A1(n6753), .A2(n6752), .ZN(n6751) );
  NAND2_X1 U6627 ( .A1(n6751), .A2(n5125), .ZN(n6811) );
  NAND2_X1 U6628 ( .A1(n4287), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n5134) );
  NAND2_X1 U6629 ( .A1(n5127), .A2(n5126), .ZN(n5128) );
  XNOR2_X1 U6630 ( .A(n5129), .B(n5128), .ZN(n6630) );
  NAND2_X1 U6631 ( .A1(n5130), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5131) );
  XNOR2_X1 U6632 ( .A(n5131), .B(P1_IR_REG_3__SCAN_IN), .ZN(n6622) );
  NAND2_X1 U6633 ( .A1(n6579), .A2(n6622), .ZN(n5132) );
  OR2_X1 U6634 ( .A1(n5166), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n5139) );
  NAND2_X1 U6635 ( .A1(n5586), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5136) );
  NAND2_X1 U6636 ( .A1(n5446), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5135) );
  OAI22_X1 U6637 ( .A1(n9823), .A2(n5570), .B1(n5093), .B2(n9783), .ZN(n5140)
         );
  XNOR2_X1 U6638 ( .A(n5140), .B(n4286), .ZN(n5160) );
  OR2_X1 U6639 ( .A1(n5171), .A2(n9783), .ZN(n5142) );
  INV_X2 U6640 ( .A(n5093), .ZN(n5695) );
  NAND2_X1 U6641 ( .A1(n7294), .A2(n5695), .ZN(n5141) );
  NAND2_X1 U6642 ( .A1(n5142), .A2(n5141), .ZN(n5158) );
  XNOR2_X1 U6643 ( .A(n5160), .B(n5158), .ZN(n6812) );
  NAND2_X1 U6644 ( .A1(n6811), .A2(n6812), .ZN(n6810) );
  NAND2_X1 U6645 ( .A1(n4287), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n5150) );
  OR2_X1 U6646 ( .A1(n5108), .A2(n6632), .ZN(n5149) );
  NAND2_X1 U6647 ( .A1(n5144), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5145) );
  MUX2_X1 U6648 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5145), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n5147) );
  AND2_X1 U6649 ( .A1(n5147), .A2(n5146), .ZN(n6602) );
  NAND2_X1 U6650 ( .A1(n6579), .A2(n6602), .ZN(n5148) );
  XNOR2_X1 U6651 ( .A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n9793) );
  OR2_X1 U6652 ( .A1(n5166), .A2(n9793), .ZN(n5154) );
  NAND2_X1 U6653 ( .A1(n4289), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5153) );
  NAND2_X1 U6654 ( .A1(n4290), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5152) );
  NAND2_X1 U6655 ( .A1(n5586), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5151) );
  NAND4_X1 U6656 ( .A1(n5154), .A2(n5153), .A3(n5152), .A4(n5151), .ZN(n9159)
         );
  OAI22_X1 U6657 ( .A1(n9829), .A2(n5570), .B1(n5093), .B2(n9767), .ZN(n5155)
         );
  XNOR2_X1 U6658 ( .A(n5155), .B(n7124), .ZN(n5164) );
  OR2_X1 U6659 ( .A1(n5171), .A2(n9767), .ZN(n5157) );
  NAND2_X1 U6660 ( .A1(n7116), .A2(n5621), .ZN(n5156) );
  AND2_X1 U6661 ( .A1(n5157), .A2(n5156), .ZN(n5162) );
  XNOR2_X1 U6662 ( .A(n5164), .B(n5162), .ZN(n6887) );
  INV_X1 U6663 ( .A(n5158), .ZN(n5159) );
  NAND2_X1 U6664 ( .A1(n5160), .A2(n5159), .ZN(n6885) );
  AND2_X1 U6665 ( .A1(n6887), .A2(n6885), .ZN(n5161) );
  INV_X1 U6666 ( .A(n5162), .ZN(n5163) );
  NAND2_X1 U6667 ( .A1(n5164), .A2(n5163), .ZN(n7218) );
  INV_X1 U6668 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n7281) );
  NAND2_X1 U6669 ( .A1(n5188), .A2(n7281), .ZN(n5165) );
  NAND2_X1 U6670 ( .A1(n5217), .A2(n5165), .ZN(n9743) );
  OR2_X1 U6671 ( .A1(n5166), .A2(n9743), .ZN(n5170) );
  NAND2_X1 U6672 ( .A1(n4288), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5169) );
  NAND2_X1 U6673 ( .A1(n5586), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5168) );
  NAND2_X1 U6674 ( .A1(n5446), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5167) );
  OR2_X1 U6675 ( .A1(n4285), .A2(n5181), .ZN(n5180) );
  NAND2_X1 U6676 ( .A1(n5213), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n5178) );
  XNOR2_X1 U6677 ( .A(n5172), .B(n5173), .ZN(n6641) );
  OR2_X1 U6678 ( .A1(n5108), .A2(n6641), .ZN(n5177) );
  INV_X1 U6679 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9493) );
  OR2_X1 U6680 ( .A1(n5174), .A2(n9493), .ZN(n5175) );
  XNOR2_X1 U6681 ( .A(n5175), .B(P1_IR_REG_6__SCAN_IN), .ZN(n6640) );
  NAND2_X1 U6682 ( .A1(n6579), .A2(n6640), .ZN(n5176) );
  AND3_X2 U6683 ( .A1(n5178), .A2(n5177), .A3(n5176), .ZN(n9841) );
  INV_X1 U6684 ( .A(n9841), .ZN(n7284) );
  NAND2_X1 U6685 ( .A1(n7284), .A2(n5621), .ZN(n5179) );
  AND2_X1 U6686 ( .A1(n5180), .A2(n5179), .ZN(n5184) );
  OAI22_X1 U6687 ( .A1(n9841), .A2(n5570), .B1(n5093), .B2(n5181), .ZN(n5182)
         );
  XNOR2_X1 U6688 ( .A(n5182), .B(n5247), .ZN(n5183) );
  NAND2_X1 U6689 ( .A1(n5183), .A2(n5184), .ZN(n5207) );
  OAI21_X1 U6690 ( .B1(n5184), .B2(n5183), .A(n5207), .ZN(n7274) );
  INV_X1 U6691 ( .A(n7274), .ZN(n5201) );
  NAND2_X1 U6692 ( .A1(n4289), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5191) );
  INV_X1 U6693 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5186) );
  NAND2_X1 U6694 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n5185) );
  NAND2_X1 U6695 ( .A1(n5186), .A2(n5185), .ZN(n5187) );
  NAND2_X1 U6696 ( .A1(n5188), .A2(n5187), .ZN(n7225) );
  OR2_X1 U6697 ( .A1(n5166), .A2(n7225), .ZN(n5190) );
  NAND2_X1 U6699 ( .A1(n4287), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n5197) );
  XNOR2_X1 U6700 ( .A(n5192), .B(n5193), .ZN(n6627) );
  OR2_X1 U6701 ( .A1(n5108), .A2(n6627), .ZN(n5196) );
  NAND2_X1 U6702 ( .A1(n5146), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5194) );
  XNOR2_X1 U6703 ( .A(n5194), .B(P1_IR_REG_5__SCAN_IN), .ZN(n6625) );
  NAND2_X1 U6704 ( .A1(n6579), .A2(n6625), .ZN(n5195) );
  OR2_X1 U6705 ( .A1(n5171), .A2(n9782), .ZN(n5200) );
  INV_X1 U6706 ( .A(n9836), .ZN(n9752) );
  NAND2_X1 U6707 ( .A1(n9752), .A2(n5621), .ZN(n5199) );
  AND2_X1 U6708 ( .A1(n5200), .A2(n5199), .ZN(n7217) );
  INV_X1 U6709 ( .A(n5206), .ZN(n5202) );
  AND2_X1 U6710 ( .A1(n7218), .A2(n5202), .ZN(n5203) );
  NAND2_X1 U6711 ( .A1(n5204), .A2(n7217), .ZN(n5205) );
  OR2_X1 U6712 ( .A1(n5206), .A2(n5205), .ZN(n7278) );
  AND2_X1 U6713 ( .A1(n5207), .A2(n7278), .ZN(n5208) );
  NAND2_X1 U6714 ( .A1(n5174), .A2(n5211), .ZN(n5233) );
  NAND2_X1 U6715 ( .A1(n5233), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5212) );
  XNOR2_X1 U6716 ( .A(n5212), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6647) );
  AOI22_X1 U6717 ( .A1(n4287), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n6579), .B2(
        n6647), .ZN(n5214) );
  NAND2_X1 U6718 ( .A1(n5215), .A2(n5214), .ZN(n7106) );
  INV_X1 U6719 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5216) );
  NAND2_X1 U6720 ( .A1(n5217), .A2(n5216), .ZN(n5218) );
  NAND2_X1 U6721 ( .A1(n5261), .A2(n5218), .ZN(n8312) );
  OR2_X1 U6722 ( .A1(n5166), .A2(n8312), .ZN(n5222) );
  NAND2_X1 U6723 ( .A1(n4289), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5221) );
  NAND2_X1 U6724 ( .A1(n5586), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5220) );
  NAND2_X1 U6725 ( .A1(n4290), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5219) );
  NAND4_X1 U6726 ( .A1(n5222), .A2(n5221), .A3(n5220), .A4(n5219), .ZN(n9735)
         );
  OAI22_X1 U6727 ( .A1(n9849), .A2(n5570), .B1(n7315), .B2(n5093), .ZN(n5223)
         );
  XNOR2_X1 U6728 ( .A(n5223), .B(n5247), .ZN(n5225) );
  OR2_X1 U6729 ( .A1(n5171), .A2(n7315), .ZN(n5224) );
  OAI21_X1 U6730 ( .B1(n9849), .B2(n5093), .A(n5224), .ZN(n5226) );
  XNOR2_X1 U6731 ( .A(n5225), .B(n5226), .ZN(n8310) );
  INV_X1 U6732 ( .A(n5225), .ZN(n5227) );
  OR2_X1 U6733 ( .A1(n5227), .A2(n5226), .ZN(n7304) );
  NAND2_X1 U6734 ( .A1(n5231), .A2(n5230), .ZN(n5232) );
  NOR2_X1 U6735 ( .A1(n5255), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n5277) );
  OR2_X1 U6736 ( .A1(n5277), .A2(n9493), .ZN(n5234) );
  XNOR2_X1 U6737 ( .A(n5234), .B(P1_IR_REG_9__SCAN_IN), .ZN(n6775) );
  AOI22_X1 U6738 ( .A1(n4287), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n6579), .B2(
        n6775), .ZN(n5235) );
  NAND2_X1 U6739 ( .A1(n5586), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5246) );
  INV_X1 U6740 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n5238) );
  OR2_X1 U6741 ( .A1(n5237), .A2(n5238), .ZN(n5245) );
  NAND2_X1 U6742 ( .A1(n5263), .A2(n5239), .ZN(n5240) );
  NAND2_X1 U6743 ( .A1(n5281), .A2(n5240), .ZN(n7486) );
  OR2_X1 U6744 ( .A1(n5166), .A2(n7486), .ZN(n5244) );
  INV_X1 U6745 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n5242) );
  OR2_X1 U6746 ( .A1(n5241), .A2(n5242), .ZN(n5243) );
  OAI22_X1 U6747 ( .A1(n9864), .A2(n5570), .B1(n7207), .B2(n5093), .ZN(n5248)
         );
  XNOR2_X1 U6748 ( .A(n5248), .B(n4286), .ZN(n5292) );
  OAI22_X1 U6749 ( .A1(n9864), .A2(n5093), .B1(n7207), .B2(n5451), .ZN(n5291)
         );
  INV_X1 U6750 ( .A(n5291), .ZN(n5249) );
  NAND2_X1 U6751 ( .A1(n5292), .A2(n5249), .ZN(n5251) );
  AND2_X1 U6752 ( .A1(n7304), .A2(n5251), .ZN(n5250) );
  INV_X1 U6753 ( .A(n5251), .ZN(n5293) );
  INV_X1 U6754 ( .A(n5252), .ZN(n5253) );
  XNOR2_X1 U6755 ( .A(n5254), .B(n5253), .ZN(n5863) );
  INV_X1 U6756 ( .A(n5277), .ZN(n5258) );
  NAND2_X1 U6757 ( .A1(n5255), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5256) );
  MUX2_X1 U6758 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5256), .S(
        P1_IR_REG_8__SCAN_IN), .Z(n5257) );
  NAND2_X1 U6759 ( .A1(n6314), .A2(n5621), .ZN(n5270) );
  NAND2_X1 U6760 ( .A1(n4288), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5268) );
  INV_X1 U6761 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n6592) );
  OR2_X1 U6762 ( .A1(n5111), .A2(n6592), .ZN(n5267) );
  INV_X1 U6763 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6744) );
  NAND2_X1 U6764 ( .A1(n5261), .A2(n6744), .ZN(n5262) );
  NAND2_X1 U6765 ( .A1(n5263), .A2(n5262), .ZN(n7186) );
  OR2_X1 U6766 ( .A1(n5166), .A2(n7186), .ZN(n5266) );
  INV_X1 U6767 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n5264) );
  OR2_X1 U6768 ( .A1(n5241), .A2(n5264), .ZN(n5265) );
  OR2_X1 U6769 ( .A1(n5451), .A2(n8315), .ZN(n5269) );
  AND2_X1 U6770 ( .A1(n5270), .A2(n5269), .ZN(n7305) );
  NAND2_X1 U6771 ( .A1(n6314), .A2(n5700), .ZN(n5272) );
  OR2_X1 U6772 ( .A1(n8315), .A2(n5093), .ZN(n5271) );
  NAND2_X1 U6773 ( .A1(n5272), .A2(n5271), .ZN(n5273) );
  XNOR2_X1 U6774 ( .A(n5273), .B(n4286), .ZN(n7307) );
  AND2_X1 U6775 ( .A1(n8310), .A2(n7307), .ZN(n5274) );
  INV_X1 U6776 ( .A(n7304), .ZN(n5275) );
  NAND2_X1 U6777 ( .A1(n6657), .A2(n6416), .ZN(n5280) );
  INV_X1 U6778 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n5276) );
  NAND2_X1 U6779 ( .A1(n5277), .A2(n5276), .ZN(n5299) );
  NAND2_X1 U6780 ( .A1(n5299), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5278) );
  XNOR2_X1 U6781 ( .A(n5278), .B(P1_IR_REG_10__SCAN_IN), .ZN(n6776) );
  AOI22_X1 U6782 ( .A1(n4287), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6579), .B2(
        n6776), .ZN(n5279) );
  NAND2_X1 U6783 ( .A1(n5280), .A2(n5279), .ZN(n7503) );
  NAND2_X1 U6784 ( .A1(n7503), .A2(n5700), .ZN(n5288) );
  NAND2_X1 U6785 ( .A1(n5281), .A2(n7268), .ZN(n5282) );
  NAND2_X1 U6786 ( .A1(n5304), .A2(n5282), .ZN(n7211) );
  OR2_X1 U6787 ( .A1(n5166), .A2(n7211), .ZN(n5286) );
  NAND2_X1 U6788 ( .A1(n5446), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5285) );
  NAND2_X1 U6789 ( .A1(n4288), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5284) );
  NAND2_X1 U6790 ( .A1(n5586), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5283) );
  NAND4_X1 U6791 ( .A1(n5286), .A2(n5285), .A3(n5284), .A4(n5283), .ZN(n9155)
         );
  INV_X1 U6792 ( .A(n9155), .ZN(n7490) );
  OR2_X1 U6793 ( .A1(n7490), .A2(n5093), .ZN(n5287) );
  NAND2_X1 U6794 ( .A1(n5288), .A2(n5287), .ZN(n5289) );
  XNOR2_X1 U6795 ( .A(n5289), .B(n5247), .ZN(n5296) );
  NOR2_X1 U6796 ( .A1(n5451), .A2(n7490), .ZN(n5290) );
  AOI21_X1 U6797 ( .B1(n7503), .B2(n5695), .A(n5290), .ZN(n5295) );
  OR2_X1 U6798 ( .A1(n5296), .A2(n5295), .ZN(n7264) );
  XNOR2_X1 U6799 ( .A(n5292), .B(n5291), .ZN(n7484) );
  OR2_X1 U6800 ( .A1(n5293), .A2(n7484), .ZN(n7261) );
  AND2_X1 U6801 ( .A1(n7264), .A2(n7261), .ZN(n5294) );
  NAND2_X1 U6802 ( .A1(n5296), .A2(n5295), .ZN(n7263) );
  XNOR2_X1 U6803 ( .A(n5297), .B(n5298), .ZN(n6666) );
  NAND2_X1 U6804 ( .A1(n6666), .A2(n6416), .ZN(n5302) );
  OAI21_X1 U6805 ( .B1(n5299), .B2(P1_IR_REG_10__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5300) );
  XNOR2_X1 U6806 ( .A(n5300), .B(P1_IR_REG_11__SCAN_IN), .ZN(n8334) );
  AOI22_X1 U6807 ( .A1(n5213), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n6579), .B2(
        n8334), .ZN(n5301) );
  NAND2_X1 U6808 ( .A1(n5302), .A2(n5301), .ZN(n9470) );
  NAND2_X1 U6809 ( .A1(n9470), .A2(n5700), .ZN(n5311) );
  INV_X1 U6810 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5303) );
  NAND2_X1 U6811 ( .A1(n5304), .A2(n5303), .ZN(n5305) );
  NAND2_X1 U6812 ( .A1(n5326), .A2(n5305), .ZN(n7159) );
  OR2_X1 U6813 ( .A1(n5166), .A2(n7159), .ZN(n5309) );
  NAND2_X1 U6814 ( .A1(n4290), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5308) );
  NAND2_X1 U6815 ( .A1(n4289), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5307) );
  NAND2_X1 U6816 ( .A1(n5586), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5306) );
  NAND4_X1 U6817 ( .A1(n5309), .A2(n5308), .A3(n5307), .A4(n5306), .ZN(n9559)
         );
  INV_X1 U6818 ( .A(n9559), .ZN(n7655) );
  OR2_X1 U6819 ( .A1(n7655), .A2(n5093), .ZN(n5310) );
  NAND2_X1 U6820 ( .A1(n5311), .A2(n5310), .ZN(n5312) );
  XNOR2_X1 U6821 ( .A(n5312), .B(n4286), .ZN(n5315) );
  NOR2_X1 U6822 ( .A1(n5451), .A2(n7655), .ZN(n5313) );
  AOI21_X1 U6823 ( .B1(n9470), .B2(n5621), .A(n5313), .ZN(n5314) );
  XNOR2_X1 U6824 ( .A(n5315), .B(n5314), .ZN(n7643) );
  OR2_X1 U6825 ( .A1(n5315), .A2(n5314), .ZN(n5316) );
  XNOR2_X1 U6826 ( .A(n5318), .B(n5317), .ZN(n6674) );
  NAND2_X1 U6827 ( .A1(n6674), .A2(n6416), .ZN(n5324) );
  NOR2_X1 U6828 ( .A1(n5319), .A2(n9493), .ZN(n5320) );
  MUX2_X1 U6829 ( .A(n9493), .B(n5320), .S(P1_IR_REG_12__SCAN_IN), .Z(n5322)
         );
  OR2_X1 U6830 ( .A1(n5322), .A2(n5321), .ZN(n8291) );
  INV_X1 U6831 ( .A(n8291), .ZN(n8271) );
  AOI22_X1 U6832 ( .A1(n4287), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6579), .B2(
        n8271), .ZN(n5323) );
  NAND2_X1 U6833 ( .A1(n5324), .A2(n5323), .ZN(n9571) );
  NAND2_X1 U6834 ( .A1(n9571), .A2(n5700), .ZN(n5334) );
  NAND2_X1 U6835 ( .A1(n4290), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5332) );
  INV_X1 U6836 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5325) );
  NAND2_X1 U6837 ( .A1(n5326), .A2(n5325), .ZN(n5327) );
  NAND2_X1 U6838 ( .A1(n5349), .A2(n5327), .ZN(n9566) );
  OR2_X1 U6839 ( .A1(n5166), .A2(n9566), .ZN(n5331) );
  INV_X1 U6840 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n5328) );
  OR2_X1 U6841 ( .A1(n5237), .A2(n5328), .ZN(n5330) );
  INV_X1 U6842 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n6771) );
  OR2_X1 U6843 ( .A1(n5111), .A2(n6771), .ZN(n5329) );
  OR2_X1 U6844 ( .A1(n7674), .A2(n5093), .ZN(n5333) );
  NAND2_X1 U6845 ( .A1(n5334), .A2(n5333), .ZN(n5335) );
  XNOR2_X1 U6846 ( .A(n5335), .B(n4286), .ZN(n5340) );
  NOR2_X1 U6847 ( .A1(n5451), .A2(n7674), .ZN(n5336) );
  AOI21_X1 U6848 ( .B1(n9571), .B2(n5695), .A(n5336), .ZN(n5339) );
  XNOR2_X1 U6849 ( .A(n5340), .B(n5339), .ZN(n7653) );
  INV_X1 U6850 ( .A(n7653), .ZN(n5337) );
  NAND2_X1 U6851 ( .A1(n5340), .A2(n5339), .ZN(n5341) );
  XNOR2_X1 U6852 ( .A(n5343), .B(n5342), .ZN(n6679) );
  NAND2_X1 U6853 ( .A1(n6679), .A2(n6416), .ZN(n5347) );
  NAND2_X1 U6854 ( .A1(n5344), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5345) );
  XNOR2_X1 U6855 ( .A(n5345), .B(P1_IR_REG_13__SCAN_IN), .ZN(n9645) );
  AOI22_X1 U6856 ( .A1(n4287), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n6579), .B2(
        n9645), .ZN(n5346) );
  NAND2_X1 U6857 ( .A1(n7823), .A2(n5700), .ZN(n5356) );
  NAND2_X1 U6858 ( .A1(n5349), .A2(n5348), .ZN(n5350) );
  NAND2_X1 U6859 ( .A1(n5370), .A2(n5350), .ZN(n7677) );
  OR2_X1 U6860 ( .A1(n5166), .A2(n7677), .ZN(n5354) );
  NAND2_X1 U6861 ( .A1(n4288), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5353) );
  NAND2_X1 U6862 ( .A1(n5446), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5352) );
  NAND2_X1 U6863 ( .A1(n5586), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5351) );
  NAND4_X1 U6864 ( .A1(n5354), .A2(n5353), .A3(n5352), .A4(n5351), .ZN(n9153)
         );
  OR2_X1 U6865 ( .A1(n9561), .A2(n5093), .ZN(n5355) );
  NAND2_X1 U6866 ( .A1(n5356), .A2(n5355), .ZN(n5357) );
  XNOR2_X1 U6867 ( .A(n5357), .B(n5247), .ZN(n7671) );
  NOR2_X1 U6868 ( .A1(n5451), .A2(n9561), .ZN(n5358) );
  AOI21_X1 U6869 ( .B1(n7823), .B2(n5695), .A(n5358), .ZN(n7670) );
  AND2_X1 U6870 ( .A1(n7671), .A2(n7670), .ZN(n5362) );
  INV_X1 U6871 ( .A(n7671), .ZN(n5360) );
  INV_X1 U6872 ( .A(n7670), .ZN(n5359) );
  NAND2_X1 U6873 ( .A1(n5360), .A2(n5359), .ZN(n5361) );
  XNOR2_X1 U6874 ( .A(n5364), .B(n5363), .ZN(n6683) );
  NAND2_X1 U6875 ( .A1(n6683), .A2(n6416), .ZN(n5369) );
  INV_X1 U6876 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5365) );
  NAND2_X1 U6877 ( .A1(n5321), .A2(n5365), .ZN(n5366) );
  NAND2_X1 U6878 ( .A1(n5366), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5387) );
  XNOR2_X1 U6879 ( .A(n5387), .B(n5386), .ZN(n9660) );
  INV_X1 U6880 ( .A(n9660), .ZN(n5367) );
  AOI22_X1 U6881 ( .A1(n5213), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n6579), .B2(
        n5367), .ZN(n5368) );
  NAND2_X1 U6882 ( .A1(n7877), .A2(n5700), .ZN(n5377) );
  INV_X1 U6883 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n7872) );
  NAND2_X1 U6884 ( .A1(n5370), .A2(n7872), .ZN(n5371) );
  NAND2_X1 U6885 ( .A1(n5393), .A2(n5371), .ZN(n7875) );
  OR2_X1 U6886 ( .A1(n5166), .A2(n7875), .ZN(n5375) );
  NAND2_X1 U6887 ( .A1(n5446), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5374) );
  NAND2_X1 U6888 ( .A1(n4289), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5373) );
  NAND2_X1 U6889 ( .A1(n5586), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5372) );
  NAND4_X1 U6890 ( .A1(n5375), .A2(n5374), .A3(n5373), .A4(n5372), .ZN(n9152)
         );
  INV_X1 U6891 ( .A(n9152), .ZN(n7963) );
  OR2_X1 U6892 ( .A1(n7963), .A2(n5093), .ZN(n5376) );
  NAND2_X1 U6893 ( .A1(n5377), .A2(n5376), .ZN(n5378) );
  XNOR2_X1 U6894 ( .A(n5378), .B(n7124), .ZN(n7869) );
  INV_X1 U6895 ( .A(n7869), .ZN(n5381) );
  NAND2_X1 U6896 ( .A1(n7877), .A2(n5621), .ZN(n5380) );
  OR2_X1 U6897 ( .A1(n5451), .A2(n7963), .ZN(n5379) );
  NAND2_X1 U6898 ( .A1(n5380), .A2(n5379), .ZN(n5402) );
  INV_X1 U6899 ( .A(n5402), .ZN(n7868) );
  NAND2_X1 U6900 ( .A1(n5381), .A2(n7868), .ZN(n5405) );
  NAND2_X1 U6901 ( .A1(n5383), .A2(n5382), .ZN(n5384) );
  NAND2_X1 U6902 ( .A1(n6749), .A2(n6416), .ZN(n5391) );
  NAND2_X1 U6903 ( .A1(n5387), .A2(n5386), .ZN(n5388) );
  NAND2_X1 U6904 ( .A1(n5388), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5389) );
  XNOR2_X1 U6905 ( .A(n5389), .B(P1_IR_REG_15__SCAN_IN), .ZN(n9674) );
  AOI22_X1 U6906 ( .A1(n4287), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n6579), .B2(
        n9674), .ZN(n5390) );
  NAND2_X1 U6907 ( .A1(n7912), .A2(n5700), .ZN(n5400) );
  NAND2_X1 U6908 ( .A1(n5393), .A2(n5392), .ZN(n5394) );
  NAND2_X1 U6909 ( .A1(n5414), .A2(n5394), .ZN(n7964) );
  OR2_X1 U6910 ( .A1(n5166), .A2(n7964), .ZN(n5398) );
  NAND2_X1 U6911 ( .A1(n4290), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5397) );
  NAND2_X1 U6912 ( .A1(n4289), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5396) );
  NAND2_X1 U6913 ( .A1(n5586), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5395) );
  NAND4_X1 U6914 ( .A1(n5398), .A2(n5397), .A3(n5396), .A4(n5395), .ZN(n9151)
         );
  OR2_X1 U6915 ( .A1(n7913), .A2(n5093), .ZN(n5399) );
  NAND2_X1 U6916 ( .A1(n5400), .A2(n5399), .ZN(n5401) );
  XNOR2_X1 U6917 ( .A(n5401), .B(n7124), .ZN(n5406) );
  AND2_X1 U6918 ( .A1(n7869), .A2(n5402), .ZN(n5404) );
  NOR2_X1 U6919 ( .A1(n5451), .A2(n7913), .ZN(n5403) );
  AOI21_X1 U6920 ( .B1(n7912), .B2(n5695), .A(n5403), .ZN(n7959) );
  XNOR2_X1 U6921 ( .A(n5407), .B(n5408), .ZN(n6881) );
  NAND2_X1 U6922 ( .A1(n6881), .A2(n6416), .ZN(n5412) );
  OR2_X1 U6923 ( .A1(n5409), .A2(n9493), .ZN(n5410) );
  XNOR2_X1 U6924 ( .A(n5410), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9687) );
  AOI22_X1 U6925 ( .A1(n5213), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n6579), .B2(
        n9687), .ZN(n5411) );
  NAND2_X1 U6926 ( .A1(n9465), .A2(n5700), .ZN(n5423) );
  INV_X1 U6927 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n5413) );
  NAND2_X1 U6928 ( .A1(n5414), .A2(n5413), .ZN(n5415) );
  NAND2_X1 U6929 ( .A1(n5416), .A2(n5415), .ZN(n8024) );
  OR2_X1 U6930 ( .A1(n8024), .A2(n5166), .ZN(n5421) );
  INV_X1 U6931 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n5417) );
  OR2_X1 U6932 ( .A1(n5241), .A2(n5417), .ZN(n5420) );
  INV_X1 U6933 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n8296) );
  OR2_X1 U6934 ( .A1(n5237), .A2(n8296), .ZN(n5419) );
  INV_X1 U6935 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n7917) );
  OR2_X1 U6936 ( .A1(n5111), .A2(n7917), .ZN(n5418) );
  OR2_X1 U6937 ( .A1(n7982), .A2(n5093), .ZN(n5422) );
  NAND2_X1 U6938 ( .A1(n5423), .A2(n5422), .ZN(n5424) );
  XNOR2_X1 U6939 ( .A(n5424), .B(n4286), .ZN(n5427) );
  NOR2_X1 U6940 ( .A1(n5451), .A2(n7982), .ZN(n5425) );
  AOI21_X1 U6941 ( .B1(n9465), .B2(n5621), .A(n5425), .ZN(n5426) );
  NAND2_X1 U6942 ( .A1(n5427), .A2(n5426), .ZN(n5429) );
  OR2_X1 U6943 ( .A1(n5427), .A2(n5426), .ZN(n5428) );
  NAND2_X1 U6944 ( .A1(n5429), .A2(n5428), .ZN(n8018) );
  INV_X1 U6945 ( .A(n5429), .ZN(n5430) );
  NOR2_X1 U6946 ( .A1(n8023), .A2(n5430), .ZN(n9081) );
  XNOR2_X1 U6947 ( .A(n5432), .B(n5431), .ZN(n9080) );
  XNOR2_X1 U6948 ( .A(n5436), .B(n5435), .ZN(n7039) );
  NAND2_X1 U6949 ( .A1(n7039), .A2(n6416), .ZN(n5442) );
  NAND2_X1 U6950 ( .A1(n5438), .A2(n5437), .ZN(n5439) );
  NAND2_X1 U6951 ( .A1(n5439), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5440) );
  XNOR2_X1 U6952 ( .A(n5440), .B(P1_IR_REG_18__SCAN_IN), .ZN(n8287) );
  AOI22_X1 U6953 ( .A1(n4287), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n6579), .B2(
        n8287), .ZN(n5441) );
  NAND2_X2 U6954 ( .A1(n5442), .A2(n5441), .ZN(n9453) );
  INV_X1 U6955 ( .A(n9453), .ZN(n8046) );
  INV_X1 U6956 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n5443) );
  NAND2_X1 U6957 ( .A1(n5444), .A2(n5443), .ZN(n5445) );
  NAND2_X1 U6958 ( .A1(n5456), .A2(n5445), .ZN(n9126) );
  OR2_X1 U6959 ( .A1(n9126), .A2(n5166), .ZN(n5449) );
  AOI22_X1 U6960 ( .A1(n4289), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n5446), .B2(
        P1_REG0_REG_18__SCAN_IN), .ZN(n5448) );
  NAND2_X1 U6961 ( .A1(n5586), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n5447) );
  OAI22_X1 U6962 ( .A1(n8046), .A2(n5570), .B1(n9083), .B2(n5093), .ZN(n5450)
         );
  INV_X1 U6963 ( .A(n5451), .ZN(n5696) );
  AOI22_X1 U6964 ( .A1(n9453), .A2(n5621), .B1(n5696), .B2(n9380), .ZN(n9121)
         );
  XNOR2_X1 U6965 ( .A(n5453), .B(n5452), .ZN(n7351) );
  NAND2_X1 U6966 ( .A1(n7351), .A2(n6416), .ZN(n5455) );
  AOI22_X1 U6967 ( .A1(n5213), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9757), .B2(
        n6579), .ZN(n5454) );
  NAND2_X1 U6968 ( .A1(n9447), .A2(n5700), .ZN(n5464) );
  INV_X1 U6969 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n7450) );
  NAND2_X1 U6970 ( .A1(n5456), .A2(n7450), .ZN(n5457) );
  NAND2_X1 U6971 ( .A1(n5474), .A2(n5457), .ZN(n9374) );
  OR2_X1 U6972 ( .A1(n9374), .A2(n5166), .ZN(n5462) );
  INV_X1 U6973 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n8300) );
  NAND2_X1 U6974 ( .A1(n5446), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5459) );
  NAND2_X1 U6975 ( .A1(n5586), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n5458) );
  OAI211_X1 U6976 ( .C1(n5237), .C2(n8300), .A(n5459), .B(n5458), .ZN(n5460)
         );
  INV_X1 U6977 ( .A(n5460), .ZN(n5461) );
  NAND2_X1 U6978 ( .A1(n5462), .A2(n5461), .ZN(n9174) );
  NAND2_X1 U6979 ( .A1(n9174), .A2(n5621), .ZN(n5463) );
  NAND2_X1 U6980 ( .A1(n5464), .A2(n5463), .ZN(n5465) );
  XNOR2_X1 U6981 ( .A(n5465), .B(n4286), .ZN(n5468) );
  AND2_X1 U6982 ( .A1(n5696), .A2(n9174), .ZN(n5466) );
  AOI21_X1 U6983 ( .B1(n9447), .B2(n5695), .A(n5466), .ZN(n5467) );
  NAND2_X1 U6984 ( .A1(n5468), .A2(n5467), .ZN(n5469) );
  OAI21_X1 U6985 ( .B1(n5468), .B2(n5467), .A(n5469), .ZN(n9063) );
  INV_X1 U6986 ( .A(n5469), .ZN(n9100) );
  XNOR2_X1 U6987 ( .A(n5471), .B(n5470), .ZN(n7495) );
  NAND2_X1 U6988 ( .A1(n7495), .A2(n6416), .ZN(n5473) );
  NAND2_X1 U6989 ( .A1(n4287), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n5472) );
  NAND2_X1 U6990 ( .A1(n9442), .A2(n5700), .ZN(n5483) );
  NAND2_X1 U6991 ( .A1(n5474), .A2(n9104), .ZN(n5475) );
  NAND2_X1 U6992 ( .A1(n5497), .A2(n5475), .ZN(n9354) );
  OR2_X1 U6993 ( .A1(n9354), .A2(n5166), .ZN(n5481) );
  INV_X1 U6994 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n5478) );
  NAND2_X1 U6995 ( .A1(n4289), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n5477) );
  NAND2_X1 U6996 ( .A1(n5446), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n5476) );
  OAI211_X1 U6997 ( .C1(n5111), .C2(n5478), .A(n5477), .B(n5476), .ZN(n5479)
         );
  INV_X1 U6998 ( .A(n5479), .ZN(n5480) );
  NAND2_X1 U6999 ( .A1(n5481), .A2(n5480), .ZN(n9381) );
  NAND2_X1 U7000 ( .A1(n9381), .A2(n5621), .ZN(n5482) );
  NAND2_X1 U7001 ( .A1(n5483), .A2(n5482), .ZN(n5484) );
  XNOR2_X1 U7002 ( .A(n5484), .B(n5247), .ZN(n5486) );
  AND2_X1 U7003 ( .A1(n9381), .A2(n5696), .ZN(n5485) );
  AOI21_X1 U7004 ( .B1(n9442), .B2(n5621), .A(n5485), .ZN(n5487) );
  NAND2_X1 U7005 ( .A1(n5486), .A2(n5487), .ZN(n5491) );
  INV_X1 U7006 ( .A(n5486), .ZN(n5489) );
  INV_X1 U7007 ( .A(n5487), .ZN(n5488) );
  NAND2_X1 U7008 ( .A1(n5489), .A2(n5488), .ZN(n5490) );
  AND2_X1 U7009 ( .A1(n5491), .A2(n5490), .ZN(n9099) );
  XNOR2_X1 U7010 ( .A(n5493), .B(n5492), .ZN(n7498) );
  NAND2_X1 U7011 ( .A1(n7498), .A2(n6416), .ZN(n5495) );
  NAND2_X1 U7012 ( .A1(n5213), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n5494) );
  NAND2_X1 U7013 ( .A1(n5497), .A2(n5496), .ZN(n5498) );
  AND2_X1 U7014 ( .A1(n5514), .A2(n5498), .ZN(n9339) );
  NAND2_X1 U7015 ( .A1(n9339), .A2(n5087), .ZN(n5504) );
  INV_X1 U7016 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n5501) );
  NAND2_X1 U7017 ( .A1(n4290), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5500) );
  NAND2_X1 U7018 ( .A1(n4289), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n5499) );
  OAI211_X1 U7019 ( .C1(n5501), .C2(n5111), .A(n5500), .B(n5499), .ZN(n5502)
         );
  INV_X1 U7020 ( .A(n5502), .ZN(n5503) );
  OAI22_X1 U7021 ( .A1(n9341), .A2(n5093), .B1(n9363), .B2(n5451), .ZN(n5508)
         );
  NAND2_X1 U7022 ( .A1(n9438), .A2(n5700), .ZN(n5506) );
  INV_X1 U7023 ( .A(n9363), .ZN(n9328) );
  NAND2_X1 U7024 ( .A1(n9328), .A2(n5695), .ZN(n5505) );
  NAND2_X1 U7025 ( .A1(n5506), .A2(n5505), .ZN(n5507) );
  XNOR2_X1 U7026 ( .A(n5507), .B(n7124), .ZN(n5509) );
  XOR2_X1 U7027 ( .A(n5508), .B(n5509), .Z(n9073) );
  XNOR2_X1 U7028 ( .A(n5511), .B(n5510), .ZN(n7647) );
  NAND2_X1 U7029 ( .A1(n7647), .A2(n6416), .ZN(n5513) );
  NAND2_X1 U7030 ( .A1(n4287), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n5512) );
  INV_X1 U7031 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9113) );
  NAND2_X1 U7032 ( .A1(n5514), .A2(n9113), .ZN(n5515) );
  NAND2_X1 U7033 ( .A1(n5516), .A2(n5515), .ZN(n9322) );
  OR2_X1 U7034 ( .A1(n9322), .A2(n5166), .ZN(n5522) );
  INV_X1 U7035 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n5519) );
  NAND2_X1 U7036 ( .A1(n4290), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5518) );
  NAND2_X1 U7037 ( .A1(n4289), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n5517) );
  OAI211_X1 U7038 ( .C1(n5519), .C2(n5111), .A(n5518), .B(n5517), .ZN(n5520)
         );
  INV_X1 U7039 ( .A(n5520), .ZN(n5521) );
  NAND2_X1 U7040 ( .A1(n5522), .A2(n5521), .ZN(n9346) );
  AOI22_X1 U7041 ( .A1(n9432), .A2(n5695), .B1(n5696), .B2(n9346), .ZN(n5526)
         );
  OAI22_X1 U7042 ( .A1(n9325), .A2(n5570), .B1(n9315), .B2(n5093), .ZN(n5523)
         );
  XNOR2_X1 U7043 ( .A(n5523), .B(n7124), .ZN(n9112) );
  OAI22_X1 U7044 ( .A1(n9307), .A2(n5570), .B1(n9179), .B2(n5093), .ZN(n5524)
         );
  XNOR2_X1 U7045 ( .A(n5524), .B(n4286), .ZN(n5527) );
  NAND2_X1 U7046 ( .A1(n5531), .A2(n5530), .ZN(n5549) );
  INV_X1 U7047 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7894) );
  MUX2_X1 U7048 ( .A(n7867), .B(n7894), .S(n4278), .Z(n5551) );
  XNOR2_X1 U7049 ( .A(n5551), .B(SI_24_), .ZN(n5550) );
  XNOR2_X1 U7050 ( .A(n5549), .B(n5550), .ZN(n7893) );
  NAND2_X1 U7051 ( .A1(n7893), .A2(n6416), .ZN(n5533) );
  NAND2_X1 U7052 ( .A1(n5213), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n5532) );
  NAND2_X1 U7053 ( .A1(n9423), .A2(n5700), .ZN(n5543) );
  INV_X1 U7054 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n5534) );
  NAND2_X1 U7055 ( .A1(n5535), .A2(n5534), .ZN(n5536) );
  AND2_X1 U7056 ( .A1(n5562), .A2(n5536), .ZN(n9297) );
  NAND2_X1 U7057 ( .A1(n9297), .A2(n5087), .ZN(n5541) );
  INV_X1 U7058 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n9300) );
  NAND2_X1 U7059 ( .A1(n4289), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n5538) );
  NAND2_X1 U7060 ( .A1(n5446), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5537) );
  OAI211_X1 U7061 ( .C1(n9300), .C2(n5111), .A(n5538), .B(n5537), .ZN(n5539)
         );
  INV_X1 U7062 ( .A(n5539), .ZN(n5540) );
  NAND2_X1 U7063 ( .A1(n5541), .A2(n5540), .ZN(n9283) );
  NAND2_X1 U7064 ( .A1(n9283), .A2(n5695), .ZN(n5542) );
  NAND2_X1 U7065 ( .A1(n5543), .A2(n5542), .ZN(n5544) );
  XNOR2_X1 U7066 ( .A(n5544), .B(n7124), .ZN(n5548) );
  NAND2_X1 U7067 ( .A1(n9423), .A2(n5621), .ZN(n5546) );
  NAND2_X1 U7068 ( .A1(n9283), .A2(n5696), .ZN(n5545) );
  NAND2_X1 U7069 ( .A1(n5546), .A2(n5545), .ZN(n5547) );
  NOR2_X1 U7070 ( .A1(n5548), .A2(n5547), .ZN(n5572) );
  AOI21_X1 U7071 ( .B1(n5548), .B2(n5547), .A(n5572), .ZN(n9091) );
  INV_X1 U7072 ( .A(n5551), .ZN(n5552) );
  NAND2_X1 U7073 ( .A1(n5552), .A2(SI_24_), .ZN(n5553) );
  MUX2_X1 U7074 ( .A(n7946), .B(n7942), .S(n4278), .Z(n5555) );
  INV_X1 U7075 ( .A(SI_25_), .ZN(n5554) );
  NAND2_X1 U7076 ( .A1(n5555), .A2(n5554), .ZN(n5575) );
  INV_X1 U7077 ( .A(n5555), .ZN(n5556) );
  NAND2_X1 U7078 ( .A1(n5556), .A2(SI_25_), .ZN(n5557) );
  NAND2_X1 U7079 ( .A1(n5575), .A2(n5557), .ZN(n5576) );
  NAND2_X1 U7080 ( .A1(n7940), .A2(n6416), .ZN(n5559) );
  NAND2_X1 U7081 ( .A1(n4287), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n5558) );
  INV_X1 U7082 ( .A(n5562), .ZN(n5560) );
  NAND2_X1 U7083 ( .A1(n5560), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n5584) );
  INV_X1 U7084 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n5561) );
  NAND2_X1 U7085 ( .A1(n5562), .A2(n5561), .ZN(n5563) );
  NAND2_X1 U7086 ( .A1(n5584), .A2(n5563), .ZN(n9277) );
  OR2_X1 U7087 ( .A1(n9277), .A2(n5166), .ZN(n5569) );
  INV_X1 U7088 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n5566) );
  NAND2_X1 U7089 ( .A1(n4289), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n5565) );
  NAND2_X1 U7090 ( .A1(n5446), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5564) );
  OAI211_X1 U7091 ( .C1(n5111), .C2(n5566), .A(n5565), .B(n5564), .ZN(n5567)
         );
  INV_X1 U7092 ( .A(n5567), .ZN(n5568) );
  NAND2_X1 U7093 ( .A1(n5569), .A2(n5568), .ZN(n9293) );
  OAI22_X1 U7094 ( .A1(n9280), .A2(n5093), .B1(n9266), .B2(n5451), .ZN(n5597)
         );
  OAI22_X1 U7095 ( .A1(n9280), .A2(n5570), .B1(n9266), .B2(n5093), .ZN(n5571)
         );
  XNOR2_X1 U7096 ( .A(n5571), .B(n7124), .ZN(n5596) );
  XOR2_X1 U7097 ( .A(n5597), .B(n5596), .Z(n8322) );
  AND2_X1 U7098 ( .A1(n9091), .A2(n8322), .ZN(n5574) );
  INV_X1 U7099 ( .A(n8322), .ZN(n5573) );
  INV_X1 U7100 ( .A(n5572), .ZN(n8320) );
  INV_X1 U7101 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n8015) );
  MUX2_X1 U7102 ( .A(n8015), .B(n8013), .S(n4278), .Z(n5579) );
  INV_X1 U7103 ( .A(SI_26_), .ZN(n5578) );
  NAND2_X1 U7104 ( .A1(n5579), .A2(n5578), .ZN(n5603) );
  INV_X1 U7105 ( .A(n5579), .ZN(n5580) );
  NAND2_X1 U7106 ( .A1(n5580), .A2(SI_26_), .ZN(n5581) );
  XNOR2_X1 U7107 ( .A(n5602), .B(n5601), .ZN(n8012) );
  NAND2_X1 U7108 ( .A1(n8012), .A2(n6416), .ZN(n5583) );
  NAND2_X1 U7109 ( .A1(n4287), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n5582) );
  NAND2_X1 U7110 ( .A1(n9412), .A2(n5700), .ZN(n5593) );
  INV_X1 U7111 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9143) );
  NAND2_X1 U7112 ( .A1(n5584), .A2(n9143), .ZN(n5585) );
  NAND2_X1 U7113 ( .A1(n9260), .A2(n5087), .ZN(n5591) );
  INV_X1 U7114 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n7437) );
  NAND2_X1 U7115 ( .A1(n4290), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5588) );
  NAND2_X1 U7116 ( .A1(n5586), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n5587) );
  OAI211_X1 U7117 ( .C1(n5237), .C2(n7437), .A(n5588), .B(n5587), .ZN(n5589)
         );
  INV_X1 U7118 ( .A(n5589), .ZN(n5590) );
  NAND2_X1 U7119 ( .A1(n9284), .A2(n5695), .ZN(n5592) );
  NAND2_X1 U7120 ( .A1(n5593), .A2(n5592), .ZN(n5594) );
  XNOR2_X1 U7121 ( .A(n5594), .B(n7124), .ZN(n5628) );
  NOR2_X1 U7122 ( .A1(n6472), .A2(n5451), .ZN(n5595) );
  AOI21_X1 U7123 ( .B1(n9412), .B2(n5695), .A(n5595), .ZN(n5626) );
  XNOR2_X1 U7124 ( .A(n5628), .B(n5626), .ZN(n9137) );
  INV_X1 U7125 ( .A(n5596), .ZN(n5599) );
  INV_X1 U7126 ( .A(n5597), .ZN(n5598) );
  NAND2_X1 U7127 ( .A1(n5599), .A2(n5598), .ZN(n9133) );
  INV_X1 U7128 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n8052) );
  INV_X1 U7129 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n5605) );
  MUX2_X1 U7130 ( .A(n8052), .B(n5605), .S(n4283), .Z(n5606) );
  INV_X1 U7131 ( .A(SI_27_), .ZN(n7425) );
  NAND2_X1 U7132 ( .A1(n5606), .A2(n7425), .ZN(n5692) );
  INV_X1 U7133 ( .A(n5606), .ZN(n5607) );
  NAND2_X1 U7134 ( .A1(n5607), .A2(SI_27_), .ZN(n5608) );
  NAND2_X1 U7135 ( .A1(n8029), .A2(n6416), .ZN(n5610) );
  NAND2_X1 U7136 ( .A1(n5213), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n5609) );
  NAND2_X1 U7137 ( .A1(n9248), .A2(n5700), .ZN(n5618) );
  XNOR2_X1 U7138 ( .A(n5673), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n9247) );
  NAND2_X1 U7139 ( .A1(n9247), .A2(n5087), .ZN(n5616) );
  INV_X1 U7140 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n5613) );
  NAND2_X1 U7141 ( .A1(n4288), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n5612) );
  NAND2_X1 U7142 ( .A1(n5446), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5611) );
  OAI211_X1 U7143 ( .C1(n5111), .C2(n5613), .A(n5612), .B(n5611), .ZN(n5614)
         );
  INV_X1 U7144 ( .A(n5614), .ZN(n5615) );
  NAND2_X1 U7145 ( .A1(n9228), .A2(n5621), .ZN(n5617) );
  NAND2_X1 U7146 ( .A1(n5618), .A2(n5617), .ZN(n5619) );
  XNOR2_X1 U7147 ( .A(n5619), .B(n4286), .ZN(n5623) );
  INV_X1 U7148 ( .A(n5623), .ZN(n5625) );
  NOR2_X1 U7149 ( .A1(n9267), .A2(n5451), .ZN(n5620) );
  AOI21_X1 U7150 ( .B1(n9248), .B2(n5695), .A(n5620), .ZN(n5622) );
  INV_X1 U7151 ( .A(n5622), .ZN(n5624) );
  INV_X1 U7152 ( .A(n5626), .ZN(n5627) );
  NAND2_X1 U7153 ( .A1(n5628), .A2(n5627), .ZN(n5630) );
  AOI21_X1 U7154 ( .B1(n9135), .B2(n5630), .A(n5629), .ZN(n5657) );
  NAND2_X1 U7155 ( .A1(n7648), .A2(n7499), .ZN(n7029) );
  INV_X1 U7156 ( .A(n7029), .ZN(n6710) );
  NAND2_X1 U7157 ( .A1(n7941), .A2(P1_B_REG_SCAN_IN), .ZN(n5635) );
  MUX2_X1 U7158 ( .A(n5635), .B(P1_B_REG_SCAN_IN), .S(n5634), .Z(n5636) );
  INV_X1 U7159 ( .A(n5637), .ZN(n8014) );
  NAND2_X1 U7160 ( .A1(n8014), .A2(n7941), .ZN(n6643) );
  OAI21_X1 U7161 ( .B1(n6701), .B2(P1_D_REG_1__SCAN_IN), .A(n6643), .ZN(n6706)
         );
  INV_X1 U7162 ( .A(n6706), .ZN(n7014) );
  NOR4_X1 U7163 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_15__SCAN_IN), .A3(
        P1_D_REG_16__SCAN_IN), .A4(P1_D_REG_18__SCAN_IN), .ZN(n5641) );
  NOR4_X1 U7164 ( .A1(P1_D_REG_12__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_11__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n5640) );
  NOR4_X1 U7165 ( .A1(P1_D_REG_24__SCAN_IN), .A2(P1_D_REG_25__SCAN_IN), .A3(
        P1_D_REG_26__SCAN_IN), .A4(P1_D_REG_29__SCAN_IN), .ZN(n5639) );
  NOR4_X1 U7166 ( .A1(P1_D_REG_19__SCAN_IN), .A2(P1_D_REG_20__SCAN_IN), .A3(
        P1_D_REG_21__SCAN_IN), .A4(P1_D_REG_22__SCAN_IN), .ZN(n5638) );
  AND4_X1 U7167 ( .A1(n5641), .A2(n5640), .A3(n5639), .A4(n5638), .ZN(n5647)
         );
  NOR2_X1 U7168 ( .A1(P1_D_REG_23__SCAN_IN), .A2(P1_D_REG_17__SCAN_IN), .ZN(
        n5645) );
  NOR4_X1 U7169 ( .A1(P1_D_REG_27__SCAN_IN), .A2(P1_D_REG_28__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_4__SCAN_IN), .ZN(n5644) );
  NOR4_X1 U7170 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_7__SCAN_IN), .ZN(n5643) );
  NOR4_X1 U7171 ( .A1(P1_D_REG_8__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_31__SCAN_IN), .A4(P1_D_REG_6__SCAN_IN), .ZN(n5642) );
  AND4_X1 U7172 ( .A1(n5645), .A2(n5644), .A3(n5643), .A4(n5642), .ZN(n5646)
         );
  NAND2_X1 U7173 ( .A1(n5647), .A2(n5646), .ZN(n6699) );
  INV_X1 U7174 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n7428) );
  NOR2_X1 U7175 ( .A1(n6699), .A2(n7428), .ZN(n5648) );
  NAND2_X1 U7176 ( .A1(n8014), .A2(n7896), .ZN(n9491) );
  OAI21_X1 U7177 ( .B1(n6701), .B2(n5648), .A(n9491), .ZN(n6715) );
  INV_X1 U7178 ( .A(n6715), .ZN(n5649) );
  NAND2_X1 U7179 ( .A1(n7014), .A2(n5649), .ZN(n5667) );
  INV_X1 U7180 ( .A(n5650), .ZN(n5651) );
  NAND2_X1 U7181 ( .A1(n5651), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5653) );
  INV_X1 U7182 ( .A(n6688), .ZN(n6563) );
  OR2_X1 U7183 ( .A1(n5667), .A2(n6563), .ZN(n5659) );
  INV_X1 U7184 ( .A(n6708), .ZN(n7025) );
  NOR2_X1 U7185 ( .A1(n5659), .A2(n7025), .ZN(n5656) );
  NOR2_X1 U7186 ( .A1(n7029), .A2(n5658), .ZN(n9753) );
  INV_X1 U7187 ( .A(n5659), .ZN(n5670) );
  NAND2_X1 U7188 ( .A1(n9753), .A2(n5670), .ZN(n5662) );
  NAND2_X1 U7189 ( .A1(n7499), .A2(n6688), .ZN(n5661) );
  OR2_X1 U7190 ( .A1(n6708), .A2(n5663), .ZN(n6689) );
  AND3_X1 U7191 ( .A1(n6689), .A2(n6568), .A3(n6558), .ZN(n5665) );
  INV_X1 U7192 ( .A(n5667), .ZN(n5664) );
  OR2_X1 U7193 ( .A1(n9856), .A2(n5664), .ZN(n6690) );
  NAND2_X1 U7194 ( .A1(n5665), .A2(n6690), .ZN(n5666) );
  NAND2_X1 U7195 ( .A1(n5666), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5669) );
  AND2_X1 U7196 ( .A1(n5667), .A2(n6688), .ZN(n5668) );
  NAND2_X1 U7197 ( .A1(n9753), .A2(n5668), .ZN(n6692) );
  OR2_X1 U7198 ( .A1(n7017), .A2(n5064), .ZN(n7125) );
  INV_X1 U7199 ( .A(n7125), .ZN(n6709) );
  NAND2_X1 U7200 ( .A1(n5670), .A2(n6709), .ZN(n5683) );
  INV_X1 U7201 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n5672) );
  OAI22_X1 U7202 ( .A1(n6472), .A2(n9114), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n5672), .ZN(n5685) );
  INV_X1 U7203 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n5710) );
  OAI21_X1 U7204 ( .B1(n5673), .B2(n5672), .A(n5710), .ZN(n5676) );
  INV_X1 U7205 ( .A(n5673), .ZN(n5675) );
  AND2_X1 U7206 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n5674) );
  NAND2_X1 U7207 ( .A1(n5675), .A2(n5674), .ZN(n9213) );
  NAND2_X1 U7208 ( .A1(n5676), .A2(n9213), .ZN(n9223) );
  OR2_X1 U7209 ( .A1(n9223), .A2(n5166), .ZN(n5682) );
  INV_X1 U7210 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n5679) );
  NAND2_X1 U7211 ( .A1(n4289), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n5678) );
  NAND2_X1 U7212 ( .A1(n5446), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5677) );
  OAI211_X1 U7213 ( .C1(n5679), .C2(n5111), .A(n5678), .B(n5677), .ZN(n5680)
         );
  INV_X1 U7214 ( .A(n5680), .ZN(n5681) );
  NOR2_X1 U7215 ( .A1(n9245), .A2(n9123), .ZN(n5684) );
  AOI211_X1 U7216 ( .C1(n9247), .C2(n9140), .A(n5685), .B(n5684), .ZN(n5686)
         );
  INV_X1 U7217 ( .A(n5687), .ZN(n5688) );
  NAND2_X1 U7218 ( .A1(n5689), .A2(n5688), .ZN(P1_U3212) );
  INV_X1 U7219 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8461) );
  INV_X1 U7220 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n8056) );
  MUX2_X1 U7221 ( .A(n8461), .B(n8056), .S(n4283), .Z(n6386) );
  XNOR2_X1 U7222 ( .A(n6386), .B(SI_28_), .ZN(n6383) );
  NAND2_X1 U7223 ( .A1(n8459), .A2(n6416), .ZN(n5694) );
  NAND2_X1 U7224 ( .A1(n5213), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n5693) );
  NAND2_X1 U7225 ( .A1(n9401), .A2(n5621), .ZN(n5698) );
  NAND2_X1 U7226 ( .A1(n9208), .A2(n5696), .ZN(n5697) );
  NAND2_X1 U7227 ( .A1(n5698), .A2(n5697), .ZN(n5699) );
  XNOR2_X1 U7228 ( .A(n5699), .B(n7124), .ZN(n5702) );
  AOI22_X1 U7229 ( .A1(n9401), .A2(n5700), .B1(n5621), .B2(n9208), .ZN(n5701)
         );
  XNOR2_X1 U7230 ( .A(n5702), .B(n5701), .ZN(n5704) );
  AND2_X1 U7231 ( .A1(n5704), .A2(n9136), .ZN(n5716) );
  NAND3_X1 U7232 ( .A1(n5704), .A2(n5703), .A3(n9136), .ZN(n5715) );
  OR2_X1 U7233 ( .A1(n9213), .A2(n5166), .ZN(n5709) );
  INV_X1 U7234 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n7460) );
  NAND2_X1 U7235 ( .A1(n4289), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n5706) );
  NAND2_X1 U7236 ( .A1(n5446), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n5705) );
  OAI211_X1 U7237 ( .C1(n7460), .C2(n5111), .A(n5706), .B(n5705), .ZN(n5707)
         );
  INV_X1 U7238 ( .A(n5707), .ZN(n5708) );
  NAND2_X1 U7239 ( .A1(n5709), .A2(n5708), .ZN(n9229) );
  OAI22_X1 U7240 ( .A1(n9223), .A2(n9127), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n5710), .ZN(n5711) );
  AOI21_X1 U7241 ( .B1(n9145), .B2(n9229), .A(n5711), .ZN(n5712) );
  OAI21_X1 U7242 ( .B1(n9267), .B2(n9114), .A(n5712), .ZN(n5713) );
  AOI21_X1 U7243 ( .B1(n9401), .B2(n9129), .A(n5713), .ZN(n5714) );
  NAND3_X1 U7244 ( .A1(n5943), .A2(n5946), .A3(n5720), .ZN(n5975) );
  NOR2_X1 U7245 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n5725) );
  NOR2_X1 U7246 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_25__SCAN_IN), .ZN(
        n5724) );
  NOR2_X1 U7247 ( .A1(P2_IR_REG_26__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .ZN(
        n5723) );
  NAND4_X1 U7248 ( .A1(n5726), .A2(n5725), .A3(n5724), .A4(n5723), .ZN(n5727)
         );
  INV_X1 U7249 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5728) );
  NAND2_X1 U7250 ( .A1(n5731), .A2(n5730), .ZN(n5733) );
  XNOR2_X2 U7251 ( .A(n5734), .B(P2_IR_REG_30__SCAN_IN), .ZN(n5736) );
  NAND2_X1 U7252 ( .A1(n4275), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6917) );
  INV_X1 U7253 ( .A(n5736), .ZN(n8059) );
  AND2_X2 U7254 ( .A1(n5736), .A2(n9050), .ZN(n6148) );
  NAND2_X1 U7255 ( .A1(n6148), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n6915) );
  INV_X1 U7256 ( .A(n6008), .ZN(n5739) );
  NAND2_X1 U7257 ( .A1(n5741), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5743) );
  INV_X1 U7258 ( .A(n5744), .ZN(n5745) );
  NAND2_X1 U7259 ( .A1(n5750), .A2(n5746), .ZN(n5747) );
  NAND2_X1 U7260 ( .A1(n5747), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5749) );
  INV_X1 U7261 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6633) );
  XNOR2_X1 U7262 ( .A(n6108), .B(n8414), .ZN(n5762) );
  XNOR2_X1 U7263 ( .A(n5764), .B(n5762), .ZN(n8417) );
  NAND2_X1 U7264 ( .A1(n4275), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6925) );
  NAND2_X1 U7265 ( .A1(n6148), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6922) );
  NAND4_X1 U7266 ( .A1(n6923), .A2(n6925), .A3(n6922), .A4(n6924), .ZN(n5759)
         );
  NAND2_X1 U7267 ( .A1(n4873), .A2(SI_0_), .ZN(n5758) );
  XNOR2_X1 U7268 ( .A(n5758), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n9052) );
  NAND2_X1 U7269 ( .A1(n7067), .A2(n5760), .ZN(n8407) );
  OR2_X1 U7270 ( .A1(n6108), .A2(n9952), .ZN(n5761) );
  AND2_X1 U7271 ( .A1(n8407), .A2(n5761), .ZN(n8416) );
  NAND2_X1 U7272 ( .A1(n8417), .A2(n8416), .ZN(n8415) );
  INV_X1 U7273 ( .A(n5762), .ZN(n5763) );
  NAND2_X1 U7274 ( .A1(n5764), .A2(n5763), .ZN(n5765) );
  AND2_X1 U7275 ( .A1(n8415), .A2(n5765), .ZN(n8377) );
  NAND2_X1 U7276 ( .A1(n4275), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5769) );
  NAND2_X1 U7277 ( .A1(n5792), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5768) );
  NAND2_X1 U7278 ( .A1(n5806), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5767) );
  NAND2_X1 U7279 ( .A1(n6148), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5766) );
  OR2_X1 U7280 ( .A1(n7072), .A2(n7043), .ZN(n5775) );
  OR2_X1 U7281 ( .A1(n5757), .A2(n5728), .ZN(n5771) );
  INV_X1 U7282 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5770) );
  XNOR2_X1 U7283 ( .A(n8373), .B(n6152), .ZN(n5776) );
  NAND2_X1 U7284 ( .A1(n5775), .A2(n5776), .ZN(n5774) );
  NAND2_X1 U7285 ( .A1(n8377), .A2(n5774), .ZN(n8378) );
  INV_X1 U7286 ( .A(n5775), .ZN(n5777) );
  INV_X1 U7287 ( .A(n5776), .ZN(n8371) );
  NAND2_X1 U7288 ( .A1(n5777), .A2(n8371), .ZN(n8376) );
  NAND2_X1 U7289 ( .A1(n5806), .A2(n9924), .ZN(n5781) );
  NAND2_X1 U7290 ( .A1(n4275), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5780) );
  NAND2_X1 U7291 ( .A1(n5792), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5779) );
  NAND2_X1 U7292 ( .A1(n6148), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5778) );
  NOR2_X1 U7293 ( .A1(n7074), .A2(n7043), .ZN(n5786) );
  OR3_X1 U7294 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .A3(
        P2_IR_REG_0__SCAN_IN), .ZN(n5782) );
  NAND2_X1 U7295 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n5782), .ZN(n5783) );
  XNOR2_X1 U7296 ( .A(n5783), .B(P2_IR_REG_3__SCAN_IN), .ZN(n6254) );
  INV_X1 U7297 ( .A(n6254), .ZN(n7006) );
  OR2_X1 U7298 ( .A1(n5797), .A2(n6630), .ZN(n5784) );
  XNOR2_X1 U7299 ( .A(n9932), .B(n6108), .ZN(n7045) );
  NAND2_X1 U7300 ( .A1(n5786), .A2(n7045), .ZN(n5803) );
  INV_X1 U7301 ( .A(n5786), .ZN(n5788) );
  INV_X1 U7302 ( .A(n7045), .ZN(n5787) );
  NAND2_X1 U7303 ( .A1(n5788), .A2(n5787), .ZN(n5789) );
  AND2_X1 U7304 ( .A1(n5803), .A2(n5789), .ZN(n8482) );
  INV_X1 U7305 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n5790) );
  NAND2_X1 U7306 ( .A1(n9924), .A2(n5790), .ZN(n5791) );
  NAND2_X1 U7307 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5808) );
  AND2_X1 U7308 ( .A1(n5791), .A2(n5808), .ZN(n7522) );
  NAND2_X1 U7309 ( .A1(n6093), .A2(n7522), .ZN(n5796) );
  NAND2_X1 U7310 ( .A1(n6068), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5795) );
  NAND2_X1 U7311 ( .A1(n6148), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5794) );
  NAND2_X1 U7312 ( .A1(n6722), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5793) );
  NAND2_X1 U7313 ( .A1(n8619), .A2(n5760), .ZN(n5805) );
  OR2_X1 U7314 ( .A1(n6082), .A2(n6631), .ZN(n5802) );
  OR2_X1 U7315 ( .A1(n5797), .A2(n6632), .ZN(n5801) );
  NAND2_X1 U7316 ( .A1(n5798), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5799) );
  XNOR2_X1 U7317 ( .A(n5799), .B(n4806), .ZN(n6958) );
  OR2_X1 U7318 ( .A1(n6286), .A2(n6958), .ZN(n5800) );
  XNOR2_X1 U7319 ( .A(n7531), .B(n6152), .ZN(n7342) );
  XNOR2_X1 U7320 ( .A(n5805), .B(n7342), .ZN(n7044) );
  INV_X1 U7321 ( .A(n7342), .ZN(n5804) );
  INV_X1 U7322 ( .A(n5808), .ZN(n5807) );
  NAND2_X1 U7323 ( .A1(n5807), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5836) );
  INV_X1 U7324 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n7341) );
  NAND2_X1 U7325 ( .A1(n5808), .A2(n7341), .ZN(n5809) );
  AND2_X1 U7326 ( .A1(n5836), .A2(n5809), .ZN(n7663) );
  NAND2_X1 U7327 ( .A1(n6093), .A2(n7663), .ZN(n5813) );
  NAND2_X1 U7328 ( .A1(n6068), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5812) );
  NAND2_X1 U7329 ( .A1(n6148), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5811) );
  NAND2_X1 U7330 ( .A1(n6722), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5810) );
  OR2_X1 U7331 ( .A1(n7079), .A2(n7043), .ZN(n5818) );
  OR2_X1 U7332 ( .A1(n5814), .A2(n5728), .ZN(n5824) );
  XNOR2_X1 U7333 ( .A(n5824), .B(P2_IR_REG_5__SCAN_IN), .ZN(n6252) );
  INV_X1 U7334 ( .A(n6252), .ZN(n6982) );
  OR2_X1 U7335 ( .A1(n5797), .A2(n6627), .ZN(n5816) );
  OR2_X1 U7336 ( .A1(n6082), .A2(n6628), .ZN(n5815) );
  OAI211_X1 U7337 ( .C1(n6286), .C2(n6982), .A(n5816), .B(n5815), .ZN(n7661)
         );
  XNOR2_X1 U7338 ( .A(n7661), .B(n6108), .ZN(n8391) );
  XNOR2_X1 U7339 ( .A(n5818), .B(n8391), .ZN(n7344) );
  INV_X1 U7340 ( .A(n8391), .ZN(n5817) );
  NAND2_X1 U7341 ( .A1(n5818), .A2(n5817), .ZN(n5819) );
  NAND2_X1 U7342 ( .A1(n8402), .A2(n5819), .ZN(n5828) );
  XNOR2_X1 U7343 ( .A(n5836), .B(P2_REG3_REG_6__SCAN_IN), .ZN(n8394) );
  NAND2_X1 U7344 ( .A1(n6093), .A2(n8394), .ZN(n5823) );
  NAND2_X1 U7345 ( .A1(n6068), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5822) );
  NAND2_X1 U7346 ( .A1(n6148), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5821) );
  NAND2_X1 U7347 ( .A1(n6722), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5820) );
  OR2_X1 U7348 ( .A1(n7727), .A2(n7043), .ZN(n5831) );
  NAND2_X1 U7349 ( .A1(n5824), .A2(n4715), .ZN(n5825) );
  NAND2_X1 U7350 ( .A1(n5825), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5842) );
  XNOR2_X1 U7351 ( .A(n5842), .B(P2_IR_REG_6__SCAN_IN), .ZN(n6250) );
  INV_X1 U7352 ( .A(n6250), .ZN(n6946) );
  OR2_X1 U7353 ( .A1(n5797), .A2(n6641), .ZN(n5827) );
  OR2_X1 U7354 ( .A1(n6082), .A2(n6639), .ZN(n5826) );
  OAI211_X1 U7355 ( .C1(n6286), .C2(n6946), .A(n5827), .B(n5826), .ZN(n8398)
         );
  XNOR2_X1 U7356 ( .A(n6108), .B(n8398), .ZN(n5829) );
  XNOR2_X1 U7357 ( .A(n5831), .B(n5829), .ZN(n8392) );
  INV_X1 U7358 ( .A(n5829), .ZN(n5830) );
  NAND2_X1 U7359 ( .A1(n5831), .A2(n5830), .ZN(n5832) );
  INV_X1 U7360 ( .A(n5836), .ZN(n5834) );
  AND2_X1 U7361 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_REG3_REG_6__SCAN_IN), 
        .ZN(n5833) );
  NAND2_X1 U7362 ( .A1(n5834), .A2(n5833), .ZN(n5854) );
  INV_X1 U7363 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n6940) );
  INV_X1 U7364 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5835) );
  OAI21_X1 U7365 ( .B1(n5836), .B2(n6940), .A(n5835), .ZN(n5837) );
  AND2_X1 U7366 ( .A1(n5854), .A2(n5837), .ZN(n7735) );
  NAND2_X1 U7367 ( .A1(n6093), .A2(n7735), .ZN(n5841) );
  NAND2_X1 U7368 ( .A1(n6068), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5840) );
  NAND2_X1 U7369 ( .A1(n6721), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5839) );
  NAND2_X1 U7370 ( .A1(n6722), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5838) );
  NOR2_X1 U7371 ( .A1(n8396), .A2(n7043), .ZN(n5847) );
  NAND2_X1 U7372 ( .A1(n5842), .A2(n4716), .ZN(n5843) );
  NAND2_X1 U7373 ( .A1(n5843), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5844) );
  XNOR2_X1 U7374 ( .A(n5844), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6248) );
  INV_X1 U7375 ( .A(n6248), .ZN(n6970) );
  OR2_X1 U7376 ( .A1(n5797), .A2(n6648), .ZN(n5846) );
  OR2_X1 U7377 ( .A1(n6082), .A2(n6646), .ZN(n5845) );
  OAI211_X1 U7378 ( .C1(n6286), .C2(n6970), .A(n5846), .B(n5845), .ZN(n7734)
         );
  XNOR2_X1 U7379 ( .A(n7734), .B(n6108), .ZN(n7599) );
  NAND2_X1 U7380 ( .A1(n5847), .A2(n7599), .ZN(n5852) );
  INV_X1 U7381 ( .A(n5847), .ZN(n5849) );
  INV_X1 U7382 ( .A(n7599), .ZN(n5848) );
  NAND2_X1 U7383 ( .A1(n5849), .A2(n5848), .ZN(n5850) );
  NAND2_X1 U7384 ( .A1(n5852), .A2(n5850), .ZN(n6570) );
  NAND2_X1 U7385 ( .A1(n6569), .A2(n5852), .ZN(n7534) );
  INV_X1 U7386 ( .A(n5854), .ZN(n5853) );
  NAND2_X1 U7387 ( .A1(n5853), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5884) );
  INV_X1 U7388 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n6831) );
  NAND2_X1 U7389 ( .A1(n5854), .A2(n6831), .ZN(n5855) );
  AND2_X1 U7390 ( .A1(n5884), .A2(n5855), .ZN(n7692) );
  NAND2_X1 U7391 ( .A1(n6093), .A2(n7692), .ZN(n5859) );
  NAND2_X1 U7392 ( .A1(n6068), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5858) );
  NAND2_X1 U7393 ( .A1(n6721), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5857) );
  NAND2_X1 U7394 ( .A1(n6722), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5856) );
  NOR2_X1 U7395 ( .A1(n7726), .A2(n7043), .ZN(n5866) );
  NAND2_X1 U7396 ( .A1(n5860), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5861) );
  MUX2_X1 U7397 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5861), .S(
        P2_IR_REG_8__SCAN_IN), .Z(n5862) );
  NAND2_X1 U7398 ( .A1(n5862), .A2(n4300), .ZN(n6843) );
  OR2_X1 U7399 ( .A1(n5797), .A2(n5863), .ZN(n5865) );
  OR2_X1 U7400 ( .A1(n6082), .A2(n6652), .ZN(n5864) );
  OAI211_X1 U7401 ( .C1(n6286), .C2(n6843), .A(n5865), .B(n5864), .ZN(n7702)
         );
  XNOR2_X1 U7402 ( .A(n7702), .B(n6108), .ZN(n7536) );
  NAND2_X1 U7403 ( .A1(n5866), .A2(n7536), .ZN(n5898) );
  INV_X1 U7404 ( .A(n5866), .ZN(n5868) );
  INV_X1 U7405 ( .A(n7536), .ZN(n5867) );
  NAND2_X1 U7406 ( .A1(n5868), .A2(n5867), .ZN(n5869) );
  AND2_X1 U7407 ( .A1(n5898), .A2(n5869), .ZN(n7600) );
  INV_X1 U7408 ( .A(n5886), .ZN(n5870) );
  NAND2_X1 U7409 ( .A1(n5870), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5919) );
  INV_X1 U7410 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n6893) );
  NAND2_X1 U7411 ( .A1(n5886), .A2(n6893), .ZN(n5871) );
  AND2_X1 U7412 ( .A1(n5919), .A2(n5871), .ZN(n7884) );
  NAND2_X1 U7413 ( .A1(n6093), .A2(n7884), .ZN(n5875) );
  NAND2_X1 U7414 ( .A1(n6068), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5874) );
  NAND2_X1 U7415 ( .A1(n6721), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5873) );
  NAND2_X1 U7416 ( .A1(n6722), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5872) );
  NOR2_X1 U7417 ( .A1(n7779), .A2(n7043), .ZN(n5880) );
  OR2_X1 U7418 ( .A1(n4300), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n5876) );
  NAND2_X1 U7419 ( .A1(n5876), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5877) );
  XNOR2_X1 U7420 ( .A(n5877), .B(P2_IR_REG_10__SCAN_IN), .ZN(n6659) );
  AOI22_X1 U7421 ( .A1(n6023), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6022), .B2(
        n6659), .ZN(n5879) );
  NAND2_X1 U7422 ( .A1(n6657), .A2(n8084), .ZN(n5878) );
  XNOR2_X1 U7423 ( .A(n7887), .B(n6108), .ZN(n5881) );
  INV_X1 U7424 ( .A(n5900), .ZN(n5894) );
  INV_X1 U7425 ( .A(n5880), .ZN(n5882) );
  INV_X1 U7426 ( .A(n5881), .ZN(n7760) );
  NAND2_X1 U7427 ( .A1(n5884), .A2(n5883), .ZN(n5885) );
  AND2_X1 U7428 ( .A1(n5886), .A2(n5885), .ZN(n7718) );
  NAND2_X1 U7429 ( .A1(n6093), .A2(n7718), .ZN(n5890) );
  NAND2_X1 U7430 ( .A1(n6068), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5889) );
  NAND2_X1 U7431 ( .A1(n6721), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5888) );
  NAND2_X1 U7432 ( .A1(n6722), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5887) );
  OR2_X1 U7433 ( .A1(n7889), .A2(n7043), .ZN(n5897) );
  NAND2_X1 U7434 ( .A1(n4300), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5891) );
  XNOR2_X1 U7435 ( .A(n5891), .B(P2_IR_REG_9__SCAN_IN), .ZN(n6264) );
  INV_X1 U7436 ( .A(n6264), .ZN(n6994) );
  OR2_X1 U7437 ( .A1(n6082), .A2(n6653), .ZN(n5892) );
  XNOR2_X1 U7438 ( .A(n7721), .B(n6152), .ZN(n5896) );
  NAND2_X1 U7439 ( .A1(n5897), .A2(n5896), .ZN(n7758) );
  OR2_X1 U7440 ( .A1(n5894), .A2(n5893), .ZN(n5895) );
  XNOR2_X1 U7441 ( .A(n5897), .B(n5896), .ZN(n7538) );
  INV_X1 U7442 ( .A(n5898), .ZN(n5899) );
  NOR2_X1 U7443 ( .A1(n7538), .A2(n5899), .ZN(n7535) );
  NAND2_X1 U7444 ( .A1(n6666), .A2(n8084), .ZN(n5904) );
  NAND2_X1 U7445 ( .A1(n5901), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5902) );
  XNOR2_X1 U7446 ( .A(n5902), .B(P2_IR_REG_11__SCAN_IN), .ZN(n6265) );
  AOI22_X1 U7447 ( .A1(n6023), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6022), .B2(
        n6265), .ZN(n5903) );
  NAND2_X1 U7448 ( .A1(n5904), .A2(n5903), .ZN(n7988) );
  XNOR2_X1 U7449 ( .A(n7988), .B(n6108), .ZN(n5910) );
  XNOR2_X1 U7450 ( .A(n5919), .B(P2_REG3_REG_11__SCAN_IN), .ZN(n7764) );
  NAND2_X1 U7451 ( .A1(n6093), .A2(n7764), .ZN(n5908) );
  NAND2_X1 U7452 ( .A1(n6068), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5907) );
  NAND2_X1 U7453 ( .A1(n6721), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n5906) );
  NAND2_X1 U7454 ( .A1(n6722), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5905) );
  OR2_X1 U7455 ( .A1(n7904), .A2(n7043), .ZN(n5909) );
  INV_X1 U7456 ( .A(n5909), .ZN(n5911) );
  NAND2_X1 U7457 ( .A1(n6674), .A2(n8084), .ZN(n5915) );
  OR2_X1 U7458 ( .A1(n5912), .A2(n5728), .ZN(n5913) );
  XNOR2_X1 U7459 ( .A(n5913), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7240) );
  AOI22_X1 U7460 ( .A1(n6023), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6022), .B2(
        n7240), .ZN(n5914) );
  XNOR2_X1 U7461 ( .A(n10020), .B(n6108), .ZN(n5926) );
  INV_X1 U7462 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n5917) );
  INV_X1 U7463 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n5916) );
  OAI21_X1 U7464 ( .B1(n5919), .B2(n5917), .A(n5916), .ZN(n5920) );
  NAND2_X1 U7465 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_REG3_REG_11__SCAN_IN), 
        .ZN(n5918) );
  AND2_X1 U7466 ( .A1(n5920), .A2(n5933), .ZN(n9904) );
  NAND2_X1 U7467 ( .A1(n6093), .A2(n9904), .ZN(n5924) );
  NAND2_X1 U7468 ( .A1(n6068), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5923) );
  NAND2_X1 U7469 ( .A1(n6721), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5922) );
  NAND2_X1 U7470 ( .A1(n6722), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5921) );
  NAND4_X1 U7471 ( .A1(n5924), .A2(n5923), .A3(n5922), .A4(n5921), .ZN(n8611)
         );
  NAND2_X1 U7472 ( .A1(n8611), .A2(n5760), .ZN(n5927) );
  NAND2_X1 U7473 ( .A1(n5926), .A2(n5927), .ZN(n5925) );
  NAND2_X1 U7474 ( .A1(n7900), .A2(n5925), .ZN(n7897) );
  INV_X1 U7475 ( .A(n5926), .ZN(n7902) );
  INV_X1 U7476 ( .A(n5927), .ZN(n5928) );
  NAND2_X1 U7477 ( .A1(n7902), .A2(n5928), .ZN(n7898) );
  NAND2_X1 U7478 ( .A1(n6679), .A2(n8084), .ZN(n5931) );
  NAND2_X1 U7479 ( .A1(n5976), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5944) );
  XNOR2_X1 U7480 ( .A(n5944), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7629) );
  AOI22_X1 U7481 ( .A1(n6023), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6022), .B2(
        n7629), .ZN(n5930) );
  XNOR2_X1 U7482 ( .A(n8426), .B(n6108), .ZN(n5939) );
  INV_X1 U7483 ( .A(n5933), .ZN(n5932) );
  NAND2_X1 U7484 ( .A1(n5932), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5968) );
  INV_X1 U7485 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n7630) );
  NAND2_X1 U7486 ( .A1(n5933), .A2(n7630), .ZN(n5934) );
  AND2_X1 U7487 ( .A1(n5968), .A2(n5934), .ZN(n8006) );
  NAND2_X1 U7488 ( .A1(n6093), .A2(n8006), .ZN(n5938) );
  NAND2_X1 U7489 ( .A1(n6068), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n5937) );
  NAND2_X1 U7490 ( .A1(n6721), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5936) );
  NAND2_X1 U7491 ( .A1(n6722), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5935) );
  NAND4_X1 U7492 ( .A1(n5938), .A2(n5937), .A3(n5936), .A4(n5935), .ZN(n8610)
         );
  AND2_X1 U7493 ( .A1(n8610), .A2(n5760), .ZN(n5940) );
  NAND2_X1 U7494 ( .A1(n5939), .A2(n5940), .ZN(n5955) );
  INV_X1 U7495 ( .A(n5939), .ZN(n7926) );
  INV_X1 U7496 ( .A(n5940), .ZN(n5941) );
  NAND2_X1 U7497 ( .A1(n7926), .A2(n5941), .ZN(n5942) );
  AND2_X1 U7498 ( .A1(n5955), .A2(n5942), .ZN(n7773) );
  NAND2_X1 U7499 ( .A1(n6683), .A2(n8084), .ZN(n5950) );
  NAND2_X1 U7500 ( .A1(n5944), .A2(n5943), .ZN(n5945) );
  NAND2_X1 U7501 ( .A1(n5945), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5947) );
  NAND2_X1 U7502 ( .A1(n5947), .A2(n5946), .ZN(n5961) );
  OR2_X1 U7503 ( .A1(n5947), .A2(n5946), .ZN(n5948) );
  AOI22_X1 U7504 ( .A1(n6023), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6022), .B2(
        n7751), .ZN(n5949) );
  XNOR2_X1 U7505 ( .A(n8927), .B(n6152), .ZN(n5959) );
  XNOR2_X1 U7506 ( .A(n5968), .B(P2_REG3_REG_14__SCAN_IN), .ZN(n8931) );
  NAND2_X1 U7507 ( .A1(n6093), .A2(n8931), .ZN(n5954) );
  NAND2_X1 U7508 ( .A1(n6068), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n5953) );
  NAND2_X1 U7509 ( .A1(n5792), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5952) );
  NAND2_X1 U7510 ( .A1(n6721), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n5951) );
  NOR2_X1 U7511 ( .A1(n8904), .A2(n7043), .ZN(n5957) );
  XNOR2_X1 U7512 ( .A(n5959), .B(n5957), .ZN(n7939) );
  AND2_X1 U7513 ( .A1(n7939), .A2(n5955), .ZN(n5956) );
  NAND2_X1 U7514 ( .A1(n7925), .A2(n5956), .ZN(n7934) );
  INV_X1 U7515 ( .A(n5957), .ZN(n5958) );
  NAND2_X1 U7516 ( .A1(n5959), .A2(n5958), .ZN(n5960) );
  NAND2_X1 U7517 ( .A1(n5961), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5962) );
  XNOR2_X1 U7518 ( .A(n5962), .B(P2_IR_REG_15__SCAN_IN), .ZN(n6270) );
  AOI22_X1 U7519 ( .A1(n6023), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n6022), .B2(
        n6270), .ZN(n5963) );
  XNOR2_X1 U7520 ( .A(n8911), .B(n6152), .ZN(n5964) );
  INV_X1 U7521 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n5967) );
  OAI21_X1 U7522 ( .B1(n5968), .B2(n5967), .A(n7952), .ZN(n5969) );
  AND2_X1 U7523 ( .A1(n5969), .A2(n5982), .ZN(n8910) );
  NAND2_X1 U7524 ( .A1(n6093), .A2(n8910), .ZN(n5973) );
  NAND2_X1 U7525 ( .A1(n4275), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n5972) );
  NAND2_X1 U7526 ( .A1(n6721), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n5971) );
  NAND2_X1 U7527 ( .A1(n6722), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5970) );
  NAND2_X1 U7528 ( .A1(n6881), .A2(n8084), .ZN(n5980) );
  OR2_X1 U7529 ( .A1(n5976), .A2(n5975), .ZN(n5977) );
  NAND2_X1 U7530 ( .A1(n5977), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5978) );
  XNOR2_X1 U7531 ( .A(n5978), .B(P2_IR_REG_16__SCAN_IN), .ZN(n8628) );
  AOI22_X1 U7532 ( .A1(n6023), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6022), .B2(
        n8628), .ZN(n5979) );
  XNOR2_X1 U7533 ( .A(n9015), .B(n6152), .ZN(n5989) );
  INV_X1 U7534 ( .A(n5982), .ZN(n5981) );
  NAND2_X1 U7535 ( .A1(n5981), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5997) );
  INV_X1 U7536 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n8626) );
  NAND2_X1 U7537 ( .A1(n5982), .A2(n8626), .ZN(n5983) );
  AND2_X1 U7538 ( .A1(n5997), .A2(n5983), .ZN(n8890) );
  NAND2_X1 U7539 ( .A1(n6093), .A2(n8890), .ZN(n5987) );
  NAND2_X1 U7540 ( .A1(n4275), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n5986) );
  NAND2_X1 U7541 ( .A1(n6721), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n5985) );
  NAND2_X1 U7542 ( .A1(n6722), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5984) );
  NAND4_X1 U7543 ( .A1(n5987), .A2(n5986), .A3(n5985), .A4(n5984), .ZN(n8860)
         );
  NAND2_X1 U7544 ( .A1(n8860), .A2(n5760), .ZN(n5988) );
  XNOR2_X1 U7545 ( .A(n5989), .B(n5988), .ZN(n8524) );
  NAND2_X1 U7546 ( .A1(n5989), .A2(n5988), .ZN(n5990) );
  NAND2_X1 U7547 ( .A1(n7009), .A2(n8084), .ZN(n5995) );
  AND2_X1 U7548 ( .A1(n5929), .A2(n5991), .ZN(n5992) );
  OR2_X1 U7549 ( .A1(n5992), .A2(n5728), .ZN(n5993) );
  XNOR2_X1 U7550 ( .A(n5993), .B(P2_IR_REG_17__SCAN_IN), .ZN(n6246) );
  AOI22_X1 U7551 ( .A1(n6023), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6022), .B2(
        n6246), .ZN(n5994) );
  XNOR2_X1 U7552 ( .A(n9012), .B(n6108), .ZN(n6003) );
  INV_X1 U7553 ( .A(n5997), .ZN(n5996) );
  NAND2_X1 U7554 ( .A1(n5996), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n6012) );
  INV_X1 U7555 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8533) );
  NAND2_X1 U7556 ( .A1(n5997), .A2(n8533), .ZN(n5998) );
  AND2_X1 U7557 ( .A1(n6012), .A2(n5998), .ZN(n8869) );
  NAND2_X1 U7558 ( .A1(n6093), .A2(n8869), .ZN(n6002) );
  NAND2_X1 U7559 ( .A1(n4275), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n6001) );
  NAND2_X1 U7560 ( .A1(n6148), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n6000) );
  NAND2_X1 U7561 ( .A1(n6722), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5999) );
  NAND4_X1 U7562 ( .A1(n6002), .A2(n6001), .A3(n6000), .A4(n5999), .ZN(n8850)
         );
  AND2_X1 U7563 ( .A1(n8850), .A2(n5760), .ZN(n6004) );
  NAND2_X1 U7564 ( .A1(n6003), .A2(n6004), .ZN(n6007) );
  INV_X1 U7565 ( .A(n6003), .ZN(n8574) );
  INV_X1 U7566 ( .A(n6004), .ZN(n6005) );
  NAND2_X1 U7567 ( .A1(n8574), .A2(n6005), .ZN(n6006) );
  NAND2_X1 U7568 ( .A1(n6007), .A2(n6006), .ZN(n8530) );
  NAND2_X1 U7569 ( .A1(n7039), .A2(n8084), .ZN(n6011) );
  NAND2_X1 U7570 ( .A1(n6008), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6009) );
  XNOR2_X1 U7571 ( .A(n6009), .B(P2_IR_REG_18__SCAN_IN), .ZN(n6245) );
  AOI22_X1 U7572 ( .A1(n6023), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6022), .B2(
        n6245), .ZN(n6010) );
  XNOR2_X1 U7573 ( .A(n9005), .B(n6108), .ZN(n6018) );
  INV_X1 U7574 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n8577) );
  NAND2_X1 U7575 ( .A1(n6012), .A2(n8577), .ZN(n6013) );
  AND2_X1 U7576 ( .A1(n6042), .A2(n6013), .ZN(n8844) );
  NAND2_X1 U7577 ( .A1(n6093), .A2(n8844), .ZN(n6017) );
  NAND2_X1 U7578 ( .A1(n4275), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n6016) );
  NAND2_X1 U7579 ( .A1(n6148), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n6015) );
  NAND2_X1 U7580 ( .A1(n6722), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n6014) );
  NOR2_X1 U7581 ( .A1(n8832), .A2(n7043), .ZN(n6019) );
  NAND2_X1 U7582 ( .A1(n6018), .A2(n6019), .ZN(n6030) );
  INV_X1 U7583 ( .A(n6018), .ZN(n8492) );
  INV_X1 U7584 ( .A(n6019), .ZN(n6020) );
  NAND2_X1 U7585 ( .A1(n8492), .A2(n6020), .ZN(n6021) );
  AND2_X1 U7586 ( .A1(n6030), .A2(n6021), .ZN(n8572) );
  NAND2_X1 U7587 ( .A1(n7351), .A2(n8084), .ZN(n6025) );
  AOI22_X1 U7588 ( .A1(n6023), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n4284), .B2(
        n6022), .ZN(n6024) );
  XNOR2_X1 U7589 ( .A(n9002), .B(n6152), .ZN(n6034) );
  XNOR2_X1 U7590 ( .A(n6042), .B(P2_REG3_REG_19__SCAN_IN), .ZN(n8837) );
  NAND2_X1 U7591 ( .A1(n6093), .A2(n8837), .ZN(n6029) );
  NAND2_X1 U7592 ( .A1(n4275), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n6028) );
  NAND2_X1 U7593 ( .A1(n6148), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n6027) );
  NAND2_X1 U7594 ( .A1(n6722), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n6026) );
  NOR2_X1 U7595 ( .A1(n8578), .A2(n7043), .ZN(n6032) );
  XNOR2_X1 U7596 ( .A(n6034), .B(n6032), .ZN(n8493) );
  AND2_X1 U7597 ( .A1(n8493), .A2(n6030), .ZN(n6031) );
  INV_X1 U7598 ( .A(n6032), .ZN(n6033) );
  NAND2_X1 U7599 ( .A1(n6034), .A2(n6033), .ZN(n6035) );
  NAND2_X1 U7600 ( .A1(n7495), .A2(n8084), .ZN(n6037) );
  OR2_X1 U7601 ( .A1(n6082), .A2(n7497), .ZN(n6036) );
  XNOR2_X1 U7602 ( .A(n8993), .B(n6108), .ZN(n6048) );
  INV_X1 U7603 ( .A(n6042), .ZN(n6039) );
  AND2_X1 U7604 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_REG3_REG_20__SCAN_IN), 
        .ZN(n6038) );
  NAND2_X1 U7605 ( .A1(n6039), .A2(n6038), .ZN(n6056) );
  INV_X1 U7606 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n6041) );
  INV_X1 U7607 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n6040) );
  OAI21_X1 U7608 ( .B1(n6042), .B2(n6041), .A(n6040), .ZN(n6043) );
  AND2_X1 U7609 ( .A1(n6056), .A2(n6043), .ZN(n8810) );
  NAND2_X1 U7610 ( .A1(n6093), .A2(n8810), .ZN(n6047) );
  NAND2_X1 U7611 ( .A1(n4275), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n6046) );
  NAND2_X1 U7612 ( .A1(n6148), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n6045) );
  NAND2_X1 U7613 ( .A1(n6722), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n6044) );
  NOR2_X1 U7614 ( .A1(n8833), .A2(n7043), .ZN(n6049) );
  NAND2_X1 U7615 ( .A1(n6048), .A2(n6049), .ZN(n6052) );
  INV_X1 U7616 ( .A(n6048), .ZN(n8501) );
  INV_X1 U7617 ( .A(n6049), .ZN(n6050) );
  NAND2_X1 U7618 ( .A1(n8501), .A2(n6050), .ZN(n6051) );
  NAND2_X1 U7619 ( .A1(n6052), .A2(n6051), .ZN(n8553) );
  NAND2_X1 U7620 ( .A1(n7498), .A2(n8084), .ZN(n6054) );
  OR2_X1 U7621 ( .A1(n6082), .A2(n7511), .ZN(n6053) );
  XNOR2_X1 U7622 ( .A(n8988), .B(n6152), .ZN(n6073) );
  INV_X1 U7623 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n6055) );
  NAND2_X1 U7624 ( .A1(n6056), .A2(n6055), .ZN(n6057) );
  AND2_X1 U7625 ( .A1(n6066), .A2(n6057), .ZN(n8794) );
  NAND2_X1 U7626 ( .A1(n6093), .A2(n8794), .ZN(n6061) );
  NAND2_X1 U7627 ( .A1(n4275), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n6060) );
  NAND2_X1 U7628 ( .A1(n6148), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n6059) );
  NAND2_X1 U7629 ( .A1(n6722), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n6058) );
  NOR2_X1 U7630 ( .A1(n8431), .A2(n7043), .ZN(n6074) );
  XNOR2_X1 U7631 ( .A(n6073), .B(n6074), .ZN(n8499) );
  NAND2_X1 U7632 ( .A1(n7647), .A2(n8084), .ZN(n6063) );
  OR2_X1 U7633 ( .A1(n6082), .A2(n8058), .ZN(n6062) );
  XNOR2_X1 U7634 ( .A(n8983), .B(n6108), .ZN(n6077) );
  INV_X1 U7635 ( .A(n6066), .ZN(n6064) );
  NAND2_X1 U7636 ( .A1(n6064), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6090) );
  INV_X1 U7637 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n6065) );
  NAND2_X1 U7638 ( .A1(n6066), .A2(n6065), .ZN(n6067) );
  AND2_X1 U7639 ( .A1(n6090), .A2(n6067), .ZN(n8774) );
  NAND2_X1 U7640 ( .A1(n6093), .A2(n8774), .ZN(n6072) );
  NAND2_X1 U7641 ( .A1(n6068), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n6071) );
  NAND2_X1 U7642 ( .A1(n6148), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n6070) );
  NAND2_X1 U7643 ( .A1(n6722), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n6069) );
  NOR2_X1 U7644 ( .A1(n8757), .A2(n7043), .ZN(n8563) );
  INV_X1 U7645 ( .A(n6073), .ZN(n6075) );
  AND2_X1 U7646 ( .A1(n6075), .A2(n6074), .ZN(n8558) );
  AOI21_X1 U7647 ( .B1(n6077), .B2(n8563), .A(n8558), .ZN(n6076) );
  INV_X1 U7648 ( .A(n6077), .ZN(n8560) );
  INV_X1 U7649 ( .A(n8563), .ZN(n6078) );
  NAND2_X1 U7650 ( .A1(n8560), .A2(n6078), .ZN(n6079) );
  NAND2_X1 U7651 ( .A1(n7769), .A2(n8084), .ZN(n6081) );
  OR2_X1 U7652 ( .A1(n6082), .A2(n7771), .ZN(n6080) );
  XNOR2_X1 U7653 ( .A(n8975), .B(n6108), .ZN(n8537) );
  XNOR2_X1 U7654 ( .A(n6101), .B(n8537), .ZN(n8470) );
  NAND2_X1 U7655 ( .A1(n7893), .A2(n8084), .ZN(n6084) );
  OR2_X1 U7656 ( .A1(n6082), .A2(n7867), .ZN(n6083) );
  XNOR2_X1 U7657 ( .A(n8970), .B(n6152), .ZN(n6100) );
  INV_X1 U7658 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8473) );
  INV_X1 U7659 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n8546) );
  NAND2_X1 U7660 ( .A1(n6092), .A2(n8546), .ZN(n6085) );
  AND2_X1 U7661 ( .A1(n6111), .A2(n6085), .ZN(n8738) );
  NAND2_X1 U7662 ( .A1(n6093), .A2(n8738), .ZN(n6089) );
  NAND2_X1 U7663 ( .A1(n6068), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n6088) );
  NAND2_X1 U7664 ( .A1(n6721), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n6087) );
  NAND2_X1 U7665 ( .A1(n5792), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n6086) );
  NAND2_X1 U7666 ( .A1(n6090), .A2(n8473), .ZN(n6091) );
  AND2_X1 U7667 ( .A1(n6092), .A2(n6091), .ZN(n8765) );
  NAND2_X1 U7668 ( .A1(n6093), .A2(n8765), .ZN(n6097) );
  NAND2_X1 U7669 ( .A1(n6068), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n6096) );
  NAND2_X1 U7670 ( .A1(n6148), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n6095) );
  NAND2_X1 U7671 ( .A1(n6722), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n6094) );
  OR2_X1 U7672 ( .A1(n8746), .A2(n7043), .ZN(n8471) );
  AOI21_X1 U7673 ( .B1(n6100), .B2(n8756), .A(n8471), .ZN(n6099) );
  NOR2_X1 U7674 ( .A1(n8756), .A2(n7043), .ZN(n6103) );
  INV_X1 U7675 ( .A(n6103), .ZN(n8544) );
  INV_X1 U7676 ( .A(n6100), .ZN(n8541) );
  INV_X1 U7677 ( .A(n6101), .ZN(n8538) );
  AND2_X1 U7678 ( .A1(n8538), .A2(n8537), .ZN(n6102) );
  OAI21_X1 U7679 ( .B1(n8541), .B2(n6103), .A(n6102), .ZN(n6104) );
  NAND2_X1 U7680 ( .A1(n7940), .A2(n8084), .ZN(n6107) );
  OR2_X1 U7681 ( .A1(n6082), .A2(n7946), .ZN(n6106) );
  XNOR2_X1 U7682 ( .A(n8966), .B(n6108), .ZN(n8515) );
  INV_X1 U7683 ( .A(n6111), .ZN(n6109) );
  NAND2_X1 U7684 ( .A1(n6109), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6125) );
  INV_X1 U7685 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n6110) );
  NAND2_X1 U7686 ( .A1(n6111), .A2(n6110), .ZN(n6112) );
  AND2_X1 U7687 ( .A1(n6125), .A2(n6112), .ZN(n8726) );
  NAND2_X1 U7688 ( .A1(n8726), .A2(n6093), .ZN(n6116) );
  NAND2_X1 U7689 ( .A1(n6068), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n6115) );
  NAND2_X1 U7690 ( .A1(n5792), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6114) );
  NAND2_X1 U7691 ( .A1(n6148), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n6113) );
  NOR2_X1 U7692 ( .A1(n8745), .A2(n7043), .ZN(n6117) );
  AND2_X1 U7693 ( .A1(n8515), .A2(n6117), .ZN(n8512) );
  INV_X1 U7694 ( .A(n8515), .ZN(n6119) );
  INV_X1 U7695 ( .A(n6117), .ZN(n6118) );
  NAND2_X1 U7696 ( .A1(n6119), .A2(n6118), .ZN(n8517) );
  OAI21_X2 U7697 ( .B1(n8518), .B2(n8512), .A(n8517), .ZN(n8583) );
  NAND2_X1 U7698 ( .A1(n8012), .A2(n8084), .ZN(n6121) );
  XNOR2_X1 U7699 ( .A(n8961), .B(n6152), .ZN(n6131) );
  NAND2_X1 U7700 ( .A1(n5792), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6123) );
  NAND2_X1 U7701 ( .A1(n6148), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n6122) );
  AND2_X1 U7702 ( .A1(n6123), .A2(n6122), .ZN(n6129) );
  INV_X1 U7703 ( .A(n6093), .ZN(n6202) );
  INV_X1 U7704 ( .A(n6125), .ZN(n6124) );
  NAND2_X1 U7705 ( .A1(n6124), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6134) );
  INV_X1 U7706 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8584) );
  NAND2_X1 U7707 ( .A1(n6125), .A2(n8584), .ZN(n6126) );
  NAND2_X1 U7708 ( .A1(n6134), .A2(n6126), .ZN(n8717) );
  OR2_X1 U7709 ( .A1(n6202), .A2(n8717), .ZN(n6128) );
  NAND2_X1 U7710 ( .A1(n6068), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n6127) );
  INV_X1 U7711 ( .A(n8693), .ZN(n8606) );
  NAND2_X1 U7712 ( .A1(n8606), .A2(n5760), .ZN(n6130) );
  XNOR2_X1 U7713 ( .A(n6131), .B(n6130), .ZN(n8582) );
  NAND2_X1 U7714 ( .A1(n8029), .A2(n8084), .ZN(n6133) );
  XNOR2_X1 U7715 ( .A(n8957), .B(n6152), .ZN(n6139) );
  INV_X1 U7716 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n8464) );
  NAND2_X1 U7717 ( .A1(n6134), .A2(n8464), .ZN(n6135) );
  NAND2_X1 U7718 ( .A1(n8698), .A2(n6093), .ZN(n6138) );
  AOI22_X1 U7719 ( .A1(n5792), .A2(P2_REG0_REG_27__SCAN_IN), .B1(n6148), .B2(
        P2_REG2_REG_27__SCAN_IN), .ZN(n6137) );
  NAND2_X1 U7720 ( .A1(n6068), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n6136) );
  NOR2_X1 U7721 ( .A1(n8586), .A2(n7043), .ZN(n6140) );
  XNOR2_X1 U7722 ( .A(n6139), .B(n6140), .ZN(n8462) );
  INV_X1 U7723 ( .A(n6139), .ZN(n6141) );
  NAND2_X1 U7724 ( .A1(n8459), .A2(n8084), .ZN(n6143) );
  OR2_X1 U7725 ( .A1(n6082), .A2(n8461), .ZN(n6142) );
  INV_X1 U7726 ( .A(n8950), .ZN(n8679) );
  INV_X1 U7727 ( .A(n6146), .ZN(n6144) );
  NAND2_X1 U7728 ( .A1(n6144), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n8452) );
  INV_X1 U7729 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n6145) );
  NAND2_X1 U7730 ( .A1(n6146), .A2(n6145), .ZN(n6147) );
  NAND2_X1 U7731 ( .A1(n8452), .A2(n6147), .ZN(n8676) );
  OR2_X1 U7732 ( .A1(n8676), .A2(n6202), .ZN(n6151) );
  AOI22_X1 U7733 ( .A1(n5792), .A2(P2_REG0_REG_28__SCAN_IN), .B1(n6148), .B2(
        P2_REG2_REG_28__SCAN_IN), .ZN(n6150) );
  NAND2_X1 U7734 ( .A1(n6068), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6149) );
  NOR2_X1 U7735 ( .A1(n8694), .A2(n7043), .ZN(n6153) );
  XNOR2_X1 U7736 ( .A(n6153), .B(n6152), .ZN(n6193) );
  INV_X1 U7737 ( .A(n6193), .ZN(n6194) );
  NAND3_X1 U7738 ( .A1(n6161), .A2(n6164), .A3(n6166), .ZN(n6154) );
  NOR2_X1 U7739 ( .A1(n6159), .A2(n5728), .ZN(n6156) );
  MUX2_X1 U7740 ( .A(n5728), .B(n6156), .S(P2_IR_REG_25__SCAN_IN), .Z(n6157)
         );
  INV_X1 U7741 ( .A(n6157), .ZN(n6160) );
  NAND2_X1 U7742 ( .A1(n6159), .A2(n6158), .ZN(n6169) );
  NAND2_X1 U7743 ( .A1(n6187), .A2(n6164), .ZN(n6165) );
  XOR2_X1 U7744 ( .A(n6237), .B(P2_B_REG_SCAN_IN), .Z(n6168) );
  NAND2_X1 U7745 ( .A1(n6169), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6170) );
  MUX2_X1 U7746 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6170), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n6172) );
  INV_X1 U7747 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n9949) );
  NOR2_X1 U7748 ( .A1(n6186), .A2(n7943), .ZN(n9951) );
  INV_X1 U7749 ( .A(n6186), .ZN(n8017) );
  INV_X1 U7750 ( .A(n9947), .ZN(n6175) );
  INV_X1 U7751 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n9946) );
  NAND2_X1 U7752 ( .A1(n9938), .A2(n9946), .ZN(n6174) );
  NOR4_X1 U7753 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_4__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_6__SCAN_IN), .ZN(n6184) );
  INV_X1 U7754 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n9940) );
  INV_X1 U7755 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n9942) );
  INV_X1 U7756 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n9941) );
  INV_X1 U7757 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n9943) );
  NAND4_X1 U7758 ( .A1(n9940), .A2(n9942), .A3(n9941), .A4(n9943), .ZN(n6181)
         );
  NOR4_X1 U7759 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n6179) );
  NOR4_X1 U7760 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_14__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n6178) );
  NOR4_X1 U7761 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n6177) );
  NOR4_X1 U7762 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n6176) );
  NAND4_X1 U7763 ( .A1(n6179), .A2(n6178), .A3(n6177), .A4(n6176), .ZN(n6180)
         );
  NOR4_X1 U7764 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        n6181), .A4(n6180), .ZN(n6183) );
  NOR4_X1 U7765 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_8__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_10__SCAN_IN), .ZN(n6182) );
  NAND3_X1 U7766 ( .A1(n6184), .A2(n6183), .A3(n6182), .ZN(n6185) );
  NAND3_X1 U7767 ( .A1(n7515), .A2(n7514), .A3(n7517), .ZN(n6208) );
  NAND2_X1 U7768 ( .A1(n6186), .A2(n7943), .ZN(n6238) );
  INV_X1 U7769 ( .A(n9945), .ZN(n6188) );
  INV_X1 U7770 ( .A(n7496), .ZN(n8259) );
  NAND2_X1 U7771 ( .A1(n9953), .A2(n8259), .ZN(n7527) );
  INV_X1 U7772 ( .A(n7527), .ZN(n6190) );
  NAND2_X1 U7773 ( .A1(n6201), .A2(n6190), .ZN(n6191) );
  NAND2_X1 U7774 ( .A1(n9913), .A2(n4284), .ZN(n6905) );
  NOR3_X1 U7775 ( .A1(n8679), .A2(n6194), .A3(n8589), .ZN(n6192) );
  AOI21_X1 U7776 ( .B1(n8679), .B2(n6194), .A(n6192), .ZN(n6200) );
  NOR3_X1 U7777 ( .A1(n8679), .A2(n6193), .A3(n8589), .ZN(n6196) );
  NOR2_X1 U7778 ( .A1(n8950), .A2(n6194), .ZN(n6195) );
  INV_X1 U7779 ( .A(n8265), .ZN(n6911) );
  NOR2_X1 U7780 ( .A1(n9016), .A2(n6236), .ZN(n6198) );
  OAI21_X1 U7781 ( .B1(n8679), .B2(n8604), .A(n8593), .ZN(n6199) );
  OR2_X1 U7782 ( .A1(n8452), .A2(n6202), .ZN(n6205) );
  AOI22_X1 U7783 ( .A1(P2_REG1_REG_29__SCAN_IN), .A2(n6068), .B1(n5792), .B2(
        P2_REG0_REG_29__SCAN_IN), .ZN(n6204) );
  NAND2_X1 U7784 ( .A1(n6148), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n6203) );
  OR2_X1 U7785 ( .A1(n8586), .A2(n8905), .ZN(n6207) );
  OAI21_X1 U7786 ( .B1(n8081), .B2(n8907), .A(n6207), .ZN(n8682) );
  AOI22_X1 U7787 ( .A1(n8509), .A2(n8682), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3152), .ZN(n6213) );
  NAND2_X1 U7788 ( .A1(n6208), .A2(n6905), .ZN(n6211) );
  OR2_X1 U7789 ( .A1(n6912), .A2(n8265), .ZN(n7512) );
  AND2_X1 U7790 ( .A1(n6209), .A2(n7512), .ZN(n6210) );
  NAND2_X1 U7791 ( .A1(n6211), .A2(n6210), .ZN(n8418) );
  NAND2_X1 U7792 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n8628), .ZN(n6214) );
  OAI21_X1 U7793 ( .B1(n8628), .B2(P2_REG2_REG_16__SCAN_IN), .A(n6214), .ZN(
        n8633) );
  INV_X1 U7794 ( .A(n6270), .ZN(n7955) );
  XNOR2_X1 U7795 ( .A(n7240), .B(P2_REG2_REG_12__SCAN_IN), .ZN(n7232) );
  INV_X1 U7796 ( .A(n6843), .ZN(n6224) );
  INV_X1 U7797 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6215) );
  XNOR2_X1 U7798 ( .A(n6958), .B(n6215), .ZN(n6950) );
  INV_X1 U7799 ( .A(n6638), .ZN(n9521) );
  INV_X1 U7800 ( .A(n6635), .ZN(n9509) );
  INV_X1 U7801 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6216) );
  MUX2_X1 U7802 ( .A(n6216), .B(P2_REG2_REG_1__SCAN_IN), .S(n6635), .Z(n6217)
         );
  NAND2_X1 U7803 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n9507) );
  INV_X1 U7804 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6218) );
  MUX2_X1 U7805 ( .A(n6218), .B(P2_REG2_REG_2__SCAN_IN), .S(n6638), .Z(n6219)
         );
  INV_X1 U7806 ( .A(n6219), .ZN(n9519) );
  NAND2_X1 U7807 ( .A1(n6254), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6220) );
  OAI21_X1 U7808 ( .B1(n6254), .B2(P2_REG2_REG_3__SCAN_IN), .A(n6220), .ZN(
        n6998) );
  NOR2_X1 U7809 ( .A1(n6999), .A2(n6998), .ZN(n6997) );
  NOR2_X1 U7810 ( .A1(n6950), .A2(n6951), .ZN(n6949) );
  NAND2_X1 U7811 ( .A1(P2_REG2_REG_5__SCAN_IN), .A2(n6252), .ZN(n6221) );
  OAI21_X1 U7812 ( .B1(n6252), .B2(P2_REG2_REG_5__SCAN_IN), .A(n6221), .ZN(
        n6974) );
  NAND2_X1 U7813 ( .A1(P2_REG2_REG_6__SCAN_IN), .A2(n6250), .ZN(n6222) );
  OAI21_X1 U7814 ( .B1(n6250), .B2(P2_REG2_REG_6__SCAN_IN), .A(n6222), .ZN(
        n6938) );
  NAND2_X1 U7815 ( .A1(n6248), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6223) );
  OAI21_X1 U7816 ( .B1(n6248), .B2(P2_REG2_REG_7__SCAN_IN), .A(n6223), .ZN(
        n6962) );
  NOR2_X1 U7817 ( .A1(n6963), .A2(n6962), .ZN(n6961) );
  XOR2_X1 U7818 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n6843), .Z(n6836) );
  NAND2_X1 U7819 ( .A1(P2_REG2_REG_9__SCAN_IN), .A2(n6264), .ZN(n6225) );
  OAI21_X1 U7820 ( .B1(n6264), .B2(P2_REG2_REG_9__SCAN_IN), .A(n6225), .ZN(
        n6986) );
  XNOR2_X1 U7821 ( .A(n6659), .B(P2_REG2_REG_10__SCAN_IN), .ZN(n6898) );
  INV_X1 U7822 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n6226) );
  MUX2_X1 U7823 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n6226), .S(n6265), .Z(n7062)
         );
  INV_X1 U7824 ( .A(n7231), .ZN(n6227) );
  NAND2_X1 U7825 ( .A1(n7629), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n6228) );
  OAI21_X1 U7826 ( .B1(n7629), .B2(P2_REG2_REG_13__SCAN_IN), .A(n6228), .ZN(
        n7626) );
  INV_X1 U7827 ( .A(n7751), .ZN(n6685) );
  INV_X1 U7828 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n6229) );
  AOI22_X1 U7829 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n7751), .B1(n6685), .B2(
        n6229), .ZN(n7745) );
  OAI21_X1 U7830 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n7751), .A(n7744), .ZN(
        n6230) );
  NAND2_X1 U7831 ( .A1(n7955), .A2(n6230), .ZN(n6231) );
  XNOR2_X1 U7832 ( .A(n6230), .B(n6270), .ZN(n7949) );
  INV_X1 U7833 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n7948) );
  NAND2_X1 U7834 ( .A1(n7949), .A2(n7948), .ZN(n7947) );
  NAND2_X1 U7835 ( .A1(n6246), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n6232) );
  OAI21_X1 U7836 ( .B1(n6246), .B2(P2_REG2_REG_17__SCAN_IN), .A(n6232), .ZN(
        n8638) );
  INV_X1 U7837 ( .A(n6245), .ZN(n8654) );
  INV_X1 U7838 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8651) );
  NAND2_X1 U7839 ( .A1(n6233), .A2(n8654), .ZN(n6234) );
  INV_X1 U7840 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n6235) );
  INV_X1 U7841 ( .A(n6284), .ZN(n6281) );
  OR2_X1 U7842 ( .A1(n9939), .A2(n6236), .ZN(n6240) );
  OR2_X1 U7843 ( .A1(n6237), .A2(P2_U3152), .ZN(n7865) );
  NAND2_X1 U7844 ( .A1(n9945), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8270) );
  AND2_X1 U7845 ( .A1(n6241), .A2(n8270), .ZN(n6239) );
  NAND2_X1 U7846 ( .A1(n6240), .A2(n6239), .ZN(n6279) );
  NAND2_X1 U7847 ( .A1(n6279), .A2(n6286), .ZN(n6242) );
  NAND2_X1 U7848 ( .A1(n6242), .A2(n6760), .ZN(n6244) );
  NOR2_X1 U7849 ( .A1(n6206), .A2(n8264), .ZN(n6243) );
  NAND2_X1 U7850 ( .A1(n6244), .A2(n6206), .ZN(n9893) );
  INV_X1 U7851 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n6276) );
  AOI22_X1 U7852 ( .A1(n6245), .A2(n6276), .B1(P2_REG1_REG_18__SCAN_IN), .B2(
        n8654), .ZN(n8649) );
  INV_X1 U7853 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n6275) );
  INV_X1 U7854 ( .A(n6246), .ZN(n8644) );
  XNOR2_X1 U7855 ( .A(n8644), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n8641) );
  OR2_X1 U7856 ( .A1(n8628), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n6274) );
  XNOR2_X1 U7857 ( .A(n8628), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n8624) );
  INV_X1 U7858 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n9540) );
  AOI22_X1 U7859 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n6685), .B1(n7751), .B2(
        n9540), .ZN(n7743) );
  INV_X1 U7860 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n9547) );
  INV_X1 U7861 ( .A(n7629), .ZN(n6681) );
  INV_X1 U7862 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n10043) );
  MUX2_X1 U7863 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n10043), .S(n7240), .Z(n7235) );
  INV_X1 U7864 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n10040) );
  INV_X1 U7865 ( .A(n6265), .ZN(n7066) );
  INV_X1 U7866 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n10038) );
  MUX2_X1 U7867 ( .A(n10038), .B(P2_REG1_REG_10__SCAN_IN), .S(n6659), .Z(n6895) );
  INV_X1 U7868 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6247) );
  MUX2_X1 U7869 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n6247), .S(n6264), .Z(n6990)
         );
  INV_X1 U7870 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6262) );
  NAND2_X1 U7871 ( .A1(n6248), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6260) );
  INV_X1 U7872 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6249) );
  MUX2_X1 U7873 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n6249), .S(n6248), .Z(n6966)
         );
  NAND2_X1 U7874 ( .A1(P2_REG1_REG_6__SCAN_IN), .A2(n6250), .ZN(n6259) );
  INV_X1 U7875 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6251) );
  MUX2_X1 U7876 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n6251), .S(n6250), .Z(n6942)
         );
  NAND2_X1 U7877 ( .A1(P2_REG1_REG_5__SCAN_IN), .A2(n6252), .ZN(n6258) );
  INV_X1 U7878 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6253) );
  MUX2_X1 U7879 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n6253), .S(n6252), .Z(n6979)
         );
  INV_X1 U7880 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6257) );
  NAND2_X1 U7881 ( .A1(n6254), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6256) );
  INV_X1 U7882 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6255) );
  MUX2_X1 U7883 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n6255), .S(n6254), .Z(n7003)
         );
  INV_X1 U7884 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10031) );
  MUX2_X1 U7885 ( .A(n10031), .B(P2_REG1_REG_2__SCAN_IN), .S(n6638), .Z(n9524)
         );
  INV_X1 U7886 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6936) );
  MUX2_X1 U7887 ( .A(n6936), .B(P2_REG1_REG_1__SCAN_IN), .S(n6635), .Z(n9512)
         );
  NAND3_X1 U7888 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .A3(n9512), .ZN(n9511) );
  OAI21_X1 U7889 ( .B1(n6635), .B2(n6936), .A(n9511), .ZN(n9525) );
  NAND2_X1 U7890 ( .A1(n9524), .A2(n9525), .ZN(n9523) );
  OAI21_X1 U7891 ( .B1(n6638), .B2(n10031), .A(n9523), .ZN(n7002) );
  NAND2_X1 U7892 ( .A1(n7003), .A2(n7002), .ZN(n7001) );
  NAND2_X1 U7893 ( .A1(n6256), .A2(n7001), .ZN(n6955) );
  MUX2_X1 U7894 ( .A(n6257), .B(P2_REG1_REG_4__SCAN_IN), .S(n6958), .Z(n6954)
         );
  NAND2_X1 U7895 ( .A1(n6955), .A2(n6954), .ZN(n6953) );
  OAI21_X1 U7896 ( .B1(n6958), .B2(n6257), .A(n6953), .ZN(n6978) );
  NAND2_X1 U7897 ( .A1(n6979), .A2(n6978), .ZN(n6977) );
  NAND2_X1 U7898 ( .A1(n6258), .A2(n6977), .ZN(n6943) );
  NAND2_X1 U7899 ( .A1(n6942), .A2(n6943), .ZN(n6941) );
  NAND2_X1 U7900 ( .A1(n6259), .A2(n6941), .ZN(n6967) );
  NAND2_X1 U7901 ( .A1(n6966), .A2(n6967), .ZN(n6965) );
  AND2_X1 U7902 ( .A1(n6260), .A2(n6965), .ZN(n6834) );
  MUX2_X1 U7903 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n6262), .S(n6843), .Z(n6833)
         );
  NOR2_X1 U7904 ( .A1(n6834), .A2(n6833), .ZN(n6832) );
  INV_X1 U7905 ( .A(n6832), .ZN(n6261) );
  OAI21_X1 U7906 ( .B1(n6262), .B2(n6843), .A(n6261), .ZN(n6991) );
  NAND2_X1 U7907 ( .A1(n6990), .A2(n6991), .ZN(n6989) );
  INV_X1 U7908 ( .A(n6989), .ZN(n6263) );
  AOI21_X1 U7909 ( .B1(n6264), .B2(P2_REG1_REG_9__SCAN_IN), .A(n6263), .ZN(
        n6896) );
  NOR2_X1 U7910 ( .A1(n6895), .A2(n6896), .ZN(n6894) );
  AOI21_X1 U7911 ( .B1(n6659), .B2(P2_REG1_REG_10__SCAN_IN), .A(n6894), .ZN(
        n7057) );
  MUX2_X1 U7912 ( .A(n10040), .B(P2_REG1_REG_11__SCAN_IN), .S(n6265), .Z(n7056) );
  OR2_X1 U7913 ( .A1(n7057), .A2(n7056), .ZN(n6266) );
  OAI21_X1 U7914 ( .B1(n10040), .B2(n7066), .A(n6266), .ZN(n6267) );
  INV_X1 U7915 ( .A(n6267), .ZN(n7234) );
  NAND2_X1 U7916 ( .A1(n7235), .A2(n7234), .ZN(n7233) );
  INV_X1 U7917 ( .A(n7240), .ZN(n6676) );
  NAND2_X1 U7918 ( .A1(n6676), .A2(n10043), .ZN(n6268) );
  NAND2_X1 U7919 ( .A1(n7233), .A2(n6268), .ZN(n7628) );
  MUX2_X1 U7920 ( .A(n9547), .B(P2_REG1_REG_13__SCAN_IN), .S(n7629), .Z(n7627)
         );
  OR2_X1 U7921 ( .A1(n7628), .A2(n7627), .ZN(n6269) );
  OAI21_X1 U7922 ( .B1(n9547), .B2(n6681), .A(n6269), .ZN(n7742) );
  NOR2_X1 U7923 ( .A1(n7743), .A2(n7742), .ZN(n7741) );
  AOI21_X1 U7924 ( .B1(n9540), .B2(n6685), .A(n7741), .ZN(n6271) );
  NAND2_X1 U7925 ( .A1(n6270), .A2(n6271), .ZN(n6272) );
  XNOR2_X1 U7926 ( .A(n6271), .B(n7955), .ZN(n7951) );
  NAND2_X1 U7927 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n7951), .ZN(n7950) );
  NAND2_X1 U7928 ( .A1(n6272), .A2(n7950), .ZN(n8625) );
  NOR2_X1 U7929 ( .A1(n8624), .A2(n8625), .ZN(n8623) );
  INV_X1 U7930 ( .A(n8623), .ZN(n6273) );
  NAND2_X1 U7931 ( .A1(n8641), .A2(n4846), .ZN(n8640) );
  OAI21_X1 U7932 ( .B1(n6275), .B2(n8644), .A(n8640), .ZN(n8648) );
  NOR2_X1 U7933 ( .A1(n8649), .A2(n8648), .ZN(n8647) );
  AOI21_X1 U7934 ( .B1(n8654), .B2(n6276), .A(n8647), .ZN(n6277) );
  XNOR2_X1 U7935 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n6277), .ZN(n6283) );
  AND2_X1 U7936 ( .A1(n6286), .A2(n8264), .ZN(n6278) );
  NAND2_X1 U7937 ( .A1(n6283), .A2(n9888), .ZN(n6280) );
  OAI211_X1 U7938 ( .C1(n6281), .C2(n9895), .A(n9893), .B(n6280), .ZN(n6282)
         );
  NAND2_X1 U7939 ( .A1(n6282), .A2(n4284), .ZN(n6294) );
  OAI22_X1 U7940 ( .A1(n6284), .A2(n9895), .B1(n6283), .B2(n9894), .ZN(n6292)
         );
  OR2_X1 U7941 ( .A1(n8270), .A2(n6286), .ZN(n6285) );
  NAND2_X1 U7942 ( .A1(n9939), .A2(n6285), .ZN(n6288) );
  NAND2_X1 U7943 ( .A1(n6912), .A2(n6286), .ZN(n6287) );
  NAND2_X1 U7944 ( .A1(n6288), .A2(n6287), .ZN(n7749) );
  NAND2_X1 U7945 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_U3152), .ZN(n6289) );
  INV_X2 U7946 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  INV_X1 U7947 ( .A(n6430), .ZN(n6418) );
  NAND2_X1 U7948 ( .A1(n9229), .A2(n6418), .ZN(n6424) );
  NOR2_X1 U7949 ( .A1(n9429), .A2(n9179), .ZN(n9192) );
  INV_X1 U7950 ( .A(n9192), .ZN(n6295) );
  INV_X1 U7951 ( .A(n9283), .ZN(n9316) );
  OR2_X1 U7952 ( .A1(n9423), .A2(n9316), .ZN(n6494) );
  AND2_X1 U7953 ( .A1(n6295), .A2(n6494), .ZN(n6469) );
  INV_X1 U7954 ( .A(n6469), .ZN(n6296) );
  NAND2_X1 U7955 ( .A1(n9423), .A2(n9316), .ZN(n9193) );
  AND2_X1 U7956 ( .A1(n6296), .A2(n9193), .ZN(n6297) );
  NOR2_X1 U7957 ( .A1(n9194), .A2(n6297), .ZN(n6300) );
  NAND2_X1 U7958 ( .A1(n9429), .A2(n9179), .ZN(n6298) );
  NAND2_X1 U7959 ( .A1(n9193), .A2(n6298), .ZN(n6364) );
  AND2_X1 U7960 ( .A1(n6364), .A2(n6494), .ZN(n6299) );
  NOR2_X1 U7961 ( .A1(n9196), .A2(n6299), .ZN(n6475) );
  MUX2_X1 U7962 ( .A(n6300), .B(n6475), .S(n6418), .Z(n6367) );
  NAND2_X1 U7963 ( .A1(n9453), .A2(n9083), .ZN(n9185) );
  NAND2_X1 U7964 ( .A1(n9458), .A2(n8037), .ZN(n6302) );
  AND2_X1 U7965 ( .A1(n9185), .A2(n6302), .ZN(n6459) );
  OR2_X1 U7966 ( .A1(n9453), .A2(n9083), .ZN(n6497) );
  NAND2_X1 U7967 ( .A1(n6497), .A2(n8032), .ZN(n6467) );
  INV_X1 U7968 ( .A(n6467), .ZN(n6301) );
  MUX2_X1 U7969 ( .A(n6459), .B(n6301), .S(n6430), .Z(n6349) );
  NAND2_X1 U7970 ( .A1(n8032), .A2(n6302), .ZN(n7980) );
  INV_X1 U7971 ( .A(n7980), .ZN(n7973) );
  OR2_X1 U7972 ( .A1(n9465), .A2(n7982), .ZN(n6457) );
  NAND2_X1 U7973 ( .A1(n9465), .A2(n7982), .ZN(n6460) );
  MUX2_X1 U7974 ( .A(n6457), .B(n6460), .S(n6430), .Z(n6347) );
  INV_X1 U7975 ( .A(n7969), .ZN(n6345) );
  NAND2_X1 U7976 ( .A1(n7912), .A2(n7913), .ZN(n7920) );
  AND2_X1 U7977 ( .A1(n9588), .A2(n9152), .ZN(n7836) );
  OR2_X1 U7978 ( .A1(n7823), .A2(n9561), .ZN(n6500) );
  INV_X1 U7979 ( .A(n6500), .ZN(n6303) );
  OR2_X1 U7980 ( .A1(n7836), .A2(n6303), .ZN(n6304) );
  NAND2_X1 U7981 ( .A1(n7877), .A2(n7963), .ZN(n6334) );
  NAND2_X1 U7982 ( .A1(n6304), .A2(n6334), .ZN(n6342) );
  AND2_X1 U7983 ( .A1(n7176), .A2(n5092), .ZN(n7022) );
  NAND2_X1 U7984 ( .A1(n7034), .A2(n6693), .ZN(n6306) );
  NAND2_X1 U7985 ( .A1(n7021), .A2(n6306), .ZN(n7247) );
  NAND2_X1 U7986 ( .A1(n7255), .A2(n9161), .ZN(n6524) );
  NAND2_X1 U7987 ( .A1(n7247), .A2(n7248), .ZN(n7246) );
  NAND2_X1 U7988 ( .A1(n9823), .A2(n9160), .ZN(n6438) );
  NAND2_X1 U7989 ( .A1(n6438), .A2(n6441), .ZN(n7112) );
  INV_X1 U7990 ( .A(n7112), .ZN(n7288) );
  NAND2_X1 U7991 ( .A1(n7116), .A2(n9767), .ZN(n9761) );
  INV_X1 U7992 ( .A(n9761), .ZN(n9758) );
  NAND2_X1 U7993 ( .A1(n9836), .A2(n9733), .ZN(n7119) );
  NAND2_X1 U7994 ( .A1(n9829), .A2(n9159), .ZN(n7115) );
  NAND2_X1 U7995 ( .A1(n7119), .A2(n7115), .ZN(n6442) );
  INV_X1 U7996 ( .A(n6442), .ZN(n6308) );
  NAND2_X1 U7997 ( .A1(n9752), .A2(n9782), .ZN(n7118) );
  NAND2_X1 U7998 ( .A1(n9779), .A2(n7115), .ZN(n9763) );
  AND2_X1 U7999 ( .A1(n7118), .A2(n9761), .ZN(n6533) );
  INV_X1 U8000 ( .A(n7119), .ZN(n6309) );
  AOI21_X1 U8001 ( .B1(n9763), .B2(n6533), .A(n6309), .ZN(n6310) );
  MUX2_X1 U8002 ( .A(n9737), .B(n6310), .S(n6430), .Z(n6311) );
  NAND2_X1 U8003 ( .A1(n9841), .A2(n9158), .ZN(n6440) );
  NAND2_X1 U8004 ( .A1(n7284), .A2(n5181), .ZN(n6530) );
  NAND2_X1 U8005 ( .A1(n6311), .A2(n9738), .ZN(n6323) );
  NAND2_X1 U8006 ( .A1(n9849), .A2(n9735), .ZN(n6526) );
  AND2_X1 U8007 ( .A1(n6526), .A2(n6440), .ZN(n6313) );
  NAND2_X1 U8008 ( .A1(n6314), .A2(n8315), .ZN(n7165) );
  AND2_X1 U8009 ( .A1(n7163), .A2(n7165), .ZN(n6448) );
  INV_X1 U8010 ( .A(n6448), .ZN(n6312) );
  AOI21_X1 U8011 ( .B1(n6323), .B2(n6313), .A(n6312), .ZN(n6318) );
  OR2_X1 U8012 ( .A1(n7503), .A2(n7490), .ZN(n6315) );
  OR2_X1 U8013 ( .A1(n7334), .A2(n7207), .ZN(n7202) );
  AND2_X1 U8014 ( .A1(n6315), .A2(n7202), .ZN(n7167) );
  AND2_X1 U8015 ( .A1(n6503), .A2(n7167), .ZN(n6456) );
  INV_X1 U8016 ( .A(n6456), .ZN(n6317) );
  NAND2_X1 U8017 ( .A1(n7503), .A2(n7490), .ZN(n6326) );
  NAND2_X1 U8018 ( .A1(n7334), .A2(n7207), .ZN(n7201) );
  NAND2_X1 U8019 ( .A1(n6326), .A2(n7201), .ZN(n6316) );
  NAND2_X1 U8020 ( .A1(n6316), .A2(n6315), .ZN(n7168) );
  OAI21_X1 U8021 ( .B1(n6318), .B2(n6317), .A(n7168), .ZN(n6321) );
  NOR2_X1 U8022 ( .A1(n9470), .A2(n9559), .ZN(n7546) );
  NAND2_X1 U8023 ( .A1(n9470), .A2(n9559), .ZN(n7547) );
  INV_X1 U8024 ( .A(n7547), .ZN(n6319) );
  OR2_X1 U8025 ( .A1(n7546), .A2(n6319), .ZN(n7170) );
  OR2_X1 U8026 ( .A1(n9571), .A2(n7674), .ZN(n7553) );
  NAND2_X1 U8027 ( .A1(n7170), .A2(n7553), .ZN(n6328) );
  NOR2_X1 U8028 ( .A1(n6328), .A2(n6430), .ZN(n6320) );
  OR2_X1 U8029 ( .A1(n7912), .A2(n7913), .ZN(n6499) );
  INV_X1 U8030 ( .A(n6499), .ZN(n6451) );
  NAND2_X1 U8031 ( .A1(n6451), .A2(n6430), .ZN(n6322) );
  NAND3_X1 U8032 ( .A1(n6323), .A2(n7163), .A3(n6530), .ZN(n6324) );
  NAND3_X1 U8033 ( .A1(n6324), .A2(n6503), .A3(n6526), .ZN(n6325) );
  NAND3_X1 U8034 ( .A1(n6325), .A2(n7165), .A3(n7201), .ZN(n6330) );
  NAND2_X1 U8035 ( .A1(n9571), .A2(n7674), .ZN(n7554) );
  NAND3_X1 U8036 ( .A1(n7554), .A2(n6430), .A3(n6326), .ZN(n6327) );
  OR2_X1 U8037 ( .A1(n6328), .A2(n6327), .ZN(n6329) );
  AOI21_X1 U8038 ( .B1(n6330), .B2(n7167), .A(n6329), .ZN(n6338) );
  OR2_X1 U8039 ( .A1(n9470), .A2(n7655), .ZN(n7550) );
  NAND2_X1 U8040 ( .A1(n7553), .A2(n7550), .ZN(n6331) );
  NAND2_X1 U8041 ( .A1(n6331), .A2(n7554), .ZN(n6332) );
  NAND2_X1 U8042 ( .A1(n6500), .A2(n6332), .ZN(n6452) );
  OAI21_X1 U8043 ( .B1(n7836), .B2(n6452), .A(n6430), .ZN(n6333) );
  INV_X1 U8044 ( .A(n6333), .ZN(n6337) );
  NAND2_X1 U8045 ( .A1(n7823), .A2(n9561), .ZN(n7825) );
  NAND2_X1 U8046 ( .A1(n6334), .A2(n7825), .ZN(n6447) );
  INV_X1 U8047 ( .A(n6447), .ZN(n6453) );
  OR2_X1 U8048 ( .A1(n6453), .A2(n7836), .ZN(n6335) );
  AND2_X1 U8049 ( .A1(n6335), .A2(n7920), .ZN(n6336) );
  OAI21_X1 U8050 ( .B1(n6338), .B2(n6337), .A(n6336), .ZN(n6344) );
  AND2_X1 U8051 ( .A1(n9470), .A2(n7655), .ZN(n7551) );
  INV_X1 U8052 ( .A(n7551), .ZN(n6339) );
  NAND2_X1 U8053 ( .A1(n7554), .A2(n6339), .ZN(n6445) );
  AND2_X1 U8054 ( .A1(n6445), .A2(n7553), .ZN(n6340) );
  OR2_X1 U8055 ( .A1(n6447), .A2(n6340), .ZN(n6341) );
  NAND4_X1 U8056 ( .A1(n6342), .A2(n6418), .A3(n6341), .A4(n6499), .ZN(n6343)
         );
  NAND3_X1 U8057 ( .A1(n7973), .A2(n6347), .A3(n6346), .ZN(n6348) );
  NAND2_X1 U8058 ( .A1(n6349), .A2(n6348), .ZN(n6351) );
  INV_X1 U8059 ( .A(n9174), .ZN(n9362) );
  OR2_X1 U8060 ( .A1(n9447), .A2(n9362), .ZN(n6498) );
  NAND3_X1 U8061 ( .A1(n6351), .A2(n6497), .A3(n6498), .ZN(n6350) );
  NAND2_X1 U8062 ( .A1(n9447), .A2(n9362), .ZN(n9187) );
  INV_X1 U8063 ( .A(n9381), .ZN(n9177) );
  NAND2_X1 U8064 ( .A1(n9442), .A2(n9177), .ZN(n6496) );
  NAND3_X1 U8065 ( .A1(n6350), .A2(n9187), .A3(n6496), .ZN(n6355) );
  NAND2_X1 U8066 ( .A1(n9342), .A2(n6498), .ZN(n6466) );
  INV_X1 U8067 ( .A(n6466), .ZN(n6353) );
  AND2_X1 U8068 ( .A1(n9187), .A2(n9185), .ZN(n6468) );
  NAND2_X1 U8069 ( .A1(n6351), .A2(n6468), .ZN(n6352) );
  NAND2_X1 U8070 ( .A1(n6353), .A2(n6352), .ZN(n6354) );
  MUX2_X1 U8071 ( .A(n6355), .B(n6354), .S(n6430), .Z(n6362) );
  NAND2_X1 U8072 ( .A1(n9438), .A2(n9363), .ZN(n9189) );
  INV_X1 U8073 ( .A(n9189), .ZN(n6356) );
  AOI21_X1 U8074 ( .B1(n6362), .B2(n9342), .A(n6356), .ZN(n6357) );
  OR2_X1 U8075 ( .A1(n9432), .A2(n9315), .ZN(n9191) );
  OR2_X1 U8076 ( .A1(n9438), .A2(n9363), .ZN(n6495) );
  NAND2_X1 U8077 ( .A1(n9191), .A2(n6495), .ZN(n6465) );
  AND2_X1 U8078 ( .A1(n9432), .A2(n9315), .ZN(n9190) );
  OAI21_X1 U8079 ( .B1(n6357), .B2(n6465), .A(n4674), .ZN(n6366) );
  INV_X1 U8080 ( .A(n6496), .ZN(n6358) );
  NAND2_X1 U8081 ( .A1(n6495), .A2(n6358), .ZN(n6359) );
  NAND2_X1 U8082 ( .A1(n6359), .A2(n9189), .ZN(n6360) );
  OR2_X1 U8083 ( .A1(n9190), .A2(n6360), .ZN(n6436) );
  AND2_X1 U8084 ( .A1(n6436), .A2(n9191), .ZN(n6470) );
  INV_X1 U8085 ( .A(n6470), .ZN(n6361) );
  OAI21_X1 U8086 ( .B1(n6465), .B2(n6362), .A(n6361), .ZN(n6363) );
  NOR2_X1 U8087 ( .A1(n6364), .A2(n6363), .ZN(n6365) );
  INV_X1 U8088 ( .A(n9196), .ZN(n6368) );
  NAND2_X1 U8089 ( .A1(n6369), .A2(n6472), .ZN(n6372) );
  NAND2_X1 U8090 ( .A1(n9412), .A2(n6472), .ZN(n6493) );
  OAI21_X1 U8091 ( .B1(n9194), .B2(n9284), .A(n6493), .ZN(n6370) );
  MUX2_X1 U8092 ( .A(n9262), .B(n6370), .S(n6418), .Z(n6371) );
  NAND2_X1 U8093 ( .A1(n6372), .A2(n6371), .ZN(n6378) );
  NAND2_X1 U8094 ( .A1(n9248), .A2(n9267), .ZN(n6479) );
  NAND2_X1 U8095 ( .A1(n9199), .A2(n6479), .ZN(n9238) );
  OAI21_X1 U8096 ( .B1(n9262), .B2(n9194), .A(n6479), .ZN(n6374) );
  OAI21_X1 U8097 ( .B1(n6472), .B2(n9196), .A(n9199), .ZN(n6373) );
  OAI21_X1 U8098 ( .B1(n6376), .B2(n9238), .A(n6375), .ZN(n6377) );
  NAND2_X1 U8099 ( .A1(n6378), .A2(n6377), .ZN(n6380) );
  NAND2_X1 U8100 ( .A1(n9401), .A2(n9245), .ZN(n9203) );
  MUX2_X1 U8101 ( .A(n9199), .B(n6479), .S(n6430), .Z(n6379) );
  NAND3_X1 U8102 ( .A1(n6380), .A2(n9227), .A3(n6379), .ZN(n6382) );
  MUX2_X1 U8103 ( .A(n9203), .B(n9200), .S(n6430), .Z(n6381) );
  INV_X1 U8104 ( .A(n6426), .ZN(n6423) );
  INV_X1 U8105 ( .A(n9229), .ZN(n6480) );
  NAND2_X1 U8106 ( .A1(n6423), .A2(n6480), .ZN(n6390) );
  INV_X1 U8107 ( .A(SI_28_), .ZN(n6385) );
  INV_X1 U8108 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n9048) );
  INV_X1 U8109 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n9501) );
  MUX2_X1 U8110 ( .A(n9048), .B(n9501), .S(n4283), .Z(n6392) );
  XNOR2_X1 U8111 ( .A(n6392), .B(SI_29_), .ZN(n6387) );
  NAND2_X1 U8112 ( .A1(n9046), .A2(n6416), .ZN(n6389) );
  NAND2_X1 U8113 ( .A1(n5213), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n6388) );
  OR2_X2 U8114 ( .A1(n6390), .A2(n9398), .ZN(n6421) );
  INV_X1 U8115 ( .A(SI_29_), .ZN(n6391) );
  AND2_X1 U8116 ( .A1(n6392), .A2(n6391), .ZN(n6395) );
  INV_X1 U8117 ( .A(n6392), .ZN(n6393) );
  NAND2_X1 U8118 ( .A1(n6393), .A2(SI_29_), .ZN(n6394) );
  MUX2_X1 U8119 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .S(n4278), .Z(n6408) );
  NAND2_X1 U8120 ( .A1(n8060), .A2(n6416), .ZN(n6398) );
  INV_X1 U8121 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8387) );
  OR2_X1 U8122 ( .A1(n6414), .A2(n8387), .ZN(n6397) );
  INV_X1 U8123 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n6401) );
  NAND2_X1 U8124 ( .A1(n4289), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n6400) );
  NAND2_X1 U8125 ( .A1(n5446), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n6399) );
  OAI211_X1 U8126 ( .C1(n5111), .C2(n6401), .A(n6400), .B(n6399), .ZN(n9206)
         );
  INV_X1 U8127 ( .A(n9206), .ZN(n6489) );
  OR2_X1 U8128 ( .A1(n9169), .A2(n6489), .ZN(n6492) );
  INV_X1 U8129 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n6405) );
  NAND2_X1 U8130 ( .A1(n4289), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6404) );
  INV_X1 U8131 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n6402) );
  OR2_X1 U8132 ( .A1(n5241), .A2(n6402), .ZN(n6403) );
  OAI211_X1 U8133 ( .C1(n5111), .C2(n6405), .A(n6404), .B(n6403), .ZN(n9165)
         );
  NAND2_X1 U8134 ( .A1(n6492), .A2(n9165), .ZN(n6417) );
  INV_X1 U8135 ( .A(SI_30_), .ZN(n6406) );
  NAND2_X1 U8136 ( .A1(n6409), .A2(n6408), .ZN(n6410) );
  MUX2_X1 U8137 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n4283), .Z(n6411) );
  XNOR2_X1 U8138 ( .A(n6411), .B(SI_31_), .ZN(n6412) );
  INV_X1 U8139 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n6413) );
  NOR2_X1 U8140 ( .A1(n6414), .A2(n6413), .ZN(n6415) );
  OAI21_X1 U8141 ( .B1(n6424), .B2(n6423), .A(n6422), .ZN(n6433) );
  NAND2_X1 U8142 ( .A1(n9206), .A2(n9165), .ZN(n6425) );
  NAND2_X1 U8143 ( .A1(n9169), .A2(n6425), .ZN(n6483) );
  NAND3_X1 U8144 ( .A1(n6487), .A2(n6426), .A3(n9398), .ZN(n6427) );
  NAND2_X1 U8145 ( .A1(n6427), .A2(n6483), .ZN(n6429) );
  INV_X1 U8146 ( .A(n9165), .ZN(n6428) );
  INV_X1 U8147 ( .A(n6517), .ZN(n6546) );
  NAND2_X1 U8148 ( .A1(n6429), .A2(n6546), .ZN(n6431) );
  MUX2_X1 U8149 ( .A(n6487), .B(n6431), .S(n6430), .Z(n6432) );
  AND2_X1 U8150 ( .A1(n6434), .A2(n9165), .ZN(n6556) );
  NAND2_X1 U8151 ( .A1(n6705), .A2(n5660), .ZN(n7019) );
  OR2_X1 U8152 ( .A1(n9398), .A2(n6480), .ZN(n6435) );
  AND2_X1 U8153 ( .A1(n6435), .A2(n9200), .ZN(n6542) );
  INV_X1 U8154 ( .A(n6542), .ZN(n6485) );
  INV_X1 U8155 ( .A(n6436), .ZN(n6437) );
  NAND2_X1 U8156 ( .A1(n6475), .A2(n6437), .ZN(n6536) );
  AND2_X1 U8157 ( .A1(n6440), .A2(n7119), .ZN(n6529) );
  AND2_X1 U8158 ( .A1(n7115), .A2(n6438), .ZN(n6439) );
  NAND2_X1 U8159 ( .A1(n6529), .A2(n6439), .ZN(n6531) );
  INV_X1 U8160 ( .A(n6440), .ZN(n6444) );
  NAND3_X1 U8161 ( .A1(n6533), .A2(n6530), .A3(n6441), .ZN(n7098) );
  NAND3_X1 U8162 ( .A1(n6442), .A2(n6530), .A3(n7118), .ZN(n6443) );
  NAND2_X1 U8163 ( .A1(n7098), .A2(n6443), .ZN(n6504) );
  OAI22_X1 U8164 ( .A1(n4656), .A2(n6531), .B1(n6444), .B2(n6504), .ZN(n6449)
         );
  AND2_X1 U8165 ( .A1(n6460), .A2(n7920), .ZN(n7978) );
  INV_X1 U8166 ( .A(n7168), .ZN(n6446) );
  NOR3_X1 U8167 ( .A1(n6447), .A2(n6446), .A3(n6445), .ZN(n6450) );
  NAND4_X1 U8168 ( .A1(n6459), .A2(n7978), .A3(n6448), .A4(n6450), .ZN(n6534)
         );
  AOI21_X1 U8169 ( .B1(n6526), .B2(n6449), .A(n6534), .ZN(n6464) );
  INV_X1 U8170 ( .A(n6450), .ZN(n6455) );
  AOI211_X1 U8171 ( .C1(n6453), .C2(n6452), .A(n7836), .B(n6451), .ZN(n6454)
         );
  OAI21_X1 U8172 ( .B1(n6456), .B2(n6455), .A(n6454), .ZN(n6458) );
  INV_X1 U8173 ( .A(n6457), .ZN(n7977) );
  AOI21_X1 U8174 ( .B1(n6458), .B2(n7920), .A(n7977), .ZN(n6463) );
  INV_X1 U8175 ( .A(n6459), .ZN(n6462) );
  INV_X1 U8176 ( .A(n6460), .ZN(n6461) );
  NOR3_X1 U8177 ( .A1(n6463), .A2(n6462), .A3(n6461), .ZN(n6538) );
  OAI21_X1 U8178 ( .B1(n6464), .B2(n6538), .A(n9187), .ZN(n6476) );
  AOI211_X1 U8179 ( .C1(n6468), .C2(n6467), .A(n6466), .B(n6465), .ZN(n6471)
         );
  OAI21_X1 U8180 ( .B1(n6471), .B2(n6470), .A(n6469), .ZN(n6474) );
  INV_X1 U8181 ( .A(n9198), .ZN(n6473) );
  AOI211_X1 U8182 ( .C1(n6475), .C2(n6474), .A(n9194), .B(n6473), .ZN(n6541)
         );
  OAI211_X1 U8183 ( .C1(n6536), .C2(n6476), .A(n6541), .B(n9199), .ZN(n6484)
         );
  INV_X1 U8184 ( .A(n6493), .ZN(n6477) );
  NAND2_X1 U8185 ( .A1(n9199), .A2(n6477), .ZN(n6478) );
  NAND3_X1 U8186 ( .A1(n9203), .A2(n6479), .A3(n6478), .ZN(n6482) );
  AND2_X1 U8187 ( .A1(n9398), .A2(n6480), .ZN(n6481) );
  AOI21_X1 U8188 ( .B1(n6542), .B2(n6482), .A(n6481), .ZN(n6545) );
  OAI211_X1 U8189 ( .C1(n6485), .C2(n6484), .A(n6483), .B(n6545), .ZN(n6486)
         );
  AOI211_X1 U8190 ( .C1(n6487), .C2(n6486), .A(n7499), .B(n6556), .ZN(n6488)
         );
  NOR3_X1 U8191 ( .A1(n6488), .A2(n9757), .A3(n5658), .ZN(n6520) );
  AND2_X1 U8192 ( .A1(n5660), .A2(n9757), .ZN(n6554) );
  INV_X1 U8193 ( .A(n6556), .ZN(n6491) );
  NAND2_X1 U8194 ( .A1(n9169), .A2(n6489), .ZN(n6490) );
  NAND2_X1 U8195 ( .A1(n6491), .A2(n6490), .ZN(n6547) );
  INV_X1 U8196 ( .A(n6492), .ZN(n6543) );
  XNOR2_X1 U8197 ( .A(n9398), .B(n9229), .ZN(n9204) );
  INV_X1 U8198 ( .A(n9281), .ZN(n9274) );
  NAND2_X1 U8199 ( .A1(n9198), .A2(n6493), .ZN(n9264) );
  NAND2_X1 U8200 ( .A1(n6495), .A2(n9189), .ZN(n9335) );
  NAND2_X1 U8201 ( .A1(n7553), .A2(n7554), .ZN(n9557) );
  INV_X1 U8202 ( .A(n7022), .ZN(n6501) );
  INV_X1 U8203 ( .A(n7176), .ZN(n7031) );
  NAND2_X1 U8204 ( .A1(n7031), .A2(n7011), .ZN(n6521) );
  AND2_X1 U8205 ( .A1(n6501), .A2(n6521), .ZN(n6711) );
  NAND3_X1 U8206 ( .A1(n6711), .A2(n7023), .A3(n7248), .ZN(n6502) );
  NOR2_X1 U8207 ( .A1(n6502), .A2(n6531), .ZN(n6505) );
  NAND2_X1 U8208 ( .A1(n6526), .A2(n7163), .ZN(n7123) );
  INV_X1 U8209 ( .A(n7123), .ZN(n7148) );
  NAND4_X1 U8210 ( .A1(n6505), .A2(n7148), .A3(n7194), .A4(n6504), .ZN(n6506)
         );
  NAND2_X1 U8211 ( .A1(n7202), .A2(n7201), .ZN(n7323) );
  NOR2_X1 U8212 ( .A1(n6506), .A2(n7323), .ZN(n6507) );
  XNOR2_X1 U8213 ( .A(n7503), .B(n9155), .ZN(n7204) );
  NAND3_X1 U8214 ( .A1(n7170), .A2(n6507), .A3(n7204), .ZN(n6508) );
  NOR2_X1 U8215 ( .A1(n9557), .A2(n6508), .ZN(n6509) );
  XNOR2_X1 U8216 ( .A(n7877), .B(n9152), .ZN(n7837) );
  NAND4_X1 U8217 ( .A1(n7842), .A2(n7556), .A3(n6509), .A4(n7837), .ZN(n6510)
         );
  NOR3_X1 U8218 ( .A1(n7980), .A2(n7969), .A3(n6510), .ZN(n6511) );
  NAND4_X1 U8219 ( .A1(n9359), .A2(n8041), .A3(n9378), .A4(n6511), .ZN(n6512)
         );
  NOR2_X1 U8220 ( .A1(n9335), .A2(n6512), .ZN(n6513) );
  XNOR2_X1 U8221 ( .A(n9429), .B(n9329), .ZN(n9312) );
  NAND4_X1 U8222 ( .A1(n9291), .A2(n9326), .A3(n6513), .A4(n9312), .ZN(n6514)
         );
  NOR4_X1 U8223 ( .A1(n9238), .A2(n9274), .A3(n9264), .A4(n6514), .ZN(n6515)
         );
  NAND3_X1 U8224 ( .A1(n9204), .A2(n6515), .A3(n9227), .ZN(n6516) );
  NOR2_X1 U8225 ( .A1(n6518), .A2(n6705), .ZN(n6519) );
  MUX2_X1 U8226 ( .A(n6520), .B(n6554), .S(n6519), .Z(n6552) );
  INV_X1 U8227 ( .A(n9238), .ZN(n9241) );
  OAI211_X1 U8228 ( .C1(n6693), .C2(n7034), .A(n6521), .B(n6705), .ZN(n6523)
         );
  NAND2_X1 U8229 ( .A1(n6523), .A2(n6522), .ZN(n6525) );
  OAI21_X1 U8230 ( .B1(n7247), .B2(n6525), .A(n6524), .ZN(n6528) );
  INV_X1 U8231 ( .A(n6526), .ZN(n6527) );
  AOI21_X1 U8232 ( .B1(n6528), .B2(n4655), .A(n6527), .ZN(n6535) );
  INV_X1 U8233 ( .A(n6529), .ZN(n6532) );
  OAI211_X1 U8234 ( .C1(n6533), .C2(n6532), .A(n6531), .B(n6530), .ZN(n7099)
         );
  AOI21_X1 U8235 ( .B1(n6535), .B2(n7099), .A(n6534), .ZN(n6539) );
  INV_X1 U8236 ( .A(n6536), .ZN(n6537) );
  OAI211_X1 U8237 ( .C1(n6539), .C2(n6538), .A(n6537), .B(n9187), .ZN(n6540)
         );
  NAND4_X1 U8238 ( .A1(n6542), .A2(n9241), .A3(n6541), .A4(n6540), .ZN(n6544)
         );
  AOI21_X1 U8239 ( .B1(n6545), .B2(n6544), .A(n6543), .ZN(n6548) );
  OAI21_X1 U8240 ( .B1(n6548), .B2(n6547), .A(n6546), .ZN(n6549) );
  XNOR2_X1 U8241 ( .A(n6549), .B(n9298), .ZN(n6550) );
  NOR2_X1 U8242 ( .A1(n6550), .A2(n5660), .ZN(n6551) );
  INV_X1 U8243 ( .A(n6553), .ZN(n6557) );
  INV_X1 U8244 ( .A(n6554), .ZN(n6555) );
  NOR4_X1 U8245 ( .A1(n6557), .A2(n6556), .A3(n6708), .A4(n6555), .ZN(n6560)
         );
  NAND2_X1 U8246 ( .A1(n6577), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7755) );
  INV_X1 U8247 ( .A(n7755), .ZN(n6559) );
  OAI21_X1 U8248 ( .B1(n6561), .B2(n6560), .A(n6559), .ZN(n6567) );
  OR2_X1 U8249 ( .A1(n4280), .A2(P1_U3084), .ZN(n8031) );
  NOR4_X1 U8250 ( .A1(n7125), .A2(n5671), .A3(n6563), .A4(n8031), .ZN(n6565)
         );
  OAI21_X1 U8251 ( .B1(n5655), .B2(n7755), .A(P1_B_REG_SCAN_IN), .ZN(n6564) );
  OR2_X1 U8252 ( .A1(n6565), .A2(n6564), .ZN(n6566) );
  NAND2_X1 U8253 ( .A1(n6567), .A2(n6566), .ZN(P1_U3240) );
  INV_X1 U8254 ( .A(n6569), .ZN(n7601) );
  AOI211_X1 U8255 ( .C1(n6571), .C2(n6570), .A(n8593), .B(n7601), .ZN(n6576)
         );
  NOR2_X1 U8256 ( .A1(n8598), .A2(n7727), .ZN(n6575) );
  INV_X1 U8257 ( .A(n7735), .ZN(n6572) );
  OAI22_X1 U8258 ( .A1(n8597), .A2(n7726), .B1(n8585), .B2(n6572), .ZN(n6574)
         );
  INV_X1 U8259 ( .A(n7734), .ZN(n9979) );
  OAI22_X1 U8260 ( .A1(n8604), .A2(n9979), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5835), .ZN(n6573) );
  OR4_X1 U8261 ( .A1(n6576), .A2(n6575), .A3(n6574), .A4(n6573), .ZN(P2_U3215)
         );
  OR2_X1 U8262 ( .A1(n6708), .A2(n6577), .ZN(n6578) );
  NAND2_X1 U8263 ( .A1(n6578), .A2(n6613), .ZN(n6597) );
  OR2_X1 U8264 ( .A1(n6597), .A2(n6579), .ZN(n9616) );
  NAND2_X1 U8265 ( .A1(n9616), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  AND2_X1 U8266 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7487) );
  OR2_X1 U8267 ( .A1(n6775), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6581) );
  NAND2_X1 U8268 ( .A1(n6775), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6580) );
  NAND2_X1 U8269 ( .A1(n6581), .A2(n6580), .ZN(n6595) );
  INV_X1 U8270 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6582) );
  MUX2_X1 U8271 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n6582), .S(n6864), .Z(n6867)
         );
  AND2_X1 U8272 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n6866) );
  NAND2_X1 U8273 ( .A1(n6867), .A2(n6866), .ZN(n6865) );
  NAND2_X1 U8274 ( .A1(n6864), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6583) );
  NAND2_X1 U8275 ( .A1(n6865), .A2(n6583), .ZN(n6850) );
  NAND2_X1 U8276 ( .A1(n6855), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6584) );
  INV_X1 U8277 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6585) );
  XNOR2_X1 U8278 ( .A(n6622), .B(n6585), .ZN(n6827) );
  NAND2_X1 U8279 ( .A1(n6622), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6586) );
  NAND2_X1 U8280 ( .A1(n6825), .A2(n6586), .ZN(n6793) );
  XNOR2_X1 U8281 ( .A(n6602), .B(P1_REG2_REG_4__SCAN_IN), .ZN(n6792) );
  OR2_X1 U8282 ( .A1(n6793), .A2(n6792), .ZN(n6795) );
  INV_X1 U8283 ( .A(n6602), .ZN(n6804) );
  INV_X1 U8284 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n9794) );
  NAND2_X1 U8285 ( .A1(n6804), .A2(n9794), .ZN(n6587) );
  NAND2_X1 U8286 ( .A1(n6795), .A2(n6587), .ZN(n6872) );
  INV_X1 U8287 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n6588) );
  XNOR2_X1 U8288 ( .A(n6625), .B(n6588), .ZN(n6871) );
  NOR2_X1 U8289 ( .A1(n6625), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6589) );
  AOI21_X1 U8290 ( .B1(n6872), .B2(n6871), .A(n6589), .ZN(n9622) );
  INV_X1 U8291 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n9744) );
  XNOR2_X1 U8292 ( .A(n6640), .B(n9744), .ZN(n9623) );
  NAND2_X1 U8293 ( .A1(n6640), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6590) );
  XNOR2_X1 U8294 ( .A(n6647), .B(P1_REG2_REG_7__SCAN_IN), .ZN(n8359) );
  OR2_X1 U8295 ( .A1(n6647), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6591) );
  XNOR2_X1 U8296 ( .A(n6745), .B(n6592), .ZN(n6737) );
  NAND2_X1 U8297 ( .A1(n6736), .A2(n6737), .ZN(n6735) );
  INV_X1 U8298 ( .A(n6745), .ZN(n6650) );
  NAND2_X1 U8299 ( .A1(n6650), .A2(n6592), .ZN(n6593) );
  NAND2_X1 U8300 ( .A1(n6735), .A2(n6593), .ZN(n6594) );
  NOR2_X1 U8301 ( .A1(n6594), .A2(n6595), .ZN(n6774) );
  AOI211_X1 U8302 ( .C1(n6595), .C2(n6594), .A(n6774), .B(n9681), .ZN(n6616)
         );
  NAND2_X1 U8303 ( .A1(n4280), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6596) );
  INV_X1 U8304 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n9875) );
  MUX2_X1 U8305 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n9875), .S(n6855), .Z(n6846)
         );
  INV_X1 U8306 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n9873) );
  MUX2_X1 U8307 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n9873), .S(n6864), .Z(n6861)
         );
  AND2_X1 U8308 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n6860) );
  NAND2_X1 U8309 ( .A1(n6861), .A2(n6860), .ZN(n6859) );
  NAND2_X1 U8310 ( .A1(n6864), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6598) );
  NAND2_X1 U8311 ( .A1(n6859), .A2(n6598), .ZN(n6845) );
  NAND2_X1 U8312 ( .A1(n6846), .A2(n6845), .ZN(n6844) );
  NAND2_X1 U8313 ( .A1(n6855), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6599) );
  NAND2_X1 U8314 ( .A1(n6844), .A2(n6599), .ZN(n6819) );
  INV_X1 U8315 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6600) );
  XNOR2_X1 U8316 ( .A(n6622), .B(n6600), .ZN(n6820) );
  NAND2_X1 U8317 ( .A1(n6819), .A2(n6820), .ZN(n6818) );
  NAND2_X1 U8318 ( .A1(n6622), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6601) );
  NAND2_X1 U8319 ( .A1(n6818), .A2(n6601), .ZN(n6798) );
  XNOR2_X1 U8320 ( .A(n6602), .B(P1_REG1_REG_4__SCAN_IN), .ZN(n6797) );
  OR2_X1 U8321 ( .A1(n6798), .A2(n6797), .ZN(n6800) );
  INV_X1 U8322 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6603) );
  NAND2_X1 U8323 ( .A1(n6804), .A2(n6603), .ZN(n6604) );
  AND2_X1 U8324 ( .A1(n6800), .A2(n6604), .ZN(n6874) );
  OR2_X1 U8325 ( .A1(n6625), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6605) );
  NAND2_X1 U8326 ( .A1(n6625), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n9627) );
  AND2_X1 U8327 ( .A1(n6605), .A2(n9627), .ZN(n6873) );
  NAND2_X1 U8328 ( .A1(n6874), .A2(n6873), .ZN(n9628) );
  INV_X1 U8329 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6606) );
  XNOR2_X1 U8330 ( .A(n6640), .B(n6606), .ZN(n9626) );
  AND2_X1 U8331 ( .A1(n9626), .A2(n9627), .ZN(n6607) );
  NAND2_X1 U8332 ( .A1(n9628), .A2(n6607), .ZN(n9625) );
  OAI21_X1 U8333 ( .B1(n6640), .B2(P1_REG1_REG_6__SCAN_IN), .A(n9625), .ZN(
        n8361) );
  XOR2_X1 U8334 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n6647), .Z(n8362) );
  NAND2_X1 U8335 ( .A1(n8361), .A2(n8362), .ZN(n8360) );
  OAI21_X1 U8336 ( .B1(P1_REG1_REG_7__SCAN_IN), .B2(n6647), .A(n8360), .ZN(
        n6740) );
  NAND2_X1 U8337 ( .A1(n6745), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6738) );
  INV_X1 U8338 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6608) );
  NAND2_X1 U8339 ( .A1(n6650), .A2(n6608), .ZN(n6739) );
  INV_X1 U8340 ( .A(n6739), .ZN(n6609) );
  AOI21_X1 U8341 ( .B1(n6740), .B2(n6738), .A(n6609), .ZN(n6611) );
  INV_X1 U8342 ( .A(n6775), .ZN(n6654) );
  AOI22_X1 U8343 ( .A1(n6775), .A2(n5238), .B1(P1_REG1_REG_9__SCAN_IN), .B2(
        n6654), .ZN(n6610) );
  NOR2_X1 U8344 ( .A1(n6611), .A2(n6610), .ZN(n6761) );
  AOI21_X1 U8345 ( .B1(n6611), .B2(n6610), .A(n6761), .ZN(n6612) );
  NOR2_X1 U8346 ( .A1(n9724), .A2(n6612), .ZN(n6615) );
  INV_X1 U8347 ( .A(n6613), .ZN(n6790) );
  INV_X1 U8348 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10086) );
  OAI22_X1 U8349 ( .A1(n9727), .A2(n10086), .B1(n6654), .B2(n9717), .ZN(n6614)
         );
  OR4_X1 U8350 ( .A1(n7487), .A2(n6616), .A3(n6615), .A4(n6614), .ZN(P1_U3250)
         );
  INV_X1 U8351 ( .A(n6617), .ZN(n6618) );
  NAND2_X1 U8352 ( .A1(P1_STATE_REG_SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n6788) );
  OAI21_X1 U8353 ( .B1(n6618), .B2(P1_STATE_REG_SCAN_IN), .A(n6788), .ZN(
        P1_U3353) );
  AOI22_X1 U8354 ( .A1(P2_DATAO_REG_2__SCAN_IN), .A2(n9496), .B1(n6855), .B2(
        P1_STATE_REG_SCAN_IN), .ZN(n6619) );
  OAI21_X1 U8355 ( .B1(n6637), .B2(n4282), .A(n6619), .ZN(P1_U3351) );
  INV_X1 U8356 ( .A(n9496), .ZN(n9502) );
  INV_X1 U8357 ( .A(n6864), .ZN(n6620) );
  OAI222_X1 U8358 ( .A1(n9502), .A2(n6621), .B1(n4282), .B2(n6634), .C1(
        P1_U3084), .C2(n6620), .ZN(P1_U3352) );
  INV_X1 U8359 ( .A(n6622), .ZN(n6823) );
  OAI222_X1 U8360 ( .A1(n9502), .A2(n6623), .B1(n4282), .B2(n6630), .C1(
        P1_U3084), .C2(n6823), .ZN(P1_U3350) );
  OAI222_X1 U8361 ( .A1(n9502), .A2(n6624), .B1(n4282), .B2(n6632), .C1(
        P1_U3084), .C2(n6804), .ZN(P1_U3349) );
  INV_X1 U8362 ( .A(n6625), .ZN(n6876) );
  OAI222_X1 U8363 ( .A1(n9502), .A2(n6626), .B1(n4282), .B2(n6627), .C1(
        P1_U3084), .C2(n6876), .ZN(P1_U3348) );
  NAND2_X1 U8364 ( .A1(n4283), .A2(P2_U3152), .ZN(n9047) );
  INV_X1 U8365 ( .A(n9047), .ZN(n7350) );
  INV_X1 U8366 ( .A(n7350), .ZN(n9041) );
  NOR2_X1 U8367 ( .A1(n4278), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9044) );
  INV_X2 U8368 ( .A(n9044), .ZN(n9049) );
  OAI222_X1 U8369 ( .A1(n9041), .A2(n6628), .B1(n9049), .B2(n6627), .C1(
        P2_U3152), .C2(n6982), .ZN(P2_U3353) );
  OAI222_X1 U8370 ( .A1(P2_U3152), .A2(n7006), .B1(n9049), .B2(n6630), .C1(
        n6629), .C2(n9041), .ZN(P2_U3355) );
  OAI222_X1 U8371 ( .A1(P2_U3152), .A2(n6958), .B1(n9049), .B2(n6632), .C1(
        n6631), .C2(n9041), .ZN(P2_U3354) );
  OAI222_X1 U8372 ( .A1(P2_U3152), .A2(n6635), .B1(n9049), .B2(n6634), .C1(
        n6633), .C2(n9041), .ZN(P2_U3357) );
  OAI222_X1 U8373 ( .A1(P2_U3152), .A2(n6638), .B1(n9049), .B2(n6637), .C1(
        n6636), .C2(n9041), .ZN(P2_U3356) );
  INV_X1 U8374 ( .A(n6640), .ZN(n9635) );
  INV_X1 U8375 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n6645) );
  INV_X1 U8376 ( .A(n6643), .ZN(n6644) );
  AOI22_X1 U8377 ( .A1(n9809), .A2(n6645), .B1(n6688), .B2(n6644), .ZN(
        P1_U3441) );
  OAI222_X1 U8378 ( .A1(n9041), .A2(n6646), .B1(n9049), .B2(n6648), .C1(
        P2_U3152), .C2(n6970), .ZN(P2_U3351) );
  INV_X1 U8379 ( .A(n6647), .ZN(n8363) );
  OAI222_X1 U8380 ( .A1(n9502), .A2(n6649), .B1(n4282), .B2(n6648), .C1(
        P1_U3084), .C2(n8363), .ZN(P1_U3346) );
  OAI222_X1 U8381 ( .A1(n9502), .A2(n6651), .B1(n4282), .B2(n5863), .C1(
        P1_U3084), .C2(n6650), .ZN(P1_U3345) );
  OAI222_X1 U8382 ( .A1(n9041), .A2(n6652), .B1(n9049), .B2(n5863), .C1(
        P2_U3152), .C2(n6843), .ZN(P2_U3350) );
  OAI222_X1 U8383 ( .A1(n9041), .A2(n6653), .B1(n9049), .B2(n6655), .C1(n6994), 
        .C2(P2_U3152), .ZN(P2_U3349) );
  OAI222_X1 U8384 ( .A1(n9502), .A2(n6656), .B1(n4282), .B2(n6655), .C1(n6654), 
        .C2(P1_U3084), .ZN(P1_U3344) );
  INV_X1 U8385 ( .A(n6657), .ZN(n6661) );
  INV_X1 U8386 ( .A(n6776), .ZN(n8348) );
  OAI222_X1 U8387 ( .A1(n9502), .A2(n6658), .B1(n4282), .B2(n6661), .C1(n8348), 
        .C2(P1_U3084), .ZN(P1_U3343) );
  INV_X1 U8388 ( .A(n6659), .ZN(n6904) );
  OAI222_X1 U8389 ( .A1(P2_U3152), .A2(n6904), .B1(n9049), .B2(n6661), .C1(
        n6660), .C2(n9041), .ZN(P2_U3348) );
  INV_X1 U8390 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n6663) );
  NAND2_X1 U8391 ( .A1(n4281), .A2(n7011), .ZN(n6662) );
  OAI21_X1 U8392 ( .B1(n4281), .B2(n6663), .A(n6662), .ZN(P1_U3555) );
  INV_X1 U8393 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6665) );
  NAND2_X1 U8394 ( .A1(n4281), .A2(n9165), .ZN(n6664) );
  OAI21_X1 U8395 ( .B1(n4281), .B2(n6665), .A(n6664), .ZN(P1_U3586) );
  INV_X1 U8396 ( .A(n6666), .ZN(n6668) );
  INV_X1 U8397 ( .A(n8334), .ZN(n6773) );
  OAI222_X1 U8398 ( .A1(n9502), .A2(n6667), .B1(n4282), .B2(n6668), .C1(n6773), 
        .C2(P1_U3084), .ZN(P1_U3342) );
  OAI222_X1 U8399 ( .A1(n9041), .A2(n6669), .B1(n9049), .B2(n6668), .C1(n7066), 
        .C2(P2_U3152), .ZN(P2_U3347) );
  NAND2_X1 U8400 ( .A1(n4275), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n6672) );
  NAND2_X1 U8401 ( .A1(n6148), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n6671) );
  NAND2_X1 U8402 ( .A1(n6722), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n6670) );
  NAND2_X1 U8403 ( .A1(n6760), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n6673) );
  OAI21_X1 U8404 ( .B1(n6760), .B2(n8449), .A(n6673), .ZN(P2_U3582) );
  INV_X1 U8405 ( .A(n6674), .ZN(n6677) );
  OAI222_X1 U8406 ( .A1(n9502), .A2(n6675), .B1(n4282), .B2(n6677), .C1(
        P1_U3084), .C2(n8291), .ZN(P1_U3341) );
  OAI222_X1 U8407 ( .A1(n9047), .A2(n6678), .B1(n9049), .B2(n6677), .C1(
        P2_U3152), .C2(n6676), .ZN(P2_U3346) );
  INV_X1 U8408 ( .A(n6679), .ZN(n6682) );
  AOI22_X1 U8409 ( .A1(n9645), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n9496), .ZN(n6680) );
  OAI21_X1 U8410 ( .B1(n6682), .B2(n4282), .A(n6680), .ZN(P1_U3340) );
  OAI222_X1 U8411 ( .A1(n9047), .A2(n7440), .B1(n9049), .B2(n6682), .C1(n6681), 
        .C2(P2_U3152), .ZN(P2_U3345) );
  INV_X1 U8412 ( .A(n6683), .ZN(n6686) );
  OAI222_X1 U8413 ( .A1(n9502), .A2(n6684), .B1(n4282), .B2(n6686), .C1(n9660), 
        .C2(P1_U3084), .ZN(P1_U3339) );
  OAI222_X1 U8414 ( .A1(n9047), .A2(n6687), .B1(n9049), .B2(n6686), .C1(n6685), 
        .C2(P2_U3152), .ZN(P2_U3344) );
  NOR2_X1 U8415 ( .A1(n9892), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U8416 ( .A(n6716), .ZN(n6691) );
  AND3_X1 U8417 ( .A1(n6692), .A2(n6691), .A3(n6690), .ZN(n6754) );
  INV_X1 U8418 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n7178) );
  INV_X1 U8419 ( .A(n6693), .ZN(n9162) );
  AOI22_X1 U8420 ( .A1(n7176), .A2(n9129), .B1(n9145), .B2(n9162), .ZN(n6698)
         );
  OAI21_X1 U8421 ( .B1(n6696), .B2(n6695), .A(n6694), .ZN(n6784) );
  NAND2_X1 U8422 ( .A1(n6784), .A2(n9136), .ZN(n6697) );
  OAI211_X1 U8423 ( .C1(n6754), .C2(n7178), .A(n6698), .B(n6697), .ZN(P1_U3230) );
  INV_X1 U8424 ( .A(n6699), .ZN(n6700) );
  NOR2_X1 U8425 ( .A1(n6701), .A2(n6700), .ZN(n6704) );
  OAI21_X1 U8426 ( .B1(n6701), .B2(P1_D_REG_0__SCAN_IN), .A(n9491), .ZN(n6702)
         );
  INV_X1 U8427 ( .A(n6702), .ZN(n6703) );
  OR2_X1 U8428 ( .A1(n9818), .A2(n6705), .ZN(n6707) );
  INV_X1 U8429 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6714) );
  NOR3_X1 U8430 ( .A1(n6711), .A2(n6710), .A3(n6709), .ZN(n6712) );
  AOI21_X1 U8431 ( .B1(n9736), .B2(n9162), .A(n6712), .ZN(n7177) );
  OAI21_X1 U8432 ( .B1(n7031), .B2(n7029), .A(n7177), .ZN(n6719) );
  NAND2_X1 U8433 ( .A1(n6719), .A2(n9872), .ZN(n6713) );
  OAI21_X1 U8434 ( .B1(n9872), .B2(n6714), .A(n6713), .ZN(P1_U3454) );
  NOR2_X1 U8435 ( .A1(n6716), .A2(n6715), .ZN(n6717) );
  NAND2_X1 U8436 ( .A1(n6719), .A2(n9887), .ZN(n6720) );
  OAI21_X1 U8437 ( .B1(n9887), .B2(n5098), .A(n6720), .ZN(P1_U3523) );
  NAND2_X1 U8438 ( .A1(n4275), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n6725) );
  NAND2_X1 U8439 ( .A1(n6721), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n6724) );
  NAND2_X1 U8440 ( .A1(n6722), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n6723) );
  NAND3_X1 U8441 ( .A1(n6725), .A2(n6724), .A3(n6723), .ZN(n8662) );
  NAND2_X1 U8442 ( .A1(P2_U3966), .A2(n8662), .ZN(n6726) );
  OAI21_X1 U8443 ( .B1(P2_U3966), .B2(n6413), .A(n6726), .ZN(P2_U3583) );
  XNOR2_X1 U8444 ( .A(n6728), .B(n6727), .ZN(n6729) );
  XOR2_X1 U8445 ( .A(n6730), .B(n6729), .Z(n6734) );
  OAI22_X1 U8446 ( .A1(n5092), .A2(n9114), .B1(n9123), .B2(n6307), .ZN(n6732)
         );
  NOR2_X1 U8447 ( .A1(n6754), .A2(n7032), .ZN(n6731) );
  AOI211_X1 U8448 ( .C1(n7034), .C2(n9129), .A(n6732), .B(n6731), .ZN(n6733)
         );
  OAI21_X1 U8449 ( .B1(n9131), .B2(n6734), .A(n6733), .ZN(P1_U3220) );
  INV_X1 U8450 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n6748) );
  OAI21_X1 U8451 ( .B1(n6737), .B2(n6736), .A(n6735), .ZN(n6743) );
  NAND2_X1 U8452 ( .A1(n6739), .A2(n6738), .ZN(n6741) );
  XOR2_X1 U8453 ( .A(n6741), .B(n6740), .Z(n6742) );
  AOI22_X1 U8454 ( .A1(n9714), .A2(n6743), .B1(n9704), .B2(n6742), .ZN(n6747)
         );
  NOR2_X1 U8455 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6744), .ZN(n7312) );
  AOI21_X1 U8456 ( .B1(n9688), .B2(n6745), .A(n7312), .ZN(n6746) );
  OAI211_X1 U8457 ( .C1(n9727), .C2(n6748), .A(n6747), .B(n6746), .ZN(P1_U3249) );
  INV_X1 U8458 ( .A(n6749), .ZN(n6808) );
  AOI22_X1 U8459 ( .A1(n9674), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n9496), .ZN(n6750) );
  OAI21_X1 U8460 ( .B1(n6808), .B2(n4282), .A(n6750), .ZN(P1_U3338) );
  OAI21_X1 U8461 ( .B1(n6753), .B2(n6752), .A(n6751), .ZN(n6757) );
  OAI22_X1 U8462 ( .A1(n6693), .A2(n9114), .B1(n9123), .B2(n9783), .ZN(n6756)
         );
  INV_X1 U8463 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n6848) );
  OAI22_X1 U8464 ( .A1(n6754), .A2(n6848), .B1(n7255), .B2(n9148), .ZN(n6755)
         );
  AOI211_X1 U8465 ( .C1(n6757), .C2(n9136), .A(n6756), .B(n6755), .ZN(n6758)
         );
  INV_X1 U8466 ( .A(n6758), .ZN(P1_U3235) );
  NAND2_X1 U8467 ( .A1(n6760), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n6759) );
  OAI21_X1 U8468 ( .B1(n6760), .B2(n8081), .A(n6759), .ZN(P2_U3581) );
  INV_X1 U8469 ( .A(n9727), .ZN(n8367) );
  NAND2_X1 U8470 ( .A1(P1_U3084), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7654) );
  MUX2_X1 U8471 ( .A(n5328), .B(P1_REG1_REG_12__SCAN_IN), .S(n8291), .Z(n6768)
         );
  INV_X1 U8472 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n6765) );
  NOR2_X1 U8473 ( .A1(n6775), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6762) );
  NOR2_X1 U8474 ( .A1(n6762), .A2(n6761), .ZN(n8345) );
  INV_X1 U8475 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6763) );
  MUX2_X1 U8476 ( .A(n6763), .B(P1_REG1_REG_10__SCAN_IN), .S(n6776), .Z(n8344)
         );
  OR2_X1 U8477 ( .A1(n8345), .A2(n8344), .ZN(n8342) );
  OR2_X1 U8478 ( .A1(n6776), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6764) );
  AND2_X1 U8479 ( .A1(n8342), .A2(n6764), .ZN(n8330) );
  AOI22_X1 U8480 ( .A1(P1_REG1_REG_11__SCAN_IN), .A2(n6773), .B1(n8334), .B2(
        n6765), .ZN(n8329) );
  NOR2_X1 U8481 ( .A1(n8330), .A2(n8329), .ZN(n8328) );
  AOI21_X1 U8482 ( .B1(n6765), .B2(n6773), .A(n8328), .ZN(n6766) );
  INV_X1 U8483 ( .A(n6766), .ZN(n6767) );
  NAND2_X1 U8484 ( .A1(n6768), .A2(n6767), .ZN(n8289) );
  OAI21_X1 U8485 ( .B1(n6768), .B2(n6767), .A(n8289), .ZN(n6769) );
  NAND2_X1 U8486 ( .A1(n9704), .A2(n6769), .ZN(n6770) );
  OAI211_X1 U8487 ( .C1(n9717), .C2(n8291), .A(n7654), .B(n6770), .ZN(n6782)
         );
  XNOR2_X1 U8488 ( .A(n8291), .B(n6771), .ZN(n6780) );
  OR2_X1 U8489 ( .A1(n8334), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6777) );
  INV_X1 U8490 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n6772) );
  AOI22_X1 U8491 ( .A1(P1_REG2_REG_11__SCAN_IN), .A2(n8334), .B1(n6773), .B2(
        n6772), .ZN(n8332) );
  AOI21_X1 U8492 ( .B1(n6775), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6774), .ZN(
        n8351) );
  XNOR2_X1 U8493 ( .A(n6776), .B(P1_REG2_REG_10__SCAN_IN), .ZN(n8350) );
  NOR2_X1 U8494 ( .A1(n8351), .A2(n8350), .ZN(n8349) );
  INV_X1 U8495 ( .A(n8273), .ZN(n6778) );
  AOI211_X1 U8496 ( .C1(n6780), .C2(n6779), .A(n6778), .B(n9681), .ZN(n6781)
         );
  AOI211_X1 U8497 ( .C1(P1_ADDR_REG_12__SCAN_IN), .C2(n8367), .A(n6782), .B(
        n6781), .ZN(n6783) );
  INV_X1 U8498 ( .A(n6783), .ZN(P1_U3253) );
  INV_X1 U8499 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n6807) );
  INV_X1 U8500 ( .A(n6784), .ZN(n6786) );
  INV_X1 U8501 ( .A(n4280), .ZN(n9164) );
  NOR2_X1 U8502 ( .A1(n4280), .A2(n6866), .ZN(n6785) );
  NOR2_X1 U8503 ( .A1(n6785), .A2(n5671), .ZN(n9612) );
  OAI21_X1 U8504 ( .B1(n6786), .B2(n9164), .A(n9612), .ZN(n6791) );
  NAND2_X1 U8505 ( .A1(n7024), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8054) );
  NOR2_X1 U8506 ( .A1(n4280), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6787) );
  OR2_X1 U8507 ( .A1(n8054), .A2(n6787), .ZN(n6789) );
  NAND2_X1 U8508 ( .A1(n6789), .A2(n6788), .ZN(n9614) );
  NAND3_X1 U8509 ( .A1(n6791), .A2(n6790), .A3(n9614), .ZN(n6856) );
  NAND2_X1 U8510 ( .A1(n6793), .A2(n6792), .ZN(n6794) );
  NAND2_X1 U8511 ( .A1(n6795), .A2(n6794), .ZN(n6796) );
  NAND2_X1 U8512 ( .A1(n9714), .A2(n6796), .ZN(n6803) );
  NAND2_X1 U8513 ( .A1(n6798), .A2(n6797), .ZN(n6799) );
  NAND2_X1 U8514 ( .A1(n6800), .A2(n6799), .ZN(n6801) );
  AND2_X1 U8515 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n6890) );
  AOI21_X1 U8516 ( .B1(n9704), .B2(n6801), .A(n6890), .ZN(n6802) );
  OAI211_X1 U8517 ( .C1(n9717), .C2(n6804), .A(n6803), .B(n6802), .ZN(n6805)
         );
  INV_X1 U8518 ( .A(n6805), .ZN(n6806) );
  OAI211_X1 U8519 ( .C1(n6807), .C2(n9727), .A(n6856), .B(n6806), .ZN(P1_U3245) );
  OAI222_X1 U8520 ( .A1(n9047), .A2(n6809), .B1(n9049), .B2(n6808), .C1(
        P2_U3152), .C2(n7955), .ZN(P2_U3343) );
  OAI21_X1 U8521 ( .B1(n6812), .B2(n6811), .A(n6810), .ZN(n6813) );
  NAND2_X1 U8522 ( .A1(n6813), .A2(n9136), .ZN(n6817) );
  OAI22_X1 U8523 ( .A1(n9823), .A2(n9148), .B1(n9114), .B2(n6307), .ZN(n6815)
         );
  INV_X1 U8524 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n7298) );
  OR2_X1 U8525 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7298), .ZN(n6821) );
  OAI21_X1 U8526 ( .B1(n9123), .B2(n9767), .A(n6821), .ZN(n6814) );
  NOR2_X1 U8527 ( .A1(n6815), .A2(n6814), .ZN(n6816) );
  OAI211_X1 U8528 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n9127), .A(n6817), .B(
        n6816), .ZN(P1_U3216) );
  INV_X1 U8529 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n6830) );
  OAI211_X1 U8530 ( .C1(n6820), .C2(n6819), .A(n9704), .B(n6818), .ZN(n6822)
         );
  OAI211_X1 U8531 ( .C1(n9717), .C2(n6823), .A(n6822), .B(n6821), .ZN(n6824)
         );
  INV_X1 U8532 ( .A(n6824), .ZN(n6829) );
  OAI211_X1 U8533 ( .C1(n6827), .C2(n6826), .A(n9714), .B(n6825), .ZN(n6828)
         );
  OAI211_X1 U8534 ( .C1(n6830), .C2(n9727), .A(n6829), .B(n6828), .ZN(P1_U3244) );
  NOR2_X1 U8535 ( .A1(n6831), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7607) );
  AOI211_X1 U8536 ( .C1(n6834), .C2(n6833), .A(n6832), .B(n9894), .ZN(n6835)
         );
  AOI211_X1 U8537 ( .C1(n9892), .C2(P2_ADDR_REG_8__SCAN_IN), .A(n7607), .B(
        n6835), .ZN(n6842) );
  INV_X1 U8538 ( .A(n6836), .ZN(n6840) );
  INV_X1 U8539 ( .A(n6837), .ZN(n6839) );
  OAI211_X1 U8540 ( .C1(n6840), .C2(n6839), .A(n9889), .B(n6838), .ZN(n6841)
         );
  OAI211_X1 U8541 ( .C1(n9893), .C2(n6843), .A(n6842), .B(n6841), .ZN(P2_U3253) );
  INV_X1 U8542 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n6858) );
  OAI211_X1 U8543 ( .C1(n6846), .C2(n6845), .A(n9704), .B(n6844), .ZN(n6847)
         );
  OAI21_X1 U8544 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n6848), .A(n6847), .ZN(n6854) );
  OAI211_X1 U8545 ( .C1(n6851), .C2(n6850), .A(n9714), .B(n6849), .ZN(n6852)
         );
  INV_X1 U8546 ( .A(n6852), .ZN(n6853) );
  AOI211_X1 U8547 ( .C1(n9688), .C2(n6855), .A(n6854), .B(n6853), .ZN(n6857)
         );
  OAI211_X1 U8548 ( .C1(n6858), .C2(n9727), .A(n6857), .B(n6856), .ZN(P1_U3243) );
  INV_X1 U8549 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n6870) );
  OAI211_X1 U8550 ( .C1(n6861), .C2(n6860), .A(n9704), .B(n6859), .ZN(n6862)
         );
  OAI21_X1 U8551 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n7032), .A(n6862), .ZN(n6863) );
  AOI21_X1 U8552 ( .B1(n6864), .B2(n9688), .A(n6863), .ZN(n6869) );
  OAI211_X1 U8553 ( .C1(n6867), .C2(n6866), .A(n9714), .B(n6865), .ZN(n6868)
         );
  OAI211_X1 U8554 ( .C1(n6870), .C2(n9727), .A(n6869), .B(n6868), .ZN(P1_U3242) );
  INV_X1 U8555 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n6880) );
  XNOR2_X1 U8556 ( .A(n6872), .B(n6871), .ZN(n6878) );
  OAI211_X1 U8557 ( .C1(n6874), .C2(n6873), .A(n9704), .B(n9628), .ZN(n6875)
         );
  NAND2_X1 U8558 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n7222) );
  OAI211_X1 U8559 ( .C1(n9717), .C2(n6876), .A(n6875), .B(n7222), .ZN(n6877)
         );
  AOI21_X1 U8560 ( .B1(n9714), .B2(n6878), .A(n6877), .ZN(n6879) );
  OAI21_X1 U8561 ( .B1(n9727), .B2(n6880), .A(n6879), .ZN(P1_U3246) );
  INV_X1 U8562 ( .A(n6881), .ZN(n6884) );
  AOI22_X1 U8563 ( .A1(n8628), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n7350), .ZN(n6882) );
  OAI21_X1 U8564 ( .B1(n6884), .B2(n9049), .A(n6882), .ZN(P2_U3342) );
  AOI22_X1 U8565 ( .A1(n9687), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n9496), .ZN(n6883) );
  OAI21_X1 U8566 ( .B1(n6884), .B2(n4282), .A(n6883), .ZN(P1_U3337) );
  AND2_X1 U8567 ( .A1(n6810), .A2(n6885), .ZN(n6888) );
  OAI211_X1 U8568 ( .C1(n6888), .C2(n6887), .A(n9136), .B(n6886), .ZN(n6892)
         );
  OAI22_X1 U8569 ( .A1(n9829), .A2(n9148), .B1(n9114), .B2(n9783), .ZN(n6889)
         );
  AOI211_X1 U8570 ( .C1(n9145), .C2(n9733), .A(n6890), .B(n6889), .ZN(n6891)
         );
  OAI211_X1 U8571 ( .C1(n9127), .C2(n9793), .A(n6892), .B(n6891), .ZN(P1_U3228) );
  NOR2_X1 U8572 ( .A1(n6893), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7886) );
  AOI211_X1 U8573 ( .C1(n6896), .C2(n6895), .A(n6894), .B(n9894), .ZN(n6897)
         );
  AOI211_X1 U8574 ( .C1(n9892), .C2(P2_ADDR_REG_10__SCAN_IN), .A(n7886), .B(
        n6897), .ZN(n6903) );
  INV_X1 U8575 ( .A(n6898), .ZN(n6901) );
  OAI211_X1 U8576 ( .C1(n6901), .C2(n4500), .A(n9889), .B(n6900), .ZN(n6902)
         );
  OAI211_X1 U8577 ( .C1(n9893), .C2(n6904), .A(n6903), .B(n6902), .ZN(P2_U3255) );
  INV_X1 U8578 ( .A(n7515), .ZN(n6909) );
  NAND2_X1 U8579 ( .A1(n6905), .A2(n7512), .ZN(n6906) );
  INV_X1 U8580 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n6932) );
  INV_X1 U8581 ( .A(n9953), .ZN(n6913) );
  NAND3_X1 U8582 ( .A1(n6914), .A2(n6913), .A3(n6912), .ZN(n8883) );
  AND2_X1 U8583 ( .A1(n7496), .A2(n4284), .ZN(n7528) );
  NAND2_X1 U8584 ( .A1(n8122), .A2(n7528), .ZN(n9541) );
  INV_X1 U8585 ( .A(n8143), .ZN(n6919) );
  INV_X1 U8586 ( .A(n8414), .ZN(n7585) );
  NAND4_X1 U8587 ( .A1(n6918), .A2(n6917), .A3(n6916), .A4(n6915), .ZN(n8621)
         );
  NAND2_X1 U8588 ( .A1(n7585), .A2(n8621), .ZN(n8134) );
  INV_X1 U8589 ( .A(n8134), .ZN(n8144) );
  NOR2_X1 U8590 ( .A1(n6919), .A2(n8144), .ZN(n6926) );
  INV_X1 U8591 ( .A(n6926), .ZN(n6920) );
  XOR2_X1 U8592 ( .A(n7067), .B(n6920), .Z(n7588) );
  INV_X1 U8593 ( .A(n7588), .ZN(n6930) );
  NAND2_X1 U8594 ( .A1(n8414), .A2(n9952), .ZN(n6921) );
  AND3_X1 U8595 ( .A1(n7615), .A2(n9913), .A3(n6921), .ZN(n7583) );
  NAND2_X1 U8596 ( .A1(n8268), .A2(n4284), .ZN(n8120) );
  OAI21_X1 U8597 ( .B1(n6926), .B2(n7590), .A(n9922), .ZN(n6928) );
  NOR2_X1 U8598 ( .A1(n7081), .A2(n8144), .ZN(n8094) );
  INV_X1 U8599 ( .A(n8425), .ZN(n8622) );
  AOI22_X1 U8600 ( .A1(n8861), .A2(n8622), .B1(n7071), .B2(n8862), .ZN(n6927)
         );
  OAI21_X1 U8601 ( .B1(n6928), .B2(n8094), .A(n6927), .ZN(n7582) );
  AOI211_X1 U8602 ( .C1(n9016), .C2(n8414), .A(n7583), .B(n7582), .ZN(n6929)
         );
  OAI21_X1 U8603 ( .B1(n10001), .B2(n6930), .A(n6929), .ZN(n6934) );
  NAND2_X1 U8604 ( .A1(n6934), .A2(n10028), .ZN(n6931) );
  OAI21_X1 U8605 ( .B1(n10028), .B2(n6932), .A(n6931), .ZN(P2_U3454) );
  NAND2_X1 U8606 ( .A1(n6934), .A2(n10045), .ZN(n6935) );
  OAI21_X1 U8607 ( .B1(n10045), .B2(n6936), .A(n6935), .ZN(P2_U3521) );
  AOI211_X1 U8608 ( .C1(n6939), .C2(n6938), .A(n6937), .B(n9895), .ZN(n6948)
         );
  NOR2_X1 U8609 ( .A1(n6940), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8397) );
  AOI21_X1 U8610 ( .B1(n9892), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n8397), .ZN(
        n6945) );
  OAI211_X1 U8611 ( .C1(n6943), .C2(n6942), .A(n9888), .B(n6941), .ZN(n6944)
         );
  OAI211_X1 U8612 ( .C1(n9893), .C2(n6946), .A(n6945), .B(n6944), .ZN(n6947)
         );
  OR2_X1 U8613 ( .A1(n6948), .A2(n6947), .ZN(P2_U3251) );
  AOI211_X1 U8614 ( .C1(n6951), .C2(n6950), .A(n6949), .B(n9895), .ZN(n6960)
         );
  AND2_X1 U8615 ( .A1(P2_U3152), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n6952) );
  AOI21_X1 U8616 ( .B1(n9892), .B2(P2_ADDR_REG_4__SCAN_IN), .A(n6952), .ZN(
        n6957) );
  OAI211_X1 U8617 ( .C1(n6955), .C2(n6954), .A(n9888), .B(n6953), .ZN(n6956)
         );
  OAI211_X1 U8618 ( .C1(n9893), .C2(n6958), .A(n6957), .B(n6956), .ZN(n6959)
         );
  OR2_X1 U8619 ( .A1(n6960), .A2(n6959), .ZN(P2_U3249) );
  AOI211_X1 U8620 ( .C1(n6963), .C2(n6962), .A(n6961), .B(n9895), .ZN(n6972)
         );
  NOR2_X1 U8621 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5835), .ZN(n6964) );
  AOI21_X1 U8622 ( .B1(n9892), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n6964), .ZN(
        n6969) );
  OAI211_X1 U8623 ( .C1(n6967), .C2(n6966), .A(n9888), .B(n6965), .ZN(n6968)
         );
  OAI211_X1 U8624 ( .C1(n9893), .C2(n6970), .A(n6969), .B(n6968), .ZN(n6971)
         );
  OR2_X1 U8625 ( .A1(n6972), .A2(n6971), .ZN(P2_U3252) );
  AOI211_X1 U8626 ( .C1(n6975), .C2(n6974), .A(n6973), .B(n9895), .ZN(n6984)
         );
  NOR2_X1 U8627 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7341), .ZN(n6976) );
  AOI21_X1 U8628 ( .B1(n9892), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n6976), .ZN(
        n6981) );
  OAI211_X1 U8629 ( .C1(n6979), .C2(n6978), .A(n9888), .B(n6977), .ZN(n6980)
         );
  OAI211_X1 U8630 ( .C1(n9893), .C2(n6982), .A(n6981), .B(n6980), .ZN(n6983)
         );
  OR2_X1 U8631 ( .A1(n6984), .A2(n6983), .ZN(P2_U3250) );
  AOI211_X1 U8632 ( .C1(n6987), .C2(n6986), .A(n6985), .B(n9895), .ZN(n6996)
         );
  NAND2_X1 U8633 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3152), .ZN(n7541) );
  INV_X1 U8634 ( .A(n7541), .ZN(n6988) );
  AOI21_X1 U8635 ( .B1(n9892), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n6988), .ZN(
        n6993) );
  OAI211_X1 U8636 ( .C1(n6991), .C2(n6990), .A(n9888), .B(n6989), .ZN(n6992)
         );
  OAI211_X1 U8637 ( .C1(n9893), .C2(n6994), .A(n6993), .B(n6992), .ZN(n6995)
         );
  OR2_X1 U8638 ( .A1(n6996), .A2(n6995), .ZN(P2_U3254) );
  AOI211_X1 U8639 ( .C1(n6999), .C2(n6998), .A(n6997), .B(n9895), .ZN(n7008)
         );
  INV_X1 U8640 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n9924) );
  NOR2_X1 U8641 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9924), .ZN(n7000) );
  AOI21_X1 U8642 ( .B1(n9892), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n7000), .ZN(
        n7005) );
  OAI211_X1 U8643 ( .C1(n7003), .C2(n7002), .A(n9888), .B(n7001), .ZN(n7004)
         );
  OAI211_X1 U8644 ( .C1(n9893), .C2(n7006), .A(n7005), .B(n7004), .ZN(n7007)
         );
  OR2_X1 U8645 ( .A1(n7008), .A2(n7007), .ZN(P2_U3248) );
  INV_X1 U8646 ( .A(n7009), .ZN(n7037) );
  AOI22_X1 U8647 ( .A1(n8288), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n9496), .ZN(n7010) );
  OAI21_X1 U8648 ( .B1(n7037), .B2(n4282), .A(n7010), .ZN(P1_U3336) );
  NAND2_X1 U8649 ( .A1(n7012), .A2(n7013), .ZN(n7108) );
  NAND2_X1 U8650 ( .A1(n7015), .A2(n7014), .ZN(n7103) );
  NOR2_X1 U8651 ( .A1(n5064), .A2(n9298), .ZN(n7016) );
  AND2_X1 U8652 ( .A1(n9797), .A2(n7016), .ZN(n9778) );
  INV_X1 U8653 ( .A(n9778), .ZN(n7337) );
  NAND2_X1 U8654 ( .A1(n7648), .A2(n9298), .ZN(n7018) );
  MUX2_X1 U8655 ( .A(n7018), .B(n7017), .S(n5064), .Z(n9789) );
  NAND2_X1 U8656 ( .A1(n5655), .A2(n9757), .ZN(n7020) );
  OAI21_X1 U8657 ( .B1(n7023), .B2(n7022), .A(n7021), .ZN(n7027) );
  OAI22_X1 U8658 ( .A1(n9784), .A2(n5092), .B1(n6307), .B2(n9781), .ZN(n7026)
         );
  AOI21_X1 U8659 ( .B1(n9786), .B2(n7027), .A(n7026), .ZN(n7028) );
  OAI21_X1 U8660 ( .B1(n9789), .B2(n9810), .A(n7028), .ZN(n9812) );
  INV_X1 U8661 ( .A(n7254), .ZN(n7030) );
  OAI211_X1 U8662 ( .C1(n4568), .C2(n7031), .A(n7030), .B(n9857), .ZN(n9811)
         );
  OAI22_X1 U8663 ( .A1(n9811), .A2(n9757), .B1(n9792), .B2(n7032), .ZN(n7033)
         );
  OAI21_X1 U8664 ( .B1(n9812), .B2(n7033), .A(n9797), .ZN(n7036) );
  AOI22_X1 U8665 ( .A1(n9569), .A2(n7034), .B1(n9568), .B2(
        P1_REG2_REG_1__SCAN_IN), .ZN(n7035) );
  OAI211_X1 U8666 ( .C1(n9810), .C2(n7337), .A(n7036), .B(n7035), .ZN(P1_U3290) );
  OAI222_X1 U8667 ( .A1(n9047), .A2(n7038), .B1(n9049), .B2(n7037), .C1(n8644), 
        .C2(P2_U3152), .ZN(P2_U3341) );
  INV_X1 U8668 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7040) );
  INV_X1 U8669 ( .A(n7039), .ZN(n7041) );
  OAI222_X1 U8670 ( .A1(n9047), .A2(n7040), .B1(n9049), .B2(n7041), .C1(
        P2_U3152), .C2(n8654), .ZN(P2_U3340) );
  INV_X1 U8671 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n7042) );
  INV_X1 U8672 ( .A(n8287), .ZN(n9718) );
  OAI222_X1 U8673 ( .A1(n9502), .A2(n7042), .B1(n4282), .B2(n7041), .C1(
        P1_U3084), .C2(n9718), .ZN(P1_U3335) );
  OAI21_X1 U8674 ( .B1(n7044), .B2(n8481), .A(n7343), .ZN(n7054) );
  INV_X1 U8675 ( .A(n7044), .ZN(n7046) );
  NAND3_X1 U8676 ( .A1(n7046), .A2(n7045), .A3(n8620), .ZN(n7048) );
  INV_X1 U8677 ( .A(n7522), .ZN(n7047) );
  OAI22_X1 U8678 ( .A1(n8592), .A2(n7048), .B1(n7047), .B2(n8585), .ZN(n7053)
         );
  OR2_X1 U8679 ( .A1(n7079), .A2(n8907), .ZN(n7050) );
  OR2_X1 U8680 ( .A1(n7074), .A2(n8905), .ZN(n7049) );
  NAND2_X1 U8681 ( .A1(n7050), .A2(n7049), .ZN(n7136) );
  AOI22_X1 U8682 ( .A1(n8509), .A2(n7136), .B1(P2_REG3_REG_4__SCAN_IN), .B2(
        P2_U3152), .ZN(n7051) );
  OAI21_X1 U8683 ( .B1(n8604), .B2(n7531), .A(n7051), .ZN(n7052) );
  AOI211_X1 U8684 ( .C1(n8488), .C2(n7054), .A(n7053), .B(n7052), .ZN(n7055)
         );
  INV_X1 U8685 ( .A(n7055), .ZN(P2_U3232) );
  NOR2_X1 U8686 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5917), .ZN(n7060) );
  XNOR2_X1 U8687 ( .A(n7057), .B(n7056), .ZN(n7058) );
  NOR2_X1 U8688 ( .A1(n9894), .A2(n7058), .ZN(n7059) );
  AOI211_X1 U8689 ( .C1(n9892), .C2(P2_ADDR_REG_11__SCAN_IN), .A(n7060), .B(
        n7059), .ZN(n7065) );
  OAI21_X1 U8690 ( .B1(n4323), .B2(n7062), .A(n7061), .ZN(n7063) );
  NAND2_X1 U8691 ( .A1(n9889), .A2(n7063), .ZN(n7064) );
  OAI211_X1 U8692 ( .C1(n9893), .C2(n7066), .A(n7065), .B(n7064), .ZN(P2_U3256) );
  INV_X1 U8693 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n7095) );
  OAI21_X1 U8694 ( .B1(n8621), .B2(n8414), .A(n7067), .ZN(n7069) );
  NAND2_X1 U8695 ( .A1(n8621), .A2(n8414), .ZN(n7068) );
  AND2_X1 U8696 ( .A1(n7069), .A2(n7068), .ZN(n7614) );
  NAND2_X2 U8697 ( .A1(n8146), .A2(n9918), .ZN(n7612) );
  NAND2_X1 U8698 ( .A1(n7614), .A2(n7612), .ZN(n7613) );
  NAND2_X1 U8699 ( .A1(n7072), .A2(n7070), .ZN(n7073) );
  NAND2_X1 U8700 ( .A1(n7613), .A2(n7073), .ZN(n9926) );
  NAND2_X1 U8701 ( .A1(n7074), .A2(n9932), .ZN(n8137) );
  NAND2_X1 U8702 ( .A1(n8620), .A2(n9966), .ZN(n8128) );
  INV_X1 U8703 ( .A(n9919), .ZN(n7075) );
  NAND2_X1 U8704 ( .A1(n9926), .A2(n7075), .ZN(n7077) );
  NAND2_X1 U8705 ( .A1(n7074), .A2(n9966), .ZN(n7076) );
  NAND2_X1 U8706 ( .A1(n7077), .A2(n7076), .ZN(n7128) );
  NAND2_X1 U8707 ( .A1(n8619), .A2(n7531), .ZN(n8129) );
  NAND2_X1 U8708 ( .A1(n4860), .A2(n8129), .ZN(n8095) );
  NAND2_X1 U8709 ( .A1(n7128), .A2(n8095), .ZN(n7130) );
  INV_X1 U8710 ( .A(n8619), .ZN(n8480) );
  NAND2_X1 U8711 ( .A1(n8480), .A2(n7531), .ZN(n7078) );
  NAND2_X1 U8712 ( .A1(n7130), .A2(n7078), .ZN(n7080) );
  NAND2_X1 U8713 ( .A1(n7079), .A2(n7661), .ZN(n8142) );
  INV_X1 U8714 ( .A(n7079), .ZN(n8618) );
  NAND2_X1 U8715 ( .A1(n8142), .A2(n8126), .ZN(n8091) );
  OAI21_X1 U8716 ( .B1(n7080), .B2(n8091), .A(n7569), .ZN(n7662) );
  INV_X1 U8717 ( .A(n7662), .ZN(n7093) );
  NAND2_X1 U8718 ( .A1(n7081), .A2(n8134), .ZN(n7620) );
  INV_X1 U8719 ( .A(n7620), .ZN(n7083) );
  INV_X1 U8720 ( .A(n7612), .ZN(n7082) );
  NAND2_X1 U8721 ( .A1(n7083), .A2(n7082), .ZN(n7618) );
  AND2_X1 U8722 ( .A1(n9918), .A2(n8137), .ZN(n7084) );
  NAND2_X1 U8723 ( .A1(n7618), .A2(n7084), .ZN(n7086) );
  NAND2_X1 U8724 ( .A1(n7086), .A2(n7085), .ZN(n7131) );
  NAND2_X1 U8725 ( .A1(n7131), .A2(n4860), .ZN(n7133) );
  XNOR2_X1 U8726 ( .A(n7570), .B(n8091), .ZN(n7089) );
  OR2_X1 U8727 ( .A1(n7727), .A2(n8907), .ZN(n7088) );
  NAND2_X1 U8728 ( .A1(n8619), .A2(n8861), .ZN(n7087) );
  NAND2_X1 U8729 ( .A1(n7088), .A2(n7087), .ZN(n7338) );
  AOI21_X1 U8730 ( .B1(n7089), .B2(n9922), .A(n7338), .ZN(n7669) );
  NAND2_X1 U8731 ( .A1(n9927), .A2(n9966), .ZN(n9928) );
  INV_X1 U8732 ( .A(n7531), .ZN(n7140) );
  NAND2_X1 U8733 ( .A1(n7138), .A2(n7661), .ZN(n7090) );
  NAND2_X1 U8734 ( .A1(n7090), .A2(n9913), .ZN(n7091) );
  NOR2_X1 U8735 ( .A1(n7574), .A2(n7091), .ZN(n7664) );
  AOI21_X1 U8736 ( .B1(n9016), .B2(n7661), .A(n7664), .ZN(n7092) );
  OAI211_X1 U8737 ( .C1(n10001), .C2(n7093), .A(n7669), .B(n7092), .ZN(n7096)
         );
  NAND2_X1 U8738 ( .A1(n7096), .A2(n10028), .ZN(n7094) );
  OAI21_X1 U8739 ( .B1(n10028), .B2(n7095), .A(n7094), .ZN(P2_U3466) );
  NAND2_X1 U8740 ( .A1(n7096), .A2(n10045), .ZN(n7097) );
  OAI21_X1 U8741 ( .B1(n10045), .B2(n6253), .A(n7097), .ZN(P2_U3525) );
  OAI21_X1 U8742 ( .B1(n7148), .B2(n4374), .A(n7164), .ZN(n7100) );
  INV_X1 U8743 ( .A(n8315), .ZN(n9157) );
  AOI222_X1 U8744 ( .A1(n9786), .A2(n7100), .B1(n9157), .B2(n9736), .C1(n9158), 
        .C2(n9734), .ZN(n9848) );
  INV_X1 U8745 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7101) );
  OAI22_X1 U8746 ( .A1(n9797), .A2(n7101), .B1(n8312), .B2(n9792), .ZN(n7105)
         );
  NAND2_X1 U8747 ( .A1(n7254), .A2(n7255), .ZN(n7295) );
  INV_X1 U8748 ( .A(n9731), .ZN(n7102) );
  OAI211_X1 U8749 ( .C1(n7102), .C2(n9849), .A(n9857), .B(n7185), .ZN(n9847)
         );
  NOR2_X1 U8750 ( .A1(n7103), .A2(n9757), .ZN(n9575) );
  INV_X1 U8751 ( .A(n9575), .ZN(n7831) );
  NOR2_X1 U8752 ( .A1(n9847), .A2(n7831), .ZN(n7104) );
  AOI211_X1 U8753 ( .C1(n9569), .C2(n7106), .A(n7105), .B(n7104), .ZN(n7127)
         );
  NAND2_X1 U8754 ( .A1(n6305), .A2(n9162), .ZN(n7107) );
  NAND2_X1 U8755 ( .A1(n7108), .A2(n7107), .ZN(n7243) );
  INV_X1 U8756 ( .A(n7243), .ZN(n7110) );
  NAND2_X1 U8757 ( .A1(n7255), .A2(n6307), .ZN(n7111) );
  NAND2_X1 U8758 ( .A1(n7245), .A2(n7111), .ZN(n7287) );
  NAND2_X1 U8759 ( .A1(n7287), .A2(n7112), .ZN(n7114) );
  NAND2_X1 U8760 ( .A1(n9823), .A2(n9783), .ZN(n7113) );
  NAND2_X1 U8761 ( .A1(n7114), .A2(n7113), .ZN(n9771) );
  NAND2_X1 U8762 ( .A1(n7115), .A2(n9761), .ZN(n9780) );
  NOR2_X1 U8763 ( .A1(n7116), .A2(n9159), .ZN(n7117) );
  AOI21_X1 U8764 ( .B1(n9771), .B2(n9780), .A(n7117), .ZN(n9749) );
  NAND2_X1 U8765 ( .A1(n7119), .A2(n7118), .ZN(n9760) );
  NAND2_X1 U8766 ( .A1(n9749), .A2(n9760), .ZN(n7121) );
  NAND2_X1 U8767 ( .A1(n9752), .A2(n9733), .ZN(n7120) );
  NAND2_X1 U8768 ( .A1(n7121), .A2(n7120), .ZN(n9729) );
  NOR2_X1 U8769 ( .A1(n9729), .A2(n9738), .ZN(n7155) );
  INV_X1 U8770 ( .A(n7155), .ZN(n9730) );
  NAND2_X1 U8771 ( .A1(n9841), .A2(n5181), .ZN(n7146) );
  NAND2_X1 U8772 ( .A1(n9730), .A2(n7146), .ZN(n7122) );
  XNOR2_X1 U8773 ( .A(n7123), .B(n7122), .ZN(n9851) );
  INV_X1 U8774 ( .A(n9387), .ZN(n8042) );
  NAND2_X1 U8775 ( .A1(n9851), .A2(n8042), .ZN(n7126) );
  OAI211_X1 U8776 ( .C1(n9568), .C2(n9848), .A(n7127), .B(n7126), .ZN(P1_U3284) );
  OR2_X1 U8777 ( .A1(n7128), .A2(n8095), .ZN(n7129) );
  AND2_X1 U8778 ( .A1(n7130), .A2(n7129), .ZN(n7530) );
  INV_X1 U8779 ( .A(n8129), .ZN(n7132) );
  NOR2_X1 U8780 ( .A1(n7133), .A2(n7132), .ZN(n7134) );
  AOI211_X1 U8781 ( .C1(n8095), .C2(n7135), .A(n8920), .B(n7134), .ZN(n7137)
         );
  NOR2_X1 U8782 ( .A1(n7137), .A2(n7136), .ZN(n7526) );
  INV_X1 U8783 ( .A(n7138), .ZN(n7139) );
  AOI211_X1 U8784 ( .C1(n7140), .C2(n9928), .A(n10004), .B(n7139), .ZN(n7523)
         );
  AOI21_X1 U8785 ( .B1(n9016), .B2(n7140), .A(n7523), .ZN(n7141) );
  OAI211_X1 U8786 ( .C1(n10001), .C2(n7530), .A(n7526), .B(n7141), .ZN(n7143)
         );
  NAND2_X1 U8787 ( .A1(n7143), .A2(n10045), .ZN(n7142) );
  OAI21_X1 U8788 ( .B1(n10045), .B2(n6257), .A(n7142), .ZN(P2_U3524) );
  INV_X1 U8789 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n7145) );
  NAND2_X1 U8790 ( .A1(n7143), .A2(n10028), .ZN(n7144) );
  OAI21_X1 U8791 ( .B1(n10028), .B2(n7145), .A(n7144), .ZN(P2_U3463) );
  NAND2_X1 U8792 ( .A1(n9849), .A2(n7315), .ZN(n7147) );
  AND2_X1 U8793 ( .A1(n7146), .A2(n7147), .ZN(n7191) );
  INV_X1 U8794 ( .A(n7194), .ZN(n7149) );
  AND2_X1 U8795 ( .A1(n7191), .A2(n7149), .ZN(n7189) );
  NAND2_X1 U8796 ( .A1(n9864), .A2(n7207), .ZN(n7152) );
  NAND2_X1 U8797 ( .A1(n7189), .A2(n7152), .ZN(n7154) );
  INV_X1 U8798 ( .A(n7193), .ZN(n7150) );
  NAND2_X1 U8799 ( .A1(n6314), .A2(n9157), .ZN(n7151) );
  INV_X1 U8800 ( .A(n7207), .ZN(n9156) );
  OAI21_X1 U8801 ( .B1(n7155), .B2(n7154), .A(n7153), .ZN(n7200) );
  OR2_X1 U8802 ( .A1(n7503), .A2(n9155), .ZN(n7157) );
  XNOR2_X1 U8803 ( .A(n7548), .B(n7170), .ZN(n9473) );
  INV_X1 U8804 ( .A(n7503), .ZN(n7214) );
  NAND2_X1 U8805 ( .A1(n7331), .A2(n7214), .ZN(n7208) );
  AOI21_X1 U8806 ( .B1(n7208), .B2(n9470), .A(n9865), .ZN(n7158) );
  AND2_X1 U8807 ( .A1(n7158), .A2(n9570), .ZN(n9469) );
  NAND2_X1 U8808 ( .A1(n9569), .A2(n9470), .ZN(n7161) );
  INV_X1 U8809 ( .A(n9792), .ZN(n9755) );
  INV_X1 U8810 ( .A(n7159), .ZN(n7636) );
  NAND2_X1 U8811 ( .A1(n9755), .A2(n7636), .ZN(n7160) );
  OAI211_X1 U8812 ( .C1(n9797), .C2(n6772), .A(n7161), .B(n7160), .ZN(n7162)
         );
  AOI21_X1 U8813 ( .B1(n9469), .B2(n9350), .A(n7162), .ZN(n7175) );
  NAND2_X1 U8814 ( .A1(n7164), .A2(n7163), .ZN(n7183) );
  NAND2_X1 U8815 ( .A1(n7183), .A2(n7194), .ZN(n7166) );
  NAND2_X1 U8816 ( .A1(n7166), .A2(n7165), .ZN(n7324) );
  NAND2_X1 U8817 ( .A1(n7324), .A2(n7167), .ZN(n7169) );
  NAND2_X1 U8818 ( .A1(n7169), .A2(n7168), .ZN(n7552) );
  XNOR2_X1 U8819 ( .A(n7552), .B(n7170), .ZN(n7171) );
  NAND2_X1 U8820 ( .A1(n7171), .A2(n9786), .ZN(n7173) );
  INV_X1 U8821 ( .A(n7674), .ZN(n9154) );
  AOI22_X1 U8822 ( .A1(n9736), .A2(n9154), .B1(n9734), .B2(n9155), .ZN(n7172)
         );
  NAND2_X1 U8823 ( .A1(n7173), .A2(n7172), .ZN(n9468) );
  NAND2_X1 U8824 ( .A1(n9468), .A2(n9797), .ZN(n7174) );
  OAI211_X1 U8825 ( .C1(n9473), .C2(n9387), .A(n7175), .B(n7174), .ZN(P1_U3280) );
  INV_X1 U8826 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n7182) );
  OAI21_X1 U8827 ( .B1(n9777), .B2(n9569), .A(n7176), .ZN(n7181) );
  OAI21_X1 U8828 ( .B1(n7178), .B2(n9792), .A(n7177), .ZN(n7179) );
  NAND2_X1 U8829 ( .A1(n7179), .A2(n9797), .ZN(n7180) );
  OAI211_X1 U8830 ( .C1(n7182), .C2(n9797), .A(n7181), .B(n7180), .ZN(P1_U3291) );
  XNOR2_X1 U8831 ( .A(n7194), .B(n7183), .ZN(n7184) );
  AOI222_X1 U8832 ( .A1(n9786), .A2(n7184), .B1(n9735), .B2(n9734), .C1(n9156), 
        .C2(n9736), .ZN(n9860) );
  AOI21_X1 U8833 ( .B1(n6314), .B2(n7185), .A(n7329), .ZN(n9858) );
  INV_X1 U8834 ( .A(n7186), .ZN(n7311) );
  AOI22_X1 U8835 ( .A1(n9568), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n7311), .B2(
        n9755), .ZN(n7187) );
  OAI21_X1 U8836 ( .B1(n9791), .B2(n4574), .A(n7187), .ZN(n7188) );
  AOI21_X1 U8837 ( .B1(n9858), .B2(n9777), .A(n7188), .ZN(n7197) );
  NAND2_X1 U8838 ( .A1(n9730), .A2(n7189), .ZN(n7321) );
  AND2_X1 U8839 ( .A1(n7190), .A2(n7321), .ZN(n9855) );
  NAND2_X1 U8840 ( .A1(n9730), .A2(n7191), .ZN(n7192) );
  AND2_X1 U8841 ( .A1(n7193), .A2(n7192), .ZN(n7195) );
  NAND2_X1 U8842 ( .A1(n7195), .A2(n7194), .ZN(n9854) );
  NAND3_X1 U8843 ( .A1(n9855), .A2(n9854), .A3(n8042), .ZN(n7196) );
  OAI211_X1 U8844 ( .C1(n9860), .C2(n9568), .A(n7197), .B(n7196), .ZN(P1_U3283) );
  INV_X1 U8845 ( .A(n7198), .ZN(n7199) );
  AOI21_X1 U8846 ( .B1(n7204), .B2(n7200), .A(n7199), .ZN(n7505) );
  INV_X1 U8847 ( .A(n7201), .ZN(n7203) );
  OAI21_X1 U8848 ( .B1(n7324), .B2(n7203), .A(n7202), .ZN(n7205) );
  XNOR2_X1 U8849 ( .A(n7205), .B(n7204), .ZN(n7206) );
  OAI222_X1 U8850 ( .A1(n9781), .A2(n7655), .B1(n9784), .B2(n7207), .C1(n7206), 
        .C2(n9766), .ZN(n7502) );
  INV_X1 U8851 ( .A(n7331), .ZN(n7210) );
  INV_X1 U8852 ( .A(n7208), .ZN(n7209) );
  AOI211_X1 U8853 ( .C1(n7503), .C2(n7210), .A(n9865), .B(n7209), .ZN(n7501)
         );
  NAND2_X1 U8854 ( .A1(n7501), .A2(n9575), .ZN(n7213) );
  INV_X1 U8855 ( .A(n7211), .ZN(n7267) );
  AOI22_X1 U8856 ( .A1(n9568), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n7267), .B2(
        n9755), .ZN(n7212) );
  OAI211_X1 U8857 ( .C1(n7214), .C2(n9791), .A(n7213), .B(n7212), .ZN(n7215)
         );
  AOI21_X1 U8858 ( .B1(n9797), .B2(n7502), .A(n7215), .ZN(n7216) );
  OAI21_X1 U8859 ( .B1(n7505), .B2(n9387), .A(n7216), .ZN(P1_U3281) );
  INV_X1 U8860 ( .A(n7217), .ZN(n7221) );
  AND2_X1 U8861 ( .A1(n6886), .A2(n7218), .ZN(n7219) );
  NAND2_X1 U8862 ( .A1(n7219), .A2(n5204), .ZN(n7275) );
  OAI21_X1 U8863 ( .B1(n7219), .B2(n5204), .A(n7275), .ZN(n7220) );
  NOR2_X1 U8864 ( .A1(n7220), .A2(n7221), .ZN(n7277) );
  AOI21_X1 U8865 ( .B1(n7221), .B2(n7220), .A(n7277), .ZN(n7228) );
  OAI22_X1 U8866 ( .A1(n9836), .A2(n9148), .B1(n9114), .B2(n9767), .ZN(n7224)
         );
  OAI21_X1 U8867 ( .B1(n9123), .B2(n5181), .A(n7222), .ZN(n7223) );
  NOR2_X1 U8868 ( .A1(n7224), .A2(n7223), .ZN(n7227) );
  INV_X1 U8869 ( .A(n7225), .ZN(n9754) );
  NAND2_X1 U8870 ( .A1(n9140), .A2(n9754), .ZN(n7226) );
  OAI211_X1 U8871 ( .C1(n7228), .C2(n9131), .A(n7227), .B(n7226), .ZN(P1_U3225) );
  INV_X1 U8872 ( .A(n7351), .ZN(n7229) );
  OAI222_X1 U8873 ( .A1(n9502), .A2(n7230), .B1(n4282), .B2(n7229), .C1(
        P1_U3084), .C2(n9298), .ZN(P1_U3334) );
  XNOR2_X1 U8874 ( .A(n7232), .B(n7231), .ZN(n7242) );
  INV_X1 U8875 ( .A(n9893), .ZN(n9522) );
  INV_X1 U8876 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7238) );
  OAI21_X1 U8877 ( .B1(n7235), .B2(n7234), .A(n7233), .ZN(n7236) );
  NAND2_X1 U8878 ( .A1(n9888), .A2(n7236), .ZN(n7237) );
  NAND2_X1 U8879 ( .A1(P2_U3152), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n7905) );
  OAI211_X1 U8880 ( .C1(n7749), .C2(n7238), .A(n7237), .B(n7905), .ZN(n7239)
         );
  AOI21_X1 U8881 ( .B1(n7240), .B2(n9522), .A(n7239), .ZN(n7241) );
  OAI21_X1 U8882 ( .B1(n7242), .B2(n9895), .A(n7241), .ZN(P2_U3257) );
  NAND2_X1 U8883 ( .A1(n7243), .A2(n7248), .ZN(n7244) );
  NAND2_X1 U8884 ( .A1(n7245), .A2(n7244), .ZN(n7253) );
  INV_X1 U8885 ( .A(n9789), .ZN(n9565) );
  NAND2_X1 U8886 ( .A1(n7253), .A2(n9565), .ZN(n7252) );
  OAI21_X1 U8887 ( .B1(n7248), .B2(n7247), .A(n7246), .ZN(n7249) );
  NAND2_X1 U8888 ( .A1(n7249), .A2(n9786), .ZN(n7251) );
  AOI22_X1 U8889 ( .A1(n9736), .A2(n9160), .B1(n9734), .B2(n9162), .ZN(n7250)
         );
  NAND3_X1 U8890 ( .A1(n7252), .A2(n7251), .A3(n7250), .ZN(n9820) );
  MUX2_X1 U8891 ( .A(n9820), .B(P1_REG2_REG_2__SCAN_IN), .S(n9568), .Z(n7260)
         );
  INV_X1 U8892 ( .A(n7253), .ZN(n9819) );
  OR2_X1 U8893 ( .A1(n7255), .A2(n7254), .ZN(n7256) );
  AND2_X1 U8894 ( .A1(n7256), .A2(n7295), .ZN(n9816) );
  NAND2_X1 U8895 ( .A1(n9777), .A2(n9816), .ZN(n7258) );
  AOI22_X1 U8896 ( .A1(n9569), .A2(n9815), .B1(n9755), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n7257) );
  OAI211_X1 U8897 ( .C1(n9819), .C2(n7337), .A(n7258), .B(n7257), .ZN(n7259)
         );
  OR2_X1 U8898 ( .A1(n7260), .A2(n7259), .ZN(P1_U3289) );
  AND2_X1 U8899 ( .A1(n7262), .A2(n7261), .ZN(n7266) );
  NAND2_X1 U8900 ( .A1(n7264), .A2(n7263), .ZN(n7265) );
  XNOR2_X1 U8901 ( .A(n7266), .B(n7265), .ZN(n7273) );
  NAND2_X1 U8902 ( .A1(n9140), .A2(n7267), .ZN(n7270) );
  NOR2_X1 U8903 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7268), .ZN(n8346) );
  AOI21_X1 U8904 ( .B1(n9139), .B2(n9156), .A(n8346), .ZN(n7269) );
  OAI211_X1 U8905 ( .C1(n7655), .C2(n9123), .A(n7270), .B(n7269), .ZN(n7271)
         );
  AOI21_X1 U8906 ( .B1(n7503), .B2(n9129), .A(n7271), .ZN(n7272) );
  OAI21_X1 U8907 ( .B1(n7273), .B2(n9131), .A(n7272), .ZN(P1_U3215) );
  INV_X1 U8908 ( .A(n7275), .ZN(n7276) );
  NOR3_X1 U8909 ( .A1(n7277), .A2(n5201), .A3(n7276), .ZN(n7280) );
  OAI21_X1 U8910 ( .B1(n7280), .B2(n4373), .A(n9136), .ZN(n7286) );
  NOR2_X1 U8911 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7281), .ZN(n9624) );
  AOI21_X1 U8912 ( .B1(n9139), .B2(n9733), .A(n9624), .ZN(n7282) );
  OAI21_X1 U8913 ( .B1(n7315), .B2(n9123), .A(n7282), .ZN(n7283) );
  AOI21_X1 U8914 ( .B1(n7284), .B2(n9129), .A(n7283), .ZN(n7285) );
  OAI211_X1 U8915 ( .C1(n9127), .C2(n9743), .A(n7286), .B(n7285), .ZN(P1_U3237) );
  XNOR2_X1 U8916 ( .A(n7287), .B(n7288), .ZN(n7293) );
  XNOR2_X1 U8917 ( .A(n7289), .B(n7288), .ZN(n7291) );
  OAI22_X1 U8918 ( .A1(n9784), .A2(n6307), .B1(n9767), .B2(n9781), .ZN(n7290)
         );
  AOI21_X1 U8919 ( .B1(n7291), .B2(n9786), .A(n7290), .ZN(n7292) );
  OAI21_X1 U8920 ( .B1(n7293), .B2(n9789), .A(n7292), .ZN(n9825) );
  INV_X1 U8921 ( .A(n9825), .ZN(n7303) );
  INV_X1 U8922 ( .A(n7293), .ZN(n9827) );
  NAND2_X1 U8923 ( .A1(n7295), .A2(n7294), .ZN(n7296) );
  NAND2_X1 U8924 ( .A1(n9772), .A2(n7296), .ZN(n9824) );
  INV_X1 U8925 ( .A(n9824), .ZN(n7297) );
  NAND2_X1 U8926 ( .A1(n9777), .A2(n7297), .ZN(n7300) );
  AOI22_X1 U8927 ( .A1(n9383), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n9755), .B2(
        n7298), .ZN(n7299) );
  OAI211_X1 U8928 ( .C1(n9823), .C2(n9791), .A(n7300), .B(n7299), .ZN(n7301)
         );
  AOI21_X1 U8929 ( .B1(n9778), .B2(n9827), .A(n7301), .ZN(n7302) );
  OAI21_X1 U8930 ( .B1(n9568), .B2(n7303), .A(n7302), .ZN(P1_U3288) );
  INV_X1 U8931 ( .A(n7481), .ZN(n7310) );
  NAND2_X1 U8932 ( .A1(n8309), .A2(n7304), .ZN(n7306) );
  NAND2_X1 U8933 ( .A1(n7306), .A2(n7305), .ZN(n7480) );
  OR2_X1 U8934 ( .A1(n7306), .A2(n7305), .ZN(n7308) );
  AOI21_X1 U8935 ( .B1(n7308), .B2(n7480), .A(n7307), .ZN(n7309) );
  AOI21_X1 U8936 ( .B1(n7310), .B2(n7480), .A(n7309), .ZN(n7318) );
  NAND2_X1 U8937 ( .A1(n9140), .A2(n7311), .ZN(n7314) );
  AOI21_X1 U8938 ( .B1(n9145), .B2(n9156), .A(n7312), .ZN(n7313) );
  OAI211_X1 U8939 ( .C1(n7315), .C2(n9114), .A(n7314), .B(n7313), .ZN(n7316)
         );
  AOI21_X1 U8940 ( .B1(n6314), .B2(n9129), .A(n7316), .ZN(n7317) );
  OAI21_X1 U8941 ( .B1(n7318), .B2(n9131), .A(n7317), .ZN(P1_U3219) );
  INV_X1 U8942 ( .A(n7319), .ZN(n7320) );
  NAND2_X1 U8943 ( .A1(n7321), .A2(n7320), .ZN(n7322) );
  XNOR2_X1 U8944 ( .A(n7322), .B(n7323), .ZN(n9862) );
  XOR2_X1 U8945 ( .A(n7324), .B(n7323), .Z(n7326) );
  OAI22_X1 U8946 ( .A1(n9784), .A2(n8315), .B1(n7490), .B2(n9781), .ZN(n7325)
         );
  AOI21_X1 U8947 ( .B1(n7326), .B2(n9786), .A(n7325), .ZN(n7327) );
  OAI21_X1 U8948 ( .B1(n9862), .B2(n9789), .A(n7327), .ZN(n9867) );
  NAND2_X1 U8949 ( .A1(n9867), .A2(n9797), .ZN(n7336) );
  INV_X1 U8950 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n7328) );
  OAI22_X1 U8951 ( .A1(n9797), .A2(n7328), .B1(n7486), .B2(n9792), .ZN(n7333)
         );
  NOR2_X1 U8952 ( .A1(n7329), .A2(n9864), .ZN(n7330) );
  OR2_X1 U8953 ( .A1(n7331), .A2(n7330), .ZN(n9866) );
  INV_X1 U8954 ( .A(n9777), .ZN(n9251) );
  NOR2_X1 U8955 ( .A1(n9866), .A2(n9251), .ZN(n7332) );
  AOI211_X1 U8956 ( .C1(n9569), .C2(n7334), .A(n7333), .B(n7332), .ZN(n7335)
         );
  OAI211_X1 U8957 ( .C1(n9862), .C2(n7337), .A(n7336), .B(n7335), .ZN(P1_U3282) );
  NAND2_X1 U8958 ( .A1(n8589), .A2(n7661), .ZN(n7340) );
  NAND2_X1 U8959 ( .A1(n8509), .A2(n7338), .ZN(n7339) );
  OAI211_X1 U8960 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n7341), .A(n7340), .B(n7339), .ZN(n7348) );
  AOI22_X1 U8961 ( .A1(n8514), .A2(n8619), .B1(n8488), .B2(n7342), .ZN(n7346)
         );
  INV_X1 U8962 ( .A(n7343), .ZN(n7345) );
  NOR3_X1 U8963 ( .A1(n7346), .A2(n7345), .A3(n7344), .ZN(n7347) );
  AOI211_X1 U8964 ( .C1(n8601), .C2(n7663), .A(n7348), .B(n7347), .ZN(n7349)
         );
  OAI21_X1 U8965 ( .B1(n8402), .B2(n8593), .A(n7349), .ZN(P2_U3229) );
  AOI222_X1 U8966 ( .A1(n7351), .A2(n9044), .B1(P1_DATAO_REG_19__SCAN_IN), 
        .B2(n7350), .C1(n4284), .C2(P2_STATE_REG_SCAN_IN), .ZN(n7479) );
  NAND4_X1 U8967 ( .A1(keyinput29), .A2(keyinput33), .A3(keyinput21), .A4(
        keyinput49), .ZN(n7355) );
  NAND4_X1 U8968 ( .A1(keyinput41), .A2(keyinput61), .A3(keyinput20), .A4(
        keyinput4), .ZN(n7354) );
  NAND4_X1 U8969 ( .A1(keyinput16), .A2(keyinput28), .A3(keyinput60), .A4(
        keyinput58), .ZN(n7353) );
  NAND4_X1 U8970 ( .A1(keyinput50), .A2(keyinput55), .A3(keyinput30), .A4(
        keyinput19), .ZN(n7352) );
  NOR4_X1 U8971 ( .A1(n7355), .A2(n7354), .A3(n7353), .A4(n7352), .ZN(n7477)
         );
  NAND4_X1 U8972 ( .A1(keyinput27), .A2(keyinput14), .A3(keyinput42), .A4(
        keyinput40), .ZN(n7375) );
  NAND2_X1 U8973 ( .A1(keyinput51), .A2(keyinput31), .ZN(n7356) );
  NOR3_X1 U8974 ( .A1(keyinput2), .A2(keyinput24), .A3(n7356), .ZN(n7360) );
  NOR3_X1 U8975 ( .A1(keyinput46), .A2(keyinput62), .A3(keyinput3), .ZN(n7359)
         );
  NAND2_X1 U8976 ( .A1(keyinput63), .A2(keyinput18), .ZN(n7357) );
  NOR3_X1 U8977 ( .A1(keyinput59), .A2(keyinput38), .A3(n7357), .ZN(n7358) );
  NAND4_X1 U8978 ( .A1(n7360), .A2(keyinput10), .A3(n7359), .A4(n7358), .ZN(
        n7374) );
  NOR3_X1 U8979 ( .A1(keyinput1), .A2(keyinput11), .A3(keyinput7), .ZN(n7366)
         );
  NOR4_X1 U8980 ( .A1(keyinput39), .A2(keyinput37), .A3(keyinput44), .A4(
        keyinput25), .ZN(n7365) );
  NAND3_X1 U8981 ( .A1(keyinput43), .A2(keyinput22), .A3(keyinput23), .ZN(
        n7363) );
  INV_X1 U8982 ( .A(keyinput56), .ZN(n7361) );
  NAND3_X1 U8983 ( .A1(keyinput32), .A2(keyinput6), .A3(n7361), .ZN(n7362) );
  NOR4_X1 U8984 ( .A1(keyinput48), .A2(keyinput45), .A3(n7363), .A4(n7362), 
        .ZN(n7364) );
  NAND4_X1 U8985 ( .A1(keyinput12), .A2(n7366), .A3(n7365), .A4(n7364), .ZN(
        n7373) );
  NOR4_X1 U8986 ( .A1(keyinput13), .A2(keyinput5), .A3(keyinput17), .A4(
        keyinput53), .ZN(n7371) );
  NOR4_X1 U8987 ( .A1(keyinput57), .A2(keyinput8), .A3(keyinput36), .A4(
        keyinput52), .ZN(n7370) );
  NOR4_X1 U8988 ( .A1(keyinput0), .A2(keyinput47), .A3(keyinput34), .A4(
        keyinput35), .ZN(n7369) );
  INV_X1 U8989 ( .A(keyinput9), .ZN(n7367) );
  NOR4_X1 U8990 ( .A1(keyinput54), .A2(keyinput15), .A3(keyinput26), .A4(n7367), .ZN(n7368) );
  NAND4_X1 U8991 ( .A1(n7371), .A2(n7370), .A3(n7369), .A4(n7368), .ZN(n7372)
         );
  NOR4_X1 U8992 ( .A1(n7375), .A2(n7374), .A3(n7373), .A4(n7372), .ZN(n7476)
         );
  INV_X1 U8993 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n9802) );
  INV_X1 U8994 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n8283) );
  AOI22_X1 U8995 ( .A1(n9802), .A2(keyinput31), .B1(keyinput2), .B2(n8283), 
        .ZN(n7376) );
  OAI221_X1 U8996 ( .B1(n9802), .B2(keyinput31), .C1(n8283), .C2(keyinput2), 
        .A(n7376), .ZN(n7385) );
  INV_X1 U8997 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n9828) );
  AOI22_X1 U8998 ( .A1(n8056), .A2(keyinput51), .B1(keyinput24), .B2(n9828), 
        .ZN(n7377) );
  OAI221_X1 U8999 ( .B1(n8056), .B2(keyinput51), .C1(n9828), .C2(keyinput24), 
        .A(n7377), .ZN(n7384) );
  INV_X1 U9000 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n9550) );
  AOI22_X1 U9001 ( .A1(n9550), .A2(keyinput27), .B1(n9940), .B2(keyinput14), 
        .ZN(n7378) );
  OAI221_X1 U9002 ( .B1(n9550), .B2(keyinput27), .C1(n9940), .C2(keyinput14), 
        .A(n7378), .ZN(n7383) );
  INV_X1 U9003 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n7381) );
  INV_X1 U9004 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n7380) );
  AOI22_X1 U9005 ( .A1(n7381), .A2(keyinput42), .B1(keyinput40), .B2(n7380), 
        .ZN(n7379) );
  OAI221_X1 U9006 ( .B1(n7381), .B2(keyinput42), .C1(n7380), .C2(keyinput40), 
        .A(n7379), .ZN(n7382) );
  NOR4_X1 U9007 ( .A1(n7385), .A2(n7384), .A3(n7383), .A4(n7382), .ZN(n7422)
         );
  AOI22_X1 U9008 ( .A1(n10043), .A2(keyinput46), .B1(n7387), .B2(keyinput62), 
        .ZN(n7386) );
  OAI221_X1 U9009 ( .B1(n10043), .B2(keyinput46), .C1(n7387), .C2(keyinput62), 
        .A(n7386), .ZN(n7396) );
  INV_X1 U9010 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n9971) );
  AOI22_X1 U9011 ( .A1(n9971), .A2(keyinput3), .B1(n7757), .B2(keyinput10), 
        .ZN(n7388) );
  OAI221_X1 U9012 ( .B1(n9971), .B2(keyinput3), .C1(n7757), .C2(keyinput10), 
        .A(n7388), .ZN(n7395) );
  INV_X1 U9013 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n7391) );
  INV_X1 U9014 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n7390) );
  AOI22_X1 U9015 ( .A1(n7391), .A2(keyinput59), .B1(n7390), .B2(keyinput18), 
        .ZN(n7389) );
  OAI221_X1 U9016 ( .B1(n7391), .B2(keyinput59), .C1(n7390), .C2(keyinput18), 
        .A(n7389), .ZN(n7394) );
  INV_X1 U9017 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n9803) );
  INV_X1 U9018 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n9804) );
  AOI22_X1 U9019 ( .A1(n9803), .A2(keyinput38), .B1(keyinput63), .B2(n9804), 
        .ZN(n7392) );
  OAI221_X1 U9020 ( .B1(n9803), .B2(keyinput38), .C1(n9804), .C2(keyinput63), 
        .A(n7392), .ZN(n7393) );
  NOR4_X1 U9021 ( .A1(n7396), .A2(n7395), .A3(n7394), .A4(n7393), .ZN(n7421)
         );
  INV_X1 U9022 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10029) );
  INV_X1 U9023 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n7398) );
  AOI22_X1 U9024 ( .A1(n10029), .A2(keyinput48), .B1(n7398), .B2(keyinput43), 
        .ZN(n7397) );
  OAI221_X1 U9025 ( .B1(n10029), .B2(keyinput48), .C1(n7398), .C2(keyinput43), 
        .A(n7397), .ZN(n7409) );
  INV_X1 U9026 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n7400) );
  AOI22_X1 U9027 ( .A1(n7400), .A2(keyinput12), .B1(n6608), .B2(keyinput7), 
        .ZN(n7399) );
  OAI221_X1 U9028 ( .B1(n7400), .B2(keyinput12), .C1(n6608), .C2(keyinput7), 
        .A(n7399), .ZN(n7408) );
  INV_X1 U9029 ( .A(SI_6_), .ZN(n7402) );
  AOI22_X1 U9030 ( .A1(n6257), .A2(keyinput22), .B1(n7402), .B2(keyinput23), 
        .ZN(n7401) );
  OAI221_X1 U9031 ( .B1(n6257), .B2(keyinput22), .C1(n7402), .C2(keyinput23), 
        .A(n7401), .ZN(n7407) );
  INV_X1 U9032 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n7403) );
  XOR2_X1 U9033 ( .A(n7403), .B(keyinput11), .Z(n7405) );
  XNOR2_X1 U9034 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(keyinput1), .ZN(n7404) );
  NAND2_X1 U9035 ( .A1(n7405), .A2(n7404), .ZN(n7406) );
  NOR4_X1 U9036 ( .A1(n7409), .A2(n7408), .A3(n7407), .A4(n7406), .ZN(n7420)
         );
  INV_X1 U9037 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n9805) );
  AOI22_X1 U9038 ( .A1(n9941), .A2(keyinput6), .B1(n9805), .B2(keyinput32), 
        .ZN(n7410) );
  OAI221_X1 U9039 ( .B1(n9941), .B2(keyinput6), .C1(n9805), .C2(keyinput32), 
        .A(n7410), .ZN(n7418) );
  AOI22_X1 U9040 ( .A1(n7946), .A2(keyinput39), .B1(keyinput37), .B2(n4715), 
        .ZN(n7411) );
  OAI221_X1 U9041 ( .B1(n7946), .B2(keyinput39), .C1(n4715), .C2(keyinput37), 
        .A(n7411), .ZN(n7417) );
  INV_X1 U9042 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n9807) );
  AOI22_X1 U9043 ( .A1(n9942), .A2(keyinput44), .B1(n9807), .B2(keyinput25), 
        .ZN(n7412) );
  OAI221_X1 U9044 ( .B1(n9942), .B2(keyinput44), .C1(n9807), .C2(keyinput25), 
        .A(n7412), .ZN(n7416) );
  XNOR2_X1 U9045 ( .A(P2_IR_REG_17__SCAN_IN), .B(keyinput45), .ZN(n7414) );
  XNOR2_X1 U9046 ( .A(P1_REG0_REG_29__SCAN_IN), .B(keyinput56), .ZN(n7413) );
  NAND2_X1 U9047 ( .A1(n7414), .A2(n7413), .ZN(n7415) );
  NOR4_X1 U9048 ( .A1(n7418), .A2(n7417), .A3(n7416), .A4(n7415), .ZN(n7419)
         );
  NAND4_X1 U9049 ( .A1(n7422), .A2(n7421), .A3(n7420), .A4(n7419), .ZN(n7475)
         );
  INV_X1 U9050 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n10082) );
  AOI22_X1 U9051 ( .A1(n9943), .A2(keyinput8), .B1(keyinput30), .B2(n10082), 
        .ZN(n7423) );
  OAI221_X1 U9052 ( .B1(n9943), .B2(keyinput8), .C1(n10082), .C2(keyinput30), 
        .A(n7423), .ZN(n7434) );
  AOI22_X1 U9053 ( .A1(n7425), .A2(keyinput34), .B1(keyinput60), .B2(n6251), 
        .ZN(n7424) );
  OAI221_X1 U9054 ( .B1(n7425), .B2(keyinput34), .C1(n6251), .C2(keyinput60), 
        .A(n7424), .ZN(n7433) );
  INV_X1 U9055 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n7427) );
  AOI22_X1 U9056 ( .A1(n7428), .A2(keyinput36), .B1(keyinput61), .B2(n7427), 
        .ZN(n7426) );
  OAI221_X1 U9057 ( .B1(n7428), .B2(keyinput36), .C1(n7427), .C2(keyinput61), 
        .A(n7426), .ZN(n7432) );
  XNOR2_X1 U9058 ( .A(P2_REG1_REG_30__SCAN_IN), .B(keyinput58), .ZN(n7430) );
  XNOR2_X1 U9059 ( .A(P1_IR_REG_14__SCAN_IN), .B(keyinput53), .ZN(n7429) );
  NAND2_X1 U9060 ( .A1(n7430), .A2(n7429), .ZN(n7431) );
  NOR4_X1 U9061 ( .A1(n7434), .A2(n7433), .A3(n7432), .A4(n7431), .ZN(n7473)
         );
  INV_X1 U9062 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n7436) );
  AOI22_X1 U9063 ( .A1(n7437), .A2(keyinput15), .B1(keyinput21), .B2(n7436), 
        .ZN(n7435) );
  OAI221_X1 U9064 ( .B1(n7437), .B2(keyinput15), .C1(n7436), .C2(keyinput21), 
        .A(n7435), .ZN(n7446) );
  INV_X1 U9065 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n8298) );
  AOI22_X1 U9066 ( .A1(n8298), .A2(keyinput52), .B1(n9104), .B2(keyinput20), 
        .ZN(n7438) );
  OAI221_X1 U9067 ( .B1(n8298), .B2(keyinput52), .C1(n9104), .C2(keyinput20), 
        .A(n7438), .ZN(n7445) );
  INV_X1 U9068 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7441) );
  AOI22_X1 U9069 ( .A1(n7441), .A2(keyinput17), .B1(n7440), .B2(keyinput26), 
        .ZN(n7439) );
  OAI221_X1 U9070 ( .B1(n7441), .B2(keyinput17), .C1(n7440), .C2(keyinput26), 
        .A(n7439), .ZN(n7444) );
  INV_X1 U9071 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n9668) );
  AOI22_X1 U9072 ( .A1(n9668), .A2(keyinput29), .B1(P2_U3152), .B2(keyinput19), 
        .ZN(n7442) );
  OAI221_X1 U9073 ( .B1(n9668), .B2(keyinput29), .C1(P2_U3152), .C2(keyinput19), .A(n7442), .ZN(n7443) );
  NOR4_X1 U9074 ( .A1(n7446), .A2(n7445), .A3(n7444), .A4(n7443), .ZN(n7472)
         );
  INV_X1 U9075 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n9800) );
  INV_X1 U9076 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9709) );
  AOI22_X1 U9077 ( .A1(n9800), .A2(keyinput47), .B1(keyinput16), .B2(n9709), 
        .ZN(n7447) );
  OAI221_X1 U9078 ( .B1(n9800), .B2(keyinput47), .C1(n9709), .C2(keyinput16), 
        .A(n7447), .ZN(n7456) );
  INV_X1 U9079 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7449) );
  AOI22_X1 U9080 ( .A1(n7450), .A2(keyinput0), .B1(keyinput54), .B2(n7449), 
        .ZN(n7448) );
  OAI221_X1 U9081 ( .B1(n7450), .B2(keyinput0), .C1(n7449), .C2(keyinput54), 
        .A(n7448), .ZN(n7455) );
  INV_X1 U9082 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n9598) );
  INV_X1 U9083 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n9806) );
  AOI22_X1 U9084 ( .A1(n9598), .A2(keyinput4), .B1(n9806), .B2(keyinput55), 
        .ZN(n7451) );
  OAI221_X1 U9085 ( .B1(n9598), .B2(keyinput4), .C1(n9806), .C2(keyinput55), 
        .A(n7451), .ZN(n7454) );
  AOI22_X1 U9086 ( .A1(n6255), .A2(keyinput13), .B1(n5652), .B2(keyinput57), 
        .ZN(n7452) );
  OAI221_X1 U9087 ( .B1(n6255), .B2(keyinput13), .C1(n5652), .C2(keyinput57), 
        .A(n7452), .ZN(n7453) );
  NOR4_X1 U9088 ( .A1(n7456), .A2(n7455), .A3(n7454), .A4(n7453), .ZN(n7471)
         );
  INV_X1 U9089 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n9801) );
  AOI22_X1 U9090 ( .A1(n9801), .A2(keyinput33), .B1(keyinput50), .B2(n5328), 
        .ZN(n7457) );
  OAI221_X1 U9091 ( .B1(n9801), .B2(keyinput33), .C1(n5328), .C2(keyinput50), 
        .A(n7457), .ZN(n7469) );
  INV_X1 U9092 ( .A(keyinput28), .ZN(n7459) );
  AOI22_X1 U9093 ( .A1(n7460), .A2(keyinput5), .B1(P1_WR_REG_SCAN_IN), .B2(
        n7459), .ZN(n7458) );
  OAI221_X1 U9094 ( .B1(n7460), .B2(keyinput5), .C1(n7459), .C2(
        P1_WR_REG_SCAN_IN), .A(n7458), .ZN(n7468) );
  INV_X1 U9095 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7463) );
  AOI22_X1 U9096 ( .A1(n7463), .A2(keyinput9), .B1(n7462), .B2(keyinput41), 
        .ZN(n7461) );
  OAI221_X1 U9097 ( .B1(n7463), .B2(keyinput9), .C1(n7462), .C2(keyinput41), 
        .A(n7461), .ZN(n7467) );
  XNOR2_X1 U9098 ( .A(P1_REG3_REG_6__SCAN_IN), .B(keyinput49), .ZN(n7465) );
  XNOR2_X1 U9099 ( .A(P1_IR_REG_0__SCAN_IN), .B(keyinput35), .ZN(n7464) );
  NAND2_X1 U9100 ( .A1(n7465), .A2(n7464), .ZN(n7466) );
  NOR4_X1 U9101 ( .A1(n7469), .A2(n7468), .A3(n7467), .A4(n7466), .ZN(n7470)
         );
  NAND4_X1 U9102 ( .A1(n7473), .A2(n7472), .A3(n7471), .A4(n7470), .ZN(n7474)
         );
  AOI211_X1 U9103 ( .C1(n7477), .C2(n7476), .A(n7475), .B(n7474), .ZN(n7478)
         );
  XNOR2_X1 U9104 ( .A(n7479), .B(n7478), .ZN(P2_U3339) );
  NAND2_X1 U9105 ( .A1(n7481), .A2(n7480), .ZN(n7483) );
  NAND2_X1 U9106 ( .A1(n7483), .A2(n7484), .ZN(n7482) );
  OAI21_X1 U9107 ( .B1(n7484), .B2(n7483), .A(n7482), .ZN(n7485) );
  NAND2_X1 U9108 ( .A1(n7485), .A2(n9136), .ZN(n7494) );
  INV_X1 U9109 ( .A(n7486), .ZN(n7492) );
  OR2_X1 U9110 ( .A1(n9114), .A2(n8315), .ZN(n7489) );
  INV_X1 U9111 ( .A(n7487), .ZN(n7488) );
  OAI211_X1 U9112 ( .C1(n7490), .C2(n9123), .A(n7489), .B(n7488), .ZN(n7491)
         );
  AOI21_X1 U9113 ( .B1(n7492), .B2(n9140), .A(n7491), .ZN(n7493) );
  OAI211_X1 U9114 ( .C1(n9864), .C2(n9148), .A(n7494), .B(n7493), .ZN(P1_U3229) );
  INV_X1 U9115 ( .A(n7495), .ZN(n8385) );
  OAI222_X1 U9116 ( .A1(n9047), .A2(n7497), .B1(P2_U3152), .B2(n7496), .C1(
        n9049), .C2(n8385), .ZN(P2_U3338) );
  INV_X1 U9117 ( .A(n7498), .ZN(n7510) );
  OAI222_X1 U9118 ( .A1(n9502), .A2(n7500), .B1(n4282), .B2(n7510), .C1(n7499), 
        .C2(P1_U3084), .ZN(P1_U3332) );
  INV_X1 U9119 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n7507) );
  AOI211_X1 U9120 ( .C1(n9856), .C2(n7503), .A(n7502), .B(n7501), .ZN(n7504)
         );
  OAI21_X1 U9121 ( .B1(n7505), .B2(n9472), .A(n7504), .ZN(n7508) );
  NAND2_X1 U9122 ( .A1(n7508), .A2(n9872), .ZN(n7506) );
  OAI21_X1 U9123 ( .B1(n9872), .B2(n7507), .A(n7506), .ZN(P1_U3484) );
  NAND2_X1 U9124 ( .A1(n7508), .A2(n9887), .ZN(n7509) );
  OAI21_X1 U9125 ( .B1(n9887), .B2(n6763), .A(n7509), .ZN(P1_U3533) );
  OAI222_X1 U9126 ( .A1(n9041), .A2(n7511), .B1(P2_U3152), .B2(n8133), .C1(
        n9049), .C2(n7510), .ZN(P2_U3337) );
  INV_X1 U9127 ( .A(n7512), .ZN(n7513) );
  NOR3_X1 U9128 ( .A1(n7514), .A2(n7513), .A3(n9939), .ZN(n7516) );
  AND2_X1 U9129 ( .A1(n7516), .A2(n7515), .ZN(n7521) );
  NAND2_X1 U9130 ( .A1(n7521), .A2(n7517), .ZN(n7518) );
  NOR2_X1 U9131 ( .A1(n7519), .A2(n4284), .ZN(n7520) );
  INV_X2 U9132 ( .A(n8718), .ZN(n9925) );
  AOI22_X1 U9133 ( .A1(n7523), .A2(n9933), .B1(n7522), .B2(n9925), .ZN(n7525)
         );
  NAND2_X1 U9134 ( .A1(n9937), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n7524) );
  OAI211_X1 U9135 ( .C1(n7526), .C2(n8932), .A(n7525), .B(n7524), .ZN(n7533)
         );
  NAND2_X1 U9136 ( .A1(n7528), .A2(n8118), .ZN(n7707) );
  AND2_X1 U9137 ( .A1(n8883), .A2(n7707), .ZN(n7529) );
  OAI22_X1 U9138 ( .A1(n7531), .A2(n9906), .B1(n8918), .B2(n7530), .ZN(n7532)
         );
  OR2_X1 U9139 ( .A1(n7533), .A2(n7532), .ZN(P2_U3292) );
  NAND2_X1 U9140 ( .A1(n7534), .A2(n7600), .ZN(n7602) );
  NAND2_X1 U9141 ( .A1(n7602), .A2(n7535), .ZN(n7759) );
  NAND3_X1 U9142 ( .A1(n8514), .A2(n7536), .A3(n8615), .ZN(n7537) );
  OAI21_X1 U9143 ( .B1(n7602), .B2(n8593), .A(n7537), .ZN(n7539) );
  NAND2_X1 U9144 ( .A1(n7539), .A2(n7538), .ZN(n7545) );
  INV_X1 U9145 ( .A(n8597), .ZN(n8565) );
  INV_X1 U9146 ( .A(n7718), .ZN(n7540) );
  OAI22_X1 U9147 ( .A1(n8598), .A2(n7726), .B1(n7540), .B2(n8585), .ZN(n7543)
         );
  INV_X1 U9148 ( .A(n7721), .ZN(n9994) );
  OAI21_X1 U9149 ( .B1(n8604), .B2(n9994), .A(n7541), .ZN(n7542) );
  AOI211_X1 U9150 ( .C1(n8565), .C2(n8613), .A(n7543), .B(n7542), .ZN(n7544)
         );
  OAI211_X1 U9151 ( .C1(n8593), .C2(n7759), .A(n7545), .B(n7544), .ZN(P2_U3233) );
  NAND2_X1 U9152 ( .A1(n9555), .A2(n9557), .ZN(n9554) );
  NAND2_X1 U9153 ( .A1(n9571), .A2(n9154), .ZN(n7549) );
  NAND2_X1 U9154 ( .A1(n9554), .A2(n7549), .ZN(n7822) );
  XNOR2_X1 U9155 ( .A(n7822), .B(n7556), .ZN(n9595) );
  INV_X1 U9156 ( .A(n7553), .ZN(n7555) );
  OAI21_X1 U9157 ( .B1(n9558), .B2(n7555), .A(n7554), .ZN(n7557) );
  NOR2_X1 U9158 ( .A1(n7557), .A2(n7556), .ZN(n7558) );
  OAI21_X1 U9159 ( .B1(n7558), .B2(n7827), .A(n9786), .ZN(n7560) );
  AOI22_X1 U9160 ( .A1(n9736), .A2(n9152), .B1(n9734), .B2(n9154), .ZN(n7559)
         );
  NAND2_X1 U9161 ( .A1(n7560), .A2(n7559), .ZN(n7561) );
  AOI21_X1 U9162 ( .B1(n9595), .B2(n9565), .A(n7561), .ZN(n9597) );
  OR2_X1 U9163 ( .A1(n9570), .A2(n9571), .ZN(n9572) );
  AND2_X1 U9164 ( .A1(n9572), .A2(n7823), .ZN(n7562) );
  NOR2_X2 U9165 ( .A1(n9572), .A2(n7823), .ZN(n7829) );
  OR2_X1 U9166 ( .A1(n7562), .A2(n7829), .ZN(n9593) );
  OAI22_X1 U9167 ( .A1(n9797), .A2(n7441), .B1(n7677), .B2(n9792), .ZN(n7563)
         );
  AOI21_X1 U9168 ( .B1(n7823), .B2(n9569), .A(n7563), .ZN(n7564) );
  OAI21_X1 U9169 ( .B1(n9593), .B2(n9251), .A(n7564), .ZN(n7565) );
  AOI21_X1 U9170 ( .B1(n9595), .B2(n9778), .A(n7565), .ZN(n7566) );
  OAI21_X1 U9171 ( .B1(n9597), .B2(n9383), .A(n7566), .ZN(P1_U3278) );
  NAND2_X1 U9172 ( .A1(n7727), .A2(n8398), .ZN(n8154) );
  INV_X1 U9173 ( .A(n7727), .ZN(n8617) );
  INV_X1 U9174 ( .A(n8398), .ZN(n9972) );
  NAND2_X1 U9175 ( .A1(n8617), .A2(n9972), .ZN(n8149) );
  NAND2_X1 U9176 ( .A1(n7079), .A2(n7567), .ZN(n7568) );
  XOR2_X1 U9177 ( .A(n8092), .B(n7686), .Z(n9976) );
  INV_X1 U9178 ( .A(n9976), .ZN(n7581) );
  OAI21_X1 U9179 ( .B1(n8092), .B2(n7571), .A(n7681), .ZN(n7572) );
  INV_X1 U9180 ( .A(n8396), .ZN(n8616) );
  AOI222_X1 U9181 ( .A1(n9922), .A2(n7572), .B1(n8616), .B2(n8862), .C1(n8618), 
        .C2(n8861), .ZN(n7573) );
  INV_X1 U9182 ( .A(n7573), .ZN(n9974) );
  AOI22_X1 U9183 ( .A1(n8932), .A2(P2_REG2_REG_6__SCAN_IN), .B1(n8394), .B2(
        n9925), .ZN(n7578) );
  NOR2_X1 U9184 ( .A1(n7574), .A2(n9972), .ZN(n7575) );
  OR2_X1 U9185 ( .A1(n7733), .A2(n7575), .ZN(n9973) );
  INV_X1 U9186 ( .A(n9973), .ZN(n7576) );
  NAND2_X1 U9187 ( .A1(n8896), .A2(n7576), .ZN(n7577) );
  OAI211_X1 U9188 ( .C1(n9906), .C2(n9972), .A(n7578), .B(n7577), .ZN(n7579)
         );
  AOI21_X1 U9189 ( .B1(n9974), .B2(n8916), .A(n7579), .ZN(n7580) );
  OAI21_X1 U9190 ( .B1(n7581), .B2(n8918), .A(n7580), .ZN(P2_U3290) );
  MUX2_X1 U9191 ( .A(n7582), .B(P2_REG2_REG_1__SCAN_IN), .S(n9937), .Z(n7587)
         );
  AOI22_X1 U9192 ( .A1(n9933), .A2(n7583), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n9925), .ZN(n7584) );
  OAI21_X1 U9193 ( .B1(n9906), .B2(n7585), .A(n7584), .ZN(n7586) );
  AOI211_X1 U9194 ( .C1(n9934), .C2(n7588), .A(n7587), .B(n7586), .ZN(n7589)
         );
  INV_X1 U9195 ( .A(n7589), .ZN(P2_U3295) );
  NOR2_X1 U9196 ( .A1(n8425), .A2(n9952), .ZN(n8145) );
  INV_X1 U9197 ( .A(n7590), .ZN(n7591) );
  OR2_X1 U9198 ( .A1(n8145), .A2(n7591), .ZN(n9954) );
  NOR2_X1 U9199 ( .A1(n8413), .A2(n8907), .ZN(n7592) );
  AOI21_X1 U9200 ( .B1(n9954), .B2(n9922), .A(n7592), .ZN(n9956) );
  INV_X1 U9201 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n7593) );
  OAI22_X1 U9202 ( .A1(n9937), .A2(n9956), .B1(n7593), .B2(n8718), .ZN(n7596)
         );
  INV_X1 U9203 ( .A(n9954), .ZN(n7594) );
  NOR2_X1 U9204 ( .A1(n8918), .A2(n7594), .ZN(n7595) );
  AOI211_X1 U9205 ( .C1(n9937), .C2(P2_REG2_REG_0__SCAN_IN), .A(n7596), .B(
        n7595), .ZN(n7598) );
  OAI21_X1 U9206 ( .B1(n9931), .B2(n8896), .A(n9952), .ZN(n7597) );
  NAND2_X1 U9207 ( .A1(n7598), .A2(n7597), .ZN(P2_U3296) );
  NAND3_X1 U9208 ( .A1(n8514), .A2(n7599), .A3(n8616), .ZN(n7605) );
  OAI21_X1 U9209 ( .B1(n7601), .B2(n7600), .A(n8488), .ZN(n7604) );
  INV_X1 U9210 ( .A(n7602), .ZN(n7603) );
  AOI21_X1 U9211 ( .B1(n7605), .B2(n7604), .A(n7603), .ZN(n7611) );
  INV_X1 U9212 ( .A(n7692), .ZN(n7606) );
  OAI22_X1 U9213 ( .A1(n8597), .A2(n7889), .B1(n8585), .B2(n7606), .ZN(n7610)
         );
  AOI21_X1 U9214 ( .B1(n8589), .B2(n7702), .A(n7607), .ZN(n7608) );
  OAI21_X1 U9215 ( .B1(n8598), .B2(n8396), .A(n7608), .ZN(n7609) );
  OR3_X1 U9216 ( .A1(n7611), .A2(n7610), .A3(n7609), .ZN(P2_U3223) );
  OAI21_X1 U9217 ( .B1(n7614), .B2(n7612), .A(n7613), .ZN(n9962) );
  AND2_X1 U9218 ( .A1(n7615), .A2(n8373), .ZN(n7616) );
  NOR2_X1 U9219 ( .A1(n9927), .A2(n7616), .ZN(n9958) );
  AOI22_X1 U9220 ( .A1(n8896), .A2(n9958), .B1(P2_REG3_REG_2__SCAN_IN), .B2(
        n9925), .ZN(n7617) );
  OAI21_X1 U9221 ( .B1(n7070), .B2(n9906), .A(n7617), .ZN(n7623) );
  INV_X1 U9222 ( .A(n7618), .ZN(n7619) );
  AOI21_X1 U9223 ( .B1(n7612), .B2(n7620), .A(n7619), .ZN(n7621) );
  OAI222_X1 U9224 ( .A1(n8907), .A2(n7074), .B1(n8905), .B2(n8413), .C1(n8920), 
        .C2(n7621), .ZN(n9960) );
  MUX2_X1 U9225 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n9960), .S(n8916), .Z(n7622)
         );
  AOI211_X1 U9226 ( .C1(n9934), .C2(n9962), .A(n7623), .B(n7622), .ZN(n7624)
         );
  INV_X1 U9227 ( .A(n7624), .ZN(P2_U3294) );
  AOI211_X1 U9228 ( .C1(n7626), .C2(n7625), .A(n4371), .B(n9895), .ZN(n7635)
         );
  XNOR2_X1 U9229 ( .A(n7628), .B(n7627), .ZN(n7633) );
  NAND2_X1 U9230 ( .A1(n9522), .A2(n7629), .ZN(n7632) );
  NOR2_X1 U9231 ( .A1(n7630), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7775) );
  AOI21_X1 U9232 ( .B1(n9892), .B2(P2_ADDR_REG_13__SCAN_IN), .A(n7775), .ZN(
        n7631) );
  OAI211_X1 U9233 ( .C1(n7633), .C2(n9894), .A(n7632), .B(n7631), .ZN(n7634)
         );
  OR2_X1 U9234 ( .A1(n7635), .A2(n7634), .ZN(P2_U3258) );
  NAND2_X1 U9235 ( .A1(n9140), .A2(n7636), .ZN(n7639) );
  NAND2_X1 U9236 ( .A1(P1_U3084), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n8336) );
  INV_X1 U9237 ( .A(n8336), .ZN(n7637) );
  AOI21_X1 U9238 ( .B1(n9139), .B2(n9155), .A(n7637), .ZN(n7638) );
  OAI211_X1 U9239 ( .C1(n7674), .C2(n9123), .A(n7639), .B(n7638), .ZN(n7645)
         );
  INV_X1 U9240 ( .A(n7640), .ZN(n7641) );
  AOI211_X1 U9241 ( .C1(n7643), .C2(n7642), .A(n9131), .B(n7641), .ZN(n7644)
         );
  AOI211_X1 U9242 ( .C1(n9470), .C2(n9129), .A(n7645), .B(n7644), .ZN(n7646)
         );
  INV_X1 U9243 ( .A(n7646), .ZN(P1_U3234) );
  INV_X1 U9244 ( .A(n7647), .ZN(n8057) );
  OAI222_X1 U9245 ( .A1(n9502), .A2(n7649), .B1(n4282), .B2(n8057), .C1(
        P1_U3084), .C2(n7648), .ZN(P1_U3331) );
  INV_X1 U9246 ( .A(n7650), .ZN(n7651) );
  AOI21_X1 U9247 ( .B1(n7653), .B2(n7652), .A(n7651), .ZN(n7660) );
  OAI21_X1 U9248 ( .B1(n9114), .B2(n7655), .A(n7654), .ZN(n7657) );
  NOR2_X1 U9249 ( .A1(n9127), .A2(n9566), .ZN(n7656) );
  AOI211_X1 U9250 ( .C1(n9145), .C2(n9153), .A(n7657), .B(n7656), .ZN(n7659)
         );
  NAND2_X1 U9251 ( .A1(n9571), .A2(n9129), .ZN(n7658) );
  OAI211_X1 U9252 ( .C1(n7660), .C2(n9131), .A(n7659), .B(n7658), .ZN(P1_U3222) );
  AOI22_X1 U9253 ( .A1(n7662), .A2(n9934), .B1(n9931), .B2(n7661), .ZN(n7667)
         );
  AOI22_X1 U9254 ( .A1(n8932), .A2(P2_REG2_REG_5__SCAN_IN), .B1(n7663), .B2(
        n9925), .ZN(n7666) );
  NOR2_X1 U9255 ( .A1(n8932), .A2(n4284), .ZN(n8868) );
  NAND2_X1 U9256 ( .A1(n8868), .A2(n7664), .ZN(n7665) );
  AND3_X1 U9257 ( .A1(n7667), .A2(n7666), .A3(n7665), .ZN(n7668) );
  OAI21_X1 U9258 ( .B1(n9937), .B2(n7669), .A(n7668), .ZN(P2_U3291) );
  XNOR2_X1 U9259 ( .A(n7671), .B(n7670), .ZN(n7672) );
  XNOR2_X1 U9260 ( .A(n7673), .B(n7672), .ZN(n7680) );
  AND2_X1 U9261 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9644) );
  NOR2_X1 U9262 ( .A1(n9114), .A2(n7674), .ZN(n7675) );
  AOI211_X1 U9263 ( .C1(n9145), .C2(n9152), .A(n9644), .B(n7675), .ZN(n7676)
         );
  OAI21_X1 U9264 ( .B1(n9127), .B2(n7677), .A(n7676), .ZN(n7678) );
  AOI21_X1 U9265 ( .B1(n7823), .B2(n9129), .A(n7678), .ZN(n7679) );
  OAI21_X1 U9266 ( .B1(n7680), .B2(n9131), .A(n7679), .ZN(P1_U3232) );
  NAND2_X1 U9267 ( .A1(n7726), .A2(n7702), .ZN(n8156) );
  INV_X1 U9268 ( .A(n7702), .ZN(n9986) );
  NAND2_X1 U9269 ( .A1(n8615), .A2(n9986), .ZN(n8163) );
  NAND2_X1 U9270 ( .A1(n8156), .A2(n8163), .ZN(n7689) );
  NAND2_X1 U9271 ( .A1(n8396), .A2(n7734), .ZN(n8161) );
  NAND2_X1 U9272 ( .A1(n8616), .A2(n9979), .ZN(n8155) );
  INV_X1 U9273 ( .A(n7684), .ZN(n7683) );
  NAND2_X1 U9274 ( .A1(n7683), .A2(n7682), .ZN(n7710) );
  INV_X1 U9275 ( .A(n7710), .ZN(n7709) );
  AOI21_X1 U9276 ( .B1(n7689), .B2(n7684), .A(n7709), .ZN(n7685) );
  OAI222_X1 U9277 ( .A1(n8907), .A2(n7889), .B1(n8905), .B2(n8396), .C1(n8920), 
        .C2(n7685), .ZN(n9988) );
  NAND2_X1 U9278 ( .A1(n7732), .A2(n7731), .ZN(n7688) );
  NAND2_X1 U9279 ( .A1(n8396), .A2(n9979), .ZN(n7687) );
  INV_X1 U9280 ( .A(n9990), .ZN(n7691) );
  AND2_X1 U9281 ( .A1(n7690), .A2(n7682), .ZN(n9985) );
  NOR3_X1 U9282 ( .A1(n7691), .A2(n9985), .A3(n8918), .ZN(n7700) );
  AOI22_X1 U9283 ( .A1(n8932), .A2(P2_REG2_REG_8__SCAN_IN), .B1(n7692), .B2(
        n9925), .ZN(n7698) );
  NAND2_X1 U9284 ( .A1(n7733), .A2(n9979), .ZN(n7693) );
  NAND2_X1 U9285 ( .A1(n7693), .A2(n7702), .ZN(n7695) );
  NOR2_X1 U9286 ( .A1(n7702), .A2(n7734), .ZN(n7694) );
  NAND2_X1 U9287 ( .A1(n7695), .A2(n7716), .ZN(n9987) );
  INV_X1 U9288 ( .A(n9987), .ZN(n7696) );
  NAND2_X1 U9289 ( .A1(n8896), .A2(n7696), .ZN(n7697) );
  OAI211_X1 U9290 ( .C1(n9906), .C2(n9986), .A(n7698), .B(n7697), .ZN(n7699)
         );
  AOI211_X1 U9291 ( .C1(n9988), .C2(n8916), .A(n7700), .B(n7699), .ZN(n7701)
         );
  INV_X1 U9292 ( .A(n7701), .ZN(P2_U3288) );
  NAND2_X1 U9293 ( .A1(n7889), .A2(n7721), .ZN(n8173) );
  INV_X1 U9294 ( .A(n7889), .ZN(n8614) );
  NAND2_X1 U9295 ( .A1(n8614), .A2(n9994), .ZN(n8164) );
  NAND2_X1 U9296 ( .A1(n8615), .A2(n7702), .ZN(n7703) );
  INV_X1 U9297 ( .A(n7706), .ZN(n7704) );
  INV_X1 U9298 ( .A(n7784), .ZN(n7705) );
  AOI21_X1 U9299 ( .B1(n8100), .B2(n7706), .A(n7705), .ZN(n9993) );
  AOI22_X1 U9300 ( .A1(n8861), .A2(n8615), .B1(n8613), .B2(n8862), .ZN(n7715)
         );
  INV_X1 U9301 ( .A(n8156), .ZN(n7708) );
  NOR3_X1 U9302 ( .A1(n7709), .A2(n8100), .A3(n7708), .ZN(n7713) );
  NAND2_X1 U9303 ( .A1(n7710), .A2(n8156), .ZN(n7711) );
  INV_X1 U9304 ( .A(n7778), .ZN(n7712) );
  OAI21_X1 U9305 ( .B1(n7713), .B2(n7712), .A(n9922), .ZN(n7714) );
  OAI211_X1 U9306 ( .C1(n9993), .C2(n8883), .A(n7715), .B(n7714), .ZN(n9996)
         );
  NAND2_X1 U9307 ( .A1(n9996), .A2(n8916), .ZN(n7723) );
  INV_X1 U9308 ( .A(n8896), .ZN(n8914) );
  INV_X1 U9309 ( .A(n7716), .ZN(n7717) );
  OAI21_X1 U9310 ( .B1(n7717), .B2(n9994), .A(n7858), .ZN(n9995) );
  AOI22_X1 U9311 ( .A1(n9937), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n7718), .B2(
        n9925), .ZN(n7719) );
  OAI21_X1 U9312 ( .B1(n8914), .B2(n9995), .A(n7719), .ZN(n7720) );
  AOI21_X1 U9313 ( .B1(n9931), .B2(n7721), .A(n7720), .ZN(n7722) );
  OAI211_X1 U9314 ( .C1(n9993), .C2(n8893), .A(n7723), .B(n7722), .ZN(P2_U3287) );
  XNOR2_X1 U9315 ( .A(n7724), .B(n4588), .ZN(n7725) );
  NAND2_X1 U9316 ( .A1(n7725), .A2(n9922), .ZN(n7730) );
  OAI22_X1 U9317 ( .A1(n7727), .A2(n8905), .B1(n7726), .B2(n8907), .ZN(n7728)
         );
  INV_X1 U9318 ( .A(n7728), .ZN(n7729) );
  NAND2_X1 U9319 ( .A1(n7730), .A2(n7729), .ZN(n9983) );
  INV_X1 U9320 ( .A(n9983), .ZN(n7740) );
  XNOR2_X1 U9321 ( .A(n7732), .B(n7731), .ZN(n9978) );
  XNOR2_X1 U9322 ( .A(n7733), .B(n9979), .ZN(n9980) );
  NAND2_X1 U9323 ( .A1(n9931), .A2(n7734), .ZN(n7737) );
  AOI22_X1 U9324 ( .A1(n8932), .A2(P2_REG2_REG_7__SCAN_IN), .B1(n7735), .B2(
        n9925), .ZN(n7736) );
  OAI211_X1 U9325 ( .C1(n8914), .C2(n9980), .A(n7737), .B(n7736), .ZN(n7738)
         );
  AOI21_X1 U9326 ( .B1(n9978), .B2(n9934), .A(n7738), .ZN(n7739) );
  OAI21_X1 U9327 ( .B1(n7740), .B2(n9937), .A(n7739), .ZN(P2_U3289) );
  AOI21_X1 U9328 ( .B1(n7743), .B2(n7742), .A(n7741), .ZN(n7754) );
  OAI21_X1 U9329 ( .B1(n7746), .B2(n7745), .A(n7744), .ZN(n7747) );
  NAND2_X1 U9330 ( .A1(n7747), .A2(n9889), .ZN(n7753) );
  INV_X1 U9331 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7748) );
  NAND2_X1 U9332 ( .A1(P2_U3152), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n7931) );
  OAI21_X1 U9333 ( .B1(n7749), .B2(n7748), .A(n7931), .ZN(n7750) );
  AOI21_X1 U9334 ( .B1(n9522), .B2(n7751), .A(n7750), .ZN(n7752) );
  OAI211_X1 U9335 ( .C1(n7754), .C2(n9894), .A(n7753), .B(n7752), .ZN(P2_U3259) );
  NAND2_X1 U9336 ( .A1(n7769), .A2(n8053), .ZN(n7756) );
  OAI211_X1 U9337 ( .C1(n7757), .C2(n9502), .A(n7756), .B(n7755), .ZN(P1_U3330) );
  NAND2_X1 U9338 ( .A1(n7759), .A2(n7758), .ZN(n7882) );
  OR2_X1 U9339 ( .A1(n7882), .A2(n7883), .ZN(n7880) );
  AOI21_X1 U9340 ( .B1(n7880), .B2(n4375), .A(n8593), .ZN(n7763) );
  NOR3_X1 U9341 ( .A1(n8592), .A2(n7779), .A3(n7760), .ZN(n7762) );
  OAI21_X1 U9342 ( .B1(n7763), .B2(n7762), .A(n7761), .ZN(n7768) );
  INV_X1 U9343 ( .A(n8598), .ZN(n8566) );
  INV_X1 U9344 ( .A(n8611), .ZN(n7998) );
  INV_X1 U9345 ( .A(n7764), .ZN(n7857) );
  OAI22_X1 U9346 ( .A1(n8597), .A2(n7998), .B1(n8585), .B2(n7857), .ZN(n7766)
         );
  OAI22_X1 U9347 ( .A1(n8604), .A2(n10013), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5917), .ZN(n7765) );
  AOI211_X1 U9348 ( .C1(n8566), .C2(n8613), .A(n7766), .B(n7765), .ZN(n7767)
         );
  NAND2_X1 U9349 ( .A1(n7768), .A2(n7767), .ZN(P2_U3238) );
  NAND2_X1 U9350 ( .A1(n7769), .A2(n9044), .ZN(n7770) );
  OAI211_X1 U9351 ( .C1(n7771), .C2(n9041), .A(n7770), .B(n8270), .ZN(P2_U3335) );
  OAI211_X1 U9352 ( .C1(n7773), .C2(n7772), .A(n7925), .B(n8488), .ZN(n7777)
         );
  OAI22_X1 U9353 ( .A1(n7998), .A2(n8598), .B1(n8597), .B2(n8904), .ZN(n7774)
         );
  AOI211_X1 U9354 ( .C1(n8601), .C2(n8006), .A(n7775), .B(n7774), .ZN(n7776)
         );
  OAI211_X1 U9355 ( .C1(n8003), .C2(n8604), .A(n7777), .B(n7776), .ZN(P2_U3236) );
  NAND2_X1 U9356 ( .A1(n7779), .A2(n7887), .ZN(n8157) );
  INV_X1 U9357 ( .A(n7887), .ZN(n10003) );
  NAND2_X1 U9358 ( .A1(n8613), .A2(n10003), .ZN(n8166) );
  NAND2_X1 U9359 ( .A1(n8157), .A2(n8166), .ZN(n7852) );
  XNOR2_X1 U9360 ( .A(n7853), .B(n7852), .ZN(n7780) );
  OAI222_X1 U9361 ( .A1(n8907), .A2(n7904), .B1(n8905), .B2(n7889), .C1(n7780), 
        .C2(n8920), .ZN(n10006) );
  XNOR2_X1 U9362 ( .A(n7858), .B(n7887), .ZN(n10005) );
  NAND2_X1 U9363 ( .A1(n9931), .A2(n7887), .ZN(n7782) );
  AOI22_X1 U9364 ( .A1(n8932), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n7884), .B2(
        n9925), .ZN(n7781) );
  OAI211_X1 U9365 ( .C1(n10005), .C2(n8914), .A(n7782), .B(n7781), .ZN(n7788)
         );
  NAND2_X1 U9366 ( .A1(n7889), .A2(n9994), .ZN(n7783) );
  INV_X1 U9367 ( .A(n7852), .ZN(n8103) );
  INV_X1 U9368 ( .A(n10008), .ZN(n7786) );
  AND2_X1 U9369 ( .A1(n7785), .A2(n8103), .ZN(n10002) );
  NOR3_X1 U9370 ( .A1(n7786), .A2(n10002), .A3(n8918), .ZN(n7787) );
  AOI211_X1 U9371 ( .C1(n8916), .C2(n10006), .A(n7788), .B(n7787), .ZN(n7789)
         );
  INV_X1 U9372 ( .A(n7789), .ZN(P2_U3286) );
  INV_X1 U9373 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10080) );
  NOR2_X1 U9374 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7790) );
  AOI21_X1 U9375 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n7790), .ZN(n10052) );
  NOR2_X1 U9376 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7791) );
  AOI21_X1 U9377 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n7791), .ZN(n10055) );
  NOR2_X1 U9378 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7792) );
  AOI21_X1 U9379 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n7792), .ZN(n10058) );
  NOR2_X1 U9380 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7793) );
  AOI21_X1 U9381 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n7793), .ZN(n10061) );
  NOR2_X1 U9382 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7794) );
  AOI21_X1 U9383 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n7794), .ZN(n10064) );
  NOR2_X1 U9384 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7801) );
  XNOR2_X1 U9385 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10093) );
  NAND2_X1 U9386 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7799) );
  XOR2_X1 U9387 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10091) );
  NAND2_X1 U9388 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n7797) );
  XOR2_X1 U9389 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(P1_ADDR_REG_2__SCAN_IN), .Z(
        n10088) );
  AOI21_X1 U9390 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10046) );
  INV_X1 U9391 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n7795) );
  NAND3_X1 U9392 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n10048) );
  OAI21_X1 U9393 ( .B1(n10046), .B2(n7795), .A(n10048), .ZN(n10087) );
  NAND2_X1 U9394 ( .A1(n10088), .A2(n10087), .ZN(n7796) );
  NAND2_X1 U9395 ( .A1(n7797), .A2(n7796), .ZN(n10090) );
  NAND2_X1 U9396 ( .A1(n10091), .A2(n10090), .ZN(n7798) );
  NAND2_X1 U9397 ( .A1(n7799), .A2(n7798), .ZN(n10092) );
  NOR2_X1 U9398 ( .A1(n10093), .A2(n10092), .ZN(n7800) );
  NOR2_X1 U9399 ( .A1(n7801), .A2(n7800), .ZN(n7802) );
  NOR2_X1 U9400 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n7802), .ZN(n10076) );
  AND2_X1 U9401 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n7802), .ZN(n10075) );
  NOR2_X1 U9402 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10075), .ZN(n7803) );
  NOR2_X1 U9403 ( .A1(n10076), .A2(n7803), .ZN(n7804) );
  NAND2_X1 U9404 ( .A1(n7804), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n7806) );
  XOR2_X1 U9405 ( .A(n7804), .B(P1_ADDR_REG_6__SCAN_IN), .Z(n10074) );
  NAND2_X1 U9406 ( .A1(n10074), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n7805) );
  NAND2_X1 U9407 ( .A1(n7806), .A2(n7805), .ZN(n7807) );
  NAND2_X1 U9408 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n7807), .ZN(n7809) );
  XOR2_X1 U9409 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n7807), .Z(n10083) );
  NAND2_X1 U9410 ( .A1(n10083), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n7808) );
  NAND2_X1 U9411 ( .A1(n7809), .A2(n7808), .ZN(n7810) );
  NAND2_X1 U9412 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n7810), .ZN(n7812) );
  XOR2_X1 U9413 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n7810), .Z(n10089) );
  NAND2_X1 U9414 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10089), .ZN(n7811) );
  NAND2_X1 U9415 ( .A1(n7812), .A2(n7811), .ZN(n7813) );
  AND2_X1 U9416 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n7813), .ZN(n7814) );
  XNOR2_X1 U9417 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n7813), .ZN(n10085) );
  NOR2_X1 U9418 ( .A1(n10086), .A2(n10085), .ZN(n10084) );
  NAND2_X1 U9419 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n7815) );
  OAI21_X1 U9420 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n7815), .ZN(n10072) );
  NAND2_X1 U9421 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n7816) );
  OAI21_X1 U9422 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n7816), .ZN(n10069) );
  NOR2_X1 U9423 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7817) );
  AOI21_X1 U9424 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n7817), .ZN(n10066) );
  NAND2_X1 U9425 ( .A1(n10067), .A2(n10066), .ZN(n10065) );
  NAND2_X1 U9426 ( .A1(n10064), .A2(n10063), .ZN(n10062) );
  NAND2_X1 U9427 ( .A1(n10061), .A2(n10060), .ZN(n10059) );
  OAI21_X1 U9428 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10059), .ZN(n10057) );
  NAND2_X1 U9429 ( .A1(n10058), .A2(n10057), .ZN(n10056) );
  OAI21_X1 U9430 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10056), .ZN(n10054) );
  NAND2_X1 U9431 ( .A1(n10055), .A2(n10054), .ZN(n10053) );
  OAI21_X1 U9432 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10053), .ZN(n10051) );
  NAND2_X1 U9433 ( .A1(n10052), .A2(n10051), .ZN(n10050) );
  OAI21_X1 U9434 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10050), .ZN(n10079) );
  NOR2_X1 U9435 ( .A1(n10080), .A2(n10079), .ZN(n7818) );
  NAND2_X1 U9436 ( .A1(n10080), .A2(n10079), .ZN(n10078) );
  OAI21_X1 U9437 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n7818), .A(n10078), .ZN(
        n7820) );
  XNOR2_X1 U9438 ( .A(n8307), .B(P2_ADDR_REG_19__SCAN_IN), .ZN(n7819) );
  XNOR2_X1 U9439 ( .A(n7820), .B(n7819), .ZN(ADD_1071_U4) );
  NAND2_X1 U9440 ( .A1(n7822), .A2(n7821), .ZN(n7824) );
  INV_X1 U9441 ( .A(n7823), .ZN(n9592) );
  NAND2_X1 U9442 ( .A1(n7824), .A2(n4841), .ZN(n7841) );
  XNOR2_X1 U9443 ( .A(n7841), .B(n7837), .ZN(n9590) );
  INV_X1 U9444 ( .A(n9590), .ZN(n7835) );
  INV_X1 U9445 ( .A(n7825), .ZN(n7826) );
  XOR2_X1 U9446 ( .A(n7837), .B(n7838), .Z(n7828) );
  AOI222_X1 U9447 ( .A1(n9786), .A2(n7828), .B1(n9151), .B2(n9736), .C1(n9153), 
        .C2(n9734), .ZN(n9587) );
  OAI21_X1 U9448 ( .B1(n7875), .B2(n9792), .A(n9587), .ZN(n7833) );
  OAI211_X1 U9449 ( .C1(n7829), .C2(n9588), .A(n7844), .B(n9857), .ZN(n9586)
         );
  AOI22_X1 U9450 ( .A1(n7877), .A2(n9569), .B1(P1_REG2_REG_14__SCAN_IN), .B2(
        n9383), .ZN(n7830) );
  OAI21_X1 U9451 ( .B1(n9586), .B2(n7831), .A(n7830), .ZN(n7832) );
  AOI21_X1 U9452 ( .B1(n7833), .B2(n9797), .A(n7832), .ZN(n7834) );
  OAI21_X1 U9453 ( .B1(n7835), .B2(n9387), .A(n7834), .ZN(P1_U3277) );
  OAI21_X1 U9454 ( .B1(n7839), .B2(n7842), .A(n7979), .ZN(n7840) );
  AOI222_X1 U9455 ( .A1(n9786), .A2(n7840), .B1(n9150), .B2(n9736), .C1(n9152), 
        .C2(n9734), .ZN(n9579) );
  XNOR2_X1 U9456 ( .A(n7915), .B(n7842), .ZN(n9584) );
  NAND2_X1 U9457 ( .A1(n9584), .A2(n8042), .ZN(n7849) );
  INV_X1 U9458 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n7843) );
  OAI22_X1 U9459 ( .A1(n9797), .A2(n7843), .B1(n7964), .B2(n9792), .ZN(n7847)
         );
  INV_X1 U9460 ( .A(n7844), .ZN(n7845) );
  OAI21_X1 U9461 ( .B1(n7845), .B2(n9580), .A(n7916), .ZN(n9581) );
  NOR2_X1 U9462 ( .A1(n9581), .A2(n9251), .ZN(n7846) );
  AOI211_X1 U9463 ( .C1(n9569), .C2(n7912), .A(n7847), .B(n7846), .ZN(n7848)
         );
  OAI211_X1 U9464 ( .C1(n9383), .C2(n9579), .A(n7849), .B(n7848), .ZN(P1_U3276) );
  NAND2_X1 U9465 ( .A1(n8613), .A2(n7887), .ZN(n7850) );
  NAND2_X1 U9466 ( .A1(n10008), .A2(n7850), .ZN(n7851) );
  NAND2_X1 U9467 ( .A1(n7904), .A2(n7988), .ZN(n8177) );
  INV_X1 U9468 ( .A(n7904), .ZN(n8612) );
  NAND2_X1 U9469 ( .A1(n10013), .A2(n8612), .ZN(n8175) );
  NAND2_X1 U9470 ( .A1(n8177), .A2(n8175), .ZN(n8102) );
  OAI21_X1 U9471 ( .B1(n7851), .B2(n8102), .A(n7990), .ZN(n10011) );
  XNOR2_X1 U9472 ( .A(n7995), .B(n8102), .ZN(n7854) );
  NAND2_X1 U9473 ( .A1(n7854), .A2(n9922), .ZN(n7856) );
  AOI22_X1 U9474 ( .A1(n8613), .A2(n8861), .B1(n8862), .B2(n8611), .ZN(n7855)
         );
  NAND2_X1 U9475 ( .A1(n7856), .A2(n7855), .ZN(n10014) );
  NAND2_X1 U9476 ( .A1(n10014), .A2(n8916), .ZN(n7864) );
  OAI22_X1 U9477 ( .A1(n8916), .A2(n6226), .B1(n7857), .B2(n8718), .ZN(n7862)
         );
  OAI211_X1 U9478 ( .C1(n7859), .C2(n10013), .A(n9911), .B(n9913), .ZN(n10012)
         );
  INV_X1 U9479 ( .A(n9933), .ZN(n7860) );
  NOR2_X1 U9480 ( .A1(n10012), .A2(n7860), .ZN(n7861) );
  AOI211_X1 U9481 ( .C1(n9931), .C2(n7988), .A(n7862), .B(n7861), .ZN(n7863)
         );
  OAI211_X1 U9482 ( .C1(n8918), .C2(n10011), .A(n7864), .B(n7863), .ZN(
        P2_U3285) );
  NAND2_X1 U9483 ( .A1(n7893), .A2(n9044), .ZN(n7866) );
  OAI211_X1 U9484 ( .C1(n9047), .C2(n7867), .A(n7866), .B(n7865), .ZN(P2_U3334) );
  XNOR2_X1 U9485 ( .A(n7869), .B(n7868), .ZN(n7870) );
  XNOR2_X1 U9486 ( .A(n7871), .B(n7870), .ZN(n7879) );
  NOR2_X1 U9487 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7872), .ZN(n9657) );
  NOR2_X1 U9488 ( .A1(n9114), .A2(n9561), .ZN(n7873) );
  AOI211_X1 U9489 ( .C1(n9145), .C2(n9151), .A(n9657), .B(n7873), .ZN(n7874)
         );
  OAI21_X1 U9490 ( .B1(n9127), .B2(n7875), .A(n7874), .ZN(n7876) );
  AOI21_X1 U9491 ( .B1(n7877), .B2(n9129), .A(n7876), .ZN(n7878) );
  OAI21_X1 U9492 ( .B1(n7879), .B2(n9131), .A(n7878), .ZN(P1_U3213) );
  INV_X1 U9493 ( .A(n7880), .ZN(n7881) );
  AOI211_X1 U9494 ( .C1(n7883), .C2(n7882), .A(n8593), .B(n7881), .ZN(n7892)
         );
  INV_X1 U9495 ( .A(n7884), .ZN(n7885) );
  OAI22_X1 U9496 ( .A1(n8597), .A2(n7904), .B1(n8585), .B2(n7885), .ZN(n7891)
         );
  AOI21_X1 U9497 ( .B1(n8589), .B2(n7887), .A(n7886), .ZN(n7888) );
  OAI21_X1 U9498 ( .B1(n8598), .B2(n7889), .A(n7888), .ZN(n7890) );
  OR3_X1 U9499 ( .A1(n7892), .A2(n7891), .A3(n7890), .ZN(P2_U3219) );
  INV_X1 U9500 ( .A(n7893), .ZN(n7895) );
  OAI222_X1 U9501 ( .A1(P1_U3084), .A2(n7896), .B1(n4282), .B2(n7895), .C1(
        n7894), .C2(n9502), .ZN(P1_U3329) );
  INV_X1 U9502 ( .A(n7772), .ZN(n7903) );
  INV_X1 U9503 ( .A(n7897), .ZN(n7899) );
  NAND2_X1 U9504 ( .A1(n7899), .A2(n7898), .ZN(n7901) );
  AOI22_X1 U9505 ( .A1(n7903), .A2(n7902), .B1(n7901), .B2(n7900), .ZN(n7911)
         );
  INV_X1 U9506 ( .A(n9904), .ZN(n7907) );
  INV_X1 U9507 ( .A(n8610), .ZN(n8067) );
  OAI22_X1 U9508 ( .A1(n8067), .A2(n8907), .B1(n7904), .B2(n8905), .ZN(n9902)
         );
  NAND2_X1 U9509 ( .A1(n8509), .A2(n9902), .ZN(n7906) );
  OAI211_X1 U9510 ( .C1(n8585), .C2(n7907), .A(n7906), .B(n7905), .ZN(n7909)
         );
  NOR3_X1 U9511 ( .A1(n7772), .A2(n7998), .A3(n8592), .ZN(n7908) );
  AOI211_X1 U9512 ( .C1(n8002), .C2(n8589), .A(n7909), .B(n7908), .ZN(n7910)
         );
  OAI21_X1 U9513 ( .B1(n7911), .B2(n8593), .A(n7910), .ZN(P2_U3226) );
  NAND2_X1 U9514 ( .A1(n9580), .A2(n7913), .ZN(n7914) );
  XNOR2_X1 U9515 ( .A(n7970), .B(n7969), .ZN(n9467) );
  AOI211_X1 U9516 ( .C1(n9465), .C2(n7916), .A(n9865), .B(n7975), .ZN(n9464)
         );
  NOR2_X1 U9517 ( .A1(n4571), .A2(n9791), .ZN(n7919) );
  OAI22_X1 U9518 ( .A1(n9797), .A2(n7917), .B1(n8024), .B2(n9792), .ZN(n7918)
         );
  AOI211_X1 U9519 ( .C1(n9464), .C2(n9575), .A(n7919), .B(n7918), .ZN(n7924)
         );
  NAND2_X1 U9520 ( .A1(n7979), .A2(n7920), .ZN(n7921) );
  XNOR2_X1 U9521 ( .A(n7921), .B(n7969), .ZN(n7922) );
  OAI222_X1 U9522 ( .A1(n9781), .A2(n8037), .B1(n9784), .B2(n7913), .C1(n7922), 
        .C2(n9766), .ZN(n9463) );
  NAND2_X1 U9523 ( .A1(n9463), .A2(n9797), .ZN(n7923) );
  OAI211_X1 U9524 ( .C1(n9467), .C2(n9387), .A(n7924), .B(n7923), .ZN(P1_U3275) );
  INV_X1 U9525 ( .A(n7925), .ZN(n7928) );
  NOR3_X1 U9526 ( .A1(n8592), .A2(n8067), .A3(n7926), .ZN(n7927) );
  AOI21_X1 U9527 ( .B1(n7928), .B2(n8488), .A(n7927), .ZN(n7938) );
  INV_X1 U9528 ( .A(n8931), .ZN(n7933) );
  OR2_X1 U9529 ( .A1(n8877), .A2(n8907), .ZN(n7930) );
  NAND2_X1 U9530 ( .A1(n8610), .A2(n8861), .ZN(n7929) );
  NAND2_X1 U9531 ( .A1(n7930), .A2(n7929), .ZN(n8921) );
  NAND2_X1 U9532 ( .A1(n8509), .A2(n8921), .ZN(n7932) );
  OAI211_X1 U9533 ( .C1(n8585), .C2(n7933), .A(n7932), .B(n7931), .ZN(n7936)
         );
  NOR2_X1 U9534 ( .A1(n7934), .A2(n8593), .ZN(n7935) );
  AOI211_X1 U9535 ( .C1(n8927), .C2(n8589), .A(n7936), .B(n7935), .ZN(n7937)
         );
  OAI21_X1 U9536 ( .B1(n7939), .B2(n7938), .A(n7937), .ZN(P2_U3217) );
  INV_X1 U9537 ( .A(n7940), .ZN(n7945) );
  OAI222_X1 U9538 ( .A1(n9502), .A2(n7942), .B1(n4282), .B2(n7945), .C1(
        P1_U3084), .C2(n7941), .ZN(P1_U3328) );
  INV_X1 U9539 ( .A(n7943), .ZN(n7944) );
  OAI222_X1 U9540 ( .A1(n9047), .A2(n7946), .B1(n9049), .B2(n7945), .C1(
        P2_U3152), .C2(n7944), .ZN(P2_U3333) );
  OAI21_X1 U9541 ( .B1(n7949), .B2(n7948), .A(n7947), .ZN(n7957) );
  OAI211_X1 U9542 ( .C1(n7951), .C2(P2_REG1_REG_15__SCAN_IN), .A(n9888), .B(
        n7950), .ZN(n7954) );
  NOR2_X1 U9543 ( .A1(n7952), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8600) );
  AOI21_X1 U9544 ( .B1(n9892), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n8600), .ZN(
        n7953) );
  OAI211_X1 U9545 ( .C1(n9893), .C2(n7955), .A(n7954), .B(n7953), .ZN(n7956)
         );
  AOI21_X1 U9546 ( .B1(n9889), .B2(n7957), .A(n7956), .ZN(n7958) );
  INV_X1 U9547 ( .A(n7958), .ZN(P2_U3260) );
  INV_X1 U9548 ( .A(n8020), .ZN(n7962) );
  OAI21_X1 U9549 ( .B1(n7960), .B2(n8019), .A(n7959), .ZN(n7961) );
  OAI211_X1 U9550 ( .C1(n7962), .C2(n8019), .A(n9136), .B(n7961), .ZN(n7968)
         );
  NAND2_X1 U9551 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9669) );
  OAI21_X1 U9552 ( .B1(n9114), .B2(n7963), .A(n9669), .ZN(n7966) );
  NOR2_X1 U9553 ( .A1(n9127), .A2(n7964), .ZN(n7965) );
  AOI211_X1 U9554 ( .C1(n9145), .C2(n9150), .A(n7966), .B(n7965), .ZN(n7967)
         );
  OAI211_X1 U9555 ( .C1(n9580), .C2(n9148), .A(n7968), .B(n7967), .ZN(P1_U3239) );
  NAND2_X1 U9556 ( .A1(n7970), .A2(n7969), .ZN(n7972) );
  XNOR2_X1 U9557 ( .A(n7974), .B(n7973), .ZN(n9462) );
  AOI21_X1 U9558 ( .B1(n9458), .B2(n4573), .A(n8043), .ZN(n9459) );
  AOI22_X1 U9559 ( .A1(n9383), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9087), .B2(
        n9755), .ZN(n7976) );
  OAI21_X1 U9560 ( .B1(n9084), .B2(n9791), .A(n7976), .ZN(n7986) );
  NOR2_X1 U9561 ( .A1(n7981), .A2(n7980), .ZN(n8034) );
  AOI211_X1 U9562 ( .C1(n7981), .C2(n7980), .A(n9766), .B(n8034), .ZN(n7984)
         );
  OAI22_X1 U9563 ( .A1(n9784), .A2(n7982), .B1(n9083), .B2(n9781), .ZN(n7983)
         );
  NOR2_X1 U9564 ( .A1(n7984), .A2(n7983), .ZN(n9461) );
  NOR2_X1 U9565 ( .A1(n9461), .A2(n9383), .ZN(n7985) );
  AOI211_X1 U9566 ( .C1(n9459), .C2(n9777), .A(n7986), .B(n7985), .ZN(n7987)
         );
  OAI21_X1 U9567 ( .B1(n9462), .B2(n9387), .A(n7987), .ZN(P1_U3274) );
  NAND2_X1 U9568 ( .A1(n7988), .A2(n8612), .ZN(n7989) );
  AND2_X1 U9569 ( .A1(n10020), .A2(n8611), .ZN(n7997) );
  NAND2_X1 U9570 ( .A1(n8002), .A2(n7998), .ZN(n8178) );
  XNOR2_X1 U9571 ( .A(n8426), .B(n8610), .ZN(n8182) );
  NAND2_X1 U9572 ( .A1(n7992), .A2(n8182), .ZN(n7993) );
  NAND2_X1 U9573 ( .A1(n7994), .A2(n7993), .ZN(n9542) );
  NAND2_X1 U9574 ( .A1(n7996), .A2(n8175), .ZN(n9901) );
  OAI21_X1 U9575 ( .B1(n9901), .B2(n7997), .A(n8178), .ZN(n8066) );
  XNOR2_X1 U9576 ( .A(n8066), .B(n8182), .ZN(n8000) );
  OAI22_X1 U9577 ( .A1(n7998), .A2(n8905), .B1(n8904), .B2(n8907), .ZN(n7999)
         );
  AOI21_X1 U9578 ( .B1(n8000), .B2(n9922), .A(n7999), .ZN(n8001) );
  OAI21_X1 U9579 ( .B1(n9542), .B2(n8883), .A(n8001), .ZN(n9544) );
  NAND2_X1 U9580 ( .A1(n9544), .A2(n8916), .ZN(n8011) );
  NAND2_X1 U9581 ( .A1(n9912), .A2(n8426), .ZN(n8005) );
  NAND2_X1 U9582 ( .A1(n8928), .A2(n8005), .ZN(n9543) );
  INV_X1 U9583 ( .A(n9543), .ZN(n8009) );
  AOI22_X1 U9584 ( .A1(n8932), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n8006), .B2(
        n9925), .ZN(n8007) );
  OAI21_X1 U9585 ( .B1(n9906), .B2(n8003), .A(n8007), .ZN(n8008) );
  AOI21_X1 U9586 ( .B1(n8009), .B2(n8896), .A(n8008), .ZN(n8010) );
  OAI211_X1 U9587 ( .C1(n9542), .C2(n8893), .A(n8011), .B(n8010), .ZN(P2_U3283) );
  INV_X1 U9588 ( .A(n8012), .ZN(n8016) );
  OAI222_X1 U9589 ( .A1(P1_U3084), .A2(n8014), .B1(n4282), .B2(n8016), .C1(
        n8013), .C2(n9502), .ZN(P1_U3327) );
  OAI222_X1 U9590 ( .A1(P2_U3152), .A2(n8017), .B1(n9049), .B2(n8016), .C1(
        n8015), .C2(n9041), .ZN(P2_U3332) );
  OAI21_X1 U9591 ( .B1(n8020), .B2(n8019), .A(n8018), .ZN(n8021) );
  INV_X1 U9592 ( .A(n8021), .ZN(n8022) );
  OAI21_X1 U9593 ( .B1(n8023), .B2(n8022), .A(n9136), .ZN(n8028) );
  NAND2_X1 U9594 ( .A1(P1_U3084), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9680) );
  OAI21_X1 U9595 ( .B1(n9114), .B2(n7913), .A(n9680), .ZN(n8026) );
  NOR2_X1 U9596 ( .A1(n9127), .A2(n8024), .ZN(n8025) );
  AOI211_X1 U9597 ( .C1(n9145), .C2(n9149), .A(n8026), .B(n8025), .ZN(n8027)
         );
  OAI211_X1 U9598 ( .C1(n4571), .C2(n9148), .A(n8028), .B(n8027), .ZN(P1_U3224) );
  INV_X1 U9599 ( .A(n8029), .ZN(n8051) );
  NAND2_X1 U9600 ( .A1(n9496), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n8030) );
  OAI211_X1 U9601 ( .C1(n8051), .C2(n4282), .A(n8031), .B(n8030), .ZN(P1_U3326) );
  INV_X1 U9602 ( .A(n8032), .ZN(n8033) );
  NOR2_X1 U9603 ( .A1(n8034), .A2(n8033), .ZN(n8035) );
  OAI21_X1 U9604 ( .B1(n8041), .B2(n8035), .A(n9186), .ZN(n8036) );
  AOI222_X1 U9605 ( .A1(n9786), .A2(n8036), .B1(n9149), .B2(n9734), .C1(n9174), 
        .C2(n9736), .ZN(n9456) );
  OAI22_X1 U9606 ( .A1(n8039), .A2(n8038), .B1(n9458), .B2(n9149), .ZN(n8040)
         );
  AOI21_X1 U9607 ( .B1(n8041), .B2(n8040), .A(n9173), .ZN(n9452) );
  NAND2_X1 U9608 ( .A1(n9452), .A2(n8042), .ZN(n8050) );
  INV_X1 U9609 ( .A(n8043), .ZN(n8045) );
  NAND2_X1 U9610 ( .A1(n8043), .A2(n8046), .ZN(n9373) );
  INV_X1 U9611 ( .A(n9373), .ZN(n8044) );
  AOI21_X1 U9612 ( .B1(n9453), .B2(n8045), .A(n8044), .ZN(n9454) );
  NOR2_X1 U9613 ( .A1(n8046), .A2(n9791), .ZN(n8048) );
  OAI22_X1 U9614 ( .A1(n9797), .A2(n8283), .B1(n9126), .B2(n9792), .ZN(n8047)
         );
  AOI211_X1 U9615 ( .C1(n9454), .C2(n9777), .A(n8048), .B(n8047), .ZN(n8049)
         );
  OAI211_X1 U9616 ( .C1(n9568), .C2(n9456), .A(n8050), .B(n8049), .ZN(P1_U3273) );
  OAI222_X1 U9617 ( .A1(n9047), .A2(n8052), .B1(P2_U3152), .B2(n8264), .C1(
        n9049), .C2(n8051), .ZN(P2_U3331) );
  NAND2_X1 U9618 ( .A1(n8459), .A2(n8053), .ZN(n8055) );
  OAI211_X1 U9619 ( .C1(n9502), .C2(n8056), .A(n8055), .B(n8054), .ZN(P1_U3325) );
  OAI222_X1 U9620 ( .A1(n9047), .A2(n8058), .B1(n9049), .B2(n8057), .C1(n8122), 
        .C2(P2_U3152), .ZN(P2_U3336) );
  INV_X1 U9621 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8061) );
  INV_X1 U9622 ( .A(n8060), .ZN(n8388) );
  OAI222_X1 U9623 ( .A1(n9041), .A2(n8061), .B1(n9049), .B2(n8388), .C1(n8059), 
        .C2(P2_U3152), .ZN(P2_U3328) );
  NAND2_X1 U9624 ( .A1(n8060), .A2(n8084), .ZN(n8063) );
  OR2_X1 U9625 ( .A1(n6082), .A2(n8061), .ZN(n8062) );
  NOR2_X1 U9626 ( .A1(n8662), .A2(n8133), .ZN(n8082) );
  NAND2_X1 U9627 ( .A1(n9046), .A2(n8084), .ZN(n8065) );
  OR2_X1 U9628 ( .A1(n6082), .A2(n9048), .ZN(n8064) );
  NAND2_X1 U9629 ( .A1(n8947), .A2(n8081), .ZN(n8251) );
  NAND2_X1 U9630 ( .A1(n8066), .A2(n8182), .ZN(n8068) );
  NAND2_X1 U9631 ( .A1(n8426), .A2(n8067), .ZN(n8185) );
  NAND2_X1 U9632 ( .A1(n8068), .A2(n8185), .ZN(n8899) );
  NAND2_X1 U9633 ( .A1(n8927), .A2(n8904), .ZN(n8184) );
  NAND2_X1 U9634 ( .A1(n8911), .A2(n8877), .ZN(n8105) );
  INV_X1 U9635 ( .A(n8105), .ZN(n8190) );
  INV_X1 U9636 ( .A(n8191), .ZN(n8106) );
  NAND2_X1 U9637 ( .A1(n9015), .A2(n8860), .ZN(n8430) );
  OR2_X1 U9638 ( .A1(n9015), .A2(n8860), .ZN(n8069) );
  INV_X1 U9639 ( .A(n8860), .ZN(n8906) );
  AND2_X1 U9640 ( .A1(n9015), .A2(n8906), .ZN(n8193) );
  XNOR2_X1 U9641 ( .A(n9012), .B(n8850), .ZN(n8858) );
  NAND2_X1 U9642 ( .A1(n9005), .A2(n8832), .ZN(n8199) );
  AND2_X1 U9643 ( .A1(n8858), .A2(n8199), .ZN(n8070) );
  INV_X1 U9644 ( .A(n8850), .ZN(n8878) );
  OR2_X1 U9645 ( .A1(n9012), .A2(n8878), .ZN(n8847) );
  OR2_X1 U9646 ( .A1(n9005), .A2(n8832), .ZN(n8201) );
  AND2_X1 U9647 ( .A1(n8847), .A2(n8201), .ZN(n8071) );
  OR2_X1 U9648 ( .A1(n8200), .A2(n8071), .ZN(n8825) );
  OR2_X1 U9649 ( .A1(n9002), .A2(n8578), .ZN(n8202) );
  NAND2_X1 U9650 ( .A1(n9002), .A2(n8578), .ZN(n8806) );
  NAND2_X1 U9651 ( .A1(n8202), .A2(n8806), .ZN(n8829) );
  INV_X1 U9652 ( .A(n8829), .ZN(n8112) );
  AND2_X1 U9653 ( .A1(n8825), .A2(n8112), .ZN(n8072) );
  NAND2_X1 U9654 ( .A1(n8993), .A2(n8833), .ZN(n8210) );
  NAND2_X1 U9655 ( .A1(n8212), .A2(n8210), .ZN(n8090) );
  NOR2_X1 U9656 ( .A1(n8090), .A2(n4539), .ZN(n8073) );
  NAND2_X1 U9657 ( .A1(n8827), .A2(n8073), .ZN(n8074) );
  OR2_X1 U9658 ( .A1(n8988), .A2(n8431), .ZN(n8215) );
  NAND2_X1 U9659 ( .A1(n8988), .A2(n8431), .ZN(n8777) );
  NAND2_X1 U9660 ( .A1(n8215), .A2(n8777), .ZN(n8797) );
  NAND2_X1 U9661 ( .A1(n8983), .A2(n8757), .ZN(n8204) );
  NAND2_X1 U9662 ( .A1(n8214), .A2(n8204), .ZN(n8772) );
  INV_X1 U9663 ( .A(n8777), .ZN(n8211) );
  NOR2_X1 U9664 ( .A1(n8772), .A2(n8211), .ZN(n8075) );
  OR2_X1 U9665 ( .A1(n8975), .A2(n8746), .ZN(n8218) );
  NAND2_X1 U9666 ( .A1(n8975), .A2(n8746), .ZN(n8742) );
  NAND2_X1 U9667 ( .A1(n8218), .A2(n8742), .ZN(n8752) );
  OR2_X1 U9668 ( .A1(n8970), .A2(n8756), .ZN(n8224) );
  NAND2_X1 U9669 ( .A1(n8970), .A2(n8756), .ZN(n8225) );
  NAND2_X1 U9670 ( .A1(n8224), .A2(n8225), .ZN(n8736) );
  INV_X1 U9671 ( .A(n8742), .ZN(n8077) );
  NOR2_X1 U9672 ( .A1(n8736), .A2(n8077), .ZN(n8078) );
  NAND2_X1 U9673 ( .A1(n8966), .A2(n8745), .ZN(n8229) );
  INV_X1 U9674 ( .A(n8228), .ZN(n8079) );
  OR2_X1 U9675 ( .A1(n8961), .A2(n8693), .ZN(n8234) );
  NAND2_X1 U9676 ( .A1(n8961), .A2(n8693), .ZN(n8231) );
  NAND2_X1 U9677 ( .A1(n8709), .A2(n8710), .ZN(n8708) );
  NAND2_X1 U9678 ( .A1(n8708), .A2(n8231), .ZN(n8691) );
  OAI22_X1 U9679 ( .A1(n8691), .A2(n8690), .B1(n8586), .B2(n8957), .ZN(n8681)
         );
  NAND2_X1 U9680 ( .A1(n8950), .A2(n8694), .ZN(n8241) );
  NAND2_X1 U9681 ( .A1(n8681), .A2(n8238), .ZN(n8080) );
  NAND2_X1 U9682 ( .A1(n8080), .A2(n8242), .ZN(n8446) );
  OR2_X1 U9683 ( .A1(n8947), .A2(n8081), .ZN(n8244) );
  AOI211_X1 U9684 ( .C1(n8082), .C2(n8666), .A(n4531), .B(n8445), .ZN(n8083)
         );
  NAND2_X1 U9685 ( .A1(n9039), .A2(n8084), .ZN(n8086) );
  OR2_X1 U9686 ( .A1(n6082), .A2(n6665), .ZN(n8085) );
  INV_X1 U9687 ( .A(n8662), .ZN(n8087) );
  OR2_X1 U9688 ( .A1(n8938), .A2(n8087), .ZN(n8256) );
  NAND2_X1 U9689 ( .A1(n8666), .A2(n8449), .ZN(n8250) );
  NAND2_X1 U9690 ( .A1(n8938), .A2(n8087), .ZN(n8246) );
  NAND2_X1 U9691 ( .A1(n5760), .A2(n8089), .ZN(n8263) );
  AND2_X1 U9692 ( .A1(n8246), .A2(n4302), .ZN(n8253) );
  INV_X1 U9693 ( .A(n8736), .ZN(n8741) );
  NAND2_X1 U9694 ( .A1(n8201), .A2(n8199), .ZN(n8848) );
  INV_X1 U9695 ( .A(n8926), .ZN(n8109) );
  INV_X1 U9696 ( .A(n8091), .ZN(n8093) );
  NAND3_X1 U9697 ( .A1(n8094), .A2(n8093), .A3(n8092), .ZN(n8099) );
  NOR2_X1 U9698 ( .A1(n8095), .A2(n7612), .ZN(n8097) );
  INV_X1 U9699 ( .A(n8145), .ZN(n8096) );
  NAND4_X1 U9700 ( .A1(n8097), .A2(n9919), .A3(n8259), .A4(n8096), .ZN(n8098)
         );
  NOR2_X1 U9701 ( .A1(n8099), .A2(n8098), .ZN(n8101) );
  AND4_X1 U9702 ( .A1(n8101), .A2(n8100), .A3(n7682), .A4(n4588), .ZN(n8104)
         );
  NAND4_X1 U9703 ( .A1(n8104), .A2(n9908), .A3(n4834), .A4(n8103), .ZN(n8107)
         );
  NAND2_X1 U9704 ( .A1(n8106), .A2(n8105), .ZN(n8902) );
  NOR2_X1 U9705 ( .A1(n8107), .A2(n8902), .ZN(n8108) );
  NAND4_X1 U9706 ( .A1(n8875), .A2(n8109), .A3(n8108), .A4(n8182), .ZN(n8110)
         );
  NOR2_X1 U9707 ( .A1(n8848), .A2(n8110), .ZN(n8111) );
  NAND4_X1 U9708 ( .A1(n8817), .A2(n8112), .A3(n8111), .A4(n8858), .ZN(n8113)
         );
  NOR4_X1 U9709 ( .A1(n8752), .A2(n8772), .A3(n8797), .A4(n8113), .ZN(n8114)
         );
  NAND4_X1 U9710 ( .A1(n8710), .A2(n8437), .A3(n8741), .A4(n8114), .ZN(n8115)
         );
  NOR4_X1 U9711 ( .A1(n8447), .A2(n8680), .A3(n8690), .A4(n8115), .ZN(n8116)
         );
  NAND3_X1 U9712 ( .A1(n4330), .A2(n8253), .A3(n8116), .ZN(n8117) );
  XNOR2_X1 U9713 ( .A(n8117), .B(n5751), .ZN(n8119) );
  OAI22_X1 U9714 ( .A1(n8119), .A2(n8118), .B1(n8259), .B2(n8120), .ZN(n8262)
         );
  INV_X1 U9715 ( .A(n8120), .ZN(n8121) );
  NOR2_X1 U9716 ( .A1(n8121), .A2(n9953), .ZN(n8261) );
  NOR2_X1 U9717 ( .A1(n8133), .A2(n5751), .ZN(n8123) );
  INV_X1 U9718 ( .A(n8204), .ZN(n8207) );
  INV_X1 U9719 ( .A(n8875), .ZN(n8879) );
  AND2_X1 U9720 ( .A1(n8173), .A2(n8157), .ZN(n8124) );
  MUX2_X1 U9721 ( .A(n8164), .B(n8124), .S(n8257), .Z(n8125) );
  NAND2_X1 U9722 ( .A1(n8125), .A2(n8166), .ZN(n8174) );
  INV_X1 U9723 ( .A(n8149), .ZN(n8130) );
  NOR3_X1 U9724 ( .A1(n8132), .A2(n8131), .A3(n8130), .ZN(n8153) );
  NOR2_X1 U9725 ( .A1(n8145), .A2(n8133), .ZN(n8135) );
  OAI211_X1 U9726 ( .C1(n8135), .C2(n7081), .A(n8146), .B(n8134), .ZN(n8136)
         );
  NAND3_X1 U9727 ( .A1(n8136), .A2(n9918), .A3(n8257), .ZN(n8139) );
  NAND2_X1 U9728 ( .A1(n4860), .A2(n8137), .ZN(n8138) );
  AOI22_X1 U9729 ( .A1(n8139), .A2(n9919), .B1(n8257), .B2(n8138), .ZN(n8141)
         );
  NOR2_X1 U9730 ( .A1(n8141), .A2(n8140), .ZN(n8151) );
  AOI21_X1 U9731 ( .B1(n8142), .B2(n8154), .A(n8127), .ZN(n8150) );
  OAI211_X1 U9732 ( .C1(n8145), .C2(n8144), .A(n9918), .B(n8143), .ZN(n8147)
         );
  NAND3_X1 U9733 ( .A1(n8147), .A2(n8127), .A3(n8146), .ZN(n8148) );
  OAI211_X1 U9734 ( .C1(n8151), .C2(n8150), .A(n8149), .B(n8148), .ZN(n8152)
         );
  INV_X1 U9735 ( .A(n8177), .ZN(n8159) );
  INV_X1 U9736 ( .A(n8157), .ZN(n8158) );
  NOR3_X1 U9737 ( .A1(n8160), .A2(n8159), .A3(n8158), .ZN(n8171) );
  NAND2_X1 U9738 ( .A1(n8162), .A2(n4849), .ZN(n8165) );
  NAND3_X1 U9739 ( .A1(n8165), .A2(n8164), .A3(n8163), .ZN(n8169) );
  INV_X1 U9740 ( .A(n8174), .ZN(n8168) );
  INV_X1 U9741 ( .A(n8175), .ZN(n8167) );
  AOI211_X1 U9742 ( .C1(n8169), .C2(n8168), .A(n8167), .B(n4595), .ZN(n8170)
         );
  MUX2_X1 U9743 ( .A(n8171), .B(n8170), .S(n8257), .Z(n8172) );
  OAI21_X1 U9744 ( .B1(n8174), .B2(n8173), .A(n8172), .ZN(n8179) );
  NAND3_X1 U9745 ( .A1(n8179), .A2(n8180), .A3(n8175), .ZN(n8176) );
  NAND3_X1 U9746 ( .A1(n8179), .A2(n8178), .A3(n8177), .ZN(n8181) );
  INV_X1 U9747 ( .A(n8182), .ZN(n8183) );
  OAI21_X1 U9748 ( .B1(n8926), .B2(n8185), .A(n8184), .ZN(n8188) );
  NAND2_X1 U9749 ( .A1(n8003), .A2(n8610), .ZN(n8186) );
  OAI21_X1 U9750 ( .B1(n8926), .B2(n8186), .A(n8900), .ZN(n8187) );
  MUX2_X1 U9751 ( .A(n8188), .B(n8187), .S(n8257), .Z(n8189) );
  MUX2_X1 U9752 ( .A(n8191), .B(n8190), .S(n8257), .Z(n8192) );
  INV_X1 U9753 ( .A(n8847), .ZN(n8196) );
  INV_X1 U9754 ( .A(n9012), .ZN(n8872) );
  NAND2_X1 U9755 ( .A1(n8858), .A2(n8193), .ZN(n8194) );
  OAI211_X1 U9756 ( .C1(n8872), .C2(n8850), .A(n8199), .B(n8194), .ZN(n8195)
         );
  MUX2_X1 U9757 ( .A(n8196), .B(n8195), .S(n8127), .Z(n8197) );
  INV_X1 U9758 ( .A(n8199), .ZN(n8200) );
  NOR2_X1 U9759 ( .A1(n8209), .A2(n8200), .ZN(n8203) );
  NAND2_X1 U9760 ( .A1(n8202), .A2(n8201), .ZN(n8208) );
  MUX2_X1 U9761 ( .A(n8207), .B(n8206), .S(n8257), .Z(n8223) );
  OAI21_X1 U9762 ( .B1(n8209), .B2(n8208), .A(n8806), .ZN(n8213) );
  AOI211_X1 U9763 ( .C1(n8213), .C2(n8212), .A(n8211), .B(n4540), .ZN(n8217)
         );
  INV_X1 U9764 ( .A(n8215), .ZN(n8216) );
  NAND2_X1 U9765 ( .A1(n8741), .A2(n8218), .ZN(n8220) );
  NAND2_X1 U9766 ( .A1(n8225), .A2(n8742), .ZN(n8219) );
  MUX2_X1 U9767 ( .A(n8220), .B(n8219), .S(n8257), .Z(n8221) );
  MUX2_X1 U9768 ( .A(n8225), .B(n8224), .S(n8257), .Z(n8226) );
  OAI211_X1 U9769 ( .C1(n8228), .C2(n8257), .A(n8227), .B(n8234), .ZN(n8232)
         );
  NAND2_X1 U9770 ( .A1(n8231), .A2(n8229), .ZN(n8230) );
  AOI22_X1 U9771 ( .A1(n8232), .A2(n8231), .B1(n8257), .B2(n8230), .ZN(n8240)
         );
  INV_X1 U9772 ( .A(n8690), .ZN(n8233) );
  OAI21_X1 U9773 ( .B1(n8127), .B2(n8234), .A(n8233), .ZN(n8239) );
  INV_X1 U9774 ( .A(n8586), .ZN(n8712) );
  NAND2_X1 U9775 ( .A1(n8712), .A2(n8127), .ZN(n8236) );
  NAND2_X1 U9776 ( .A1(n8586), .A2(n8257), .ZN(n8235) );
  MUX2_X1 U9777 ( .A(n8236), .B(n8235), .S(n8957), .Z(n8237) );
  MUX2_X1 U9778 ( .A(n8242), .B(n8241), .S(n8127), .Z(n8243) );
  NAND2_X1 U9779 ( .A1(n8252), .A2(n8245), .ZN(n8248) );
  INV_X1 U9780 ( .A(n8246), .ZN(n8247) );
  AOI21_X1 U9781 ( .B1(n8248), .B2(n4330), .A(n8247), .ZN(n8249) );
  INV_X1 U9782 ( .A(n8256), .ZN(n8258) );
  NAND2_X1 U9783 ( .A1(n8258), .A2(n8257), .ZN(n8260) );
  INV_X1 U9784 ( .A(n9939), .ZN(n8266) );
  INV_X1 U9785 ( .A(n8264), .ZN(n8443) );
  NAND4_X1 U9786 ( .A1(n8266), .A2(n8265), .A3(n8443), .A4(n8861), .ZN(n8267)
         );
  OAI211_X1 U9787 ( .C1(n8268), .C2(n8270), .A(n8267), .B(P2_B_REG_SCAN_IN), 
        .ZN(n8269) );
  NAND2_X1 U9788 ( .A1(n8271), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n8272) );
  NAND2_X1 U9789 ( .A1(n8273), .A2(n8272), .ZN(n9640) );
  OR2_X1 U9790 ( .A1(n9645), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n8275) );
  NAND2_X1 U9791 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n9645), .ZN(n8274) );
  AND2_X1 U9792 ( .A1(n8275), .A2(n8274), .ZN(n9639) );
  AOI21_X1 U9793 ( .B1(n9645), .B2(P1_REG2_REG_13__SCAN_IN), .A(n9642), .ZN(
        n8276) );
  NOR2_X1 U9794 ( .A1(n8276), .A2(n9660), .ZN(n8277) );
  INV_X1 U9795 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n9654) );
  XNOR2_X1 U9796 ( .A(n9660), .B(n8276), .ZN(n9655) );
  NOR2_X1 U9797 ( .A1(n9654), .A2(n9655), .ZN(n9653) );
  INV_X1 U9798 ( .A(n8278), .ZN(n8279) );
  NAND2_X1 U9799 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n9687), .ZN(n8280) );
  OAI21_X1 U9800 ( .B1(n9687), .B2(P1_REG2_REG_16__SCAN_IN), .A(n8280), .ZN(
        n9683) );
  NOR2_X1 U9801 ( .A1(n9684), .A2(n9683), .ZN(n9682) );
  AOI21_X1 U9802 ( .B1(n9687), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9682), .ZN(
        n9696) );
  OR2_X1 U9803 ( .A1(n8288), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n8282) );
  NAND2_X1 U9804 ( .A1(n8288), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n8281) );
  NAND2_X1 U9805 ( .A1(n8282), .A2(n8281), .ZN(n9697) );
  NOR2_X1 U9806 ( .A1(n9696), .A2(n9697), .ZN(n9695) );
  AOI21_X1 U9807 ( .B1(n8288), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9695), .ZN(
        n9711) );
  OR2_X1 U9808 ( .A1(n8287), .A2(n8283), .ZN(n8285) );
  NAND2_X1 U9809 ( .A1(n8287), .A2(n8283), .ZN(n8284) );
  AND2_X1 U9810 ( .A1(n8285), .A2(n8284), .ZN(n9712) );
  NOR2_X1 U9811 ( .A1(n9711), .A2(n9712), .ZN(n9710) );
  AOI21_X1 U9812 ( .B1(P1_REG2_REG_18__SCAN_IN), .B2(n8287), .A(n9710), .ZN(
        n8286) );
  XNOR2_X1 U9813 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n8286), .ZN(n8306) );
  INV_X1 U9814 ( .A(n8306), .ZN(n8302) );
  INV_X1 U9815 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n8299) );
  XNOR2_X1 U9816 ( .A(n8287), .B(P1_REG1_REG_18__SCAN_IN), .ZN(n9722) );
  INV_X1 U9817 ( .A(n8288), .ZN(n9701) );
  XNOR2_X1 U9818 ( .A(n9701), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9706) );
  INV_X1 U9819 ( .A(n9687), .ZN(n8297) );
  XOR2_X1 U9820 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9687), .Z(n9691) );
  INV_X1 U9821 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9591) );
  INV_X1 U9822 ( .A(n9645), .ZN(n8293) );
  INV_X1 U9823 ( .A(n8289), .ZN(n8290) );
  AOI21_X1 U9824 ( .B1(n5328), .B2(n8291), .A(n8290), .ZN(n9648) );
  NOR2_X1 U9825 ( .A1(n9645), .A2(n9598), .ZN(n8292) );
  AOI21_X1 U9826 ( .B1(n9645), .B2(n9598), .A(n8292), .ZN(n9647) );
  NOR2_X1 U9827 ( .A1(n9648), .A2(n9647), .ZN(n9646) );
  AOI21_X1 U9828 ( .B1(n9598), .B2(n8293), .A(n9646), .ZN(n9664) );
  MUX2_X1 U9829 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9591), .S(n9660), .Z(n9663)
         );
  NOR2_X1 U9830 ( .A1(n9664), .A2(n9663), .ZN(n9662) );
  AOI21_X1 U9831 ( .B1(n9660), .B2(n9591), .A(n9662), .ZN(n8294) );
  XOR2_X1 U9832 ( .A(n9674), .B(n8294), .Z(n9675) );
  AOI22_X1 U9833 ( .A1(n9675), .A2(P1_REG1_REG_15__SCAN_IN), .B1(n9674), .B2(
        n8294), .ZN(n8295) );
  INV_X1 U9834 ( .A(n8295), .ZN(n9690) );
  NAND2_X1 U9835 ( .A1(n9691), .A2(n9690), .ZN(n9689) );
  OAI21_X1 U9836 ( .B1(n8297), .B2(n8296), .A(n9689), .ZN(n9705) );
  NAND2_X1 U9837 ( .A1(n9706), .A2(n9705), .ZN(n9703) );
  OAI21_X1 U9838 ( .B1(n9701), .B2(n8298), .A(n9703), .ZN(n9721) );
  NOR2_X1 U9839 ( .A1(n9722), .A2(n9721), .ZN(n9720) );
  AOI21_X1 U9840 ( .B1(n8299), .B2(n9718), .A(n9720), .ZN(n8301) );
  XOR2_X1 U9841 ( .A(n8301), .B(n8300), .Z(n8303) );
  AOI21_X1 U9842 ( .B1(n8303), .B2(n9704), .A(n9688), .ZN(n8304) );
  NAND2_X1 U9843 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9065) );
  OAI21_X1 U9844 ( .B1(n8310), .B2(n8308), .A(n8309), .ZN(n8311) );
  NAND2_X1 U9845 ( .A1(n8311), .A2(n9136), .ZN(n8319) );
  INV_X1 U9846 ( .A(n8312), .ZN(n8317) );
  OR2_X1 U9847 ( .A1(n9114), .A2(n5181), .ZN(n8314) );
  AND2_X1 U9848 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n8365) );
  INV_X1 U9849 ( .A(n8365), .ZN(n8313) );
  OAI211_X1 U9850 ( .C1(n8315), .C2(n9123), .A(n8314), .B(n8313), .ZN(n8316)
         );
  AOI21_X1 U9851 ( .B1(n8317), .B2(n9140), .A(n8316), .ZN(n8318) );
  OAI211_X1 U9852 ( .C1(n9849), .C2(n9148), .A(n8319), .B(n8318), .ZN(P1_U3211) );
  NAND2_X1 U9853 ( .A1(n9092), .A2(n9091), .ZN(n9090) );
  NAND2_X1 U9854 ( .A1(n9090), .A2(n8320), .ZN(n8321) );
  OAI21_X1 U9855 ( .B1(n8322), .B2(n8321), .A(n9134), .ZN(n8323) );
  NAND2_X1 U9856 ( .A1(n8323), .A2(n9136), .ZN(n8327) );
  AOI22_X1 U9857 ( .A1(n9283), .A2(n9139), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3084), .ZN(n8324) );
  OAI21_X1 U9858 ( .B1(n9127), .B2(n9277), .A(n8324), .ZN(n8325) );
  AOI21_X1 U9859 ( .B1(n9284), .B2(n9145), .A(n8325), .ZN(n8326) );
  OAI211_X1 U9860 ( .C1(n9280), .C2(n9148), .A(n8327), .B(n8326), .ZN(P1_U3223) );
  AOI21_X1 U9861 ( .B1(n8330), .B2(n8329), .A(n8328), .ZN(n8341) );
  OAI21_X1 U9862 ( .B1(n8333), .B2(n8332), .A(n8331), .ZN(n8339) );
  INV_X1 U9863 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n8337) );
  NAND2_X1 U9864 ( .A1(n9688), .A2(n8334), .ZN(n8335) );
  OAI211_X1 U9865 ( .C1(n9727), .C2(n8337), .A(n8336), .B(n8335), .ZN(n8338)
         );
  AOI21_X1 U9866 ( .B1(n8339), .B2(n9714), .A(n8338), .ZN(n8340) );
  OAI21_X1 U9867 ( .B1(n8341), .B2(n9724), .A(n8340), .ZN(P1_U3252) );
  INV_X1 U9868 ( .A(n8342), .ZN(n8343) );
  AOI21_X1 U9869 ( .B1(n8345), .B2(n8344), .A(n8343), .ZN(n8355) );
  INV_X1 U9870 ( .A(n8346), .ZN(n8347) );
  OAI21_X1 U9871 ( .B1(n9717), .B2(n8348), .A(n8347), .ZN(n8353) );
  AOI211_X1 U9872 ( .C1(n8351), .C2(n8350), .A(n9681), .B(n8349), .ZN(n8352)
         );
  AOI211_X1 U9873 ( .C1(n8367), .C2(P1_ADDR_REG_10__SCAN_IN), .A(n8353), .B(
        n8352), .ZN(n8354) );
  OAI21_X1 U9874 ( .B1(n8355), .B2(n9724), .A(n8354), .ZN(P1_U3251) );
  INV_X1 U9875 ( .A(n8356), .ZN(n8357) );
  AOI21_X1 U9876 ( .B1(n8359), .B2(n8358), .A(n8357), .ZN(n8370) );
  OAI21_X1 U9877 ( .B1(n8362), .B2(n8361), .A(n8360), .ZN(n8366) );
  NOR2_X1 U9878 ( .A1(n9717), .A2(n8363), .ZN(n8364) );
  AOI211_X1 U9879 ( .C1(n9704), .C2(n8366), .A(n8365), .B(n8364), .ZN(n8369)
         );
  NAND2_X1 U9880 ( .A1(n8367), .A2(P1_ADDR_REG_7__SCAN_IN), .ZN(n8368) );
  OAI211_X1 U9881 ( .C1(n8370), .C2(n9681), .A(n8369), .B(n8368), .ZN(P1_U3248) );
  AOI22_X1 U9882 ( .A1(n8514), .A2(n7071), .B1(n8488), .B2(n8371), .ZN(n8384)
         );
  AND2_X1 U9883 ( .A1(P2_U3152), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n9517) );
  AOI21_X1 U9884 ( .B1(n8418), .B2(P2_REG3_REG_2__SCAN_IN), .A(n9517), .ZN(
        n8375) );
  NAND2_X1 U9885 ( .A1(n8589), .A2(n8373), .ZN(n8374) );
  OAI211_X1 U9886 ( .C1(n8597), .C2(n7074), .A(n8375), .B(n8374), .ZN(n8382)
         );
  INV_X1 U9887 ( .A(n8376), .ZN(n8379) );
  OAI211_X1 U9888 ( .C1(n8379), .C2(n8378), .A(n8488), .B(n8377), .ZN(n8380)
         );
  OAI21_X1 U9889 ( .B1(n8598), .B2(n8413), .A(n8380), .ZN(n8381) );
  NOR2_X1 U9890 ( .A1(n8382), .A2(n8381), .ZN(n8383) );
  OAI21_X1 U9891 ( .B1(n8384), .B2(n8372), .A(n8383), .ZN(P2_U3239) );
  OAI222_X1 U9892 ( .A1(n9502), .A2(n8386), .B1(n4282), .B2(n8385), .C1(n5658), 
        .C2(P1_U3084), .ZN(P1_U3333) );
  OAI222_X1 U9893 ( .A1(P1_U3084), .A2(n8389), .B1(n4282), .B2(n8388), .C1(
        n8387), .C2(n9502), .ZN(P1_U3323) );
  AOI22_X1 U9894 ( .A1(n8514), .A2(n8618), .B1(n8488), .B2(n8391), .ZN(n8393)
         );
  NOR2_X1 U9895 ( .A1(n8393), .A2(n8392), .ZN(n8403) );
  INV_X1 U9896 ( .A(n8394), .ZN(n8395) );
  OAI22_X1 U9897 ( .A1(n8597), .A2(n8396), .B1(n8585), .B2(n8395), .ZN(n8401)
         );
  AOI21_X1 U9898 ( .B1(n8589), .B2(n8398), .A(n8397), .ZN(n8399) );
  OAI21_X1 U9899 ( .B1(n8598), .B2(n7079), .A(n8399), .ZN(n8400) );
  AOI211_X1 U9900 ( .C1(n8403), .C2(n8402), .A(n8401), .B(n8400), .ZN(n8404)
         );
  OAI21_X1 U9901 ( .B1(n8405), .B2(n8593), .A(n8404), .ZN(P2_U3241) );
  INV_X1 U9902 ( .A(n9952), .ZN(n8406) );
  OAI22_X1 U9903 ( .A1(n8592), .A2(n8425), .B1(n8406), .B2(n8593), .ZN(n8408)
         );
  NAND2_X1 U9904 ( .A1(n8408), .A2(n8407), .ZN(n8412) );
  NAND2_X1 U9905 ( .A1(n8418), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n8409) );
  NAND2_X1 U9906 ( .A1(P2_U3152), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n9890) );
  NAND2_X1 U9907 ( .A1(n8409), .A2(n9890), .ZN(n8410) );
  AOI21_X1 U9908 ( .B1(n8589), .B2(n9952), .A(n8410), .ZN(n8411) );
  OAI211_X1 U9909 ( .C1(n8413), .C2(n8597), .A(n8412), .B(n8411), .ZN(P2_U3234) );
  AOI22_X1 U9910 ( .A1(n8565), .A2(n7071), .B1(n8414), .B2(n8589), .ZN(n8424)
         );
  OAI21_X1 U9911 ( .B1(n8417), .B2(n8416), .A(n8415), .ZN(n8422) );
  INV_X1 U9912 ( .A(n8418), .ZN(n8420) );
  INV_X1 U9913 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n8419) );
  NAND2_X1 U9914 ( .A1(P2_U3152), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n9503) );
  OAI21_X1 U9915 ( .B1(n8420), .B2(n8419), .A(n9503), .ZN(n8421) );
  AOI21_X1 U9916 ( .B1(n8488), .B2(n8422), .A(n8421), .ZN(n8423) );
  OAI211_X1 U9917 ( .C1(n8425), .C2(n8598), .A(n8424), .B(n8423), .ZN(P2_U3224) );
  NAND2_X1 U9918 ( .A1(n8924), .A2(n8926), .ZN(n8925) );
  INV_X1 U9919 ( .A(n8904), .ZN(n8609) );
  OR2_X1 U9920 ( .A1(n8927), .A2(n8609), .ZN(n8428) );
  NAND2_X1 U9921 ( .A1(n8925), .A2(n8428), .ZN(n8898) );
  INV_X1 U9922 ( .A(n8877), .ZN(n8608) );
  NOR2_X1 U9923 ( .A1(n8911), .A2(n8608), .ZN(n8429) );
  AOI21_X1 U9924 ( .B1(n8898), .B2(n8902), .A(n8429), .ZN(n8880) );
  NAND2_X1 U9925 ( .A1(n8880), .A2(n8879), .ZN(n8882) );
  NAND2_X1 U9926 ( .A1(n8882), .A2(n8430), .ZN(n8856) );
  NOR2_X1 U9927 ( .A1(n9005), .A2(n8863), .ZN(n8821) );
  OR2_X1 U9928 ( .A1(n8821), .A2(n4854), .ZN(n8814) );
  OR2_X1 U9929 ( .A1(n8814), .A2(n8817), .ZN(n8786) );
  OR2_X1 U9930 ( .A1(n8786), .A2(n4859), .ZN(n8436) );
  NAND2_X1 U9931 ( .A1(n9005), .A2(n8863), .ZN(n8822) );
  AND2_X1 U9932 ( .A1(n4853), .A2(n8822), .ZN(n8432) );
  OR2_X1 U9933 ( .A1(n4854), .A2(n8432), .ZN(n8815) );
  OR2_X1 U9934 ( .A1(n8817), .A2(n8815), .ZN(n8787) );
  INV_X1 U9935 ( .A(n8833), .ZN(n8800) );
  NAND2_X1 U9936 ( .A1(n8993), .A2(n8800), .ZN(n8789) );
  NAND2_X1 U9937 ( .A1(n8988), .A2(n8808), .ZN(n8433) );
  AND2_X1 U9938 ( .A1(n8789), .A2(n8433), .ZN(n8434) );
  AND2_X1 U9939 ( .A1(n8787), .A2(n8434), .ZN(n8435) );
  INV_X1 U9940 ( .A(n8772), .ZN(n8778) );
  INV_X1 U9941 ( .A(n8757), .ZN(n8801) );
  OAI21_X1 U9942 ( .B1(n8767), .B2(n8746), .A(n8762), .ZN(n8735) );
  INV_X1 U9943 ( .A(n8756), .ZN(n8607) );
  NAND2_X1 U9944 ( .A1(n8723), .A2(n8728), .ZN(n8722) );
  INV_X1 U9945 ( .A(n8745), .ZN(n8711) );
  NAND2_X1 U9946 ( .A1(n8722), .A2(n8438), .ZN(n8706) );
  NAND2_X1 U9947 ( .A1(n8671), .A2(n8680), .ZN(n8672) );
  INV_X1 U9948 ( .A(n8694), .ZN(n8605) );
  NAND2_X1 U9949 ( .A1(n8672), .A2(n8440), .ZN(n8442) );
  XNOR2_X1 U9950 ( .A(n8442), .B(n8441), .ZN(n8949) );
  NAND2_X1 U9951 ( .A1(n8443), .A2(P2_B_REG_SCAN_IN), .ZN(n8444) );
  NAND2_X1 U9952 ( .A1(n8862), .A2(n8444), .ZN(n8660) );
  AOI21_X1 U9953 ( .B1(n8447), .B2(n8446), .A(n8445), .ZN(n8448) );
  OAI222_X1 U9954 ( .A1(n8905), .A2(n8694), .B1(n8660), .B2(n8449), .C1(n8448), 
        .C2(n8920), .ZN(n8948) );
  INV_X1 U9955 ( .A(n8947), .ZN(n8456) );
  INV_X1 U9956 ( .A(n9015), .ZN(n8892) );
  INV_X1 U9957 ( .A(n9002), .ZN(n8450) );
  NAND2_X1 U9958 ( .A1(n8773), .A2(n8767), .ZN(n8763) );
  INV_X1 U9959 ( .A(n8957), .ZN(n8701) );
  NAND2_X1 U9960 ( .A1(n8714), .A2(n8701), .ZN(n8695) );
  NOR2_X2 U9961 ( .A1(n8674), .A2(n8947), .ZN(n8665) );
  AOI211_X1 U9962 ( .C1(n8947), .C2(n8674), .A(n10004), .B(n8665), .ZN(n8946)
         );
  NAND2_X1 U9963 ( .A1(n8946), .A2(n9933), .ZN(n8455) );
  INV_X1 U9964 ( .A(n8452), .ZN(n8453) );
  AOI22_X1 U9965 ( .A1(n9937), .A2(P2_REG2_REG_29__SCAN_IN), .B1(n8453), .B2(
        n9925), .ZN(n8454) );
  OAI211_X1 U9966 ( .C1(n8456), .C2(n9906), .A(n8455), .B(n8454), .ZN(n8457)
         );
  AOI21_X1 U9967 ( .B1(n8948), .B2(n8916), .A(n8457), .ZN(n8458) );
  OAI21_X1 U9968 ( .B1(n8949), .B2(n8918), .A(n8458), .ZN(P2_U3267) );
  INV_X1 U9969 ( .A(n8459), .ZN(n8460) );
  XNOR2_X1 U9970 ( .A(n8463), .B(n8462), .ZN(n8469) );
  INV_X1 U9971 ( .A(n8698), .ZN(n8465) );
  OAI22_X1 U9972 ( .A1(n8585), .A2(n8465), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8464), .ZN(n8467) );
  OAI22_X1 U9973 ( .A1(n8693), .A2(n8598), .B1(n8597), .B2(n8694), .ZN(n8466)
         );
  AOI211_X1 U9974 ( .C1(n8957), .C2(n8589), .A(n8467), .B(n8466), .ZN(n8468)
         );
  OAI21_X1 U9975 ( .B1(n8469), .B2(n8593), .A(n8468), .ZN(P2_U3216) );
  INV_X1 U9976 ( .A(n8746), .ZN(n8780) );
  AOI22_X1 U9977 ( .A1(n8470), .A2(n8488), .B1(n8514), .B2(n8780), .ZN(n8479)
         );
  INV_X1 U9978 ( .A(n8471), .ZN(n8472) );
  NAND2_X1 U9979 ( .A1(n8470), .A2(n8472), .ZN(n8540) );
  INV_X1 U9980 ( .A(n8540), .ZN(n8478) );
  INV_X1 U9981 ( .A(n8765), .ZN(n8474) );
  OAI22_X1 U9982 ( .A1(n8585), .A2(n8474), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8473), .ZN(n8476) );
  OAI22_X1 U9983 ( .A1(n8757), .A2(n8598), .B1(n8597), .B2(n8756), .ZN(n8475)
         );
  AOI211_X1 U9984 ( .C1(n8975), .C2(n8589), .A(n8476), .B(n8475), .ZN(n8477)
         );
  OAI21_X1 U9985 ( .B1(n8479), .B2(n8478), .A(n8477), .ZN(P2_U3218) );
  OAI22_X1 U9986 ( .A1(n8480), .A2(n8907), .B1(n7072), .B2(n8905), .ZN(n9921)
         );
  AOI22_X1 U9987 ( .A1(n9932), .A2(n8589), .B1(n8509), .B2(n9921), .ZN(n8485)
         );
  MUX2_X1 U9988 ( .A(n8585), .B(P2_STATE_REG_SCAN_IN), .S(
        P2_REG3_REG_3__SCAN_IN), .Z(n8484) );
  OAI211_X1 U9989 ( .C1(n8482), .C2(n8372), .A(n8488), .B(n8481), .ZN(n8483)
         );
  NAND3_X1 U9990 ( .A1(n8485), .A2(n8484), .A3(n8483), .ZN(P2_U3220) );
  OAI21_X1 U9991 ( .B1(n8493), .B2(n8486), .A(n8487), .ZN(n8489) );
  NAND2_X1 U9992 ( .A1(n8489), .A2(n8488), .ZN(n8497) );
  AOI22_X1 U9993 ( .A1(n8601), .A2(n8837), .B1(P2_REG3_REG_19__SCAN_IN), .B2(
        P2_U3152), .ZN(n8490) );
  OAI21_X1 U9994 ( .B1(n8833), .B2(n8597), .A(n8490), .ZN(n8491) );
  AOI21_X1 U9995 ( .B1(n9002), .B2(n8589), .A(n8491), .ZN(n8496) );
  NOR3_X1 U9996 ( .A1(n8493), .A2(n8492), .A3(n8592), .ZN(n8494) );
  OAI21_X1 U9997 ( .B1(n8494), .B2(n8566), .A(n8863), .ZN(n8495) );
  NAND3_X1 U9998 ( .A1(n8497), .A2(n8496), .A3(n8495), .ZN(P2_U3221) );
  INV_X1 U9999 ( .A(n8499), .ZN(n8500) );
  AOI21_X1 U10000 ( .B1(n8498), .B2(n8500), .A(n8593), .ZN(n8504) );
  NOR3_X1 U10001 ( .A1(n8501), .A2(n8833), .A3(n8592), .ZN(n8503) );
  OAI21_X1 U10002 ( .B1(n8504), .B2(n8503), .A(n8502), .ZN(n8508) );
  AOI22_X1 U10003 ( .A1(n8601), .A2(n8794), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3152), .ZN(n8507) );
  AOI22_X1 U10004 ( .A1(n8566), .A2(n8800), .B1(n8565), .B2(n8801), .ZN(n8506)
         );
  NAND2_X1 U10005 ( .A1(n8988), .A2(n8589), .ZN(n8505) );
  NAND4_X1 U10006 ( .A1(n8508), .A2(n8507), .A3(n8506), .A4(n8505), .ZN(
        P2_U3225) );
  INV_X1 U10007 ( .A(n8726), .ZN(n8511) );
  OAI22_X1 U10008 ( .A1(n8693), .A2(n8907), .B1(n8756), .B2(n8905), .ZN(n8730)
         );
  AOI22_X1 U10009 ( .A1(n8509), .A2(n8730), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3152), .ZN(n8510) );
  OAI21_X1 U10010 ( .B1(n8511), .B2(n8585), .A(n8510), .ZN(n8520) );
  INV_X1 U10011 ( .A(n8517), .ZN(n8513) );
  NAND3_X1 U10012 ( .A1(n8515), .A2(n8514), .A3(n8711), .ZN(n8516) );
  OAI21_X1 U10013 ( .B1(n8517), .B2(n8593), .A(n8516), .ZN(n8519) );
  INV_X1 U10014 ( .A(n8521), .ZN(n8522) );
  AOI21_X1 U10015 ( .B1(n8524), .B2(n8523), .A(n8522), .ZN(n8529) );
  INV_X1 U10016 ( .A(n8890), .ZN(n8525) );
  OAI22_X1 U10017 ( .A1(n8585), .A2(n8525), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8626), .ZN(n8527) );
  OAI22_X1 U10018 ( .A1(n8877), .A2(n8598), .B1(n8597), .B2(n8878), .ZN(n8526)
         );
  AOI211_X1 U10019 ( .C1(n9015), .C2(n8589), .A(n8527), .B(n8526), .ZN(n8528)
         );
  OAI21_X1 U10020 ( .B1(n8529), .B2(n8593), .A(n8528), .ZN(P2_U3228) );
  NAND2_X1 U10021 ( .A1(n8532), .A2(n8531), .ZN(n8536) );
  NOR2_X1 U10022 ( .A1(n8533), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8639) );
  OAI22_X1 U10023 ( .A1(n8906), .A2(n8598), .B1(n8597), .B2(n8832), .ZN(n8534)
         );
  AOI211_X1 U10024 ( .C1(n8601), .C2(n8869), .A(n8639), .B(n8534), .ZN(n8535)
         );
  OAI211_X1 U10025 ( .C1(n8872), .C2(n8604), .A(n8536), .B(n8535), .ZN(
        P2_U3230) );
  NAND2_X1 U10026 ( .A1(n8538), .A2(n8537), .ZN(n8539) );
  NAND2_X1 U10027 ( .A1(n8540), .A2(n8539), .ZN(n8542) );
  XNOR2_X1 U10028 ( .A(n8542), .B(n8541), .ZN(n8545) );
  OAI22_X1 U10029 ( .A1(n8545), .A2(n8593), .B1(n8756), .B2(n8592), .ZN(n8543)
         );
  OAI21_X1 U10030 ( .B1(n8545), .B2(n8544), .A(n8543), .ZN(n8550) );
  NOR2_X1 U10031 ( .A1(n8546), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8548) );
  OAI22_X1 U10032 ( .A1(n8746), .A2(n8598), .B1(n8597), .B2(n8745), .ZN(n8547)
         );
  AOI211_X1 U10033 ( .C1(n8601), .C2(n8738), .A(n8548), .B(n8547), .ZN(n8549)
         );
  OAI211_X1 U10034 ( .C1(n4480), .C2(n8604), .A(n8550), .B(n8549), .ZN(
        P2_U3231) );
  INV_X1 U10035 ( .A(n8498), .ZN(n8551) );
  AOI211_X1 U10036 ( .C1(n8553), .C2(n8552), .A(n8593), .B(n8551), .ZN(n8557)
         );
  INV_X1 U10037 ( .A(n8993), .ZN(n8812) );
  AOI22_X1 U10038 ( .A1(n8601), .A2(n8810), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3152), .ZN(n8555) );
  AOI22_X1 U10039 ( .A1(n8565), .A2(n8808), .B1(n8566), .B2(n8851), .ZN(n8554)
         );
  OAI211_X1 U10040 ( .C1(n8812), .C2(n8604), .A(n8555), .B(n8554), .ZN(n8556)
         );
  OR2_X1 U10041 ( .A1(n8557), .A2(n8556), .ZN(P2_U3235) );
  INV_X1 U10042 ( .A(n8558), .ZN(n8559) );
  NAND2_X1 U10043 ( .A1(n8502), .A2(n8559), .ZN(n8561) );
  XNOR2_X1 U10044 ( .A(n8561), .B(n8560), .ZN(n8562) );
  NOR3_X1 U10045 ( .A1(n8562), .A2(n8757), .A3(n8592), .ZN(n8571) );
  INV_X1 U10046 ( .A(n8562), .ZN(n8564) );
  NOR3_X1 U10047 ( .A1(n8564), .A2(n8563), .A3(n8593), .ZN(n8570) );
  INV_X1 U10048 ( .A(n8983), .ZN(n8776) );
  AOI22_X1 U10049 ( .A1(n8601), .A2(n8774), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3152), .ZN(n8568) );
  AOI22_X1 U10050 ( .A1(n8566), .A2(n8808), .B1(n8565), .B2(n8780), .ZN(n8567)
         );
  OAI211_X1 U10051 ( .C1(n8776), .C2(n8604), .A(n8568), .B(n8567), .ZN(n8569)
         );
  OR3_X1 U10052 ( .A1(n8571), .A2(n8570), .A3(n8569), .ZN(P2_U3237) );
  INV_X1 U10053 ( .A(n9005), .ZN(n8846) );
  INV_X1 U10054 ( .A(n8572), .ZN(n8573) );
  AOI21_X1 U10055 ( .B1(n8531), .B2(n8573), .A(n8593), .ZN(n8576) );
  NOR3_X1 U10056 ( .A1(n8574), .A2(n8878), .A3(n8592), .ZN(n8575) );
  OAI21_X1 U10057 ( .B1(n8576), .B2(n8575), .A(n8486), .ZN(n8581) );
  NOR2_X1 U10058 ( .A1(n8577), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8656) );
  OAI22_X1 U10059 ( .A1(n8878), .A2(n8598), .B1(n8597), .B2(n8578), .ZN(n8579)
         );
  AOI211_X1 U10060 ( .C1(n8601), .C2(n8844), .A(n8656), .B(n8579), .ZN(n8580)
         );
  OAI211_X1 U10061 ( .C1(n8846), .C2(n8604), .A(n8581), .B(n8580), .ZN(
        P2_U3240) );
  XNOR2_X1 U10062 ( .A(n8583), .B(n8582), .ZN(n8591) );
  OAI22_X1 U10063 ( .A1(n8585), .A2(n8717), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8584), .ZN(n8588) );
  OAI22_X1 U10064 ( .A1(n8745), .A2(n8598), .B1(n8597), .B2(n8586), .ZN(n8587)
         );
  AOI211_X1 U10065 ( .C1(n8961), .C2(n8589), .A(n8588), .B(n8587), .ZN(n8590)
         );
  OAI21_X1 U10066 ( .B1(n8591), .B2(n8593), .A(n8590), .ZN(P2_U3242) );
  OAI22_X1 U10067 ( .A1(n8594), .A2(n8593), .B1(n8877), .B2(n8592), .ZN(n8596)
         );
  NAND2_X1 U10068 ( .A1(n8596), .A2(n8595), .ZN(n8603) );
  OAI22_X1 U10069 ( .A1(n8904), .A2(n8598), .B1(n8597), .B2(n8906), .ZN(n8599)
         );
  AOI211_X1 U10070 ( .C1(n8601), .C2(n8910), .A(n8600), .B(n8599), .ZN(n8602)
         );
  OAI211_X1 U10071 ( .C1(n9529), .C2(n8604), .A(n8603), .B(n8602), .ZN(
        P2_U3243) );
  MUX2_X1 U10072 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n8605), .S(P2_U3966), .Z(
        P2_U3580) );
  MUX2_X1 U10073 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8712), .S(P2_U3966), .Z(
        P2_U3579) );
  MUX2_X1 U10074 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n8606), .S(P2_U3966), .Z(
        P2_U3578) );
  MUX2_X1 U10075 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8711), .S(P2_U3966), .Z(
        P2_U3577) );
  MUX2_X1 U10076 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8607), .S(P2_U3966), .Z(
        P2_U3576) );
  MUX2_X1 U10077 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n8780), .S(P2_U3966), .Z(
        P2_U3575) );
  MUX2_X1 U10078 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8801), .S(P2_U3966), .Z(
        P2_U3574) );
  MUX2_X1 U10079 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8808), .S(P2_U3966), .Z(
        P2_U3573) );
  MUX2_X1 U10080 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8800), .S(P2_U3966), .Z(
        P2_U3572) );
  MUX2_X1 U10081 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8851), .S(P2_U3966), .Z(
        P2_U3571) );
  MUX2_X1 U10082 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8863), .S(P2_U3966), .Z(
        P2_U3570) );
  MUX2_X1 U10083 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8850), .S(P2_U3966), .Z(
        P2_U3569) );
  MUX2_X1 U10084 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8860), .S(P2_U3966), .Z(
        P2_U3568) );
  MUX2_X1 U10085 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8608), .S(P2_U3966), .Z(
        P2_U3567) );
  MUX2_X1 U10086 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8609), .S(P2_U3966), .Z(
        P2_U3566) );
  MUX2_X1 U10087 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n8610), .S(P2_U3966), .Z(
        P2_U3565) );
  MUX2_X1 U10088 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n8611), .S(P2_U3966), .Z(
        P2_U3564) );
  MUX2_X1 U10089 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n8612), .S(P2_U3966), .Z(
        P2_U3563) );
  MUX2_X1 U10090 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n8613), .S(P2_U3966), .Z(
        P2_U3562) );
  MUX2_X1 U10091 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n8614), .S(P2_U3966), .Z(
        P2_U3561) );
  MUX2_X1 U10092 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n8615), .S(P2_U3966), .Z(
        P2_U3560) );
  MUX2_X1 U10093 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n8616), .S(P2_U3966), .Z(
        P2_U3559) );
  MUX2_X1 U10094 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n8617), .S(P2_U3966), .Z(
        P2_U3558) );
  MUX2_X1 U10095 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n8618), .S(P2_U3966), .Z(
        P2_U3557) );
  MUX2_X1 U10096 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n8619), .S(P2_U3966), .Z(
        P2_U3556) );
  MUX2_X1 U10097 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n8620), .S(P2_U3966), .Z(
        P2_U3555) );
  MUX2_X1 U10098 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n7071), .S(P2_U3966), .Z(
        P2_U3554) );
  MUX2_X1 U10099 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n8621), .S(P2_U3966), .Z(
        P2_U3553) );
  MUX2_X1 U10100 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n8622), .S(P2_U3966), .Z(
        P2_U3552) );
  AOI21_X1 U10101 ( .B1(n8625), .B2(n8624), .A(n8623), .ZN(n8631) );
  NOR2_X1 U10102 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8626), .ZN(n8627) );
  AOI21_X1 U10103 ( .B1(n9892), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n8627), .ZN(
        n8630) );
  NAND2_X1 U10104 ( .A1(n9522), .A2(n8628), .ZN(n8629) );
  OAI211_X1 U10105 ( .C1(n8631), .C2(n9894), .A(n8630), .B(n8629), .ZN(n8636)
         );
  AOI211_X1 U10106 ( .C1(n8634), .C2(n8633), .A(n8632), .B(n9895), .ZN(n8635)
         );
  OR2_X1 U10107 ( .A1(n8636), .A2(n8635), .ZN(P2_U3261) );
  AOI211_X1 U10108 ( .C1(n4367), .C2(n8638), .A(n8637), .B(n9895), .ZN(n8646)
         );
  AOI21_X1 U10109 ( .B1(n9892), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n8639), .ZN(
        n8643) );
  OAI211_X1 U10110 ( .C1(n8641), .C2(n4846), .A(n9888), .B(n8640), .ZN(n8642)
         );
  OAI211_X1 U10111 ( .C1(n9893), .C2(n8644), .A(n8643), .B(n8642), .ZN(n8645)
         );
  OR2_X1 U10112 ( .A1(n8646), .A2(n8645), .ZN(P2_U3262) );
  AOI21_X1 U10113 ( .B1(n8649), .B2(n8648), .A(n8647), .ZN(n8659) );
  OAI21_X1 U10114 ( .B1(n8652), .B2(n8651), .A(n8650), .ZN(n8653) );
  NAND2_X1 U10115 ( .A1(n8653), .A2(n9889), .ZN(n8658) );
  NOR2_X1 U10116 ( .A1(n9893), .A2(n8654), .ZN(n8655) );
  AOI211_X1 U10117 ( .C1(n9892), .C2(P2_ADDR_REG_18__SCAN_IN), .A(n8656), .B(
        n8655), .ZN(n8657) );
  OAI211_X1 U10118 ( .C1(n8659), .C2(n9894), .A(n8658), .B(n8657), .ZN(
        P2_U3263) );
  NAND2_X1 U10119 ( .A1(n8665), .A2(n8945), .ZN(n8942) );
  XNOR2_X1 U10120 ( .A(n8942), .B(n8938), .ZN(n8940) );
  INV_X1 U10121 ( .A(n8660), .ZN(n8661) );
  NAND2_X1 U10122 ( .A1(n8662), .A2(n8661), .ZN(n8943) );
  NOR2_X1 U10123 ( .A1(n9937), .A2(n8943), .ZN(n8668) );
  AOI21_X1 U10124 ( .B1(n9937), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8668), .ZN(
        n8664) );
  NAND2_X1 U10125 ( .A1(n8938), .A2(n9931), .ZN(n8663) );
  OAI211_X1 U10126 ( .C1(n8940), .C2(n8914), .A(n8664), .B(n8663), .ZN(
        P2_U3265) );
  INV_X1 U10127 ( .A(n8665), .ZN(n8667) );
  NAND2_X1 U10128 ( .A1(n8667), .A2(n8666), .ZN(n8941) );
  NAND3_X1 U10129 ( .A1(n8942), .A2(n8896), .A3(n8941), .ZN(n8670) );
  AOI21_X1 U10130 ( .B1(n9937), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8668), .ZN(
        n8669) );
  OAI211_X1 U10131 ( .C1(n8945), .C2(n9906), .A(n8670), .B(n8669), .ZN(
        P2_U3266) );
  OAI21_X1 U10132 ( .B1(n8671), .B2(n8680), .A(n8672), .ZN(n8673) );
  INV_X1 U10133 ( .A(n8673), .ZN(n8954) );
  INV_X1 U10134 ( .A(n8674), .ZN(n8675) );
  AOI21_X1 U10135 ( .B1(n8950), .B2(n8695), .A(n8675), .ZN(n8951) );
  INV_X1 U10136 ( .A(n8676), .ZN(n8677) );
  AOI22_X1 U10137 ( .A1(n8932), .A2(P2_REG2_REG_28__SCAN_IN), .B1(n8677), .B2(
        n9925), .ZN(n8678) );
  OAI21_X1 U10138 ( .B1(n8679), .B2(n9906), .A(n8678), .ZN(n8685) );
  XNOR2_X1 U10139 ( .A(n8681), .B(n8680), .ZN(n8683) );
  AOI21_X1 U10140 ( .B1(n8683), .B2(n9922), .A(n8682), .ZN(n8953) );
  NOR2_X1 U10141 ( .A1(n8953), .A2(n8932), .ZN(n8684) );
  AOI211_X1 U10142 ( .C1(n8951), .C2(n8896), .A(n8685), .B(n8684), .ZN(n8686)
         );
  OAI21_X1 U10143 ( .B1(n8954), .B2(n8918), .A(n8686), .ZN(P2_U3268) );
  OAI21_X1 U10144 ( .B1(n8688), .B2(n8690), .A(n8687), .ZN(n8689) );
  INV_X1 U10145 ( .A(n8689), .ZN(n8959) );
  XNOR2_X1 U10146 ( .A(n8691), .B(n8690), .ZN(n8692) );
  OAI222_X1 U10147 ( .A1(n8907), .A2(n8694), .B1(n8905), .B2(n8693), .C1(n8920), .C2(n8692), .ZN(n8955) );
  INV_X1 U10148 ( .A(n8714), .ZN(n8697) );
  INV_X1 U10149 ( .A(n8695), .ZN(n8696) );
  AOI211_X1 U10150 ( .C1(n8957), .C2(n8697), .A(n10004), .B(n8696), .ZN(n8956)
         );
  NAND2_X1 U10151 ( .A1(n8956), .A2(n9933), .ZN(n8700) );
  AOI22_X1 U10152 ( .A1(n8932), .A2(P2_REG2_REG_27__SCAN_IN), .B1(n8698), .B2(
        n9925), .ZN(n8699) );
  OAI211_X1 U10153 ( .C1(n8701), .C2(n9906), .A(n8700), .B(n8699), .ZN(n8702)
         );
  AOI21_X1 U10154 ( .B1(n8955), .B2(n8916), .A(n8702), .ZN(n8703) );
  OAI21_X1 U10155 ( .B1(n8959), .B2(n8918), .A(n8703), .ZN(P2_U3269) );
  OAI21_X1 U10156 ( .B1(n8706), .B2(n8705), .A(n8704), .ZN(n8707) );
  INV_X1 U10157 ( .A(n8707), .ZN(n8964) );
  AOI22_X1 U10158 ( .A1(n8961), .A2(n9931), .B1(n9937), .B2(
        P2_REG2_REG_26__SCAN_IN), .ZN(n8721) );
  OAI21_X1 U10159 ( .B1(n8710), .B2(n8709), .A(n8708), .ZN(n8713) );
  AOI222_X1 U10160 ( .A1(n9922), .A2(n8713), .B1(n8712), .B2(n8862), .C1(n8711), .C2(n8861), .ZN(n8963) );
  INV_X1 U10161 ( .A(n8725), .ZN(n8715) );
  AOI211_X1 U10162 ( .C1(n8961), .C2(n8715), .A(n10004), .B(n8714), .ZN(n8960)
         );
  NAND2_X1 U10163 ( .A1(n8960), .A2(n5751), .ZN(n8716) );
  OAI211_X1 U10164 ( .C1(n8718), .C2(n8717), .A(n8963), .B(n8716), .ZN(n8719)
         );
  NAND2_X1 U10165 ( .A1(n8719), .A2(n8916), .ZN(n8720) );
  OAI211_X1 U10166 ( .C1(n8964), .C2(n8918), .A(n8721), .B(n8720), .ZN(
        P2_U3270) );
  OAI21_X1 U10167 ( .B1(n8723), .B2(n8728), .A(n8722), .ZN(n8724) );
  INV_X1 U10168 ( .A(n8724), .ZN(n8969) );
  AOI211_X1 U10169 ( .C1(n8966), .C2(n8737), .A(n10004), .B(n8725), .ZN(n8965)
         );
  AOI22_X1 U10170 ( .A1(n8932), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n8726), .B2(
        n9925), .ZN(n8727) );
  OAI21_X1 U10171 ( .B1(n4481), .B2(n9906), .A(n8727), .ZN(n8733) );
  XNOR2_X1 U10172 ( .A(n8729), .B(n8728), .ZN(n8731) );
  AOI21_X1 U10173 ( .B1(n8731), .B2(n9922), .A(n8730), .ZN(n8968) );
  NOR2_X1 U10174 ( .A1(n8968), .A2(n9937), .ZN(n8732) );
  AOI211_X1 U10175 ( .C1(n8965), .C2(n8868), .A(n8733), .B(n8732), .ZN(n8734)
         );
  OAI21_X1 U10176 ( .B1(n8969), .B2(n8918), .A(n8734), .ZN(P2_U3271) );
  XNOR2_X1 U10177 ( .A(n8735), .B(n8736), .ZN(n8974) );
  AOI21_X1 U10178 ( .B1(n8970), .B2(n8763), .A(n8451), .ZN(n8971) );
  AOI22_X1 U10179 ( .A1(n8932), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n8738), .B2(
        n9925), .ZN(n8739) );
  OAI21_X1 U10180 ( .B1(n4480), .B2(n9906), .A(n8739), .ZN(n8750) );
  INV_X1 U10181 ( .A(n8740), .ZN(n8744) );
  AOI21_X1 U10182 ( .B1(n8755), .B2(n8742), .A(n8741), .ZN(n8743) );
  NOR3_X1 U10183 ( .A1(n8744), .A2(n8743), .A3(n8920), .ZN(n8748) );
  OAI22_X1 U10184 ( .A1(n8746), .A2(n8905), .B1(n8745), .B2(n8907), .ZN(n8747)
         );
  NOR2_X1 U10185 ( .A1(n8748), .A2(n8747), .ZN(n8973) );
  NOR2_X1 U10186 ( .A1(n8973), .A2(n9937), .ZN(n8749) );
  AOI211_X1 U10187 ( .C1(n8971), .C2(n8896), .A(n8750), .B(n8749), .ZN(n8751)
         );
  OAI21_X1 U10188 ( .B1(n8918), .B2(n8974), .A(n8751), .ZN(P2_U3272) );
  NAND2_X1 U10189 ( .A1(n8753), .A2(n8752), .ZN(n8754) );
  NAND2_X1 U10190 ( .A1(n8755), .A2(n8754), .ZN(n8759) );
  OAI22_X1 U10191 ( .A1(n8757), .A2(n8905), .B1(n8756), .B2(n8907), .ZN(n8758)
         );
  AOI21_X1 U10192 ( .B1(n8759), .B2(n9922), .A(n8758), .ZN(n8978) );
  NAND2_X1 U10193 ( .A1(n8760), .A2(n8076), .ZN(n8761) );
  AND2_X1 U10194 ( .A1(n8762), .A2(n8761), .ZN(n8980) );
  NAND2_X1 U10195 ( .A1(n8980), .A2(n9934), .ZN(n8770) );
  OR2_X1 U10196 ( .A1(n8773), .A2(n8767), .ZN(n8764) );
  AND2_X1 U10197 ( .A1(n8764), .A2(n8763), .ZN(n8976) );
  AOI22_X1 U10198 ( .A1(n9937), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n8765), .B2(
        n9925), .ZN(n8766) );
  OAI21_X1 U10199 ( .B1(n8767), .B2(n9906), .A(n8766), .ZN(n8768) );
  AOI21_X1 U10200 ( .B1(n8976), .B2(n8896), .A(n8768), .ZN(n8769) );
  OAI211_X1 U10201 ( .C1(n9937), .C2(n8978), .A(n8770), .B(n8769), .ZN(
        P2_U3273) );
  XNOR2_X1 U10202 ( .A(n8771), .B(n8772), .ZN(n8987) );
  AOI21_X1 U10203 ( .B1(n8983), .B2(n8792), .A(n8773), .ZN(n8984) );
  AOI22_X1 U10204 ( .A1(n8932), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8774), .B2(
        n9925), .ZN(n8775) );
  OAI21_X1 U10205 ( .B1(n8776), .B2(n9906), .A(n8775), .ZN(n8783) );
  NAND2_X1 U10206 ( .A1(n8798), .A2(n8777), .ZN(n8779) );
  XNOR2_X1 U10207 ( .A(n8779), .B(n8778), .ZN(n8781) );
  AOI222_X1 U10208 ( .A1(n9922), .A2(n8781), .B1(n8780), .B2(n8862), .C1(n8808), .C2(n8861), .ZN(n8986) );
  NOR2_X1 U10209 ( .A1(n8986), .A2(n9937), .ZN(n8782) );
  AOI211_X1 U10210 ( .C1(n8984), .C2(n8896), .A(n8783), .B(n8782), .ZN(n8784)
         );
  OAI21_X1 U10211 ( .B1(n8918), .B2(n8987), .A(n8784), .ZN(P2_U3274) );
  OR2_X1 U10212 ( .A1(n8785), .A2(n8786), .ZN(n8788) );
  NAND2_X1 U10213 ( .A1(n8996), .A2(n8789), .ZN(n8790) );
  XNOR2_X1 U10214 ( .A(n8790), .B(n8797), .ZN(n8992) );
  INV_X1 U10215 ( .A(n8792), .ZN(n8793) );
  AOI21_X1 U10216 ( .B1(n8988), .B2(n4475), .A(n8793), .ZN(n8989) );
  INV_X1 U10217 ( .A(n8988), .ZN(n8796) );
  AOI22_X1 U10218 ( .A1(n8932), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8794), .B2(
        n9925), .ZN(n8795) );
  OAI21_X1 U10219 ( .B1(n8796), .B2(n9906), .A(n8795), .ZN(n8804) );
  INV_X1 U10220 ( .A(n8797), .ZN(n8799) );
  OAI21_X1 U10221 ( .B1(n4334), .B2(n8799), .A(n8798), .ZN(n8802) );
  AOI222_X1 U10222 ( .A1(n9922), .A2(n8802), .B1(n8801), .B2(n8862), .C1(n8800), .C2(n8861), .ZN(n8991) );
  NOR2_X1 U10223 ( .A1(n8991), .A2(n9937), .ZN(n8803) );
  AOI211_X1 U10224 ( .C1(n8989), .C2(n8896), .A(n8804), .B(n8803), .ZN(n8805)
         );
  OAI21_X1 U10225 ( .B1(n8918), .B2(n8992), .A(n8805), .ZN(P2_U3275) );
  NAND2_X1 U10226 ( .A1(n8827), .A2(n8806), .ZN(n8807) );
  XNOR2_X1 U10227 ( .A(n8807), .B(n8817), .ZN(n8809) );
  AOI222_X1 U10228 ( .A1(n9922), .A2(n8809), .B1(n8851), .B2(n8861), .C1(n8808), .C2(n8862), .ZN(n8999) );
  AOI21_X1 U10229 ( .B1(n8993), .B2(n8834), .A(n8791), .ZN(n8994) );
  AOI22_X1 U10230 ( .A1(n8932), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8810), .B2(
        n9925), .ZN(n8811) );
  OAI21_X1 U10231 ( .B1(n8812), .B2(n9906), .A(n8811), .ZN(n8813) );
  AOI21_X1 U10232 ( .B1(n8994), .B2(n8896), .A(n8813), .ZN(n8820) );
  OR2_X1 U10233 ( .A1(n8785), .A2(n8814), .ZN(n8816) );
  AND2_X1 U10234 ( .A1(n8816), .A2(n8815), .ZN(n8818) );
  NAND2_X1 U10235 ( .A1(n8818), .A2(n8817), .ZN(n8995) );
  NAND3_X1 U10236 ( .A1(n8996), .A2(n8995), .A3(n9934), .ZN(n8819) );
  OAI211_X1 U10237 ( .C1(n8999), .C2(n8932), .A(n8820), .B(n8819), .ZN(
        P2_U3276) );
  OR2_X1 U10238 ( .A1(n8785), .A2(n8821), .ZN(n8823) );
  NAND2_X1 U10239 ( .A1(n8823), .A2(n8822), .ZN(n8824) );
  XNOR2_X1 U10240 ( .A(n8824), .B(n8829), .ZN(n9004) );
  NAND2_X1 U10241 ( .A1(n8826), .A2(n8825), .ZN(n8830) );
  INV_X1 U10242 ( .A(n8827), .ZN(n8828) );
  AOI21_X1 U10243 ( .B1(n8830), .B2(n8829), .A(n8828), .ZN(n8831) );
  OAI222_X1 U10244 ( .A1(n8907), .A2(n8833), .B1(n8905), .B2(n8832), .C1(n8920), .C2(n8831), .ZN(n9000) );
  INV_X1 U10245 ( .A(n9000), .ZN(n8839) );
  INV_X1 U10246 ( .A(n8843), .ZN(n8836) );
  INV_X1 U10247 ( .A(n8834), .ZN(n8835) );
  AOI211_X1 U10248 ( .C1(n9002), .C2(n8836), .A(n10004), .B(n8835), .ZN(n9001)
         );
  AOI22_X1 U10249 ( .A1(n9001), .A2(n5751), .B1(n9925), .B2(n8837), .ZN(n8838)
         );
  OAI211_X1 U10250 ( .C1(n8883), .C2(n9004), .A(n8839), .B(n8838), .ZN(n8840)
         );
  NAND2_X1 U10251 ( .A1(n8840), .A2(n8916), .ZN(n8842) );
  AOI22_X1 U10252 ( .A1(n9002), .A2(n9931), .B1(n9937), .B2(
        P2_REG2_REG_19__SCAN_IN), .ZN(n8841) );
  OAI211_X1 U10253 ( .C1(n9004), .C2(n8893), .A(n8842), .B(n8841), .ZN(
        P2_U3277) );
  XOR2_X1 U10254 ( .A(n8848), .B(n8785), .Z(n9009) );
  AOI21_X1 U10255 ( .B1(n9005), .B2(n8866), .A(n8843), .ZN(n9006) );
  AOI22_X1 U10256 ( .A1(n8932), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8844), .B2(
        n9925), .ZN(n8845) );
  OAI21_X1 U10257 ( .B1(n8846), .B2(n9906), .A(n8845), .ZN(n8854) );
  NAND2_X1 U10258 ( .A1(n8859), .A2(n8858), .ZN(n8857) );
  NAND2_X1 U10259 ( .A1(n8857), .A2(n8847), .ZN(n8849) );
  XNOR2_X1 U10260 ( .A(n8849), .B(n8848), .ZN(n8852) );
  AOI222_X1 U10261 ( .A1(n9922), .A2(n8852), .B1(n8851), .B2(n8862), .C1(n8850), .C2(n8861), .ZN(n9008) );
  NOR2_X1 U10262 ( .A1(n9008), .A2(n8932), .ZN(n8853) );
  AOI211_X1 U10263 ( .C1(n9006), .C2(n8896), .A(n8854), .B(n8853), .ZN(n8855)
         );
  OAI21_X1 U10264 ( .B1(n9009), .B2(n8918), .A(n8855), .ZN(P2_U3278) );
  XOR2_X1 U10265 ( .A(n8856), .B(n8858), .Z(n9014) );
  OAI211_X1 U10266 ( .C1(n8859), .C2(n8858), .A(n8857), .B(n9922), .ZN(n8865)
         );
  AOI22_X1 U10267 ( .A1(n8863), .A2(n8862), .B1(n8861), .B2(n8860), .ZN(n8864)
         );
  NAND2_X1 U10268 ( .A1(n8865), .A2(n8864), .ZN(n9010) );
  INV_X1 U10269 ( .A(n8866), .ZN(n8867) );
  AOI211_X1 U10270 ( .C1(n9012), .C2(n8887), .A(n10004), .B(n8867), .ZN(n9011)
         );
  NAND2_X1 U10271 ( .A1(n9011), .A2(n8868), .ZN(n8871) );
  AOI22_X1 U10272 ( .A1(n8932), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n8869), .B2(
        n9925), .ZN(n8870) );
  OAI211_X1 U10273 ( .C1(n8872), .C2(n9906), .A(n8871), .B(n8870), .ZN(n8873)
         );
  AOI21_X1 U10274 ( .B1(n9010), .B2(n8916), .A(n8873), .ZN(n8874) );
  OAI21_X1 U10275 ( .B1(n9014), .B2(n8918), .A(n8874), .ZN(P2_U3279) );
  XNOR2_X1 U10276 ( .A(n8876), .B(n8875), .ZN(n8886) );
  OAI22_X1 U10277 ( .A1(n8878), .A2(n8907), .B1(n8877), .B2(n8905), .ZN(n8885)
         );
  OR2_X1 U10278 ( .A1(n8880), .A2(n8879), .ZN(n8881) );
  NAND2_X1 U10279 ( .A1(n8882), .A2(n8881), .ZN(n9020) );
  NOR2_X1 U10280 ( .A1(n9020), .A2(n8883), .ZN(n8884) );
  AOI211_X1 U10281 ( .C1(n9922), .C2(n8886), .A(n8885), .B(n8884), .ZN(n9019)
         );
  INV_X1 U10282 ( .A(n8909), .ZN(n8889) );
  INV_X1 U10283 ( .A(n8887), .ZN(n8888) );
  AOI21_X1 U10284 ( .B1(n9015), .B2(n8889), .A(n8888), .ZN(n9017) );
  AOI22_X1 U10285 ( .A1(n8932), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n8890), .B2(
        n9925), .ZN(n8891) );
  OAI21_X1 U10286 ( .B1(n8892), .B2(n9906), .A(n8891), .ZN(n8895) );
  NOR2_X1 U10287 ( .A1(n9020), .A2(n8893), .ZN(n8894) );
  AOI211_X1 U10288 ( .C1(n9017), .C2(n8896), .A(n8895), .B(n8894), .ZN(n8897)
         );
  OAI21_X1 U10289 ( .B1(n9019), .B2(n8932), .A(n8897), .ZN(P2_U3280) );
  XNOR2_X1 U10290 ( .A(n8898), .B(n8902), .ZN(n9533) );
  INV_X1 U10291 ( .A(n9533), .ZN(n8919) );
  OR2_X1 U10292 ( .A1(n8899), .A2(n8926), .ZN(n8922) );
  NAND2_X1 U10293 ( .A1(n8922), .A2(n8900), .ZN(n8901) );
  XOR2_X1 U10294 ( .A(n8902), .B(n8901), .Z(n8903) );
  OAI222_X1 U10295 ( .A1(n8907), .A2(n8906), .B1(n8905), .B2(n8904), .C1(n8920), .C2(n8903), .ZN(n9531) );
  NOR2_X1 U10296 ( .A1(n8929), .A2(n9529), .ZN(n8908) );
  OR2_X1 U10297 ( .A1(n8909), .A2(n8908), .ZN(n9530) );
  AOI22_X1 U10298 ( .A1(n8932), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n8910), .B2(
        n9925), .ZN(n8913) );
  NAND2_X1 U10299 ( .A1(n9931), .A2(n8911), .ZN(n8912) );
  OAI211_X1 U10300 ( .C1(n9530), .C2(n8914), .A(n8913), .B(n8912), .ZN(n8915)
         );
  AOI21_X1 U10301 ( .B1(n9531), .B2(n8916), .A(n8915), .ZN(n8917) );
  OAI21_X1 U10302 ( .B1(n8919), .B2(n8918), .A(n8917), .ZN(P2_U3281) );
  AOI21_X1 U10303 ( .B1(n8899), .B2(n8926), .A(n8920), .ZN(n8923) );
  AOI21_X1 U10304 ( .B1(n8923), .B2(n8922), .A(n8921), .ZN(n9536) );
  OAI21_X1 U10305 ( .B1(n8924), .B2(n8926), .A(n8925), .ZN(n9539) );
  NAND2_X1 U10306 ( .A1(n9539), .A2(n9934), .ZN(n8937) );
  INV_X1 U10307 ( .A(n8927), .ZN(n9537) );
  INV_X1 U10308 ( .A(n8928), .ZN(n8930) );
  OAI211_X1 U10309 ( .C1(n9537), .C2(n8930), .A(n4471), .B(n9913), .ZN(n9535)
         );
  INV_X1 U10310 ( .A(n9535), .ZN(n8935) );
  AOI22_X1 U10311 ( .A1(n8932), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n8931), .B2(
        n9925), .ZN(n8933) );
  OAI21_X1 U10312 ( .B1(n9906), .B2(n9537), .A(n8933), .ZN(n8934) );
  AOI21_X1 U10313 ( .B1(n8935), .B2(n9933), .A(n8934), .ZN(n8936) );
  OAI211_X1 U10314 ( .C1(n9536), .C2(n9937), .A(n8937), .B(n8936), .ZN(
        P2_U3282) );
  NAND2_X1 U10315 ( .A1(n8938), .A2(n9016), .ZN(n8939) );
  OAI211_X1 U10316 ( .C1(n8940), .C2(n10004), .A(n8939), .B(n8943), .ZN(n9021)
         );
  MUX2_X1 U10317 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n9021), .S(n10045), .Z(
        P2_U3551) );
  NAND3_X1 U10318 ( .A1(n8942), .A2(n9913), .A3(n8941), .ZN(n8944) );
  OAI211_X1 U10319 ( .C1(n8945), .C2(n10019), .A(n8944), .B(n8943), .ZN(n9022)
         );
  MUX2_X1 U10320 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n9022), .S(n10045), .Z(
        P2_U3550) );
  MUX2_X1 U10321 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n9023), .S(n10045), .Z(
        P2_U3549) );
  AOI22_X1 U10322 ( .A1(n8951), .A2(n9913), .B1(n9016), .B2(n8950), .ZN(n8952)
         );
  OAI211_X1 U10323 ( .C1(n8954), .C2(n10001), .A(n8953), .B(n8952), .ZN(n9024)
         );
  MUX2_X1 U10324 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n9024), .S(n10045), .Z(
        P2_U3548) );
  AOI211_X1 U10325 ( .C1(n9016), .C2(n8957), .A(n8956), .B(n8955), .ZN(n8958)
         );
  OAI21_X1 U10326 ( .B1(n8959), .B2(n10001), .A(n8958), .ZN(n9025) );
  MUX2_X1 U10327 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n9025), .S(n10045), .Z(
        P2_U3547) );
  AOI21_X1 U10328 ( .B1(n9016), .B2(n8961), .A(n8960), .ZN(n8962) );
  OAI211_X1 U10329 ( .C1(n8964), .C2(n10001), .A(n8963), .B(n8962), .ZN(n9026)
         );
  MUX2_X1 U10330 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n9026), .S(n10045), .Z(
        P2_U3546) );
  AOI21_X1 U10331 ( .B1(n9016), .B2(n8966), .A(n8965), .ZN(n8967) );
  OAI211_X1 U10332 ( .C1(n8969), .C2(n10001), .A(n8968), .B(n8967), .ZN(n9027)
         );
  MUX2_X1 U10333 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n9027), .S(n10045), .Z(
        P2_U3545) );
  AOI22_X1 U10334 ( .A1(n8971), .A2(n9913), .B1(n9016), .B2(n8970), .ZN(n8972)
         );
  OAI211_X1 U10335 ( .C1(n8974), .C2(n10001), .A(n8973), .B(n8972), .ZN(n9028)
         );
  MUX2_X1 U10336 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n9028), .S(n10045), .Z(
        P2_U3544) );
  INV_X1 U10337 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8981) );
  AOI22_X1 U10338 ( .A1(n8976), .A2(n9913), .B1(n9016), .B2(n8975), .ZN(n8977)
         );
  NAND2_X1 U10339 ( .A1(n8978), .A2(n8977), .ZN(n8979) );
  AOI21_X1 U10340 ( .B1(n8980), .B2(n10025), .A(n8979), .ZN(n9029) );
  MUX2_X1 U10341 ( .A(n8981), .B(n9029), .S(n10045), .Z(n8982) );
  INV_X1 U10342 ( .A(n8982), .ZN(P2_U3543) );
  AOI22_X1 U10343 ( .A1(n8984), .A2(n9913), .B1(n9016), .B2(n8983), .ZN(n8985)
         );
  OAI211_X1 U10344 ( .C1(n10001), .C2(n8987), .A(n8986), .B(n8985), .ZN(n9032)
         );
  MUX2_X1 U10345 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n9032), .S(n10045), .Z(
        P2_U3542) );
  AOI22_X1 U10346 ( .A1(n8989), .A2(n9913), .B1(n9016), .B2(n8988), .ZN(n8990)
         );
  OAI211_X1 U10347 ( .C1(n10001), .C2(n8992), .A(n8991), .B(n8990), .ZN(n9033)
         );
  MUX2_X1 U10348 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n9033), .S(n10045), .Z(
        P2_U3541) );
  AOI22_X1 U10349 ( .A1(n8994), .A2(n9913), .B1(n9016), .B2(n8993), .ZN(n8998)
         );
  NAND3_X1 U10350 ( .A1(n8996), .A2(n10025), .A3(n8995), .ZN(n8997) );
  NAND3_X1 U10351 ( .A1(n8999), .A2(n8998), .A3(n8997), .ZN(n9034) );
  MUX2_X1 U10352 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n9034), .S(n10045), .Z(
        P2_U3540) );
  AOI211_X1 U10353 ( .C1(n9016), .C2(n9002), .A(n9001), .B(n9000), .ZN(n9003)
         );
  OAI21_X1 U10354 ( .B1(n10001), .B2(n9004), .A(n9003), .ZN(n9035) );
  MUX2_X1 U10355 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n9035), .S(n10045), .Z(
        P2_U3539) );
  AOI22_X1 U10356 ( .A1(n9006), .A2(n9913), .B1(n9016), .B2(n9005), .ZN(n9007)
         );
  OAI211_X1 U10357 ( .C1(n9009), .C2(n10001), .A(n9008), .B(n9007), .ZN(n9036)
         );
  MUX2_X1 U10358 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n9036), .S(n10045), .Z(
        P2_U3538) );
  AOI211_X1 U10359 ( .C1(n9016), .C2(n9012), .A(n9011), .B(n9010), .ZN(n9013)
         );
  OAI21_X1 U10360 ( .B1(n10001), .B2(n9014), .A(n9013), .ZN(n9037) );
  MUX2_X1 U10361 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n9037), .S(n10045), .Z(
        P2_U3537) );
  AOI22_X1 U10362 ( .A1(n9017), .A2(n9913), .B1(n9016), .B2(n9015), .ZN(n9018)
         );
  OAI211_X1 U10363 ( .C1(n9541), .C2(n9020), .A(n9019), .B(n9018), .ZN(n9038)
         );
  MUX2_X1 U10364 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n9038), .S(n10045), .Z(
        P2_U3536) );
  MUX2_X1 U10365 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n9021), .S(n10028), .Z(
        P2_U3519) );
  MUX2_X1 U10366 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n9022), .S(n10028), .Z(
        P2_U3518) );
  MUX2_X1 U10367 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n9023), .S(n10028), .Z(
        P2_U3517) );
  MUX2_X1 U10368 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n9024), .S(n10028), .Z(
        P2_U3516) );
  MUX2_X1 U10369 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n9025), .S(n10028), .Z(
        P2_U3515) );
  MUX2_X1 U10370 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n9026), .S(n10028), .Z(
        P2_U3514) );
  MUX2_X1 U10371 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n9027), .S(n10028), .Z(
        P2_U3513) );
  MUX2_X1 U10372 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n9028), .S(n10028), .Z(
        P2_U3512) );
  INV_X1 U10373 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n9030) );
  MUX2_X1 U10374 ( .A(n9030), .B(n9029), .S(n10028), .Z(n9031) );
  INV_X1 U10375 ( .A(n9031), .ZN(P2_U3511) );
  MUX2_X1 U10376 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n9032), .S(n10028), .Z(
        P2_U3510) );
  MUX2_X1 U10377 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n9033), .S(n10028), .Z(
        P2_U3509) );
  MUX2_X1 U10378 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n9034), .S(n10028), .Z(
        P2_U3508) );
  MUX2_X1 U10379 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n9035), .S(n10028), .Z(
        P2_U3507) );
  MUX2_X1 U10380 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n9036), .S(n10028), .Z(
        P2_U3505) );
  MUX2_X1 U10381 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n9037), .S(n10028), .Z(
        P2_U3502) );
  MUX2_X1 U10382 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n9038), .S(n10028), .Z(
        P2_U3499) );
  INV_X1 U10383 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n9040) );
  NAND3_X1 U10384 ( .A1(n9040), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n9042) );
  OAI22_X1 U10385 ( .A1(n5733), .A2(n9042), .B1(n6665), .B2(n9041), .ZN(n9043)
         );
  AOI21_X1 U10386 ( .B1(n9039), .B2(n9044), .A(n9043), .ZN(n9045) );
  INV_X1 U10387 ( .A(n9045), .ZN(P2_U3327) );
  INV_X1 U10388 ( .A(n9046), .ZN(n9500) );
  OAI222_X1 U10389 ( .A1(P2_U3152), .A2(n9050), .B1(n9049), .B2(n9500), .C1(
        n9048), .C2(n9047), .ZN(P2_U3329) );
  MUX2_X1 U10390 ( .A(n9052), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  INV_X1 U10391 ( .A(n9053), .ZN(n9055) );
  NOR2_X1 U10392 ( .A1(n9055), .A2(n9054), .ZN(n9057) );
  XNOR2_X1 U10393 ( .A(n9057), .B(n9056), .ZN(n9062) );
  NAND2_X1 U10394 ( .A1(n9283), .A2(n9145), .ZN(n9059) );
  AOI22_X1 U10395 ( .A1(n9346), .A2(n9139), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3084), .ZN(n9058) );
  OAI211_X1 U10396 ( .C1(n9127), .C2(n9308), .A(n9059), .B(n9058), .ZN(n9060)
         );
  AOI21_X1 U10397 ( .B1(n9429), .B2(n9129), .A(n9060), .ZN(n9061) );
  OAI21_X1 U10398 ( .B1(n9062), .B2(n9131), .A(n9061), .ZN(P1_U3214) );
  AOI21_X1 U10399 ( .B1(n9064), .B2(n9063), .A(n9101), .ZN(n9070) );
  OAI21_X1 U10400 ( .B1(n9123), .B2(n9177), .A(n9065), .ZN(n9066) );
  AOI21_X1 U10401 ( .B1(n9139), .B2(n9380), .A(n9066), .ZN(n9067) );
  OAI21_X1 U10402 ( .B1(n9127), .B2(n9374), .A(n9067), .ZN(n9068) );
  AOI21_X1 U10403 ( .B1(n9447), .B2(n9129), .A(n9068), .ZN(n9069) );
  OAI21_X1 U10404 ( .B1(n9070), .B2(n9131), .A(n9069), .ZN(P1_U3217) );
  OAI21_X1 U10405 ( .B1(n9073), .B2(n9072), .A(n9071), .ZN(n9074) );
  NAND2_X1 U10406 ( .A1(n9074), .A2(n9136), .ZN(n9078) );
  AOI22_X1 U10407 ( .A1(n9139), .A2(n9381), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3084), .ZN(n9075) );
  OAI21_X1 U10408 ( .B1(n9315), .B2(n9123), .A(n9075), .ZN(n9076) );
  AOI21_X1 U10409 ( .B1(n9339), .B2(n9140), .A(n9076), .ZN(n9077) );
  OAI211_X1 U10410 ( .C1(n9341), .C2(n9148), .A(n9078), .B(n9077), .ZN(
        P1_U3221) );
  AOI21_X1 U10411 ( .B1(n9081), .B2(n9080), .A(n9079), .ZN(n9089) );
  NAND2_X1 U10412 ( .A1(n9139), .A2(n9150), .ZN(n9082) );
  NAND2_X1 U10413 ( .A1(P1_U3084), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9699) );
  OAI211_X1 U10414 ( .C1(n9083), .C2(n9123), .A(n9082), .B(n9699), .ZN(n9086)
         );
  NOR2_X1 U10415 ( .A1(n9084), .A2(n9148), .ZN(n9085) );
  AOI211_X1 U10416 ( .C1(n9087), .C2(n9140), .A(n9086), .B(n9085), .ZN(n9088)
         );
  OAI21_X1 U10417 ( .B1(n9089), .B2(n9131), .A(n9088), .ZN(P1_U3226) );
  INV_X1 U10418 ( .A(n9423), .ZN(n9301) );
  OAI21_X1 U10419 ( .B1(n9092), .B2(n9091), .A(n9090), .ZN(n9093) );
  NAND2_X1 U10420 ( .A1(n9093), .A2(n9136), .ZN(n9097) );
  AOI22_X1 U10421 ( .A1(n9329), .A2(n9139), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3084), .ZN(n9094) );
  OAI21_X1 U10422 ( .B1(n9266), .B2(n9123), .A(n9094), .ZN(n9095) );
  AOI21_X1 U10423 ( .B1(n9297), .B2(n9140), .A(n9095), .ZN(n9096) );
  OAI211_X1 U10424 ( .C1(n9301), .C2(n9148), .A(n9097), .B(n9096), .ZN(
        P1_U3227) );
  INV_X1 U10425 ( .A(n9442), .ZN(n9357) );
  INV_X1 U10426 ( .A(n9098), .ZN(n9103) );
  NOR3_X1 U10427 ( .A1(n9101), .A2(n9100), .A3(n9099), .ZN(n9102) );
  OAI21_X1 U10428 ( .B1(n9103), .B2(n9102), .A(n9136), .ZN(n9108) );
  OAI22_X1 U10429 ( .A1(n9363), .A2(n9123), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9104), .ZN(n9106) );
  NOR2_X1 U10430 ( .A1(n9127), .A2(n9354), .ZN(n9105) );
  AOI211_X1 U10431 ( .C1(n9139), .C2(n9174), .A(n9106), .B(n9105), .ZN(n9107)
         );
  OAI211_X1 U10432 ( .C1(n9357), .C2(n9148), .A(n9108), .B(n9107), .ZN(
        P1_U3231) );
  NAND2_X1 U10433 ( .A1(n9109), .A2(n9110), .ZN(n9111) );
  XOR2_X1 U10434 ( .A(n9112), .B(n9111), .Z(n9119) );
  OAI22_X1 U10435 ( .A1(n9363), .A2(n9114), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9113), .ZN(n9115) );
  AOI21_X1 U10436 ( .B1(n9329), .B2(n9145), .A(n9115), .ZN(n9116) );
  OAI21_X1 U10437 ( .B1(n9127), .B2(n9322), .A(n9116), .ZN(n9117) );
  AOI21_X1 U10438 ( .B1(n9432), .B2(n9129), .A(n9117), .ZN(n9118) );
  OAI21_X1 U10439 ( .B1(n9119), .B2(n9131), .A(n9118), .ZN(P1_U3233) );
  NAND2_X1 U10440 ( .A1(n4370), .A2(n9120), .ZN(n9122) );
  XNOR2_X1 U10441 ( .A(n9122), .B(n9121), .ZN(n9132) );
  NAND2_X1 U10442 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9715) );
  OAI21_X1 U10443 ( .B1(n9123), .B2(n9362), .A(n9715), .ZN(n9124) );
  AOI21_X1 U10444 ( .B1(n9139), .B2(n9149), .A(n9124), .ZN(n9125) );
  OAI21_X1 U10445 ( .B1(n9127), .B2(n9126), .A(n9125), .ZN(n9128) );
  AOI21_X1 U10446 ( .B1(n9453), .B2(n9129), .A(n9128), .ZN(n9130) );
  OAI21_X1 U10447 ( .B1(n9132), .B2(n9131), .A(n9130), .ZN(P1_U3236) );
  AND2_X1 U10448 ( .A1(n9134), .A2(n9133), .ZN(n9138) );
  OAI211_X1 U10449 ( .C1(n9138), .C2(n9137), .A(n9136), .B(n9135), .ZN(n9147)
         );
  NAND2_X1 U10450 ( .A1(n9293), .A2(n9139), .ZN(n9142) );
  NAND2_X1 U10451 ( .A1(n9260), .A2(n9140), .ZN(n9141) );
  OAI211_X1 U10452 ( .C1(P1_STATE_REG_SCAN_IN), .C2(n9143), .A(n9142), .B(
        n9141), .ZN(n9144) );
  AOI21_X1 U10453 ( .B1(n9228), .B2(n9145), .A(n9144), .ZN(n9146) );
  OAI211_X1 U10454 ( .C1(n9262), .C2(n9148), .A(n9147), .B(n9146), .ZN(
        P1_U3238) );
  MUX2_X1 U10455 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9206), .S(n4281), .Z(
        P1_U3585) );
  MUX2_X1 U10456 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9229), .S(n4281), .Z(
        P1_U3584) );
  MUX2_X1 U10457 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9208), .S(n4281), .Z(
        P1_U3583) );
  MUX2_X1 U10458 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9228), .S(n4281), .Z(
        P1_U3582) );
  MUX2_X1 U10459 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9284), .S(n4281), .Z(
        P1_U3581) );
  MUX2_X1 U10460 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9293), .S(n4281), .Z(
        P1_U3580) );
  MUX2_X1 U10461 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9283), .S(n4281), .Z(
        P1_U3579) );
  MUX2_X1 U10462 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9329), .S(n4281), .Z(
        P1_U3578) );
  MUX2_X1 U10463 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9346), .S(n4281), .Z(
        P1_U3577) );
  MUX2_X1 U10464 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9328), .S(n4281), .Z(
        P1_U3576) );
  MUX2_X1 U10465 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9381), .S(n4281), .Z(
        P1_U3575) );
  MUX2_X1 U10466 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9174), .S(n4281), .Z(
        P1_U3574) );
  MUX2_X1 U10467 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9380), .S(n4281), .Z(
        P1_U3573) );
  MUX2_X1 U10468 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9149), .S(n4281), .Z(
        P1_U3572) );
  MUX2_X1 U10469 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9150), .S(n4281), .Z(
        P1_U3571) );
  MUX2_X1 U10470 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9151), .S(n4281), .Z(
        P1_U3570) );
  MUX2_X1 U10471 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9152), .S(n4281), .Z(
        P1_U3569) );
  MUX2_X1 U10472 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9153), .S(n4281), .Z(
        P1_U3568) );
  MUX2_X1 U10473 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9154), .S(n4281), .Z(
        P1_U3567) );
  MUX2_X1 U10474 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9559), .S(n4281), .Z(
        P1_U3566) );
  MUX2_X1 U10475 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9155), .S(n4281), .Z(
        P1_U3565) );
  MUX2_X1 U10476 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9156), .S(n4281), .Z(
        P1_U3564) );
  MUX2_X1 U10477 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9157), .S(n4281), .Z(
        P1_U3563) );
  MUX2_X1 U10478 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9735), .S(n4281), .Z(
        P1_U3562) );
  MUX2_X1 U10479 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9158), .S(n4281), .Z(
        P1_U3561) );
  MUX2_X1 U10480 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9733), .S(n4281), .Z(
        P1_U3560) );
  MUX2_X1 U10481 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9159), .S(n4281), .Z(
        P1_U3559) );
  MUX2_X1 U10482 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9160), .S(n4281), .Z(
        P1_U3558) );
  MUX2_X1 U10483 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n9161), .S(n4281), .Z(
        P1_U3557) );
  MUX2_X1 U10484 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n9162), .S(n4281), .Z(
        P1_U3556) );
  OR2_X2 U10485 ( .A1(n9373), .A2(n9447), .ZN(n9371) );
  OR2_X2 U10486 ( .A1(n9306), .A2(n9423), .ZN(n9295) );
  NOR2_X2 U10487 ( .A1(n9295), .A2(n9417), .ZN(n9276) );
  AND2_X2 U10488 ( .A1(n9262), .A2(n9276), .ZN(n9258) );
  XNOR2_X1 U10489 ( .A(n6434), .B(n9391), .ZN(n9388) );
  NAND2_X1 U10490 ( .A1(n9388), .A2(n9777), .ZN(n9167) );
  AOI21_X1 U10491 ( .B1(P1_B_REG_SCAN_IN), .B2(n9164), .A(n9781), .ZN(n9207)
         );
  NAND2_X1 U10492 ( .A1(n9207), .A2(n9165), .ZN(n9392) );
  NOR2_X1 U10493 ( .A1(n9568), .A2(n9392), .ZN(n9170) );
  AOI21_X1 U10494 ( .B1(n9383), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9170), .ZN(
        n9166) );
  OAI211_X1 U10495 ( .C1(n6434), .C2(n9791), .A(n9167), .B(n9166), .ZN(
        P1_U3261) );
  INV_X1 U10496 ( .A(n9212), .ZN(n9168) );
  NAND2_X1 U10497 ( .A1(n9169), .A2(n9168), .ZN(n9390) );
  NAND3_X1 U10498 ( .A1(n9391), .A2(n9777), .A3(n9390), .ZN(n9172) );
  AOI21_X1 U10499 ( .B1(n9568), .B2(P1_REG2_REG_30__SCAN_IN), .A(n9170), .ZN(
        n9171) );
  OAI211_X1 U10500 ( .C1(n9394), .C2(n9791), .A(n9172), .B(n9171), .ZN(
        P1_U3262) );
  NOR2_X1 U10501 ( .A1(n9447), .A2(n9174), .ZN(n9175) );
  INV_X1 U10502 ( .A(n9447), .ZN(n9377) );
  AOI21_X1 U10503 ( .B1(n9357), .B2(n9177), .A(n9176), .ZN(n9336) );
  NAND2_X1 U10504 ( .A1(n9336), .A2(n9335), .ZN(n9334) );
  NAND2_X1 U10505 ( .A1(n9334), .A2(n4840), .ZN(n9319) );
  NOR2_X1 U10506 ( .A1(n9307), .A2(n9179), .ZN(n9180) );
  OAI22_X1 U10507 ( .A1(n9275), .A2(n9281), .B1(n9293), .B2(n9417), .ZN(n9256)
         );
  NAND2_X1 U10508 ( .A1(n9256), .A2(n9264), .ZN(n9255) );
  NAND2_X1 U10509 ( .A1(n9255), .A2(n9181), .ZN(n9239) );
  INV_X1 U10510 ( .A(n9227), .ZN(n9183) );
  XNOR2_X1 U10511 ( .A(n9184), .B(n9204), .ZN(n9395) );
  INV_X1 U10512 ( .A(n9395), .ZN(n9218) );
  AOI22_X1 U10513 ( .A1(n9398), .A2(n9569), .B1(P1_REG2_REG_29__SCAN_IN), .B2(
        n9383), .ZN(n9217) );
  INV_X1 U10514 ( .A(n9187), .ZN(n9188) );
  INV_X1 U10515 ( .A(n9335), .ZN(n9344) );
  NAND3_X1 U10516 ( .A1(n9365), .A2(n9344), .A3(n9342), .ZN(n9343) );
  NAND2_X1 U10517 ( .A1(n9343), .A2(n9189), .ZN(n9327) );
  INV_X1 U10518 ( .A(n9194), .ZN(n9195) );
  OAI21_X1 U10519 ( .B1(n9282), .B2(n9196), .A(n9195), .ZN(n9263) );
  INV_X1 U10520 ( .A(n9264), .ZN(n9197) );
  NAND2_X1 U10521 ( .A1(n9263), .A2(n9197), .ZN(n9269) );
  INV_X1 U10522 ( .A(n9200), .ZN(n9201) );
  OAI21_X1 U10523 ( .B1(n9226), .B2(n9201), .A(n9203), .ZN(n9202) );
  MUX2_X1 U10524 ( .A(n9202), .B(n9201), .S(n9204), .Z(n9211) );
  NAND2_X1 U10525 ( .A1(n9205), .A2(n9786), .ZN(n9210) );
  AOI22_X1 U10526 ( .A1(n9208), .A2(n9734), .B1(n9207), .B2(n9206), .ZN(n9209)
         );
  OAI21_X1 U10527 ( .B1(n9211), .B2(n9210), .A(n9209), .ZN(n9396) );
  AOI211_X1 U10528 ( .C1(n9398), .C2(n9221), .A(n9865), .B(n9212), .ZN(n9397)
         );
  INV_X1 U10529 ( .A(n9397), .ZN(n9214) );
  OAI22_X1 U10530 ( .A1(n9214), .A2(n9757), .B1(n9792), .B2(n9213), .ZN(n9215)
         );
  OAI21_X1 U10531 ( .B1(n9396), .B2(n9215), .A(n9797), .ZN(n9216) );
  OAI211_X1 U10532 ( .C1(n9218), .C2(n9387), .A(n9217), .B(n9216), .ZN(
        P1_U3355) );
  OAI21_X1 U10533 ( .B1(n9220), .B2(n9183), .A(n9219), .ZN(n9405) );
  INV_X1 U10534 ( .A(n9221), .ZN(n9222) );
  AOI21_X1 U10535 ( .B1(n9401), .B2(n9246), .A(n9222), .ZN(n9402) );
  INV_X1 U10536 ( .A(n9223), .ZN(n9224) );
  AOI22_X1 U10537 ( .A1(n9224), .A2(n9755), .B1(P1_REG2_REG_28__SCAN_IN), .B2(
        n9383), .ZN(n9225) );
  OAI21_X1 U10538 ( .B1(n4585), .B2(n9791), .A(n9225), .ZN(n9235) );
  XOR2_X1 U10539 ( .A(n9227), .B(n9226), .Z(n9233) );
  NAND2_X1 U10540 ( .A1(n9229), .A2(n9736), .ZN(n9230) );
  AOI211_X1 U10541 ( .C1(n9777), .C2(n9402), .A(n9235), .B(n9234), .ZN(n9236)
         );
  OAI21_X1 U10542 ( .B1(n9405), .B2(n9387), .A(n9236), .ZN(P1_U3263) );
  OAI21_X1 U10543 ( .B1(n9239), .B2(n9238), .A(n9237), .ZN(n9410) );
  INV_X1 U10544 ( .A(n9410), .ZN(n9254) );
  OAI211_X1 U10545 ( .C1(n9242), .C2(n9241), .A(n9240), .B(n9786), .ZN(n9244)
         );
  NAND2_X1 U10546 ( .A1(n9284), .A2(n9734), .ZN(n9243) );
  OAI211_X1 U10547 ( .C1(n9245), .C2(n9781), .A(n9244), .B(n9243), .ZN(n9409)
         );
  OAI21_X1 U10548 ( .B1(n9406), .B2(n9258), .A(n9246), .ZN(n9407) );
  AOI22_X1 U10549 ( .A1(n9247), .A2(n9755), .B1(P1_REG2_REG_27__SCAN_IN), .B2(
        n9383), .ZN(n9250) );
  NAND2_X1 U10550 ( .A1(n9248), .A2(n9569), .ZN(n9249) );
  OAI211_X1 U10551 ( .C1(n9407), .C2(n9251), .A(n9250), .B(n9249), .ZN(n9252)
         );
  AOI21_X1 U10552 ( .B1(n9409), .B2(n9797), .A(n9252), .ZN(n9253) );
  OAI21_X1 U10553 ( .B1(n9254), .B2(n9387), .A(n9253), .ZN(P1_U3264) );
  OAI21_X1 U10554 ( .B1(n9256), .B2(n9264), .A(n9255), .ZN(n9257) );
  INV_X1 U10555 ( .A(n9257), .ZN(n9416) );
  INV_X1 U10556 ( .A(n9276), .ZN(n9259) );
  AOI21_X1 U10557 ( .B1(n9412), .B2(n9259), .A(n9258), .ZN(n9413) );
  AOI22_X1 U10558 ( .A1(n9260), .A2(n9755), .B1(P1_REG2_REG_26__SCAN_IN), .B2(
        n9383), .ZN(n9261) );
  OAI21_X1 U10559 ( .B1(n9262), .B2(n9791), .A(n9261), .ZN(n9272) );
  INV_X1 U10560 ( .A(n9263), .ZN(n9265) );
  AOI21_X1 U10561 ( .B1(n9265), .B2(n9264), .A(n9766), .ZN(n9270) );
  OAI22_X1 U10562 ( .A1(n9267), .A2(n9781), .B1(n9266), .B2(n9784), .ZN(n9268)
         );
  AOI21_X1 U10563 ( .B1(n9270), .B2(n9269), .A(n9268), .ZN(n9415) );
  NOR2_X1 U10564 ( .A1(n9415), .A2(n9568), .ZN(n9271) );
  AOI211_X1 U10565 ( .C1(n9413), .C2(n9777), .A(n9272), .B(n9271), .ZN(n9273)
         );
  OAI21_X1 U10566 ( .B1(n9416), .B2(n9387), .A(n9273), .ZN(P1_U3265) );
  XNOR2_X1 U10567 ( .A(n9275), .B(n9274), .ZN(n9421) );
  AOI21_X1 U10568 ( .B1(n9417), .B2(n9295), .A(n9276), .ZN(n9418) );
  INV_X1 U10569 ( .A(n9277), .ZN(n9278) );
  AOI22_X1 U10570 ( .A1(n9278), .A2(n9755), .B1(P1_REG2_REG_25__SCAN_IN), .B2(
        n9383), .ZN(n9279) );
  OAI21_X1 U10571 ( .B1(n9280), .B2(n9791), .A(n9279), .ZN(n9287) );
  XNOR2_X1 U10572 ( .A(n9282), .B(n9281), .ZN(n9285) );
  AOI222_X1 U10573 ( .A1(n9786), .A2(n9285), .B1(n9284), .B2(n9736), .C1(n9283), .C2(n9734), .ZN(n9420) );
  NOR2_X1 U10574 ( .A1(n9420), .A2(n9568), .ZN(n9286) );
  AOI211_X1 U10575 ( .C1(n9418), .C2(n9777), .A(n9287), .B(n9286), .ZN(n9288)
         );
  OAI21_X1 U10576 ( .B1(n9421), .B2(n9387), .A(n9288), .ZN(P1_U3266) );
  XNOR2_X1 U10577 ( .A(n9289), .B(n9291), .ZN(n9426) );
  OAI21_X1 U10578 ( .B1(n9292), .B2(n9291), .A(n9290), .ZN(n9294) );
  AOI222_X1 U10579 ( .A1(n9786), .A2(n9294), .B1(n9293), .B2(n9736), .C1(n9329), .C2(n9734), .ZN(n9425) );
  INV_X1 U10580 ( .A(n9295), .ZN(n9296) );
  AOI211_X1 U10581 ( .C1(n9423), .C2(n9306), .A(n9865), .B(n9296), .ZN(n9422)
         );
  AOI22_X1 U10582 ( .A1(n9422), .A2(n9298), .B1(n9755), .B2(n9297), .ZN(n9299)
         );
  AOI21_X1 U10583 ( .B1(n9425), .B2(n9299), .A(n9568), .ZN(n9303) );
  OAI22_X1 U10584 ( .A1(n9301), .A2(n9791), .B1(n9300), .B2(n9797), .ZN(n9302)
         );
  NOR2_X1 U10585 ( .A1(n9303), .A2(n9302), .ZN(n9304) );
  OAI21_X1 U10586 ( .B1(n9426), .B2(n9387), .A(n9304), .ZN(P1_U3267) );
  XOR2_X1 U10587 ( .A(n9305), .B(n9312), .Z(n9431) );
  AOI211_X1 U10588 ( .C1(n9429), .C2(n9320), .A(n9865), .B(n4581), .ZN(n9428)
         );
  NOR2_X1 U10589 ( .A1(n9307), .A2(n9791), .ZN(n9311) );
  OAI22_X1 U10590 ( .A1(n9797), .A2(n9309), .B1(n9308), .B2(n9792), .ZN(n9310)
         );
  AOI211_X1 U10591 ( .C1(n9428), .C2(n9350), .A(n9311), .B(n9310), .ZN(n9318)
         );
  XNOR2_X1 U10592 ( .A(n9313), .B(n9312), .ZN(n9314) );
  OAI222_X1 U10593 ( .A1(n9781), .A2(n9316), .B1(n9784), .B2(n9315), .C1(n9766), .C2(n9314), .ZN(n9427) );
  NAND2_X1 U10594 ( .A1(n9427), .A2(n9797), .ZN(n9317) );
  OAI211_X1 U10595 ( .C1(n9431), .C2(n9387), .A(n9318), .B(n9317), .ZN(
        P1_U3268) );
  XOR2_X1 U10596 ( .A(n9319), .B(n9326), .Z(n9436) );
  INV_X1 U10597 ( .A(n9337), .ZN(n9321) );
  AOI21_X1 U10598 ( .B1(n9432), .B2(n9321), .A(n4577), .ZN(n9433) );
  INV_X1 U10599 ( .A(n9322), .ZN(n9323) );
  AOI22_X1 U10600 ( .A1(n9568), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n9323), .B2(
        n9755), .ZN(n9324) );
  OAI21_X1 U10601 ( .B1(n9325), .B2(n9791), .A(n9324), .ZN(n9332) );
  XNOR2_X1 U10602 ( .A(n9327), .B(n9326), .ZN(n9330) );
  AOI222_X1 U10603 ( .A1(n9786), .A2(n9330), .B1(n9329), .B2(n9736), .C1(n9328), .C2(n9734), .ZN(n9435) );
  NOR2_X1 U10604 ( .A1(n9435), .A2(n9568), .ZN(n9331) );
  AOI211_X1 U10605 ( .C1(n9433), .C2(n9777), .A(n9332), .B(n9331), .ZN(n9333)
         );
  OAI21_X1 U10606 ( .B1(n9436), .B2(n9387), .A(n9333), .ZN(P1_U3269) );
  OAI21_X1 U10607 ( .B1(n9336), .B2(n9335), .A(n9334), .ZN(n9441) );
  INV_X1 U10608 ( .A(n9353), .ZN(n9338) );
  AOI211_X1 U10609 ( .C1(n9438), .C2(n9338), .A(n9865), .B(n9337), .ZN(n9437)
         );
  AOI22_X1 U10610 ( .A1(n9383), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n9339), .B2(
        n9755), .ZN(n9340) );
  OAI21_X1 U10611 ( .B1(n9341), .B2(n9791), .A(n9340), .ZN(n9349) );
  AND2_X1 U10612 ( .A1(n9365), .A2(n9342), .ZN(n9345) );
  OAI21_X1 U10613 ( .B1(n9345), .B2(n9344), .A(n9343), .ZN(n9347) );
  AOI222_X1 U10614 ( .A1(n9786), .A2(n9347), .B1(n9381), .B2(n9734), .C1(n9346), .C2(n9736), .ZN(n9440) );
  NOR2_X1 U10615 ( .A1(n9440), .A2(n9568), .ZN(n9348) );
  AOI211_X1 U10616 ( .C1(n9437), .C2(n9350), .A(n9349), .B(n9348), .ZN(n9351)
         );
  OAI21_X1 U10617 ( .B1(n9441), .B2(n9387), .A(n9351), .ZN(P1_U3270) );
  XOR2_X1 U10618 ( .A(n9359), .B(n9352), .Z(n9446) );
  AOI21_X1 U10619 ( .B1(n9442), .B2(n9371), .A(n9353), .ZN(n9443) );
  INV_X1 U10620 ( .A(n9354), .ZN(n9355) );
  AOI22_X1 U10621 ( .A1(n9568), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9355), .B2(
        n9755), .ZN(n9356) );
  OAI21_X1 U10622 ( .B1(n9357), .B2(n9791), .A(n9356), .ZN(n9368) );
  INV_X1 U10623 ( .A(n9358), .ZN(n9361) );
  INV_X1 U10624 ( .A(n9359), .ZN(n9360) );
  AOI21_X1 U10625 ( .B1(n9361), .B2(n9360), .A(n9766), .ZN(n9366) );
  OAI22_X1 U10626 ( .A1(n9363), .A2(n9781), .B1(n9362), .B2(n9784), .ZN(n9364)
         );
  AOI21_X1 U10627 ( .B1(n9366), .B2(n9365), .A(n9364), .ZN(n9445) );
  NOR2_X1 U10628 ( .A1(n9445), .A2(n9568), .ZN(n9367) );
  AOI211_X1 U10629 ( .C1(n9443), .C2(n9777), .A(n9368), .B(n9367), .ZN(n9369)
         );
  OAI21_X1 U10630 ( .B1(n9446), .B2(n9387), .A(n9369), .ZN(P1_U3271) );
  XNOR2_X1 U10631 ( .A(n9370), .B(n9378), .ZN(n9451) );
  INV_X1 U10632 ( .A(n9371), .ZN(n9372) );
  AOI21_X1 U10633 ( .B1(n9447), .B2(n9373), .A(n9372), .ZN(n9448) );
  INV_X1 U10634 ( .A(n9374), .ZN(n9375) );
  AOI22_X1 U10635 ( .A1(n9568), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9375), .B2(
        n9755), .ZN(n9376) );
  OAI21_X1 U10636 ( .B1(n9377), .B2(n9791), .A(n9376), .ZN(n9385) );
  XNOR2_X1 U10637 ( .A(n9379), .B(n9378), .ZN(n9382) );
  AOI222_X1 U10638 ( .A1(n9786), .A2(n9382), .B1(n9381), .B2(n9736), .C1(n9380), .C2(n9734), .ZN(n9450) );
  NOR2_X1 U10639 ( .A1(n9450), .A2(n9383), .ZN(n9384) );
  AOI211_X1 U10640 ( .C1(n9448), .C2(n9777), .A(n9385), .B(n9384), .ZN(n9386)
         );
  OAI21_X1 U10641 ( .B1(n9451), .B2(n9387), .A(n9386), .ZN(P1_U3272) );
  NAND2_X1 U10642 ( .A1(n9388), .A2(n9857), .ZN(n9389) );
  OAI211_X1 U10643 ( .C1(n6434), .C2(n9863), .A(n9389), .B(n9392), .ZN(n9474)
         );
  MUX2_X1 U10644 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9474), .S(n9887), .Z(
        P1_U3554) );
  NAND3_X1 U10645 ( .A1(n9391), .A2(n9857), .A3(n9390), .ZN(n9393) );
  OAI211_X1 U10646 ( .C1(n9394), .C2(n9863), .A(n9393), .B(n9392), .ZN(n9475)
         );
  MUX2_X1 U10647 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n9475), .S(n9887), .Z(
        P1_U3553) );
  NAND2_X1 U10648 ( .A1(n9395), .A2(n9853), .ZN(n9400) );
  AOI211_X2 U10649 ( .C1(n9856), .C2(n9398), .A(n9397), .B(n9396), .ZN(n9399)
         );
  NAND2_X1 U10650 ( .A1(n9400), .A2(n9399), .ZN(n9476) );
  MUX2_X1 U10651 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9476), .S(n9887), .Z(
        P1_U3552) );
  AOI22_X1 U10652 ( .A1(n9402), .A2(n9857), .B1(n9856), .B2(n9401), .ZN(n9403)
         );
  OAI211_X1 U10653 ( .C1(n9405), .C2(n9472), .A(n9404), .B(n9403), .ZN(n9477)
         );
  MUX2_X1 U10654 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9477), .S(n9887), .Z(
        P1_U3551) );
  OAI22_X1 U10655 ( .A1(n9407), .A2(n9865), .B1(n9406), .B2(n9863), .ZN(n9408)
         );
  AOI211_X1 U10656 ( .C1(n9410), .C2(n9853), .A(n9409), .B(n9408), .ZN(n9411)
         );
  INV_X1 U10657 ( .A(n9411), .ZN(n9478) );
  MUX2_X1 U10658 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9478), .S(n9887), .Z(
        P1_U3550) );
  AOI22_X1 U10659 ( .A1(n9413), .A2(n9857), .B1(n9856), .B2(n9412), .ZN(n9414)
         );
  OAI211_X1 U10660 ( .C1(n9416), .C2(n9472), .A(n9415), .B(n9414), .ZN(n9479)
         );
  MUX2_X1 U10661 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9479), .S(n9887), .Z(
        P1_U3549) );
  AOI22_X1 U10662 ( .A1(n9418), .A2(n9857), .B1(n9856), .B2(n9417), .ZN(n9419)
         );
  OAI211_X1 U10663 ( .C1(n9421), .C2(n9472), .A(n9420), .B(n9419), .ZN(n9480)
         );
  MUX2_X1 U10664 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9480), .S(n9887), .Z(
        P1_U3548) );
  AOI21_X1 U10665 ( .B1(n9856), .B2(n9423), .A(n9422), .ZN(n9424) );
  OAI211_X1 U10666 ( .C1(n9426), .C2(n9472), .A(n9425), .B(n9424), .ZN(n9481)
         );
  MUX2_X1 U10667 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9481), .S(n9887), .Z(
        P1_U3547) );
  AOI211_X1 U10668 ( .C1(n9856), .C2(n9429), .A(n9428), .B(n9427), .ZN(n9430)
         );
  OAI21_X1 U10669 ( .B1(n9431), .B2(n9472), .A(n9430), .ZN(n9482) );
  MUX2_X1 U10670 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9482), .S(n9887), .Z(
        P1_U3546) );
  AOI22_X1 U10671 ( .A1(n9433), .A2(n9857), .B1(n9856), .B2(n9432), .ZN(n9434)
         );
  OAI211_X1 U10672 ( .C1(n9436), .C2(n9472), .A(n9435), .B(n9434), .ZN(n9483)
         );
  MUX2_X1 U10673 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9483), .S(n9887), .Z(
        P1_U3545) );
  AOI21_X1 U10674 ( .B1(n9856), .B2(n9438), .A(n9437), .ZN(n9439) );
  OAI211_X1 U10675 ( .C1(n9441), .C2(n9472), .A(n9440), .B(n9439), .ZN(n9484)
         );
  MUX2_X1 U10676 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9484), .S(n9887), .Z(
        P1_U3544) );
  AOI22_X1 U10677 ( .A1(n9443), .A2(n9857), .B1(n9856), .B2(n9442), .ZN(n9444)
         );
  OAI211_X1 U10678 ( .C1(n9446), .C2(n9472), .A(n9445), .B(n9444), .ZN(n9485)
         );
  MUX2_X1 U10679 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9485), .S(n9887), .Z(
        P1_U3543) );
  AOI22_X1 U10680 ( .A1(n9448), .A2(n9857), .B1(n9856), .B2(n9447), .ZN(n9449)
         );
  OAI211_X1 U10681 ( .C1(n9451), .C2(n9472), .A(n9450), .B(n9449), .ZN(n9486)
         );
  MUX2_X1 U10682 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9486), .S(n9887), .Z(
        P1_U3542) );
  INV_X1 U10683 ( .A(n9452), .ZN(n9457) );
  AOI22_X1 U10684 ( .A1(n9454), .A2(n9857), .B1(n9856), .B2(n9453), .ZN(n9455)
         );
  OAI211_X1 U10685 ( .C1(n9457), .C2(n9472), .A(n9456), .B(n9455), .ZN(n9487)
         );
  MUX2_X1 U10686 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9487), .S(n9887), .Z(
        P1_U3541) );
  AOI22_X1 U10687 ( .A1(n9459), .A2(n9857), .B1(n9856), .B2(n9458), .ZN(n9460)
         );
  OAI211_X1 U10688 ( .C1(n9462), .C2(n9472), .A(n9461), .B(n9460), .ZN(n9488)
         );
  MUX2_X1 U10689 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9488), .S(n9887), .Z(
        P1_U3540) );
  AOI211_X1 U10690 ( .C1(n9856), .C2(n9465), .A(n9464), .B(n9463), .ZN(n9466)
         );
  OAI21_X1 U10691 ( .B1(n9467), .B2(n9472), .A(n9466), .ZN(n9489) );
  MUX2_X1 U10692 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9489), .S(n9887), .Z(
        P1_U3539) );
  AOI211_X1 U10693 ( .C1(n9856), .C2(n9470), .A(n9469), .B(n9468), .ZN(n9471)
         );
  OAI21_X1 U10694 ( .B1(n9473), .B2(n9472), .A(n9471), .ZN(n9490) );
  MUX2_X1 U10695 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n9490), .S(n9887), .Z(
        P1_U3534) );
  MUX2_X1 U10696 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9474), .S(n9872), .Z(
        P1_U3522) );
  MUX2_X1 U10697 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n9475), .S(n9872), .Z(
        P1_U3521) );
  MUX2_X1 U10698 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9476), .S(n9872), .Z(
        P1_U3520) );
  MUX2_X1 U10699 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9477), .S(n9872), .Z(
        P1_U3519) );
  MUX2_X1 U10700 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9478), .S(n9872), .Z(
        P1_U3518) );
  MUX2_X1 U10701 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9479), .S(n9872), .Z(
        P1_U3517) );
  MUX2_X1 U10702 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9480), .S(n9872), .Z(
        P1_U3516) );
  MUX2_X1 U10703 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9481), .S(n9872), .Z(
        P1_U3515) );
  MUX2_X1 U10704 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9482), .S(n9872), .Z(
        P1_U3514) );
  MUX2_X1 U10705 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9483), .S(n9872), .Z(
        P1_U3513) );
  MUX2_X1 U10706 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9484), .S(n9872), .Z(
        P1_U3512) );
  MUX2_X1 U10707 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9485), .S(n9872), .Z(
        P1_U3511) );
  MUX2_X1 U10708 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9486), .S(n9872), .Z(
        P1_U3510) );
  MUX2_X1 U10709 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9487), .S(n9872), .Z(
        P1_U3508) );
  MUX2_X1 U10710 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9488), .S(n9872), .Z(
        P1_U3505) );
  MUX2_X1 U10711 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9489), .S(n9872), .Z(
        P1_U3502) );
  MUX2_X1 U10712 ( .A(P1_REG0_REG_11__SCAN_IN), .B(n9490), .S(n9872), .Z(
        P1_U3487) );
  MUX2_X1 U10713 ( .A(n9491), .B(P1_D_REG_0__SCAN_IN), .S(n9809), .Z(P1_U3440)
         );
  INV_X1 U10714 ( .A(n9039), .ZN(n9498) );
  INV_X1 U10715 ( .A(n9492), .ZN(n9494) );
  NOR4_X1 U10716 ( .A1(n9494), .A2(P1_IR_REG_30__SCAN_IN), .A3(n9493), .A4(
        P1_U3084), .ZN(n9495) );
  AOI21_X1 U10717 ( .B1(n9496), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9495), .ZN(
        n9497) );
  OAI21_X1 U10718 ( .B1(n9498), .B2(n4282), .A(n9497), .ZN(P1_U3322) );
  OAI222_X1 U10719 ( .A1(n9502), .A2(n9501), .B1(n4282), .B2(n9500), .C1(n9499), .C2(P1_U3084), .ZN(P1_U3324) );
  INV_X1 U10720 ( .A(n9503), .ZN(n9504) );
  AOI21_X1 U10721 ( .B1(n9892), .B2(P2_ADDR_REG_1__SCAN_IN), .A(n9504), .ZN(
        n9516) );
  AOI211_X1 U10722 ( .C1(n9507), .C2(n9506), .A(n9505), .B(n9895), .ZN(n9508)
         );
  AOI21_X1 U10723 ( .B1(n9522), .B2(n9509), .A(n9508), .ZN(n9515) );
  INV_X1 U10724 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n9510) );
  NOR2_X1 U10725 ( .A1(n9510), .A2(n10029), .ZN(n9513) );
  OAI211_X1 U10726 ( .C1(n9513), .C2(n9512), .A(n9888), .B(n9511), .ZN(n9514)
         );
  NAND3_X1 U10727 ( .A1(n9516), .A2(n9515), .A3(n9514), .ZN(P2_U3246) );
  AOI21_X1 U10728 ( .B1(n9892), .B2(P2_ADDR_REG_2__SCAN_IN), .A(n9517), .ZN(
        n9528) );
  AOI211_X1 U10729 ( .C1(n4321), .C2(n9519), .A(n9518), .B(n9895), .ZN(n9520)
         );
  AOI21_X1 U10730 ( .B1(n9522), .B2(n9521), .A(n9520), .ZN(n9527) );
  OAI211_X1 U10731 ( .C1(n9525), .C2(n9524), .A(n9888), .B(n9523), .ZN(n9526)
         );
  NAND3_X1 U10732 ( .A1(n9528), .A2(n9527), .A3(n9526), .ZN(P2_U3247) );
  OAI22_X1 U10733 ( .A1(n9530), .A2(n10004), .B1(n9529), .B2(n10019), .ZN(
        n9532) );
  AOI211_X1 U10734 ( .C1(n10025), .C2(n9533), .A(n9532), .B(n9531), .ZN(n9549)
         );
  INV_X1 U10735 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n9534) );
  AOI22_X1 U10736 ( .A1(n10045), .A2(n9549), .B1(n9534), .B2(n10042), .ZN(
        P2_U3535) );
  OAI211_X1 U10737 ( .C1(n9537), .C2(n10019), .A(n9536), .B(n9535), .ZN(n9538)
         );
  AOI21_X1 U10738 ( .B1(n10025), .B2(n9539), .A(n9538), .ZN(n9551) );
  AOI22_X1 U10739 ( .A1(n10045), .A2(n9551), .B1(n9540), .B2(n10042), .ZN(
        P2_U3534) );
  INV_X1 U10740 ( .A(n9541), .ZN(n9999) );
  INV_X1 U10741 ( .A(n9542), .ZN(n9546) );
  OAI22_X1 U10742 ( .A1(n9543), .A2(n10004), .B1(n8003), .B2(n10019), .ZN(
        n9545) );
  AOI211_X1 U10743 ( .C1(n9999), .C2(n9546), .A(n9545), .B(n9544), .ZN(n9553)
         );
  AOI22_X1 U10744 ( .A1(n10045), .A2(n9553), .B1(n9547), .B2(n10042), .ZN(
        P2_U3533) );
  INV_X1 U10745 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n9548) );
  AOI22_X1 U10746 ( .A1(n10028), .A2(n9549), .B1(n9548), .B2(n10026), .ZN(
        P2_U3496) );
  AOI22_X1 U10747 ( .A1(n10028), .A2(n9551), .B1(n9550), .B2(n10026), .ZN(
        P2_U3493) );
  INV_X1 U10748 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n9552) );
  AOI22_X1 U10749 ( .A1(n10028), .A2(n9553), .B1(n9552), .B2(n10026), .ZN(
        P2_U3490) );
  OAI21_X1 U10750 ( .B1(n9555), .B2(n9557), .A(n9554), .ZN(n9556) );
  INV_X1 U10751 ( .A(n9556), .ZN(n9603) );
  XNOR2_X1 U10752 ( .A(n9558), .B(n9557), .ZN(n9563) );
  NAND2_X1 U10753 ( .A1(n9734), .A2(n9559), .ZN(n9560) );
  OAI21_X1 U10754 ( .B1(n9561), .B2(n9781), .A(n9560), .ZN(n9562) );
  AOI21_X1 U10755 ( .B1(n9563), .B2(n9786), .A(n9562), .ZN(n9600) );
  INV_X1 U10756 ( .A(n9600), .ZN(n9564) );
  AOI21_X1 U10757 ( .B1(n9603), .B2(n9565), .A(n9564), .ZN(n9578) );
  INV_X1 U10758 ( .A(n9566), .ZN(n9567) );
  AOI222_X1 U10759 ( .A1(n9571), .A2(n9569), .B1(P1_REG2_REG_12__SCAN_IN), 
        .B2(n9568), .C1(n9755), .C2(n9567), .ZN(n9577) );
  INV_X1 U10760 ( .A(n9570), .ZN(n9573) );
  INV_X1 U10761 ( .A(n9571), .ZN(n9601) );
  OAI211_X1 U10762 ( .C1(n9573), .C2(n9601), .A(n9857), .B(n9572), .ZN(n9599)
         );
  INV_X1 U10763 ( .A(n9599), .ZN(n9574) );
  AOI22_X1 U10764 ( .A1(n9603), .A2(n9778), .B1(n9575), .B2(n9574), .ZN(n9576)
         );
  OAI211_X1 U10765 ( .C1(n9383), .C2(n9578), .A(n9577), .B(n9576), .ZN(
        P1_U3279) );
  INV_X1 U10766 ( .A(n9579), .ZN(n9583) );
  OAI22_X1 U10767 ( .A1(n9581), .A2(n9865), .B1(n9580), .B2(n9863), .ZN(n9582)
         );
  AOI211_X1 U10768 ( .C1(n9584), .C2(n9853), .A(n9583), .B(n9582), .ZN(n9605)
         );
  INV_X1 U10769 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9585) );
  AOI22_X1 U10770 ( .A1(n9887), .A2(n9605), .B1(n9585), .B2(n9885), .ZN(
        P1_U3538) );
  OAI211_X1 U10771 ( .C1(n9588), .C2(n9863), .A(n9587), .B(n9586), .ZN(n9589)
         );
  AOI21_X1 U10772 ( .B1(n9853), .B2(n9590), .A(n9589), .ZN(n9607) );
  AOI22_X1 U10773 ( .A1(n9887), .A2(n9607), .B1(n9591), .B2(n9885), .ZN(
        P1_U3537) );
  INV_X1 U10774 ( .A(n9818), .ZN(n9870) );
  OAI22_X1 U10775 ( .A1(n9593), .A2(n9865), .B1(n9592), .B2(n9863), .ZN(n9594)
         );
  AOI21_X1 U10776 ( .B1(n9595), .B2(n9870), .A(n9594), .ZN(n9596) );
  AND2_X1 U10777 ( .A1(n9597), .A2(n9596), .ZN(n9609) );
  AOI22_X1 U10778 ( .A1(n9887), .A2(n9609), .B1(n9598), .B2(n9885), .ZN(
        P1_U3536) );
  OAI211_X1 U10779 ( .C1(n9601), .C2(n9863), .A(n9600), .B(n9599), .ZN(n9602)
         );
  AOI21_X1 U10780 ( .B1(n9603), .B2(n9853), .A(n9602), .ZN(n9611) );
  AOI22_X1 U10781 ( .A1(n9887), .A2(n9611), .B1(n5328), .B2(n9885), .ZN(
        P1_U3535) );
  INV_X1 U10782 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n9604) );
  AOI22_X1 U10783 ( .A1(n9872), .A2(n9605), .B1(n9604), .B2(n9871), .ZN(
        P1_U3499) );
  INV_X1 U10784 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n9606) );
  AOI22_X1 U10785 ( .A1(n9872), .A2(n9607), .B1(n9606), .B2(n9871), .ZN(
        P1_U3496) );
  INV_X1 U10786 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n9608) );
  AOI22_X1 U10787 ( .A1(n9872), .A2(n9609), .B1(n9608), .B2(n9871), .ZN(
        P1_U3493) );
  INV_X1 U10788 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n9610) );
  AOI22_X1 U10789 ( .A1(n9872), .A2(n9611), .B1(n9610), .B2(n9871), .ZN(
        P1_U3490) );
  XNOR2_X1 U10790 ( .A(P1_WR_REG_SCAN_IN), .B(P2_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U10791 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  INV_X1 U10792 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n9617) );
  OAI21_X1 U10793 ( .B1(P1_IR_REG_0__SCAN_IN), .B2(n5098), .A(n9612), .ZN(
        n9613) );
  NAND2_X1 U10794 ( .A1(n9614), .A2(n9613), .ZN(n9615) );
  OAI22_X1 U10795 ( .A1(n9727), .A2(n9617), .B1(n9616), .B2(n9615), .ZN(n9618)
         );
  INV_X1 U10796 ( .A(n9618), .ZN(n9620) );
  NAND3_X1 U10797 ( .A1(n9704), .A2(P1_IR_REG_0__SCAN_IN), .A3(n5098), .ZN(
        n9619) );
  OAI211_X1 U10798 ( .C1(P1_STATE_REG_SCAN_IN), .C2(n7178), .A(n9620), .B(
        n9619), .ZN(P1_U3241) );
  OAI21_X1 U10799 ( .B1(n9623), .B2(n9622), .A(n9621), .ZN(n9633) );
  INV_X1 U10800 ( .A(n9624), .ZN(n9632) );
  INV_X1 U10801 ( .A(n9625), .ZN(n9630) );
  AOI21_X1 U10802 ( .B1(n9628), .B2(n9627), .A(n9626), .ZN(n9629) );
  OAI21_X1 U10803 ( .B1(n9630), .B2(n9629), .A(n9704), .ZN(n9631) );
  OAI211_X1 U10804 ( .C1(n9681), .C2(n9633), .A(n9632), .B(n9631), .ZN(n9634)
         );
  INV_X1 U10805 ( .A(n9634), .ZN(n9638) );
  OAI22_X1 U10806 ( .A1(n9727), .A2(n7403), .B1(n9635), .B2(n9717), .ZN(n9636)
         );
  INV_X1 U10807 ( .A(n9636), .ZN(n9637) );
  NAND2_X1 U10808 ( .A1(n9638), .A2(n9637), .ZN(P1_U3247) );
  INV_X1 U10809 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n9652) );
  NOR2_X1 U10810 ( .A1(n9640), .A2(n9639), .ZN(n9641) );
  NOR3_X1 U10811 ( .A1(n9681), .A2(n9642), .A3(n9641), .ZN(n9643) );
  AOI211_X1 U10812 ( .C1(n9688), .C2(n9645), .A(n9644), .B(n9643), .ZN(n9651)
         );
  AOI21_X1 U10813 ( .B1(n9648), .B2(n9647), .A(n9646), .ZN(n9649) );
  OR2_X1 U10814 ( .A1(n9724), .A2(n9649), .ZN(n9650) );
  OAI211_X1 U10815 ( .C1(n9652), .C2(n9727), .A(n9651), .B(n9650), .ZN(
        P1_U3254) );
  AOI21_X1 U10816 ( .B1(n9655), .B2(n9654), .A(n9653), .ZN(n9656) );
  NAND2_X1 U10817 ( .A1(n9714), .A2(n9656), .ZN(n9659) );
  INV_X1 U10818 ( .A(n9657), .ZN(n9658) );
  OAI211_X1 U10819 ( .C1(n9717), .C2(n9660), .A(n9659), .B(n9658), .ZN(n9661)
         );
  INV_X1 U10820 ( .A(n9661), .ZN(n9667) );
  AOI21_X1 U10821 ( .B1(n9664), .B2(n9663), .A(n9662), .ZN(n9665) );
  OR2_X1 U10822 ( .A1(n9724), .A2(n9665), .ZN(n9666) );
  OAI211_X1 U10823 ( .C1(n9668), .C2(n9727), .A(n9667), .B(n9666), .ZN(
        P1_U3255) );
  INV_X1 U10824 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n9679) );
  INV_X1 U10825 ( .A(n9669), .ZN(n9673) );
  AOI211_X1 U10826 ( .C1(n7843), .C2(n9671), .A(n9681), .B(n9670), .ZN(n9672)
         );
  AOI211_X1 U10827 ( .C1(n9688), .C2(n9674), .A(n9673), .B(n9672), .ZN(n9678)
         );
  XOR2_X1 U10828 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9675), .Z(n9676) );
  NAND2_X1 U10829 ( .A1(n9704), .A2(n9676), .ZN(n9677) );
  OAI211_X1 U10830 ( .C1(n9679), .C2(n9727), .A(n9678), .B(n9677), .ZN(
        P1_U3256) );
  INV_X1 U10831 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n9694) );
  INV_X1 U10832 ( .A(n9680), .ZN(n9686) );
  AOI211_X1 U10833 ( .C1(n9684), .C2(n9683), .A(n9682), .B(n9681), .ZN(n9685)
         );
  AOI211_X1 U10834 ( .C1(n9688), .C2(n9687), .A(n9686), .B(n9685), .ZN(n9693)
         );
  OAI211_X1 U10835 ( .C1(n9691), .C2(n9690), .A(n9704), .B(n9689), .ZN(n9692)
         );
  OAI211_X1 U10836 ( .C1(n9694), .C2(n9727), .A(n9693), .B(n9692), .ZN(
        P1_U3257) );
  AOI21_X1 U10837 ( .B1(n9697), .B2(n9696), .A(n9695), .ZN(n9698) );
  NAND2_X1 U10838 ( .A1(n9714), .A2(n9698), .ZN(n9700) );
  OAI211_X1 U10839 ( .C1(n9717), .C2(n9701), .A(n9700), .B(n9699), .ZN(n9702)
         );
  INV_X1 U10840 ( .A(n9702), .ZN(n9708) );
  OAI211_X1 U10841 ( .C1(n9706), .C2(n9705), .A(n9704), .B(n9703), .ZN(n9707)
         );
  OAI211_X1 U10842 ( .C1(n9709), .C2(n9727), .A(n9708), .B(n9707), .ZN(
        P1_U3258) );
  INV_X1 U10843 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n9728) );
  AOI21_X1 U10844 ( .B1(n9712), .B2(n9711), .A(n9710), .ZN(n9713) );
  NAND2_X1 U10845 ( .A1(n9714), .A2(n9713), .ZN(n9716) );
  OAI211_X1 U10846 ( .C1(n9718), .C2(n9717), .A(n9716), .B(n9715), .ZN(n9719)
         );
  INV_X1 U10847 ( .A(n9719), .ZN(n9726) );
  AOI21_X1 U10848 ( .B1(n9722), .B2(n9721), .A(n9720), .ZN(n9723) );
  OR2_X1 U10849 ( .A1(n9724), .A2(n9723), .ZN(n9725) );
  OAI211_X1 U10850 ( .C1(n9728), .C2(n9727), .A(n9726), .B(n9725), .ZN(
        P1_U3259) );
  AOI21_X1 U10851 ( .B1(n9738), .B2(n9729), .A(n7155), .ZN(n9742) );
  INV_X1 U10852 ( .A(n9742), .ZN(n9845) );
  OAI21_X1 U10853 ( .B1(n9750), .B2(n9841), .A(n9731), .ZN(n9842) );
  INV_X1 U10854 ( .A(n9842), .ZN(n9732) );
  AOI22_X1 U10855 ( .A1(n9845), .A2(n9778), .B1(n9777), .B2(n9732), .ZN(n9748)
         );
  AOI22_X1 U10856 ( .A1(n9736), .A2(n9735), .B1(n9734), .B2(n9733), .ZN(n9741)
         );
  XOR2_X1 U10857 ( .A(n9738), .B(n9737), .Z(n9739) );
  NAND2_X1 U10858 ( .A1(n9739), .A2(n9786), .ZN(n9740) );
  OAI211_X1 U10859 ( .C1(n9742), .C2(n9789), .A(n9741), .B(n9740), .ZN(n9843)
         );
  NOR2_X1 U10860 ( .A1(n9791), .A2(n9841), .ZN(n9746) );
  OAI22_X1 U10861 ( .A1(n9797), .A2(n9744), .B1(n9743), .B2(n9792), .ZN(n9745)
         );
  AOI211_X1 U10862 ( .C1(n9843), .C2(n9797), .A(n9746), .B(n9745), .ZN(n9747)
         );
  NAND2_X1 U10863 ( .A1(n9748), .A2(n9747), .ZN(P1_U3285) );
  XOR2_X1 U10864 ( .A(n9749), .B(n9760), .Z(n9839) );
  OAI21_X1 U10865 ( .B1(n9773), .B2(n9836), .A(n9857), .ZN(n9751) );
  OR2_X1 U10866 ( .A1(n9751), .A2(n9750), .ZN(n9835) );
  AOI22_X1 U10867 ( .A1(n9755), .A2(n9754), .B1(n9753), .B2(n9752), .ZN(n9756)
         );
  OAI21_X1 U10868 ( .B1(n9835), .B2(n9757), .A(n9756), .ZN(n9768) );
  INV_X1 U10869 ( .A(n9760), .ZN(n9759) );
  NOR2_X1 U10870 ( .A1(n9759), .A2(n9758), .ZN(n9764) );
  AOI21_X1 U10871 ( .B1(n9763), .B2(n9761), .A(n9760), .ZN(n9762) );
  AOI21_X1 U10872 ( .B1(n9764), .B2(n9763), .A(n9762), .ZN(n9765) );
  OAI222_X1 U10873 ( .A1(n9781), .A2(n5181), .B1(n9784), .B2(n9767), .C1(n9766), .C2(n9765), .ZN(n9837) );
  AOI211_X1 U10874 ( .C1(n9769), .C2(n9839), .A(n9768), .B(n9837), .ZN(n9770)
         );
  AOI22_X1 U10875 ( .A1(n9383), .A2(n6588), .B1(n9770), .B2(n9797), .ZN(
        P1_U3286) );
  XOR2_X1 U10876 ( .A(n9771), .B(n9780), .Z(n9790) );
  INV_X1 U10877 ( .A(n9790), .ZN(n9833) );
  INV_X1 U10878 ( .A(n9772), .ZN(n9775) );
  INV_X1 U10879 ( .A(n9773), .ZN(n9774) );
  OAI21_X1 U10880 ( .B1(n9829), .B2(n9775), .A(n9774), .ZN(n9830) );
  INV_X1 U10881 ( .A(n9830), .ZN(n9776) );
  AOI22_X1 U10882 ( .A1(n9833), .A2(n9778), .B1(n9777), .B2(n9776), .ZN(n9799)
         );
  XOR2_X1 U10883 ( .A(n9780), .B(n9779), .Z(n9787) );
  OAI22_X1 U10884 ( .A1(n9784), .A2(n9783), .B1(n9782), .B2(n9781), .ZN(n9785)
         );
  AOI21_X1 U10885 ( .B1(n9787), .B2(n9786), .A(n9785), .ZN(n9788) );
  OAI21_X1 U10886 ( .B1(n9790), .B2(n9789), .A(n9788), .ZN(n9831) );
  NOR2_X1 U10887 ( .A1(n9791), .A2(n9829), .ZN(n9796) );
  OAI22_X1 U10888 ( .A1(n9797), .A2(n9794), .B1(n9793), .B2(n9792), .ZN(n9795)
         );
  AOI211_X1 U10889 ( .C1(n9831), .C2(n9797), .A(n9796), .B(n9795), .ZN(n9798)
         );
  NAND2_X1 U10890 ( .A1(n9799), .A2(n9798), .ZN(P1_U3287) );
  NOR2_X1 U10891 ( .A1(n9808), .A2(n9800), .ZN(P1_U3292) );
  NOR2_X1 U10892 ( .A1(n9808), .A2(n9801), .ZN(P1_U3293) );
  AND2_X1 U10893 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9809), .ZN(P1_U3294) );
  AND2_X1 U10894 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9809), .ZN(P1_U3295) );
  AND2_X1 U10895 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9809), .ZN(P1_U3296) );
  AND2_X1 U10896 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9809), .ZN(P1_U3297) );
  AND2_X1 U10897 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9809), .ZN(P1_U3298) );
  AND2_X1 U10898 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9809), .ZN(P1_U3299) );
  NOR2_X1 U10899 ( .A1(n9808), .A2(n9802), .ZN(P1_U3300) );
  AND2_X1 U10900 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9809), .ZN(P1_U3301) );
  AND2_X1 U10901 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9809), .ZN(P1_U3302) );
  AND2_X1 U10902 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9809), .ZN(P1_U3303) );
  AND2_X1 U10903 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9809), .ZN(P1_U3304) );
  AND2_X1 U10904 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9809), .ZN(P1_U3305) );
  NOR2_X1 U10905 ( .A1(n9808), .A2(n9803), .ZN(P1_U3306) );
  AND2_X1 U10906 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9809), .ZN(P1_U3307) );
  AND2_X1 U10907 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9809), .ZN(P1_U3308) );
  AND2_X1 U10908 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9809), .ZN(P1_U3309) );
  AND2_X1 U10909 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9809), .ZN(P1_U3310) );
  AND2_X1 U10910 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9809), .ZN(P1_U3311) );
  AND2_X1 U10911 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9809), .ZN(P1_U3312) );
  AND2_X1 U10912 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9809), .ZN(P1_U3313) );
  NOR2_X1 U10913 ( .A1(n9808), .A2(n9804), .ZN(P1_U3314) );
  NOR2_X1 U10914 ( .A1(n9808), .A2(n9805), .ZN(P1_U3315) );
  AND2_X1 U10915 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9809), .ZN(P1_U3316) );
  NOR2_X1 U10916 ( .A1(n9808), .A2(n9806), .ZN(P1_U3317) );
  AND2_X1 U10917 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9809), .ZN(P1_U3318) );
  NOR2_X1 U10918 ( .A1(n9808), .A2(n9807), .ZN(P1_U3319) );
  AND2_X1 U10919 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9809), .ZN(P1_U3320) );
  AND2_X1 U10920 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9809), .ZN(P1_U3321) );
  INV_X1 U10921 ( .A(n9810), .ZN(n9814) );
  OAI21_X1 U10922 ( .B1(n4568), .B2(n9863), .A(n9811), .ZN(n9813) );
  AOI211_X1 U10923 ( .C1(n9870), .C2(n9814), .A(n9813), .B(n9812), .ZN(n9874)
         );
  AOI22_X1 U10924 ( .A1(n9872), .A2(n9874), .B1(n5112), .B2(n9871), .ZN(
        P1_U3457) );
  AOI22_X1 U10925 ( .A1(n9816), .A2(n9857), .B1(n9856), .B2(n9815), .ZN(n9817)
         );
  OAI21_X1 U10926 ( .B1(n9819), .B2(n9818), .A(n9817), .ZN(n9821) );
  NOR2_X1 U10927 ( .A1(n9821), .A2(n9820), .ZN(n9876) );
  INV_X1 U10928 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9822) );
  AOI22_X1 U10929 ( .A1(n9872), .A2(n9876), .B1(n9822), .B2(n9871), .ZN(
        P1_U3460) );
  OAI22_X1 U10930 ( .A1(n9824), .A2(n9865), .B1(n9823), .B2(n9863), .ZN(n9826)
         );
  AOI211_X1 U10931 ( .C1(n9870), .C2(n9827), .A(n9826), .B(n9825), .ZN(n9877)
         );
  AOI22_X1 U10932 ( .A1(n9872), .A2(n9877), .B1(n9828), .B2(n9871), .ZN(
        P1_U3463) );
  OAI22_X1 U10933 ( .A1(n9830), .A2(n9865), .B1(n9829), .B2(n9863), .ZN(n9832)
         );
  AOI211_X1 U10934 ( .C1(n9870), .C2(n9833), .A(n9832), .B(n9831), .ZN(n9878)
         );
  INV_X1 U10935 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n9834) );
  AOI22_X1 U10936 ( .A1(n9872), .A2(n9878), .B1(n9834), .B2(n9871), .ZN(
        P1_U3466) );
  OAI21_X1 U10937 ( .B1(n9836), .B2(n9863), .A(n9835), .ZN(n9838) );
  AOI211_X1 U10938 ( .C1(n9853), .C2(n9839), .A(n9838), .B(n9837), .ZN(n9880)
         );
  INV_X1 U10939 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n9840) );
  AOI22_X1 U10940 ( .A1(n9872), .A2(n9880), .B1(n9840), .B2(n9871), .ZN(
        P1_U3469) );
  OAI22_X1 U10941 ( .A1(n9842), .A2(n9865), .B1(n9841), .B2(n9863), .ZN(n9844)
         );
  AOI211_X1 U10942 ( .C1(n9870), .C2(n9845), .A(n9844), .B(n9843), .ZN(n9881)
         );
  INV_X1 U10943 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9846) );
  AOI22_X1 U10944 ( .A1(n9872), .A2(n9881), .B1(n9846), .B2(n9871), .ZN(
        P1_U3472) );
  OAI211_X1 U10945 ( .C1(n9849), .C2(n9863), .A(n9848), .B(n9847), .ZN(n9850)
         );
  AOI21_X1 U10946 ( .B1(n9853), .B2(n9851), .A(n9850), .ZN(n9883) );
  INV_X1 U10947 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9852) );
  AOI22_X1 U10948 ( .A1(n9872), .A2(n9883), .B1(n9852), .B2(n9871), .ZN(
        P1_U3475) );
  NAND3_X1 U10949 ( .A1(n9855), .A2(n9854), .A3(n9853), .ZN(n9861) );
  AOI22_X1 U10950 ( .A1(n9858), .A2(n9857), .B1(n9856), .B2(n6314), .ZN(n9859)
         );
  AND3_X1 U10951 ( .A1(n9861), .A2(n9860), .A3(n9859), .ZN(n9884) );
  AOI22_X1 U10952 ( .A1(n9872), .A2(n9884), .B1(n5264), .B2(n9871), .ZN(
        P1_U3478) );
  INV_X1 U10953 ( .A(n9862), .ZN(n9869) );
  OAI22_X1 U10954 ( .A1(n9866), .A2(n9865), .B1(n9864), .B2(n9863), .ZN(n9868)
         );
  AOI211_X1 U10955 ( .C1(n9870), .C2(n9869), .A(n9868), .B(n9867), .ZN(n9886)
         );
  AOI22_X1 U10956 ( .A1(n9872), .A2(n9886), .B1(n5242), .B2(n9871), .ZN(
        P1_U3481) );
  AOI22_X1 U10957 ( .A1(n9887), .A2(n9874), .B1(n9873), .B2(n9885), .ZN(
        P1_U3524) );
  AOI22_X1 U10958 ( .A1(n9887), .A2(n9876), .B1(n9875), .B2(n9885), .ZN(
        P1_U3525) );
  AOI22_X1 U10959 ( .A1(n9887), .A2(n9877), .B1(n6600), .B2(n9885), .ZN(
        P1_U3526) );
  AOI22_X1 U10960 ( .A1(n9887), .A2(n9878), .B1(n6603), .B2(n9885), .ZN(
        P1_U3527) );
  INV_X1 U10961 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n9879) );
  AOI22_X1 U10962 ( .A1(n9887), .A2(n9880), .B1(n9879), .B2(n9885), .ZN(
        P1_U3528) );
  AOI22_X1 U10963 ( .A1(n9887), .A2(n9881), .B1(n6606), .B2(n9885), .ZN(
        P1_U3529) );
  INV_X1 U10964 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n9882) );
  AOI22_X1 U10965 ( .A1(n9887), .A2(n9883), .B1(n9882), .B2(n9885), .ZN(
        P1_U3530) );
  AOI22_X1 U10966 ( .A1(n9887), .A2(n9884), .B1(n6608), .B2(n9885), .ZN(
        P1_U3531) );
  AOI22_X1 U10967 ( .A1(n9887), .A2(n9886), .B1(n5238), .B2(n9885), .ZN(
        P1_U3532) );
  AOI22_X1 U10968 ( .A1(n9889), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n9888), .ZN(n9900) );
  INV_X1 U10969 ( .A(n9890), .ZN(n9891) );
  AOI21_X1 U10970 ( .B1(n9892), .B2(P2_ADDR_REG_0__SCAN_IN), .A(n9891), .ZN(
        n9899) );
  OAI21_X1 U10971 ( .B1(n9894), .B2(P2_REG1_REG_0__SCAN_IN), .A(n9893), .ZN(
        n9897) );
  NOR2_X1 U10972 ( .A1(n9895), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n9896) );
  OAI21_X1 U10973 ( .B1(n9897), .B2(n9896), .A(P2_IR_REG_0__SCAN_IN), .ZN(
        n9898) );
  OAI211_X1 U10974 ( .C1(P2_IR_REG_0__SCAN_IN), .C2(n9900), .A(n9899), .B(
        n9898), .ZN(P2_U3245) );
  XOR2_X1 U10975 ( .A(n9901), .B(n9908), .Z(n9903) );
  AOI21_X1 U10976 ( .B1(n9903), .B2(n9922), .A(n9902), .ZN(n10021) );
  AOI22_X1 U10977 ( .A1(n9937), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n9904), .B2(
        n9925), .ZN(n9905) );
  OAI21_X1 U10978 ( .B1(n9906), .B2(n10020), .A(n9905), .ZN(n9907) );
  INV_X1 U10979 ( .A(n9907), .ZN(n9917) );
  OAI21_X1 U10980 ( .B1(n9910), .B2(n7991), .A(n9909), .ZN(n10024) );
  INV_X1 U10981 ( .A(n9911), .ZN(n9914) );
  OAI211_X1 U10982 ( .C1(n9914), .C2(n10020), .A(n9913), .B(n9912), .ZN(n10018) );
  INV_X1 U10983 ( .A(n10018), .ZN(n9915) );
  AOI22_X1 U10984 ( .A1(n10024), .A2(n9934), .B1(n9933), .B2(n9915), .ZN(n9916) );
  OAI211_X1 U10985 ( .C1(n9937), .C2(n10021), .A(n9917), .B(n9916), .ZN(
        P2_U3284) );
  NAND2_X1 U10986 ( .A1(n7618), .A2(n9918), .ZN(n9920) );
  XNOR2_X1 U10987 ( .A(n9920), .B(n9919), .ZN(n9923) );
  AOI21_X1 U10988 ( .B1(n9923), .B2(n9922), .A(n9921), .ZN(n9967) );
  AOI22_X1 U10989 ( .A1(n9925), .A2(n9924), .B1(P2_REG2_REG_3__SCAN_IN), .B2(
        n9937), .ZN(n9936) );
  XNOR2_X1 U10990 ( .A(n9926), .B(n7075), .ZN(n9970) );
  INV_X1 U10991 ( .A(n9927), .ZN(n9930) );
  INV_X1 U10992 ( .A(n9928), .ZN(n9929) );
  AOI211_X1 U10993 ( .C1(n9932), .C2(n9930), .A(n10004), .B(n9929), .ZN(n9964)
         );
  AOI222_X1 U10994 ( .A1(n9970), .A2(n9934), .B1(n9933), .B2(n9964), .C1(n9932), .C2(n9931), .ZN(n9935) );
  OAI211_X1 U10995 ( .C1(n9937), .C2(n9967), .A(n9936), .B(n9935), .ZN(
        P2_U3293) );
  AND2_X1 U10996 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n9948), .ZN(P2_U3297) );
  AND2_X1 U10997 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n9948), .ZN(P2_U3298) );
  AND2_X1 U10998 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n9948), .ZN(P2_U3299) );
  AND2_X1 U10999 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n9948), .ZN(P2_U3300) );
  AND2_X1 U11000 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n9948), .ZN(P2_U3301) );
  AND2_X1 U11001 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n9948), .ZN(P2_U3302) );
  AND2_X1 U11002 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n9948), .ZN(P2_U3303) );
  AND2_X1 U11003 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n9948), .ZN(P2_U3304) );
  AND2_X1 U11004 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n9948), .ZN(P2_U3305) );
  AND2_X1 U11005 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n9948), .ZN(P2_U3306) );
  AND2_X1 U11006 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n9948), .ZN(P2_U3307) );
  AND2_X1 U11007 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n9948), .ZN(P2_U3308) );
  AND2_X1 U11008 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n9948), .ZN(P2_U3309) );
  AND2_X1 U11009 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n9948), .ZN(P2_U3310) );
  AND2_X1 U11010 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n9948), .ZN(P2_U3311) );
  NOR2_X1 U11011 ( .A1(n9944), .A2(n9940), .ZN(P2_U3312) );
  AND2_X1 U11012 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n9948), .ZN(P2_U3313) );
  AND2_X1 U11013 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n9948), .ZN(P2_U3314) );
  NOR2_X1 U11014 ( .A1(n9944), .A2(n9941), .ZN(P2_U3315) );
  NOR2_X1 U11015 ( .A1(n9944), .A2(n9942), .ZN(P2_U3316) );
  AND2_X1 U11016 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n9948), .ZN(P2_U3317) );
  AND2_X1 U11017 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n9948), .ZN(P2_U3318) );
  AND2_X1 U11018 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n9948), .ZN(P2_U3319) );
  AND2_X1 U11019 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n9948), .ZN(P2_U3320) );
  AND2_X1 U11020 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n9948), .ZN(P2_U3321) );
  AND2_X1 U11021 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n9948), .ZN(P2_U3322) );
  AND2_X1 U11022 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n9948), .ZN(P2_U3323) );
  AND2_X1 U11023 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n9948), .ZN(P2_U3324) );
  NOR2_X1 U11024 ( .A1(n9944), .A2(n9943), .ZN(P2_U3325) );
  AND2_X1 U11025 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n9948), .ZN(P2_U3326) );
  NOR2_X1 U11026 ( .A1(n9945), .A2(P2_U3152), .ZN(n9950) );
  AOI22_X1 U11027 ( .A1(n9947), .A2(n9950), .B1(n9946), .B2(n9948), .ZN(
        P2_U3437) );
  AOI22_X1 U11028 ( .A1(n9951), .A2(n9950), .B1(n9949), .B2(n9948), .ZN(
        P2_U3438) );
  AOI22_X1 U11029 ( .A1(n9954), .A2(n10025), .B1(n9953), .B2(n9952), .ZN(n9955) );
  AND2_X1 U11030 ( .A1(n9956), .A2(n9955), .ZN(n10030) );
  INV_X1 U11031 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n9957) );
  AOI22_X1 U11032 ( .A1(n10028), .A2(n10030), .B1(n9957), .B2(n10026), .ZN(
        P2_U3451) );
  INV_X1 U11033 ( .A(n9958), .ZN(n9959) );
  OAI22_X1 U11034 ( .A1(n9959), .A2(n10004), .B1(n7070), .B2(n10019), .ZN(
        n9961) );
  AOI211_X1 U11035 ( .C1(n10025), .C2(n9962), .A(n9961), .B(n9960), .ZN(n10032) );
  INV_X1 U11036 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n9963) );
  AOI22_X1 U11037 ( .A1(n10028), .A2(n10032), .B1(n9963), .B2(n10026), .ZN(
        P2_U3457) );
  INV_X1 U11038 ( .A(n9964), .ZN(n9965) );
  OAI21_X1 U11039 ( .B1(n9966), .B2(n10019), .A(n9965), .ZN(n9969) );
  INV_X1 U11040 ( .A(n9967), .ZN(n9968) );
  AOI211_X1 U11041 ( .C1(n10025), .C2(n9970), .A(n9969), .B(n9968), .ZN(n10033) );
  AOI22_X1 U11042 ( .A1(n10028), .A2(n10033), .B1(n9971), .B2(n10026), .ZN(
        P2_U3460) );
  OAI22_X1 U11043 ( .A1(n9973), .A2(n10004), .B1(n9972), .B2(n10019), .ZN(
        n9975) );
  AOI211_X1 U11044 ( .C1(n10025), .C2(n9976), .A(n9975), .B(n9974), .ZN(n10034) );
  INV_X1 U11045 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n9977) );
  AOI22_X1 U11046 ( .A1(n10028), .A2(n10034), .B1(n9977), .B2(n10026), .ZN(
        P2_U3469) );
  AND2_X1 U11047 ( .A1(n9978), .A2(n10025), .ZN(n9982) );
  OAI22_X1 U11048 ( .A1(n9980), .A2(n10004), .B1(n9979), .B2(n10019), .ZN(
        n9981) );
  NOR3_X1 U11049 ( .A1(n9983), .A2(n9982), .A3(n9981), .ZN(n10035) );
  INV_X1 U11050 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n9984) );
  AOI22_X1 U11051 ( .A1(n10028), .A2(n10035), .B1(n9984), .B2(n10026), .ZN(
        P2_U3472) );
  NOR2_X1 U11052 ( .A1(n9985), .A2(n10001), .ZN(n9991) );
  OAI22_X1 U11053 ( .A1(n9987), .A2(n10004), .B1(n9986), .B2(n10019), .ZN(
        n9989) );
  AOI211_X1 U11054 ( .C1(n9991), .C2(n9990), .A(n9989), .B(n9988), .ZN(n10036)
         );
  INV_X1 U11055 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n9992) );
  AOI22_X1 U11056 ( .A1(n10028), .A2(n10036), .B1(n9992), .B2(n10026), .ZN(
        P2_U3475) );
  INV_X1 U11057 ( .A(n9993), .ZN(n9998) );
  OAI22_X1 U11058 ( .A1(n9995), .A2(n10004), .B1(n9994), .B2(n10019), .ZN(
        n9997) );
  AOI211_X1 U11059 ( .C1(n9999), .C2(n9998), .A(n9997), .B(n9996), .ZN(n10037)
         );
  INV_X1 U11060 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10000) );
  AOI22_X1 U11061 ( .A1(n10028), .A2(n10037), .B1(n10000), .B2(n10026), .ZN(
        P2_U3478) );
  NOR2_X1 U11062 ( .A1(n10002), .A2(n10001), .ZN(n10009) );
  OAI22_X1 U11063 ( .A1(n10005), .A2(n10004), .B1(n10003), .B2(n10019), .ZN(
        n10007) );
  AOI211_X1 U11064 ( .C1(n10009), .C2(n10008), .A(n10007), .B(n10006), .ZN(
        n10039) );
  INV_X1 U11065 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10010) );
  AOI22_X1 U11066 ( .A1(n10028), .A2(n10039), .B1(n10010), .B2(n10026), .ZN(
        P2_U3481) );
  INV_X1 U11067 ( .A(n10011), .ZN(n10016) );
  OAI21_X1 U11068 ( .B1(n10013), .B2(n10019), .A(n10012), .ZN(n10015) );
  AOI211_X1 U11069 ( .C1(n10016), .C2(n10025), .A(n10015), .B(n10014), .ZN(
        n10041) );
  INV_X1 U11070 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10017) );
  AOI22_X1 U11071 ( .A1(n10028), .A2(n10041), .B1(n10017), .B2(n10026), .ZN(
        P2_U3484) );
  OAI21_X1 U11072 ( .B1(n10020), .B2(n10019), .A(n10018), .ZN(n10023) );
  INV_X1 U11073 ( .A(n10021), .ZN(n10022) );
  AOI211_X1 U11074 ( .C1(n10025), .C2(n10024), .A(n10023), .B(n10022), .ZN(
        n10044) );
  INV_X1 U11075 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10027) );
  AOI22_X1 U11076 ( .A1(n10028), .A2(n10044), .B1(n10027), .B2(n10026), .ZN(
        P2_U3487) );
  AOI22_X1 U11077 ( .A1(n10045), .A2(n10030), .B1(n10029), .B2(n10042), .ZN(
        P2_U3520) );
  AOI22_X1 U11078 ( .A1(n10045), .A2(n10032), .B1(n10031), .B2(n10042), .ZN(
        P2_U3522) );
  AOI22_X1 U11079 ( .A1(n10045), .A2(n10033), .B1(n6255), .B2(n10042), .ZN(
        P2_U3523) );
  AOI22_X1 U11080 ( .A1(n10045), .A2(n10034), .B1(n6251), .B2(n10042), .ZN(
        P2_U3526) );
  AOI22_X1 U11081 ( .A1(n10045), .A2(n10035), .B1(n6249), .B2(n10042), .ZN(
        P2_U3527) );
  AOI22_X1 U11082 ( .A1(n10045), .A2(n10036), .B1(n6262), .B2(n10042), .ZN(
        P2_U3528) );
  AOI22_X1 U11083 ( .A1(n10045), .A2(n10037), .B1(n6247), .B2(n10042), .ZN(
        P2_U3529) );
  AOI22_X1 U11084 ( .A1(n10045), .A2(n10039), .B1(n10038), .B2(n10042), .ZN(
        P2_U3530) );
  AOI22_X1 U11085 ( .A1(n10045), .A2(n10041), .B1(n10040), .B2(n10042), .ZN(
        P2_U3531) );
  AOI22_X1 U11086 ( .A1(n10045), .A2(n10044), .B1(n10043), .B2(n10042), .ZN(
        P2_U3532) );
  INV_X1 U11087 ( .A(n10046), .ZN(n10047) );
  NAND2_X1 U11088 ( .A1(n10048), .A2(n10047), .ZN(n10049) );
  XNOR2_X1 U11089 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n10049), .ZN(ADD_1071_U5)
         );
  XOR2_X1 U11090 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  OAI21_X1 U11091 ( .B1(n10052), .B2(n10051), .A(n10050), .ZN(ADD_1071_U56) );
  OAI21_X1 U11092 ( .B1(n10055), .B2(n10054), .A(n10053), .ZN(ADD_1071_U57) );
  OAI21_X1 U11093 ( .B1(n10058), .B2(n10057), .A(n10056), .ZN(ADD_1071_U58) );
  OAI21_X1 U11094 ( .B1(n10061), .B2(n10060), .A(n10059), .ZN(ADD_1071_U59) );
  OAI21_X1 U11095 ( .B1(n10064), .B2(n10063), .A(n10062), .ZN(ADD_1071_U60) );
  OAI21_X1 U11096 ( .B1(n10067), .B2(n10066), .A(n10065), .ZN(ADD_1071_U61) );
  AOI21_X1 U11097 ( .B1(n10070), .B2(n10069), .A(n10068), .ZN(ADD_1071_U62) );
  AOI21_X1 U11098 ( .B1(n10073), .B2(n10072), .A(n10071), .ZN(ADD_1071_U63) );
  XOR2_X1 U11099 ( .A(n10074), .B(P2_ADDR_REG_6__SCAN_IN), .Z(ADD_1071_U50) );
  NOR2_X1 U11100 ( .A1(n10076), .A2(n10075), .ZN(n10077) );
  XOR2_X1 U11101 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n10077), .Z(ADD_1071_U51) );
  OAI21_X1 U11102 ( .B1(n10080), .B2(n10079), .A(n10078), .ZN(n10081) );
  XNOR2_X1 U11103 ( .A(n10081), .B(P1_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  XNOR2_X1 U11104 ( .A(n10083), .B(n10082), .ZN(ADD_1071_U49) );
  AOI21_X1 U11105 ( .B1(n10086), .B2(n10085), .A(n10084), .ZN(ADD_1071_U47) );
  XOR2_X1 U11106 ( .A(n10088), .B(n10087), .Z(ADD_1071_U54) );
  XOR2_X1 U11107 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n10089), .Z(ADD_1071_U48) );
  XOR2_X1 U11108 ( .A(n10091), .B(n10090), .Z(ADD_1071_U53) );
  XNOR2_X1 U11109 ( .A(n10093), .B(n10092), .ZN(ADD_1071_U52) );
  XNOR2_X1 U6532 ( .A(n5037), .B(P1_IR_REG_30__SCAN_IN), .ZN(n5035) );
  NAND2_X1 U6698 ( .A1(n5191), .A2(n4313), .ZN(n9733) );
  CLKBUF_X1 U4811 ( .A(n6148), .Z(n6721) );
  XOR2_X1 U4924 ( .A(n4995), .B(P1_IR_REG_27__SCAN_IN), .Z(n10096) );
endmodule

