

module b21_C_AntiSAT_k_128_6 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3, 
        keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, 
        keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, 
        keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, 
        keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, 
        keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, 
        keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, 
        keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, 
        keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, 
        keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, 
        keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, 
        keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, 
        keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, 
        keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, 
        keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, 
        keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, 
        keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, 
        keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, 
        keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, 
        keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, 
        keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, 
        keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, 
        keyinput125, keyinput126, keyinput127, ADD_1071_U4, ADD_1071_U55, 
        ADD_1071_U56, ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, 
        ADD_1071_U61, ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, 
        ADD_1071_U49, ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, 
        ADD_1071_U54, ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3323, P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, 
        P1_U3454, P1_U3457, P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, 
        P1_U3475, P1_U3478, P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, 
        P1_U3496, P1_U3499, P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, 
        P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, 
        P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, 
        P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, 
        P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, 
        P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, 
        P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, 
        P1_U3554, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3264, P1_U3263, P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, 
        P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, 
        P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, 
        P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, 
        P1_U3586, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3212, P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, 
        P2_U3357, P2_U3356, P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, 
        P2_U3350, P2_U3349, P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, 
        P2_U3343, P2_U3342, P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, 
        P2_U3336, P2_U3335, P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, 
        P2_U3329, P2_U3328, P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, 
        P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, 
        P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, 
        P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, 
        P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, 
        P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, 
        P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, 
        P2_U3493, P2_U3496, P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, 
        P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, 
        P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, 
        P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, 
        P2_U3530, P2_U3531, P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, 
        P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, 
        P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, 
        P2_U3551, P2_U3296, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, 
        P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, 
        P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, 
        P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, 
        P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, 
        P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, 
        P2_U3562, P2_U3563, P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, 
        P2_U3569, P2_U3570, P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, 
        P2_U3576, P2_U3577, P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, 
        P2_U3583, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, 
        P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, 
        P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, 
        P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, 
        P2_U3217, P2_U3216, P2_U3215, P2_U3152, P2_U3151, P2_U3966 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
         n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
         n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
         n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
         n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
         n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
         n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
         n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
         n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
         n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
         n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
         n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
         n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
         n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294,
         n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304,
         n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314,
         n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324,
         n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334,
         n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344,
         n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354,
         n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364,
         n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374,
         n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384,
         n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394,
         n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404,
         n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414,
         n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424,
         n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434,
         n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444,
         n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454,
         n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464,
         n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474,
         n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484,
         n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494,
         n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504,
         n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514,
         n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524,
         n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534,
         n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544,
         n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554,
         n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564,
         n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574,
         n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584,
         n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594,
         n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604,
         n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614,
         n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624,
         n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634,
         n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644,
         n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654,
         n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664,
         n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674,
         n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684,
         n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694,
         n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704,
         n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714,
         n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724,
         n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734,
         n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744,
         n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754,
         n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764,
         n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774,
         n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784,
         n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794,
         n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804,
         n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814,
         n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824,
         n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834,
         n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844,
         n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854,
         n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864,
         n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874,
         n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884,
         n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894,
         n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904,
         n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914,
         n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924,
         n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934,
         n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944,
         n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954,
         n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964,
         n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974,
         n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984,
         n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994,
         n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004,
         n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014,
         n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024,
         n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034,
         n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044,
         n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054,
         n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064,
         n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074,
         n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084,
         n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094,
         n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104,
         n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114,
         n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124,
         n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134,
         n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144,
         n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154,
         n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164,
         n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174,
         n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184,
         n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194,
         n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204,
         n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214,
         n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224,
         n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234,
         n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244,
         n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254,
         n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264,
         n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274,
         n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284,
         n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294,
         n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304,
         n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314,
         n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324,
         n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334,
         n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344,
         n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354,
         n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364,
         n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
         n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
         n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
         n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
         n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414,
         n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
         n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434,
         n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444,
         n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454,
         n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
         n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
         n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484,
         n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494,
         n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504,
         n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514,
         n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
         n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
         n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
         n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
         n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
         n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
         n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
         n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
         n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
         n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
         n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624,
         n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634,
         n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644,
         n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654,
         n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664,
         n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674,
         n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684,
         n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694,
         n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704,
         n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714,
         n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724,
         n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734,
         n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744,
         n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754,
         n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764,
         n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774,
         n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784,
         n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794,
         n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804,
         n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814,
         n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824,
         n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834,
         n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844,
         n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854,
         n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864,
         n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874,
         n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884,
         n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894,
         n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904,
         n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914,
         n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924,
         n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934,
         n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944,
         n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954,
         n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964,
         n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974,
         n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984,
         n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994,
         n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004,
         n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014,
         n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024,
         n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034,
         n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044,
         n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054,
         n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064,
         n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074,
         n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084,
         n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094,
         n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104,
         n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114,
         n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124,
         n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134,
         n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144,
         n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154,
         n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164,
         n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174,
         n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184,
         n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194,
         n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204,
         n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214,
         n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224,
         n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234,
         n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244,
         n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254,
         n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264,
         n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274,
         n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284,
         n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294,
         n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304,
         n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314,
         n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324,
         n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334,
         n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344,
         n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354,
         n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364,
         n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374,
         n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384,
         n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394,
         n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404,
         n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414,
         n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424,
         n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434,
         n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444,
         n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454,
         n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464,
         n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474,
         n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484,
         n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494,
         n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504,
         n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514,
         n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524,
         n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534,
         n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544,
         n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554,
         n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564,
         n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574,
         n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584,
         n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594,
         n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604,
         n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614,
         n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624,
         n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634,
         n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644,
         n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654,
         n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664,
         n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674,
         n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684,
         n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694,
         n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704,
         n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714,
         n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724,
         n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734,
         n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744,
         n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754,
         n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764,
         n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774,
         n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784,
         n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794,
         n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804,
         n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814,
         n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824,
         n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834,
         n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844,
         n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854,
         n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864,
         n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874,
         n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884,
         n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894,
         n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904,
         n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914,
         n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924,
         n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934,
         n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944,
         n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954,
         n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964,
         n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974,
         n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984,
         n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994,
         n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004,
         n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014,
         n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024,
         n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034,
         n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044,
         n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054,
         n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064,
         n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074,
         n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084,
         n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094,
         n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104,
         n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114,
         n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124,
         n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134,
         n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144,
         n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154,
         n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164,
         n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174,
         n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184,
         n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194,
         n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204,
         n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214,
         n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224,
         n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234,
         n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244,
         n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254,
         n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264,
         n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274,
         n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284,
         n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294,
         n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304,
         n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314,
         n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324,
         n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334,
         n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344,
         n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354,
         n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364,
         n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374,
         n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384,
         n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394,
         n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404,
         n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414,
         n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424,
         n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434,
         n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444,
         n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454,
         n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464,
         n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474,
         n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484,
         n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494,
         n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504,
         n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514,
         n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524,
         n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534,
         n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544,
         n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554,
         n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564,
         n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574,
         n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584,
         n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594,
         n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604,
         n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614,
         n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624,
         n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634,
         n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644,
         n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654,
         n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664,
         n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674,
         n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684,
         n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694,
         n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704,
         n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714,
         n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724,
         n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734,
         n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744,
         n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754,
         n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764,
         n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774,
         n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784,
         n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794,
         n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804,
         n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814,
         n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824,
         n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834,
         n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844,
         n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854,
         n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864,
         n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874,
         n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884,
         n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894,
         n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904,
         n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914,
         n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924,
         n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934,
         n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944,
         n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954,
         n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964,
         n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974,
         n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984,
         n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994,
         n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004,
         n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014,
         n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024,
         n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034,
         n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044,
         n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054,
         n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064,
         n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074,
         n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084,
         n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094,
         n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104,
         n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114,
         n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124,
         n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134,
         n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144,
         n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154,
         n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164,
         n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174,
         n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184,
         n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194,
         n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204,
         n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214,
         n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224,
         n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234,
         n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244,
         n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254,
         n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264,
         n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274,
         n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284,
         n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294,
         n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304,
         n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314,
         n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324,
         n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334,
         n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344,
         n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354,
         n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364,
         n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374,
         n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384,
         n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394,
         n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404,
         n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414,
         n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424,
         n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434,
         n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444,
         n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454,
         n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464,
         n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474,
         n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484,
         n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494,
         n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504,
         n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514,
         n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524,
         n9525, n9526, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535,
         n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545,
         n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555,
         n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565,
         n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575,
         n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585,
         n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595,
         n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605,
         n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615,
         n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625,
         n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635,
         n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645,
         n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655,
         n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665,
         n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675,
         n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685,
         n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695,
         n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705,
         n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715,
         n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725,
         n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735,
         n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745,
         n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755,
         n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765,
         n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775,
         n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785,
         n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795,
         n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805,
         n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815,
         n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825,
         n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835,
         n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845,
         n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855,
         n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865,
         n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875,
         n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885,
         n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895,
         n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905,
         n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915,
         n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925,
         n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935,
         n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945,
         n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955,
         n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965,
         n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975,
         n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985,
         n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995,
         n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004,
         n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012,
         n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020,
         n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028,
         n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036,
         n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044,
         n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052,
         n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060,
         n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068,
         n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076,
         n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084,
         n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092,
         n10093, n10094, n10095, n10096, n10097;

  NAND2_X1 U4820 ( .A1(n8791), .A2(n4767), .ZN(n4766) );
  OAI22_X1 U4821 ( .A1(n7692), .A2(n8187), .B1(n7691), .B2(n8373), .ZN(n7722)
         );
  CLKBUF_X2 U4822 ( .A(n5873), .Z(n6197) );
  INV_X1 U4824 ( .A(n6290), .ZN(n6302) );
  AND4_X1 U4825 ( .A1(n5768), .A2(n5767), .A3(n5766), .A4(n5765), .ZN(n7134)
         );
  INV_X1 U4826 ( .A(n7026), .ZN(n8826) );
  OR3_X2 U4827 ( .A1(n7933), .A2(n7802), .A3(n7828), .ZN(n6543) );
  NAND2_X2 U4828 ( .A1(n5620), .A2(n8364), .ZN(n6875) );
  INV_X1 U4829 ( .A(n8569), .ZN(n8356) );
  NAND2_X1 U4830 ( .A1(n4324), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4915) );
  CLKBUF_X1 U4831 ( .A(n8137), .Z(n4315) );
  NOR4_X1 U4832 ( .A1(n5617), .A2(n6860), .A3(n9802), .A4(n9759), .ZN(n8137)
         );
  AOI22_X1 U4833 ( .A1(n8705), .A2(n8704), .B1(n8889), .B2(n8698), .ZN(n4316)
         );
  AOI22_X1 U4834 ( .A1(n8705), .A2(n8704), .B1(n8889), .B2(n8698), .ZN(n8688)
         );
  OAI21_X1 U4835 ( .B1(n4527), .B2(n8026), .A(n8007), .ZN(n8705) );
  NOR2_X1 U4836 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n5671) );
  INV_X1 U4837 ( .A(n6209), .ZN(n5873) );
  NAND2_X2 U4838 ( .A1(n6642), .A2(n5755), .ZN(n6215) );
  AND2_X1 U4839 ( .A1(n4826), .A2(n4827), .ZN(n4825) );
  NAND2_X1 U4840 ( .A1(n8138), .A2(n4351), .ZN(n8063) );
  INV_X1 U4841 ( .A(n6215), .ZN(n6179) );
  NAND2_X1 U4842 ( .A1(n4432), .A2(n4793), .ZN(n5650) );
  NAND2_X1 U4843 ( .A1(n7936), .A2(n6775), .ZN(n6639) );
  INV_X1 U4844 ( .A(n7234), .ZN(n6618) );
  NAND2_X1 U4845 ( .A1(n8140), .A2(n8139), .ZN(n8138) );
  XNOR2_X1 U4846 ( .A(n5589), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8365) );
  AND2_X1 U4847 ( .A1(n5704), .A2(n5703), .ZN(n5743) );
  AND4_X1 U4848 ( .A1(n5783), .A2(n5782), .A3(n5781), .A4(n5780), .ZN(n7262)
         );
  INV_X1 U4849 ( .A(n5704), .ZN(n7937) );
  AOI21_X2 U4850 ( .B1(n6393), .B2(n6392), .A(n6391), .ZN(n6395) );
  INV_X1 U4851 ( .A(n7440), .ZN(n7296) );
  INV_X1 U4852 ( .A(n6246), .ZN(n4317) );
  AND2_X1 U4854 ( .A1(n5704), .A2(n5703), .ZN(n4319) );
  NAND2_X2 U4856 ( .A1(n4703), .A2(n4702), .ZN(n5513) );
  OR2_X1 U4857 ( .A1(n9414), .A2(n9413), .ZN(n9415) );
  NAND2_X1 U4858 ( .A1(n8636), .A2(n8640), .ZN(n8635) );
  AND2_X1 U4859 ( .A1(n6126), .A2(n4427), .ZN(n9066) );
  NAND2_X1 U4860 ( .A1(n9368), .A2(n7966), .ZN(n9350) );
  NAND2_X1 U4861 ( .A1(n4766), .A2(n4764), .ZN(n8744) );
  NAND2_X1 U4862 ( .A1(n7813), .A2(n5266), .ZN(n8093) );
  NAND2_X1 U4863 ( .A1(n7713), .A2(n4350), .ZN(n7813) );
  NAND2_X1 U4864 ( .A1(n7292), .A2(n6500), .ZN(n7387) );
  NAND2_X1 U4865 ( .A1(n5140), .A2(n5139), .ZN(n7772) );
  NAND2_X1 U4866 ( .A1(n5865), .A2(n5864), .ZN(n7520) );
  INV_X1 U4867 ( .A(n7487), .ZN(n7469) );
  NAND2_X1 U4868 ( .A1(n9130), .A2(n7173), .ZN(n6379) );
  NAND2_X1 U4871 ( .A1(n5036), .A2(n5035), .ZN(n5060) );
  OAI211_X1 U4872 ( .C1(n4987), .C2(n6671), .A(n4972), .B(n4971), .ZN(n7355)
         );
  NAND2_X1 U4873 ( .A1(n5801), .A2(n5655), .ZN(n6290) );
  INV_X1 U4874 ( .A(n5044), .ZN(n4321) );
  OR2_X1 U4875 ( .A1(n8199), .A2(n8356), .ZN(n8363) );
  NAND2_X4 U4876 ( .A1(n4493), .A2(n4492), .ZN(n4994) );
  INV_X2 U4877 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  AND2_X1 U4878 ( .A1(P2_ADDR_REG_19__SCAN_IN), .A2(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n7576) );
  OAI21_X1 U4879 ( .B1(n8360), .B2(n4464), .A(n4850), .ZN(n4560) );
  NAND2_X1 U4880 ( .A1(n8057), .A2(n5484), .ZN(n5491) );
  AND2_X1 U4881 ( .A1(n5487), .A2(n5486), .ZN(n8111) );
  AND2_X1 U4882 ( .A1(n8985), .A2(n8987), .ZN(n4660) );
  AOI21_X1 U4883 ( .B1(n4590), .B2(n4589), .A(n4587), .ZN(n8337) );
  NOR2_X1 U4884 ( .A1(n6485), .A2(n9282), .ZN(n4737) );
  NOR3_X1 U4885 ( .A1(n9064), .A2(n9066), .A3(n6130), .ZN(n8984) );
  NAND2_X1 U4886 ( .A1(n8635), .A2(n8010), .ZN(n8621) );
  NAND3_X1 U4887 ( .A1(n4473), .A2(n4472), .A3(n8319), .ZN(n8600) );
  NAND2_X1 U4888 ( .A1(n8744), .A2(n8003), .ZN(n8728) );
  OR2_X1 U4889 ( .A1(n9420), .A2(n9210), .ZN(n7977) );
  OAI21_X1 U4890 ( .B1(n7907), .B2(n7906), .A(n7908), .ZN(n7909) );
  NAND2_X1 U4891 ( .A1(n4439), .A2(n4440), .ZN(n7897) );
  NAND2_X1 U4892 ( .A1(n7872), .A2(n7871), .ZN(n7907) );
  NAND2_X1 U4893 ( .A1(n7715), .A2(n7714), .ZN(n7713) );
  NAND2_X1 U4894 ( .A1(n7745), .A2(n4674), .ZN(n4441) );
  OR2_X1 U4895 ( .A1(n7841), .A2(n7840), .ZN(n7872) );
  NAND2_X1 U4896 ( .A1(n6166), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n6204) );
  NAND2_X1 U4897 ( .A1(n4677), .A2(n4675), .ZN(n7715) );
  NAND2_X1 U4898 ( .A1(n7781), .A2(n7780), .ZN(n7837) );
  NOR2_X1 U4899 ( .A1(n9390), .A2(n9465), .ZN(n9375) );
  INV_X1 U4900 ( .A(n4862), .ZN(n4861) );
  NAND2_X1 U4901 ( .A1(n5460), .A2(n5459), .ZN(n5465) );
  OAI21_X1 U4902 ( .B1(n5449), .B2(n5448), .A(n5450), .ZN(n5460) );
  NAND2_X1 U4903 ( .A1(n7808), .A2(n8259), .ZN(n7696) );
  AND2_X1 U4904 ( .A1(n4747), .A2(n7452), .ZN(n4746) );
  AND2_X1 U4905 ( .A1(n7449), .A2(n7657), .ZN(n7450) );
  NOR2_X2 U4906 ( .A1(n7706), .A2(n9825), .ZN(n7043) );
  NOR2_X2 U4907 ( .A1(n6910), .A2(P2_U3152), .ZN(n5616) );
  OR2_X1 U4908 ( .A1(n7255), .A2(n7440), .ZN(n7390) );
  OAI21_X1 U4909 ( .B1(n6935), .B2(n6934), .A(n6495), .ZN(n7116) );
  INV_X1 U4910 ( .A(n7403), .ZN(n9794) );
  AND4_X1 U4911 ( .A1(n5835), .A2(n5834), .A3(n5833), .A4(n5832), .ZN(n7300)
         );
  AND4_X1 U4912 ( .A1(n5800), .A2(n5799), .A3(n5798), .A4(n5797), .ZN(n7441)
         );
  AND3_X1 U4913 ( .A1(n5043), .A2(n4466), .A3(n5042), .ZN(n7403) );
  AND3_X1 U4914 ( .A1(n5024), .A2(n5023), .A3(n4891), .ZN(n7195) );
  NAND4_X1 U4915 ( .A1(n5051), .A2(n5050), .A3(n5049), .A4(n5048), .ZN(n8810)
         );
  OAI211_X1 U4916 ( .C1(n4987), .C2(n6654), .A(n5000), .B(n4999), .ZN(n9749)
         );
  NAND2_X1 U4917 ( .A1(n5006), .A2(n5005), .ZN(n8379) );
  OAI211_X2 U4918 ( .C1(n6290), .C2(n6666), .A(n5734), .B(n5733), .ZN(n7234)
         );
  NAND2_X2 U4919 ( .A1(n5721), .A2(n6639), .ZN(n7304) );
  OR2_X1 U4920 ( .A1(n5929), .A2(n5928), .ZN(n5947) );
  AND2_X1 U4921 ( .A1(n4948), .A2(n4751), .ZN(n7026) );
  INV_X2 U4922 ( .A(n5801), .ZN(n6057) );
  INV_X1 U4923 ( .A(n5044), .ZN(n4320) );
  INV_X2 U4925 ( .A(n5044), .ZN(n8035) );
  NAND2_X1 U4926 ( .A1(n8202), .A2(n6820), .ZN(n8338) );
  NAND2_X4 U4927 ( .A1(n6249), .A2(n7983), .ZN(n5801) );
  XNOR2_X1 U4928 ( .A(n5662), .B(n5661), .ZN(n7933) );
  INV_X1 U4929 ( .A(n7930), .ZN(n5703) );
  NAND2_X1 U4930 ( .A1(n5702), .A2(n5701), .ZN(n7930) );
  OR2_X1 U4931 ( .A1(n5885), .A2(n5884), .ZN(n5904) );
  INV_X1 U4932 ( .A(n8365), .ZN(n6820) );
  NAND2_X1 U4933 ( .A1(n5654), .A2(n5653), .ZN(n4592) );
  NAND2_X1 U4934 ( .A1(n4942), .A2(n4941), .ZN(n8364) );
  XNOR2_X1 U4935 ( .A(n4932), .B(P2_IR_REG_20__SCAN_IN), .ZN(n8199) );
  XNOR2_X1 U4936 ( .A(n4929), .B(n4928), .ZN(n8201) );
  NAND2_X1 U4937 ( .A1(n5701), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5697) );
  AND2_X1 U4938 ( .A1(n5319), .A2(n5281), .ZN(n5317) );
  NAND2_X1 U4939 ( .A1(n4454), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5589) );
  OR2_X2 U4940 ( .A1(n4994), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8967) );
  AND2_X1 U4941 ( .A1(n5642), .A2(n5633), .ZN(n4434) );
  AND2_X1 U4942 ( .A1(n4435), .A2(n5646), .ZN(n4433) );
  NOR2_X2 U4943 ( .A1(n5016), .A2(n4856), .ZN(n5039) );
  AND2_X1 U4944 ( .A1(n4417), .A2(n4416), .ZN(n4926) );
  AND2_X1 U4945 ( .A1(n5643), .A2(n5674), .ZN(n4619) );
  AND2_X1 U4946 ( .A1(n4790), .A2(n5637), .ZN(n4639) );
  AND3_X1 U4947 ( .A1(n4638), .A2(n5634), .A3(n5635), .ZN(n5636) );
  NOR2_X1 U4948 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n4638) );
  NOR2_X2 U4949 ( .A1(P2_ADDR_REG_19__SCAN_IN), .A2(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n7577) );
  INV_X1 U4950 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n9959) );
  NOR2_X1 U4951 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n5644) );
  INV_X1 U4952 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5973) );
  NOR2_X1 U4953 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n4790) );
  NOR2_X1 U4954 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n5752) );
  INV_X1 U4955 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5182) );
  INV_X1 U4956 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5181) );
  INV_X1 U4957 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5591) );
  INV_X1 U4958 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n9893) );
  INV_X1 U4959 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5085) );
  INV_X4 U4960 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  INV_X1 U4961 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n4924) );
  INV_X1 U4962 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5251) );
  NOR2_X1 U4963 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n5631) );
  NAND2_X2 U4964 ( .A1(n6817), .A2(n7026), .ZN(n8224) );
  NAND2_X2 U4965 ( .A1(n7046), .A2(n8224), .ZN(n6818) );
  NAND2_X2 U4966 ( .A1(n7025), .A2(n8826), .ZN(n7046) );
  AND2_X4 U4967 ( .A1(n4919), .A2(n4918), .ZN(n5213) );
  NAND2_X2 U4968 ( .A1(n5649), .A2(n5648), .ZN(n6249) );
  AOI21_X2 U4969 ( .B1(n8621), .B2(n8628), .A(n8011), .ZN(n8606) );
  OAI211_X2 U4970 ( .C1(n6290), .C2(n6672), .A(n5754), .B(n5753), .ZN(n6308)
         );
  AND2_X2 U4971 ( .A1(n4919), .A2(n8970), .ZN(n4974) );
  AOI21_X2 U4972 ( .B1(n8728), .B2(n8005), .A(n8004), .ZN(n8716) );
  NAND3_X4 U4973 ( .A1(n4922), .A2(n4921), .A3(n4920), .ZN(n6817) );
  OAI21_X2 U4974 ( .B1(n8606), .B2(n8614), .A(n4770), .ZN(n8594) );
  INV_X1 U4975 ( .A(n4320), .ZN(n4322) );
  NOR2_X1 U4976 ( .A1(n8970), .A2(n4919), .ZN(n4973) );
  AND2_X1 U4977 ( .A1(n8965), .A2(n8970), .ZN(n4323) );
  AND2_X4 U4978 ( .A1(n8965), .A2(n8970), .ZN(n5020) );
  NOR2_X1 U4979 ( .A1(n4500), .A2(n5343), .ZN(n4499) );
  INV_X1 U4980 ( .A(n4706), .ZN(n4500) );
  AND2_X1 U4981 ( .A1(n4374), .A2(n4924), .ZN(n4704) );
  OAI21_X1 U4982 ( .B1(n8345), .B2(n8344), .A(n8343), .ZN(n8361) );
  OR2_X1 U4983 ( .A1(n5610), .A2(n8199), .ZN(n9825) );
  OR2_X1 U4984 ( .A1(n9429), .A2(n9278), .ZN(n9244) );
  NAND2_X1 U4985 ( .A1(n4459), .A2(n4573), .ZN(n8223) );
  NAND2_X1 U4986 ( .A1(n4574), .A2(n8322), .ZN(n4573) );
  NAND2_X1 U4987 ( .A1(n8207), .A2(n8209), .ZN(n4572) );
  AOI21_X1 U4988 ( .B1(n4365), .B2(n4578), .A(n4582), .ZN(n4577) );
  NAND2_X1 U4989 ( .A1(n8678), .A2(n8297), .ZN(n4582) );
  INV_X1 U4990 ( .A(n4579), .ZN(n4578) );
  OAI211_X1 U4991 ( .C1(n8305), .C2(n8322), .A(n8307), .B(n4463), .ZN(n4462)
         );
  AND2_X1 U4992 ( .A1(n8655), .A2(n4342), .ZN(n4463) );
  AND2_X1 U4993 ( .A1(n8309), .A2(n8308), .ZN(n4461) );
  AOI22_X1 U4994 ( .A1(n8318), .A2(n8317), .B1(n8316), .B2(n8338), .ZN(n4470)
         );
  NAND2_X1 U4995 ( .A1(n4563), .A2(n4561), .ZN(n8318) );
  INV_X1 U4996 ( .A(n4562), .ZN(n4561) );
  AND2_X1 U4997 ( .A1(n4861), .A2(n4408), .ZN(n4407) );
  NAND2_X1 U4998 ( .A1(n7697), .A2(n4409), .ZN(n4408) );
  INV_X1 U4999 ( .A(n7945), .ZN(n4802) );
  NAND2_X1 U5000 ( .A1(n5206), .A2(n5205), .ZN(n5222) );
  INV_X1 U5001 ( .A(n4479), .ZN(n4478) );
  OAI21_X1 U5002 ( .B1(n4481), .B2(n4480), .A(n5156), .ZN(n4479) );
  INV_X1 U5003 ( .A(n4451), .ZN(n4450) );
  OAI21_X1 U5004 ( .B1(n4699), .B2(n4336), .A(n4453), .ZN(n4451) );
  OR2_X1 U5005 ( .A1(n5176), .A2(n5175), .ZN(n4453) );
  NOR2_X1 U5006 ( .A1(n8858), .A2(n8630), .ZN(n4773) );
  NOR2_X1 U5007 ( .A1(n8863), .A2(n8867), .ZN(n4532) );
  OR2_X1 U5008 ( .A1(n6204), .A2(n6203), .ZN(n6243) );
  NOR2_X1 U5009 ( .A1(n7959), .A2(n4824), .ZN(n4823) );
  INV_X1 U5010 ( .A(n7957), .ZN(n4824) );
  NOR2_X1 U5011 ( .A1(n4838), .A2(n4843), .ZN(n4832) );
  NAND2_X1 U5012 ( .A1(n4339), .A2(n7953), .ZN(n4838) );
  AND2_X1 U5013 ( .A1(n6450), .A2(n6449), .ZN(n7970) );
  OR2_X1 U5014 ( .A1(n9317), .A2(n9452), .ZN(n4606) );
  OR2_X1 U5015 ( .A1(n9455), .A2(n9330), .ZN(n7967) );
  OR2_X1 U5016 ( .A1(n9452), .A2(n9055), .ZN(n9302) );
  OR2_X1 U5017 ( .A1(n7685), .A2(n7620), .ZN(n7618) );
  NAND2_X1 U5018 ( .A1(n4510), .A2(n5495), .ZN(n5519) );
  AOI21_X1 U5019 ( .B1(n4496), .B2(n4498), .A(n5362), .ZN(n4495) );
  NAND2_X1 U5020 ( .A1(n5250), .A2(n5249), .ZN(n5272) );
  NAND2_X1 U5021 ( .A1(n5248), .A2(n5247), .ZN(n5250) );
  NAND2_X1 U5022 ( .A1(n5161), .A2(n5160), .ZN(n5179) );
  NAND2_X1 U5023 ( .A1(n5108), .A2(n5107), .ZN(n5129) );
  NAND2_X1 U5024 ( .A1(n8093), .A2(n5308), .ZN(n5316) );
  NAND2_X1 U5025 ( .A1(n5527), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5564) );
  AND2_X1 U5026 ( .A1(n4926), .A2(n4928), .ZN(n4455) );
  INV_X1 U5027 ( .A(n5020), .ZN(n5627) );
  NOR2_X1 U5028 ( .A1(n8842), .A2(n8584), .ZN(n8577) );
  OR2_X1 U5029 ( .A1(n8847), .A2(n8595), .ZN(n8584) );
  OR2_X1 U5030 ( .A1(n8863), .A2(n8150), .ZN(n8314) );
  AND2_X1 U5031 ( .A1(n8319), .A2(n8317), .ZN(n8614) );
  NAND2_X1 U5032 ( .A1(n8314), .A2(n8315), .ZN(n8628) );
  AOI21_X1 U5033 ( .B1(n4761), .B2(n4325), .A(n4360), .ZN(n4760) );
  OR2_X1 U5034 ( .A1(n8879), .A2(n10075), .ZN(n8292) );
  NOR2_X1 U5035 ( .A1(n8706), .A2(n8884), .ZN(n8669) );
  NOR2_X1 U5036 ( .A1(n8794), .A2(n8783), .ZN(n8781) );
  NOR2_X1 U5037 ( .A1(n8765), .A2(n4768), .ZN(n4767) );
  INV_X1 U5038 ( .A(n8002), .ZN(n4768) );
  INV_X1 U5039 ( .A(n8754), .ZN(n9744) );
  NAND2_X1 U5040 ( .A1(n4935), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4932) );
  NAND2_X1 U5041 ( .A1(n4441), .A2(n4328), .ZN(n4439) );
  OAI21_X1 U5042 ( .B1(n9064), .B2(n9066), .A(n6130), .ZN(n8985) );
  XNOR2_X1 U5043 ( .A(n5737), .B(n6212), .ZN(n6833) );
  NAND2_X1 U5044 ( .A1(n5873), .A2(n9133), .ZN(n5736) );
  NAND3_X1 U5045 ( .A1(n9099), .A2(n4349), .A3(n9021), .ZN(n4652) );
  AND2_X1 U5046 ( .A1(n5726), .A2(n4896), .ZN(n6802) );
  AND2_X1 U5047 ( .A1(n9061), .A2(n9065), .ZN(n9064) );
  NAND2_X1 U5048 ( .A1(n6282), .A2(n6281), .ZN(n9193) );
  NOR2_X1 U5049 ( .A1(n4594), .A2(n7986), .ZN(n4593) );
  NAND2_X1 U5050 ( .A1(n4596), .A2(n4828), .ZN(n4594) );
  OAI21_X1 U5051 ( .B1(n9229), .B2(n4631), .A(n4629), .ZN(n7981) );
  NAND2_X1 U5052 ( .A1(n7959), .A2(n7978), .ZN(n4631) );
  NAND2_X1 U5053 ( .A1(n4630), .A2(n7978), .ZN(n4629) );
  INV_X1 U5054 ( .A(n4632), .ZN(n4630) );
  NAND2_X1 U5055 ( .A1(n4828), .A2(n9210), .ZN(n4827) );
  OR2_X1 U5056 ( .A1(n9429), .A2(n9248), .ZN(n7955) );
  AND2_X1 U5057 ( .A1(n4788), .A2(n7785), .ZN(n4787) );
  AOI21_X1 U5058 ( .B1(n6619), .B2(n7224), .A(n4359), .ZN(n6930) );
  AND2_X1 U5059 ( .A1(n6631), .A2(n6803), .ZN(n9401) );
  NAND2_X1 U5060 ( .A1(n6165), .A2(n6164), .ZN(n9424) );
  NAND2_X1 U5061 ( .A1(n7888), .A2(n5751), .ZN(n6165) );
  NAND2_X1 U5062 ( .A1(n4506), .A2(n4503), .ZN(n7823) );
  NAND2_X1 U5063 ( .A1(n4510), .A2(n4504), .ZN(n4503) );
  NOR2_X1 U5064 ( .A1(n5518), .A2(n4505), .ZN(n4504) );
  AND2_X1 U5065 ( .A1(n5678), .A2(n5676), .ZN(n6775) );
  XNOR2_X1 U5066 ( .A(n5061), .B(n5037), .ZN(n5059) );
  AOI21_X1 U5067 ( .B1(n8562), .B2(n8563), .A(n8561), .ZN(n8564) );
  OR2_X1 U5068 ( .A1(n6875), .A2(n6892), .ZN(n4971) );
  NAND2_X1 U5069 ( .A1(n6175), .A2(n6174), .ZN(n9264) );
  OR2_X1 U5070 ( .A1(n9090), .A2(n6095), .ZN(n6175) );
  AND2_X1 U5071 ( .A1(n8239), .A2(n8238), .ZN(n8240) );
  NAND2_X1 U5072 ( .A1(n4340), .A2(n8235), .ZN(n4468) );
  OAI21_X1 U5073 ( .B1(n8264), .B2(n4569), .A(n8261), .ZN(n4568) );
  INV_X1 U5074 ( .A(n8259), .ZN(n4569) );
  NOR2_X1 U5075 ( .A1(n8260), .A2(n8338), .ZN(n4567) );
  NAND2_X1 U5076 ( .A1(n8265), .A2(n8338), .ZN(n4570) );
  NAND2_X1 U5077 ( .A1(n4363), .A2(n4580), .ZN(n4579) );
  NAND2_X1 U5078 ( .A1(n8295), .A2(n4581), .ZN(n4580) );
  INV_X1 U5079 ( .A(n8291), .ZN(n4581) );
  OR2_X1 U5080 ( .A1(n8319), .A2(n8322), .ZN(n8320) );
  AOI21_X1 U5081 ( .B1(n4869), .B2(n8194), .A(n4873), .ZN(n4867) );
  NAND2_X1 U5082 ( .A1(n4608), .A2(n7227), .ZN(n6494) );
  INV_X1 U5083 ( .A(n6266), .ZN(n4734) );
  AOI21_X1 U5084 ( .B1(n4733), .B2(n6266), .A(n4387), .ZN(n4732) );
  INV_X1 U5085 ( .A(n5605), .ZN(n4733) );
  NAND2_X1 U5086 ( .A1(n5274), .A2(n5273), .ZN(n5277) );
  INV_X1 U5087 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5637) );
  NAND2_X1 U5088 ( .A1(n8198), .A2(n4446), .ZN(n4447) );
  AND2_X1 U5089 ( .A1(n5610), .A2(n8201), .ZN(n4446) );
  INV_X1 U5090 ( .A(n8201), .ZN(n8346) );
  AND2_X1 U5091 ( .A1(n4865), .A2(n4871), .ZN(n4864) );
  NAND2_X1 U5092 ( .A1(n4872), .A2(n8350), .ZN(n4871) );
  NAND2_X1 U5093 ( .A1(n4867), .A2(n4868), .ZN(n4865) );
  INV_X1 U5094 ( .A(n8351), .ZN(n4872) );
  INV_X1 U5095 ( .A(SI_11_), .ZN(n10058) );
  AND2_X1 U5096 ( .A1(n8034), .A2(n8325), .ZN(n4869) );
  NAND2_X1 U5097 ( .A1(n4471), .A2(n8321), .ZN(n8588) );
  NAND2_X1 U5098 ( .A1(n8600), .A2(n4779), .ZN(n4471) );
  OR2_X1 U5099 ( .A1(n8852), .A2(n8149), .ZN(n8321) );
  AND2_X1 U5100 ( .A1(n8614), .A2(n4847), .ZN(n4846) );
  NAND2_X1 U5101 ( .A1(n8628), .A2(n8314), .ZN(n4847) );
  INV_X1 U5102 ( .A(n4761), .ZN(n4755) );
  OR2_X1 U5103 ( .A1(n8867), .A2(n8088), .ZN(n8311) );
  NOR2_X1 U5104 ( .A1(n8677), .A2(n4762), .ZN(n4761) );
  NOR2_X1 U5105 ( .A1(n4325), .A2(n8008), .ZN(n4762) );
  NAND2_X1 U5106 ( .A1(n4877), .A2(n8769), .ZN(n4875) );
  NOR2_X1 U5107 ( .A1(n8899), .A2(n8905), .ZN(n4528) );
  NOR2_X1 U5108 ( .A1(n8753), .A2(n4878), .ZN(n4877) );
  INV_X1 U5109 ( .A(n8285), .ZN(n4878) );
  OR2_X1 U5110 ( .A1(n5327), .A2(n8533), .ZN(n5350) );
  AOI21_X1 U5111 ( .B1(n4861), .B2(n4863), .A(n4860), .ZN(n4859) );
  NAND2_X1 U5112 ( .A1(n4407), .A2(n4410), .ZN(n4406) );
  NOR2_X1 U5113 ( .A1(n8925), .A2(n4537), .ZN(n4535) );
  OR2_X1 U5114 ( .A1(n8918), .A2(n8001), .ZN(n8278) );
  NAND2_X1 U5115 ( .A1(n8928), .A2(n4534), .ZN(n4537) );
  AOI21_X1 U5116 ( .B1(n8247), .B2(n4403), .A(n4402), .ZN(n4401) );
  INV_X1 U5117 ( .A(n8246), .ZN(n4403) );
  INV_X1 U5118 ( .A(n8212), .ZN(n4398) );
  NAND2_X1 U5119 ( .A1(n7359), .A2(n9749), .ZN(n8212) );
  OAI21_X1 U5120 ( .B1(n7405), .B2(n8211), .A(n8214), .ZN(n8809) );
  NOR2_X1 U5121 ( .A1(n9005), .A2(n4650), .ZN(n4649) );
  INV_X1 U5122 ( .A(n6089), .ZN(n4650) );
  OR2_X1 U5123 ( .A1(n9214), .A2(n9231), .ZN(n6374) );
  INV_X1 U5124 ( .A(n6168), .ZN(n6166) );
  AND2_X1 U5125 ( .A1(n6441), .A2(n9260), .ZN(n7973) );
  NOR2_X1 U5126 ( .A1(n4801), .A2(n4797), .ZN(n4796) );
  INV_X1 U5127 ( .A(n7943), .ZN(n4797) );
  INV_X1 U5128 ( .A(n9381), .ZN(n4799) );
  AND2_X1 U5129 ( .A1(n6426), .A2(n7966), .ZN(n7964) );
  NAND2_X1 U5130 ( .A1(n9132), .A2(n6933), .ZN(n6492) );
  INV_X1 U5131 ( .A(n4606), .ZN(n4605) );
  INV_X1 U5132 ( .A(n9436), .ZN(n4604) );
  INV_X1 U5133 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5638) );
  NAND2_X1 U5134 ( .A1(n5604), .A2(n5603), .ZN(n5606) );
  OAI21_X1 U5135 ( .B1(n5519), .B2(n4727), .A(n4724), .ZN(n5604) );
  AOI21_X1 U5136 ( .B1(n4728), .B2(n4726), .A(n4725), .ZN(n4724) );
  INV_X1 U5137 ( .A(n4728), .ZN(n4727) );
  INV_X1 U5138 ( .A(n5543), .ZN(n4725) );
  AND2_X1 U5139 ( .A1(n5543), .A2(n5524), .ZN(n5541) );
  NAND2_X1 U5140 ( .A1(n5465), .A2(n4508), .ZN(n4510) );
  NAND4_X1 U5141 ( .A1(n4619), .A2(n6233), .A3(n5644), .A4(n5671), .ZN(n4794)
         );
  NAND2_X1 U5142 ( .A1(n5673), .A2(n4648), .ZN(n4647) );
  NAND2_X1 U5143 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), 
        .ZN(n4648) );
  AND2_X1 U5144 ( .A1(n5409), .A2(n5391), .ZN(n5407) );
  AOI21_X1 U5145 ( .B1(n4499), .B2(n4497), .A(n4380), .ZN(n4496) );
  INV_X1 U5146 ( .A(n4709), .ZN(n4497) );
  INV_X1 U5147 ( .A(n4499), .ZN(n4498) );
  AOI21_X1 U5148 ( .B1(n4709), .B2(n4712), .A(n4707), .ZN(n4706) );
  INV_X1 U5149 ( .A(n4714), .ZN(n4712) );
  INV_X1 U5150 ( .A(n5319), .ZN(n4707) );
  AOI21_X1 U5151 ( .B1(n4714), .B2(n4711), .A(n4710), .ZN(n4709) );
  INV_X1 U5152 ( .A(n4716), .ZN(n4711) );
  INV_X1 U5153 ( .A(n5317), .ZN(n4710) );
  AND2_X1 U5154 ( .A1(n5270), .A2(n4717), .ZN(n4716) );
  INV_X1 U5155 ( .A(n5300), .ZN(n4717) );
  AOI21_X1 U5156 ( .B1(n5271), .B2(n4716), .A(n4715), .ZN(n4714) );
  INV_X1 U5157 ( .A(n5277), .ZN(n4715) );
  INV_X1 U5158 ( .A(n5267), .ZN(n5271) );
  XNOR2_X1 U5159 ( .A(n5268), .B(SI_14_), .ZN(n5267) );
  AOI21_X1 U5160 ( .B1(n4485), .B2(n4487), .A(n4484), .ZN(n4483) );
  INV_X1 U5161 ( .A(n4487), .ZN(n4486) );
  INV_X1 U5162 ( .A(n5222), .ZN(n4484) );
  AND2_X1 U5163 ( .A1(n5249), .A2(n5228), .ZN(n5247) );
  NOR2_X1 U5164 ( .A1(n5202), .A2(n4491), .ZN(n4490) );
  INV_X1 U5165 ( .A(n5179), .ZN(n4491) );
  INV_X1 U5166 ( .A(n5199), .ZN(n5202) );
  XNOR2_X1 U5167 ( .A(n5200), .B(n10058), .ZN(n5199) );
  AOI21_X1 U5168 ( .B1(n4478), .B2(n4480), .A(n4476), .ZN(n4475) );
  INV_X1 U5169 ( .A(n5158), .ZN(n4476) );
  AND2_X1 U5170 ( .A1(n5179), .A2(n5163), .ZN(n5177) );
  OR2_X1 U5171 ( .A1(n5852), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n5859) );
  INV_X1 U5172 ( .A(n5062), .ZN(n4719) );
  INV_X1 U5173 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5632) );
  NAND2_X1 U5174 ( .A1(n5717), .A2(n4960), .ZN(n4966) );
  NAND2_X1 U5175 ( .A1(n7577), .A2(n4723), .ZN(n4493) );
  INV_X1 U5176 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4723) );
  NAND2_X1 U5177 ( .A1(n7576), .A2(n4722), .ZN(n4492) );
  INV_X1 U5178 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4722) );
  OR2_X1 U5179 ( .A1(n5169), .A2(n5168), .ZN(n5189) );
  AND2_X1 U5180 ( .A1(n8847), .A2(n8146), .ZN(n5612) );
  INV_X1 U5181 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n5116) );
  NAND2_X1 U5182 ( .A1(n5469), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5505) );
  INV_X1 U5183 ( .A(n5476), .ZN(n5469) );
  NAND2_X1 U5184 ( .A1(n7100), .A2(n7101), .ZN(n4700) );
  OR2_X1 U5185 ( .A1(n5117), .A2(n5116), .ZN(n5143) );
  NOR2_X1 U5186 ( .A1(n8119), .A2(n4698), .ZN(n4697) );
  INV_X1 U5187 ( .A(n5382), .ZN(n4698) );
  NAND2_X1 U5188 ( .A1(n4450), .A2(n4336), .ZN(n4448) );
  AOI21_X1 U5189 ( .B1(n7527), .B2(n4680), .A(n4679), .ZN(n4678) );
  INV_X1 U5190 ( .A(n7525), .ZN(n4680) );
  INV_X1 U5191 ( .A(n7580), .ZN(n4679) );
  INV_X1 U5192 ( .A(n7527), .ZN(n4681) );
  NOR2_X1 U5193 ( .A1(n8083), .A2(n4688), .ZN(n4687) );
  INV_X1 U5194 ( .A(n5489), .ZN(n4688) );
  NOR2_X1 U5195 ( .A1(n8388), .A2(n8387), .ZN(n8386) );
  NOR2_X1 U5196 ( .A1(n8386), .A2(n4548), .ZN(n8401) );
  AND2_X1 U5197 ( .A1(n8385), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n4548) );
  OR2_X1 U5198 ( .A1(n8401), .A2(n8402), .ZN(n4547) );
  NOR2_X1 U5199 ( .A1(n8414), .A2(n4378), .ZN(n8429) );
  OR2_X1 U5200 ( .A1(n8429), .A2(n8430), .ZN(n4549) );
  NOR2_X1 U5201 ( .A1(n8443), .A2(n8444), .ZN(n8442) );
  OR2_X1 U5202 ( .A1(n8457), .A2(n8458), .ZN(n4544) );
  AND2_X1 U5203 ( .A1(n4544), .A2(n4543), .ZN(n8471) );
  NAND2_X1 U5204 ( .A1(n8455), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n4543) );
  OR2_X1 U5205 ( .A1(n8471), .A2(n8472), .ZN(n4542) );
  AND2_X1 U5206 ( .A1(n5565), .A2(n8019), .ZN(n8586) );
  NAND2_X1 U5207 ( .A1(n8658), .A2(n4348), .ZN(n8595) );
  INV_X1 U5208 ( .A(n4773), .ZN(n4770) );
  INV_X1 U5209 ( .A(n8628), .ZN(n8620) );
  AND2_X1 U5210 ( .A1(n4880), .A2(n8032), .ZN(n4879) );
  OR2_X1 U5211 ( .A1(n4393), .A2(n8028), .ZN(n4390) );
  NAND2_X1 U5212 ( .A1(n4316), .A2(n4761), .ZN(n4759) );
  AND2_X1 U5213 ( .A1(n8670), .A2(n8663), .ZN(n8658) );
  NAND2_X1 U5214 ( .A1(n8676), .A2(n8031), .ZN(n8675) );
  NAND2_X1 U5215 ( .A1(n8675), .A2(n4882), .ZN(n8652) );
  AND2_X1 U5216 ( .A1(n8292), .A2(n8306), .ZN(n8677) );
  AND2_X1 U5217 ( .A1(n8669), .A2(n8674), .ZN(n8670) );
  NAND2_X1 U5218 ( .A1(n8693), .A2(n8029), .ZN(n8676) );
  OR2_X1 U5219 ( .A1(n8896), .A2(n8739), .ZN(n8006) );
  NAND2_X1 U5220 ( .A1(n8024), .A2(n8765), .ZN(n8772) );
  OR2_X1 U5221 ( .A1(n8925), .A2(n8161), .ZN(n8272) );
  NAND2_X1 U5222 ( .A1(n7726), .A2(n7700), .ZN(n8023) );
  NAND2_X1 U5223 ( .A1(n7724), .A2(n7697), .ZN(n7726) );
  NOR2_X1 U5224 ( .A1(n9748), .A2(n9749), .ZN(n4520) );
  AND2_X1 U5225 ( .A1(n4520), .A2(n9788), .ZN(n7400) );
  INV_X1 U5226 ( .A(n8379), .ZN(n7359) );
  NAND3_X1 U5227 ( .A1(n8217), .A2(n4855), .A3(n8224), .ZN(n9740) );
  OR2_X1 U5228 ( .A1(n6696), .A2(n5621), .ZN(n8754) );
  NAND2_X1 U5229 ( .A1(n8016), .A2(n8015), .ZN(n8842) );
  AND2_X1 U5230 ( .A1(n8780), .A2(n9809), .ZN(n9797) );
  AND2_X1 U5231 ( .A1(n5599), .A2(n5595), .ZN(n9758) );
  OR2_X1 U5232 ( .A1(n7824), .A2(n5594), .ZN(n5595) );
  NAND2_X1 U5233 ( .A1(n4941), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4525) );
  INV_X1 U5234 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n4417) );
  NAND2_X1 U5235 ( .A1(n4899), .A2(n4857), .ZN(n4856) );
  INV_X1 U5236 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n4857) );
  NAND2_X1 U5237 ( .A1(n7434), .A2(n5823), .ZN(n4672) );
  NAND2_X1 U5238 ( .A1(n4652), .A2(n4355), .ZN(n6054) );
  NAND2_X1 U5239 ( .A1(n9034), .A2(n4654), .ZN(n4653) );
  INV_X1 U5240 ( .A(n6020), .ZN(n4654) );
  INV_X1 U5241 ( .A(n4422), .ZN(n4421) );
  OAI21_X1 U5242 ( .B1(n5845), .B2(n5858), .A(n7536), .ZN(n4422) );
  NAND2_X1 U5243 ( .A1(n5693), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n6111) );
  INV_X1 U5244 ( .A(n6093), .ZN(n5693) );
  AOI21_X1 U5245 ( .B1(n4649), .B2(n4430), .A(n4377), .ZN(n4429) );
  INV_X1 U5246 ( .A(n6086), .ZN(n4430) );
  INV_X1 U5247 ( .A(n4649), .ZN(n4431) );
  AOI21_X1 U5248 ( .B1(n4643), .B2(n4645), .A(n4347), .ZN(n4640) );
  AND2_X1 U5249 ( .A1(n4666), .A2(n4662), .ZN(n4661) );
  NAND2_X1 U5250 ( .A1(n4660), .A2(n4657), .ZN(n4656) );
  NAND2_X1 U5251 ( .A1(n5992), .A2(n5991), .ZN(n9099) );
  NAND2_X1 U5252 ( .A1(n4439), .A2(n4436), .ZN(n5992) );
  NOR2_X1 U5253 ( .A1(n4438), .A2(n4437), .ZN(n4436) );
  AND4_X1 U5254 ( .A1(n5816), .A2(n5815), .A3(n5814), .A4(n5813), .ZN(n7297)
         );
  NAND2_X1 U5255 ( .A1(n4830), .A2(n4823), .ZN(n4829) );
  NAND2_X1 U5256 ( .A1(n9233), .A2(n7977), .ZN(n9207) );
  NAND2_X1 U5257 ( .A1(n9261), .A2(n7973), .ZN(n9245) );
  NAND2_X1 U5258 ( .A1(n9273), .A2(n7972), .ZN(n9261) );
  AOI21_X1 U5259 ( .B1(n4339), .B2(n4836), .A(n4835), .ZN(n4834) );
  NOR2_X1 U5260 ( .A1(n9436), .A2(n9265), .ZN(n4835) );
  NOR2_X1 U5261 ( .A1(n7954), .A2(n4840), .ZN(n4839) );
  INV_X1 U5262 ( .A(n7951), .ZN(n4840) );
  INV_X1 U5263 ( .A(n7953), .ZN(n4837) );
  NAND2_X1 U5264 ( .A1(n7970), .A2(n4626), .ZN(n4625) );
  INV_X1 U5265 ( .A(n7968), .ZN(n4626) );
  NAND2_X1 U5266 ( .A1(n7970), .A2(n4356), .ZN(n4624) );
  INV_X1 U5267 ( .A(n7969), .ZN(n4628) );
  NOR2_X1 U5268 ( .A1(n9344), .A2(n9452), .ZN(n9334) );
  OAI21_X1 U5269 ( .B1(n9343), .B2(n7948), .A(n7947), .ZN(n9325) );
  NAND2_X1 U5270 ( .A1(n7944), .A2(n7943), .ZN(n9374) );
  NAND2_X1 U5271 ( .A1(n7941), .A2(n7940), .ZN(n9389) );
  AND2_X1 U5272 ( .A1(n6418), .A2(n9397), .ZN(n7913) );
  OR2_X1 U5273 ( .A1(n7831), .A2(n4812), .ZN(n4807) );
  AOI21_X1 U5274 ( .B1(n4811), .B2(n4809), .A(n4366), .ZN(n4808) );
  INV_X1 U5275 ( .A(n4816), .ZN(n4809) );
  NOR2_X1 U5276 ( .A1(n7878), .A2(n4817), .ZN(n4816) );
  INV_X1 U5277 ( .A(n7829), .ZN(n4817) );
  OAI21_X1 U5278 ( .B1(n7878), .B2(n4815), .A(n7877), .ZN(n4814) );
  NAND2_X1 U5279 ( .A1(n7830), .A2(n7829), .ZN(n4815) );
  NAND2_X1 U5280 ( .A1(n4618), .A2(n7618), .ZN(n7759) );
  NAND2_X1 U5281 ( .A1(n7386), .A2(n4338), .ZN(n7365) );
  NAND2_X1 U5282 ( .A1(n7252), .A2(n6624), .ZN(n7290) );
  NOR2_X1 U5283 ( .A1(n7387), .A2(n4612), .ZN(n4613) );
  NOR2_X1 U5284 ( .A1(n7289), .A2(n4615), .ZN(n4612) );
  NAND2_X1 U5285 ( .A1(n7249), .A2(n4783), .ZN(n7299) );
  NOR2_X1 U5286 ( .A1(n6627), .A2(n4784), .ZN(n4783) );
  INV_X1 U5287 ( .A(n6626), .ZN(n4784) );
  AND2_X1 U5288 ( .A1(n7132), .A2(n6622), .ZN(n7250) );
  NAND2_X1 U5289 ( .A1(n6304), .A2(n6303), .ZN(n7986) );
  NAND2_X1 U5290 ( .A1(n6059), .A2(n6058), .ZN(n9460) );
  NAND2_X1 U5291 ( .A1(n6041), .A2(n6040), .ZN(n9465) );
  NAND2_X1 U5292 ( .A1(n5927), .A2(n5926), .ZN(n9482) );
  INV_X1 U5293 ( .A(n7538), .ZN(n7411) );
  AND2_X1 U5294 ( .A1(n6932), .A2(n6527), .ZN(n9483) );
  INV_X1 U5295 ( .A(n7247), .ZN(n9717) );
  AND2_X1 U5296 ( .A1(n7342), .A2(n6241), .ZN(n6932) );
  XNOR2_X1 U5297 ( .A(n6289), .B(n6288), .ZN(n8172) );
  NAND2_X1 U5298 ( .A1(n5659), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5666) );
  XNOR2_X1 U5299 ( .A(n5496), .B(n5492), .ZN(n7769) );
  NAND2_X1 U5300 ( .A1(n5465), .A2(n5464), .ZN(n5496) );
  NAND2_X1 U5301 ( .A1(n5106), .A2(n4481), .ZN(n4477) );
  XNOR2_X1 U5302 ( .A(n5082), .B(SI_6_), .ZN(n5080) );
  NAND2_X1 U5303 ( .A1(n5463), .A2(n5462), .ZN(n8873) );
  NAND2_X1 U5304 ( .A1(n5412), .A2(n5411), .ZN(n8884) );
  NAND2_X1 U5305 ( .A1(n5503), .A2(n5502), .ZN(n8863) );
  NAND2_X1 U5306 ( .A1(n7823), .A2(n8171), .ZN(n5503) );
  NAND2_X1 U5307 ( .A1(n5286), .A2(n5285), .ZN(n8783) );
  XNOR2_X1 U5308 ( .A(n8113), .B(n8115), .ZN(n4457) );
  NAND2_X1 U5309 ( .A1(n5434), .A2(n5433), .ZN(n8879) );
  NAND2_X1 U5310 ( .A1(n4465), .A2(n4851), .ZN(n4464) );
  NAND2_X1 U5311 ( .A1(n4853), .A2(n4852), .ZN(n4851) );
  NAND2_X1 U5312 ( .A1(n8361), .A2(n8362), .ZN(n4465) );
  NAND2_X1 U5313 ( .A1(n5513), .A2(n8358), .ZN(n4852) );
  NAND2_X1 U5314 ( .A1(n8198), .A2(n5610), .ZN(n8359) );
  NAND2_X1 U5315 ( .A1(n8565), .A2(n4557), .ZN(n4556) );
  INV_X1 U5316 ( .A(n4558), .ZN(n4557) );
  OAI21_X1 U5317 ( .B1(n8566), .B2(n9732), .A(n9730), .ZN(n4558) );
  NAND2_X1 U5318 ( .A1(n4555), .A2(n4554), .ZN(n4553) );
  INV_X1 U5319 ( .A(n8571), .ZN(n4554) );
  NAND2_X1 U5320 ( .A1(n9734), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n4555) );
  NAND2_X1 U5321 ( .A1(n4778), .A2(n4775), .ZN(n4774) );
  AND2_X1 U5322 ( .A1(n4776), .A2(n4772), .ZN(n4771) );
  AND2_X1 U5323 ( .A1(n4515), .A2(n4513), .ZN(n8845) );
  AOI21_X1 U5324 ( .B1(n8601), .B2(n9743), .A(n4514), .ZN(n4513) );
  NAND2_X1 U5325 ( .A1(n4516), .A2(n8813), .ZN(n4515) );
  AND2_X1 U5326 ( .A1(n8369), .A2(n8572), .ZN(n4514) );
  AND2_X1 U5327 ( .A1(n4414), .A2(n4411), .ZN(n8850) );
  AND2_X1 U5328 ( .A1(n4413), .A2(n4412), .ZN(n4411) );
  NAND2_X1 U5329 ( .A1(n4415), .A2(n8813), .ZN(n4414) );
  NAND2_X1 U5330 ( .A1(n8590), .A2(n9744), .ZN(n4412) );
  OR2_X1 U5331 ( .A1(n6653), .A2(n4987), .ZN(n4466) );
  NAND2_X1 U5332 ( .A1(n7042), .A2(n7668), .ZN(n8830) );
  NAND2_X1 U5333 ( .A1(n4884), .A2(n4913), .ZN(n4883) );
  INV_X1 U5334 ( .A(n4886), .ZN(n4884) );
  NAND2_X1 U5335 ( .A1(n4782), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4940) );
  AND4_X1 U5336 ( .A1(n5851), .A2(n5850), .A3(n5849), .A4(n5848), .ZN(n7480)
         );
  NAND2_X1 U5337 ( .A1(n7514), .A2(n7515), .ZN(n4642) );
  AND2_X1 U5338 ( .A1(n6157), .A2(n6156), .ZN(n9278) );
  OR2_X1 U5339 ( .A1(n9256), .A2(n6095), .ZN(n6157) );
  NAND2_X1 U5340 ( .A1(n4445), .A2(n4444), .ZN(n4443) );
  AOI21_X1 U5341 ( .B1(n4664), .B2(n4667), .A(n9089), .ZN(n4444) );
  NAND2_X1 U5342 ( .A1(n4670), .A2(n4665), .ZN(n4445) );
  AND2_X1 U5343 ( .A1(n4667), .A2(n4668), .ZN(n4665) );
  AND2_X1 U5344 ( .A1(n9088), .A2(n9087), .ZN(n4442) );
  INV_X1 U5345 ( .A(n9697), .ZN(n6767) );
  NOR2_X1 U5346 ( .A1(n4737), .A2(n7936), .ZN(n4736) );
  NAND2_X1 U5347 ( .A1(n4739), .A2(n9282), .ZN(n4738) );
  INV_X1 U5348 ( .A(n7480), .ZN(n9126) );
  INV_X1 U5349 ( .A(n7297), .ZN(n9128) );
  NAND2_X1 U5350 ( .A1(n6284), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5729) );
  NAND3_X1 U5351 ( .A1(n7937), .A2(n5703), .A3(P1_REG1_REG_0__SCAN_IN), .ZN(
        n5711) );
  OR2_X1 U5352 ( .A1(n5744), .A2(n5710), .ZN(n5712) );
  XNOR2_X1 U5353 ( .A(n7961), .B(n7980), .ZN(n7997) );
  AOI21_X1 U5354 ( .B1(n4825), .B2(n4821), .A(n4361), .ZN(n4820) );
  OR3_X1 U5355 ( .A1(n9238), .A2(n4822), .A3(n7958), .ZN(n4819) );
  AND2_X1 U5356 ( .A1(n4598), .A2(n4597), .ZN(n7996) );
  NAND2_X1 U5357 ( .A1(n4341), .A2(n7986), .ZN(n4598) );
  AND2_X1 U5358 ( .A1(n4637), .A2(n4636), .ZN(n7994) );
  AOI22_X1 U5359 ( .A1(n7960), .A2(n9401), .B1(n9194), .B2(n9117), .ZN(n4636)
         );
  NAND2_X1 U5360 ( .A1(n7985), .A2(n9406), .ZN(n4637) );
  INV_X1 U5361 ( .A(n6638), .ZN(n9321) );
  NAND3_X1 U5362 ( .A1(n9717), .A2(n9697), .A3(n7342), .ZN(n9692) );
  NAND2_X1 U5363 ( .A1(n8214), .A2(n8213), .ZN(n4574) );
  NOR2_X1 U5364 ( .A1(n8215), .A2(n4571), .ZN(n8216) );
  OAI21_X1 U5365 ( .B1(n8223), .B2(n4332), .A(n8214), .ZN(n4571) );
  NOR2_X1 U5366 ( .A1(n4458), .A2(n8210), .ZN(n8236) );
  OAI21_X1 U5367 ( .B1(n8223), .B2(n4358), .A(n8207), .ZN(n4458) );
  NAND2_X1 U5368 ( .A1(n8250), .A2(n8249), .ZN(n4565) );
  AND2_X1 U5369 ( .A1(n8247), .A2(n8241), .ZN(n4467) );
  NAND2_X1 U5370 ( .A1(n4570), .A2(n4566), .ZN(n8271) );
  NAND2_X1 U5371 ( .A1(n4568), .A2(n4567), .ZN(n4566) );
  NAND2_X1 U5372 ( .A1(n4576), .A2(n4575), .ZN(n8293) );
  AOI21_X1 U5373 ( .B1(n4577), .B2(n4579), .A(n4364), .ZN(n4575) );
  OAI21_X1 U5374 ( .B1(n8314), .B2(n8338), .A(n8319), .ZN(n4562) );
  NAND2_X1 U5375 ( .A1(n4460), .A2(n4564), .ZN(n4563) );
  AND2_X1 U5376 ( .A1(n8620), .A2(n8313), .ZN(n4564) );
  NAND2_X1 U5377 ( .A1(n4462), .A2(n4354), .ZN(n4460) );
  INV_X1 U5378 ( .A(n4869), .ZN(n4868) );
  NAND2_X1 U5379 ( .A1(n4591), .A2(n8329), .ZN(n4590) );
  NAND2_X1 U5380 ( .A1(n4779), .A2(n8320), .ZN(n4469) );
  NAND2_X1 U5381 ( .A1(n8034), .A2(n4588), .ZN(n4587) );
  NAND2_X1 U5382 ( .A1(n8331), .A2(n8338), .ZN(n4588) );
  NAND2_X1 U5383 ( .A1(n8328), .A2(n8338), .ZN(n4589) );
  OR2_X1 U5384 ( .A1(n8838), .A2(n8175), .ZN(n8351) );
  OR2_X1 U5385 ( .A1(n8842), .A2(n8017), .ZN(n8333) );
  INV_X1 U5386 ( .A(n7697), .ZN(n4410) );
  OAI21_X1 U5387 ( .B1(n7700), .B2(n4863), .A(n8275), .ZN(n4862) );
  INV_X1 U5388 ( .A(n8272), .ZN(n4863) );
  INV_X1 U5389 ( .A(n8278), .ZN(n4860) );
  AND2_X1 U5390 ( .A1(n7986), .A2(n9209), .ZN(n6366) );
  NOR2_X1 U5391 ( .A1(n9476), .A2(n9113), .ZN(n4601) );
  OR2_X1 U5392 ( .A1(n7764), .A2(n9482), .ZN(n7792) );
  AOI21_X1 U5393 ( .B1(n4732), .B2(n4734), .A(SI_29_), .ZN(n4731) );
  INV_X1 U5394 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5639) );
  AND2_X1 U5395 ( .A1(n4729), .A2(n5541), .ZN(n4728) );
  NAND2_X1 U5396 ( .A1(n5518), .A2(n5520), .ZN(n4729) );
  INV_X1 U5397 ( .A(n5520), .ZN(n4726) );
  INV_X1 U5398 ( .A(n5518), .ZN(n4507) );
  NOR2_X1 U5399 ( .A1(n5223), .A2(n4488), .ZN(n4487) );
  INV_X1 U5400 ( .A(n5201), .ZN(n4488) );
  INV_X1 U5401 ( .A(n4490), .ZN(n4485) );
  INV_X1 U5402 ( .A(n5129), .ZN(n4480) );
  AND2_X1 U5403 ( .A1(n5154), .A2(n5126), .ZN(n4699) );
  INV_X1 U5404 ( .A(n5155), .ZN(n4452) );
  INV_X1 U5405 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n4539) );
  NOR2_X1 U5406 ( .A1(n8858), .A2(n4531), .ZN(n4530) );
  INV_X1 U5407 ( .A(n4532), .ZN(n4531) );
  INV_X1 U5408 ( .A(n4393), .ZN(n4392) );
  NAND2_X1 U5409 ( .A1(n4882), .A2(n8029), .ZN(n4393) );
  NAND2_X1 U5410 ( .A1(n4882), .A2(n4881), .ZN(n4880) );
  INV_X1 U5411 ( .A(n8031), .ZN(n4881) );
  OR2_X1 U5412 ( .A1(n8889), .A2(n8077), .ZN(n8301) );
  NAND2_X1 U5413 ( .A1(n5348), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5373) );
  INV_X1 U5414 ( .A(n5350), .ZN(n5348) );
  NAND2_X1 U5415 ( .A1(n5289), .A2(n5288), .ZN(n5327) );
  INV_X1 U5416 ( .A(n5295), .ZN(n5289) );
  NAND2_X1 U5417 ( .A1(n5256), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5295) );
  INV_X1 U5418 ( .A(n5257), .ZN(n5256) );
  NAND2_X1 U5419 ( .A1(n7696), .A2(n8262), .ZN(n7724) );
  NAND2_X1 U5420 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5046) );
  OR2_X1 U5421 ( .A1(n6665), .A2(n4994), .ZN(n4750) );
  NAND2_X1 U5422 ( .A1(n4994), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n4749) );
  INV_X1 U5423 ( .A(n8380), .ZN(n6822) );
  NOR2_X1 U5424 ( .A1(n7666), .A2(n7772), .ZN(n7665) );
  NAND2_X1 U5425 ( .A1(n4518), .A2(n4517), .ZN(n7666) );
  INV_X1 U5426 ( .A(n7279), .ZN(n4518) );
  NAND2_X1 U5427 ( .A1(n4519), .A2(n7329), .ZN(n7279) );
  INV_X1 U5428 ( .A(n8816), .ZN(n4519) );
  INV_X1 U5429 ( .A(n5880), .ZN(n4645) );
  INV_X1 U5430 ( .A(n4644), .ZN(n4643) );
  OAI21_X1 U5431 ( .B1(n7515), .B2(n4645), .A(n7683), .ZN(n4644) );
  NOR2_X1 U5432 ( .A1(n4664), .A2(n9042), .ZN(n4657) );
  AND2_X1 U5433 ( .A1(n9089), .A2(n4667), .ZN(n4666) );
  NAND2_X1 U5434 ( .A1(n9013), .A2(n4663), .ZN(n4662) );
  INV_X1 U5435 ( .A(n4668), .ZN(n4663) );
  INV_X1 U5436 ( .A(n4367), .ZN(n4438) );
  INV_X1 U5437 ( .A(n4440), .ZN(n4437) );
  NOR2_X1 U5438 ( .A1(n4826), .A2(n4633), .ZN(n4632) );
  INV_X1 U5439 ( .A(n7977), .ZN(n4633) );
  AND2_X1 U5440 ( .A1(n6446), .A2(n9272), .ZN(n7972) );
  NOR2_X1 U5441 ( .A1(n4839), .A2(n4837), .ZN(n4836) );
  INV_X1 U5442 ( .A(n7949), .ZN(n4844) );
  NAND2_X1 U5443 ( .A1(n5689), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n5980) );
  INV_X1 U5444 ( .A(n5960), .ZN(n5689) );
  NAND2_X1 U5445 ( .A1(n7756), .A2(n7757), .ZN(n4788) );
  NOR2_X1 U5446 ( .A1(n6343), .A2(n7497), .ZN(n4617) );
  OR2_X1 U5447 ( .A1(n5846), .A2(n6759), .ZN(n5867) );
  AOI21_X1 U5448 ( .B1(n7289), .B2(n4616), .A(n4615), .ZN(n4611) );
  INV_X1 U5449 ( .A(n6624), .ZN(n4616) );
  NAND2_X1 U5450 ( .A1(n7832), .A2(n4601), .ZN(n7919) );
  OR2_X1 U5451 ( .A1(n7254), .A2(n9680), .ZN(n7255) );
  INV_X1 U5452 ( .A(n5495), .ZN(n4505) );
  NOR2_X1 U5453 ( .A1(n4507), .A2(n4509), .ZN(n4502) );
  NOR2_X1 U5454 ( .A1(n5127), .A2(n4482), .ZN(n4481) );
  INV_X1 U5455 ( .A(n5105), .ZN(n4482) );
  AND2_X1 U5456 ( .A1(n5158), .A2(n5134), .ZN(n5156) );
  OR2_X1 U5457 ( .A1(n4333), .A2(n4684), .ZN(n4683) );
  INV_X1 U5458 ( .A(n5540), .ZN(n4684) );
  OR2_X1 U5459 ( .A1(n8113), .A2(n8115), .ZN(n5489) );
  NAND2_X1 U5460 ( .A1(n5141), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5169) );
  OAI21_X1 U5461 ( .B1(n4700), .B2(n4336), .A(n4450), .ZN(n7524) );
  NAND2_X1 U5462 ( .A1(n7524), .A2(n7525), .ZN(n7523) );
  AND2_X1 U5463 ( .A1(n5315), .A2(n5338), .ZN(n4701) );
  AND2_X1 U5464 ( .A1(n8365), .A2(n8346), .ZN(n6860) );
  INV_X1 U5465 ( .A(n8811), .ZN(n7203) );
  INV_X1 U5466 ( .A(n8615), .ZN(n8149) );
  INV_X1 U5467 ( .A(n8363), .ZN(n4703) );
  XNOR2_X1 U5468 ( .A(n8357), .B(n8569), .ZN(n4853) );
  AOI21_X1 U5469 ( .B1(n8355), .B2(n8354), .A(n8353), .ZN(n8357) );
  NAND2_X1 U5470 ( .A1(n4866), .A2(n4864), .ZN(n8355) );
  XNOR2_X1 U5471 ( .A(n4947), .B(n4539), .ZN(n9516) );
  AND2_X1 U5472 ( .A1(n4547), .A2(n6866), .ZN(n8415) );
  AND2_X1 U5473 ( .A1(n4549), .A2(n6869), .ZN(n8443) );
  OR2_X1 U5474 ( .A1(n5111), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n5184) );
  NAND2_X1 U5475 ( .A1(n8469), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n4541) );
  NOR2_X1 U5476 ( .A1(n7015), .A2(n4551), .ZN(n7019) );
  AND2_X1 U5477 ( .A1(n7016), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n4551) );
  NOR2_X1 U5478 ( .A1(n7018), .A2(n7019), .ZN(n7161) );
  NOR2_X1 U5479 ( .A1(n7161), .A2(n4550), .ZN(n8485) );
  AND2_X1 U5480 ( .A1(n7162), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n4550) );
  NAND2_X1 U5481 ( .A1(n8485), .A2(n8486), .ZN(n8484) );
  NAND2_X1 U5482 ( .A1(n8534), .A2(n4546), .ZN(n8537) );
  OR2_X1 U5483 ( .A1(n8535), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n4546) );
  NOR2_X1 U5484 ( .A1(n8537), .A2(n8536), .ZN(n8548) );
  NOR2_X1 U5485 ( .A1(n8548), .A2(n4545), .ZN(n8562) );
  AND2_X1 U5486 ( .A1(n8549), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n4545) );
  NAND2_X1 U5487 ( .A1(n4778), .A2(n4773), .ZN(n4772) );
  INV_X1 U5488 ( .A(n4777), .ZN(n4776) );
  OAI21_X1 U5489 ( .B1(n8589), .B2(n4781), .A(n8012), .ZN(n4777) );
  OR2_X1 U5490 ( .A1(n8847), .A2(n8601), .ZN(n8012) );
  NOR2_X1 U5491 ( .A1(n8589), .A2(n4779), .ZN(n4778) );
  INV_X1 U5492 ( .A(n8614), .ZN(n4775) );
  OAI21_X1 U5493 ( .B1(n8033), .B2(n8034), .A(n8349), .ZN(n4516) );
  AND2_X1 U5494 ( .A1(n4870), .A2(n8325), .ZN(n8033) );
  NAND2_X1 U5495 ( .A1(n4870), .A2(n4869), .ZN(n8349) );
  XNOR2_X1 U5496 ( .A(n8588), .B(n8194), .ZN(n4415) );
  NAND2_X1 U5497 ( .A1(n8615), .A2(n9743), .ZN(n4413) );
  INV_X1 U5498 ( .A(n8314), .ZN(n4848) );
  NAND2_X1 U5499 ( .A1(n8658), .A2(n4530), .ZN(n8607) );
  AOI21_X1 U5500 ( .B1(n4756), .B2(n4755), .A(n4763), .ZN(n4754) );
  NAND2_X1 U5501 ( .A1(n8311), .A2(n8312), .ZN(n8640) );
  NAND2_X1 U5502 ( .A1(n4394), .A2(n8028), .ZN(n8693) );
  INV_X1 U5503 ( .A(n8710), .ZN(n4394) );
  NAND2_X1 U5504 ( .A1(n8781), .A2(n4331), .ZN(n8706) );
  NAND2_X1 U5505 ( .A1(n8781), .A2(n4326), .ZN(n8721) );
  INV_X1 U5506 ( .A(n4877), .ZN(n4876) );
  AND2_X1 U5507 ( .A1(n8025), .A2(n4875), .ZN(n4874) );
  NAND2_X1 U5508 ( .A1(n8781), .A2(n4528), .ZN(n8729) );
  AND2_X1 U5509 ( .A1(n8781), .A2(n8750), .ZN(n8746) );
  NOR2_X1 U5510 ( .A1(n8282), .A2(n4769), .ZN(n4764) );
  NAND2_X1 U5511 ( .A1(n4536), .A2(n4330), .ZN(n8794) );
  NAND2_X1 U5512 ( .A1(n4536), .A2(n4535), .ZN(n8796) );
  NOR2_X1 U5513 ( .A1(n7645), .A2(n4537), .ZN(n7737) );
  NAND2_X1 U5514 ( .A1(n5188), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5235) );
  INV_X1 U5515 ( .A(n5189), .ZN(n5188) );
  OR3_X1 U5516 ( .A1(n5235), .A2(n5234), .A3(n7167), .ZN(n5257) );
  NOR2_X1 U5517 ( .A1(n7645), .A2(n7691), .ZN(n7735) );
  NAND2_X1 U5518 ( .A1(n7665), .A2(n9817), .ZN(n7804) );
  INV_X1 U5519 ( .A(n8376), .ZN(n7456) );
  NAND2_X1 U5520 ( .A1(n4401), .A2(n4404), .ZN(n4400) );
  OAI21_X1 U5521 ( .B1(n7276), .B2(n4404), .A(n4401), .ZN(n7654) );
  INV_X1 U5522 ( .A(n8377), .ZN(n7656) );
  NAND2_X1 U5523 ( .A1(n7205), .A2(n4404), .ZN(n7658) );
  NAND2_X1 U5524 ( .A1(n7276), .A2(n8246), .ZN(n7213) );
  NAND2_X1 U5525 ( .A1(n7213), .A2(n8247), .ZN(n7454) );
  AND2_X1 U5526 ( .A1(n8241), .A2(n8246), .ZN(n8239) );
  NAND2_X1 U5527 ( .A1(n8214), .A2(n8207), .ZN(n8180) );
  NAND2_X1 U5528 ( .A1(n9753), .A2(n4397), .ZN(n4395) );
  INV_X1 U5529 ( .A(n4397), .ZN(n4396) );
  NAND2_X1 U5530 ( .A1(n9742), .A2(n8212), .ZN(n7211) );
  NAND2_X1 U5531 ( .A1(n4854), .A2(n8220), .ZN(n9742) );
  NOR2_X1 U5532 ( .A1(n8826), .A2(n9770), .ZN(n7352) );
  AND2_X1 U5533 ( .A1(n4759), .A2(n4756), .ZN(n8878) );
  INV_X1 U5534 ( .A(n7355), .ZN(n9776) );
  OR2_X1 U5535 ( .A1(n5615), .A2(P2_U3152), .ZN(n9759) );
  NOR2_X1 U5536 ( .A1(n4885), .A2(P2_IR_REG_25__SCAN_IN), .ZN(n4521) );
  NAND2_X1 U5537 ( .A1(n4912), .A2(n4887), .ZN(n4885) );
  XNOR2_X1 U5538 ( .A(n5593), .B(n4906), .ZN(n6540) );
  NAND2_X1 U5539 ( .A1(n4931), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4933) );
  OR2_X1 U5540 ( .A1(n7859), .A2(n7858), .ZN(n4440) );
  OR2_X1 U5541 ( .A1(n6113), .A2(n8989), .ZN(n6133) );
  OR2_X1 U5542 ( .A1(n6133), .A2(n9044), .ZN(n6150) );
  NAND2_X1 U5543 ( .A1(n6148), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n6168) );
  INV_X1 U5544 ( .A(n6150), .ZN(n6148) );
  NAND2_X1 U5545 ( .A1(n5690), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n6007) );
  INV_X1 U5546 ( .A(n5980), .ZN(n5690) );
  OR2_X1 U5547 ( .A1(n6007), .A2(n6006), .ZN(n6025) );
  NAND2_X1 U5548 ( .A1(n5692), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n6078) );
  INV_X1 U5549 ( .A(n6061), .ZN(n5692) );
  OR2_X1 U5550 ( .A1(n6078), .A2(n9054), .ZN(n6093) );
  AOI21_X1 U5551 ( .B1(n4674), .B2(n7746), .A(n4357), .ZN(n4673) );
  NAND2_X1 U5552 ( .A1(n5694), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n6113) );
  INV_X1 U5553 ( .A(n6111), .ZN(n5694) );
  NAND2_X1 U5554 ( .A1(n4428), .A2(n4426), .ZN(n9061) );
  AOI21_X1 U5555 ( .B1(n4429), .B2(n4431), .A(n4427), .ZN(n4426) );
  NAND2_X1 U5556 ( .A1(n4423), .A2(n6056), .ZN(n9077) );
  INV_X1 U5557 ( .A(n6054), .ZN(n4423) );
  NAND2_X1 U5558 ( .A1(n6054), .A2(n6055), .ZN(n9076) );
  NAND2_X1 U5559 ( .A1(n5691), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n6043) );
  INV_X1 U5560 ( .A(n6025), .ZN(n5691) );
  OR2_X1 U5561 ( .A1(n6043), .A2(n6042), .ZN(n6061) );
  NAND2_X1 U5562 ( .A1(n5791), .A2(n7080), .ZN(n7434) );
  INV_X1 U5563 ( .A(n6768), .ZN(n6841) );
  NAND2_X1 U5564 ( .A1(n4669), .A2(n6144), .ZN(n4668) );
  INV_X1 U5565 ( .A(n6145), .ZN(n4669) );
  NAND2_X1 U5566 ( .A1(n4659), .A2(n4658), .ZN(n4670) );
  INV_X1 U5567 ( .A(n9042), .ZN(n4658) );
  NOR2_X1 U5568 ( .A1(n6003), .A2(n4792), .ZN(n5651) );
  NAND2_X1 U5569 ( .A1(n4741), .A2(n4740), .ZN(n4739) );
  INV_X1 U5570 ( .A(n6484), .ZN(n4740) );
  NAND2_X1 U5571 ( .A1(n6486), .A2(n6631), .ZN(n4741) );
  OR2_X1 U5572 ( .A1(n9193), .A2(n6367), .ZN(n6487) );
  AND3_X1 U5573 ( .A1(n6098), .A2(n6097), .A3(n6096), .ZN(n9055) );
  INV_X1 U5574 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5836) );
  NAND2_X1 U5575 ( .A1(n6292), .A2(n6291), .ZN(n9198) );
  INV_X1 U5576 ( .A(n4597), .ZN(n9199) );
  INV_X1 U5577 ( .A(n4825), .ZN(n4822) );
  INV_X1 U5578 ( .A(n4823), .ZN(n4821) );
  AND2_X1 U5579 ( .A1(n4596), .A2(n4828), .ZN(n4595) );
  AND2_X1 U5580 ( .A1(n6205), .A2(n6243), .ZN(n9216) );
  NAND2_X1 U5581 ( .A1(n7976), .A2(n7975), .ZN(n9229) );
  NAND2_X1 U5582 ( .A1(n9244), .A2(n6441), .ZN(n9263) );
  NAND2_X1 U5583 ( .A1(n4623), .A2(n4621), .ZN(n9273) );
  AOI21_X1 U5584 ( .B1(n4625), .B2(n4624), .A(n4622), .ZN(n4621) );
  NOR2_X1 U5585 ( .A1(n9344), .A2(n4606), .ZN(n9312) );
  NAND2_X1 U5586 ( .A1(n4627), .A2(n7967), .ZN(n9327) );
  OR2_X1 U5587 ( .A1(n9350), .A2(n7968), .ZN(n4627) );
  OR2_X1 U5588 ( .A1(n6448), .A2(n7968), .ZN(n9351) );
  AOI21_X1 U5589 ( .B1(n4800), .B2(n4799), .A(n4379), .ZN(n4798) );
  NAND2_X1 U5590 ( .A1(n7832), .A2(n4327), .ZN(n9392) );
  AND2_X1 U5591 ( .A1(n9379), .A2(n6421), .ZN(n9399) );
  AND2_X1 U5592 ( .A1(n7832), .A2(n7835), .ZN(n7882) );
  AND2_X1 U5593 ( .A1(n6350), .A2(n7838), .ZN(n7836) );
  NAND2_X1 U5594 ( .A1(n5688), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5929) );
  INV_X1 U5595 ( .A(n5904), .ZN(n5688) );
  NAND2_X1 U5596 ( .A1(n7759), .A2(n7758), .ZN(n7779) );
  NAND2_X1 U5597 ( .A1(n5883), .A2(n5882), .ZN(n7685) );
  NOR2_X1 U5598 ( .A1(n7505), .A2(n7685), .ZN(n7626) );
  INV_X1 U5599 ( .A(n4805), .ZN(n4804) );
  OAI22_X1 U5600 ( .A1(n4338), .A2(n4806), .B1(n7520), .B2(n9125), .ZN(n4805)
         );
  NAND2_X1 U5601 ( .A1(n4362), .A2(n7364), .ZN(n4806) );
  NAND2_X1 U5602 ( .A1(n5687), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n5885) );
  INV_X1 U5603 ( .A(n5867), .ZN(n5687) );
  OR2_X1 U5604 ( .A1(n7375), .A2(n7520), .ZN(n7505) );
  NAND2_X1 U5605 ( .A1(n7369), .A2(n7368), .ZN(n7498) );
  NAND2_X1 U5606 ( .A1(n5685), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5830) );
  NAND2_X1 U5607 ( .A1(n5686), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5846) );
  INV_X1 U5608 ( .A(n5830), .ZN(n5686) );
  NAND2_X1 U5609 ( .A1(n7299), .A2(n7298), .ZN(n7388) );
  AND2_X1 U5610 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n5792) );
  AND2_X1 U5611 ( .A1(n6624), .A2(n6623), .ZN(n7251) );
  NAND2_X1 U5612 ( .A1(n4610), .A2(n7116), .ZN(n4609) );
  INV_X1 U5613 ( .A(n7144), .ZN(n7173) );
  NAND2_X1 U5614 ( .A1(n6377), .A2(n6496), .ZN(n7115) );
  AND4_X2 U5615 ( .A1(n5749), .A2(n5748), .A3(n5747), .A4(n5746), .ZN(n6309)
         );
  OR2_X1 U5616 ( .A1(n5744), .A2(n6973), .ZN(n5747) );
  NAND2_X1 U5617 ( .A1(n6932), .A2(n5684), .ZN(n6642) );
  AND2_X1 U5618 ( .A1(n6631), .A2(n6527), .ZN(n6768) );
  AND2_X1 U5619 ( .A1(n7248), .A2(n7247), .ZN(n9561) );
  OR2_X1 U5620 ( .A1(n6471), .A2(n6615), .ZN(n7247) );
  INV_X1 U5621 ( .A(n9559), .ZN(n9707) );
  OAI21_X1 U5622 ( .B1(n6289), .B2(n6288), .A(n6277), .ZN(n6280) );
  XNOR2_X1 U5623 ( .A(n6301), .B(n6300), .ZN(n8013) );
  XNOR2_X1 U5624 ( .A(n6267), .B(n6266), .ZN(n7926) );
  XNOR2_X1 U5625 ( .A(n5604), .B(n5603), .ZN(n7891) );
  XNOR2_X1 U5626 ( .A(n5542), .B(n5541), .ZN(n7888) );
  OR2_X1 U5627 ( .A1(n6003), .A2(n4794), .ZN(n5658) );
  NAND2_X1 U5628 ( .A1(n4735), .A2(n5365), .ZN(n5383) );
  OAI21_X1 U5629 ( .B1(n5272), .B2(n4498), .A(n4496), .ZN(n5363) );
  NAND2_X1 U5630 ( .A1(n4501), .A2(n4706), .ZN(n5344) );
  NAND2_X1 U5631 ( .A1(n5272), .A2(n4709), .ZN(n4501) );
  NAND2_X1 U5632 ( .A1(n4708), .A2(n4714), .ZN(n5318) );
  NAND2_X1 U5633 ( .A1(n5272), .A2(n4716), .ZN(n4708) );
  NAND2_X1 U5634 ( .A1(n4713), .A2(n5270), .ZN(n5301) );
  OR2_X1 U5635 ( .A1(n5272), .A2(n5271), .ZN(n4713) );
  INV_X1 U5636 ( .A(n5636), .ZN(n4789) );
  NAND2_X1 U5637 ( .A1(n4489), .A2(n5201), .ZN(n5224) );
  NAND2_X1 U5638 ( .A1(n5180), .A2(n4490), .ZN(n4489) );
  NAND2_X1 U5639 ( .A1(n5180), .A2(n5179), .ZN(n5203) );
  NAND2_X1 U5640 ( .A1(n5106), .A2(n5105), .ZN(n5128) );
  NAND2_X1 U5641 ( .A1(n5080), .A2(n4719), .ZN(n4718) );
  AND2_X1 U5642 ( .A1(n5805), .A2(n4791), .ZN(n6590) );
  NAND2_X1 U5643 ( .A1(n5633), .A2(n5632), .ZN(n5802) );
  NAND2_X1 U5644 ( .A1(n4994), .A2(n4944), .ZN(n5717) );
  NAND2_X1 U5645 ( .A1(n7713), .A2(n5246), .ZN(n7815) );
  NAND2_X1 U5646 ( .A1(n7240), .A2(n5155), .ZN(n7344) );
  NAND2_X1 U5647 ( .A1(n8138), .A2(n5361), .ZN(n8065) );
  OAI21_X1 U5648 ( .B1(n8847), .B2(n4696), .A(n4691), .ZN(n4690) );
  NAND2_X1 U5649 ( .A1(n5612), .A2(n4696), .ZN(n4691) );
  INV_X1 U5650 ( .A(n4693), .ZN(n4692) );
  OAI21_X1 U5651 ( .B1(n8847), .B2(n5573), .A(n4694), .ZN(n4693) );
  NAND2_X1 U5652 ( .A1(n5612), .A2(n5573), .ZN(n4694) );
  AOI22_X1 U5653 ( .A1(n5612), .A2(n5614), .B1(n5613), .B2(n5614), .ZN(n4695)
         );
  NAND2_X1 U5654 ( .A1(n7523), .A2(n7527), .ZN(n7582) );
  NAND2_X1 U5655 ( .A1(n5316), .A2(n5315), .ZN(n8106) );
  OR2_X1 U5656 ( .A1(n6974), .A2(n6977), .ZN(n6975) );
  NAND2_X1 U5657 ( .A1(n4700), .A2(n5126), .ZN(n7239) );
  NAND2_X1 U5658 ( .A1(n8063), .A2(n5382), .ZN(n8120) );
  AOI21_X1 U5659 ( .B1(n4678), .B2(n4681), .A(n4676), .ZN(n4675) );
  NAND2_X1 U5660 ( .A1(n4449), .A2(n4345), .ZN(n4677) );
  INV_X1 U5661 ( .A(n7581), .ZN(n4676) );
  XNOR2_X1 U5662 ( .A(n5445), .B(n5443), .ZN(n8129) );
  INV_X1 U5663 ( .A(n8124), .ZN(n8160) );
  NAND2_X1 U5664 ( .A1(n4686), .A2(n8082), .ZN(n8147) );
  INV_X1 U5665 ( .A(n8368), .ZN(n4850) );
  NAND2_X1 U5666 ( .A1(n5535), .A2(n5534), .ZN(n8630) );
  OR2_X1 U5667 ( .A1(n8609), .A2(n5627), .ZN(n5535) );
  INV_X1 U5668 ( .A(n4547), .ZN(n8400) );
  INV_X1 U5669 ( .A(n4549), .ZN(n8428) );
  INV_X1 U5670 ( .A(n4544), .ZN(n8456) );
  INV_X1 U5671 ( .A(n4542), .ZN(n8470) );
  OAI22_X1 U5672 ( .A1(n9509), .A2(n4987), .B1(n5063), .B2(n8170), .ZN(n8835)
         );
  XNOR2_X1 U5673 ( .A(n8835), .B(n8576), .ZN(n8837) );
  AND2_X1 U5674 ( .A1(n8174), .A2(n8173), .ZN(n8578) );
  NAND2_X1 U5675 ( .A1(n4845), .A2(n8314), .ZN(n8613) );
  NAND2_X1 U5676 ( .A1(n8629), .A2(n8620), .ZN(n4845) );
  NAND2_X1 U5677 ( .A1(n8658), .A2(n8009), .ZN(n8623) );
  NAND2_X1 U5678 ( .A1(n4759), .A2(n4760), .ZN(n8656) );
  AND2_X1 U5679 ( .A1(n8675), .A2(n8292), .ZN(n4894) );
  AOI21_X1 U5680 ( .B1(n4316), .B2(n8008), .A(n4325), .ZN(n8668) );
  NAND2_X1 U5681 ( .A1(n8772), .A2(n8285), .ZN(n8752) );
  INV_X1 U5682 ( .A(n4766), .ZN(n8767) );
  NAND2_X1 U5683 ( .A1(n8791), .A2(n8002), .ZN(n8766) );
  NAND2_X1 U5684 ( .A1(n8023), .A2(n8272), .ZN(n8800) );
  NAND2_X1 U5685 ( .A1(n7721), .A2(n7695), .ZN(n7998) );
  NOR2_X1 U5686 ( .A1(n7400), .A2(n4389), .ZN(n9787) );
  NAND2_X1 U5687 ( .A1(n8217), .A2(n8224), .ZN(n7357) );
  INV_X1 U5688 ( .A(n7668), .ZN(n9747) );
  NAND2_X1 U5689 ( .A1(n8845), .A2(n4511), .ZN(n8942) );
  INV_X1 U5690 ( .A(n4512), .ZN(n4511) );
  OAI21_X1 U5691 ( .B1(n8846), .B2(n9797), .A(n8844), .ZN(n4512) );
  NAND2_X1 U5692 ( .A1(n4913), .A2(n8962), .ZN(n4585) );
  OR2_X1 U5693 ( .A1(n4937), .A2(n4586), .ZN(n4584) );
  NAND2_X1 U5694 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_29__SCAN_IN), 
        .ZN(n4586) );
  NAND2_X1 U5695 ( .A1(n4523), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4522) );
  NAND2_X1 U5696 ( .A1(n4930), .A2(n4926), .ZN(n4927) );
  INV_X1 U5697 ( .A(n8199), .ZN(n8343) );
  AND2_X1 U5698 ( .A1(n5041), .A2(n5040), .ZN(n8413) );
  OR3_X1 U5699 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .A3(
        P2_IR_REG_0__SCAN_IN), .ZN(n4997) );
  AND2_X1 U5700 ( .A1(P2_U3152), .A2(n4994), .ZN(n8969) );
  NAND2_X1 U5701 ( .A1(n4742), .A2(n4958), .ZN(n4959) );
  NAND2_X1 U5702 ( .A1(n5655), .A2(SI_0_), .ZN(n4742) );
  NAND2_X1 U5703 ( .A1(n4672), .A2(n5828), .ZN(n7483) );
  INV_X1 U5704 ( .A(n9075), .ZN(n4424) );
  NOR2_X1 U5705 ( .A1(n6056), .A2(n9075), .ZN(n4425) );
  NAND2_X1 U5706 ( .A1(n7481), .A2(n4337), .ZN(n7534) );
  NAND2_X1 U5707 ( .A1(n4420), .A2(n5857), .ZN(n7533) );
  NAND2_X1 U5708 ( .A1(n7481), .A2(n5845), .ZN(n4420) );
  NAND2_X1 U5709 ( .A1(n9050), .A2(n6086), .ZN(n4651) );
  NAND2_X1 U5710 ( .A1(n4670), .A2(n4668), .ZN(n9012) );
  NAND2_X1 U5711 ( .A1(n6147), .A2(n6146), .ZN(n9429) );
  AND4_X1 U5712 ( .A1(n6048), .A2(n6047), .A3(n6046), .A4(n6045), .ZN(n9037)
         );
  AND2_X1 U5713 ( .A1(n4652), .A2(n4653), .ZN(n9033) );
  INV_X1 U5714 ( .A(n4659), .ZN(n9041) );
  AND4_X1 U5715 ( .A1(n5890), .A2(n5889), .A3(n5888), .A4(n5887), .ZN(n7620)
         );
  NAND2_X1 U5716 ( .A1(n4421), .A2(n5858), .ZN(n4418) );
  INV_X1 U5717 ( .A(n9115), .ZN(n9087) );
  NAND2_X1 U5718 ( .A1(n6077), .A2(n6076), .ZN(n9455) );
  NAND2_X1 U5719 ( .A1(n4441), .A2(n4673), .ZN(n7861) );
  AND4_X1 U5720 ( .A1(n5934), .A2(n5933), .A3(n5932), .A4(n5931), .ZN(n7787)
         );
  INV_X1 U5721 ( .A(n9092), .ZN(n9104) );
  NAND2_X1 U5722 ( .A1(n9076), .A2(n9075), .ZN(n9080) );
  NAND2_X1 U5723 ( .A1(n6252), .A2(n6236), .ZN(n9115) );
  AND4_X1 U5724 ( .A1(n6012), .A2(n6011), .A3(n6010), .A4(n6009), .ZN(n9110)
         );
  NAND2_X1 U5725 ( .A1(n6242), .A2(n9692), .ZN(n9112) );
  NOR2_X1 U5726 ( .A1(n6534), .A2(n6533), .ZN(n6537) );
  INV_X1 U5727 ( .A(n9278), .ZN(n9248) );
  INV_X1 U5728 ( .A(n7134), .ZN(n9131) );
  INV_X1 U5729 ( .A(n9198), .ZN(n9556) );
  AND2_X1 U5730 ( .A1(n9206), .A2(n9205), .ZN(n9416) );
  NAND2_X1 U5731 ( .A1(n4829), .A2(n4825), .ZN(n9206) );
  NAND2_X1 U5732 ( .A1(n4829), .A2(n4827), .ZN(n9204) );
  NAND2_X1 U5733 ( .A1(n4830), .A2(n7957), .ZN(n9222) );
  INV_X1 U5734 ( .A(n9682), .ZN(n9282) );
  NAND2_X1 U5735 ( .A1(n6132), .A2(n6131), .ZN(n9436) );
  AOI21_X1 U5736 ( .B1(n4841), .B2(n4839), .A(n4837), .ZN(n4833) );
  NAND2_X1 U5737 ( .A1(n4620), .A2(n4624), .ZN(n9289) );
  OR2_X1 U5738 ( .A1(n9350), .A2(n4625), .ZN(n4620) );
  NAND2_X1 U5739 ( .A1(n4841), .A2(n7951), .ZN(n9287) );
  NAND2_X1 U5740 ( .A1(n7950), .A2(n7949), .ZN(n9301) );
  NAND2_X1 U5741 ( .A1(n6091), .A2(n6090), .ZN(n9452) );
  NAND2_X1 U5742 ( .A1(n4803), .A2(n7945), .ZN(n9357) );
  NAND2_X1 U5743 ( .A1(n9374), .A2(n9381), .ZN(n4803) );
  NAND2_X1 U5744 ( .A1(n4807), .A2(n4808), .ZN(n7914) );
  INV_X1 U5745 ( .A(n7913), .ZN(n4818) );
  NAND2_X1 U5746 ( .A1(n4813), .A2(n4810), .ZN(n7912) );
  INV_X1 U5747 ( .A(n4814), .ZN(n4810) );
  NAND2_X1 U5748 ( .A1(n7831), .A2(n4816), .ZN(n4813) );
  OAI21_X1 U5749 ( .B1(n7831), .B2(n7830), .A(n7829), .ZN(n7879) );
  NAND2_X1 U5750 ( .A1(n5945), .A2(n5944), .ZN(n7868) );
  NAND2_X1 U5751 ( .A1(n4786), .A2(n7757), .ZN(n7786) );
  OR2_X1 U5752 ( .A1(n7755), .A2(n7756), .ZN(n4786) );
  NAND2_X1 U5753 ( .A1(n7365), .A2(n7364), .ZN(n7496) );
  NAND2_X1 U5754 ( .A1(n7290), .A2(n7289), .ZN(n7383) );
  NAND2_X1 U5755 ( .A1(n7249), .A2(n6626), .ZN(n6628) );
  OR2_X1 U5756 ( .A1(n5838), .A2(n6665), .ZN(n5734) );
  AND2_X1 U5757 ( .A1(n6543), .A2(n6235), .ZN(n9697) );
  INV_X1 U5758 ( .A(n8169), .ZN(n9509) );
  NAND2_X1 U5759 ( .A1(n5700), .A2(n5699), .ZN(n5702) );
  NAND2_X1 U5760 ( .A1(n5696), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5699) );
  NAND2_X1 U5761 ( .A1(n5678), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5679) );
  NAND2_X1 U5762 ( .A1(n4721), .A2(n5062), .ZN(n5081) );
  NAND2_X1 U5763 ( .A1(n5060), .A2(n5059), .ZN(n4721) );
  INV_X1 U5764 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n10041) );
  XNOR2_X1 U5765 ( .A(n5060), .B(n5059), .ZN(n6653) );
  NOR2_X1 U5766 ( .A1(n7571), .A2(n10080), .ZN(n9876) );
  OAI21_X1 U5767 ( .B1(n4456), .B2(n5614), .A(n4386), .ZN(P2_U3231) );
  XNOR2_X1 U5768 ( .A(n8114), .B(n4457), .ZN(n4456) );
  OR2_X1 U5769 ( .A1(n8367), .A2(n8366), .ZN(n4849) );
  NAND2_X1 U5770 ( .A1(n4559), .A2(n4552), .ZN(P2_U3264) );
  NAND2_X1 U5771 ( .A1(n8570), .A2(n8569), .ZN(n4559) );
  AOI21_X1 U5772 ( .B1(n4556), .B2(n8356), .A(n4553), .ZN(n4552) );
  NOR2_X1 U5773 ( .A1(n8850), .A2(n8804), .ZN(n8591) );
  NAND2_X1 U5774 ( .A1(n4443), .A2(n4442), .ZN(n9096) );
  OAI21_X1 U5775 ( .B1(n7994), .B2(n6638), .A(n4634), .ZN(P1_U3355) );
  AOI211_X1 U5776 ( .C1(n7996), .C2(n9409), .A(n4635), .B(n7995), .ZN(n4634)
         );
  NOR2_X1 U5777 ( .A1(n7997), .A2(n9411), .ZN(n4635) );
  OR2_X2 U5778 ( .A1(n5584), .A2(n4883), .ZN(n4324) );
  NAND2_X1 U5779 ( .A1(n7950), .A2(n4842), .ZN(n4841) );
  AND2_X1 U5780 ( .A1(n8692), .A2(n8681), .ZN(n4325) );
  INV_X1 U5781 ( .A(n8655), .ZN(n4758) );
  AND2_X1 U5782 ( .A1(n6875), .A2(n4994), .ZN(n4996) );
  AND2_X1 U5783 ( .A1(n4528), .A2(n4527), .ZN(n4326) );
  AND2_X1 U5784 ( .A1(n4601), .A2(n4600), .ZN(n4327) );
  INV_X1 U5785 ( .A(n9210), .ZN(n9249) );
  AND2_X1 U5786 ( .A1(n6192), .A2(n6191), .ZN(n9210) );
  AND2_X1 U5787 ( .A1(n8325), .A2(n8329), .ZN(n8589) );
  NAND2_X1 U5788 ( .A1(n5633), .A2(n4790), .ZN(n4791) );
  AND2_X1 U5789 ( .A1(n4673), .A2(n4353), .ZN(n4328) );
  NAND2_X1 U5790 ( .A1(n5959), .A2(n5958), .ZN(n9476) );
  OR2_X1 U5791 ( .A1(n5016), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n4329) );
  AND2_X1 U5792 ( .A1(n4538), .A2(n4535), .ZN(n4330) );
  AND2_X1 U5793 ( .A1(n4326), .A2(n4526), .ZN(n4331) );
  NAND2_X1 U5794 ( .A1(n8810), .A2(n7403), .ZN(n8207) );
  AND2_X1 U5795 ( .A1(n8212), .A2(n8213), .ZN(n4332) );
  INV_X2 U5796 ( .A(n4994), .ZN(n5655) );
  AND2_X1 U5797 ( .A1(n8655), .A2(n8292), .ZN(n4882) );
  NAND3_X1 U5798 ( .A1(n4979), .A2(n4978), .A3(n4977), .ZN(n7029) );
  NOR2_X1 U5799 ( .A1(n8148), .A2(n4685), .ZN(n4333) );
  AND2_X1 U5800 ( .A1(n4327), .A2(n4599), .ZN(n4334) );
  XNOR2_X1 U5801 ( .A(n5679), .B(n5643), .ZN(n6241) );
  NAND2_X1 U5802 ( .A1(n7747), .A2(n4674), .ZN(n7848) );
  NAND2_X1 U5803 ( .A1(n5915), .A2(n5914), .ZN(n7747) );
  AND2_X4 U5804 ( .A1(n7937), .A2(n5703), .ZN(n4335) );
  INV_X1 U5805 ( .A(n5213), .ZN(n5418) );
  XNOR2_X1 U5806 ( .A(n4946), .B(n4540), .ZN(n4947) );
  INV_X1 U5807 ( .A(n5745), .ZN(n5796) );
  INV_X2 U5808 ( .A(n5796), .ZN(n6283) );
  OR2_X1 U5809 ( .A1(n7343), .A2(n4452), .ZN(n4336) );
  NAND2_X1 U5810 ( .A1(n4911), .A2(n4521), .ZN(n4941) );
  OR2_X1 U5811 ( .A1(n8858), .A2(n8087), .ZN(n8319) );
  AND2_X1 U5812 ( .A1(n5845), .A2(n5858), .ZN(n4337) );
  AND2_X1 U5813 ( .A1(n7302), .A2(n7301), .ZN(n4338) );
  NAND2_X1 U5814 ( .A1(n5657), .A2(n5656), .ZN(n9441) );
  AND2_X1 U5815 ( .A1(n7849), .A2(n5920), .ZN(n4674) );
  AND2_X1 U5816 ( .A1(n8267), .A2(n8266), .ZN(n8188) );
  INV_X1 U5817 ( .A(n8247), .ZN(n4404) );
  OAI211_X1 U5818 ( .C1(n4987), .C2(n6662), .A(n5019), .B(n5018), .ZN(n7045)
         );
  NAND2_X1 U5819 ( .A1(n9436), .A2(n9265), .ZN(n4339) );
  NAND2_X1 U5820 ( .A1(n7937), .A2(n7930), .ZN(n5744) );
  AND2_X1 U5821 ( .A1(n8272), .A2(n8273), .ZN(n8269) );
  NAND4_X2 U5822 ( .A1(n5729), .A2(n5728), .A3(n5731), .A4(n5730), .ZN(n9133)
         );
  INV_X1 U5823 ( .A(n4974), .ZN(n5624) );
  AND2_X1 U5824 ( .A1(n4682), .A2(n4683), .ZN(n8045) );
  INV_X1 U5825 ( .A(n8242), .ZN(n4402) );
  NAND2_X1 U5826 ( .A1(n4651), .A2(n6089), .ZN(n9004) );
  INV_X1 U5827 ( .A(n4833), .ZN(n9270) );
  OR2_X1 U5828 ( .A1(n8236), .A2(n8338), .ZN(n4340) );
  NOR2_X1 U5829 ( .A1(n6330), .A2(n6366), .ZN(n7979) );
  NAND2_X1 U5830 ( .A1(n9239), .A2(n4595), .ZN(n4341) );
  NAND2_X2 U5831 ( .A1(n6543), .A2(n5677), .ZN(n6209) );
  INV_X1 U5832 ( .A(n7029), .ZN(n7030) );
  INV_X4 U5833 ( .A(n5838), .ZN(n5751) );
  NAND2_X1 U5834 ( .A1(n5550), .A2(n5549), .ZN(n8852) );
  INV_X1 U5835 ( .A(n8852), .ZN(n4529) );
  NAND2_X1 U5836 ( .A1(n6109), .A2(n6108), .ZN(n9317) );
  OR2_X1 U5837 ( .A1(n8847), .A2(n8048), .ZN(n8325) );
  OR2_X1 U5838 ( .A1(n8306), .A2(n8338), .ZN(n4342) );
  AND2_X1 U5839 ( .A1(n4542), .A2(n4541), .ZN(n4343) );
  AND2_X1 U5840 ( .A1(n7977), .A2(n6372), .ZN(n7959) );
  NAND2_X1 U5841 ( .A1(n8321), .A2(n8327), .ZN(n8599) );
  INV_X1 U5842 ( .A(n8599), .ZN(n4779) );
  AND2_X1 U5843 ( .A1(n4808), .A2(n4818), .ZN(n4344) );
  AND2_X1 U5844 ( .A1(n4678), .A2(n4448), .ZN(n4345) );
  AND2_X1 U5845 ( .A1(n9233), .A2(n4632), .ZN(n4346) );
  AND2_X1 U5846 ( .A1(n5898), .A2(n5897), .ZN(n4347) );
  INV_X1 U5847 ( .A(n4602), .ZN(n9292) );
  NOR3_X1 U5848 ( .A1(n9344), .A2(n9441), .A3(n4606), .ZN(n4602) );
  AND2_X1 U5849 ( .A1(n4530), .A2(n4529), .ZN(n4348) );
  NAND2_X1 U5850 ( .A1(n5526), .A2(n5525), .ZN(n8858) );
  NAND2_X1 U5851 ( .A1(n5255), .A2(n5254), .ZN(n8925) );
  NAND2_X1 U5852 ( .A1(n5978), .A2(n5977), .ZN(n9113) );
  NOR2_X1 U5853 ( .A1(n9344), .A2(n4603), .ZN(n4607) );
  AND2_X1 U5854 ( .A1(n9020), .A2(n9034), .ZN(n4349) );
  AND2_X1 U5855 ( .A1(n5263), .A2(n5246), .ZN(n4350) );
  AND2_X1 U5856 ( .A1(n5379), .A2(n5361), .ZN(n4351) );
  INV_X1 U5857 ( .A(n8867), .ZN(n8009) );
  NAND2_X1 U5858 ( .A1(n5468), .A2(n5467), .ZN(n8867) );
  AND2_X1 U5859 ( .A1(n4743), .A2(n7635), .ZN(n4352) );
  NAND2_X1 U5860 ( .A1(n7859), .A2(n7858), .ZN(n4353) );
  NOR2_X1 U5861 ( .A1(n4794), .A2(n4889), .ZN(n4793) );
  AND2_X1 U5862 ( .A1(n8310), .A2(n4461), .ZN(n4354) );
  INV_X1 U5863 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n4925) );
  INV_X1 U5864 ( .A(n8262), .ZN(n4409) );
  AND2_X1 U5865 ( .A1(n4653), .A2(n6038), .ZN(n4355) );
  AND2_X1 U5866 ( .A1(n7382), .A2(n6380), .ZN(n6627) );
  AND2_X1 U5867 ( .A1(n8250), .A2(n8206), .ZN(n8182) );
  NAND2_X1 U5868 ( .A1(n4628), .A2(n7967), .ZN(n4356) );
  INV_X1 U5869 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n4887) );
  AND2_X1 U5870 ( .A1(n5941), .A2(n5940), .ZN(n4357) );
  INV_X1 U5871 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n4705) );
  AOI21_X1 U5872 ( .B1(n5668), .B2(P1_IR_REG_31__SCAN_IN), .A(n4647), .ZN(
        n4646) );
  AND2_X1 U5873 ( .A1(n8209), .A2(n8208), .ZN(n4358) );
  AND2_X1 U5874 ( .A1(n6104), .A2(n6105), .ZN(n9005) );
  AND2_X1 U5875 ( .A1(n9133), .A2(n7234), .ZN(n4359) );
  NAND2_X1 U5876 ( .A1(n7198), .A2(n9794), .ZN(n8214) );
  INV_X1 U5877 ( .A(n4801), .ZN(n4800) );
  OR2_X1 U5878 ( .A1(n7946), .A2(n4802), .ZN(n4801) );
  INV_X1 U5879 ( .A(n4769), .ZN(n4765) );
  INV_X1 U5880 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n4910) );
  NOR2_X1 U5881 ( .A1(n8879), .A2(n8699), .ZN(n4360) );
  NAND2_X1 U5882 ( .A1(n6201), .A2(n6200), .ZN(n9214) );
  INV_X1 U5883 ( .A(n9214), .ZN(n4596) );
  AND2_X1 U5884 ( .A1(n9214), .A2(n7960), .ZN(n4361) );
  NAND2_X1 U5885 ( .A1(n9745), .A2(n9788), .ZN(n8209) );
  INV_X1 U5886 ( .A(n4843), .ZN(n4842) );
  OR2_X1 U5887 ( .A1(n7952), .A2(n4844), .ZN(n4843) );
  INV_X1 U5888 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n4899) );
  NAND2_X1 U5889 ( .A1(n6186), .A2(n6185), .ZN(n9420) );
  INV_X1 U5890 ( .A(n9420), .ZN(n4828) );
  INV_X1 U5891 ( .A(n4781), .ZN(n4780) );
  NAND2_X1 U5892 ( .A1(n4529), .A2(n8149), .ZN(n4781) );
  NAND2_X1 U5893 ( .A1(n7520), .A2(n9125), .ZN(n4362) );
  OAI21_X1 U5894 ( .B1(n8578), .B2(n8350), .A(n8348), .ZN(n4873) );
  AND2_X1 U5895 ( .A1(n8301), .A2(n8299), .ZN(n4363) );
  NAND2_X1 U5896 ( .A1(n8302), .A2(n8322), .ZN(n4364) );
  NAND2_X1 U5897 ( .A1(n4583), .A2(n8295), .ZN(n4365) );
  INV_X1 U5898 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n6233) );
  NAND2_X1 U5899 ( .A1(n8333), .A2(n8348), .ZN(n8330) );
  NOR2_X1 U5900 ( .A1(n9113), .A2(n9119), .ZN(n4366) );
  XNOR2_X1 U5901 ( .A(n8873), .B(n8645), .ZN(n8655) );
  NAND2_X1 U5902 ( .A1(n7895), .A2(n5989), .ZN(n4367) );
  AND2_X1 U5903 ( .A1(n4683), .A2(n8046), .ZN(n4368) );
  AND2_X1 U5904 ( .A1(n8249), .A2(n8242), .ZN(n8247) );
  AND2_X1 U5905 ( .A1(n6374), .A2(n7978), .ZN(n9203) );
  INV_X1 U5906 ( .A(n9203), .ZN(n4826) );
  AND2_X1 U5907 ( .A1(n5703), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n4369) );
  AND2_X1 U5908 ( .A1(n7699), .A2(n7695), .ZN(n4370) );
  AND2_X1 U5909 ( .A1(n4910), .A2(n4887), .ZN(n4371) );
  AND2_X1 U5910 ( .A1(n5385), .A2(n5365), .ZN(n4372) );
  AND2_X1 U5911 ( .A1(n8182), .A2(n4400), .ZN(n4373) );
  AND2_X1 U5912 ( .A1(n4925), .A2(n4705), .ZN(n4374) );
  INV_X1 U5913 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n4928) );
  OR2_X1 U5914 ( .A1(n4421), .A2(n4337), .ZN(n4375) );
  INV_X1 U5915 ( .A(n4812), .ZN(n4811) );
  OR2_X1 U5916 ( .A1(n4814), .A2(n7911), .ZN(n4812) );
  INV_X1 U5917 ( .A(n4757), .ZN(n4756) );
  NAND2_X1 U5918 ( .A1(n4760), .A2(n4758), .ZN(n4757) );
  INV_X1 U5919 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n4523) );
  INV_X1 U5920 ( .A(n5513), .ZN(n7065) );
  INV_X2 U5922 ( .A(n9688), .ZN(n6638) );
  NAND2_X1 U5923 ( .A1(n7694), .A2(n8270), .ZN(n7721) );
  INV_X1 U5924 ( .A(n9013), .ZN(n4664) );
  NAND2_X1 U5925 ( .A1(n5371), .A2(n5370), .ZN(n8896) );
  INV_X1 U5926 ( .A(n8896), .ZN(n4527) );
  NAND2_X1 U5927 ( .A1(n4807), .A2(n4344), .ZN(n7941) );
  AND2_X1 U5928 ( .A1(n8772), .A2(n4877), .ZN(n4376) );
  NAND2_X1 U5929 ( .A1(n5608), .A2(n5607), .ZN(n8847) );
  AND2_X1 U5930 ( .A1(n4639), .A2(n5636), .ZN(n4435) );
  NAND2_X1 U5931 ( .A1(n5283), .A2(n4925), .ZN(n5323) );
  OAI22_X1 U5932 ( .A1(n6054), .A2(n4425), .B1(n6055), .B2(n4424), .ZN(n8997)
         );
  INV_X1 U5933 ( .A(n6125), .ZN(n4427) );
  NAND2_X1 U5934 ( .A1(n5668), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6039) );
  INV_X1 U5935 ( .A(n7971), .ZN(n4622) );
  INV_X1 U5936 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5588) );
  NAND2_X1 U5937 ( .A1(n5326), .A2(n5325), .ZN(n8905) );
  INV_X2 U5938 ( .A(n6246), .ZN(n6293) );
  AND2_X1 U5939 ( .A1(n6107), .A2(n6106), .ZN(n4377) );
  NAND2_X1 U5940 ( .A1(n9019), .A2(n6020), .ZN(n9032) );
  INV_X1 U5941 ( .A(n8088), .ZN(n8653) );
  AND2_X1 U5942 ( .A1(n5475), .A2(n5474), .ZN(n8088) );
  NAND2_X1 U5943 ( .A1(n8658), .A2(n4532), .ZN(n4533) );
  INV_X1 U5944 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n4416) );
  AND2_X1 U5945 ( .A1(n8413), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n4378) );
  NOR2_X1 U5946 ( .A1(n9460), .A2(n9383), .ZN(n4379) );
  NAND2_X1 U5947 ( .A1(n9739), .A2(n8228), .ZN(n8176) );
  INV_X1 U5948 ( .A(n8176), .ZN(n4855) );
  NAND2_X1 U5949 ( .A1(n4435), .A2(n5633), .ZN(n5923) );
  AND2_X1 U5950 ( .A1(n5342), .A2(SI_17_), .ZN(n4380) );
  INV_X1 U5951 ( .A(n8082), .ZN(n4685) );
  INV_X1 U5952 ( .A(n8899), .ZN(n8734) );
  NAND2_X1 U5953 ( .A1(n5347), .A2(n5346), .ZN(n8899) );
  NOR2_X1 U5954 ( .A1(n4507), .A2(n5495), .ZN(n4381) );
  NOR2_X1 U5955 ( .A1(n4789), .A2(n4791), .ZN(n5921) );
  AND2_X1 U5956 ( .A1(n4687), .A2(n5540), .ZN(n4382) );
  AND2_X1 U5957 ( .A1(n4766), .A2(n4765), .ZN(n4383) );
  AND2_X1 U5958 ( .A1(n7747), .A2(n5920), .ZN(n4384) );
  NAND2_X1 U5959 ( .A1(n6005), .A2(n6004), .ZN(n7939) );
  INV_X1 U5960 ( .A(n7939), .ZN(n4600) );
  NAND2_X1 U5961 ( .A1(n5212), .A2(n5211), .ZN(n7691) );
  INV_X1 U5962 ( .A(n7691), .ZN(n4534) );
  NAND2_X1 U5963 ( .A1(n6023), .A2(n6022), .ZN(n9470) );
  INV_X1 U5964 ( .A(n9470), .ZN(n4599) );
  NAND2_X1 U5965 ( .A1(n6820), .A2(n8201), .ZN(n5610) );
  INV_X1 U5966 ( .A(n5610), .ZN(n4702) );
  OR2_X1 U5967 ( .A1(n7804), .A2(n8934), .ZN(n7645) );
  INV_X1 U5968 ( .A(n7645), .ZN(n4536) );
  INV_X1 U5969 ( .A(n4996), .ZN(n5063) );
  INV_X1 U5970 ( .A(n7382), .ZN(n4615) );
  OAI21_X1 U5971 ( .B1(n7074), .B2(n7073), .A(n5100), .ZN(n7100) );
  OAI211_X1 U5972 ( .C1(n4854), .C2(n4396), .A(n4395), .B(n8209), .ZN(n7405)
         );
  NAND2_X1 U5973 ( .A1(n4419), .A2(n4418), .ZN(n7514) );
  NAND2_X1 U5974 ( .A1(n4642), .A2(n5880), .ZN(n7682) );
  NAND2_X1 U5975 ( .A1(n5307), .A2(n5306), .ZN(n8918) );
  INV_X1 U5976 ( .A(n8918), .ZN(n4538) );
  NAND2_X1 U5977 ( .A1(n5393), .A2(n5392), .ZN(n8889) );
  INV_X1 U5978 ( .A(n8889), .ZN(n4526) );
  OR2_X1 U5979 ( .A1(n6003), .A2(n5645), .ZN(n4385) );
  AND3_X1 U5980 ( .A1(n8118), .A2(n8116), .A3(n8117), .ZN(n4386) );
  NAND2_X1 U5981 ( .A1(n4641), .A2(n4640), .ZN(n7745) );
  NAND2_X1 U5982 ( .A1(n4911), .A2(n4910), .ZN(n5584) );
  NAND2_X1 U5983 ( .A1(n4700), .A2(n4699), .ZN(n7240) );
  AND2_X1 U5984 ( .A1(n6269), .A2(n6268), .ZN(n4387) );
  INV_X1 U5985 ( .A(n4509), .ZN(n4508) );
  NAND2_X1 U5986 ( .A1(n5464), .A2(n5492), .ZN(n4509) );
  AND2_X1 U5987 ( .A1(n7386), .A2(n7301), .ZN(n4388) );
  INV_X1 U5988 ( .A(n4911), .ZN(n5586) );
  NAND2_X1 U5989 ( .A1(n4938), .A2(n4939), .ZN(n5620) );
  INV_X1 U5990 ( .A(n7448), .ZN(n4517) );
  NAND2_X1 U5991 ( .A1(n5763), .A2(n5760), .ZN(n6946) );
  OAI22_X1 U5992 ( .A1(n6986), .A2(n6987), .B1(n5008), .B2(n5007), .ZN(n6974)
         );
  NOR2_X1 U5993 ( .A1(n4520), .A2(n9788), .ZN(n4389) );
  NAND2_X1 U5994 ( .A1(n4936), .A2(n4935), .ZN(n8569) );
  XNOR2_X1 U5995 ( .A(n5670), .B(n5669), .ZN(n7936) );
  INV_X1 U5996 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n4752) );
  NAND2_X1 U5997 ( .A1(n4572), .A2(n8338), .ZN(n4459) );
  NAND2_X1 U5998 ( .A1(n4746), .A2(n7205), .ZN(n4745) );
  NAND2_X2 U5999 ( .A1(n8792), .A2(n8799), .ZN(n8791) );
  NAND2_X1 U6000 ( .A1(n4477), .A2(n5129), .ZN(n5157) );
  INV_X1 U6001 ( .A(n4753), .ZN(n8636) );
  NAND2_X1 U6002 ( .A1(n8710), .A2(n4392), .ZN(n4391) );
  NAND3_X1 U6003 ( .A1(n4391), .A2(n4879), .A3(n4390), .ZN(n8643) );
  NOR2_X1 U6004 ( .A1(n4398), .A2(n7210), .ZN(n4397) );
  NAND2_X1 U6005 ( .A1(n7276), .A2(n4401), .ZN(n4399) );
  NAND2_X1 U6006 ( .A1(n4373), .A2(n4399), .ZN(n7653) );
  NAND2_X1 U6007 ( .A1(n4407), .A2(n7696), .ZN(n4405) );
  NAND3_X1 U6008 ( .A1(n4406), .A2(n4405), .A3(n4859), .ZN(n8770) );
  OR2_X1 U6009 ( .A1(n7030), .A2(n7355), .ZN(n8228) );
  NAND4_X1 U6010 ( .A1(n4926), .A2(n5591), .A3(n4924), .A4(n4906), .ZN(n4908)
         );
  INV_X2 U6011 ( .A(n6875), .ZN(n6694) );
  NAND2_X1 U6012 ( .A1(n4369), .A2(n7937), .ZN(n5728) );
  NAND2_X1 U6013 ( .A1(n4335), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5749) );
  NAND2_X1 U6014 ( .A1(n7481), .A2(n4375), .ZN(n4419) );
  NAND2_X1 U6015 ( .A1(n8997), .A2(n8995), .ZN(n6075) );
  OAI21_X1 U6016 ( .B1(n9050), .B2(n4431), .A(n4429), .ZN(n6124) );
  NAND2_X1 U6017 ( .A1(n9050), .A2(n4429), .ZN(n4428) );
  NAND4_X1 U6018 ( .A1(n5642), .A2(n4639), .A3(n5633), .A4(n5636), .ZN(n6003)
         );
  INV_X1 U6020 ( .A(n7745), .ZN(n5915) );
  AND2_X2 U6021 ( .A1(n4447), .A2(n7040), .ZN(n4986) );
  NAND2_X1 U6022 ( .A1(n4700), .A2(n4450), .ZN(n4449) );
  NAND2_X1 U6023 ( .A1(n4930), .A2(n4455), .ZN(n4454) );
  XNOR2_X2 U6024 ( .A(n5485), .B(n5486), .ZN(n8057) );
  NOR2_X1 U6025 ( .A1(n4923), .A2(n8962), .ZN(n5282) );
  NAND2_X1 U6026 ( .A1(n4923), .A2(n4704), .ZN(n4931) );
  AND2_X1 U6027 ( .A1(n4923), .A2(n4924), .ZN(n5283) );
  NAND3_X1 U6028 ( .A1(n4493), .A2(n4492), .A3(n4943), .ZN(n4960) );
  AOI21_X1 U6029 ( .B1(n8248), .B2(n4467), .A(n4402), .ZN(n8245) );
  NAND2_X1 U6030 ( .A1(n4468), .A2(n8240), .ZN(n8248) );
  OAI21_X1 U6031 ( .B1(n4470), .B2(n4469), .A(n8326), .ZN(n4591) );
  NAND2_X1 U6032 ( .A1(n4846), .A2(n4848), .ZN(n4472) );
  NAND2_X1 U6033 ( .A1(n4846), .A2(n8629), .ZN(n4473) );
  NAND2_X1 U6034 ( .A1(n5106), .A2(n4478), .ZN(n4474) );
  NAND2_X1 U6035 ( .A1(n4474), .A2(n4475), .ZN(n5178) );
  OAI21_X1 U6036 ( .B1(n5180), .B2(n4486), .A(n4483), .ZN(n5248) );
  NAND2_X1 U6037 ( .A1(n5272), .A2(n4496), .ZN(n4494) );
  NAND2_X1 U6038 ( .A1(n4494), .A2(n4495), .ZN(n4735) );
  AOI21_X1 U6039 ( .B1(n5465), .B2(n4502), .A(n4381), .ZN(n4506) );
  NAND2_X1 U6040 ( .A1(n4524), .A2(n4522), .ZN(n4939) );
  NAND2_X1 U6041 ( .A1(n4525), .A2(P2_IR_REG_28__SCAN_IN), .ZN(n4524) );
  INV_X1 U6042 ( .A(n4533), .ZN(n8622) );
  NOR2_X1 U6043 ( .A1(n4947), .A2(n4539), .ZN(n6862) );
  MUX2_X1 U6044 ( .A(n6890), .B(P2_REG2_REG_1__SCAN_IN), .S(n4947), .Z(n9522)
         );
  INV_X1 U6045 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n4540) );
  NAND2_X1 U6046 ( .A1(n4560), .A2(n4849), .ZN(P2_U3244) );
  AND2_X2 U6047 ( .A1(n4923), .A2(n4909), .ZN(n4911) );
  AND2_X2 U6048 ( .A1(n4905), .A2(n5039), .ZN(n4923) );
  AOI21_X1 U6049 ( .B1(n8248), .B2(n4893), .A(n4565), .ZN(n8253) );
  NAND2_X1 U6050 ( .A1(n8290), .A2(n4577), .ZN(n4576) );
  NAND2_X1 U6051 ( .A1(n8290), .A2(n4583), .ZN(n8296) );
  AND2_X1 U6052 ( .A1(n8289), .A2(n8291), .ZN(n4583) );
  AND3_X2 U6053 ( .A1(n4584), .A2(n4324), .A3(n4585), .ZN(n8970) );
  NAND2_X2 U6054 ( .A1(n5801), .A2(n4994), .ZN(n5838) );
  NAND2_X2 U6055 ( .A1(n4592), .A2(n5650), .ZN(n7983) );
  NAND2_X1 U6056 ( .A1(n9239), .A2(n4593), .ZN(n4597) );
  NAND2_X1 U6057 ( .A1(n9239), .A2(n4828), .ZN(n9223) );
  NAND2_X1 U6058 ( .A1(n4334), .A2(n7832), .ZN(n9390) );
  NAND3_X1 U6059 ( .A1(n9298), .A2(n4605), .A3(n4604), .ZN(n4603) );
  INV_X1 U6060 ( .A(n4607), .ZN(n9279) );
  AND2_X1 U6061 ( .A1(n4608), .A2(n6491), .ZN(n7228) );
  NAND2_X1 U6062 ( .A1(n6305), .A2(n7234), .ZN(n4608) );
  INV_X1 U6063 ( .A(n7115), .ZN(n4610) );
  NAND2_X1 U6064 ( .A1(n4609), .A2(n6496), .ZN(n7137) );
  NAND2_X1 U6065 ( .A1(n7252), .A2(n4611), .ZN(n4614) );
  NAND2_X1 U6066 ( .A1(n4614), .A2(n4613), .ZN(n7367) );
  NAND2_X1 U6067 ( .A1(n7369), .A2(n4617), .ZN(n7617) );
  NAND2_X1 U6068 ( .A1(n7617), .A2(n7616), .ZN(n4618) );
  NAND3_X1 U6069 ( .A1(n4619), .A2(n5644), .A3(n5671), .ZN(n5645) );
  NAND2_X1 U6070 ( .A1(n9350), .A2(n4624), .ZN(n4623) );
  OR2_X1 U6071 ( .A1(n9229), .A2(n9228), .ZN(n9233) );
  NAND2_X2 U6072 ( .A1(n6492), .A2(n6495), .ZN(n6934) );
  MUX2_X1 U6073 ( .A(n8255), .B(n8254), .S(n8338), .Z(n8256) );
  NAND2_X2 U6074 ( .A1(n7135), .A2(n6379), .ZN(n7252) );
  INV_X1 U6075 ( .A(n4793), .ZN(n4792) );
  INV_X2 U6076 ( .A(n5784), .ZN(n5633) );
  NAND2_X1 U6077 ( .A1(n7514), .A2(n4643), .ZN(n4641) );
  OAI21_X1 U6078 ( .B1(n5668), .B2(P1_IR_REG_18__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5681) );
  INV_X1 U6079 ( .A(n4646), .ZN(n5675) );
  NAND3_X1 U6080 ( .A1(n9099), .A2(n9021), .A3(n9020), .ZN(n9019) );
  NAND2_X1 U6081 ( .A1(n8984), .A2(n4657), .ZN(n4655) );
  OR2_X1 U6082 ( .A1(n4660), .A2(n8984), .ZN(n4659) );
  NAND3_X1 U6083 ( .A1(n4656), .A2(n4661), .A3(n4655), .ZN(n9088) );
  NAND2_X1 U6084 ( .A1(n6163), .A2(n6162), .ZN(n4667) );
  AND2_X1 U6085 ( .A1(n5842), .A2(n5828), .ZN(n4671) );
  NAND2_X1 U6086 ( .A1(n4672), .A2(n4671), .ZN(n7481) );
  NAND3_X1 U6087 ( .A1(n5491), .A2(n5490), .A3(n4382), .ZN(n4682) );
  NAND2_X1 U6088 ( .A1(n4682), .A2(n4368), .ZN(n5561) );
  NAND3_X1 U6089 ( .A1(n5491), .A2(n5490), .A3(n4687), .ZN(n4686) );
  NAND3_X1 U6090 ( .A1(n5491), .A2(n5490), .A3(n5489), .ZN(n8085) );
  NAND2_X1 U6091 ( .A1(n5574), .A2(n4690), .ZN(n4689) );
  OAI211_X1 U6092 ( .C1(n5574), .C2(n4692), .A(n4695), .B(n4689), .ZN(n5630)
         );
  INV_X1 U6093 ( .A(n5573), .ZN(n4696) );
  NAND2_X1 U6094 ( .A1(n8063), .A2(n4697), .ZN(n8121) );
  NAND2_X2 U6095 ( .A1(n8103), .A2(n5339), .ZN(n8140) );
  NAND2_X1 U6096 ( .A1(n5316), .A2(n4701), .ZN(n8103) );
  INV_X1 U6097 ( .A(n4931), .ZN(n4930) );
  NAND3_X1 U6098 ( .A1(n4720), .A2(n5084), .A3(n4718), .ZN(n5102) );
  NAND3_X1 U6099 ( .A1(n5060), .A2(n5080), .A3(n5059), .ZN(n4720) );
  OAI21_X1 U6100 ( .B1(n5519), .B2(n5518), .A(n5520), .ZN(n5542) );
  NAND2_X1 U6101 ( .A1(n5606), .A2(n4732), .ZN(n4730) );
  OAI21_X1 U6102 ( .B1(n5606), .B2(n4734), .A(n4732), .ZN(n6301) );
  NAND2_X1 U6103 ( .A1(n4730), .A2(n4731), .ZN(n6270) );
  NAND2_X1 U6104 ( .A1(n5606), .A2(n5605), .ZN(n6267) );
  NAND2_X1 U6105 ( .A1(n4735), .A2(n4372), .ZN(n5387) );
  NAND3_X1 U6106 ( .A1(n4738), .A2(n6489), .A3(n4736), .ZN(n6538) );
  NAND2_X2 U6107 ( .A1(n5655), .A2(P1_U3084), .ZN(n9510) );
  MUX2_X1 U6108 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n5655), .Z(n5061) );
  MUX2_X1 U6109 ( .A(n10041), .B(n6658), .S(n5655), .Z(n5082) );
  MUX2_X1 U6110 ( .A(n6667), .B(n6660), .S(n5655), .Z(n5103) );
  MUX2_X1 U6111 ( .A(n6674), .B(n6676), .S(n5655), .Z(n5108) );
  MUX2_X1 U6112 ( .A(n6679), .B(n5130), .S(n5655), .Z(n5132) );
  MUX2_X1 U6113 ( .A(n5159), .B(n6685), .S(n5655), .Z(n5161) );
  MUX2_X1 U6114 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(P1_DATAO_REG_11__SCAN_IN), 
        .S(n5655), .Z(n5200) );
  MUX2_X1 U6115 ( .A(n6720), .B(n6722), .S(n5655), .Z(n5226) );
  MUX2_X1 U6116 ( .A(n6738), .B(n6737), .S(n5655), .Z(n5268) );
  MUX2_X1 U6117 ( .A(n6970), .B(n6968), .S(n5655), .Z(n5279) );
  MUX2_X1 U6118 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(P1_DATAO_REG_18__SCAN_IN), 
        .S(n5655), .Z(n5364) );
  MUX2_X1 U6119 ( .A(n7129), .B(n7131), .S(n5655), .Z(n5367) );
  MUX2_X1 U6120 ( .A(n7341), .B(n7351), .S(n5655), .Z(n5424) );
  MUX2_X1 U6121 ( .A(n10076), .B(n7989), .S(n5655), .Z(n5430) );
  MUX2_X1 U6122 ( .A(n5451), .B(n5452), .S(n5655), .Z(n5454) );
  MUX2_X1 U6123 ( .A(n7826), .B(n5497), .S(n5655), .Z(n5499) );
  MUX2_X1 U6124 ( .A(n7931), .B(n7889), .S(n5655), .Z(n5522) );
  MUX2_X1 U6125 ( .A(n5544), .B(n7928), .S(n5655), .Z(n5546) );
  MUX2_X1 U6126 ( .A(n9511), .B(n9988), .S(n5655), .Z(n6269) );
  MUX2_X1 U6127 ( .A(n7938), .B(n6272), .S(n5655), .Z(n6274) );
  MUX2_X1 U6128 ( .A(n6705), .B(n8170), .S(n5655), .Z(n6278) );
  NAND2_X2 U6129 ( .A1(P1_U3084), .A2(n4994), .ZN(n9508) );
  NAND2_X1 U6130 ( .A1(n7450), .A2(n8247), .ZN(n4747) );
  NAND2_X1 U6131 ( .A1(n4744), .A2(n7452), .ZN(n4743) );
  INV_X1 U6132 ( .A(n7450), .ZN(n4744) );
  OAI21_X1 U6133 ( .B1(n7205), .B2(n4744), .A(n4746), .ZN(n7636) );
  NAND2_X1 U6134 ( .A1(n4745), .A2(n4352), .ZN(n7803) );
  NAND2_X1 U6135 ( .A1(n7658), .A2(n7450), .ZN(n7659) );
  NAND2_X1 U6136 ( .A1(n6875), .A2(n4748), .ZN(n4751) );
  NAND2_X1 U6137 ( .A1(n4750), .A2(n4749), .ZN(n4748) );
  OAI21_X1 U6138 ( .B1(n8688), .B2(n4757), .A(n4754), .ZN(n4753) );
  AND2_X1 U6139 ( .A1(n8873), .A2(n8645), .ZN(n4763) );
  AND2_X1 U6140 ( .A1(n8783), .A2(n8801), .ZN(n4769) );
  NAND2_X1 U6141 ( .A1(n7721), .A2(n4370), .ZN(n8000) );
  OAI21_X1 U6142 ( .B1(n8606), .B2(n4774), .A(n4771), .ZN(n8018) );
  AOI21_X2 U6143 ( .B1(n8594), .B2(n8599), .A(n4780), .ZN(n8583) );
  NAND2_X1 U6144 ( .A1(n4911), .A2(n4371), .ZN(n4782) );
  NAND2_X1 U6145 ( .A1(n4785), .A2(n4787), .ZN(n7789) );
  NAND2_X1 U6146 ( .A1(n7755), .A2(n7757), .ZN(n4785) );
  INV_X1 U6147 ( .A(n4791), .ZN(n5804) );
  NAND2_X1 U6148 ( .A1(n7944), .A2(n4796), .ZN(n4795) );
  NAND2_X1 U6149 ( .A1(n4795), .A2(n4798), .ZN(n9343) );
  OAI21_X1 U6150 ( .B1(n7386), .B2(n4806), .A(n4804), .ZN(n7612) );
  OR2_X1 U6151 ( .A1(n9238), .A2(n7958), .ZN(n4830) );
  NAND2_X1 U6152 ( .A1(n4819), .A2(n4820), .ZN(n7961) );
  NAND2_X1 U6153 ( .A1(n7950), .A2(n4832), .ZN(n4831) );
  NAND2_X1 U6154 ( .A1(n4831), .A2(n4834), .ZN(n9254) );
  NAND2_X1 U6155 ( .A1(n9740), .A2(n9739), .ZN(n4854) );
  AND2_X1 U6156 ( .A1(n4956), .A2(n4955), .ZN(n4858) );
  NAND3_X1 U6157 ( .A1(n4957), .A2(n4858), .A3(n4954), .ZN(n8380) );
  NAND2_X1 U6158 ( .A1(n6822), .A2(n9770), .ZN(n7092) );
  NAND2_X1 U6159 ( .A1(n8588), .A2(n4867), .ZN(n4866) );
  NAND2_X1 U6160 ( .A1(n8588), .A2(n8589), .ZN(n4870) );
  OAI21_X1 U6161 ( .B1(n8024), .B2(n4876), .A(n4874), .ZN(n8737) );
  NOR2_X1 U6162 ( .A1(n5584), .A2(n4886), .ZN(n4937) );
  NAND3_X1 U6163 ( .A1(n4912), .A2(n4887), .A3(n4523), .ZN(n4886) );
  INV_X1 U6164 ( .A(n8970), .ZN(n4918) );
  AOI21_X1 U6165 ( .B1(n9416), .B2(n9578), .A(n9415), .ZN(n9488) );
  NAND2_X1 U6166 ( .A1(n6469), .A2(n6471), .ZN(n6483) );
  NAND2_X1 U6167 ( .A1(n6473), .A2(n6472), .ZN(n6482) );
  NAND2_X1 U6168 ( .A1(n5727), .A2(n6801), .ZN(n6832) );
  NAND2_X1 U6169 ( .A1(n5751), .A2(n5750), .ZN(n5754) );
  AND2_X1 U6170 ( .A1(n6306), .A2(n7109), .ZN(n7224) );
  NAND2_X1 U6171 ( .A1(n5736), .A2(n5735), .ZN(n5737) );
  INV_X1 U6172 ( .A(n4335), .ZN(n6296) );
  NAND2_X1 U6173 ( .A1(n6802), .A2(n6800), .ZN(n6801) );
  NAND2_X1 U6174 ( .A1(n6305), .A2(n6618), .ZN(n6619) );
  INV_X1 U6175 ( .A(n6309), .ZN(n9132) );
  XNOR2_X1 U6176 ( .A(n6280), .B(n6279), .ZN(n8169) );
  CLKBUF_X1 U6177 ( .A(n7206), .Z(n7207) );
  NOR2_X2 U6178 ( .A1(n5650), .A2(P1_IR_REG_28__SCAN_IN), .ZN(n5698) );
  XNOR2_X1 U6179 ( .A(n7981), .B(n7980), .ZN(n7985) );
  INV_X1 U6180 ( .A(n8847), .ZN(n5613) );
  AND2_X1 U6181 ( .A1(n6237), .A2(n9087), .ZN(n4888) );
  NAND3_X1 U6182 ( .A1(n5665), .A2(n5664), .A3(n5661), .ZN(n4889) );
  OR2_X1 U6183 ( .A1(n6301), .A2(n6298), .ZN(n4890) );
  AND2_X1 U6184 ( .A1(n5022), .A2(n5021), .ZN(n4891) );
  OR4_X1 U6185 ( .A1(n6767), .A2(n7305), .A3(n6249), .A4(n7983), .ZN(n4892) );
  AND2_X1 U6186 ( .A1(n8198), .A2(n8358), .ZN(n8751) );
  INV_X1 U6187 ( .A(n9231), .ZN(n7960) );
  AND2_X1 U6188 ( .A1(n8247), .A2(n8246), .ZN(n4893) );
  AND2_X1 U6189 ( .A1(n6481), .A2(n6487), .ZN(n4895) );
  NAND2_X1 U6190 ( .A1(n6467), .A2(n6297), .ZN(n6326) );
  INV_X1 U6191 ( .A(n8646), .ZN(n8150) );
  AND2_X1 U6192 ( .A1(n5725), .A2(n5724), .ZN(n4896) );
  AND2_X1 U6193 ( .A1(n5629), .A2(n5628), .ZN(n4897) );
  NAND2_X1 U6194 ( .A1(n5658), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5663) );
  NAND2_X1 U6195 ( .A1(n8215), .A2(n8322), .ZN(n8238) );
  INV_X1 U6196 ( .A(n8338), .ZN(n8322) );
  NAND2_X1 U6197 ( .A1(n8323), .A2(n8322), .ZN(n8324) );
  AND2_X1 U6198 ( .A1(n8325), .A2(n8324), .ZN(n8326) );
  INV_X1 U6199 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n4902) );
  INV_X1 U6200 ( .A(n6471), .ZN(n6472) );
  INV_X1 U6201 ( .A(n8704), .ZN(n8028) );
  INV_X1 U6202 ( .A(n5755), .ZN(n5756) );
  NAND2_X1 U6203 ( .A1(n6544), .A2(P1_IR_REG_0__SCAN_IN), .ZN(n5724) );
  INV_X1 U6204 ( .A(n6487), .ZN(n6524) );
  INV_X1 U6205 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5667) );
  XNOR2_X1 U6206 ( .A(n4986), .B(n8826), .ZN(n4952) );
  INV_X1 U6207 ( .A(n5396), .ZN(n5394) );
  OR2_X1 U6208 ( .A1(n5435), .A2(n8131), .ZN(n5476) );
  INV_X1 U6209 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n4913) );
  INV_X1 U6210 ( .A(n5283), .ZN(n5321) );
  OAI22_X1 U6211 ( .A1(n7134), .A2(n6209), .B1(n9706), .B2(n5756), .ZN(n5774)
         );
  INV_X1 U6212 ( .A(n5857), .ZN(n5858) );
  INV_X1 U6213 ( .A(n7251), .ZN(n6625) );
  INV_X1 U6214 ( .A(n7816), .ZN(n5263) );
  INV_X1 U6215 ( .A(n5143), .ZN(n5141) );
  INV_X1 U6216 ( .A(n8105), .ZN(n5338) );
  INV_X1 U6217 ( .A(n5528), .ZN(n5527) );
  OR3_X1 U6218 ( .A1(n5505), .A2(n8086), .A3(n5504), .ZN(n5528) );
  OR2_X1 U6219 ( .A1(n5413), .A2(n8076), .ZN(n5435) );
  NAND2_X1 U6220 ( .A1(n5394), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5413) );
  INV_X1 U6221 ( .A(n4318), .ZN(n5044) );
  NAND2_X1 U6222 ( .A1(n7640), .A2(n8243), .ZN(n7808) );
  OR2_X1 U6223 ( .A1(n5184), .A2(n5183), .ZN(n5209) );
  XNOR2_X1 U6224 ( .A(n5774), .B(n6212), .ZN(n5775) );
  INV_X1 U6225 ( .A(n5811), .ZN(n5685) );
  NAND2_X1 U6226 ( .A1(n5646), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5653) );
  INV_X1 U6227 ( .A(n6241), .ZN(n6614) );
  INV_X1 U6228 ( .A(n7979), .ZN(n7980) );
  NAND2_X1 U6229 ( .A1(n6241), .A2(n9282), .ZN(n6471) );
  NOR2_X1 U6230 ( .A1(n5641), .A2(n5640), .ZN(n5642) );
  NAND2_X1 U6231 ( .A1(n5226), .A2(n5225), .ZN(n5249) );
  NAND2_X1 U6232 ( .A1(n5132), .A2(n5131), .ZN(n5158) );
  INV_X1 U6233 ( .A(n8630), .ZN(n8087) );
  NAND2_X1 U6234 ( .A1(n6962), .A2(n6963), .ZN(n6961) );
  NAND2_X1 U6235 ( .A1(n8073), .A2(n5422), .ZN(n5445) );
  OR2_X1 U6236 ( .A1(n9825), .A2(n8569), .ZN(n6814) );
  INV_X1 U6237 ( .A(n8143), .ZN(n8159) );
  NAND2_X1 U6238 ( .A1(n8365), .A2(n8356), .ZN(n8198) );
  OR2_X1 U6239 ( .A1(n5373), .A2(n5372), .ZN(n5396) );
  NOR2_X1 U6240 ( .A1(n8863), .A2(n8646), .ZN(n8011) );
  NOR2_X1 U6241 ( .A1(n8371), .A2(n8899), .ZN(n8004) );
  OR2_X1 U6242 ( .A1(n9759), .A2(n6814), .ZN(n7668) );
  INV_X1 U6243 ( .A(n8578), .ZN(n8838) );
  AND2_X1 U6244 ( .A1(n8263), .A2(n8261), .ZN(n8187) );
  AND2_X1 U6245 ( .A1(n8237), .A2(n8231), .ZN(n8819) );
  INV_X1 U6246 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n8962) );
  NAND2_X1 U6247 ( .A1(n6181), .A2(n6183), .ZN(n6184) );
  NAND2_X1 U6248 ( .A1(n6532), .A2(n6531), .ZN(n6533) );
  INV_X1 U6249 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6759) );
  AND2_X1 U6250 ( .A1(n6447), .A2(n6449), .ZN(n9305) );
  OR2_X1 U6251 ( .A1(n7868), .A2(n9121), .ZN(n7829) );
  AND2_X1 U6252 ( .A1(n6614), .A2(n6775), .ZN(n6631) );
  INV_X1 U6253 ( .A(n9401), .ZN(n9331) );
  INV_X1 U6254 ( .A(n9406), .ZN(n9329) );
  INV_X1 U6255 ( .A(n9483), .ZN(n9714) );
  OAI21_X1 U6256 ( .B1(n5428), .B2(n5427), .A(n5426), .ZN(n5449) );
  NAND2_X1 U6257 ( .A1(n5222), .A2(n5208), .ZN(n5223) );
  NAND2_X1 U6258 ( .A1(n5129), .A2(n5110), .ZN(n5127) );
  NOR2_X1 U6259 ( .A1(n8068), .A2(n8754), .ZN(n8143) );
  OR2_X1 U6260 ( .A1(n5564), .A2(n5563), .ZN(n8019) );
  AND2_X1 U6261 ( .A1(n6877), .A2(n6876), .ZN(n9729) );
  INV_X1 U6262 ( .A(n9732), .ZN(n9728) );
  INV_X1 U6263 ( .A(n8677), .ZN(n8667) );
  AND2_X1 U6264 ( .A1(n8299), .A2(n8295), .ZN(n8718) );
  INV_X1 U6265 ( .A(n8756), .ZN(n9743) );
  OR2_X1 U6266 ( .A1(n9764), .A2(n5597), .ZN(n7272) );
  NOR2_X1 U6267 ( .A1(n7036), .A2(n6816), .ZN(n7274) );
  AND2_X1 U6268 ( .A1(n5138), .A2(n5164), .ZN(n8469) );
  INV_X1 U6269 ( .A(n9109), .ZN(n9094) );
  AOI21_X1 U6270 ( .B1(n9216), .B2(n4319), .A(n6208), .ZN(n9231) );
  INV_X1 U6271 ( .A(n9182), .ZN(n9673) );
  INV_X1 U6272 ( .A(n7959), .ZN(n9228) );
  INV_X1 U6273 ( .A(n9333), .ZN(n9403) );
  NAND2_X1 U6274 ( .A1(n5792), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5811) );
  INV_X1 U6275 ( .A(n9396), .ZN(n9316) );
  AND2_X1 U6276 ( .A1(n6932), .A2(n7936), .ZN(n9559) );
  AND2_X1 U6277 ( .A1(n6841), .A2(n6766), .ZN(n7393) );
  OR3_X1 U6278 ( .A1(n7933), .A2(n6220), .A3(n6219), .ZN(n6772) );
  XNOR2_X1 U6279 ( .A(n5103), .B(SI_7_), .ZN(n5101) );
  INV_X1 U6280 ( .A(n5616), .ZN(n8163) );
  INV_X1 U6281 ( .A(n8166), .ZN(n8146) );
  NAND2_X1 U6282 ( .A1(n5556), .A2(n5555), .ZN(n8615) );
  OR2_X1 U6283 ( .A1(n6859), .A2(n9762), .ZN(n8370) );
  XNOR2_X1 U6284 ( .A(n8018), .B(n8034), .ZN(n8846) );
  AND2_X1 U6285 ( .A1(n7733), .A2(n7732), .ZN(n8933) );
  INV_X1 U6286 ( .A(n9848), .ZN(n9846) );
  INV_X1 U6287 ( .A(n9833), .ZN(n9831) );
  INV_X1 U6288 ( .A(n9761), .ZN(n9765) );
  INV_X1 U6289 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6685) );
  INV_X1 U6290 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6658) );
  INV_X1 U6291 ( .A(n9112), .ZN(n9097) );
  AOI22_X1 U6292 ( .A1(n6538), .A2(n6537), .B1(n6536), .B2(n4892), .ZN(n6539)
         );
  NAND2_X1 U6293 ( .A1(n6140), .A2(n6139), .ZN(n9265) );
  NAND2_X1 U6294 ( .A1(n9321), .A2(n9681), .ZN(n9396) );
  NAND2_X1 U6295 ( .A1(n6637), .A2(n9692), .ZN(n9688) );
  INV_X1 U6296 ( .A(n9486), .ZN(n9725) );
  NAND3_X1 U6297 ( .A1(n6953), .A2(n7393), .A3(n9697), .ZN(n9721) );
  INV_X1 U6298 ( .A(n6775), .ZN(n7342) );
  INV_X1 U6299 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6679) );
  NOR2_X1 U6300 ( .A1(n9876), .A2(n9875), .ZN(n9874) );
  AND2_X1 U6301 ( .A1(n6576), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U4006) );
  INV_X1 U6302 ( .A(n6539), .ZN(P1_U3240) );
  NOR2_X2 U6303 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n4969) );
  NOR2_X1 U6304 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n4898) );
  NAND2_X1 U6305 ( .A1(n4969), .A2(n4898), .ZN(n5016) );
  NOR2_X1 U6306 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n4901) );
  NOR2_X1 U6307 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n4900) );
  NAND4_X1 U6308 ( .A1(n4901), .A2(n4900), .A3(n5085), .A4(n5182), .ZN(n4904)
         );
  NAND4_X1 U6309 ( .A1(n9893), .A2(n5251), .A3(n5181), .A4(n4902), .ZN(n4903)
         );
  NOR2_X1 U6310 ( .A1(n4904), .A2(n4903), .ZN(n4905) );
  INV_X1 U6311 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n4906) );
  NAND4_X1 U6312 ( .A1(n5588), .A2(n4928), .A3(n4705), .A4(n4925), .ZN(n4907)
         );
  NOR2_X1 U6313 ( .A1(n4908), .A2(n4907), .ZN(n4909) );
  INV_X1 U6314 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n4912) );
  INV_X1 U6315 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n4914) );
  XNOR2_X2 U6316 ( .A(n4915), .B(n4914), .ZN(n4919) );
  NAND2_X1 U6317 ( .A1(n4318), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n4917) );
  NAND2_X1 U6318 ( .A1(n4974), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n4916) );
  AND2_X2 U6319 ( .A1(n4917), .A2(n4916), .ZN(n4922) );
  INV_X1 U6320 ( .A(n4919), .ZN(n8965) );
  NAND2_X1 U6321 ( .A1(n4323), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n4921) );
  NAND2_X1 U6322 ( .A1(n5213), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n4920) );
  NAND2_X1 U6323 ( .A1(n4927), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4929) );
  NAND2_X1 U6324 ( .A1(n4933), .A2(n4416), .ZN(n4935) );
  INV_X1 U6325 ( .A(n4933), .ZN(n4934) );
  NAND2_X1 U6326 ( .A1(n4934), .A2(P2_IR_REG_19__SCAN_IN), .ZN(n4936) );
  NAND2_X1 U6327 ( .A1(n6817), .A2(n5513), .ZN(n4951) );
  INV_X1 U6328 ( .A(n4951), .ZN(n4950) );
  NAND2_X1 U6329 ( .A1(n8343), .A2(n8346), .ZN(n7040) );
  INV_X1 U6330 ( .A(n4937), .ZN(n4938) );
  MUX2_X1 U6331 ( .A(P2_IR_REG_31__SCAN_IN), .B(n4940), .S(
        P2_IR_REG_27__SCAN_IN), .Z(n4942) );
  AND2_X1 U6332 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n4943) );
  AND2_X1 U6333 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n4944) );
  INV_X1 U6334 ( .A(SI_1_), .ZN(n4945) );
  XNOR2_X1 U6335 ( .A(n4966), .B(n4945), .ZN(n4965) );
  MUX2_X1 U6336 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n4994), .Z(n4964) );
  XNOR2_X1 U6337 ( .A(n4965), .B(n4964), .ZN(n6665) );
  NAND2_X1 U6338 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n4946) );
  OR2_X1 U6339 ( .A1(n6875), .A2(n4947), .ZN(n4948) );
  INV_X1 U6340 ( .A(n4952), .ZN(n4949) );
  NAND2_X1 U6341 ( .A1(n4950), .A2(n4949), .ZN(n4953) );
  NAND2_X1 U6342 ( .A1(n4952), .A2(n4951), .ZN(n4963) );
  NAND2_X1 U6343 ( .A1(n4953), .A2(n4963), .ZN(n7003) );
  INV_X1 U6344 ( .A(n7003), .ZN(n4962) );
  NAND2_X1 U6345 ( .A1(n4974), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n4957) );
  NAND2_X1 U6346 ( .A1(n5213), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n4956) );
  NAND2_X1 U6347 ( .A1(n5020), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n4955) );
  NAND2_X1 U6348 ( .A1(n4321), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n4954) );
  INV_X1 U6349 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n4958) );
  AND2_X1 U6350 ( .A1(n4960), .A2(n4959), .ZN(n8973) );
  MUX2_X1 U6351 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8973), .S(n6875), .Z(n9770) );
  NAND2_X1 U6352 ( .A1(n8380), .A2(n9770), .ZN(n6819) );
  OAI22_X1 U6353 ( .A1(n6819), .A2(n7065), .B1(n9770), .B2(n5115), .ZN(n7002)
         );
  INV_X1 U6354 ( .A(n7002), .ZN(n4961) );
  NAND2_X1 U6355 ( .A1(n4962), .A2(n4961), .ZN(n7000) );
  NAND2_X1 U6356 ( .A1(n7000), .A2(n4963), .ZN(n6912) );
  NAND2_X1 U6357 ( .A1(n4965), .A2(n4964), .ZN(n4968) );
  NAND2_X1 U6358 ( .A1(n4966), .A2(SI_1_), .ZN(n4967) );
  NAND2_X1 U6359 ( .A1(n4968), .A2(n4967), .ZN(n4989) );
  INV_X1 U6360 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6659) );
  INV_X1 U6361 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6672) );
  MUX2_X1 U6362 ( .A(n6659), .B(n6672), .S(n4994), .Z(n4990) );
  XNOR2_X1 U6363 ( .A(n4990), .B(SI_2_), .ZN(n4988) );
  XNOR2_X1 U6364 ( .A(n4989), .B(n4988), .ZN(n6671) );
  NAND2_X1 U6365 ( .A1(n4996), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n4972) );
  OR2_X1 U6366 ( .A1(n4969), .A2(n8962), .ZN(n4970) );
  XNOR2_X1 U6367 ( .A(n4970), .B(P2_IR_REG_2__SCAN_IN), .ZN(n9533) );
  XNOR2_X1 U6368 ( .A(n4986), .B(n7355), .ZN(n4981) );
  NAND2_X1 U6369 ( .A1(n4318), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n4976) );
  NAND2_X1 U6370 ( .A1(n4974), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n4975) );
  AND2_X1 U6371 ( .A1(n4976), .A2(n4975), .ZN(n4979) );
  NAND2_X1 U6372 ( .A1(n5020), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n4978) );
  NAND2_X1 U6373 ( .A1(n5213), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n4977) );
  NAND2_X1 U6374 ( .A1(n7029), .A2(n5513), .ZN(n4980) );
  NAND2_X1 U6375 ( .A1(n4981), .A2(n4980), .ZN(n4985) );
  INV_X1 U6376 ( .A(n4980), .ZN(n4983) );
  INV_X1 U6377 ( .A(n4981), .ZN(n4982) );
  NAND2_X1 U6378 ( .A1(n4983), .A2(n4982), .ZN(n4984) );
  AND2_X1 U6379 ( .A1(n4985), .A2(n4984), .ZN(n6913) );
  NAND2_X1 U6380 ( .A1(n6912), .A2(n6913), .ZN(n6911) );
  NAND2_X1 U6381 ( .A1(n6911), .A2(n4985), .ZN(n6986) );
  NAND2_X1 U6382 ( .A1(n4989), .A2(n4988), .ZN(n4993) );
  INV_X1 U6383 ( .A(n4990), .ZN(n4991) );
  NAND2_X1 U6384 ( .A1(n4991), .A2(SI_2_), .ZN(n4992) );
  NAND2_X1 U6385 ( .A1(n4993), .A2(n4992), .ZN(n5011) );
  INV_X1 U6386 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n4995) );
  INV_X1 U6387 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6655) );
  MUX2_X1 U6388 ( .A(n4995), .B(n6655), .S(n4994), .Z(n5012) );
  XNOR2_X1 U6389 ( .A(n5012), .B(SI_3_), .ZN(n5010) );
  XNOR2_X1 U6390 ( .A(n5011), .B(n5010), .ZN(n6654) );
  NAND2_X1 U6391 ( .A1(n4996), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n5000) );
  NAND2_X1 U6392 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n4997), .ZN(n4998) );
  XNOR2_X1 U6393 ( .A(n4998), .B(P2_IR_REG_3__SCAN_IN), .ZN(n8385) );
  NAND2_X1 U6394 ( .A1(n6694), .A2(n8385), .ZN(n4999) );
  XNOR2_X1 U6395 ( .A(n4986), .B(n9749), .ZN(n5008) );
  INV_X1 U6396 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n5001) );
  NAND2_X1 U6397 ( .A1(n5020), .A2(n5001), .ZN(n5004) );
  NAND2_X1 U6398 ( .A1(n5213), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5003) );
  NAND2_X1 U6399 ( .A1(n4974), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5002) );
  AND3_X1 U6400 ( .A1(n5004), .A2(n5003), .A3(n5002), .ZN(n5006) );
  NAND2_X1 U6401 ( .A1(n8035), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5005) );
  NAND2_X1 U6402 ( .A1(n8379), .A2(n5513), .ZN(n5007) );
  XNOR2_X1 U6403 ( .A(n5008), .B(n5007), .ZN(n6987) );
  INV_X1 U6404 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n5009) );
  INV_X1 U6405 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6663) );
  MUX2_X1 U6406 ( .A(n5009), .B(n6663), .S(n4994), .Z(n5033) );
  XNOR2_X1 U6407 ( .A(n5033), .B(SI_4_), .ZN(n5031) );
  NAND2_X1 U6408 ( .A1(n5011), .A2(n5010), .ZN(n5015) );
  INV_X1 U6409 ( .A(n5012), .ZN(n5013) );
  NAND2_X1 U6410 ( .A1(n5013), .A2(SI_3_), .ZN(n5014) );
  NAND2_X1 U6411 ( .A1(n5015), .A2(n5014), .ZN(n5032) );
  XNOR2_X1 U6412 ( .A(n5031), .B(n5032), .ZN(n6662) );
  NAND2_X1 U6413 ( .A1(n4996), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n5019) );
  NAND2_X1 U6414 ( .A1(n5016), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5017) );
  XNOR2_X1 U6415 ( .A(n5017), .B(P2_IR_REG_4__SCAN_IN), .ZN(n8399) );
  NAND2_X1 U6416 ( .A1(n6694), .A2(n8399), .ZN(n5018) );
  XNOR2_X1 U6417 ( .A(n4986), .B(n7045), .ZN(n5026) );
  NAND2_X1 U6418 ( .A1(n5213), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5024) );
  OAI21_X1 U6419 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(P2_REG3_REG_4__SCAN_IN), 
        .A(n5046), .ZN(n7051) );
  INV_X1 U6420 ( .A(n7051), .ZN(n6980) );
  NAND2_X1 U6421 ( .A1(n5020), .A2(n6980), .ZN(n5023) );
  NAND2_X1 U6422 ( .A1(n4974), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5022) );
  NAND2_X1 U6423 ( .A1(n4320), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5021) );
  INV_X1 U6424 ( .A(n7195), .ZN(n9745) );
  NAND2_X1 U6425 ( .A1(n9745), .A2(n5513), .ZN(n5025) );
  NAND2_X1 U6426 ( .A1(n5026), .A2(n5025), .ZN(n5030) );
  INV_X1 U6427 ( .A(n5025), .ZN(n5028) );
  INV_X1 U6428 ( .A(n5026), .ZN(n5027) );
  NAND2_X1 U6429 ( .A1(n5028), .A2(n5027), .ZN(n5029) );
  NAND2_X1 U6430 ( .A1(n5030), .A2(n5029), .ZN(n6977) );
  NAND2_X1 U6431 ( .A1(n6975), .A2(n5030), .ZN(n6962) );
  NAND2_X1 U6432 ( .A1(n5032), .A2(n5031), .ZN(n5036) );
  INV_X1 U6433 ( .A(n5033), .ZN(n5034) );
  NAND2_X1 U6434 ( .A1(n5034), .A2(SI_4_), .ZN(n5035) );
  INV_X1 U6435 ( .A(SI_5_), .ZN(n5037) );
  INV_X2 U6436 ( .A(n5063), .ZN(n8014) );
  NAND2_X1 U6437 ( .A1(n8014), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n5043) );
  NAND2_X1 U6438 ( .A1(n4329), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5038) );
  MUX2_X1 U6439 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5038), .S(
        P2_IR_REG_5__SCAN_IN), .Z(n5041) );
  INV_X1 U6440 ( .A(n5039), .ZN(n5040) );
  NAND2_X1 U6441 ( .A1(n6694), .A2(n8413), .ZN(n5042) );
  XNOR2_X1 U6442 ( .A(n4986), .B(n9794), .ZN(n5053) );
  NAND2_X1 U6443 ( .A1(n4320), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5051) );
  INV_X2 U6444 ( .A(n5624), .ZN(n8036) );
  NAND2_X1 U6445 ( .A1(n8036), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5050) );
  INV_X1 U6446 ( .A(n5046), .ZN(n5045) );
  NAND2_X1 U6447 ( .A1(n5045), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5068) );
  INV_X1 U6448 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n8411) );
  NAND2_X1 U6449 ( .A1(n5046), .A2(n8411), .ZN(n5047) );
  AND2_X1 U6450 ( .A1(n5068), .A2(n5047), .ZN(n6958) );
  NAND2_X1 U6451 ( .A1(n5020), .A2(n6958), .ZN(n5049) );
  NAND2_X1 U6452 ( .A1(n5213), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5048) );
  NAND2_X1 U6453 ( .A1(n8810), .A2(n5513), .ZN(n5052) );
  NAND2_X1 U6454 ( .A1(n5053), .A2(n5052), .ZN(n5057) );
  INV_X1 U6455 ( .A(n5052), .ZN(n5055) );
  INV_X1 U6456 ( .A(n5053), .ZN(n5054) );
  NAND2_X1 U6457 ( .A1(n5055), .A2(n5054), .ZN(n5056) );
  AND2_X1 U6458 ( .A1(n5057), .A2(n5056), .ZN(n6963) );
  NAND2_X1 U6459 ( .A1(n6961), .A2(n5057), .ZN(n6993) );
  OR2_X1 U6460 ( .A1(n5039), .A2(n8962), .ZN(n5058) );
  XNOR2_X1 U6461 ( .A(n5058), .B(P2_IR_REG_6__SCAN_IN), .ZN(n8427) );
  INV_X1 U6462 ( .A(n8427), .ZN(n6656) );
  NAND2_X1 U6463 ( .A1(n5061), .A2(SI_5_), .ZN(n5062) );
  XNOR2_X1 U6464 ( .A(n5081), .B(n5080), .ZN(n6657) );
  OR2_X1 U6465 ( .A1(n4987), .A2(n6657), .ZN(n5065) );
  NAND2_X1 U6466 ( .A1(n8014), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n5064) );
  OAI211_X1 U6467 ( .C1(n6875), .C2(n6656), .A(n5065), .B(n5064), .ZN(n9801)
         );
  XNOR2_X1 U6468 ( .A(n9801), .B(n4986), .ZN(n5074) );
  NAND2_X1 U6469 ( .A1(n8036), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5073) );
  NAND2_X1 U6470 ( .A1(n8035), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5072) );
  INV_X1 U6471 ( .A(n5068), .ZN(n5066) );
  NAND2_X1 U6472 ( .A1(n5066), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5090) );
  INV_X1 U6473 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n5067) );
  NAND2_X1 U6474 ( .A1(n5068), .A2(n5067), .ZN(n5069) );
  AND2_X1 U6475 ( .A1(n5090), .A2(n5069), .ZN(n8817) );
  NAND2_X1 U6476 ( .A1(n5020), .A2(n8817), .ZN(n5071) );
  NAND2_X1 U6477 ( .A1(n8037), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5070) );
  NAND4_X1 U6478 ( .A1(n5073), .A2(n5072), .A3(n5071), .A4(n5070), .ZN(n8378)
         );
  NAND2_X1 U6479 ( .A1(n8378), .A2(n5513), .ZN(n5075) );
  NAND2_X1 U6480 ( .A1(n5074), .A2(n5075), .ZN(n5079) );
  INV_X1 U6481 ( .A(n5074), .ZN(n5077) );
  INV_X1 U6482 ( .A(n5075), .ZN(n5076) );
  NAND2_X1 U6483 ( .A1(n5077), .A2(n5076), .ZN(n5078) );
  AND2_X1 U6484 ( .A1(n5079), .A2(n5078), .ZN(n6994) );
  NAND2_X1 U6485 ( .A1(n6993), .A2(n6994), .ZN(n6992) );
  NAND2_X1 U6486 ( .A1(n6992), .A2(n5079), .ZN(n7074) );
  INV_X1 U6487 ( .A(n5082), .ZN(n5083) );
  NAND2_X1 U6488 ( .A1(n5083), .A2(SI_6_), .ZN(n5084) );
  INV_X1 U6489 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6660) );
  INV_X1 U6490 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6667) );
  XNOR2_X1 U6491 ( .A(n5102), .B(n5101), .ZN(n6668) );
  OR2_X1 U6492 ( .A1(n6668), .A2(n4987), .ZN(n5088) );
  NAND2_X1 U6493 ( .A1(n5039), .A2(n5085), .ZN(n5111) );
  NAND2_X1 U6494 ( .A1(n5111), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5086) );
  XNOR2_X1 U6495 ( .A(n5086), .B(P2_IR_REG_7__SCAN_IN), .ZN(n8441) );
  AOI22_X1 U6496 ( .A1(n8014), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6694), .B2(
        n8441), .ZN(n5087) );
  NAND2_X1 U6497 ( .A1(n5088), .A2(n5087), .ZN(n7281) );
  XNOR2_X1 U6498 ( .A(n7281), .B(n4986), .ZN(n5096) );
  NAND2_X1 U6499 ( .A1(n8036), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5095) );
  NAND2_X1 U6500 ( .A1(n8037), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5094) );
  INV_X1 U6501 ( .A(n5090), .ZN(n5089) );
  NAND2_X1 U6502 ( .A1(n5089), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5117) );
  INV_X1 U6503 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n8439) );
  NAND2_X1 U6504 ( .A1(n5090), .A2(n8439), .ZN(n5091) );
  AND2_X1 U6505 ( .A1(n5117), .A2(n5091), .ZN(n7331) );
  NAND2_X1 U6506 ( .A1(n5020), .A2(n7331), .ZN(n5093) );
  NAND2_X1 U6507 ( .A1(n4320), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5092) );
  NAND4_X1 U6508 ( .A1(n5095), .A2(n5094), .A3(n5093), .A4(n5092), .ZN(n8811)
         );
  NAND2_X1 U6509 ( .A1(n8811), .A2(n5513), .ZN(n5097) );
  XNOR2_X1 U6510 ( .A(n5096), .B(n5097), .ZN(n7073) );
  INV_X1 U6511 ( .A(n5096), .ZN(n5099) );
  INV_X1 U6512 ( .A(n5097), .ZN(n5098) );
  NAND2_X1 U6513 ( .A1(n5099), .A2(n5098), .ZN(n5100) );
  NAND2_X1 U6514 ( .A1(n5102), .A2(n5101), .ZN(n5106) );
  INV_X1 U6515 ( .A(n5103), .ZN(n5104) );
  NAND2_X1 U6516 ( .A1(n5104), .A2(SI_7_), .ZN(n5105) );
  INV_X1 U6517 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6676) );
  INV_X1 U6518 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6674) );
  INV_X1 U6519 ( .A(SI_8_), .ZN(n5107) );
  INV_X1 U6520 ( .A(n5108), .ZN(n5109) );
  NAND2_X1 U6521 ( .A1(n5109), .A2(SI_8_), .ZN(n5110) );
  XNOR2_X1 U6522 ( .A(n5128), .B(n5127), .ZN(n6673) );
  NAND2_X1 U6523 ( .A1(n6673), .A2(n8171), .ZN(n5114) );
  NAND2_X1 U6524 ( .A1(n5184), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5112) );
  XNOR2_X1 U6525 ( .A(n5112), .B(P2_IR_REG_8__SCAN_IN), .ZN(n8455) );
  AOI22_X1 U6526 ( .A1(n8014), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6694), .B2(
        n8455), .ZN(n5113) );
  NAND2_X1 U6527 ( .A1(n5114), .A2(n5113), .ZN(n7448) );
  XNOR2_X1 U6528 ( .A(n7448), .B(n5115), .ZN(n5125) );
  NAND2_X1 U6529 ( .A1(n8035), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5122) );
  NAND2_X1 U6530 ( .A1(n8036), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5121) );
  NAND2_X1 U6531 ( .A1(n5117), .A2(n5116), .ZN(n5118) );
  AND2_X1 U6532 ( .A1(n5143), .A2(n5118), .ZN(n7217) );
  NAND2_X1 U6533 ( .A1(n5020), .A2(n7217), .ZN(n5120) );
  NAND2_X1 U6534 ( .A1(n5213), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5119) );
  NAND4_X1 U6535 ( .A1(n5122), .A2(n5121), .A3(n5120), .A4(n5119), .ZN(n8377)
         );
  NAND2_X1 U6536 ( .A1(n8377), .A2(n5513), .ZN(n5123) );
  XNOR2_X1 U6537 ( .A(n5125), .B(n5123), .ZN(n7101) );
  INV_X1 U6538 ( .A(n5123), .ZN(n5124) );
  NAND2_X1 U6539 ( .A1(n5125), .A2(n5124), .ZN(n5126) );
  INV_X1 U6540 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n5130) );
  INV_X1 U6541 ( .A(SI_9_), .ZN(n5131) );
  INV_X1 U6542 ( .A(n5132), .ZN(n5133) );
  NAND2_X1 U6543 ( .A1(n5133), .A2(SI_9_), .ZN(n5134) );
  XNOR2_X1 U6544 ( .A(n5157), .B(n5156), .ZN(n6677) );
  NAND2_X1 U6545 ( .A1(n6677), .A2(n8171), .ZN(n5140) );
  OR2_X1 U6546 ( .A1(n5184), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n5135) );
  NAND2_X1 U6547 ( .A1(n5135), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5137) );
  INV_X1 U6548 ( .A(n5137), .ZN(n5136) );
  NAND2_X1 U6549 ( .A1(n5136), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n5138) );
  NAND2_X1 U6550 ( .A1(n5137), .A2(n9893), .ZN(n5164) );
  AOI22_X1 U6551 ( .A1(n8014), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6694), .B2(
        n8469), .ZN(n5139) );
  XNOR2_X1 U6552 ( .A(n7772), .B(n4986), .ZN(n5149) );
  NAND2_X1 U6553 ( .A1(n4320), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5148) );
  NAND2_X1 U6554 ( .A1(n8036), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5147) );
  INV_X1 U6555 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5142) );
  NAND2_X1 U6556 ( .A1(n5143), .A2(n5142), .ZN(n5144) );
  AND2_X1 U6557 ( .A1(n5169), .A2(n5144), .ZN(n7667) );
  NAND2_X1 U6558 ( .A1(n5020), .A2(n7667), .ZN(n5146) );
  NAND2_X1 U6559 ( .A1(n5213), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5145) );
  NAND4_X1 U6560 ( .A1(n5148), .A2(n5147), .A3(n5146), .A4(n5145), .ZN(n8376)
         );
  NAND2_X1 U6561 ( .A1(n8376), .A2(n5513), .ZN(n5150) );
  NAND2_X1 U6562 ( .A1(n5149), .A2(n5150), .ZN(n5155) );
  INV_X1 U6563 ( .A(n5149), .ZN(n5152) );
  INV_X1 U6564 ( .A(n5150), .ZN(n5151) );
  NAND2_X1 U6565 ( .A1(n5152), .A2(n5151), .ZN(n5153) );
  NAND2_X1 U6566 ( .A1(n5155), .A2(n5153), .ZN(n7242) );
  INV_X1 U6567 ( .A(n7242), .ZN(n5154) );
  INV_X1 U6568 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n5159) );
  INV_X1 U6569 ( .A(SI_10_), .ZN(n5160) );
  INV_X1 U6570 ( .A(n5161), .ZN(n5162) );
  NAND2_X1 U6571 ( .A1(n5162), .A2(SI_10_), .ZN(n5163) );
  XNOR2_X1 U6572 ( .A(n5178), .B(n5177), .ZN(n6682) );
  NAND2_X1 U6573 ( .A1(n6682), .A2(n8171), .ZN(n5167) );
  NAND2_X1 U6574 ( .A1(n5164), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5165) );
  XNOR2_X1 U6575 ( .A(n5165), .B(P2_IR_REG_10__SCAN_IN), .ZN(n7016) );
  AOI22_X1 U6576 ( .A1(n8014), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6694), .B2(
        n7016), .ZN(n5166) );
  NAND2_X1 U6577 ( .A1(n5167), .A2(n5166), .ZN(n7634) );
  XNOR2_X1 U6578 ( .A(n7634), .B(n4986), .ZN(n5176) );
  NAND2_X1 U6579 ( .A1(n8036), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5174) );
  NAND2_X1 U6580 ( .A1(n5213), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5173) );
  INV_X1 U6581 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n5168) );
  NAND2_X1 U6582 ( .A1(n5169), .A2(n5168), .ZN(n5170) );
  AND2_X1 U6583 ( .A1(n5189), .A2(n5170), .ZN(n7460) );
  NAND2_X1 U6584 ( .A1(n5020), .A2(n7460), .ZN(n5172) );
  NAND2_X1 U6585 ( .A1(n4320), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5171) );
  NAND4_X1 U6586 ( .A1(n5174), .A2(n5173), .A3(n5172), .A4(n5171), .ZN(n8375)
         );
  NAND2_X1 U6587 ( .A1(n8375), .A2(n5513), .ZN(n5175) );
  XNOR2_X1 U6588 ( .A(n5176), .B(n5175), .ZN(n7343) );
  NAND2_X1 U6589 ( .A1(n5178), .A2(n5177), .ZN(n5180) );
  XNOR2_X1 U6590 ( .A(n5203), .B(n5199), .ZN(n6686) );
  NAND2_X1 U6591 ( .A1(n6686), .A2(n8171), .ZN(n5187) );
  NAND3_X1 U6592 ( .A1(n9893), .A2(n5182), .A3(n5181), .ZN(n5183) );
  NAND2_X1 U6593 ( .A1(n5209), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5185) );
  XNOR2_X1 U6594 ( .A(n5185), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7162) );
  AOI22_X1 U6595 ( .A1(n8014), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6694), .B2(
        n7162), .ZN(n5186) );
  NAND2_X1 U6596 ( .A1(n5187), .A2(n5186), .ZN(n8934) );
  XNOR2_X1 U6597 ( .A(n8934), .B(n4986), .ZN(n5195) );
  NAND2_X1 U6598 ( .A1(n8036), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5194) );
  NAND2_X1 U6599 ( .A1(n8037), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5193) );
  INV_X1 U6600 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n9881) );
  NAND2_X1 U6601 ( .A1(n5189), .A2(n9881), .ZN(n5190) );
  AND2_X1 U6602 ( .A1(n5235), .A2(n5190), .ZN(n7805) );
  NAND2_X1 U6603 ( .A1(n5020), .A2(n7805), .ZN(n5192) );
  NAND2_X1 U6604 ( .A1(n8035), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n5191) );
  NAND4_X1 U6605 ( .A1(n5194), .A2(n5193), .A3(n5192), .A4(n5191), .ZN(n8374)
         );
  NAND2_X1 U6606 ( .A1(n8374), .A2(n5513), .ZN(n5196) );
  NAND2_X1 U6607 ( .A1(n5195), .A2(n5196), .ZN(n7525) );
  INV_X1 U6608 ( .A(n5195), .ZN(n5198) );
  INV_X1 U6609 ( .A(n5196), .ZN(n5197) );
  NAND2_X1 U6610 ( .A1(n5198), .A2(n5197), .ZN(n7527) );
  NAND2_X1 U6611 ( .A1(n5200), .A2(SI_11_), .ZN(n5201) );
  INV_X1 U6612 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n5204) );
  INV_X1 U6613 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6700) );
  MUX2_X1 U6614 ( .A(n5204), .B(n6700), .S(n4994), .Z(n5206) );
  INV_X1 U6615 ( .A(SI_12_), .ZN(n5205) );
  INV_X1 U6616 ( .A(n5206), .ZN(n5207) );
  NAND2_X1 U6617 ( .A1(n5207), .A2(SI_12_), .ZN(n5208) );
  XNOR2_X1 U6618 ( .A(n5224), .B(n5223), .ZN(n6692) );
  NAND2_X1 U6619 ( .A1(n6692), .A2(n8171), .ZN(n5212) );
  NOR2_X1 U6620 ( .A1(n5209), .A2(P2_IR_REG_11__SCAN_IN), .ZN(n5230) );
  OR2_X1 U6621 ( .A1(n5230), .A2(n8962), .ZN(n5210) );
  XNOR2_X1 U6622 ( .A(n5210), .B(P2_IR_REG_12__SCAN_IN), .ZN(n8483) );
  AOI22_X1 U6623 ( .A1(n8014), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6694), .B2(
        n8483), .ZN(n5211) );
  XNOR2_X1 U6624 ( .A(n7691), .B(n4986), .ZN(n5218) );
  NAND2_X1 U6625 ( .A1(n8035), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5217) );
  NAND2_X1 U6626 ( .A1(n8036), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5216) );
  XNOR2_X1 U6627 ( .A(n5235), .B(P2_REG3_REG_12__SCAN_IN), .ZN(n7647) );
  NAND2_X1 U6628 ( .A1(n5020), .A2(n7647), .ZN(n5215) );
  NAND2_X1 U6629 ( .A1(n5213), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5214) );
  NAND4_X1 U6630 ( .A1(n5217), .A2(n5216), .A3(n5215), .A4(n5214), .ZN(n8373)
         );
  NAND2_X1 U6631 ( .A1(n8373), .A2(n5513), .ZN(n5219) );
  NAND2_X1 U6632 ( .A1(n5218), .A2(n5219), .ZN(n7580) );
  INV_X1 U6633 ( .A(n5218), .ZN(n5221) );
  INV_X1 U6634 ( .A(n5219), .ZN(n5220) );
  NAND2_X1 U6635 ( .A1(n5221), .A2(n5220), .ZN(n7581) );
  INV_X1 U6636 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6722) );
  INV_X1 U6637 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n6720) );
  INV_X1 U6638 ( .A(SI_13_), .ZN(n5225) );
  INV_X1 U6639 ( .A(n5226), .ZN(n5227) );
  NAND2_X1 U6640 ( .A1(n5227), .A2(SI_13_), .ZN(n5228) );
  XNOR2_X1 U6641 ( .A(n5248), .B(n5247), .ZN(n6718) );
  NAND2_X1 U6642 ( .A1(n6718), .A2(n8171), .ZN(n5233) );
  INV_X1 U6643 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5229) );
  NAND2_X1 U6644 ( .A1(n5230), .A2(n5229), .ZN(n5231) );
  NAND2_X1 U6645 ( .A1(n5231), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5252) );
  XNOR2_X1 U6646 ( .A(n5252), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7318) );
  AOI22_X1 U6647 ( .A1(n8014), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6694), .B2(
        n7318), .ZN(n5232) );
  NAND2_X1 U6648 ( .A1(n5233), .A2(n5232), .ZN(n7739) );
  XNOR2_X1 U6649 ( .A(n7739), .B(n5115), .ZN(n5241) );
  NAND2_X1 U6650 ( .A1(n8035), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5240) );
  NAND2_X1 U6651 ( .A1(n8036), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n5239) );
  INV_X1 U6652 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n5234) );
  INV_X1 U6653 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n7167) );
  OAI21_X1 U6654 ( .B1(n5235), .B2(n5234), .A(n7167), .ZN(n5236) );
  AND2_X1 U6655 ( .A1(n5236), .A2(n5257), .ZN(n7738) );
  NAND2_X1 U6656 ( .A1(n5020), .A2(n7738), .ZN(n5238) );
  NAND2_X1 U6657 ( .A1(n8037), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5237) );
  NAND4_X1 U6658 ( .A1(n5240), .A2(n5239), .A3(n5238), .A4(n5237), .ZN(n8372)
         );
  AND2_X1 U6659 ( .A1(n8372), .A2(n5513), .ZN(n5242) );
  NAND2_X1 U6660 ( .A1(n5241), .A2(n5242), .ZN(n5246) );
  INV_X1 U6661 ( .A(n5241), .ZN(n5244) );
  INV_X1 U6662 ( .A(n5242), .ZN(n5243) );
  NAND2_X1 U6663 ( .A1(n5244), .A2(n5243), .ZN(n5245) );
  AND2_X1 U6664 ( .A1(n5246), .A2(n5245), .ZN(n7714) );
  INV_X1 U6665 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6737) );
  INV_X1 U6666 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6738) );
  XNOR2_X1 U6667 ( .A(n5272), .B(n5267), .ZN(n6736) );
  NAND2_X1 U6668 ( .A1(n6736), .A2(n8171), .ZN(n5255) );
  NAND2_X1 U6669 ( .A1(n5252), .A2(n5251), .ZN(n5253) );
  NAND2_X1 U6670 ( .A1(n5253), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5303) );
  XNOR2_X1 U6671 ( .A(n5303), .B(P2_IR_REG_14__SCAN_IN), .ZN(n8493) );
  AOI22_X1 U6672 ( .A1(n8014), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6694), .B2(
        n8493), .ZN(n5254) );
  XNOR2_X1 U6673 ( .A(n8925), .B(n4986), .ZN(n5265) );
  NAND2_X1 U6674 ( .A1(n4320), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n5262) );
  NAND2_X1 U6675 ( .A1(n8036), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n5261) );
  INV_X1 U6676 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n10059) );
  NAND2_X1 U6677 ( .A1(n5257), .A2(n10059), .ZN(n5258) );
  AND2_X1 U6678 ( .A1(n5295), .A2(n5258), .ZN(n7817) );
  NAND2_X1 U6679 ( .A1(n5020), .A2(n7817), .ZN(n5260) );
  NAND2_X1 U6680 ( .A1(n8037), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5259) );
  NAND4_X1 U6681 ( .A1(n5262), .A2(n5261), .A3(n5260), .A4(n5259), .ZN(n8802)
         );
  NAND2_X1 U6682 ( .A1(n8802), .A2(n5513), .ZN(n5264) );
  XNOR2_X1 U6683 ( .A(n5265), .B(n5264), .ZN(n7816) );
  NAND2_X1 U6684 ( .A1(n5265), .A2(n5264), .ZN(n5266) );
  INV_X1 U6685 ( .A(n5268), .ZN(n5269) );
  NAND2_X1 U6686 ( .A1(n5269), .A2(SI_14_), .ZN(n5270) );
  INV_X1 U6687 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6829) );
  INV_X1 U6688 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6830) );
  MUX2_X1 U6689 ( .A(n6829), .B(n6830), .S(n4994), .Z(n5274) );
  INV_X1 U6690 ( .A(SI_15_), .ZN(n5273) );
  INV_X1 U6691 ( .A(n5274), .ZN(n5275) );
  NAND2_X1 U6692 ( .A1(n5275), .A2(SI_15_), .ZN(n5276) );
  NAND2_X1 U6693 ( .A1(n5277), .A2(n5276), .ZN(n5300) );
  INV_X1 U6694 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n6968) );
  INV_X1 U6695 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n6970) );
  INV_X1 U6696 ( .A(SI_16_), .ZN(n5278) );
  NAND2_X1 U6697 ( .A1(n5279), .A2(n5278), .ZN(n5319) );
  INV_X1 U6698 ( .A(n5279), .ZN(n5280) );
  NAND2_X1 U6699 ( .A1(n5280), .A2(SI_16_), .ZN(n5281) );
  XNOR2_X1 U6700 ( .A(n5318), .B(n5317), .ZN(n6967) );
  NAND2_X1 U6701 ( .A1(n6967), .A2(n8171), .ZN(n5286) );
  MUX2_X1 U6702 ( .A(n8962), .B(n5282), .S(P2_IR_REG_16__SCAN_IN), .Z(n5284)
         );
  OR2_X1 U6703 ( .A1(n5284), .A2(n5283), .ZN(n8523) );
  INV_X1 U6704 ( .A(n8523), .ZN(n8535) );
  AOI22_X1 U6705 ( .A1(n8014), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6694), .B2(
        n8535), .ZN(n5285) );
  XNOR2_X1 U6706 ( .A(n8783), .B(n5115), .ZN(n8096) );
  NAND2_X1 U6707 ( .A1(n4320), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n5294) );
  NAND2_X1 U6708 ( .A1(n8036), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n5293) );
  INV_X1 U6709 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n8158) );
  INV_X1 U6710 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n5287) );
  OAI21_X1 U6711 ( .B1(n5295), .B2(n8158), .A(n5287), .ZN(n5290) );
  AND2_X1 U6712 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_REG3_REG_15__SCAN_IN), 
        .ZN(n5288) );
  AND2_X1 U6713 ( .A1(n5290), .A2(n5327), .ZN(n8784) );
  NAND2_X1 U6714 ( .A1(n5020), .A2(n8784), .ZN(n5292) );
  NAND2_X1 U6715 ( .A1(n8037), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5291) );
  NAND4_X1 U6716 ( .A1(n5294), .A2(n5293), .A3(n5292), .A4(n5291), .ZN(n8801)
         );
  AND2_X1 U6717 ( .A1(n8801), .A2(n5513), .ZN(n5310) );
  NAND2_X1 U6718 ( .A1(n8035), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n5299) );
  NAND2_X1 U6719 ( .A1(n8036), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n5298) );
  XNOR2_X1 U6720 ( .A(n5295), .B(P2_REG3_REG_15__SCAN_IN), .ZN(n8797) );
  NAND2_X1 U6721 ( .A1(n5020), .A2(n8797), .ZN(n5297) );
  NAND2_X1 U6722 ( .A1(n8037), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5296) );
  NAND4_X1 U6723 ( .A1(n5299), .A2(n5298), .A3(n5297), .A4(n5296), .ZN(n8773)
         );
  AND2_X1 U6724 ( .A1(n8773), .A2(n5513), .ZN(n8156) );
  XNOR2_X1 U6725 ( .A(n5301), .B(n5300), .ZN(n6828) );
  NAND2_X1 U6726 ( .A1(n6828), .A2(n8171), .ZN(n5307) );
  INV_X1 U6727 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5302) );
  NAND2_X1 U6728 ( .A1(n5303), .A2(n5302), .ZN(n5304) );
  NAND2_X1 U6729 ( .A1(n5304), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5305) );
  XNOR2_X1 U6730 ( .A(n5305), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8513) );
  AOI22_X1 U6731 ( .A1(n6694), .A2(n8513), .B1(n8014), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n5306) );
  XNOR2_X1 U6732 ( .A(n8918), .B(n5115), .ZN(n5309) );
  AOI22_X1 U6733 ( .A1(n8096), .A2(n5310), .B1(n8156), .B2(n5309), .ZN(n5308)
         );
  INV_X1 U6734 ( .A(n8096), .ZN(n5314) );
  OAI21_X1 U6735 ( .B1(n5309), .B2(n8156), .A(n5310), .ZN(n5313) );
  INV_X1 U6736 ( .A(n5309), .ZN(n8094) );
  INV_X1 U6737 ( .A(n8156), .ZN(n5311) );
  INV_X1 U6738 ( .A(n5310), .ZN(n8095) );
  AND2_X1 U6739 ( .A1(n5311), .A2(n8095), .ZN(n5312) );
  AOI22_X1 U6740 ( .A1(n5314), .A2(n5313), .B1(n8094), .B2(n5312), .ZN(n5315)
         );
  INV_X1 U6741 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6984) );
  INV_X1 U6742 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n5320) );
  MUX2_X1 U6743 ( .A(n6984), .B(n5320), .S(n4994), .Z(n5341) );
  XNOR2_X1 U6744 ( .A(n5341), .B(SI_17_), .ZN(n5340) );
  XNOR2_X1 U6745 ( .A(n5344), .B(n5340), .ZN(n6956) );
  NAND2_X1 U6746 ( .A1(n6956), .A2(n8171), .ZN(n5326) );
  NAND2_X1 U6747 ( .A1(n5321), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5322) );
  MUX2_X1 U6748 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5322), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n5324) );
  AND2_X1 U6749 ( .A1(n5324), .A2(n5323), .ZN(n8549) );
  AOI22_X1 U6750 ( .A1(n8014), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6694), .B2(
        n8549), .ZN(n5325) );
  XNOR2_X1 U6751 ( .A(n8905), .B(n5115), .ZN(n5333) );
  NAND2_X1 U6752 ( .A1(n4320), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n5332) );
  NAND2_X1 U6753 ( .A1(n8036), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n5331) );
  INV_X1 U6754 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8533) );
  NAND2_X1 U6755 ( .A1(n5327), .A2(n8533), .ZN(n5328) );
  AND2_X1 U6756 ( .A1(n5350), .A2(n5328), .ZN(n8748) );
  NAND2_X1 U6757 ( .A1(n5020), .A2(n8748), .ZN(n5330) );
  NAND2_X1 U6758 ( .A1(n8037), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5329) );
  NAND4_X1 U6759 ( .A1(n5332), .A2(n5331), .A3(n5330), .A4(n5329), .ZN(n8774)
         );
  AND2_X1 U6760 ( .A1(n8774), .A2(n5513), .ZN(n5334) );
  NAND2_X1 U6761 ( .A1(n5333), .A2(n5334), .ZN(n5339) );
  INV_X1 U6762 ( .A(n5333), .ZN(n5336) );
  INV_X1 U6763 ( .A(n5334), .ZN(n5335) );
  NAND2_X1 U6764 ( .A1(n5336), .A2(n5335), .ZN(n5337) );
  NAND2_X1 U6765 ( .A1(n5339), .A2(n5337), .ZN(n8105) );
  INV_X1 U6766 ( .A(n5340), .ZN(n5343) );
  INV_X1 U6767 ( .A(n5341), .ZN(n5342) );
  XNOR2_X1 U6768 ( .A(n5364), .B(SI_18_), .ZN(n5362) );
  XNOR2_X1 U6769 ( .A(n5363), .B(n5362), .ZN(n7088) );
  NAND2_X1 U6770 ( .A1(n7088), .A2(n8171), .ZN(n5347) );
  NAND2_X1 U6771 ( .A1(n5323), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5345) );
  XNOR2_X1 U6772 ( .A(n5345), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8560) );
  AOI22_X1 U6773 ( .A1(n8014), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6694), .B2(
        n8560), .ZN(n5346) );
  XNOR2_X1 U6774 ( .A(n8899), .B(n5115), .ZN(n5356) );
  NAND2_X1 U6775 ( .A1(n8035), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n5355) );
  INV_X1 U6776 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n5349) );
  NAND2_X1 U6777 ( .A1(n5350), .A2(n5349), .ZN(n5351) );
  AND2_X1 U6778 ( .A1(n5373), .A2(n5351), .ZN(n8732) );
  NAND2_X1 U6779 ( .A1(n8732), .A2(n5020), .ZN(n5354) );
  NAND2_X1 U6780 ( .A1(n8036), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n5353) );
  NAND2_X1 U6781 ( .A1(n8037), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n5352) );
  NAND4_X1 U6782 ( .A1(n5355), .A2(n5354), .A3(n5353), .A4(n5352), .ZN(n8371)
         );
  AND2_X1 U6783 ( .A1(n8371), .A2(n5513), .ZN(n5357) );
  NAND2_X1 U6784 ( .A1(n5356), .A2(n5357), .ZN(n5361) );
  INV_X1 U6785 ( .A(n5356), .ZN(n5359) );
  INV_X1 U6786 ( .A(n5357), .ZN(n5358) );
  NAND2_X1 U6787 ( .A1(n5359), .A2(n5358), .ZN(n5360) );
  AND2_X1 U6788 ( .A1(n5361), .A2(n5360), .ZN(n8139) );
  NAND2_X1 U6789 ( .A1(n5364), .A2(SI_18_), .ZN(n5365) );
  INV_X1 U6790 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7131) );
  INV_X1 U6791 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7129) );
  INV_X1 U6792 ( .A(SI_19_), .ZN(n5366) );
  NAND2_X1 U6793 ( .A1(n5367), .A2(n5366), .ZN(n5386) );
  INV_X1 U6794 ( .A(n5367), .ZN(n5368) );
  NAND2_X1 U6795 ( .A1(n5368), .A2(SI_19_), .ZN(n5369) );
  NAND2_X1 U6796 ( .A1(n5386), .A2(n5369), .ZN(n5384) );
  XNOR2_X1 U6797 ( .A(n5383), .B(n5384), .ZN(n7128) );
  NAND2_X1 U6798 ( .A1(n7128), .A2(n8171), .ZN(n5371) );
  AOI22_X1 U6799 ( .A1(n8014), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n6694), .B2(
        n8356), .ZN(n5370) );
  XNOR2_X1 U6800 ( .A(n8896), .B(n4986), .ZN(n5381) );
  INV_X1 U6801 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n5372) );
  NAND2_X1 U6802 ( .A1(n5373), .A2(n5372), .ZN(n5374) );
  NAND2_X1 U6803 ( .A1(n5396), .A2(n5374), .ZN(n8067) );
  NAND2_X1 U6804 ( .A1(n8035), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n5376) );
  NAND2_X1 U6805 ( .A1(n8036), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n5375) );
  AND2_X1 U6806 ( .A1(n5376), .A2(n5375), .ZN(n5378) );
  NAND2_X1 U6807 ( .A1(n8037), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5377) );
  OAI211_X1 U6808 ( .C1(n8067), .C2(n5627), .A(n5378), .B(n5377), .ZN(n8739)
         );
  NAND2_X1 U6809 ( .A1(n8739), .A2(n5513), .ZN(n5380) );
  XNOR2_X1 U6810 ( .A(n5381), .B(n5380), .ZN(n8066) );
  INV_X1 U6811 ( .A(n8066), .ZN(n5379) );
  NAND2_X1 U6812 ( .A1(n5381), .A2(n5380), .ZN(n5382) );
  INV_X1 U6813 ( .A(n5384), .ZN(n5385) );
  NAND2_X1 U6814 ( .A1(n5387), .A2(n5386), .ZN(n5408) );
  INV_X1 U6815 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7288) );
  INV_X1 U6816 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7934) );
  MUX2_X1 U6817 ( .A(n7288), .B(n7934), .S(n4994), .Z(n5389) );
  INV_X1 U6818 ( .A(SI_20_), .ZN(n5388) );
  NAND2_X1 U6819 ( .A1(n5389), .A2(n5388), .ZN(n5409) );
  INV_X1 U6820 ( .A(n5389), .ZN(n5390) );
  NAND2_X1 U6821 ( .A1(n5390), .A2(SI_20_), .ZN(n5391) );
  XNOR2_X1 U6822 ( .A(n5408), .B(n5407), .ZN(n7287) );
  NAND2_X1 U6823 ( .A1(n7287), .A2(n8171), .ZN(n5393) );
  NAND2_X1 U6824 ( .A1(n8014), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n5392) );
  XNOR2_X1 U6825 ( .A(n8889), .B(n5115), .ZN(n5401) );
  INV_X1 U6826 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n5400) );
  INV_X1 U6827 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n5395) );
  NAND2_X1 U6828 ( .A1(n5396), .A2(n5395), .ZN(n5397) );
  NAND2_X1 U6829 ( .A1(n5413), .A2(n5397), .ZN(n8123) );
  OR2_X1 U6830 ( .A1(n8123), .A2(n5627), .ZN(n5399) );
  AOI22_X1 U6831 ( .A1(n4321), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8036), .B2(
        P2_REG1_REG_20__SCAN_IN), .ZN(n5398) );
  OAI211_X1 U6832 ( .C1(n5418), .C2(n5400), .A(n5399), .B(n5398), .ZN(n8698)
         );
  AND2_X1 U6833 ( .A1(n8698), .A2(n5513), .ZN(n5402) );
  NAND2_X1 U6834 ( .A1(n5401), .A2(n5402), .ZN(n5406) );
  INV_X1 U6835 ( .A(n5401), .ZN(n5404) );
  INV_X1 U6836 ( .A(n5402), .ZN(n5403) );
  NAND2_X1 U6837 ( .A1(n5404), .A2(n5403), .ZN(n5405) );
  NAND2_X1 U6838 ( .A1(n5406), .A2(n5405), .ZN(n8119) );
  NAND2_X1 U6839 ( .A1(n8121), .A2(n5406), .ZN(n8075) );
  NAND2_X1 U6840 ( .A1(n5408), .A2(n5407), .ZN(n5410) );
  NAND2_X1 U6841 ( .A1(n5410), .A2(n5409), .ZN(n5428) );
  INV_X1 U6842 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7351) );
  INV_X1 U6843 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7341) );
  XNOR2_X1 U6844 ( .A(n5424), .B(SI_21_), .ZN(n5423) );
  XNOR2_X1 U6845 ( .A(n5428), .B(n5423), .ZN(n7340) );
  NAND2_X1 U6846 ( .A1(n7340), .A2(n8171), .ZN(n5412) );
  NAND2_X1 U6847 ( .A1(n8014), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n5411) );
  XNOR2_X1 U6848 ( .A(n8884), .B(n5115), .ZN(n5421) );
  INV_X1 U6849 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n5417) );
  INV_X1 U6850 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n8076) );
  NAND2_X1 U6851 ( .A1(n5413), .A2(n8076), .ZN(n5414) );
  NAND2_X1 U6852 ( .A1(n5435), .A2(n5414), .ZN(n8689) );
  OR2_X1 U6853 ( .A1(n8689), .A2(n5627), .ZN(n5416) );
  AOI22_X1 U6854 ( .A1(n8035), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8036), .B2(
        P2_REG1_REG_21__SCAN_IN), .ZN(n5415) );
  OAI211_X1 U6855 ( .C1(n5418), .C2(n5417), .A(n5416), .B(n5415), .ZN(n8711)
         );
  NAND2_X1 U6856 ( .A1(n8711), .A2(n5513), .ZN(n5419) );
  XNOR2_X1 U6857 ( .A(n5421), .B(n5419), .ZN(n8074) );
  NAND2_X1 U6858 ( .A1(n8075), .A2(n8074), .ZN(n8073) );
  INV_X1 U6859 ( .A(n5419), .ZN(n5420) );
  NAND2_X1 U6860 ( .A1(n5421), .A2(n5420), .ZN(n5422) );
  INV_X1 U6861 ( .A(n5423), .ZN(n5427) );
  INV_X1 U6862 ( .A(n5424), .ZN(n5425) );
  NAND2_X1 U6863 ( .A1(n5425), .A2(SI_21_), .ZN(n5426) );
  INV_X1 U6864 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7989) );
  INV_X1 U6865 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n10076) );
  INV_X1 U6866 ( .A(SI_22_), .ZN(n5429) );
  NAND2_X1 U6867 ( .A1(n5430), .A2(n5429), .ZN(n5450) );
  INV_X1 U6868 ( .A(n5430), .ZN(n5431) );
  NAND2_X1 U6869 ( .A1(n5431), .A2(SI_22_), .ZN(n5432) );
  NAND2_X1 U6870 ( .A1(n5450), .A2(n5432), .ZN(n5448) );
  XNOR2_X1 U6871 ( .A(n5449), .B(n5448), .ZN(n7676) );
  NAND2_X1 U6872 ( .A1(n7676), .A2(n8171), .ZN(n5434) );
  NAND2_X1 U6873 ( .A1(n8014), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n5433) );
  XNOR2_X1 U6874 ( .A(n8879), .B(n4986), .ZN(n5443) );
  INV_X1 U6875 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n8131) );
  NAND2_X1 U6876 ( .A1(n5435), .A2(n8131), .ZN(n5436) );
  AND2_X1 U6877 ( .A1(n5476), .A2(n5436), .ZN(n8672) );
  NAND2_X1 U6878 ( .A1(n8672), .A2(n5020), .ZN(n5442) );
  INV_X1 U6879 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n5439) );
  NAND2_X1 U6880 ( .A1(n8035), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n5438) );
  NAND2_X1 U6881 ( .A1(n8036), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n5437) );
  OAI211_X1 U6882 ( .C1(n5439), .C2(n5418), .A(n5438), .B(n5437), .ZN(n5440)
         );
  INV_X1 U6883 ( .A(n5440), .ZN(n5441) );
  NAND2_X1 U6884 ( .A1(n5442), .A2(n5441), .ZN(n8699) );
  NAND2_X1 U6885 ( .A1(n8699), .A2(n5513), .ZN(n8130) );
  NAND2_X1 U6886 ( .A1(n8129), .A2(n8130), .ZN(n5447) );
  INV_X1 U6887 ( .A(n5443), .ZN(n5444) );
  OR2_X1 U6888 ( .A1(n5445), .A2(n5444), .ZN(n5446) );
  NAND2_X2 U6889 ( .A1(n5447), .A2(n5446), .ZN(n5485) );
  INV_X1 U6890 ( .A(n5460), .ZN(n5457) );
  INV_X1 U6891 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n5452) );
  INV_X1 U6892 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n5451) );
  INV_X1 U6893 ( .A(SI_23_), .ZN(n5453) );
  NAND2_X1 U6894 ( .A1(n5454), .A2(n5453), .ZN(n5464) );
  INV_X1 U6895 ( .A(n5454), .ZN(n5455) );
  NAND2_X1 U6896 ( .A1(n5455), .A2(SI_23_), .ZN(n5456) );
  NAND2_X1 U6897 ( .A1(n5464), .A2(n5456), .ZN(n5458) );
  NAND2_X1 U6898 ( .A1(n5457), .A2(n5458), .ZN(n5461) );
  INV_X1 U6899 ( .A(n5458), .ZN(n5459) );
  NAND2_X1 U6900 ( .A1(n5461), .A2(n5465), .ZN(n7677) );
  NAND2_X1 U6901 ( .A1(n7677), .A2(n8171), .ZN(n5463) );
  NAND2_X1 U6902 ( .A1(n8014), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n5462) );
  XNOR2_X1 U6903 ( .A(n8873), .B(n5115), .ZN(n5486) );
  INV_X1 U6904 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n5466) );
  INV_X1 U6905 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n10055) );
  MUX2_X1 U6906 ( .A(n5466), .B(n10055), .S(n4994), .Z(n5493) );
  XNOR2_X1 U6907 ( .A(n5493), .B(SI_24_), .ZN(n5492) );
  NAND2_X1 U6908 ( .A1(n7769), .A2(n8171), .ZN(n5468) );
  NAND2_X1 U6909 ( .A1(n8014), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n5467) );
  XNOR2_X1 U6910 ( .A(n8867), .B(n4986), .ZN(n8113) );
  XNOR2_X1 U6911 ( .A(n5505), .B(P2_REG3_REG_24__SCAN_IN), .ZN(n8638) );
  NAND2_X1 U6912 ( .A1(n8638), .A2(n5020), .ZN(n5475) );
  INV_X1 U6913 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n5472) );
  NAND2_X1 U6914 ( .A1(n8035), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n5471) );
  NAND2_X1 U6915 ( .A1(n8036), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n5470) );
  OAI211_X1 U6916 ( .C1(n5472), .C2(n5418), .A(n5471), .B(n5470), .ZN(n5473)
         );
  INV_X1 U6917 ( .A(n5473), .ZN(n5474) );
  INV_X1 U6918 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8058) );
  NAND2_X1 U6919 ( .A1(n5476), .A2(n8058), .ZN(n5477) );
  NAND2_X1 U6920 ( .A1(n5505), .A2(n5477), .ZN(n8660) );
  OR2_X1 U6921 ( .A1(n8660), .A2(n5627), .ZN(n5483) );
  INV_X1 U6922 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n5480) );
  NAND2_X1 U6923 ( .A1(n4321), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n5479) );
  NAND2_X1 U6924 ( .A1(n8036), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n5478) );
  OAI211_X1 U6925 ( .C1(n5480), .C2(n5418), .A(n5479), .B(n5478), .ZN(n5481)
         );
  INV_X1 U6926 ( .A(n5481), .ZN(n5482) );
  NAND2_X1 U6927 ( .A1(n5483), .A2(n5482), .ZN(n8645) );
  NAND2_X1 U6928 ( .A1(n8645), .A2(n5513), .ZN(n8055) );
  AOI21_X1 U6929 ( .B1(n8113), .B2(n8088), .A(n8055), .ZN(n5484) );
  INV_X1 U6930 ( .A(n5485), .ZN(n5487) );
  NAND2_X1 U6931 ( .A1(n8653), .A2(n5513), .ZN(n8115) );
  NAND2_X1 U6932 ( .A1(n8113), .A2(n8115), .ZN(n5488) );
  NAND2_X1 U6933 ( .A1(n8111), .A2(n5488), .ZN(n5490) );
  INV_X1 U6934 ( .A(n5493), .ZN(n5494) );
  NAND2_X1 U6935 ( .A1(n5494), .A2(SI_24_), .ZN(n5495) );
  INV_X1 U6936 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n5497) );
  INV_X1 U6937 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7826) );
  INV_X1 U6938 ( .A(SI_25_), .ZN(n5498) );
  NAND2_X1 U6939 ( .A1(n5499), .A2(n5498), .ZN(n5520) );
  INV_X1 U6940 ( .A(n5499), .ZN(n5500) );
  NAND2_X1 U6941 ( .A1(n5500), .A2(SI_25_), .ZN(n5501) );
  NAND2_X1 U6942 ( .A1(n5520), .A2(n5501), .ZN(n5518) );
  NAND2_X1 U6943 ( .A1(n8014), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n5502) );
  XNOR2_X1 U6944 ( .A(n8863), .B(n5115), .ZN(n5514) );
  INV_X1 U6945 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n5504) );
  INV_X1 U6946 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8086) );
  OAI21_X1 U6947 ( .B1(n5505), .B2(n5504), .A(n8086), .ZN(n5506) );
  NAND2_X1 U6948 ( .A1(n5506), .A2(n5528), .ZN(n8624) );
  OR2_X1 U6949 ( .A1(n8624), .A2(n5627), .ZN(n5512) );
  INV_X1 U6950 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n5509) );
  NAND2_X1 U6951 ( .A1(n8036), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n5508) );
  NAND2_X1 U6952 ( .A1(n4321), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n5507) );
  OAI211_X1 U6953 ( .C1(n5418), .C2(n5509), .A(n5508), .B(n5507), .ZN(n5510)
         );
  INV_X1 U6954 ( .A(n5510), .ZN(n5511) );
  NAND2_X1 U6955 ( .A1(n5512), .A2(n5511), .ZN(n8646) );
  AND2_X1 U6956 ( .A1(n8646), .A2(n5513), .ZN(n5515) );
  AND2_X1 U6957 ( .A1(n5514), .A2(n5515), .ZN(n8083) );
  INV_X1 U6958 ( .A(n5514), .ZN(n5517) );
  INV_X1 U6959 ( .A(n5515), .ZN(n5516) );
  NAND2_X1 U6960 ( .A1(n5517), .A2(n5516), .ZN(n8082) );
  INV_X1 U6961 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7889) );
  INV_X1 U6962 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7931) );
  INV_X1 U6963 ( .A(SI_26_), .ZN(n5521) );
  NAND2_X1 U6964 ( .A1(n5522), .A2(n5521), .ZN(n5543) );
  INV_X1 U6965 ( .A(n5522), .ZN(n5523) );
  NAND2_X1 U6966 ( .A1(n5523), .A2(SI_26_), .ZN(n5524) );
  NAND2_X1 U6967 ( .A1(n7888), .A2(n8171), .ZN(n5526) );
  NAND2_X1 U6968 ( .A1(n8014), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n5525) );
  XNOR2_X1 U6969 ( .A(n8858), .B(n4986), .ZN(n5536) );
  INV_X1 U6970 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n9941) );
  NAND2_X1 U6971 ( .A1(n5528), .A2(n9941), .ZN(n5529) );
  NAND2_X1 U6972 ( .A1(n5564), .A2(n5529), .ZN(n8609) );
  INV_X1 U6973 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n5532) );
  NAND2_X1 U6974 ( .A1(n8036), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n5531) );
  NAND2_X1 U6975 ( .A1(n8037), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n5530) );
  OAI211_X1 U6976 ( .C1(n4322), .C2(n5532), .A(n5531), .B(n5530), .ZN(n5533)
         );
  INV_X1 U6977 ( .A(n5533), .ZN(n5534) );
  NAND2_X1 U6978 ( .A1(n8630), .A2(n5513), .ZN(n5537) );
  XNOR2_X1 U6979 ( .A(n5536), .B(n5537), .ZN(n8148) );
  INV_X1 U6980 ( .A(n5536), .ZN(n5539) );
  INV_X1 U6981 ( .A(n5537), .ZN(n5538) );
  NAND2_X1 U6982 ( .A1(n5539), .A2(n5538), .ZN(n5540) );
  INV_X1 U6983 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n7928) );
  INV_X1 U6984 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n5544) );
  INV_X1 U6985 ( .A(SI_27_), .ZN(n5545) );
  NAND2_X1 U6986 ( .A1(n5546), .A2(n5545), .ZN(n5605) );
  INV_X1 U6987 ( .A(n5546), .ZN(n5547) );
  NAND2_X1 U6988 ( .A1(n5547), .A2(SI_27_), .ZN(n5548) );
  AND2_X1 U6989 ( .A1(n5605), .A2(n5548), .ZN(n5603) );
  NAND2_X1 U6990 ( .A1(n7891), .A2(n8171), .ZN(n5550) );
  NAND2_X1 U6991 ( .A1(n8014), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n5549) );
  XNOR2_X1 U6992 ( .A(n8852), .B(n5115), .ZN(n5559) );
  XNOR2_X1 U6993 ( .A(n5564), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n8597) );
  NAND2_X1 U6994 ( .A1(n8597), .A2(n4323), .ZN(n5556) );
  INV_X1 U6995 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n5553) );
  NAND2_X1 U6996 ( .A1(n4321), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n5552) );
  NAND2_X1 U6997 ( .A1(n8036), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n5551) );
  OAI211_X1 U6998 ( .C1(n5553), .C2(n5418), .A(n5552), .B(n5551), .ZN(n5554)
         );
  INV_X1 U6999 ( .A(n5554), .ZN(n5555) );
  NAND2_X1 U7000 ( .A1(n8615), .A2(n5513), .ZN(n5557) );
  XNOR2_X1 U7001 ( .A(n5559), .B(n5557), .ZN(n8046) );
  INV_X1 U7002 ( .A(n5557), .ZN(n5558) );
  NAND2_X1 U7003 ( .A1(n5559), .A2(n5558), .ZN(n5560) );
  NAND2_X1 U7004 ( .A1(n5561), .A2(n5560), .ZN(n5574) );
  INV_X1 U7005 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n8047) );
  INV_X1 U7006 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n5562) );
  OAI21_X1 U7007 ( .B1(n5564), .B2(n8047), .A(n5562), .ZN(n5565) );
  NAND2_X1 U7008 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .ZN(n5563) );
  NAND2_X1 U7009 ( .A1(n8586), .A2(n4323), .ZN(n5571) );
  INV_X1 U7010 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n5568) );
  NAND2_X1 U7011 ( .A1(n8035), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n5567) );
  NAND2_X1 U7012 ( .A1(n8036), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n5566) );
  OAI211_X1 U7013 ( .C1(n5568), .C2(n5418), .A(n5567), .B(n5566), .ZN(n5569)
         );
  INV_X1 U7014 ( .A(n5569), .ZN(n5570) );
  NAND2_X1 U7015 ( .A1(n5571), .A2(n5570), .ZN(n8601) );
  NAND2_X1 U7016 ( .A1(n8601), .A2(n5513), .ZN(n5572) );
  XNOR2_X1 U7017 ( .A(n5572), .B(n4986), .ZN(n5573) );
  NOR4_X1 U7018 ( .A1(P2_D_REG_5__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n5583) );
  INV_X1 U7019 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n10022) );
  INV_X1 U7020 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n9760) );
  INV_X1 U7021 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n10056) );
  INV_X1 U7022 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n10047) );
  NAND4_X1 U7023 ( .A1(n10022), .A2(n9760), .A3(n10056), .A4(n10047), .ZN(
        n5580) );
  NOR4_X1 U7024 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_19__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n5578) );
  NOR4_X1 U7025 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_12__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n5577) );
  NOR4_X1 U7026 ( .A1(P2_D_REG_25__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n5576) );
  NOR4_X1 U7027 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_23__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n5575) );
  NAND4_X1 U7028 ( .A1(n5578), .A2(n5577), .A3(n5576), .A4(n5575), .ZN(n5579)
         );
  NOR4_X1 U7029 ( .A1(P2_D_REG_28__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        n5580), .A4(n5579), .ZN(n5582) );
  NOR4_X1 U7030 ( .A1(P2_D_REG_3__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_2__SCAN_IN), .A4(P2_D_REG_4__SCAN_IN), .ZN(n5581) );
  NAND3_X1 U7031 ( .A1(n5583), .A2(n5582), .A3(n5581), .ZN(n5596) );
  NAND2_X1 U7032 ( .A1(n5584), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5585) );
  XNOR2_X1 U7033 ( .A(n5585), .B(P2_IR_REG_26__SCAN_IN), .ZN(n5599) );
  NAND2_X1 U7034 ( .A1(n5586), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5587) );
  XNOR2_X1 U7035 ( .A(n5587), .B(P2_IR_REG_25__SCAN_IN), .ZN(n7824) );
  NAND2_X1 U7036 ( .A1(n5589), .A2(n5588), .ZN(n5590) );
  NAND2_X1 U7037 ( .A1(n5590), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5600) );
  NAND2_X1 U7038 ( .A1(n5600), .A2(n5591), .ZN(n5592) );
  NAND2_X1 U7039 ( .A1(n5592), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5593) );
  XOR2_X1 U7040 ( .A(P2_B_REG_SCAN_IN), .B(n6540), .Z(n5594) );
  AND2_X1 U7041 ( .A1(n5596), .A2(n9758), .ZN(n6810) );
  INV_X1 U7042 ( .A(n5599), .ZN(n7890) );
  AND2_X1 U7043 ( .A1(n6540), .A2(n7890), .ZN(n9764) );
  INV_X1 U7044 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n9763) );
  AND2_X1 U7045 ( .A1(n9758), .A2(n9763), .ZN(n5597) );
  NOR2_X1 U7046 ( .A1(n6810), .A2(n7272), .ZN(n5598) );
  INV_X1 U7047 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n9766) );
  NOR2_X1 U7048 ( .A1(n5599), .A2(n7824), .ZN(n9768) );
  AOI21_X1 U7049 ( .B1(n9758), .B2(n9766), .A(n9768), .ZN(n7037) );
  NAND2_X1 U7050 ( .A1(n5598), .A2(n7037), .ZN(n5617) );
  AND2_X2 U7051 ( .A1(n4702), .A2(n8363), .ZN(n9802) );
  NAND2_X1 U7052 ( .A1(n5599), .A2(n7824), .ZN(n6541) );
  OR2_X1 U7053 ( .A1(n6540), .A2(n6541), .ZN(n5602) );
  XNOR2_X1 U7054 ( .A(n5600), .B(P2_IR_REG_23__SCAN_IN), .ZN(n9762) );
  INV_X1 U7055 ( .A(n9762), .ZN(n5601) );
  NAND2_X1 U7056 ( .A1(n5602), .A2(n5601), .ZN(n5615) );
  INV_X1 U7057 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n9988) );
  INV_X1 U7058 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n9511) );
  XNOR2_X1 U7059 ( .A(n6269), .B(SI_28_), .ZN(n6266) );
  NAND2_X1 U7060 ( .A1(n7926), .A2(n8171), .ZN(n5608) );
  NAND2_X1 U7061 ( .A1(n8014), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n5607) );
  INV_X1 U7062 ( .A(n9759), .ZN(n5609) );
  NOR2_X1 U7063 ( .A1(n5610), .A2(n8343), .ZN(n7044) );
  NAND2_X1 U7064 ( .A1(n5609), .A2(n7044), .ZN(n5611) );
  OAI21_X2 U7065 ( .B1(n5617), .B2(n5611), .A(n7668), .ZN(n8166) );
  INV_X1 U7066 ( .A(n4315), .ZN(n5614) );
  AND2_X1 U7067 ( .A1(n6860), .A2(n8363), .ZN(n6811) );
  AOI211_X1 U7068 ( .C1(n5617), .C2(n6814), .A(n6811), .B(n5615), .ZN(n6910)
         );
  INV_X1 U7069 ( .A(n5617), .ZN(n5619) );
  NOR2_X1 U7070 ( .A1(n9759), .A2(n8363), .ZN(n5618) );
  NAND2_X1 U7071 ( .A1(n5619), .A2(n5618), .ZN(n8068) );
  INV_X1 U7072 ( .A(n6860), .ZN(n6696) );
  INV_X1 U7073 ( .A(n5620), .ZN(n5621) );
  INV_X1 U7074 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n9983) );
  NAND2_X1 U7075 ( .A1(n4321), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n5623) );
  NAND2_X1 U7076 ( .A1(n8037), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n5622) );
  OAI211_X1 U7077 ( .C1(n5624), .C2(n9983), .A(n5623), .B(n5622), .ZN(n5625)
         );
  INV_X1 U7078 ( .A(n5625), .ZN(n5626) );
  OAI21_X1 U7079 ( .B1(n8019), .B2(n5627), .A(n5626), .ZN(n8590) );
  AOI22_X1 U7080 ( .A1(n5616), .A2(n8586), .B1(n8143), .B2(n8590), .ZN(n5629)
         );
  OR2_X1 U7081 ( .A1(n6696), .A2(n5620), .ZN(n8756) );
  NOR2_X1 U7082 ( .A1(n8068), .A2(n8756), .ZN(n8124) );
  AOI22_X1 U7083 ( .A1(n8124), .A2(n8615), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3152), .ZN(n5628) );
  NAND2_X1 U7084 ( .A1(n5630), .A2(n4897), .ZN(P2_U3222) );
  NAND2_X1 U7085 ( .A1(n5752), .A2(n5631), .ZN(n5784) );
  NOR2_X1 U7086 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n5635) );
  NOR2_X1 U7087 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n5634) );
  NAND2_X1 U7088 ( .A1(n9959), .A2(n5638), .ZN(n5641) );
  NAND2_X1 U7089 ( .A1(n5973), .A2(n5639), .ZN(n5640) );
  INV_X1 U7090 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5643) );
  INV_X1 U7091 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5665) );
  INV_X1 U7092 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5664) );
  INV_X1 U7093 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5661) );
  INV_X1 U7094 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5646) );
  NAND2_X1 U7095 ( .A1(n5650), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5647) );
  MUX2_X1 U7096 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5647), .S(
        P1_IR_REG_28__SCAN_IN), .Z(n5649) );
  INV_X1 U7097 ( .A(n5698), .ZN(n5648) );
  OR2_X1 U7098 ( .A1(n5651), .A2(n9504), .ZN(n5652) );
  NAND2_X1 U7099 ( .A1(n5652), .A2(P1_IR_REG_27__SCAN_IN), .ZN(n5654) );
  NAND2_X1 U7100 ( .A1(n7677), .A2(n5751), .ZN(n5657) );
  NAND2_X1 U7101 ( .A1(n6302), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n5656) );
  NAND2_X1 U7102 ( .A1(n5663), .A2(n5664), .ZN(n5659) );
  NAND2_X1 U7103 ( .A1(n5666), .A2(n5665), .ZN(n5660) );
  NAND2_X1 U7104 ( .A1(n5660), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5662) );
  XNOR2_X1 U7105 ( .A(n5663), .B(n5664), .ZN(n7802) );
  XNOR2_X1 U7106 ( .A(n5666), .B(n5665), .ZN(n7828) );
  NAND2_X1 U7107 ( .A1(n6003), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6021) );
  NAND2_X1 U7108 ( .A1(n6021), .A2(n5667), .ZN(n5668) );
  INV_X1 U7109 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5680) );
  NAND2_X1 U7110 ( .A1(n5681), .A2(n5680), .ZN(n5683) );
  NAND2_X1 U7111 ( .A1(n5683), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5670) );
  INV_X1 U7112 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5669) );
  INV_X1 U7113 ( .A(n5671), .ZN(n5672) );
  NAND2_X1 U7114 ( .A1(n5672), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5673) );
  INV_X1 U7115 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5674) );
  NAND2_X1 U7116 ( .A1(n4646), .A2(n5674), .ZN(n5678) );
  NAND2_X1 U7117 ( .A1(n5675), .A2(P1_IR_REG_21__SCAN_IN), .ZN(n5676) );
  INV_X1 U7118 ( .A(n6639), .ZN(n5677) );
  OR2_X1 U7119 ( .A1(n5681), .A2(n5680), .ZN(n5682) );
  NAND2_X1 U7120 ( .A1(n5683), .A2(n5682), .ZN(n9682) );
  NAND2_X1 U7121 ( .A1(n7936), .A2(n9682), .ZN(n6527) );
  INV_X1 U7122 ( .A(n6527), .ZN(n5684) );
  AND2_X4 U7123 ( .A1(n6543), .A2(n6639), .ZN(n5755) );
  INV_X1 U7124 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n5884) );
  INV_X1 U7125 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5928) );
  INV_X1 U7126 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5946) );
  OR2_X2 U7127 ( .A1(n5947), .A2(n5946), .ZN(n5960) );
  INV_X1 U7128 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n6006) );
  INV_X1 U7129 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n6042) );
  INV_X1 U7130 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n9054) );
  INV_X1 U7131 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n8989) );
  NAND2_X1 U7132 ( .A1(n6113), .A2(n8989), .ZN(n5695) );
  NAND2_X1 U7133 ( .A1(n6133), .A2(n5695), .ZN(n9294) );
  INV_X1 U7134 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5696) );
  NAND2_X1 U7135 ( .A1(n5698), .A2(n5696), .ZN(n5701) );
  XNOR2_X2 U7136 ( .A(n5697), .B(P1_IR_REG_30__SCAN_IN), .ZN(n5704) );
  OAI21_X1 U7137 ( .B1(n5698), .B2(n9504), .A(P1_IR_REG_29__SCAN_IN), .ZN(
        n5700) );
  INV_X1 U7138 ( .A(n5743), .ZN(n6095) );
  OR2_X1 U7139 ( .A1(n9294), .A2(n6095), .ZN(n5709) );
  INV_X1 U7140 ( .A(n5744), .ZN(n6284) );
  INV_X1 U7141 ( .A(n6284), .ZN(n6246) );
  INV_X1 U7142 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n9973) );
  NAND2_X1 U7143 ( .A1(n4335), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n5706) );
  AND2_X2 U7144 ( .A1(n5704), .A2(n7930), .ZN(n5745) );
  NAND2_X1 U7145 ( .A1(n5745), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n5705) );
  OAI211_X1 U7146 ( .C1(n6246), .C2(n9973), .A(n5706), .B(n5705), .ZN(n5707)
         );
  INV_X1 U7147 ( .A(n5707), .ZN(n5708) );
  NAND2_X1 U7148 ( .A1(n5709), .A2(n5708), .ZN(n9308) );
  AOI22_X1 U7149 ( .A1(n9441), .A2(n6197), .B1(n6179), .B2(n9308), .ZN(n8987)
         );
  NAND2_X1 U7150 ( .A1(n5745), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5714) );
  NAND2_X1 U7151 ( .A1(n4319), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5713) );
  INV_X1 U7152 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n5710) );
  NAND4_X2 U7153 ( .A1(n5714), .A2(n5713), .A3(n5712), .A4(n5711), .ZN(n6306)
         );
  NAND2_X1 U7154 ( .A1(n6306), .A2(n5873), .ZN(n5720) );
  NAND2_X1 U7155 ( .A1(n4994), .A2(SI_0_), .ZN(n5716) );
  INV_X1 U7156 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5715) );
  NAND2_X1 U7157 ( .A1(n5716), .A2(n5715), .ZN(n5718) );
  AND2_X1 U7158 ( .A1(n5718), .A2(n5717), .ZN(n9513) );
  MUX2_X1 U7159 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9513), .S(n5801), .Z(n7109) );
  INV_X1 U7160 ( .A(n6543), .ZN(n6544) );
  AOI22_X1 U7161 ( .A1(n7109), .A2(n5755), .B1(n6544), .B2(
        P1_REG1_REG_0__SCAN_IN), .ZN(n5719) );
  NAND2_X1 U7162 ( .A1(n5720), .A2(n5719), .ZN(n6800) );
  INV_X1 U7163 ( .A(n6800), .ZN(n5722) );
  NAND2_X1 U7164 ( .A1(n6614), .A2(n9682), .ZN(n5721) );
  NAND2_X1 U7165 ( .A1(n5722), .A2(n7304), .ZN(n5727) );
  INV_X1 U7166 ( .A(n6215), .ZN(n5723) );
  NAND2_X1 U7167 ( .A1(n5723), .A2(n6306), .ZN(n5726) );
  NAND2_X1 U7168 ( .A1(n5873), .A2(n7109), .ZN(n5725) );
  NAND2_X1 U7169 ( .A1(n5745), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5731) );
  NAND2_X1 U7170 ( .A1(n4319), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5730) );
  INV_X1 U7171 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6666) );
  NAND2_X1 U7172 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5732) );
  XNOR2_X1 U7173 ( .A(n5732), .B(P1_IR_REG_1__SCAN_IN), .ZN(n6664) );
  NAND2_X1 U7174 ( .A1(n6057), .A2(n6664), .ZN(n5733) );
  NAND2_X1 U7175 ( .A1(n7234), .A2(n5755), .ZN(n5735) );
  NAND2_X1 U7176 ( .A1(n6832), .A2(n6833), .ZN(n5740) );
  NAND2_X1 U7177 ( .A1(n9133), .A2(n6179), .ZN(n5739) );
  NAND2_X1 U7178 ( .A1(n7234), .A2(n5873), .ZN(n5738) );
  NAND2_X1 U7179 ( .A1(n5739), .A2(n5738), .ZN(n6837) );
  NAND2_X1 U7180 ( .A1(n5740), .A2(n6837), .ZN(n6840) );
  INV_X1 U7181 ( .A(n6832), .ZN(n5742) );
  INV_X1 U7182 ( .A(n6833), .ZN(n5741) );
  NAND2_X1 U7183 ( .A1(n5742), .A2(n5741), .ZN(n6836) );
  NAND2_X1 U7184 ( .A1(n6840), .A2(n6836), .ZN(n6945) );
  INV_X1 U7185 ( .A(n6945), .ZN(n5762) );
  NAND2_X1 U7186 ( .A1(n4319), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5748) );
  INV_X1 U7187 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n6973) );
  NAND2_X1 U7188 ( .A1(n5745), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5746) );
  INV_X1 U7189 ( .A(n6671), .ZN(n5750) );
  OR2_X1 U7190 ( .A1(n5752), .A2(n9504), .ZN(n5769) );
  XNOR2_X1 U7191 ( .A(n5769), .B(P1_IR_REG_2__SCAN_IN), .ZN(n6670) );
  OR2_X1 U7192 ( .A1(n5801), .A2(n9608), .ZN(n5753) );
  INV_X2 U7193 ( .A(n6308), .ZN(n6933) );
  OAI22_X1 U7194 ( .A1(n6309), .A2(n6209), .B1(n6933), .B2(n5756), .ZN(n5757)
         );
  XNOR2_X1 U7195 ( .A(n5757), .B(n7304), .ZN(n5759) );
  OAI22_X1 U7196 ( .A1(n6309), .A2(n6215), .B1(n6933), .B2(n6209), .ZN(n5758)
         );
  OR2_X1 U7197 ( .A1(n5759), .A2(n5758), .ZN(n5763) );
  NAND2_X1 U7198 ( .A1(n5759), .A2(n5758), .ZN(n5760) );
  INV_X1 U7199 ( .A(n6946), .ZN(n5761) );
  NAND2_X1 U7200 ( .A1(n5762), .A2(n5761), .ZN(n6947) );
  NAND2_X1 U7201 ( .A1(n6947), .A2(n5763), .ZN(n7057) );
  NAND2_X1 U7202 ( .A1(n4335), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5768) );
  INV_X1 U7203 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n5764) );
  NAND2_X1 U7204 ( .A1(n4319), .A2(n5764), .ZN(n5767) );
  NAND2_X1 U7205 ( .A1(n5745), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5766) );
  NAND2_X1 U7206 ( .A1(n6284), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5765) );
  OR2_X1 U7207 ( .A1(n5838), .A2(n6654), .ZN(n5773) );
  INV_X1 U7208 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n9895) );
  NAND2_X1 U7209 ( .A1(n5769), .A2(n9895), .ZN(n5770) );
  NAND2_X1 U7210 ( .A1(n5770), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5771) );
  XNOR2_X1 U7211 ( .A(n5771), .B(P1_IR_REG_3__SCAN_IN), .ZN(n9150) );
  NAND2_X1 U7212 ( .A1(n6057), .A2(n9150), .ZN(n5772) );
  OAI211_X1 U7213 ( .C1(n6290), .C2(n6655), .A(n5773), .B(n5772), .ZN(n7124)
         );
  INV_X1 U7214 ( .A(n7124), .ZN(n9706) );
  OAI22_X1 U7215 ( .A1(n7134), .A2(n6215), .B1(n9706), .B2(n6209), .ZN(n5776)
         );
  XNOR2_X1 U7216 ( .A(n5775), .B(n5776), .ZN(n7058) );
  NAND2_X1 U7217 ( .A1(n7057), .A2(n7058), .ZN(n7056) );
  INV_X1 U7218 ( .A(n5775), .ZN(n5777) );
  OR2_X1 U7219 ( .A1(n5777), .A2(n5776), .ZN(n5778) );
  NAND2_X1 U7220 ( .A1(n7056), .A2(n5778), .ZN(n7082) );
  NAND2_X1 U7221 ( .A1(n4335), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5783) );
  INV_X1 U7222 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n5779) );
  XNOR2_X1 U7223 ( .A(n5779), .B(P1_REG3_REG_3__SCAN_IN), .ZN(n7174) );
  NAND2_X1 U7224 ( .A1(n5743), .A2(n7174), .ZN(n5782) );
  NAND2_X1 U7225 ( .A1(n6284), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5781) );
  NAND2_X1 U7226 ( .A1(n6283), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5780) );
  OR2_X1 U7227 ( .A1(n5838), .A2(n6662), .ZN(n5787) );
  NAND2_X1 U7228 ( .A1(n5784), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5785) );
  XNOR2_X1 U7229 ( .A(n5785), .B(P1_IR_REG_4__SCAN_IN), .ZN(n6808) );
  NAND2_X1 U7230 ( .A1(n6057), .A2(n6808), .ZN(n5786) );
  OAI211_X1 U7231 ( .C1(n6290), .C2(n6663), .A(n5787), .B(n5786), .ZN(n7144)
         );
  OAI22_X1 U7232 ( .A1(n7262), .A2(n6209), .B1(n7173), .B2(n5756), .ZN(n5788)
         );
  XNOR2_X1 U7233 ( .A(n5788), .B(n7304), .ZN(n5790) );
  OAI22_X1 U7234 ( .A1(n7262), .A2(n6215), .B1(n7173), .B2(n6209), .ZN(n5789)
         );
  NAND2_X1 U7235 ( .A1(n5790), .A2(n5789), .ZN(n7079) );
  NAND2_X1 U7236 ( .A1(n7082), .A2(n7079), .ZN(n5791) );
  OR2_X1 U7237 ( .A1(n5790), .A2(n5789), .ZN(n7080) );
  NAND2_X1 U7238 ( .A1(n4335), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5800) );
  INV_X1 U7239 ( .A(n5792), .ZN(n5794) );
  INV_X1 U7240 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5793) );
  NAND2_X1 U7241 ( .A1(n5794), .A2(n5793), .ZN(n5795) );
  NAND2_X1 U7242 ( .A1(n5811), .A2(n5795), .ZN(n9691) );
  INV_X1 U7243 ( .A(n9691), .ZN(n7265) );
  NAND2_X1 U7244 ( .A1(n5743), .A2(n7265), .ZN(n5799) );
  NAND2_X1 U7245 ( .A1(n6283), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5798) );
  NAND2_X1 U7246 ( .A1(n4317), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5797) );
  NAND2_X1 U7247 ( .A1(n5802), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5803) );
  MUX2_X1 U7248 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5803), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n5805) );
  INV_X1 U7249 ( .A(n6590), .ZN(n6744) );
  OR2_X1 U7250 ( .A1(n5838), .A2(n6653), .ZN(n5807) );
  INV_X1 U7251 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n9957) );
  OR2_X1 U7252 ( .A1(n6290), .A2(n9957), .ZN(n5806) );
  OAI211_X1 U7253 ( .C1(n5801), .C2(n6744), .A(n5807), .B(n5806), .ZN(n9680)
         );
  INV_X1 U7254 ( .A(n9680), .ZN(n6310) );
  OAI22_X1 U7255 ( .A1(n7441), .A2(n6209), .B1(n6310), .B2(n5756), .ZN(n5808)
         );
  XNOR2_X1 U7256 ( .A(n5808), .B(n7304), .ZN(n5825) );
  OR2_X1 U7257 ( .A1(n7441), .A2(n6215), .ZN(n5810) );
  NAND2_X1 U7258 ( .A1(n9680), .A2(n6197), .ZN(n5809) );
  NAND2_X1 U7259 ( .A1(n5810), .A2(n5809), .ZN(n7260) );
  NAND2_X1 U7260 ( .A1(n4335), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5816) );
  INV_X1 U7261 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6709) );
  NAND2_X1 U7262 ( .A1(n5811), .A2(n6709), .ZN(n5812) );
  AND2_X1 U7263 ( .A1(n5830), .A2(n5812), .ZN(n7444) );
  NAND2_X1 U7264 ( .A1(n5743), .A2(n7444), .ZN(n5815) );
  NAND2_X1 U7265 ( .A1(n6283), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5814) );
  NAND2_X1 U7266 ( .A1(n6293), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5813) );
  OR2_X1 U7267 ( .A1(n5804), .A2(n9504), .ZN(n5817) );
  XNOR2_X1 U7268 ( .A(n5817), .B(P1_IR_REG_6__SCAN_IN), .ZN(n6580) );
  INV_X1 U7269 ( .A(n6580), .ZN(n6710) );
  OR2_X1 U7270 ( .A1(n5838), .A2(n6657), .ZN(n5819) );
  OR2_X1 U7271 ( .A1(n6290), .A2(n10041), .ZN(n5818) );
  OAI211_X1 U7272 ( .C1(n5801), .C2(n6710), .A(n5819), .B(n5818), .ZN(n7440)
         );
  OAI22_X1 U7273 ( .A1(n7297), .A2(n6209), .B1(n7296), .B2(n5756), .ZN(n5820)
         );
  XNOR2_X1 U7274 ( .A(n5820), .B(n7304), .ZN(n5824) );
  OR2_X1 U7275 ( .A1(n7297), .A2(n6215), .ZN(n5822) );
  NAND2_X1 U7276 ( .A1(n7440), .A2(n6197), .ZN(n5821) );
  NAND2_X1 U7277 ( .A1(n5822), .A2(n5821), .ZN(n7436) );
  AOI22_X1 U7278 ( .A1(n5825), .A2(n7260), .B1(n5824), .B2(n7436), .ZN(n5823)
         );
  OAI21_X1 U7279 ( .B1(n5825), .B2(n7260), .A(n7436), .ZN(n5827) );
  INV_X1 U7280 ( .A(n5824), .ZN(n7437) );
  INV_X1 U7281 ( .A(n5825), .ZN(n7435) );
  NOR2_X1 U7282 ( .A1(n7436), .A2(n7260), .ZN(n5826) );
  AOI22_X1 U7283 ( .A1(n5827), .A2(n7437), .B1(n7435), .B2(n5826), .ZN(n5828)
         );
  NAND2_X1 U7284 ( .A1(n4335), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5835) );
  INV_X1 U7285 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5829) );
  NAND2_X1 U7286 ( .A1(n5830), .A2(n5829), .ZN(n5831) );
  AND2_X1 U7287 ( .A1(n5846), .A2(n5831), .ZN(n7477) );
  NAND2_X1 U7288 ( .A1(n5743), .A2(n7477), .ZN(n5834) );
  NAND2_X1 U7289 ( .A1(n6293), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5833) );
  NAND2_X1 U7290 ( .A1(n6283), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5832) );
  NAND2_X1 U7291 ( .A1(n5804), .A2(n5836), .ZN(n5852) );
  NAND2_X1 U7292 ( .A1(n5852), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5837) );
  XNOR2_X1 U7293 ( .A(n5837), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6732) );
  NAND2_X1 U7294 ( .A1(n6057), .A2(n6732), .ZN(n5840) );
  OR2_X1 U7295 ( .A1(n5838), .A2(n6668), .ZN(n5839) );
  OAI211_X1 U7296 ( .C1(n6290), .C2(n6667), .A(n5840), .B(n5839), .ZN(n7487)
         );
  OAI22_X1 U7297 ( .A1(n7300), .A2(n6209), .B1(n7469), .B2(n5756), .ZN(n5841)
         );
  XNOR2_X1 U7298 ( .A(n5841), .B(n7304), .ZN(n5844) );
  OAI22_X1 U7299 ( .A1(n7300), .A2(n6215), .B1(n7469), .B2(n6209), .ZN(n5843)
         );
  XNOR2_X1 U7300 ( .A(n5844), .B(n5843), .ZN(n7484) );
  INV_X1 U7301 ( .A(n7484), .ZN(n5842) );
  NAND2_X1 U7302 ( .A1(n5844), .A2(n5843), .ZN(n5845) );
  NAND2_X1 U7303 ( .A1(n4335), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5851) );
  NAND2_X1 U7304 ( .A1(n5846), .A2(n6759), .ZN(n5847) );
  AND2_X1 U7305 ( .A1(n5867), .A2(n5847), .ZN(n7539) );
  NAND2_X1 U7306 ( .A1(n5743), .A2(n7539), .ZN(n5850) );
  NAND2_X1 U7307 ( .A1(n6293), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5849) );
  NAND2_X1 U7308 ( .A1(n6283), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5848) );
  NAND2_X1 U7309 ( .A1(n5859), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5853) );
  XNOR2_X1 U7310 ( .A(n5853), .B(P1_IR_REG_8__SCAN_IN), .ZN(n6595) );
  AOI22_X1 U7311 ( .A1(n6302), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6057), .B2(
        n6595), .ZN(n5855) );
  NAND2_X1 U7312 ( .A1(n6673), .A2(n5751), .ZN(n5854) );
  NAND2_X1 U7313 ( .A1(n5855), .A2(n5854), .ZN(n7538) );
  OAI22_X1 U7314 ( .A1(n7480), .A2(n6215), .B1(n7411), .B2(n6209), .ZN(n5857)
         );
  OAI22_X1 U7315 ( .A1(n7480), .A2(n6209), .B1(n7411), .B2(n5756), .ZN(n5856)
         );
  XNOR2_X1 U7316 ( .A(n5856), .B(n6212), .ZN(n7536) );
  NAND2_X1 U7317 ( .A1(n6677), .A2(n5751), .ZN(n5865) );
  NOR2_X1 U7318 ( .A1(n5859), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n5862) );
  INV_X1 U7319 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9504) );
  OR2_X1 U7320 ( .A1(n5862), .A2(n9504), .ZN(n5860) );
  INV_X1 U7321 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n5861) );
  MUX2_X1 U7322 ( .A(n5860), .B(P1_IR_REG_31__SCAN_IN), .S(n5861), .Z(n5863)
         );
  NAND2_X1 U7323 ( .A1(n5862), .A2(n5861), .ZN(n5899) );
  NAND2_X1 U7324 ( .A1(n5863), .A2(n5899), .ZN(n6681) );
  INV_X1 U7325 ( .A(n6681), .ZN(n9624) );
  AOI22_X1 U7326 ( .A1(n6302), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n6057), .B2(
        n9624), .ZN(n5864) );
  NAND2_X1 U7327 ( .A1(n7520), .A2(n5755), .ZN(n5875) );
  INV_X1 U7328 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5866) );
  NAND2_X1 U7329 ( .A1(n5867), .A2(n5866), .ZN(n5868) );
  AND2_X1 U7330 ( .A1(n5885), .A2(n5868), .ZN(n7516) );
  NAND2_X1 U7331 ( .A1(n5743), .A2(n7516), .ZN(n5872) );
  NAND2_X1 U7332 ( .A1(n4335), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5871) );
  NAND2_X1 U7333 ( .A1(n6283), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5870) );
  NAND2_X1 U7334 ( .A1(n6293), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5869) );
  NAND4_X1 U7335 ( .A1(n5872), .A2(n5871), .A3(n5870), .A4(n5869), .ZN(n9125)
         );
  NAND2_X1 U7336 ( .A1(n9125), .A2(n6197), .ZN(n5874) );
  NAND2_X1 U7337 ( .A1(n5875), .A2(n5874), .ZN(n5876) );
  XNOR2_X1 U7338 ( .A(n5876), .B(n7304), .ZN(n5877) );
  AOI22_X1 U7339 ( .A1(n7520), .A2(n6197), .B1(n9125), .B2(n6179), .ZN(n5878)
         );
  XNOR2_X1 U7340 ( .A(n5877), .B(n5878), .ZN(n7515) );
  INV_X1 U7341 ( .A(n5877), .ZN(n5879) );
  NAND2_X1 U7342 ( .A1(n5879), .A2(n5878), .ZN(n5880) );
  NAND2_X1 U7343 ( .A1(n6682), .A2(n5751), .ZN(n5883) );
  NAND2_X1 U7344 ( .A1(n5899), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5881) );
  XNOR2_X1 U7345 ( .A(n5881), .B(P1_IR_REG_10__SCAN_IN), .ZN(n9630) );
  AOI22_X1 U7346 ( .A1(n6302), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6057), .B2(
        n9630), .ZN(n5882) );
  NAND2_X1 U7347 ( .A1(n7685), .A2(n5755), .ZN(n5892) );
  NAND2_X1 U7348 ( .A1(n4335), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5890) );
  NAND2_X1 U7349 ( .A1(n5885), .A2(n5884), .ZN(n5886) );
  AND2_X1 U7350 ( .A1(n5904), .A2(n5886), .ZN(n7688) );
  NAND2_X1 U7351 ( .A1(n5743), .A2(n7688), .ZN(n5889) );
  NAND2_X1 U7352 ( .A1(n6293), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5888) );
  NAND2_X1 U7353 ( .A1(n6283), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5887) );
  OR2_X1 U7354 ( .A1(n7620), .A2(n6209), .ZN(n5891) );
  NAND2_X1 U7355 ( .A1(n5892), .A2(n5891), .ZN(n5893) );
  XNOR2_X1 U7356 ( .A(n5893), .B(n6212), .ZN(n5898) );
  NAND2_X1 U7357 ( .A1(n7685), .A2(n6197), .ZN(n5895) );
  OR2_X1 U7358 ( .A1(n7620), .A2(n6215), .ZN(n5894) );
  NAND2_X1 U7359 ( .A1(n5895), .A2(n5894), .ZN(n5896) );
  XNOR2_X1 U7360 ( .A(n5898), .B(n5896), .ZN(n7683) );
  INV_X1 U7361 ( .A(n5896), .ZN(n5897) );
  NAND2_X1 U7362 ( .A1(n6686), .A2(n5751), .ZN(n5902) );
  OAI21_X1 U7363 ( .B1(n5899), .B2(P1_IR_REG_10__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5900) );
  XNOR2_X1 U7364 ( .A(n5900), .B(P1_IR_REG_11__SCAN_IN), .ZN(n9650) );
  AOI22_X1 U7365 ( .A1(n6302), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n6057), .B2(
        n9650), .ZN(n5901) );
  NAND2_X1 U7366 ( .A1(n5902), .A2(n5901), .ZN(n7629) );
  NAND2_X1 U7367 ( .A1(n7629), .A2(n5755), .ZN(n5911) );
  NAND2_X1 U7368 ( .A1(n4335), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5909) );
  INV_X1 U7369 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5903) );
  NAND2_X1 U7370 ( .A1(n5904), .A2(n5903), .ZN(n5905) );
  AND2_X1 U7371 ( .A1(n5929), .A2(n5905), .ZN(n7752) );
  NAND2_X1 U7372 ( .A1(n5743), .A2(n7752), .ZN(n5908) );
  NAND2_X1 U7373 ( .A1(n6293), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5907) );
  NAND2_X1 U7374 ( .A1(n6283), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5906) );
  NAND4_X1 U7375 ( .A1(n5909), .A2(n5908), .A3(n5907), .A4(n5906), .ZN(n9123)
         );
  NAND2_X1 U7376 ( .A1(n9123), .A2(n6197), .ZN(n5910) );
  NAND2_X1 U7377 ( .A1(n5911), .A2(n5910), .ZN(n5912) );
  XNOR2_X1 U7378 ( .A(n5912), .B(n6212), .ZN(n5916) );
  AND2_X1 U7379 ( .A1(n9123), .A2(n6179), .ZN(n5913) );
  AOI21_X1 U7380 ( .B1(n7629), .B2(n6197), .A(n5913), .ZN(n5917) );
  XNOR2_X1 U7381 ( .A(n5916), .B(n5917), .ZN(n7746) );
  INV_X1 U7382 ( .A(n7746), .ZN(n5914) );
  INV_X1 U7383 ( .A(n5916), .ZN(n5919) );
  INV_X1 U7384 ( .A(n5917), .ZN(n5918) );
  NAND2_X1 U7385 ( .A1(n5919), .A2(n5918), .ZN(n5920) );
  NAND2_X1 U7386 ( .A1(n6692), .A2(n5751), .ZN(n5927) );
  NOR2_X1 U7387 ( .A1(n5921), .A2(n9504), .ZN(n5922) );
  MUX2_X1 U7388 ( .A(n9504), .B(n5922), .S(P1_IR_REG_12__SCAN_IN), .Z(n5925)
         );
  INV_X1 U7389 ( .A(n5923), .ZN(n5924) );
  OR2_X1 U7390 ( .A1(n5925), .A2(n5924), .ZN(n6923) );
  INV_X1 U7391 ( .A(n6923), .ZN(n6604) );
  AOI22_X1 U7392 ( .A1(n6302), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6057), .B2(
        n6604), .ZN(n5926) );
  NAND2_X1 U7393 ( .A1(n9482), .A2(n5755), .ZN(n5936) );
  NAND2_X1 U7394 ( .A1(n4335), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5934) );
  NAND2_X1 U7395 ( .A1(n5929), .A2(n5928), .ZN(n5930) );
  AND2_X1 U7396 ( .A1(n5947), .A2(n5930), .ZN(n7854) );
  NAND2_X1 U7397 ( .A1(n5743), .A2(n7854), .ZN(n5933) );
  NAND2_X1 U7398 ( .A1(n6283), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5932) );
  NAND2_X1 U7399 ( .A1(n6293), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5931) );
  OR2_X1 U7400 ( .A1(n7787), .A2(n6209), .ZN(n5935) );
  NAND2_X1 U7401 ( .A1(n5936), .A2(n5935), .ZN(n5937) );
  XNOR2_X1 U7402 ( .A(n5937), .B(n7304), .ZN(n5939) );
  NOR2_X1 U7403 ( .A1(n7787), .A2(n6215), .ZN(n5938) );
  AOI21_X1 U7404 ( .B1(n9482), .B2(n6197), .A(n5938), .ZN(n5940) );
  XNOR2_X1 U7405 ( .A(n5939), .B(n5940), .ZN(n7849) );
  INV_X1 U7406 ( .A(n5939), .ZN(n5941) );
  NAND2_X1 U7407 ( .A1(n6718), .A2(n5751), .ZN(n5945) );
  NAND2_X1 U7408 ( .A1(n5923), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5942) );
  MUX2_X1 U7409 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5942), .S(
        P1_IR_REG_13__SCAN_IN), .Z(n5943) );
  OR2_X1 U7410 ( .A1(n5923), .A2(P1_IR_REG_13__SCAN_IN), .ZN(n5971) );
  AND2_X1 U7411 ( .A1(n5943), .A2(n5971), .ZN(n6855) );
  AOI22_X1 U7412 ( .A1(n6302), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n6057), .B2(
        n6855), .ZN(n5944) );
  NAND2_X1 U7413 ( .A1(n7868), .A2(n5755), .ZN(n5954) );
  NAND2_X1 U7414 ( .A1(n4335), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5952) );
  NAND2_X1 U7415 ( .A1(n5947), .A2(n5946), .ZN(n5948) );
  AND2_X1 U7416 ( .A1(n5960), .A2(n5948), .ZN(n7863) );
  NAND2_X1 U7417 ( .A1(n5743), .A2(n7863), .ZN(n5951) );
  NAND2_X1 U7418 ( .A1(n6283), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5950) );
  NAND2_X1 U7419 ( .A1(n6293), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5949) );
  NAND4_X1 U7420 ( .A1(n5952), .A2(n5951), .A3(n5950), .A4(n5949), .ZN(n9121)
         );
  NAND2_X1 U7421 ( .A1(n9121), .A2(n6197), .ZN(n5953) );
  NAND2_X1 U7422 ( .A1(n5954), .A2(n5953), .ZN(n5955) );
  XNOR2_X1 U7423 ( .A(n5955), .B(n6212), .ZN(n7859) );
  AND2_X1 U7424 ( .A1(n9121), .A2(n6179), .ZN(n5956) );
  AOI21_X1 U7425 ( .B1(n7868), .B2(n6197), .A(n5956), .ZN(n7858) );
  NAND2_X1 U7426 ( .A1(n6736), .A2(n5751), .ZN(n5959) );
  NAND2_X1 U7427 ( .A1(n5971), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5957) );
  XNOR2_X1 U7428 ( .A(n5957), .B(P1_IR_REG_14__SCAN_IN), .ZN(n9663) );
  AOI22_X1 U7429 ( .A1(n6302), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n6057), .B2(
        n9663), .ZN(n5958) );
  NAND2_X1 U7430 ( .A1(n9476), .A2(n5755), .ZN(n5967) );
  NAND2_X1 U7431 ( .A1(n4335), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5965) );
  INV_X1 U7432 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n7898) );
  NAND2_X1 U7433 ( .A1(n5960), .A2(n7898), .ZN(n5961) );
  AND2_X1 U7434 ( .A1(n5980), .A2(n5961), .ZN(n7899) );
  NAND2_X1 U7435 ( .A1(n5743), .A2(n7899), .ZN(n5964) );
  NAND2_X1 U7436 ( .A1(n6293), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5963) );
  NAND2_X1 U7437 ( .A1(n6283), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5962) );
  NAND4_X1 U7438 ( .A1(n5965), .A2(n5964), .A3(n5963), .A4(n5962), .ZN(n9120)
         );
  NAND2_X1 U7439 ( .A1(n9120), .A2(n6197), .ZN(n5966) );
  NAND2_X1 U7440 ( .A1(n5967), .A2(n5966), .ZN(n5968) );
  XNOR2_X1 U7441 ( .A(n5968), .B(n7304), .ZN(n7895) );
  NAND2_X1 U7442 ( .A1(n9476), .A2(n6197), .ZN(n5970) );
  NAND2_X1 U7443 ( .A1(n9120), .A2(n6179), .ZN(n5969) );
  NAND2_X1 U7444 ( .A1(n5970), .A2(n5969), .ZN(n5989) );
  NAND2_X1 U7445 ( .A1(n6828), .A2(n5751), .ZN(n5978) );
  NOR2_X1 U7446 ( .A1(n5971), .A2(P1_IR_REG_14__SCAN_IN), .ZN(n5974) );
  OR2_X1 U7447 ( .A1(n5974), .A2(n9504), .ZN(n5972) );
  MUX2_X1 U7448 ( .A(n5972), .B(P1_IR_REG_31__SCAN_IN), .S(n5973), .Z(n5975)
         );
  NAND2_X1 U7449 ( .A1(n5974), .A2(n5973), .ZN(n6000) );
  NAND2_X1 U7450 ( .A1(n5975), .A2(n6000), .ZN(n7422) );
  INV_X1 U7451 ( .A(n7422), .ZN(n5976) );
  AOI22_X1 U7452 ( .A1(n6302), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n6057), .B2(
        n5976), .ZN(n5977) );
  NAND2_X1 U7453 ( .A1(n9113), .A2(n5755), .ZN(n5987) );
  NAND2_X1 U7454 ( .A1(n4335), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5985) );
  INV_X1 U7455 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n5979) );
  NAND2_X1 U7456 ( .A1(n5980), .A2(n5979), .ZN(n5981) );
  AND2_X1 U7457 ( .A1(n6007), .A2(n5981), .ZN(n9105) );
  NAND2_X1 U7458 ( .A1(n5743), .A2(n9105), .ZN(n5984) );
  NAND2_X1 U7459 ( .A1(n6293), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5983) );
  NAND2_X1 U7460 ( .A1(n6283), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5982) );
  NAND4_X1 U7461 ( .A1(n5985), .A2(n5984), .A3(n5983), .A4(n5982), .ZN(n9119)
         );
  NAND2_X1 U7462 ( .A1(n9119), .A2(n6197), .ZN(n5986) );
  NAND2_X1 U7463 ( .A1(n5987), .A2(n5986), .ZN(n5988) );
  XNOR2_X1 U7464 ( .A(n5988), .B(n7304), .ZN(n5994) );
  INV_X1 U7465 ( .A(n7895), .ZN(n5990) );
  INV_X1 U7466 ( .A(n5989), .ZN(n7894) );
  NAND2_X1 U7467 ( .A1(n5990), .A2(n7894), .ZN(n5993) );
  AND2_X1 U7468 ( .A1(n5994), .A2(n5993), .ZN(n5991) );
  NAND2_X1 U7469 ( .A1(n7897), .A2(n5993), .ZN(n5997) );
  INV_X1 U7470 ( .A(n5994), .ZN(n5995) );
  AND2_X1 U7471 ( .A1(n5995), .A2(n4367), .ZN(n5996) );
  NAND2_X1 U7472 ( .A1(n5997), .A2(n5996), .ZN(n9098) );
  NAND2_X1 U7473 ( .A1(n9113), .A2(n6197), .ZN(n5999) );
  NAND2_X1 U7474 ( .A1(n9119), .A2(n6179), .ZN(n5998) );
  NAND2_X1 U7475 ( .A1(n5999), .A2(n5998), .ZN(n9101) );
  NAND2_X1 U7476 ( .A1(n9098), .A2(n9101), .ZN(n9021) );
  NAND2_X1 U7477 ( .A1(n6967), .A2(n5751), .ZN(n6005) );
  NAND2_X1 U7478 ( .A1(n6000), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6001) );
  MUX2_X1 U7479 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6001), .S(
        P1_IR_REG_16__SCAN_IN), .Z(n6002) );
  AND2_X1 U7480 ( .A1(n6003), .A2(n6002), .ZN(n7588) );
  AOI22_X1 U7481 ( .A1(n6302), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n6057), .B2(
        n7588), .ZN(n6004) );
  NAND2_X1 U7482 ( .A1(n7939), .A2(n5755), .ZN(n6014) );
  NAND2_X1 U7483 ( .A1(n4335), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n6012) );
  NAND2_X1 U7484 ( .A1(n6007), .A2(n6006), .ZN(n6008) );
  AND2_X1 U7485 ( .A1(n6025), .A2(n6008), .ZN(n9029) );
  NAND2_X1 U7486 ( .A1(n5743), .A2(n9029), .ZN(n6011) );
  NAND2_X1 U7487 ( .A1(n6293), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n6010) );
  NAND2_X1 U7488 ( .A1(n5745), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n6009) );
  OR2_X1 U7489 ( .A1(n9110), .A2(n6209), .ZN(n6013) );
  NAND2_X1 U7490 ( .A1(n6014), .A2(n6013), .ZN(n6015) );
  XNOR2_X1 U7491 ( .A(n6015), .B(n6212), .ZN(n6018) );
  NOR2_X1 U7492 ( .A1(n9110), .A2(n6215), .ZN(n6016) );
  AOI21_X1 U7493 ( .B1(n7939), .B2(n6197), .A(n6016), .ZN(n6017) );
  NAND2_X1 U7494 ( .A1(n6018), .A2(n6017), .ZN(n6020) );
  OR2_X1 U7495 ( .A1(n6018), .A2(n6017), .ZN(n6019) );
  AND2_X1 U7496 ( .A1(n6020), .A2(n6019), .ZN(n9020) );
  NAND2_X1 U7497 ( .A1(n6956), .A2(n5751), .ZN(n6023) );
  XNOR2_X1 U7498 ( .A(n6021), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9161) );
  AOI22_X1 U7499 ( .A1(n6302), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n6057), .B2(
        n9161), .ZN(n6022) );
  NAND2_X1 U7500 ( .A1(n9470), .A2(n5755), .ZN(n6032) );
  NAND2_X1 U7501 ( .A1(n4335), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n6030) );
  INV_X1 U7502 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n6024) );
  NAND2_X1 U7503 ( .A1(n6025), .A2(n6024), .ZN(n6026) );
  AND2_X1 U7504 ( .A1(n6043), .A2(n6026), .ZN(n9394) );
  NAND2_X1 U7505 ( .A1(n5743), .A2(n9394), .ZN(n6029) );
  NAND2_X1 U7506 ( .A1(n6293), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n6028) );
  NAND2_X1 U7507 ( .A1(n6283), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n6027) );
  NAND4_X1 U7508 ( .A1(n6030), .A2(n6029), .A3(n6028), .A4(n6027), .ZN(n9384)
         );
  NAND2_X1 U7509 ( .A1(n9384), .A2(n6197), .ZN(n6031) );
  NAND2_X1 U7510 ( .A1(n6032), .A2(n6031), .ZN(n6033) );
  XNOR2_X1 U7511 ( .A(n6033), .B(n7304), .ZN(n6035) );
  AND2_X1 U7512 ( .A1(n9384), .A2(n6179), .ZN(n6034) );
  AOI21_X1 U7513 ( .B1(n9470), .B2(n6197), .A(n6034), .ZN(n6036) );
  XNOR2_X1 U7514 ( .A(n6035), .B(n6036), .ZN(n9034) );
  INV_X1 U7515 ( .A(n6035), .ZN(n6037) );
  NAND2_X1 U7516 ( .A1(n6037), .A2(n6036), .ZN(n6038) );
  NAND2_X1 U7517 ( .A1(n7088), .A2(n5751), .ZN(n6041) );
  XNOR2_X1 U7518 ( .A(n6039), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9175) );
  AOI22_X1 U7519 ( .A1(n6302), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n6057), .B2(
        n9175), .ZN(n6040) );
  NAND2_X1 U7520 ( .A1(n9465), .A2(n5755), .ZN(n6050) );
  NAND2_X1 U7521 ( .A1(n4335), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n6048) );
  NAND2_X1 U7522 ( .A1(n6043), .A2(n6042), .ZN(n6044) );
  AND2_X1 U7523 ( .A1(n6061), .A2(n6044), .ZN(n9376) );
  NAND2_X1 U7524 ( .A1(n5743), .A2(n9376), .ZN(n6047) );
  NAND2_X1 U7525 ( .A1(n6293), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n6046) );
  NAND2_X1 U7526 ( .A1(n6283), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n6045) );
  OR2_X1 U7527 ( .A1(n9037), .A2(n6209), .ZN(n6049) );
  NAND2_X1 U7528 ( .A1(n6050), .A2(n6049), .ZN(n6051) );
  XNOR2_X1 U7529 ( .A(n6051), .B(n6212), .ZN(n6055) );
  NAND2_X1 U7530 ( .A1(n9465), .A2(n6197), .ZN(n6053) );
  OR2_X1 U7531 ( .A1(n9037), .A2(n6215), .ZN(n6052) );
  NAND2_X1 U7532 ( .A1(n6053), .A2(n6052), .ZN(n9075) );
  INV_X1 U7533 ( .A(n6055), .ZN(n6056) );
  NAND2_X1 U7534 ( .A1(n7128), .A2(n5751), .ZN(n6059) );
  AOI22_X1 U7535 ( .A1(n6302), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9282), .B2(
        n6057), .ZN(n6058) );
  NAND2_X1 U7536 ( .A1(n9460), .A2(n5755), .ZN(n6068) );
  INV_X1 U7537 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n6060) );
  NAND2_X1 U7538 ( .A1(n6061), .A2(n6060), .ZN(n6062) );
  AND2_X1 U7539 ( .A1(n6078), .A2(n6062), .ZN(n9361) );
  NAND2_X1 U7540 ( .A1(n9361), .A2(n4319), .ZN(n6066) );
  NAND2_X1 U7541 ( .A1(n4317), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n6065) );
  NAND2_X1 U7542 ( .A1(n4335), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n6064) );
  NAND2_X1 U7543 ( .A1(n5745), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n6063) );
  NAND4_X1 U7544 ( .A1(n6066), .A2(n6065), .A3(n6064), .A4(n6063), .ZN(n9383)
         );
  NAND2_X1 U7545 ( .A1(n9383), .A2(n6197), .ZN(n6067) );
  NAND2_X1 U7546 ( .A1(n6068), .A2(n6067), .ZN(n6069) );
  XNOR2_X1 U7547 ( .A(n6069), .B(n6212), .ZN(n6071) );
  AND2_X1 U7548 ( .A1(n9383), .A2(n6179), .ZN(n6070) );
  AOI21_X1 U7549 ( .B1(n9460), .B2(n6197), .A(n6070), .ZN(n6072) );
  NAND2_X1 U7550 ( .A1(n6071), .A2(n6072), .ZN(n8995) );
  INV_X1 U7551 ( .A(n6071), .ZN(n6074) );
  INV_X1 U7552 ( .A(n6072), .ZN(n6073) );
  NAND2_X1 U7553 ( .A1(n6074), .A2(n6073), .ZN(n8996) );
  NAND2_X1 U7554 ( .A1(n6075), .A2(n8996), .ZN(n9050) );
  NAND2_X1 U7555 ( .A1(n7287), .A2(n5751), .ZN(n6077) );
  NAND2_X1 U7556 ( .A1(n6302), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n6076) );
  NAND2_X1 U7557 ( .A1(n9455), .A2(n5755), .ZN(n6083) );
  NAND2_X1 U7558 ( .A1(n6078), .A2(n9054), .ZN(n6079) );
  NAND2_X1 U7559 ( .A1(n6093), .A2(n6079), .ZN(n9346) );
  AOI22_X1 U7560 ( .A1(n4335), .A2(P1_REG1_REG_20__SCAN_IN), .B1(n6293), .B2(
        P1_REG0_REG_20__SCAN_IN), .ZN(n6081) );
  NAND2_X1 U7561 ( .A1(n6283), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n6080) );
  OAI211_X1 U7562 ( .C1(n9346), .C2(n6095), .A(n6081), .B(n6080), .ZN(n9369)
         );
  NAND2_X1 U7563 ( .A1(n9369), .A2(n6197), .ZN(n6082) );
  NAND2_X1 U7564 ( .A1(n6083), .A2(n6082), .ZN(n6084) );
  XNOR2_X1 U7565 ( .A(n6084), .B(n6212), .ZN(n9052) );
  AND2_X1 U7566 ( .A1(n9369), .A2(n6179), .ZN(n6085) );
  AOI21_X1 U7567 ( .B1(n9455), .B2(n6197), .A(n6085), .ZN(n6087) );
  NAND2_X1 U7568 ( .A1(n9052), .A2(n6087), .ZN(n6086) );
  INV_X1 U7569 ( .A(n9052), .ZN(n6088) );
  INV_X1 U7570 ( .A(n6087), .ZN(n9051) );
  NAND2_X1 U7571 ( .A1(n6088), .A2(n9051), .ZN(n6089) );
  NAND2_X1 U7572 ( .A1(n7340), .A2(n5751), .ZN(n6091) );
  NAND2_X1 U7573 ( .A1(n6302), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n6090) );
  NAND2_X1 U7574 ( .A1(n9452), .A2(n5755), .ZN(n6100) );
  INV_X1 U7575 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n6092) );
  NAND2_X1 U7576 ( .A1(n6093), .A2(n6092), .ZN(n6094) );
  NAND2_X1 U7577 ( .A1(n6111), .A2(n6094), .ZN(n9336) );
  OR2_X1 U7578 ( .A1(n9336), .A2(n6095), .ZN(n6098) );
  AOI22_X1 U7579 ( .A1(n4335), .A2(P1_REG1_REG_21__SCAN_IN), .B1(n6293), .B2(
        P1_REG0_REG_21__SCAN_IN), .ZN(n6097) );
  NAND2_X1 U7580 ( .A1(n5745), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n6096) );
  OR2_X1 U7581 ( .A1(n9055), .A2(n6209), .ZN(n6099) );
  NAND2_X1 U7582 ( .A1(n6100), .A2(n6099), .ZN(n6101) );
  XNOR2_X1 U7583 ( .A(n6101), .B(n7304), .ZN(n6104) );
  NAND2_X1 U7584 ( .A1(n9452), .A2(n6197), .ZN(n6103) );
  OR2_X1 U7585 ( .A1(n9055), .A2(n6215), .ZN(n6102) );
  NAND2_X1 U7586 ( .A1(n6103), .A2(n6102), .ZN(n6105) );
  INV_X1 U7587 ( .A(n6104), .ZN(n6107) );
  INV_X1 U7588 ( .A(n6105), .ZN(n6106) );
  NAND2_X1 U7589 ( .A1(n7676), .A2(n5751), .ZN(n6109) );
  NAND2_X1 U7590 ( .A1(n6302), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n6108) );
  INV_X1 U7591 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n6110) );
  NAND2_X1 U7592 ( .A1(n6111), .A2(n6110), .ZN(n6112) );
  NAND2_X1 U7593 ( .A1(n6113), .A2(n6112), .ZN(n9314) );
  OR2_X1 U7594 ( .A1(n9314), .A2(n6095), .ZN(n6119) );
  INV_X1 U7595 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n6116) );
  NAND2_X1 U7596 ( .A1(n6293), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n6115) );
  NAND2_X1 U7597 ( .A1(n5745), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n6114) );
  OAI211_X1 U7598 ( .C1(n6296), .C2(n6116), .A(n6115), .B(n6114), .ZN(n6117)
         );
  INV_X1 U7599 ( .A(n6117), .ZN(n6118) );
  NAND2_X1 U7600 ( .A1(n6119), .A2(n6118), .ZN(n9118) );
  AND2_X1 U7601 ( .A1(n9118), .A2(n6179), .ZN(n6120) );
  AOI21_X1 U7602 ( .B1(n9317), .B2(n6197), .A(n6120), .ZN(n6125) );
  NAND2_X1 U7603 ( .A1(n9317), .A2(n5755), .ZN(n6122) );
  NAND2_X1 U7604 ( .A1(n9118), .A2(n6197), .ZN(n6121) );
  NAND2_X1 U7605 ( .A1(n6122), .A2(n6121), .ZN(n6123) );
  XNOR2_X1 U7606 ( .A(n6123), .B(n7304), .ZN(n9065) );
  INV_X1 U7607 ( .A(n6124), .ZN(n6126) );
  NAND2_X1 U7608 ( .A1(n9441), .A2(n5755), .ZN(n6128) );
  NAND2_X1 U7609 ( .A1(n9308), .A2(n6197), .ZN(n6127) );
  NAND2_X1 U7610 ( .A1(n6128), .A2(n6127), .ZN(n6129) );
  XNOR2_X1 U7611 ( .A(n6129), .B(n7304), .ZN(n6130) );
  NAND2_X1 U7612 ( .A1(n7769), .A2(n5751), .ZN(n6132) );
  NAND2_X1 U7613 ( .A1(n6302), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n6131) );
  INV_X1 U7614 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9044) );
  NAND2_X1 U7615 ( .A1(n6133), .A2(n9044), .ZN(n6134) );
  AND2_X1 U7616 ( .A1(n6150), .A2(n6134), .ZN(n9280) );
  NAND2_X1 U7617 ( .A1(n9280), .A2(n5743), .ZN(n6140) );
  INV_X1 U7618 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n6137) );
  NAND2_X1 U7619 ( .A1(n5745), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n6136) );
  NAND2_X1 U7620 ( .A1(n4317), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n6135) );
  OAI211_X1 U7621 ( .C1(n6296), .C2(n6137), .A(n6136), .B(n6135), .ZN(n6138)
         );
  INV_X1 U7622 ( .A(n6138), .ZN(n6139) );
  AOI22_X1 U7623 ( .A1(n9436), .A2(n6197), .B1(n6179), .B2(n9265), .ZN(n6144)
         );
  NAND2_X1 U7624 ( .A1(n9436), .A2(n5755), .ZN(n6142) );
  NAND2_X1 U7625 ( .A1(n9265), .A2(n6197), .ZN(n6141) );
  NAND2_X1 U7626 ( .A1(n6142), .A2(n6141), .ZN(n6143) );
  XNOR2_X1 U7627 ( .A(n6143), .B(n7304), .ZN(n6145) );
  XOR2_X1 U7628 ( .A(n6144), .B(n6145), .Z(n9042) );
  NAND2_X1 U7629 ( .A1(n7823), .A2(n5751), .ZN(n6147) );
  NAND2_X1 U7630 ( .A1(n6302), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n6146) );
  NAND2_X1 U7631 ( .A1(n9429), .A2(n5755), .ZN(n6159) );
  INV_X1 U7632 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n6149) );
  NAND2_X1 U7633 ( .A1(n6150), .A2(n6149), .ZN(n6151) );
  NAND2_X1 U7634 ( .A1(n6168), .A2(n6151), .ZN(n9256) );
  INV_X1 U7635 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n6154) );
  NAND2_X1 U7636 ( .A1(n4317), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n6153) );
  NAND2_X1 U7637 ( .A1(n5745), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n6152) );
  OAI211_X1 U7638 ( .C1(n6296), .C2(n6154), .A(n6153), .B(n6152), .ZN(n6155)
         );
  INV_X1 U7639 ( .A(n6155), .ZN(n6156) );
  NAND2_X1 U7640 ( .A1(n9248), .A2(n6197), .ZN(n6158) );
  NAND2_X1 U7641 ( .A1(n6159), .A2(n6158), .ZN(n6160) );
  XNOR2_X1 U7642 ( .A(n6160), .B(n7304), .ZN(n6161) );
  AOI22_X1 U7643 ( .A1(n9429), .A2(n6197), .B1(n6179), .B2(n9248), .ZN(n6162)
         );
  XNOR2_X1 U7644 ( .A(n6161), .B(n6162), .ZN(n9013) );
  INV_X1 U7645 ( .A(n6161), .ZN(n6163) );
  NAND2_X1 U7646 ( .A1(n6302), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n6164) );
  NAND2_X1 U7647 ( .A1(n9424), .A2(n5755), .ZN(n6177) );
  INV_X1 U7648 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n6167) );
  NAND2_X1 U7649 ( .A1(n6168), .A2(n6167), .ZN(n6169) );
  NAND2_X1 U7650 ( .A1(n6204), .A2(n6169), .ZN(n9090) );
  INV_X1 U7651 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n6172) );
  NAND2_X1 U7652 ( .A1(n6293), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n6171) );
  NAND2_X1 U7653 ( .A1(n5745), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n6170) );
  OAI211_X1 U7654 ( .C1(n6296), .C2(n6172), .A(n6171), .B(n6170), .ZN(n6173)
         );
  INV_X1 U7655 ( .A(n6173), .ZN(n6174) );
  NAND2_X1 U7656 ( .A1(n9264), .A2(n6197), .ZN(n6176) );
  NAND2_X1 U7657 ( .A1(n6177), .A2(n6176), .ZN(n6178) );
  XNOR2_X1 U7658 ( .A(n6178), .B(n7304), .ZN(n6181) );
  AND2_X1 U7659 ( .A1(n9264), .A2(n6179), .ZN(n6180) );
  AOI21_X1 U7660 ( .B1(n9424), .B2(n6197), .A(n6180), .ZN(n6182) );
  XNOR2_X1 U7661 ( .A(n6181), .B(n6182), .ZN(n9089) );
  INV_X1 U7662 ( .A(n6182), .ZN(n6183) );
  NAND2_X1 U7663 ( .A1(n9088), .A2(n6184), .ZN(n8977) );
  NAND2_X1 U7664 ( .A1(n7891), .A2(n5751), .ZN(n6186) );
  NAND2_X1 U7665 ( .A1(n6302), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n6185) );
  NAND2_X1 U7666 ( .A1(n9420), .A2(n5755), .ZN(n6194) );
  XNOR2_X1 U7667 ( .A(n6204), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n9226) );
  NAND2_X1 U7668 ( .A1(n9226), .A2(n5743), .ZN(n6192) );
  INV_X1 U7669 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n6189) );
  NAND2_X1 U7670 ( .A1(n6293), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6188) );
  NAND2_X1 U7671 ( .A1(n6283), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n6187) );
  OAI211_X1 U7672 ( .C1(n6296), .C2(n6189), .A(n6188), .B(n6187), .ZN(n6190)
         );
  INV_X1 U7673 ( .A(n6190), .ZN(n6191) );
  OR2_X1 U7674 ( .A1(n9210), .A2(n6209), .ZN(n6193) );
  NAND2_X1 U7675 ( .A1(n6194), .A2(n6193), .ZN(n6195) );
  XNOR2_X1 U7676 ( .A(n6195), .B(n7304), .ZN(n8975) );
  INV_X1 U7677 ( .A(n8975), .ZN(n6198) );
  NOR2_X1 U7678 ( .A1(n9210), .A2(n6215), .ZN(n6196) );
  AOI21_X1 U7679 ( .B1(n9420), .B2(n6197), .A(n6196), .ZN(n8974) );
  INV_X1 U7680 ( .A(n8974), .ZN(n6239) );
  NAND2_X1 U7681 ( .A1(n6198), .A2(n8974), .ZN(n6199) );
  NAND2_X1 U7682 ( .A1(n8977), .A2(n6199), .ZN(n6240) );
  INV_X1 U7683 ( .A(n6240), .ZN(n6238) );
  NAND2_X1 U7684 ( .A1(n7926), .A2(n5751), .ZN(n6201) );
  NAND2_X1 U7685 ( .A1(n6302), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n6200) );
  NAND2_X1 U7686 ( .A1(n9214), .A2(n5755), .ZN(n6211) );
  INV_X1 U7687 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n8978) );
  INV_X1 U7688 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n6202) );
  OAI21_X1 U7689 ( .B1(n6204), .B2(n8978), .A(n6202), .ZN(n6205) );
  NAND2_X1 U7690 ( .A1(P1_REG3_REG_28__SCAN_IN), .A2(P1_REG3_REG_27__SCAN_IN), 
        .ZN(n6203) );
  INV_X1 U7691 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n9417) );
  NAND2_X1 U7692 ( .A1(n6293), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6207) );
  NAND2_X1 U7693 ( .A1(n5745), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n6206) );
  OAI211_X1 U7694 ( .C1(n6296), .C2(n9417), .A(n6207), .B(n6206), .ZN(n6208)
         );
  OR2_X1 U7695 ( .A1(n9231), .A2(n6209), .ZN(n6210) );
  NAND2_X1 U7696 ( .A1(n6211), .A2(n6210), .ZN(n6213) );
  XNOR2_X1 U7697 ( .A(n6213), .B(n6212), .ZN(n6217) );
  NAND2_X1 U7698 ( .A1(n9214), .A2(n6197), .ZN(n6214) );
  OAI21_X1 U7699 ( .B1(n9231), .B2(n6215), .A(n6214), .ZN(n6216) );
  XNOR2_X1 U7700 ( .A(n6217), .B(n6216), .ZN(n6260) );
  INV_X1 U7701 ( .A(n6260), .ZN(n6237) );
  AND3_X1 U7702 ( .A1(n7828), .A2(P1_B_REG_SCAN_IN), .A3(n7802), .ZN(n6220) );
  INV_X1 U7703 ( .A(n7802), .ZN(n6218) );
  INV_X1 U7704 ( .A(P1_B_REG_SCAN_IN), .ZN(n7982) );
  AND2_X1 U7705 ( .A1(n6218), .A2(n7982), .ZN(n6219) );
  NAND2_X1 U7706 ( .A1(n7933), .A2(n7802), .ZN(n6221) );
  OAI21_X1 U7707 ( .B1(n6772), .B2(P1_D_REG_0__SCAN_IN), .A(n6221), .ZN(n6766)
         );
  NOR4_X1 U7708 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_17__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n6225) );
  NOR4_X1 U7709 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n6224) );
  NOR4_X1 U7710 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n6223) );
  NOR4_X1 U7711 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n6222) );
  AND4_X1 U7712 ( .A1(n6225), .A2(n6224), .A3(n6223), .A4(n6222), .ZN(n6231)
         );
  NOR2_X1 U7713 ( .A1(P1_D_REG_9__SCAN_IN), .A2(P1_D_REG_15__SCAN_IN), .ZN(
        n6229) );
  NOR4_X1 U7714 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_11__SCAN_IN), .A4(P1_D_REG_18__SCAN_IN), .ZN(n6228) );
  NOR4_X1 U7715 ( .A1(P1_D_REG_5__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_7__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n6227) );
  NOR4_X1 U7716 ( .A1(P1_D_REG_28__SCAN_IN), .A2(P1_D_REG_2__SCAN_IN), .A3(
        P1_D_REG_3__SCAN_IN), .A4(P1_D_REG_4__SCAN_IN), .ZN(n6226) );
  AND4_X1 U7717 ( .A1(n6229), .A2(n6228), .A3(n6227), .A4(n6226), .ZN(n6230)
         );
  NAND2_X1 U7718 ( .A1(n6231), .A2(n6230), .ZN(n6769) );
  INV_X1 U7719 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n6691) );
  NOR2_X1 U7720 ( .A1(n6769), .A2(n6691), .ZN(n6232) );
  NAND2_X1 U7721 ( .A1(n7933), .A2(n7828), .ZN(n6771) );
  OAI21_X1 U7722 ( .B1(n6772), .B2(n6232), .A(n6771), .ZN(n6636) );
  OR2_X1 U7723 ( .A1(n6766), .A2(n6636), .ZN(n6255) );
  NAND2_X1 U7724 ( .A1(n4385), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6234) );
  XNOR2_X1 U7725 ( .A(n6234), .B(n6233), .ZN(n6545) );
  AND2_X1 U7726 ( .A1(n6545), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6235) );
  NOR2_X1 U7727 ( .A1(n6255), .A2(n6767), .ZN(n6252) );
  NOR2_X1 U7728 ( .A1(n9483), .A2(n6631), .ZN(n6236) );
  NAND2_X1 U7729 ( .A1(n6238), .A2(n4888), .ZN(n6265) );
  NAND2_X1 U7730 ( .A1(n8975), .A2(n6239), .ZN(n6259) );
  NAND4_X1 U7731 ( .A1(n6240), .A2(n6260), .A3(n6259), .A4(n9087), .ZN(n6264)
         );
  INV_X1 U7732 ( .A(n7936), .ZN(n6615) );
  AND2_X1 U7733 ( .A1(n6932), .A2(n6615), .ZN(n9681) );
  NAND2_X1 U7734 ( .A1(n6252), .A2(n9681), .ZN(n6242) );
  INV_X1 U7735 ( .A(n6243), .ZN(n7991) );
  INV_X1 U7736 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n9958) );
  NAND2_X1 U7737 ( .A1(n4335), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n6245) );
  NAND2_X1 U7738 ( .A1(n5745), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6244) );
  OAI211_X1 U7739 ( .C1(n6246), .C2(n9958), .A(n6245), .B(n6244), .ZN(n6247)
         );
  AOI21_X1 U7740 ( .B1(n7991), .B2(n5743), .A(n6247), .ZN(n9209) );
  INV_X1 U7741 ( .A(n6631), .ZN(n6248) );
  OR2_X1 U7742 ( .A1(n6248), .A2(n6527), .ZN(n7305) );
  INV_X1 U7743 ( .A(n6249), .ZN(n6803) );
  NOR2_X1 U7744 ( .A1(n7305), .A2(n6803), .ZN(n6250) );
  NAND2_X1 U7745 ( .A1(n6252), .A2(n6250), .ZN(n9109) );
  NOR2_X1 U7746 ( .A1(n7305), .A2(n6249), .ZN(n6251) );
  NAND2_X1 U7747 ( .A1(n6252), .A2(n6251), .ZN(n9092) );
  NAND2_X1 U7748 ( .A1(n9249), .A2(n9104), .ZN(n6258) );
  NAND2_X1 U7749 ( .A1(n6255), .A2(n9714), .ZN(n6842) );
  NAND4_X1 U7750 ( .A1(n6842), .A2(n6543), .A3(n6545), .A4(n6841), .ZN(n6253)
         );
  NAND2_X1 U7751 ( .A1(n6253), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6256) );
  AND2_X1 U7752 ( .A1(n9681), .A2(n9697), .ZN(n6254) );
  NAND2_X1 U7753 ( .A1(n6255), .A2(n6254), .ZN(n6843) );
  NAND2_X1 U7754 ( .A1(n6256), .A2(n6843), .ZN(n9106) );
  AOI22_X1 U7755 ( .A1(n9216), .A2(n9106), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n6257) );
  OAI211_X1 U7756 ( .C1(n9209), .C2(n9109), .A(n6258), .B(n6257), .ZN(n6262)
         );
  NOR3_X1 U7757 ( .A1(n6260), .A2(n9115), .A3(n6259), .ZN(n6261) );
  AOI211_X1 U7758 ( .C1(n9214), .C2(n9112), .A(n6262), .B(n6261), .ZN(n6263)
         );
  NAND3_X1 U7759 ( .A1(n6265), .A2(n6264), .A3(n6263), .ZN(P1_U3218) );
  INV_X1 U7760 ( .A(SI_28_), .ZN(n6268) );
  INV_X1 U7761 ( .A(SI_29_), .ZN(n6298) );
  MUX2_X1 U7762 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .S(n4994), .Z(n6299) );
  NAND2_X1 U7763 ( .A1(n6270), .A2(n6299), .ZN(n6271) );
  NAND2_X1 U7764 ( .A1(n6271), .A2(n4890), .ZN(n6289) );
  INV_X1 U7765 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n6272) );
  INV_X1 U7766 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n7938) );
  INV_X1 U7767 ( .A(SI_30_), .ZN(n6273) );
  NAND2_X1 U7768 ( .A1(n6274), .A2(n6273), .ZN(n6277) );
  INV_X1 U7769 ( .A(n6274), .ZN(n6275) );
  NAND2_X1 U7770 ( .A1(n6275), .A2(SI_30_), .ZN(n6276) );
  NAND2_X1 U7771 ( .A1(n6277), .A2(n6276), .ZN(n6288) );
  INV_X1 U7772 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n8170) );
  XNOR2_X1 U7773 ( .A(n6278), .B(SI_31_), .ZN(n6279) );
  NAND2_X1 U7774 ( .A1(n8169), .A2(n5751), .ZN(n6282) );
  OR2_X1 U7775 ( .A1(n6290), .A2(n6705), .ZN(n6281) );
  NAND2_X1 U7776 ( .A1(n4335), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6287) );
  NAND2_X1 U7777 ( .A1(n6283), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6286) );
  NAND2_X1 U7778 ( .A1(n6293), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6285) );
  AND3_X1 U7779 ( .A1(n6287), .A2(n6286), .A3(n6285), .ZN(n6367) );
  NAND2_X1 U7780 ( .A1(n9193), .A2(n6367), .ZN(n6467) );
  NAND2_X1 U7781 ( .A1(n8172), .A2(n5751), .ZN(n6292) );
  OR2_X1 U7782 ( .A1(n6290), .A2(n7938), .ZN(n6291) );
  NAND2_X1 U7783 ( .A1(n5745), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n6295) );
  NAND2_X1 U7784 ( .A1(n4317), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n6294) );
  OAI211_X1 U7785 ( .C1(n6296), .C2(n9560), .A(n6295), .B(n6294), .ZN(n9117)
         );
  INV_X1 U7786 ( .A(n9117), .ZN(n6323) );
  OR2_X1 U7787 ( .A1(n9198), .A2(n6323), .ZN(n6297) );
  NAND2_X1 U7788 ( .A1(n9214), .A2(n9231), .ZN(n7978) );
  XNOR2_X1 U7789 ( .A(n6299), .B(n6298), .ZN(n6300) );
  NAND2_X1 U7790 ( .A1(n8013), .A2(n5751), .ZN(n6304) );
  NAND2_X1 U7791 ( .A1(n6302), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n6303) );
  NOR2_X1 U7792 ( .A1(n7986), .A2(n9209), .ZN(n6330) );
  NAND2_X1 U7793 ( .A1(n9420), .A2(n9210), .ZN(n6372) );
  INV_X1 U7794 ( .A(n9265), .ZN(n9291) );
  OR2_X1 U7795 ( .A1(n9436), .A2(n9291), .ZN(n6446) );
  NAND2_X1 U7796 ( .A1(n9436), .A2(n9291), .ZN(n9260) );
  AND2_X1 U7797 ( .A1(n6446), .A2(n9260), .ZN(n9274) );
  INV_X1 U7798 ( .A(n9274), .ZN(n9271) );
  NAND2_X1 U7799 ( .A1(n9429), .A2(n9278), .ZN(n6441) );
  INV_X1 U7800 ( .A(n9308), .ZN(n9277) );
  OR2_X1 U7801 ( .A1(n9441), .A2(n9277), .ZN(n9272) );
  NAND2_X1 U7802 ( .A1(n9441), .A2(n9277), .ZN(n7971) );
  AND2_X1 U7803 ( .A1(n9272), .A2(n7971), .ZN(n9288) );
  INV_X1 U7804 ( .A(n9118), .ZN(n9332) );
  OR2_X1 U7805 ( .A1(n9317), .A2(n9332), .ZN(n6447) );
  NAND2_X1 U7806 ( .A1(n9317), .A2(n9332), .ZN(n6449) );
  NAND2_X1 U7807 ( .A1(n9452), .A2(n9055), .ZN(n9304) );
  NAND2_X1 U7808 ( .A1(n9302), .A2(n9304), .ZN(n9324) );
  INV_X1 U7809 ( .A(n9324), .ZN(n9326) );
  INV_X1 U7810 ( .A(n9369), .ZN(n9330) );
  INV_X1 U7811 ( .A(n7967), .ZN(n6448) );
  AND2_X1 U7812 ( .A1(n9455), .A2(n9330), .ZN(n7968) );
  INV_X1 U7813 ( .A(n9383), .ZN(n9083) );
  OR2_X1 U7814 ( .A1(n9460), .A2(n9083), .ZN(n6426) );
  NAND2_X1 U7815 ( .A1(n9460), .A2(n9083), .ZN(n7966) );
  INV_X1 U7816 ( .A(n7964), .ZN(n9364) );
  OR2_X1 U7817 ( .A1(n9465), .A2(n9037), .ZN(n6425) );
  NAND2_X1 U7818 ( .A1(n9465), .A2(n9037), .ZN(n9365) );
  NAND2_X1 U7819 ( .A1(n6425), .A2(n9365), .ZN(n9381) );
  INV_X1 U7820 ( .A(n9384), .ZN(n9027) );
  OR2_X1 U7821 ( .A1(n9470), .A2(n9027), .ZN(n9379) );
  NAND2_X1 U7822 ( .A1(n9470), .A2(n9027), .ZN(n6421) );
  OR2_X1 U7823 ( .A1(n7939), .A2(n9110), .ZN(n6418) );
  NAND2_X1 U7824 ( .A1(n7939), .A2(n9110), .ZN(n9397) );
  INV_X1 U7825 ( .A(n9120), .ZN(n7866) );
  OR2_X1 U7826 ( .A1(n9476), .A2(n7866), .ZN(n7871) );
  NAND2_X1 U7827 ( .A1(n9476), .A2(n7866), .ZN(n6407) );
  NAND2_X1 U7828 ( .A1(n7871), .A2(n6407), .ZN(n7840) );
  INV_X1 U7829 ( .A(n9121), .ZN(n7852) );
  OR2_X1 U7830 ( .A1(n7868), .A2(n7852), .ZN(n6350) );
  NAND2_X1 U7831 ( .A1(n7868), .A2(n7852), .ZN(n7838) );
  INV_X1 U7832 ( .A(n7836), .ZN(n6317) );
  OR2_X1 U7833 ( .A1(n9482), .A2(n7787), .ZN(n6392) );
  NAND2_X1 U7834 ( .A1(n9482), .A2(n7787), .ZN(n7780) );
  NAND2_X1 U7835 ( .A1(n6392), .A2(n7780), .ZN(n7785) );
  INV_X1 U7836 ( .A(n9133), .ZN(n6305) );
  NAND2_X1 U7837 ( .A1(n9133), .A2(n6618), .ZN(n6491) );
  INV_X1 U7838 ( .A(n6306), .ZN(n6307) );
  NAND2_X1 U7839 ( .A1(n6307), .A2(n7109), .ZN(n7227) );
  AND2_X1 U7840 ( .A1(n7228), .A2(n7227), .ZN(n7229) );
  NAND2_X1 U7841 ( .A1(n6309), .A2(n6308), .ZN(n6495) );
  INV_X1 U7842 ( .A(n7262), .ZN(n9130) );
  NAND2_X1 U7843 ( .A1(n9131), .A2(n9706), .ZN(n6377) );
  NAND2_X1 U7844 ( .A1(n6379), .A2(n6377), .ZN(n6335) );
  INV_X1 U7845 ( .A(n7109), .ZN(n7225) );
  AND2_X1 U7846 ( .A1(n6306), .A2(n7225), .ZN(n6490) );
  NOR3_X1 U7847 ( .A1(n6934), .A2(n6335), .A3(n6490), .ZN(n6311) );
  INV_X1 U7848 ( .A(n7441), .ZN(n9129) );
  NAND2_X1 U7849 ( .A1(n9129), .A2(n6310), .ZN(n6623) );
  NAND2_X1 U7850 ( .A1(n9128), .A2(n7296), .ZN(n6380) );
  AND2_X1 U7851 ( .A1(n6623), .A2(n6380), .ZN(n7289) );
  NAND2_X1 U7852 ( .A1(n7300), .A2(n7487), .ZN(n7292) );
  INV_X1 U7853 ( .A(n7300), .ZN(n9127) );
  NAND2_X1 U7854 ( .A1(n9127), .A2(n7469), .ZN(n6500) );
  INV_X1 U7855 ( .A(n7387), .ZN(n7291) );
  NAND4_X1 U7856 ( .A1(n7229), .A2(n6311), .A3(n7289), .A4(n7291), .ZN(n6312)
         );
  NAND2_X1 U7857 ( .A1(n7297), .A2(n7440), .ZN(n7382) );
  NAND2_X1 U7858 ( .A1(n7441), .A2(n9680), .ZN(n6624) );
  AND2_X1 U7859 ( .A1(n7382), .A2(n6624), .ZN(n6337) );
  NAND2_X1 U7860 ( .A1(n7262), .A2(n7144), .ZN(n6378) );
  AND2_X1 U7861 ( .A1(n6337), .A2(n6378), .ZN(n6502) );
  NAND2_X1 U7862 ( .A1(n7134), .A2(n7124), .ZN(n6496) );
  NAND2_X1 U7863 ( .A1(n6502), .A2(n6496), .ZN(n6336) );
  NAND2_X1 U7864 ( .A1(n7480), .A2(n7538), .ZN(n6398) );
  NAND2_X1 U7865 ( .A1(n9126), .A2(n7411), .ZN(n7368) );
  NAND2_X1 U7866 ( .A1(n6398), .A2(n7368), .ZN(n7302) );
  NOR3_X1 U7867 ( .A1(n6312), .A2(n6336), .A3(n7302), .ZN(n6315) );
  NAND2_X1 U7868 ( .A1(n7685), .A2(n7620), .ZN(n6387) );
  NAND2_X1 U7869 ( .A1(n7618), .A2(n6387), .ZN(n7611) );
  INV_X1 U7870 ( .A(n7611), .ZN(n6314) );
  INV_X1 U7871 ( .A(n9125), .ZN(n7295) );
  NAND2_X1 U7872 ( .A1(n7295), .A2(n7520), .ZN(n7499) );
  INV_X1 U7873 ( .A(n7499), .ZN(n6400) );
  INV_X1 U7874 ( .A(n7520), .ZN(n9715) );
  AND2_X1 U7875 ( .A1(n9715), .A2(n9125), .ZN(n7497) );
  NOR2_X1 U7876 ( .A1(n6400), .A2(n7497), .ZN(n7370) );
  NOR2_X1 U7877 ( .A1(n7629), .A2(n9123), .ZN(n7756) );
  NAND2_X1 U7878 ( .A1(n7629), .A2(n9123), .ZN(n7757) );
  INV_X1 U7879 ( .A(n7757), .ZN(n6313) );
  OR2_X1 U7880 ( .A1(n7756), .A2(n6313), .ZN(n7619) );
  NAND4_X1 U7881 ( .A1(n6315), .A2(n6314), .A3(n7370), .A4(n7619), .ZN(n6316)
         );
  NOR4_X1 U7882 ( .A1(n7840), .A2(n6317), .A3(n7785), .A4(n6316), .ZN(n6318)
         );
  AND2_X1 U7883 ( .A1(n9113), .A2(n9119), .ZN(n7911) );
  OR2_X1 U7884 ( .A1(n4366), .A2(n7911), .ZN(n7880) );
  NAND4_X1 U7885 ( .A1(n9399), .A2(n7913), .A3(n6318), .A4(n7880), .ZN(n6319)
         );
  NOR4_X1 U7886 ( .A1(n9351), .A2(n9364), .A3(n9381), .A4(n6319), .ZN(n6320)
         );
  NAND4_X1 U7887 ( .A1(n9288), .A2(n9305), .A3(n9326), .A4(n6320), .ZN(n6321)
         );
  NOR4_X1 U7888 ( .A1(n9228), .A2(n9271), .A3(n9263), .A4(n6321), .ZN(n6322)
         );
  XNOR2_X1 U7889 ( .A(n9424), .B(n9264), .ZN(n9247) );
  NAND4_X1 U7890 ( .A1(n9203), .A2(n7979), .A3(n6322), .A4(n9247), .ZN(n6324)
         );
  AND2_X1 U7891 ( .A1(n9198), .A2(n6323), .ZN(n6519) );
  NOR4_X1 U7892 ( .A1(n6524), .A2(n6326), .A3(n6324), .A4(n6519), .ZN(n6325)
         );
  NOR2_X1 U7893 ( .A1(n6325), .A2(n6775), .ZN(n6484) );
  NAND2_X1 U7894 ( .A1(n6326), .A2(n9193), .ZN(n6480) );
  INV_X1 U7895 ( .A(n9264), .ZN(n9230) );
  NAND2_X1 U7896 ( .A1(n9424), .A2(n9230), .ZN(n7975) );
  INV_X1 U7897 ( .A(n7975), .ZN(n6327) );
  NAND2_X1 U7898 ( .A1(n7977), .A2(n6327), .ZN(n6328) );
  NAND3_X1 U7899 ( .A1(n7978), .A2(n6372), .A3(n6328), .ZN(n6518) );
  OR2_X1 U7900 ( .A1(n9424), .A2(n9230), .ZN(n6456) );
  AND2_X1 U7901 ( .A1(n6456), .A2(n9244), .ZN(n7974) );
  NOR2_X1 U7902 ( .A1(n6518), .A2(n7974), .ZN(n6331) );
  INV_X1 U7903 ( .A(n6374), .ZN(n6329) );
  OR3_X1 U7904 ( .A1(n6331), .A2(n6330), .A3(n6329), .ZN(n6523) );
  NAND2_X1 U7905 ( .A1(n9302), .A2(n7968), .ZN(n6332) );
  AND2_X1 U7906 ( .A1(n6332), .A2(n9304), .ZN(n6333) );
  NAND2_X1 U7907 ( .A1(n6333), .A2(n6449), .ZN(n6435) );
  INV_X1 U7908 ( .A(n7966), .ZN(n6427) );
  NOR2_X1 U7909 ( .A1(n6435), .A2(n6427), .ZN(n6508) );
  AND2_X1 U7910 ( .A1(n6421), .A2(n9397), .ZN(n7962) );
  INV_X1 U7911 ( .A(n9123), .ZN(n7763) );
  NAND2_X1 U7912 ( .A1(n7629), .A2(n7763), .ZN(n7758) );
  AND2_X1 U7913 ( .A1(n7780), .A2(n7758), .ZN(n6389) );
  AND2_X1 U7914 ( .A1(n6387), .A2(n7499), .ZN(n7616) );
  AND2_X1 U7915 ( .A1(n7292), .A2(n6398), .ZN(n7366) );
  AND2_X1 U7916 ( .A1(n7616), .A2(n7366), .ZN(n6384) );
  AND4_X1 U7917 ( .A1(n6407), .A2(n6389), .A3(n6384), .A4(n7838), .ZN(n6334)
         );
  INV_X1 U7918 ( .A(n9119), .ZN(n7902) );
  NAND2_X1 U7919 ( .A1(n9113), .A2(n7902), .ZN(n7908) );
  NAND4_X1 U7920 ( .A1(n9365), .A2(n7962), .A3(n6334), .A4(n7908), .ZN(n6506)
         );
  NAND2_X1 U7921 ( .A1(n6494), .A2(n6491), .ZN(n6935) );
  INV_X1 U7922 ( .A(n6335), .ZN(n6498) );
  NAND2_X1 U7923 ( .A1(n7116), .A2(n6498), .ZN(n6342) );
  INV_X1 U7924 ( .A(n6336), .ZN(n6341) );
  INV_X1 U7925 ( .A(n6337), .ZN(n6339) );
  AND2_X1 U7926 ( .A1(n6379), .A2(n6623), .ZN(n6338) );
  AND2_X1 U7927 ( .A1(n6500), .A2(n6380), .ZN(n6381) );
  OAI21_X1 U7928 ( .B1(n6339), .B2(n6338), .A(n6381), .ZN(n6340) );
  AOI21_X1 U7929 ( .B1(n6342), .B2(n6341), .A(n6340), .ZN(n6356) );
  INV_X1 U7930 ( .A(n6418), .ZN(n6355) );
  NOR2_X1 U7931 ( .A1(n9113), .A2(n7902), .ZN(n7906) );
  INV_X1 U7932 ( .A(n7906), .ZN(n6353) );
  INV_X1 U7933 ( .A(n7368), .ZN(n6343) );
  OR2_X1 U7934 ( .A1(n7497), .A2(n6343), .ZN(n6344) );
  NAND2_X1 U7935 ( .A1(n7616), .A2(n6344), .ZN(n6345) );
  NAND2_X1 U7936 ( .A1(n6345), .A2(n7618), .ZN(n6383) );
  INV_X1 U7937 ( .A(n6383), .ZN(n6348) );
  INV_X1 U7938 ( .A(n6389), .ZN(n6347) );
  OR2_X1 U7939 ( .A1(n7629), .A2(n7763), .ZN(n7760) );
  AND2_X1 U7940 ( .A1(n6392), .A2(n7760), .ZN(n7778) );
  INV_X1 U7941 ( .A(n7780), .ZN(n6346) );
  OR2_X1 U7942 ( .A1(n7778), .A2(n6346), .ZN(n6404) );
  OAI21_X1 U7943 ( .B1(n6348), .B2(n6347), .A(n6404), .ZN(n6349) );
  AND2_X1 U7944 ( .A1(n6349), .A2(n7838), .ZN(n6351) );
  AND2_X1 U7945 ( .A1(n7871), .A2(n6350), .ZN(n6409) );
  INV_X1 U7946 ( .A(n6409), .ZN(n6394) );
  OAI211_X1 U7947 ( .C1(n6351), .C2(n6394), .A(n7908), .B(n6407), .ZN(n6352)
         );
  NAND2_X1 U7948 ( .A1(n6353), .A2(n6352), .ZN(n6354) );
  OAI211_X1 U7949 ( .C1(n6355), .C2(n6354), .A(n9365), .B(n7962), .ZN(n6504)
         );
  OAI21_X1 U7950 ( .B1(n6506), .B2(n6356), .A(n6504), .ZN(n6362) );
  AND2_X1 U7951 ( .A1(n6425), .A2(n9379), .ZN(n7963) );
  AND2_X1 U7952 ( .A1(n7966), .A2(n9365), .ZN(n6431) );
  INV_X1 U7953 ( .A(n6431), .ZN(n6358) );
  NAND2_X1 U7954 ( .A1(n7967), .A2(n6426), .ZN(n6430) );
  INV_X1 U7955 ( .A(n6430), .ZN(n6357) );
  OAI211_X1 U7956 ( .C1(n7963), .C2(n6358), .A(n9302), .B(n6357), .ZN(n6359)
         );
  INV_X1 U7957 ( .A(n6359), .ZN(n6360) );
  OR2_X1 U7958 ( .A1(n6435), .A2(n6360), .ZN(n6361) );
  NAND2_X1 U7959 ( .A1(n6361), .A2(n6447), .ZN(n6509) );
  AOI21_X1 U7960 ( .B1(n6508), .B2(n6362), .A(n6509), .ZN(n6363) );
  OAI21_X1 U7961 ( .B1(n6363), .B2(n4622), .A(n7972), .ZN(n6364) );
  NAND2_X1 U7962 ( .A1(n7973), .A2(n6364), .ZN(n6365) );
  AOI21_X1 U7963 ( .B1(n7977), .B2(n6365), .A(n6518), .ZN(n6369) );
  INV_X1 U7964 ( .A(n6366), .ZN(n6520) );
  INV_X1 U7965 ( .A(n6367), .ZN(n9195) );
  NAND2_X1 U7966 ( .A1(n9195), .A2(n9117), .ZN(n6368) );
  NAND2_X1 U7967 ( .A1(n9198), .A2(n6368), .ZN(n6478) );
  OAI211_X1 U7968 ( .C1(n6523), .C2(n6369), .A(n6520), .B(n6478), .ZN(n6370)
         );
  AOI211_X1 U7969 ( .C1(n6480), .C2(n6370), .A(n7342), .B(n6524), .ZN(n6371)
         );
  OR2_X1 U7970 ( .A1(n6484), .A2(n6371), .ZN(n6485) );
  MUX2_X1 U7971 ( .A(n7977), .B(n6372), .S(n6472), .Z(n6373) );
  NAND2_X1 U7972 ( .A1(n9203), .A2(n6373), .ZN(n6376) );
  MUX2_X1 U7973 ( .A(n7978), .B(n6374), .S(n6472), .Z(n6375) );
  NAND2_X1 U7974 ( .A1(n6376), .A2(n6375), .ZN(n6465) );
  NAND2_X1 U7975 ( .A1(n6378), .A2(n6379), .ZN(n7138) );
  OR2_X2 U7976 ( .A1(n7137), .A2(n7138), .ZN(n7135) );
  NAND2_X1 U7977 ( .A1(n7290), .A2(n6623), .ZN(n6613) );
  NAND2_X1 U7978 ( .A1(n6613), .A2(n6627), .ZN(n6382) );
  NAND2_X1 U7979 ( .A1(n6382), .A2(n6381), .ZN(n6385) );
  AOI21_X1 U7980 ( .B1(n6385), .B2(n6384), .A(n6383), .ZN(n6386) );
  MUX2_X1 U7981 ( .A(n6387), .B(n6386), .S(n6472), .Z(n6388) );
  AND2_X1 U7982 ( .A1(n6388), .A2(n7619), .ZN(n6403) );
  INV_X1 U7983 ( .A(n6403), .ZN(n6390) );
  NAND2_X1 U7984 ( .A1(n6390), .A2(n6389), .ZN(n6393) );
  INV_X1 U7985 ( .A(n7838), .ZN(n6391) );
  OAI21_X1 U7986 ( .B1(n6395), .B2(n6394), .A(n6407), .ZN(n6412) );
  INV_X1 U7987 ( .A(n6627), .ZN(n6396) );
  OAI211_X1 U7988 ( .C1(n6613), .C2(n6396), .A(n7382), .B(n7292), .ZN(n6397)
         );
  NAND3_X1 U7989 ( .A1(n6397), .A2(n6500), .A3(n7368), .ZN(n6399) );
  AOI21_X1 U7990 ( .B1(n6399), .B2(n6398), .A(n7497), .ZN(n6401) );
  OAI21_X1 U7991 ( .B1(n6401), .B2(n6400), .A(n7618), .ZN(n6402) );
  NAND3_X1 U7992 ( .A1(n6403), .A2(n7780), .A3(n6402), .ZN(n6405) );
  NAND2_X1 U7993 ( .A1(n6405), .A2(n6404), .ZN(n6406) );
  NAND2_X1 U7994 ( .A1(n6406), .A2(n7838), .ZN(n6410) );
  INV_X1 U7995 ( .A(n6407), .ZN(n6408) );
  AOI21_X1 U7996 ( .B1(n6410), .B2(n6409), .A(n6408), .ZN(n6411) );
  MUX2_X1 U7997 ( .A(n6412), .B(n6411), .S(n6471), .Z(n6413) );
  NAND2_X1 U7998 ( .A1(n6413), .A2(n7880), .ZN(n6417) );
  INV_X1 U7999 ( .A(n7908), .ZN(n6414) );
  MUX2_X1 U8000 ( .A(n7906), .B(n6414), .S(n6472), .Z(n6415) );
  INV_X1 U8001 ( .A(n6415), .ZN(n6416) );
  NAND3_X1 U8002 ( .A1(n6417), .A2(n7913), .A3(n6416), .ZN(n6420) );
  MUX2_X1 U8003 ( .A(n6418), .B(n9397), .S(n6471), .Z(n6419) );
  NAND3_X1 U8004 ( .A1(n6420), .A2(n9399), .A3(n6419), .ZN(n6424) );
  AND2_X1 U8005 ( .A1(n9365), .A2(n6421), .ZN(n6422) );
  MUX2_X1 U8006 ( .A(n6422), .B(n7963), .S(n6471), .Z(n6423) );
  NAND2_X1 U8007 ( .A1(n6424), .A2(n6423), .ZN(n6432) );
  AND2_X1 U8008 ( .A1(n6426), .A2(n6425), .ZN(n6429) );
  OR2_X1 U8009 ( .A1(n7968), .A2(n6427), .ZN(n6428) );
  AOI21_X1 U8010 ( .B1(n6432), .B2(n6429), .A(n6428), .ZN(n6434) );
  AOI21_X1 U8011 ( .B1(n6432), .B2(n6431), .A(n6430), .ZN(n6433) );
  MUX2_X1 U8012 ( .A(n6434), .B(n6433), .S(n6471), .Z(n6452) );
  AOI21_X1 U8013 ( .B1(n6452), .B2(n9302), .A(n6435), .ZN(n6437) );
  INV_X1 U8014 ( .A(n6447), .ZN(n6436) );
  OAI211_X1 U8015 ( .C1(n6437), .C2(n6436), .A(n9274), .B(n7971), .ZN(n6440)
         );
  INV_X1 U8016 ( .A(n7972), .ZN(n6438) );
  NAND2_X1 U8017 ( .A1(n6438), .A2(n9260), .ZN(n6439) );
  NAND3_X1 U8018 ( .A1(n6440), .A2(n9244), .A3(n6439), .ZN(n6445) );
  NAND2_X1 U8019 ( .A1(n6441), .A2(n6471), .ZN(n6443) );
  AND2_X1 U8020 ( .A1(n9264), .A2(n6471), .ZN(n6459) );
  NAND2_X1 U8021 ( .A1(n6441), .A2(n6459), .ZN(n6442) );
  OAI21_X1 U8022 ( .B1(n6443), .B2(n9424), .A(n6442), .ZN(n6444) );
  NAND2_X1 U8023 ( .A1(n6445), .A2(n6444), .ZN(n6462) );
  INV_X1 U8024 ( .A(n6446), .ZN(n6455) );
  NAND2_X1 U8025 ( .A1(n6447), .A2(n9302), .ZN(n7969) );
  OR2_X1 U8026 ( .A1(n7969), .A2(n6448), .ZN(n6451) );
  OR2_X1 U8027 ( .A1(n7969), .A2(n9304), .ZN(n6450) );
  OAI21_X1 U8028 ( .B1(n6452), .B2(n6451), .A(n7970), .ZN(n6453) );
  NAND3_X1 U8029 ( .A1(n6453), .A2(n9274), .A3(n9272), .ZN(n6454) );
  OAI211_X1 U8030 ( .C1(n6455), .C2(n7971), .A(n7973), .B(n6454), .ZN(n6457)
         );
  NAND4_X1 U8031 ( .A1(n6457), .A2(n6472), .A3(n9244), .A4(n6456), .ZN(n6461)
         );
  OAI21_X1 U8032 ( .B1(n9264), .B2(n6471), .A(n9424), .ZN(n6458) );
  OAI21_X1 U8033 ( .B1(n6459), .B2(n9424), .A(n6458), .ZN(n6460) );
  NAND3_X1 U8034 ( .A1(n6462), .A2(n6461), .A3(n6460), .ZN(n6463) );
  NAND3_X1 U8035 ( .A1(n9203), .A2(n7959), .A3(n6463), .ZN(n6464) );
  AND2_X1 U8036 ( .A1(n6465), .A2(n6464), .ZN(n6475) );
  AND2_X1 U8037 ( .A1(n6475), .A2(n6478), .ZN(n6466) );
  NAND2_X1 U8038 ( .A1(n6480), .A2(n6466), .ZN(n6470) );
  INV_X1 U8039 ( .A(n7986), .ZN(n7993) );
  INV_X1 U8040 ( .A(n6467), .ZN(n6468) );
  OAI22_X1 U8041 ( .A1(n6470), .A2(n7993), .B1(n6468), .B2(n6478), .ZN(n6469)
         );
  OAI21_X1 U8042 ( .B1(n6470), .B2(n9209), .A(n6480), .ZN(n6473) );
  NOR2_X1 U8043 ( .A1(n9209), .A2(n6472), .ZN(n6474) );
  AOI21_X1 U8044 ( .B1(n7986), .B2(n6472), .A(n6474), .ZN(n6479) );
  INV_X1 U8045 ( .A(n6475), .ZN(n6476) );
  NAND3_X1 U8046 ( .A1(n6476), .A2(n7993), .A3(n9209), .ZN(n6477) );
  NAND4_X1 U8047 ( .A1(n6480), .A2(n6479), .A3(n6478), .A4(n6477), .ZN(n6481)
         );
  AND3_X2 U8048 ( .A1(n6483), .A2(n6482), .A3(n4895), .ZN(n6486) );
  INV_X1 U8049 ( .A(n6486), .ZN(n6488) );
  NAND4_X1 U8050 ( .A1(n6488), .A2(n6775), .A3(n6487), .A4(n6241), .ZN(n6489)
         );
  INV_X1 U8051 ( .A(n6326), .ZN(n6526) );
  INV_X1 U8052 ( .A(n6490), .ZN(n6779) );
  AND2_X1 U8053 ( .A1(n6779), .A2(n6775), .ZN(n6493) );
  OAI211_X1 U8054 ( .C1(n6494), .C2(n6493), .A(n6492), .B(n6491), .ZN(n6497)
         );
  NAND3_X1 U8055 ( .A1(n6497), .A2(n6496), .A3(n6495), .ZN(n6499) );
  NAND2_X1 U8056 ( .A1(n6499), .A2(n6498), .ZN(n6503) );
  OAI21_X1 U8057 ( .B1(n4615), .B2(n7289), .A(n6500), .ZN(n6501) );
  AOI21_X1 U8058 ( .B1(n6503), .B2(n6502), .A(n6501), .ZN(n6505) );
  OAI21_X1 U8059 ( .B1(n6506), .B2(n6505), .A(n6504), .ZN(n6507) );
  INV_X1 U8060 ( .A(n6507), .ZN(n6512) );
  INV_X1 U8061 ( .A(n6508), .ZN(n6511) );
  INV_X1 U8062 ( .A(n6509), .ZN(n6510) );
  OAI21_X1 U8063 ( .B1(n6512), .B2(n6511), .A(n6510), .ZN(n6513) );
  NAND2_X1 U8064 ( .A1(n6513), .A2(n7971), .ZN(n6514) );
  NAND2_X1 U8065 ( .A1(n7972), .A2(n6514), .ZN(n6515) );
  NAND2_X1 U8066 ( .A1(n7973), .A2(n6515), .ZN(n6516) );
  AND2_X1 U8067 ( .A1(n7959), .A2(n6516), .ZN(n6517) );
  NOR2_X1 U8068 ( .A1(n6518), .A2(n6517), .ZN(n6522) );
  INV_X1 U8069 ( .A(n6519), .ZN(n6521) );
  OAI211_X1 U8070 ( .C1(n6523), .C2(n6522), .A(n6521), .B(n6520), .ZN(n6525)
         );
  AOI21_X1 U8071 ( .B1(n6526), .B2(n6525), .A(n6524), .ZN(n6529) );
  INV_X1 U8072 ( .A(n6529), .ZN(n6528) );
  NOR2_X1 U8073 ( .A1(n6528), .A2(n6527), .ZN(n6534) );
  NOR2_X1 U8074 ( .A1(n6529), .A2(n9682), .ZN(n6530) );
  NAND2_X1 U8075 ( .A1(n6530), .A2(n7936), .ZN(n6532) );
  OR2_X1 U8076 ( .A1(n6545), .A2(P1_U3084), .ZN(n7678) );
  INV_X1 U8077 ( .A(n7678), .ZN(n6531) );
  NOR2_X1 U8078 ( .A1(n6614), .A2(n7678), .ZN(n6535) );
  NOR2_X1 U8079 ( .A1(n6535), .A2(n7982), .ZN(n6536) );
  OR2_X1 U8080 ( .A1(n6540), .A2(P2_U3152), .ZN(n7771) );
  OR2_X1 U8081 ( .A1(n7771), .A2(n6541), .ZN(n6859) );
  INV_X2 U8082 ( .A(n8370), .ZN(P2_U3966) );
  INV_X1 U8083 ( .A(n6545), .ZN(n6542) );
  NOR2_X1 U8084 ( .A1(n6543), .A2(n6542), .ZN(n6576) );
  OR2_X1 U8085 ( .A1(n6631), .A2(n6544), .ZN(n6546) );
  NAND2_X1 U8086 ( .A1(n6546), .A2(n6545), .ZN(n6606) );
  NAND2_X1 U8087 ( .A1(n6606), .A2(n5801), .ZN(n6547) );
  NAND2_X1 U8088 ( .A1(n6547), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  INV_X1 U8089 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7791) );
  NOR2_X1 U8090 ( .A1(n6855), .A2(n7791), .ZN(n6548) );
  AOI21_X1 U8091 ( .B1(n7791), .B2(n6855), .A(n6548), .ZN(n6852) );
  NAND2_X1 U8092 ( .A1(n9630), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6569) );
  INV_X1 U8093 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n6549) );
  MUX2_X1 U8094 ( .A(n6549), .B(P1_REG2_REG_10__SCAN_IN), .S(n9630), .Z(n6550)
         );
  INV_X1 U8095 ( .A(n6550), .ZN(n9637) );
  NAND2_X1 U8096 ( .A1(n9624), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6568) );
  INV_X1 U8097 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n6551) );
  MUX2_X1 U8098 ( .A(n6551), .B(P1_REG2_REG_9__SCAN_IN), .S(n6681), .Z(n9626)
         );
  INV_X1 U8099 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n6565) );
  INV_X1 U8100 ( .A(n6732), .ZN(n6669) );
  AOI22_X1 U8101 ( .A1(P1_REG2_REG_7__SCAN_IN), .A2(n6669), .B1(n6732), .B2(
        n6565), .ZN(n6724) );
  NAND2_X1 U8102 ( .A1(n6580), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6564) );
  NOR2_X1 U8103 ( .A1(n6590), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6561) );
  INV_X1 U8104 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6552) );
  MUX2_X1 U8105 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n6552), .S(n6670), .Z(n9613)
         );
  INV_X1 U8106 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6553) );
  MUX2_X1 U8107 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n6553), .S(n6664), .Z(n9142)
         );
  AND2_X1 U8108 ( .A1(P1_REG2_REG_0__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n9143) );
  NAND2_X1 U8109 ( .A1(n9142), .A2(n9143), .ZN(n9141) );
  NAND2_X1 U8110 ( .A1(n6664), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6554) );
  NAND2_X1 U8111 ( .A1(n9141), .A2(n6554), .ZN(n9614) );
  NAND2_X1 U8112 ( .A1(n9613), .A2(n9614), .ZN(n9612) );
  NAND2_X1 U8113 ( .A1(n6670), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n9152) );
  NAND2_X1 U8114 ( .A1(n9612), .A2(n9152), .ZN(n6557) );
  INV_X1 U8115 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6555) );
  MUX2_X1 U8116 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n6555), .S(n9150), .Z(n6556)
         );
  NAND2_X1 U8117 ( .A1(n6557), .A2(n6556), .ZN(n9154) );
  NAND2_X1 U8118 ( .A1(n9150), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6558) );
  AND2_X1 U8119 ( .A1(n9154), .A2(n6558), .ZN(n6784) );
  INV_X1 U8120 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n7176) );
  MUX2_X1 U8121 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n7176), .S(n6808), .Z(n6559)
         );
  NAND2_X1 U8122 ( .A1(n6784), .A2(n6559), .ZN(n6795) );
  INV_X1 U8123 ( .A(n6795), .ZN(n6560) );
  NOR2_X1 U8124 ( .A1(n6808), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6792) );
  NOR2_X1 U8125 ( .A1(n6560), .A2(n6792), .ZN(n6743) );
  INV_X1 U8126 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n9947) );
  AOI22_X1 U8127 ( .A1(n6590), .A2(n9947), .B1(P1_REG2_REG_5__SCAN_IN), .B2(
        n6744), .ZN(n6742) );
  NOR2_X1 U8128 ( .A1(n6743), .A2(n6742), .ZN(n6741) );
  NOR2_X1 U8129 ( .A1(n6561), .A2(n6741), .ZN(n6714) );
  INV_X1 U8130 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6562) );
  MUX2_X1 U8131 ( .A(n6562), .B(P1_REG2_REG_6__SCAN_IN), .S(n6580), .Z(n6563)
         );
  INV_X1 U8132 ( .A(n6563), .ZN(n6713) );
  NAND2_X1 U8133 ( .A1(n6714), .A2(n6713), .ZN(n6712) );
  NAND2_X1 U8134 ( .A1(n6564), .A2(n6712), .ZN(n6725) );
  NOR2_X1 U8135 ( .A1(n6724), .A2(n6725), .ZN(n6723) );
  AOI21_X1 U8136 ( .B1(n6565), .B2(n6669), .A(n6723), .ZN(n6754) );
  INV_X1 U8137 ( .A(n6595), .ZN(n6760) );
  INV_X1 U8138 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n6566) );
  AOI22_X1 U8139 ( .A1(P1_REG2_REG_8__SCAN_IN), .A2(n6760), .B1(n6595), .B2(
        n6566), .ZN(n6753) );
  NOR2_X1 U8140 ( .A1(n6754), .A2(n6753), .ZN(n6752) );
  NOR2_X1 U8141 ( .A1(n6595), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6567) );
  NOR2_X1 U8142 ( .A1(n6752), .A2(n6567), .ZN(n9627) );
  NAND2_X1 U8143 ( .A1(n9626), .A2(n9627), .ZN(n9625) );
  NAND2_X1 U8144 ( .A1(n6568), .A2(n9625), .ZN(n9638) );
  NAND2_X1 U8145 ( .A1(n9637), .A2(n9638), .ZN(n9636) );
  NAND2_X1 U8146 ( .A1(n6569), .A2(n9636), .ZN(n9657) );
  INV_X1 U8147 ( .A(n9657), .ZN(n6570) );
  INV_X1 U8148 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n9890) );
  NOR2_X1 U8149 ( .A1(n6570), .A2(n9890), .ZN(n6571) );
  OAI22_X1 U8150 ( .A1(n6571), .A2(n9650), .B1(P1_REG2_REG_11__SCAN_IN), .B2(
        n9657), .ZN(n9655) );
  NAND2_X1 U8151 ( .A1(n6604), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n6572) );
  OAI21_X1 U8152 ( .B1(n6604), .B2(P1_REG2_REG_12__SCAN_IN), .A(n6572), .ZN(
        n6925) );
  NOR2_X1 U8153 ( .A1(n9655), .A2(n6925), .ZN(n6924) );
  AOI21_X1 U8154 ( .B1(n6604), .B2(P1_REG2_REG_12__SCAN_IN), .A(n6924), .ZN(
        n6851) );
  NOR2_X1 U8155 ( .A1(n6852), .A2(n6851), .ZN(n6850) );
  AOI21_X1 U8156 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n6855), .A(n6850), .ZN(
        n6573) );
  INV_X1 U8157 ( .A(n9663), .ZN(n6740) );
  NAND2_X1 U8158 ( .A1(n6573), .A2(n6740), .ZN(n6574) );
  XNOR2_X1 U8159 ( .A(n6573), .B(n9663), .ZN(n9667) );
  INV_X1 U8160 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n9666) );
  NAND2_X1 U8161 ( .A1(n9667), .A2(n9666), .ZN(n9665) );
  NAND2_X1 U8162 ( .A1(n6574), .A2(n9665), .ZN(n7416) );
  XNOR2_X1 U8163 ( .A(n7416), .B(n7422), .ZN(n6575) );
  INV_X1 U8164 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9943) );
  NOR2_X1 U8165 ( .A1(n9943), .A2(n6575), .ZN(n7417) );
  NOR2_X1 U8166 ( .A1(n7983), .A2(P1_U3084), .ZN(n7892) );
  AND2_X1 U8167 ( .A1(n6606), .A2(n7892), .ZN(n9643) );
  NAND2_X1 U8168 ( .A1(n9643), .A2(n6803), .ZN(n9182) );
  AOI211_X1 U8169 ( .C1(n6575), .C2(n9943), .A(n7417), .B(n9182), .ZN(n6612)
         );
  OR2_X1 U8170 ( .A1(P1_U3083), .A2(n6576), .ZN(n9678) );
  INV_X1 U8171 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n6577) );
  NOR2_X1 U8172 ( .A1(n9678), .A2(n6577), .ZN(n6611) );
  INV_X1 U8173 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n6578) );
  AOI22_X1 U8174 ( .A1(n9663), .A2(P1_REG1_REG_14__SCAN_IN), .B1(n6578), .B2(
        n6740), .ZN(n9669) );
  INV_X1 U8175 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n9580) );
  INV_X1 U8176 ( .A(n6855), .ZN(n6719) );
  NOR2_X1 U8177 ( .A1(n6719), .A2(n9580), .ZN(n6579) );
  AOI21_X1 U8178 ( .B1(n9580), .B2(n6719), .A(n6579), .ZN(n6849) );
  INV_X1 U8179 ( .A(n9650), .ZN(n9654) );
  INV_X1 U8180 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n6601) );
  OR2_X1 U8181 ( .A1(n9630), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6600) );
  NOR2_X1 U8182 ( .A1(n9624), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6597) );
  INV_X1 U8183 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6596) );
  INV_X1 U8184 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6594) );
  NOR2_X1 U8185 ( .A1(n6580), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6593) );
  INV_X1 U8186 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n7191) );
  AOI22_X1 U8187 ( .A1(n6580), .A2(n7191), .B1(P1_REG1_REG_6__SCAN_IN), .B2(
        n6710), .ZN(n6708) );
  NAND2_X1 U8188 ( .A1(n6590), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6592) );
  XNOR2_X1 U8189 ( .A(n6670), .B(P1_REG1_REG_2__SCAN_IN), .ZN(n9606) );
  INV_X1 U8190 ( .A(n9606), .ZN(n6583) );
  INV_X1 U8191 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6581) );
  MUX2_X1 U8192 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n6581), .S(n6664), .Z(n9139)
         );
  AND2_X1 U8193 ( .A1(P1_REG1_REG_0__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n9140) );
  NAND2_X1 U8194 ( .A1(n9139), .A2(n9140), .ZN(n9138) );
  NAND2_X1 U8195 ( .A1(n6664), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6582) );
  NAND2_X1 U8196 ( .A1(n9138), .A2(n6582), .ZN(n9607) );
  NAND2_X1 U8197 ( .A1(n6583), .A2(n9607), .ZN(n6585) );
  NAND2_X1 U8198 ( .A1(n6670), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6584) );
  NAND2_X1 U8199 ( .A1(n6585), .A2(n6584), .ZN(n9156) );
  INV_X1 U8200 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6586) );
  MUX2_X1 U8201 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n6586), .S(n9150), .Z(n9157)
         );
  NAND2_X1 U8202 ( .A1(n9156), .A2(n9157), .ZN(n9155) );
  NAND2_X1 U8203 ( .A1(n9150), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6587) );
  NAND2_X1 U8204 ( .A1(n9155), .A2(n6587), .ZN(n6789) );
  MUX2_X1 U8205 ( .A(n10040), .B(P1_REG1_REG_4__SCAN_IN), .S(n6808), .Z(n6588)
         );
  OR2_X1 U8206 ( .A1(n6789), .A2(n6588), .ZN(n6791) );
  NOR2_X1 U8207 ( .A1(n6808), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6788) );
  INV_X1 U8208 ( .A(n6788), .ZN(n6589) );
  NAND2_X1 U8209 ( .A1(n6791), .A2(n6589), .ZN(n6747) );
  INV_X1 U8210 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n7259) );
  MUX2_X1 U8211 ( .A(n7259), .B(P1_REG1_REG_5__SCAN_IN), .S(n6590), .Z(n6746)
         );
  OR2_X1 U8212 ( .A1(n6747), .A2(n6746), .ZN(n6591) );
  NAND2_X1 U8213 ( .A1(n6592), .A2(n6591), .ZN(n6707) );
  NOR2_X1 U8214 ( .A1(n6708), .A2(n6707), .ZN(n6706) );
  NOR2_X1 U8215 ( .A1(n6593), .A2(n6706), .ZN(n6728) );
  MUX2_X1 U8216 ( .A(n6594), .B(P1_REG1_REG_7__SCAN_IN), .S(n6732), .Z(n6727)
         );
  NOR2_X1 U8217 ( .A1(n6728), .A2(n6727), .ZN(n6726) );
  AOI21_X1 U8218 ( .B1(n6594), .B2(n6669), .A(n6726), .ZN(n6757) );
  AOI22_X1 U8219 ( .A1(P1_REG1_REG_8__SCAN_IN), .A2(n6760), .B1(n6595), .B2(
        n6596), .ZN(n6756) );
  NOR2_X1 U8220 ( .A1(n6757), .A2(n6756), .ZN(n6755) );
  AOI21_X1 U8221 ( .B1(n6596), .B2(n6760), .A(n6755), .ZN(n9620) );
  INV_X1 U8222 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n9726) );
  AOI22_X1 U8223 ( .A1(n9624), .A2(n9726), .B1(P1_REG1_REG_9__SCAN_IN), .B2(
        n6681), .ZN(n9619) );
  NOR2_X1 U8224 ( .A1(n9620), .A2(n9619), .ZN(n9618) );
  NOR2_X1 U8225 ( .A1(n6597), .A2(n9618), .ZN(n9633) );
  INV_X1 U8226 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6598) );
  MUX2_X1 U8227 ( .A(n6598), .B(P1_REG1_REG_10__SCAN_IN), .S(n9630), .Z(n9632)
         );
  NOR2_X1 U8228 ( .A1(n9633), .A2(n9632), .ZN(n9631) );
  INV_X1 U8229 ( .A(n9631), .ZN(n6599) );
  NAND2_X1 U8230 ( .A1(n6600), .A2(n6599), .ZN(n9644) );
  OAI21_X1 U8231 ( .B1(n9654), .B2(n6601), .A(n9644), .ZN(n6602) );
  NAND2_X1 U8232 ( .A1(n9654), .A2(n6601), .ZN(n9652) );
  NAND2_X1 U8233 ( .A1(n6602), .A2(n9652), .ZN(n9651) );
  NOR2_X1 U8234 ( .A1(n6604), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n6603) );
  AOI21_X1 U8235 ( .B1(P1_REG1_REG_12__SCAN_IN), .B2(n6604), .A(n6603), .ZN(
        n6919) );
  NAND2_X1 U8236 ( .A1(n9651), .A2(n6919), .ZN(n6918) );
  OAI21_X1 U8237 ( .B1(n6604), .B2(P1_REG1_REG_12__SCAN_IN), .A(n6918), .ZN(
        n6848) );
  NAND2_X1 U8238 ( .A1(n6849), .A2(n6848), .ZN(n6847) );
  OAI21_X1 U8239 ( .B1(n6855), .B2(P1_REG1_REG_13__SCAN_IN), .A(n6847), .ZN(
        n9670) );
  NAND2_X1 U8240 ( .A1(n9669), .A2(n9670), .ZN(n9668) );
  OAI21_X1 U8241 ( .B1(n9663), .B2(P1_REG1_REG_14__SCAN_IN), .A(n9668), .ZN(
        n7421) );
  XNOR2_X1 U8242 ( .A(n7422), .B(n7421), .ZN(n6608) );
  INV_X1 U8243 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9573) );
  NOR2_X1 U8244 ( .A1(n9573), .A2(n6608), .ZN(n7423) );
  AND2_X1 U8245 ( .A1(n5801), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6605) );
  NAND2_X1 U8246 ( .A1(n6606), .A2(n6605), .ZN(n9604) );
  INV_X1 U8247 ( .A(n9604), .ZN(n6607) );
  NAND2_X1 U8248 ( .A1(n6607), .A2(n7983), .ZN(n9634) );
  AOI211_X1 U8249 ( .C1(n6608), .C2(n9573), .A(n7423), .B(n9634), .ZN(n6610)
         );
  NAND2_X1 U8250 ( .A1(n9643), .A2(n6249), .ZN(n9646) );
  NAND2_X1 U8251 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9102) );
  OAI21_X1 U8252 ( .B1(n9646), .B2(n7422), .A(n9102), .ZN(n6609) );
  OR4_X1 U8253 ( .A1(n6612), .A2(n6611), .A3(n6610), .A4(n6609), .ZN(P1_U3256)
         );
  XNOR2_X1 U8254 ( .A(n6613), .B(n6627), .ZN(n6635) );
  NAND2_X1 U8255 ( .A1(n6614), .A2(n9282), .ZN(n6617) );
  NAND2_X1 U8256 ( .A1(n6615), .A2(n6775), .ZN(n6616) );
  NAND2_X1 U8257 ( .A1(n6617), .A2(n6616), .ZN(n9406) );
  NAND2_X1 U8258 ( .A1(n6930), .A2(n6934), .ZN(n6929) );
  NAND2_X1 U8259 ( .A1(n6309), .A2(n6933), .ZN(n6620) );
  NAND2_X1 U8260 ( .A1(n6929), .A2(n6620), .ZN(n7114) );
  NAND2_X1 U8261 ( .A1(n7114), .A2(n7115), .ZN(n7113) );
  NAND2_X1 U8262 ( .A1(n7134), .A2(n9706), .ZN(n6621) );
  NAND2_X1 U8263 ( .A1(n7113), .A2(n6621), .ZN(n7133) );
  NAND2_X1 U8264 ( .A1(n7133), .A2(n7138), .ZN(n7132) );
  NAND2_X1 U8265 ( .A1(n7262), .A2(n7173), .ZN(n6622) );
  NAND2_X1 U8266 ( .A1(n7250), .A2(n6625), .ZN(n7249) );
  NAND2_X1 U8267 ( .A1(n9129), .A2(n9680), .ZN(n6626) );
  NAND2_X1 U8268 ( .A1(n6628), .A2(n6627), .ZN(n6629) );
  NAND2_X1 U8269 ( .A1(n7299), .A2(n6629), .ZN(n7184) );
  AOI21_X1 U8270 ( .B1(n6241), .B2(n6639), .A(n9282), .ZN(n6630) );
  NAND2_X1 U8271 ( .A1(n7305), .A2(n6630), .ZN(n7248) );
  INV_X1 U8272 ( .A(n7248), .ZN(n7625) );
  NAND2_X1 U8273 ( .A1(n7184), .A2(n7625), .ZN(n6634) );
  NAND2_X1 U8274 ( .A1(n6631), .A2(n6249), .ZN(n9333) );
  OAI22_X1 U8275 ( .A1(n7300), .A2(n9333), .B1(n7441), .B2(n9331), .ZN(n6632)
         );
  INV_X1 U8276 ( .A(n6632), .ZN(n6633) );
  OAI211_X1 U8277 ( .C1(n6635), .C2(n9329), .A(n6634), .B(n6633), .ZN(n7185)
         );
  NOR2_X1 U8278 ( .A1(n6767), .A2(n6636), .ZN(n7394) );
  NAND2_X1 U8279 ( .A1(n7394), .A2(n7393), .ZN(n6637) );
  MUX2_X1 U8280 ( .A(n7185), .B(P1_REG2_REG_6__SCAN_IN), .S(n6638), .Z(n6649)
         );
  NOR2_X1 U8281 ( .A1(n6639), .A2(n9682), .ZN(n6640) );
  NAND2_X1 U8282 ( .A1(n9321), .A2(n6640), .ZN(n7237) );
  INV_X1 U8283 ( .A(n7237), .ZN(n7632) );
  NAND2_X1 U8284 ( .A1(n7184), .A2(n7632), .ZN(n6647) );
  NAND3_X1 U8285 ( .A1(n6618), .A2(n6933), .A3(n7225), .ZN(n7120) );
  NOR2_X1 U8286 ( .A1(n7120), .A2(n7124), .ZN(n7141) );
  NAND2_X1 U8287 ( .A1(n7141), .A2(n7173), .ZN(n7254) );
  NAND2_X1 U8288 ( .A1(n7255), .A2(n7440), .ZN(n6641) );
  AND2_X1 U8289 ( .A1(n7390), .A2(n6641), .ZN(n7186) );
  INV_X1 U8290 ( .A(n6642), .ZN(n6643) );
  AND2_X1 U8291 ( .A1(n9688), .A2(n6643), .ZN(n9409) );
  INV_X1 U8292 ( .A(n7444), .ZN(n6644) );
  OAI22_X1 U8293 ( .A1(n9396), .A2(n7296), .B1(n9692), .B2(n6644), .ZN(n6645)
         );
  AOI21_X1 U8294 ( .B1(n7186), .B2(n9409), .A(n6645), .ZN(n6646) );
  NAND2_X1 U8295 ( .A1(n6647), .A2(n6646), .ZN(n6648) );
  OR2_X1 U8296 ( .A1(n6649), .A2(n6648), .ZN(P1_U3285) );
  XNOR2_X1 U8297 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  AOI22_X1 U8298 ( .A1(n8969), .A2(P1_DATAO_REG_3__SCAN_IN), .B1(n8385), .B2(
        P2_STATE_REG_SCAN_IN), .ZN(n6650) );
  OAI21_X1 U8299 ( .B1(n6654), .B2(n8967), .A(n6650), .ZN(P2_U3355) );
  AOI22_X1 U8300 ( .A1(n8399), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_4__SCAN_IN), .B2(n8969), .ZN(n6651) );
  OAI21_X1 U8301 ( .B1(n6662), .B2(n8967), .A(n6651), .ZN(P2_U3354) );
  AOI22_X1 U8302 ( .A1(n8413), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(n8969), .ZN(n6652) );
  OAI21_X1 U8303 ( .B1(n6653), .B2(n8967), .A(n6652), .ZN(P2_U3353) );
  OAI222_X1 U8304 ( .A1(n6744), .A2(P1_U3084), .B1(n9508), .B2(n6653), .C1(
        n9957), .C2(n9510), .ZN(P1_U3348) );
  INV_X1 U8305 ( .A(n9150), .ZN(n9148) );
  OAI222_X1 U8306 ( .A1(n9510), .A2(n6655), .B1(n9508), .B2(n6654), .C1(n9148), 
        .C2(P1_U3084), .ZN(P1_U3350) );
  OAI222_X1 U8307 ( .A1(n6710), .A2(P1_U3084), .B1(n9508), .B2(n6657), .C1(
        n10041), .C2(n9510), .ZN(P1_U3347) );
  INV_X1 U8308 ( .A(n8969), .ZN(n7990) );
  OAI222_X1 U8309 ( .A1(n7990), .A2(n6658), .B1(n8967), .B2(n6657), .C1(
        P2_U3152), .C2(n6656), .ZN(P2_U3352) );
  OAI222_X1 U8310 ( .A1(P2_U3152), .A2(n4947), .B1(n8967), .B2(n6665), .C1(
        n4752), .C2(n7990), .ZN(P2_U3357) );
  INV_X1 U8311 ( .A(n9533), .ZN(n6892) );
  OAI222_X1 U8312 ( .A1(P2_U3152), .A2(n6892), .B1(n8967), .B2(n6671), .C1(
        n6659), .C2(n7990), .ZN(P2_U3356) );
  INV_X1 U8313 ( .A(n8441), .ZN(n6898) );
  OAI222_X1 U8314 ( .A1(n7990), .A2(n6660), .B1(n8967), .B2(n6668), .C1(
        P2_U3152), .C2(n6898), .ZN(P2_U3351) );
  INV_X1 U8315 ( .A(n6808), .ZN(n6661) );
  OAI222_X1 U8316 ( .A1(n9510), .A2(n6663), .B1(n9508), .B2(n6662), .C1(n6661), 
        .C2(P1_U3084), .ZN(P1_U3349) );
  INV_X1 U8317 ( .A(n6664), .ZN(n9136) );
  OAI222_X1 U8318 ( .A1(n9510), .A2(n6666), .B1(n9508), .B2(n6665), .C1(n9136), 
        .C2(P1_U3084), .ZN(P1_U3352) );
  OAI222_X1 U8319 ( .A1(n6669), .A2(P1_U3084), .B1(n9508), .B2(n6668), .C1(
        n6667), .C2(n9510), .ZN(P1_U3346) );
  INV_X1 U8320 ( .A(n6670), .ZN(n9608) );
  OAI222_X1 U8321 ( .A1(n9510), .A2(n6672), .B1(n9508), .B2(n6671), .C1(n9608), 
        .C2(P1_U3084), .ZN(P1_U3351) );
  INV_X1 U8322 ( .A(n6673), .ZN(n6675) );
  OAI222_X1 U8323 ( .A1(n6760), .A2(P1_U3084), .B1(n9508), .B2(n6675), .C1(
        n6674), .C2(n9510), .ZN(P1_U3345) );
  INV_X1 U8324 ( .A(n8455), .ZN(n6899) );
  OAI222_X1 U8325 ( .A1(n7990), .A2(n6676), .B1(n8967), .B2(n6675), .C1(
        P2_U3152), .C2(n6899), .ZN(P2_U3350) );
  INV_X1 U8326 ( .A(n6677), .ZN(n6680) );
  AOI22_X1 U8327 ( .A1(n8469), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n8969), .ZN(n6678) );
  OAI21_X1 U8328 ( .B1(n6680), .B2(n8967), .A(n6678), .ZN(P2_U3349) );
  OAI222_X1 U8329 ( .A1(P1_U3084), .A2(n6681), .B1(n9508), .B2(n6680), .C1(
        n6679), .C2(n9510), .ZN(P1_U3344) );
  INV_X1 U8330 ( .A(n6682), .ZN(n6684) );
  INV_X1 U8331 ( .A(n9510), .ZN(n9506) );
  AOI22_X1 U8332 ( .A1(n9630), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n9506), .ZN(n6683) );
  OAI21_X1 U8333 ( .B1(n6684), .B2(n9508), .A(n6683), .ZN(P1_U3343) );
  INV_X1 U8334 ( .A(n7016), .ZN(n6909) );
  OAI222_X1 U8335 ( .A1(n7990), .A2(n6685), .B1(n8967), .B2(n6684), .C1(n6909), 
        .C2(P2_U3152), .ZN(P2_U3348) );
  INV_X1 U8336 ( .A(n6686), .ZN(n6688) );
  INV_X1 U8337 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6687) );
  OAI222_X1 U8338 ( .A1(P1_U3084), .A2(n9654), .B1(n9508), .B2(n6688), .C1(
        n6687), .C2(n9510), .ZN(P1_U3342) );
  INV_X1 U8339 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6689) );
  INV_X1 U8340 ( .A(n7162), .ZN(n7154) );
  OAI222_X1 U8341 ( .A1(n7990), .A2(n6689), .B1(n8967), .B2(n6688), .C1(n7154), 
        .C2(P2_U3152), .ZN(P2_U3347) );
  NAND2_X1 U8342 ( .A1(n9697), .A2(n6772), .ZN(n9694) );
  INV_X1 U8343 ( .A(n9694), .ZN(n9693) );
  OAI21_X1 U8344 ( .B1(n9693), .B2(P1_D_REG_1__SCAN_IN), .A(n6771), .ZN(n6690)
         );
  OAI21_X1 U8345 ( .B1(n9697), .B2(n6691), .A(n6690), .ZN(P1_U3441) );
  INV_X1 U8346 ( .A(n6692), .ZN(n6699) );
  AOI22_X1 U8347 ( .A1(n8483), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_12__SCAN_IN), .B2(n8969), .ZN(n6693) );
  OAI21_X1 U8348 ( .B1(n6699), .B2(n8967), .A(n6693), .ZN(P2_U3346) );
  NAND2_X1 U8349 ( .A1(n9762), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8368) );
  NAND2_X1 U8350 ( .A1(n9759), .A2(n8368), .ZN(n6695) );
  NAND2_X1 U8351 ( .A1(n6695), .A2(n6694), .ZN(n6698) );
  OR2_X1 U8352 ( .A1(n9759), .A2(n6696), .ZN(n6697) );
  NAND2_X1 U8353 ( .A1(n6698), .A2(n6697), .ZN(n9734) );
  NOR2_X1 U8354 ( .A1(n9734), .A2(P2_U3966), .ZN(P2_U3151) );
  OAI222_X1 U8355 ( .A1(n9510), .A2(n6700), .B1(n9508), .B2(n6699), .C1(n6923), 
        .C2(P1_U3084), .ZN(P1_U3341) );
  INV_X1 U8356 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n6705) );
  NAND2_X1 U8357 ( .A1(n8036), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n6703) );
  NAND2_X1 U8358 ( .A1(n8035), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n6702) );
  NAND2_X1 U8359 ( .A1(n8037), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n6701) );
  AND3_X1 U8360 ( .A1(n6703), .A2(n6702), .A3(n6701), .ZN(n8347) );
  INV_X1 U8361 ( .A(n8347), .ZN(n8573) );
  NAND2_X1 U8362 ( .A1(P2_U3966), .A2(n8573), .ZN(n6704) );
  OAI21_X1 U8363 ( .B1(P2_U3966), .B2(n6705), .A(n6704), .ZN(P2_U3583) );
  AOI21_X1 U8364 ( .B1(n6708), .B2(n6707), .A(n6706), .ZN(n6717) );
  INV_X1 U8365 ( .A(n9678), .ZN(n9648) );
  NOR2_X1 U8366 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6709), .ZN(n7443) );
  NOR2_X1 U8367 ( .A1(n9646), .A2(n6710), .ZN(n6711) );
  AOI211_X1 U8368 ( .C1(n9648), .C2(P1_ADDR_REG_6__SCAN_IN), .A(n7443), .B(
        n6711), .ZN(n6716) );
  OAI211_X1 U8369 ( .C1(n6714), .C2(n6713), .A(n9673), .B(n6712), .ZN(n6715)
         );
  OAI211_X1 U8370 ( .C1(n6717), .C2(n9634), .A(n6716), .B(n6715), .ZN(P1_U3247) );
  INV_X1 U8371 ( .A(n6718), .ZN(n6721) );
  OAI222_X1 U8372 ( .A1(n9510), .A2(n6720), .B1(n9508), .B2(n6721), .C1(
        P1_U3084), .C2(n6719), .ZN(P1_U3340) );
  INV_X1 U8373 ( .A(n7318), .ZN(n7159) );
  OAI222_X1 U8374 ( .A1(n7990), .A2(n6722), .B1(n8967), .B2(n6721), .C1(n7159), 
        .C2(P2_U3152), .ZN(P2_U3345) );
  INV_X1 U8375 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n6735) );
  AOI21_X1 U8376 ( .B1(n6725), .B2(n6724), .A(n6723), .ZN(n6730) );
  AOI21_X1 U8377 ( .B1(n6728), .B2(n6727), .A(n6726), .ZN(n6729) );
  OAI22_X1 U8378 ( .A1(n6730), .A2(n9182), .B1(n9634), .B2(n6729), .ZN(n6731)
         );
  INV_X1 U8379 ( .A(n6731), .ZN(n6734) );
  INV_X1 U8380 ( .A(n9646), .ZN(n9664) );
  AND2_X1 U8381 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7476) );
  AOI21_X1 U8382 ( .B1(n9664), .B2(n6732), .A(n7476), .ZN(n6733) );
  OAI211_X1 U8383 ( .C1(n9678), .C2(n6735), .A(n6734), .B(n6733), .ZN(P1_U3248) );
  INV_X1 U8384 ( .A(n6736), .ZN(n6739) );
  INV_X1 U8385 ( .A(n8493), .ZN(n8498) );
  OAI222_X1 U8386 ( .A1(n7990), .A2(n6737), .B1(n8967), .B2(n6739), .C1(n8498), 
        .C2(P2_U3152), .ZN(P2_U3344) );
  OAI222_X1 U8387 ( .A1(P1_U3084), .A2(n6740), .B1(n9508), .B2(n6739), .C1(
        n6738), .C2(n9510), .ZN(P1_U3339) );
  AOI21_X1 U8388 ( .B1(n6743), .B2(n6742), .A(n6741), .ZN(n6751) );
  AND2_X1 U8389 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n7264) );
  NOR2_X1 U8390 ( .A1(n9646), .A2(n6744), .ZN(n6745) );
  AOI211_X1 U8391 ( .C1(n9648), .C2(P1_ADDR_REG_5__SCAN_IN), .A(n7264), .B(
        n6745), .ZN(n6750) );
  INV_X1 U8392 ( .A(n9634), .ZN(n9672) );
  XOR2_X1 U8393 ( .A(n6747), .B(n6746), .Z(n6748) );
  NAND2_X1 U8394 ( .A1(n9672), .A2(n6748), .ZN(n6749) );
  OAI211_X1 U8395 ( .C1(n6751), .C2(n9182), .A(n6750), .B(n6749), .ZN(P1_U3246) );
  AOI21_X1 U8396 ( .B1(n6754), .B2(n6753), .A(n6752), .ZN(n6765) );
  AOI21_X1 U8397 ( .B1(n6757), .B2(n6756), .A(n6755), .ZN(n6758) );
  NOR2_X1 U8398 ( .A1(n6758), .A2(n9634), .ZN(n6763) );
  NOR2_X1 U8399 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6759), .ZN(n7537) );
  INV_X1 U8400 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n7567) );
  NOR2_X1 U8401 ( .A1(n9678), .A2(n7567), .ZN(n6762) );
  NOR2_X1 U8402 ( .A1(n9646), .A2(n6760), .ZN(n6761) );
  NOR4_X1 U8403 ( .A1(n6763), .A2(n7537), .A3(n6762), .A4(n6761), .ZN(n6764)
         );
  OAI21_X1 U8404 ( .B1(n6765), .B2(n9182), .A(n6764), .ZN(P1_U3249) );
  OR2_X1 U8405 ( .A1(n6767), .A2(n6766), .ZN(n9695) );
  NOR2_X1 U8406 ( .A1(n9695), .A2(n6768), .ZN(n6777) );
  INV_X1 U8407 ( .A(n6772), .ZN(n6770) );
  NAND2_X1 U8408 ( .A1(n6770), .A2(n6769), .ZN(n6774) );
  OAI21_X1 U8409 ( .B1(n6772), .B2(P1_D_REG_1__SCAN_IN), .A(n6771), .ZN(n6773)
         );
  OAI211_X1 U8410 ( .C1(n7247), .C2(n6775), .A(n6774), .B(n6773), .ZN(n6776)
         );
  INV_X1 U8411 ( .A(n6776), .ZN(n6953) );
  AND2_X2 U8412 ( .A1(n6777), .A2(n6953), .ZN(n9486) );
  INV_X1 U8413 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n6783) );
  INV_X1 U8414 ( .A(n6932), .ZN(n6781) );
  INV_X1 U8415 ( .A(n7305), .ZN(n6778) );
  AOI211_X1 U8416 ( .C1(n6779), .C2(n7227), .A(n6778), .B(n6932), .ZN(n6780)
         );
  AOI21_X1 U8417 ( .B1(n9403), .B2(n9133), .A(n6780), .ZN(n7106) );
  OAI21_X1 U8418 ( .B1(n7225), .B2(n6781), .A(n7106), .ZN(n6954) );
  NAND2_X1 U8419 ( .A1(n6954), .A2(n9486), .ZN(n6782) );
  OAI21_X1 U8420 ( .B1(n9486), .B2(n6783), .A(n6782), .ZN(P1_U3523) );
  INV_X1 U8421 ( .A(n6784), .ZN(n6793) );
  NAND2_X1 U8422 ( .A1(n6793), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6787) );
  NAND2_X1 U8423 ( .A1(n6789), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6785) );
  OR2_X1 U8424 ( .A1(n9634), .A2(n6785), .ZN(n6786) );
  OAI211_X1 U8425 ( .C1(n9182), .C2(n6787), .A(n6786), .B(n9646), .ZN(n6807)
         );
  NAND2_X1 U8426 ( .A1(n6789), .A2(n6788), .ZN(n6790) );
  AND2_X1 U8427 ( .A1(n6791), .A2(n6790), .ZN(n6799) );
  NAND2_X1 U8428 ( .A1(n6793), .A2(n6792), .ZN(n6794) );
  NAND2_X1 U8429 ( .A1(n6795), .A2(n6794), .ZN(n6796) );
  AND2_X1 U8430 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n7084) );
  AOI21_X1 U8431 ( .B1(n9673), .B2(n6796), .A(n7084), .ZN(n6798) );
  NAND2_X1 U8432 ( .A1(n9648), .A2(P1_ADDR_REG_4__SCAN_IN), .ZN(n6797) );
  OAI211_X1 U8433 ( .C1(n6799), .C2(n9634), .A(n6798), .B(n6797), .ZN(n6806)
         );
  OAI21_X1 U8434 ( .B1(n6802), .B2(n6800), .A(n6801), .ZN(n6942) );
  INV_X1 U8435 ( .A(n7983), .ZN(n9597) );
  OAI21_X1 U8436 ( .B1(P1_REG2_REG_0__SCAN_IN), .B2(n7983), .A(n6803), .ZN(
        n9598) );
  NOR3_X1 U8437 ( .A1(n6942), .A2(n9597), .A3(n9598), .ZN(n6805) );
  INV_X2 U8438 ( .A(P1_U4006), .ZN(n9134) );
  NOR2_X1 U8439 ( .A1(n9598), .A2(n7983), .ZN(n6804) );
  MUX2_X1 U8440 ( .A(n9598), .B(n6804), .S(P1_IR_REG_0__SCAN_IN), .Z(n9602) );
  NOR3_X1 U8441 ( .A1(n6805), .A2(n9134), .A3(n9602), .ZN(n9610) );
  AOI211_X1 U8442 ( .C1(n6808), .C2(n6807), .A(n6806), .B(n9610), .ZN(n6809)
         );
  INV_X1 U8443 ( .A(n6809), .ZN(P1_U3245) );
  INV_X1 U8444 ( .A(n6810), .ZN(n6813) );
  NOR2_X1 U8445 ( .A1(n9759), .A2(n6811), .ZN(n6812) );
  NAND2_X1 U8446 ( .A1(n6813), .A2(n6812), .ZN(n7036) );
  INV_X1 U8447 ( .A(n6814), .ZN(n6815) );
  OR2_X1 U8448 ( .A1(n7037), .A2(n6815), .ZN(n6816) );
  AND2_X2 U8449 ( .A1(n7274), .A2(n7272), .ZN(n9833) );
  INV_X1 U8450 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n6827) );
  INV_X1 U8451 ( .A(n6817), .ZN(n7025) );
  NAND2_X1 U8452 ( .A1(n6818), .A2(n6819), .ZN(n7028) );
  OAI21_X1 U8453 ( .B1(n6818), .B2(n6819), .A(n7028), .ZN(n8828) );
  INV_X1 U8454 ( .A(n8828), .ZN(n6825) );
  XNOR2_X1 U8455 ( .A(n6820), .B(n7040), .ZN(n6821) );
  OR2_X1 U8456 ( .A1(n6821), .A2(n8356), .ZN(n8780) );
  NAND3_X1 U8457 ( .A1(n8343), .A2(n6820), .A3(n8356), .ZN(n9809) );
  XNOR2_X1 U8458 ( .A(n7092), .B(n6818), .ZN(n6823) );
  NAND2_X1 U8459 ( .A1(n8346), .A2(n8199), .ZN(n8358) );
  INV_X2 U8460 ( .A(n8751), .ZN(n8813) );
  OAI22_X1 U8461 ( .A1(n6822), .A2(n8756), .B1(n7030), .B2(n8754), .ZN(n7004)
         );
  AOI21_X1 U8462 ( .B1(n6823), .B2(n8813), .A(n7004), .ZN(n8831) );
  AOI21_X1 U8463 ( .B1(n9770), .B2(n8826), .A(n7352), .ZN(n8829) );
  INV_X1 U8464 ( .A(n9825), .ZN(n9803) );
  AOI22_X1 U8465 ( .A1(n8829), .A2(n9803), .B1(n9802), .B2(n8826), .ZN(n6824)
         );
  OAI211_X1 U8466 ( .C1(n6825), .C2(n9797), .A(n8831), .B(n6824), .ZN(n8939)
         );
  NAND2_X1 U8467 ( .A1(n9833), .A2(n8939), .ZN(n6826) );
  OAI21_X1 U8468 ( .B1(n9833), .B2(n6827), .A(n6826), .ZN(P2_U3454) );
  INV_X1 U8469 ( .A(n6828), .ZN(n6831) );
  INV_X1 U8470 ( .A(n8513), .ZN(n8507) );
  OAI222_X1 U8471 ( .A1(n7990), .A2(n6829), .B1(n8967), .B2(n6831), .C1(
        P2_U3152), .C2(n8507), .ZN(P2_U3343) );
  OAI222_X1 U8472 ( .A1(n7422), .A2(P1_U3084), .B1(n9508), .B2(n6831), .C1(
        n6830), .C2(n9510), .ZN(P1_U3338) );
  XNOR2_X1 U8473 ( .A(n6833), .B(n6832), .ZN(n6835) );
  INV_X1 U8474 ( .A(n6837), .ZN(n6834) );
  NAND2_X1 U8475 ( .A1(n6835), .A2(n6834), .ZN(n6839) );
  INV_X1 U8476 ( .A(n6836), .ZN(n6838) );
  AOI22_X1 U8477 ( .A1(n6840), .A2(n6839), .B1(n6838), .B2(n6837), .ZN(n6846)
         );
  AOI22_X1 U8478 ( .A1(n9094), .A2(n9132), .B1(n9104), .B2(n6306), .ZN(n6845)
         );
  NAND4_X1 U8479 ( .A1(n6843), .A2(n6842), .A3(n9697), .A4(n6841), .ZN(n6949)
         );
  AOI22_X1 U8480 ( .A1(n9112), .A2(n7234), .B1(P1_REG3_REG_1__SCAN_IN), .B2(
        n6949), .ZN(n6844) );
  OAI211_X1 U8481 ( .C1(n6846), .C2(n9115), .A(n6845), .B(n6844), .ZN(P1_U3220) );
  INV_X1 U8482 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n6858) );
  OAI21_X1 U8483 ( .B1(n6849), .B2(n6848), .A(n6847), .ZN(n6854) );
  AOI211_X1 U8484 ( .C1(n6852), .C2(n6851), .A(n6850), .B(n9182), .ZN(n6853)
         );
  AOI21_X1 U8485 ( .B1(n9672), .B2(n6854), .A(n6853), .ZN(n6857) );
  AND2_X1 U8486 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n7862) );
  AOI21_X1 U8487 ( .B1(n9664), .B2(n6855), .A(n7862), .ZN(n6856) );
  OAI211_X1 U8488 ( .C1(n9678), .C2(n6858), .A(n6857), .B(n6856), .ZN(P1_U3254) );
  OAI211_X1 U8489 ( .C1(n9759), .C2(n6860), .A(n8368), .B(n6859), .ZN(n6877)
         );
  NAND2_X1 U8490 ( .A1(n6877), .A2(n6875), .ZN(n6861) );
  NAND2_X1 U8491 ( .A1(n6861), .A2(n8370), .ZN(n6904) );
  NAND2_X1 U8492 ( .A1(n6904), .A2(n5620), .ZN(n9730) );
  NAND2_X1 U8493 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3152), .ZN(n7345) );
  INV_X1 U8494 ( .A(n7345), .ZN(n6880) );
  INV_X1 U8495 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n9737) );
  INV_X1 U8496 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n9834) );
  NOR3_X1 U8497 ( .A1(n9737), .A2(n9834), .A3(n9516), .ZN(n9514) );
  NOR2_X1 U8498 ( .A1(n9514), .A2(n6862), .ZN(n9531) );
  NAND2_X1 U8499 ( .A1(n9533), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6863) );
  OAI21_X1 U8500 ( .B1(n9533), .B2(P2_REG1_REG_2__SCAN_IN), .A(n6863), .ZN(
        n9530) );
  NOR2_X1 U8501 ( .A1(n9531), .A2(n9530), .ZN(n9529) );
  AOI21_X1 U8502 ( .B1(n9533), .B2(P2_REG1_REG_2__SCAN_IN), .A(n9529), .ZN(
        n8388) );
  OR2_X1 U8503 ( .A1(n8385), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6865) );
  NAND2_X1 U8504 ( .A1(n8385), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6864) );
  NAND2_X1 U8505 ( .A1(n6865), .A2(n6864), .ZN(n8387) );
  OR2_X1 U8506 ( .A1(n8399), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6867) );
  NAND2_X1 U8507 ( .A1(n8399), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6866) );
  NAND2_X1 U8508 ( .A1(n6867), .A2(n6866), .ZN(n8402) );
  NAND2_X1 U8509 ( .A1(n8413), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6868) );
  OAI21_X1 U8510 ( .B1(n8413), .B2(P2_REG1_REG_5__SCAN_IN), .A(n6868), .ZN(
        n8416) );
  NOR2_X1 U8511 ( .A1(n8415), .A2(n8416), .ZN(n8414) );
  OR2_X1 U8512 ( .A1(n8427), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6870) );
  NAND2_X1 U8513 ( .A1(n8427), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6869) );
  NAND2_X1 U8514 ( .A1(n6870), .A2(n6869), .ZN(n8430) );
  INV_X1 U8515 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6871) );
  MUX2_X1 U8516 ( .A(n6871), .B(P2_REG1_REG_7__SCAN_IN), .S(n8441), .Z(n8444)
         );
  AOI21_X1 U8517 ( .B1(n8441), .B2(P2_REG1_REG_7__SCAN_IN), .A(n8442), .ZN(
        n8457) );
  INV_X1 U8518 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6872) );
  MUX2_X1 U8519 ( .A(n6872), .B(P2_REG1_REG_8__SCAN_IN), .S(n8455), .Z(n8458)
         );
  INV_X1 U8520 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6873) );
  MUX2_X1 U8521 ( .A(n6873), .B(P2_REG1_REG_9__SCAN_IN), .S(n8469), .Z(n8472)
         );
  INV_X1 U8522 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n6874) );
  MUX2_X1 U8523 ( .A(n6874), .B(P2_REG1_REG_10__SCAN_IN), .S(n7016), .Z(n6878)
         );
  NOR2_X1 U8524 ( .A1(n4343), .A2(n6878), .ZN(n7015) );
  AND2_X1 U8525 ( .A1(n6875), .A2(n8364), .ZN(n6876) );
  INV_X1 U8526 ( .A(n9729), .ZN(n9528) );
  AOI211_X1 U8527 ( .C1(n4343), .C2(n6878), .A(n7015), .B(n9528), .ZN(n6879)
         );
  AOI211_X1 U8528 ( .C1(P2_ADDR_REG_10__SCAN_IN), .C2(n9734), .A(n6880), .B(
        n6879), .ZN(n6908) );
  NAND2_X1 U8529 ( .A1(n8469), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6900) );
  INV_X1 U8530 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n6881) );
  MUX2_X1 U8531 ( .A(n6881), .B(P2_REG2_REG_9__SCAN_IN), .S(n8469), .Z(n6882)
         );
  INV_X1 U8532 ( .A(n6882), .ZN(n8466) );
  INV_X1 U8533 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n9878) );
  MUX2_X1 U8534 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n9878), .S(n8455), .Z(n8451)
         );
  INV_X1 U8535 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6897) );
  MUX2_X1 U8536 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n6897), .S(n8441), .Z(n8437)
         );
  NAND2_X1 U8537 ( .A1(n8427), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6896) );
  INV_X1 U8538 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6883) );
  MUX2_X1 U8539 ( .A(n6883), .B(P2_REG2_REG_6__SCAN_IN), .S(n8427), .Z(n6884)
         );
  INV_X1 U8540 ( .A(n6884), .ZN(n8423) );
  NAND2_X1 U8541 ( .A1(n8413), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6895) );
  INV_X1 U8542 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6885) );
  MUX2_X1 U8543 ( .A(n6885), .B(P2_REG2_REG_5__SCAN_IN), .S(n8413), .Z(n6886)
         );
  INV_X1 U8544 ( .A(n6886), .ZN(n8409) );
  NAND2_X1 U8545 ( .A1(n8399), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6894) );
  INV_X1 U8546 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6887) );
  MUX2_X1 U8547 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n6887), .S(n8399), .Z(n8395)
         );
  NAND2_X1 U8548 ( .A1(n8385), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6893) );
  INV_X1 U8549 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6888) );
  MUX2_X1 U8550 ( .A(n6888), .B(P2_REG2_REG_3__SCAN_IN), .S(n8385), .Z(n6889)
         );
  INV_X1 U8551 ( .A(n6889), .ZN(n8383) );
  INV_X1 U8552 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6891) );
  XNOR2_X1 U8553 ( .A(n6892), .B(P2_REG2_REG_2__SCAN_IN), .ZN(n9537) );
  INV_X1 U8554 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6890) );
  NAND3_X1 U8555 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .A3(n9522), .ZN(n9521) );
  OAI21_X1 U8556 ( .B1(n4947), .B2(n6890), .A(n9521), .ZN(n9536) );
  NAND2_X1 U8557 ( .A1(n9537), .A2(n9536), .ZN(n9535) );
  OAI21_X1 U8558 ( .B1(n6892), .B2(n6891), .A(n9535), .ZN(n8382) );
  NAND2_X1 U8559 ( .A1(n8383), .A2(n8382), .ZN(n8381) );
  NAND2_X1 U8560 ( .A1(n6893), .A2(n8381), .ZN(n8396) );
  NAND2_X1 U8561 ( .A1(n8395), .A2(n8396), .ZN(n8394) );
  NAND2_X1 U8562 ( .A1(n6894), .A2(n8394), .ZN(n8410) );
  NAND2_X1 U8563 ( .A1(n8409), .A2(n8410), .ZN(n8408) );
  NAND2_X1 U8564 ( .A1(n6895), .A2(n8408), .ZN(n8424) );
  NAND2_X1 U8565 ( .A1(n8423), .A2(n8424), .ZN(n8422) );
  NAND2_X1 U8566 ( .A1(n6896), .A2(n8422), .ZN(n8438) );
  NAND2_X1 U8567 ( .A1(n8437), .A2(n8438), .ZN(n8436) );
  OAI21_X1 U8568 ( .B1(n6898), .B2(n6897), .A(n8436), .ZN(n8452) );
  NAND2_X1 U8569 ( .A1(n8451), .A2(n8452), .ZN(n8450) );
  OAI21_X1 U8570 ( .B1(n6899), .B2(n9878), .A(n8450), .ZN(n8465) );
  NAND2_X1 U8571 ( .A1(n8466), .A2(n8465), .ZN(n8464) );
  NAND2_X1 U8572 ( .A1(n6900), .A2(n8464), .ZN(n6906) );
  INV_X1 U8573 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n6901) );
  MUX2_X1 U8574 ( .A(n6901), .B(P2_REG2_REG_10__SCAN_IN), .S(n7016), .Z(n6902)
         );
  INV_X1 U8575 ( .A(n6902), .ZN(n6905) );
  NOR2_X1 U8576 ( .A1(n5620), .A2(n8364), .ZN(n6903) );
  NAND2_X1 U8577 ( .A1(n6904), .A2(n6903), .ZN(n9732) );
  NAND2_X1 U8578 ( .A1(n6905), .A2(n6906), .ZN(n7010) );
  OAI211_X1 U8579 ( .C1(n6906), .C2(n6905), .A(n9728), .B(n7010), .ZN(n6907)
         );
  OAI211_X1 U8580 ( .C1(n9730), .C2(n6909), .A(n6908), .B(n6907), .ZN(P2_U3255) );
  AND2_X1 U8581 ( .A1(n6910), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7072) );
  INV_X1 U8582 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n6917) );
  AOI22_X1 U8583 ( .A1(n8124), .A2(n6817), .B1(n8143), .B2(n8379), .ZN(n6916)
         );
  OAI21_X1 U8584 ( .B1(n6913), .B2(n6912), .A(n6911), .ZN(n6914) );
  AOI22_X1 U8585 ( .A1(n4315), .A2(n6914), .B1(n7355), .B2(n8166), .ZN(n6915)
         );
  OAI211_X1 U8586 ( .C1(n7072), .C2(n6917), .A(n6916), .B(n6915), .ZN(P2_U3239) );
  OAI21_X1 U8587 ( .B1(n9651), .B2(n6919), .A(n6918), .ZN(n6920) );
  NAND2_X1 U8588 ( .A1(n9672), .A2(n6920), .ZN(n6922) );
  NAND2_X1 U8589 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3084), .ZN(n6921) );
  OAI211_X1 U8590 ( .C1(n9646), .C2(n6923), .A(n6922), .B(n6921), .ZN(n6927)
         );
  AOI211_X1 U8591 ( .C1(n9655), .C2(n6925), .A(n6924), .B(n9182), .ZN(n6926)
         );
  AOI211_X1 U8592 ( .C1(n9648), .C2(P1_ADDR_REG_12__SCAN_IN), .A(n6927), .B(
        n6926), .ZN(n6928) );
  INV_X1 U8593 ( .A(n6928), .ZN(P1_U3253) );
  OAI21_X1 U8594 ( .B1(n6930), .B2(n6934), .A(n6929), .ZN(n7494) );
  OAI21_X1 U8595 ( .B1(n7234), .B2(n7109), .A(n6308), .ZN(n6931) );
  NAND2_X1 U8596 ( .A1(n7120), .A2(n6931), .ZN(n7490) );
  OAI22_X1 U8597 ( .A1(n7490), .A2(n9707), .B1(n6933), .B2(n9714), .ZN(n6940)
         );
  NAND2_X1 U8598 ( .A1(n7494), .A2(n7625), .ZN(n6939) );
  AOI22_X1 U8599 ( .A1(n9131), .A2(n9403), .B1(n9401), .B2(n9133), .ZN(n6938)
         );
  XNOR2_X1 U8600 ( .A(n6935), .B(n6934), .ZN(n6936) );
  NAND2_X1 U8601 ( .A1(n6936), .A2(n9406), .ZN(n6937) );
  NAND3_X1 U8602 ( .A1(n6939), .A2(n6938), .A3(n6937), .ZN(n7491) );
  AOI211_X1 U8603 ( .C1(n9717), .C2(n7494), .A(n6940), .B(n7491), .ZN(n6971)
         );
  NAND2_X1 U8604 ( .A1(n9725), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6941) );
  OAI21_X1 U8605 ( .B1(n6971), .B2(n9725), .A(n6941), .ZN(P1_U3525) );
  NAND2_X1 U8606 ( .A1(n6942), .A2(n9087), .ZN(n6944) );
  AOI22_X1 U8607 ( .A1(n9094), .A2(n9133), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        n6949), .ZN(n6943) );
  OAI211_X1 U8608 ( .C1(n9097), .C2(n7225), .A(n6944), .B(n6943), .ZN(P1_U3230) );
  INV_X1 U8609 ( .A(n6947), .ZN(n6948) );
  AOI21_X1 U8610 ( .B1(n6945), .B2(n6946), .A(n6948), .ZN(n6952) );
  AOI22_X1 U8611 ( .A1(n9094), .A2(n9131), .B1(n9104), .B2(n9133), .ZN(n6951)
         );
  AOI22_X1 U8612 ( .A1(n9112), .A2(n6308), .B1(P1_REG3_REG_2__SCAN_IN), .B2(
        n6949), .ZN(n6950) );
  OAI211_X1 U8613 ( .C1(n6952), .C2(n9115), .A(n6951), .B(n6950), .ZN(P1_U3235) );
  INV_X2 U8614 ( .A(n9721), .ZN(n9722) );
  NAND2_X1 U8615 ( .A1(n6954), .A2(n9722), .ZN(n6955) );
  OAI21_X1 U8616 ( .B1(n9722), .B2(n5710), .A(n6955), .ZN(P1_U3454) );
  INV_X1 U8617 ( .A(n6956), .ZN(n6983) );
  AOI22_X1 U8618 ( .A1(n9161), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n9506), .ZN(n6957) );
  OAI21_X1 U8619 ( .B1(n6983), .B2(n9508), .A(n6957), .ZN(P1_U3336) );
  INV_X1 U8620 ( .A(n6958), .ZN(n7402) );
  INV_X1 U8621 ( .A(n8378), .ZN(n7212) );
  OAI22_X1 U8622 ( .A1(n7195), .A2(n8756), .B1(n7212), .B2(n8754), .ZN(n7406)
         );
  INV_X1 U8623 ( .A(n7406), .ZN(n6959) );
  OAI22_X1 U8624 ( .A1(n8068), .A2(n6959), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8411), .ZN(n6960) );
  AOI21_X1 U8625 ( .B1(n9794), .B2(n8166), .A(n6960), .ZN(n6966) );
  OAI21_X1 U8626 ( .B1(n6963), .B2(n6962), .A(n6961), .ZN(n6964) );
  NAND2_X1 U8627 ( .A1(n6964), .A2(n4315), .ZN(n6965) );
  OAI211_X1 U8628 ( .C1(n8163), .C2(n7402), .A(n6966), .B(n6965), .ZN(P2_U3229) );
  INV_X1 U8629 ( .A(n6967), .ZN(n6969) );
  OAI222_X1 U8630 ( .A1(n7990), .A2(n6968), .B1(n8967), .B2(n6969), .C1(n8523), 
        .C2(P2_U3152), .ZN(P2_U3342) );
  INV_X1 U8631 ( .A(n7588), .ZN(n7429) );
  OAI222_X1 U8632 ( .A1(n9510), .A2(n6970), .B1(n9508), .B2(n6969), .C1(
        P1_U3084), .C2(n7429), .ZN(P1_U3337) );
  OR2_X1 U8633 ( .A1(n6971), .A2(n9721), .ZN(n6972) );
  OAI21_X1 U8634 ( .B1(n9722), .B2(n6973), .A(n6972), .ZN(P1_U3460) );
  INV_X1 U8635 ( .A(n6975), .ZN(n6976) );
  AOI21_X1 U8636 ( .B1(n6974), .B2(n6977), .A(n6976), .ZN(n6982) );
  INV_X1 U8637 ( .A(n7045), .ZN(n9788) );
  NAND2_X1 U8638 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3152), .ZN(n8397) );
  OAI21_X1 U8639 ( .B1(n8146), .B2(n9788), .A(n8397), .ZN(n6979) );
  INV_X1 U8640 ( .A(n8810), .ZN(n7198) );
  OAI22_X1 U8641 ( .A1(n7359), .A2(n8160), .B1(n8159), .B2(n7198), .ZN(n6978)
         );
  AOI211_X1 U8642 ( .C1(n6980), .C2(n5616), .A(n6979), .B(n6978), .ZN(n6981)
         );
  OAI21_X1 U8643 ( .B1(n6982), .B2(n5614), .A(n6981), .ZN(P2_U3232) );
  INV_X1 U8644 ( .A(n8549), .ZN(n8542) );
  OAI222_X1 U8645 ( .A1(n7990), .A2(n6984), .B1(n8967), .B2(n6983), .C1(n8542), 
        .C2(P2_U3152), .ZN(P2_U3341) );
  NAND2_X1 U8646 ( .A1(n9134), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n6985) );
  OAI21_X1 U8647 ( .B1(n9209), .B2(n9134), .A(n6985), .ZN(P1_U3584) );
  XOR2_X1 U8648 ( .A(n6987), .B(n6986), .Z(n6989) );
  OAI22_X1 U8649 ( .A1(n7030), .A2(n8160), .B1(n8159), .B2(n7195), .ZN(n6988)
         );
  AOI21_X1 U8650 ( .B1(n4315), .B2(n6989), .A(n6988), .ZN(n6991) );
  AOI22_X1 U8651 ( .A1(n8166), .A2(n9749), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        P2_U3152), .ZN(n6990) );
  OAI211_X1 U8652 ( .C1(n8163), .C2(P2_REG3_REG_3__SCAN_IN), .A(n6991), .B(
        n6990), .ZN(P2_U3220) );
  OAI21_X1 U8653 ( .B1(n6994), .B2(n6993), .A(n6992), .ZN(n6998) );
  OAI22_X1 U8654 ( .A1(n7198), .A2(n8160), .B1(n8159), .B2(n7203), .ZN(n6997)
         );
  INV_X1 U8655 ( .A(n9801), .ZN(n8820) );
  NAND2_X1 U8656 ( .A1(n5616), .A2(n8817), .ZN(n6995) );
  NAND2_X1 U8657 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3152), .ZN(n8425) );
  OAI211_X1 U8658 ( .C1(n8820), .C2(n8146), .A(n6995), .B(n8425), .ZN(n6996)
         );
  AOI211_X1 U8659 ( .C1(n4315), .C2(n6998), .A(n6997), .B(n6996), .ZN(n6999)
         );
  INV_X1 U8660 ( .A(n6999), .ZN(P2_U3241) );
  INV_X1 U8661 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7009) );
  INV_X1 U8662 ( .A(n7000), .ZN(n7001) );
  AOI21_X1 U8663 ( .B1(n7003), .B2(n7002), .A(n7001), .ZN(n7006) );
  INV_X1 U8664 ( .A(n7004), .ZN(n7005) );
  OAI22_X1 U8665 ( .A1(n5614), .A2(n7006), .B1(n7005), .B2(n8068), .ZN(n7007)
         );
  AOI21_X1 U8666 ( .B1(n8826), .B2(n8166), .A(n7007), .ZN(n7008) );
  OAI21_X1 U8667 ( .B1(n7072), .B2(n7009), .A(n7008), .ZN(P2_U3224) );
  NAND2_X1 U8668 ( .A1(n7016), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n7011) );
  NAND2_X1 U8669 ( .A1(n7011), .A2(n7010), .ZN(n7014) );
  INV_X1 U8670 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7012) );
  MUX2_X1 U8671 ( .A(n7012), .B(P2_REG2_REG_11__SCAN_IN), .S(n7162), .Z(n7013)
         );
  NOR2_X1 U8672 ( .A1(n7014), .A2(n7013), .ZN(n7153) );
  AOI21_X1 U8673 ( .B1(n7014), .B2(n7013), .A(n7153), .ZN(n7024) );
  NOR2_X1 U8674 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9881), .ZN(n7021) );
  INV_X1 U8675 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n7017) );
  MUX2_X1 U8676 ( .A(n7017), .B(P2_REG1_REG_11__SCAN_IN), .S(n7162), .Z(n7018)
         );
  AOI211_X1 U8677 ( .C1(n7019), .C2(n7018), .A(n7161), .B(n9528), .ZN(n7020)
         );
  AOI211_X1 U8678 ( .C1(P2_ADDR_REG_11__SCAN_IN), .C2(n9734), .A(n7021), .B(
        n7020), .ZN(n7023) );
  INV_X1 U8679 ( .A(n9730), .ZN(n9534) );
  NAND2_X1 U8680 ( .A1(n9534), .A2(n7162), .ZN(n7022) );
  OAI211_X1 U8681 ( .C1(n7024), .C2(n9732), .A(n7023), .B(n7022), .ZN(P2_U3256) );
  NAND2_X1 U8682 ( .A1(n7025), .A2(n7026), .ZN(n7027) );
  NAND2_X1 U8683 ( .A1(n7028), .A2(n7027), .ZN(n7354) );
  NAND2_X1 U8684 ( .A1(n7030), .A2(n7355), .ZN(n9739) );
  NAND2_X1 U8685 ( .A1(n7354), .A2(n8176), .ZN(n7353) );
  NAND2_X1 U8686 ( .A1(n7030), .A2(n9776), .ZN(n7031) );
  NAND2_X1 U8687 ( .A1(n7353), .A2(n7031), .ZN(n9752) );
  INV_X1 U8688 ( .A(n9749), .ZN(n7032) );
  NAND2_X1 U8689 ( .A1(n8379), .A2(n7032), .ZN(n8208) );
  NAND2_X1 U8690 ( .A1(n8212), .A2(n8208), .ZN(n9753) );
  NAND2_X1 U8691 ( .A1(n9752), .A2(n9753), .ZN(n7034) );
  NAND2_X1 U8692 ( .A1(n7359), .A2(n7032), .ZN(n7033) );
  NAND2_X1 U8693 ( .A1(n7034), .A2(n7033), .ZN(n7035) );
  NAND2_X1 U8694 ( .A1(n7195), .A2(n7045), .ZN(n8213) );
  NAND2_X1 U8695 ( .A1(n8213), .A2(n8209), .ZN(n8178) );
  NAND2_X1 U8696 ( .A1(n7035), .A2(n8178), .ZN(n7197) );
  OAI21_X1 U8697 ( .B1(n7035), .B2(n8178), .A(n7197), .ZN(n9792) );
  INV_X1 U8698 ( .A(n9792), .ZN(n7055) );
  INV_X1 U8699 ( .A(n7036), .ZN(n7039) );
  AND2_X1 U8700 ( .A1(n7037), .A2(n7272), .ZN(n7038) );
  NAND2_X1 U8701 ( .A1(n7039), .A2(n7038), .ZN(n7042) );
  OR2_X1 U8702 ( .A1(n7040), .A2(n8569), .ZN(n7209) );
  NAND2_X1 U8703 ( .A1(n8780), .A2(n7209), .ZN(n7041) );
  NAND2_X1 U8704 ( .A1(n8830), .A2(n7041), .ZN(n8764) );
  NAND2_X1 U8705 ( .A1(n7352), .A2(n9776), .ZN(n9748) );
  OR2_X1 U8706 ( .A1(n7042), .A2(n8356), .ZN(n7706) );
  NAND2_X1 U8707 ( .A1(n8830), .A2(n7044), .ZN(n8821) );
  INV_X1 U8708 ( .A(n8821), .ZN(n8827) );
  AOI22_X1 U8709 ( .A1(n9787), .A2(n7043), .B1(n8827), .B2(n7045), .ZN(n7054)
         );
  NAND2_X1 U8710 ( .A1(n7092), .A2(n7046), .ZN(n8217) );
  INV_X1 U8711 ( .A(n9753), .ZN(n8220) );
  INV_X1 U8712 ( .A(n8178), .ZN(n7047) );
  XNOR2_X1 U8713 ( .A(n7211), .B(n7047), .ZN(n7048) );
  NAND2_X1 U8714 ( .A1(n7048), .A2(n8813), .ZN(n7050) );
  AOI22_X1 U8715 ( .A1(n9743), .A2(n8379), .B1(n8810), .B2(n9744), .ZN(n7049)
         );
  NAND2_X1 U8716 ( .A1(n7050), .A2(n7049), .ZN(n9790) );
  OAI22_X1 U8717 ( .A1(n7668), .A2(n7051), .B1(n6887), .B2(n8830), .ZN(n7052)
         );
  AOI21_X1 U8718 ( .B1(n8830), .B2(n9790), .A(n7052), .ZN(n7053) );
  OAI211_X1 U8719 ( .C1(n7055), .C2(n8764), .A(n7054), .B(n7053), .ZN(P2_U3292) );
  OAI21_X1 U8720 ( .B1(n7058), .B2(n7057), .A(n7056), .ZN(n7063) );
  INV_X1 U8721 ( .A(n9106), .ZN(n9071) );
  AOI22_X1 U8722 ( .A1(n9094), .A2(n9130), .B1(n9112), .B2(n7124), .ZN(n7061)
         );
  NAND2_X1 U8723 ( .A1(P1_U3084), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9147) );
  INV_X1 U8724 ( .A(n9147), .ZN(n7059) );
  AOI21_X1 U8725 ( .B1(n9104), .B2(n9132), .A(n7059), .ZN(n7060) );
  OAI211_X1 U8726 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n9071), .A(n7061), .B(
        n7060), .ZN(n7062) );
  AOI21_X1 U8727 ( .B1(n7063), .B2(n9087), .A(n7062), .ZN(n7064) );
  INV_X1 U8728 ( .A(n7064), .ZN(P1_U3216) );
  INV_X1 U8729 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n7071) );
  INV_X1 U8730 ( .A(n9770), .ZN(n7066) );
  NOR2_X1 U8731 ( .A1(n8146), .A2(n7066), .ZN(n7069) );
  NAND2_X1 U8732 ( .A1(n8380), .A2(n7066), .ZN(n8225) );
  MUX2_X1 U8733 ( .A(n8225), .B(n7066), .S(n7065), .Z(n7067) );
  AOI21_X1 U8734 ( .B1(n7092), .B2(n7067), .A(n5614), .ZN(n7068) );
  AOI211_X1 U8735 ( .C1(n8143), .C2(n6817), .A(n7069), .B(n7068), .ZN(n7070)
         );
  OAI21_X1 U8736 ( .B1(n7072), .B2(n7071), .A(n7070), .ZN(P2_U3234) );
  XNOR2_X1 U8737 ( .A(n7074), .B(n7073), .ZN(n7078) );
  INV_X1 U8738 ( .A(n7281), .ZN(n7329) );
  OAI22_X1 U8739 ( .A1(n8146), .A2(n7329), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8439), .ZN(n7076) );
  OAI22_X1 U8740 ( .A1(n7212), .A2(n8160), .B1(n8159), .B2(n7656), .ZN(n7075)
         );
  AOI211_X1 U8741 ( .C1(n7331), .C2(n5616), .A(n7076), .B(n7075), .ZN(n7077)
         );
  OAI21_X1 U8742 ( .B1(n7078), .B2(n5614), .A(n7077), .ZN(P2_U3215) );
  NAND2_X1 U8743 ( .A1(n7080), .A2(n7079), .ZN(n7081) );
  XNOR2_X1 U8744 ( .A(n7082), .B(n7081), .ZN(n7087) );
  AOI22_X1 U8745 ( .A1(n9094), .A2(n9129), .B1(n9112), .B2(n7144), .ZN(n7086)
         );
  NOR2_X1 U8746 ( .A1(n9092), .A2(n7134), .ZN(n7083) );
  AOI211_X1 U8747 ( .C1(n7174), .C2(n9106), .A(n7084), .B(n7083), .ZN(n7085)
         );
  OAI211_X1 U8748 ( .C1(n7087), .C2(n9115), .A(n7086), .B(n7085), .ZN(P1_U3228) );
  INV_X1 U8749 ( .A(n7088), .ZN(n7091) );
  AOI22_X1 U8750 ( .A1(n9175), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n9506), .ZN(n7089) );
  OAI21_X1 U8751 ( .B1(n7091), .B2(n9508), .A(n7089), .ZN(P1_U3335) );
  AOI22_X1 U8752 ( .A1(n8560), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n8969), .ZN(n7090) );
  OAI21_X1 U8753 ( .B1(n7091), .B2(n8967), .A(n7090), .ZN(P2_U3340) );
  INV_X1 U8754 ( .A(n7043), .ZN(n8582) );
  NAND2_X1 U8755 ( .A1(n8582), .A2(n8821), .ZN(n9755) );
  INV_X1 U8756 ( .A(n8764), .ZN(n9754) );
  NAND2_X1 U8757 ( .A1(n7092), .A2(n8225), .ZN(n9769) );
  INV_X1 U8758 ( .A(n9769), .ZN(n7097) );
  NAND2_X1 U8759 ( .A1(n9769), .A2(n8813), .ZN(n7094) );
  NAND2_X1 U8760 ( .A1(n6817), .A2(n9744), .ZN(n7093) );
  NAND2_X1 U8761 ( .A1(n7094), .A2(n7093), .ZN(n9774) );
  AOI22_X1 U8762 ( .A1(n8830), .A2(n9774), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        n9747), .ZN(n7096) );
  INV_X1 U8763 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n9955) );
  OR2_X1 U8764 ( .A1(n8830), .A2(n9955), .ZN(n7095) );
  OAI211_X1 U8765 ( .C1(n8764), .C2(n7097), .A(n7096), .B(n7095), .ZN(n7098)
         );
  AOI21_X1 U8766 ( .B1(n9755), .B2(n9770), .A(n7098), .ZN(n7099) );
  INV_X1 U8767 ( .A(n7099), .ZN(P2_U3296) );
  XNOR2_X1 U8768 ( .A(n7100), .B(n7101), .ZN(n7105) );
  NAND2_X1 U8769 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3152), .ZN(n8453) );
  OAI21_X1 U8770 ( .B1(n8146), .B2(n4517), .A(n8453), .ZN(n7103) );
  OAI22_X1 U8771 ( .A1(n7203), .A2(n8160), .B1(n8159), .B2(n7456), .ZN(n7102)
         );
  AOI211_X1 U8772 ( .C1(n7217), .C2(n5616), .A(n7103), .B(n7102), .ZN(n7104)
         );
  OAI21_X1 U8773 ( .B1(n7105), .B2(n5614), .A(n7104), .ZN(P2_U3223) );
  INV_X1 U8774 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n7112) );
  INV_X1 U8775 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n7107) );
  OAI21_X1 U8776 ( .B1(n7107), .B2(n9692), .A(n7106), .ZN(n7108) );
  NAND2_X1 U8777 ( .A1(n7108), .A2(n9688), .ZN(n7111) );
  OAI21_X1 U8778 ( .B1(n9316), .B2(n9409), .A(n7109), .ZN(n7110) );
  OAI211_X1 U8779 ( .C1(n7112), .C2(n9688), .A(n7111), .B(n7110), .ZN(P1_U3291) );
  OAI21_X1 U8780 ( .B1(n7114), .B2(n7115), .A(n7113), .ZN(n9711) );
  INV_X1 U8781 ( .A(n9711), .ZN(n7127) );
  XNOR2_X1 U8782 ( .A(n7116), .B(n7115), .ZN(n7119) );
  OAI22_X1 U8783 ( .A1(n7262), .A2(n9333), .B1(n6309), .B2(n9331), .ZN(n7117)
         );
  AOI21_X1 U8784 ( .B1(n9711), .B2(n7625), .A(n7117), .ZN(n7118) );
  OAI21_X1 U8785 ( .B1(n9329), .B2(n7119), .A(n7118), .ZN(n9709) );
  NAND2_X1 U8786 ( .A1(n9709), .A2(n9688), .ZN(n7126) );
  OAI22_X1 U8787 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(n9692), .B1(n6555), .B2(
        n9688), .ZN(n7123) );
  INV_X1 U8788 ( .A(n9409), .ZN(n9319) );
  AND2_X1 U8789 ( .A1(n7120), .A2(n7124), .ZN(n7121) );
  OR2_X1 U8790 ( .A1(n7121), .A2(n7141), .ZN(n9708) );
  NOR2_X1 U8791 ( .A1(n9319), .A2(n9708), .ZN(n7122) );
  AOI211_X1 U8792 ( .C1(n9316), .C2(n7124), .A(n7123), .B(n7122), .ZN(n7125)
         );
  OAI211_X1 U8793 ( .C1(n7127), .C2(n7237), .A(n7126), .B(n7125), .ZN(P1_U3288) );
  INV_X1 U8794 ( .A(n7128), .ZN(n7130) );
  OAI222_X1 U8795 ( .A1(P1_U3084), .A2(n9682), .B1(n9508), .B2(n7130), .C1(
        n7129), .C2(n9510), .ZN(P1_U3334) );
  OAI222_X1 U8796 ( .A1(n7990), .A2(n7131), .B1(n8967), .B2(n7130), .C1(n8569), 
        .C2(P2_U3152), .ZN(P2_U3339) );
  INV_X1 U8797 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n10040) );
  OAI21_X1 U8798 ( .B1(n7133), .B2(n7138), .A(n7132), .ZN(n7180) );
  INV_X1 U8799 ( .A(n7180), .ZN(n7146) );
  OAI22_X1 U8800 ( .A1(n7441), .A2(n9333), .B1(n7134), .B2(n9331), .ZN(n7140)
         );
  INV_X1 U8801 ( .A(n7135), .ZN(n7136) );
  AOI211_X1 U8802 ( .C1(n7138), .C2(n7137), .A(n9329), .B(n7136), .ZN(n7139)
         );
  AOI211_X1 U8803 ( .C1(n7625), .C2(n7180), .A(n7140), .B(n7139), .ZN(n7183)
         );
  INV_X1 U8804 ( .A(n7141), .ZN(n7143) );
  INV_X1 U8805 ( .A(n7254), .ZN(n7142) );
  AOI21_X1 U8806 ( .B1(n7144), .B2(n7143), .A(n7142), .ZN(n7179) );
  AOI22_X1 U8807 ( .A1(n7179), .A2(n9559), .B1(n9483), .B2(n7144), .ZN(n7145)
         );
  OAI211_X1 U8808 ( .C1(n7146), .C2(n7247), .A(n7183), .B(n7145), .ZN(n7148)
         );
  NAND2_X1 U8809 ( .A1(n7148), .A2(n9486), .ZN(n7147) );
  OAI21_X1 U8810 ( .B1(n9486), .B2(n10040), .A(n7147), .ZN(P1_U3527) );
  INV_X1 U8811 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n7150) );
  NAND2_X1 U8812 ( .A1(n7148), .A2(n9722), .ZN(n7149) );
  OAI21_X1 U8813 ( .B1(n9722), .B2(n7150), .A(n7149), .ZN(P1_U3466) );
  NAND2_X1 U8814 ( .A1(n8483), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n7155) );
  INV_X1 U8815 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7151) );
  MUX2_X1 U8816 ( .A(n7151), .B(P2_REG2_REG_12__SCAN_IN), .S(n8483), .Z(n7152)
         );
  INV_X1 U8817 ( .A(n7152), .ZN(n8479) );
  AOI21_X1 U8818 ( .B1(n7154), .B2(n7012), .A(n7153), .ZN(n8480) );
  NAND2_X1 U8819 ( .A1(n8479), .A2(n8480), .ZN(n8478) );
  NAND2_X1 U8820 ( .A1(n7155), .A2(n8478), .ZN(n7158) );
  INV_X1 U8821 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n7156) );
  AOI22_X1 U8822 ( .A1(n7318), .A2(n7156), .B1(P2_REG2_REG_13__SCAN_IN), .B2(
        n7159), .ZN(n7157) );
  NOR2_X1 U8823 ( .A1(n7158), .A2(n7157), .ZN(n7312) );
  AOI21_X1 U8824 ( .B1(n7158), .B2(n7157), .A(n7312), .ZN(n7172) );
  INV_X1 U8825 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n7160) );
  AOI22_X1 U8826 ( .A1(n7318), .A2(P2_REG1_REG_13__SCAN_IN), .B1(n7160), .B2(
        n7159), .ZN(n7165) );
  INV_X1 U8827 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7163) );
  MUX2_X1 U8828 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n7163), .S(n8483), .Z(n8486)
         );
  OAI21_X1 U8829 ( .B1(n8483), .B2(P2_REG1_REG_12__SCAN_IN), .A(n8484), .ZN(
        n7164) );
  NAND2_X1 U8830 ( .A1(n7165), .A2(n7164), .ZN(n7317) );
  OAI21_X1 U8831 ( .B1(n7165), .B2(n7164), .A(n7317), .ZN(n7166) );
  NAND2_X1 U8832 ( .A1(n7166), .A2(n9729), .ZN(n7171) );
  INV_X1 U8833 ( .A(n9734), .ZN(n7323) );
  INV_X1 U8834 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7168) );
  OAI22_X1 U8835 ( .A1(n7323), .A2(n7168), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7167), .ZN(n7169) );
  AOI21_X1 U8836 ( .B1(n9534), .B2(n7318), .A(n7169), .ZN(n7170) );
  OAI211_X1 U8837 ( .C1(n7172), .C2(n9732), .A(n7171), .B(n7170), .ZN(P2_U3258) );
  NOR2_X1 U8838 ( .A1(n9396), .A2(n7173), .ZN(n7178) );
  INV_X1 U8839 ( .A(n7174), .ZN(n7175) );
  OAI22_X1 U8840 ( .A1(n9688), .A2(n7176), .B1(n7175), .B2(n9692), .ZN(n7177)
         );
  AOI211_X1 U8841 ( .C1(n7179), .C2(n9409), .A(n7178), .B(n7177), .ZN(n7182)
         );
  NAND2_X1 U8842 ( .A1(n7180), .A2(n7632), .ZN(n7181) );
  OAI211_X1 U8843 ( .C1(n7183), .C2(n6638), .A(n7182), .B(n7181), .ZN(P1_U3287) );
  INV_X1 U8844 ( .A(n7184), .ZN(n7189) );
  INV_X1 U8845 ( .A(n7185), .ZN(n7188) );
  AOI22_X1 U8846 ( .A1(n7186), .A2(n9559), .B1(n9483), .B2(n7440), .ZN(n7187)
         );
  OAI211_X1 U8847 ( .C1(n7189), .C2(n7247), .A(n7188), .B(n7187), .ZN(n7192)
         );
  NAND2_X1 U8848 ( .A1(n7192), .A2(n9486), .ZN(n7190) );
  OAI21_X1 U8849 ( .B1(n9486), .B2(n7191), .A(n7190), .ZN(P1_U3529) );
  INV_X1 U8850 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n7194) );
  NAND2_X1 U8851 ( .A1(n7192), .A2(n9722), .ZN(n7193) );
  OAI21_X1 U8852 ( .B1(n9722), .B2(n7194), .A(n7193), .ZN(P1_U3472) );
  NAND2_X1 U8853 ( .A1(n7195), .A2(n9788), .ZN(n7196) );
  NAND2_X1 U8854 ( .A1(n7197), .A2(n7196), .ZN(n7399) );
  NAND2_X1 U8855 ( .A1(n7399), .A2(n8180), .ZN(n7200) );
  NAND2_X1 U8856 ( .A1(n7198), .A2(n7403), .ZN(n7199) );
  NAND2_X1 U8857 ( .A1(n7200), .A2(n7199), .ZN(n8818) );
  NOR2_X1 U8858 ( .A1(n8378), .A2(n9801), .ZN(n7202) );
  NAND2_X1 U8859 ( .A1(n8378), .A2(n9801), .ZN(n7201) );
  OAI21_X1 U8860 ( .B1(n8818), .B2(n7202), .A(n7201), .ZN(n7275) );
  NAND2_X1 U8861 ( .A1(n7329), .A2(n8811), .ZN(n8241) );
  NAND2_X1 U8862 ( .A1(n7203), .A2(n7281), .ZN(n8246) );
  NAND2_X1 U8863 ( .A1(n7329), .A2(n7203), .ZN(n7204) );
  OAI21_X1 U8864 ( .B1(n7275), .B2(n8239), .A(n7204), .ZN(n7206) );
  INV_X1 U8865 ( .A(n7206), .ZN(n7205) );
  OR2_X1 U8866 ( .A1(n7656), .A2(n7448), .ZN(n8249) );
  NAND2_X1 U8867 ( .A1(n7448), .A2(n7656), .ZN(n8242) );
  NAND2_X1 U8868 ( .A1(n7207), .A2(n8247), .ZN(n7208) );
  NAND2_X1 U8869 ( .A1(n7658), .A2(n7208), .ZN(n9810) );
  INV_X2 U8870 ( .A(n8830), .ZN(n8804) );
  OR2_X1 U8871 ( .A1(n8804), .A2(n7209), .ZN(n8790) );
  AOI22_X1 U8872 ( .A1(n9743), .A2(n8811), .B1(n8376), .B2(n9744), .ZN(n7216)
         );
  INV_X1 U8873 ( .A(n8213), .ZN(n7210) );
  INV_X1 U8874 ( .A(n8207), .ZN(n8211) );
  NAND2_X1 U8875 ( .A1(n7212), .A2(n9801), .ZN(n8237) );
  NAND2_X1 U8876 ( .A1(n8820), .A2(n8378), .ZN(n8231) );
  NAND2_X1 U8877 ( .A1(n8809), .A2(n8819), .ZN(n8808) );
  NAND2_X1 U8878 ( .A1(n8808), .A2(n8237), .ZN(n7277) );
  NAND2_X1 U8879 ( .A1(n7277), .A2(n8239), .ZN(n7276) );
  OAI21_X1 U8880 ( .B1(n8247), .B2(n7213), .A(n7454), .ZN(n7214) );
  NAND2_X1 U8881 ( .A1(n7214), .A2(n8813), .ZN(n7215) );
  OAI211_X1 U8882 ( .C1(n9810), .C2(n8780), .A(n7216), .B(n7215), .ZN(n9814)
         );
  NAND2_X1 U8883 ( .A1(n9814), .A2(n8830), .ZN(n7223) );
  INV_X1 U8884 ( .A(n7217), .ZN(n7218) );
  OAI22_X1 U8885 ( .A1(n8830), .A2(n9878), .B1(n7218), .B2(n7668), .ZN(n7221)
         );
  AND2_X1 U8886 ( .A1(n7400), .A2(n7403), .ZN(n8814) );
  NAND2_X1 U8887 ( .A1(n8814), .A2(n8820), .ZN(n8816) );
  NAND2_X1 U8888 ( .A1(n7279), .A2(n7448), .ZN(n7219) );
  NAND2_X1 U8889 ( .A1(n7666), .A2(n7219), .ZN(n9811) );
  NOR2_X1 U8890 ( .A1(n8582), .A2(n9811), .ZN(n7220) );
  AOI211_X1 U8891 ( .C1(n8827), .C2(n7448), .A(n7221), .B(n7220), .ZN(n7222)
         );
  OAI211_X1 U8892 ( .C1(n9810), .C2(n8790), .A(n7223), .B(n7222), .ZN(P2_U3288) );
  XNOR2_X1 U8893 ( .A(n7228), .B(n7224), .ZN(n9704) );
  INV_X1 U8894 ( .A(n9704), .ZN(n7238) );
  XNOR2_X1 U8895 ( .A(n7225), .B(n7234), .ZN(n7226) );
  NAND2_X1 U8896 ( .A1(n7226), .A2(n9559), .ZN(n9699) );
  OAI21_X1 U8897 ( .B1(n7228), .B2(n7227), .A(n9406), .ZN(n7230) );
  OAI22_X1 U8898 ( .A1(n7230), .A2(n7229), .B1(n6309), .B2(n9333), .ZN(n7231)
         );
  AOI21_X1 U8899 ( .B1(n7625), .B2(n9704), .A(n7231), .ZN(n9701) );
  INV_X1 U8900 ( .A(n9692), .ZN(n9393) );
  AND2_X1 U8901 ( .A1(n6306), .A2(n9401), .ZN(n9698) );
  AOI21_X1 U8902 ( .B1(n9393), .B2(P1_REG3_REG_1__SCAN_IN), .A(n9698), .ZN(
        n7232) );
  OAI211_X1 U8903 ( .C1(n9282), .C2(n9699), .A(n9701), .B(n7232), .ZN(n7233)
         );
  NAND2_X1 U8904 ( .A1(n7233), .A2(n9688), .ZN(n7236) );
  AOI22_X1 U8905 ( .A1(n9316), .A2(n7234), .B1(n6638), .B2(
        P1_REG2_REG_1__SCAN_IN), .ZN(n7235) );
  OAI211_X1 U8906 ( .C1(n7238), .C2(n7237), .A(n7236), .B(n7235), .ZN(P1_U3290) );
  INV_X1 U8907 ( .A(n7240), .ZN(n7241) );
  AOI21_X1 U8908 ( .B1(n7239), .B2(n7242), .A(n7241), .ZN(n7246) );
  INV_X1 U8909 ( .A(n7772), .ZN(n7672) );
  NAND2_X1 U8910 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3152), .ZN(n8467) );
  OAI21_X1 U8911 ( .B1(n8146), .B2(n7672), .A(n8467), .ZN(n7244) );
  INV_X1 U8912 ( .A(n8375), .ZN(n7655) );
  OAI22_X1 U8913 ( .A1(n7656), .A2(n8160), .B1(n8159), .B2(n7655), .ZN(n7243)
         );
  AOI211_X1 U8914 ( .C1(n7667), .C2(n5616), .A(n7244), .B(n7243), .ZN(n7245)
         );
  OAI21_X1 U8915 ( .B1(n7246), .B2(n5614), .A(n7245), .ZN(P2_U3233) );
  OAI21_X1 U8916 ( .B1(n7250), .B2(n6625), .A(n7249), .ZN(n9686) );
  XOR2_X1 U8917 ( .A(n7252), .B(n7251), .Z(n7253) );
  AOI222_X1 U8918 ( .A1(n9406), .A2(n7253), .B1(n9130), .B2(n9401), .C1(n9128), 
        .C2(n9403), .ZN(n9685) );
  AOI21_X1 U8919 ( .B1(n7254), .B2(n9680), .A(n9707), .ZN(n7256) );
  AND2_X1 U8920 ( .A1(n7256), .A2(n7255), .ZN(n9683) );
  AOI21_X1 U8921 ( .B1(n9483), .B2(n9680), .A(n9683), .ZN(n7257) );
  OAI211_X1 U8922 ( .C1(n9561), .C2(n9686), .A(n9685), .B(n7257), .ZN(n7269)
         );
  NAND2_X1 U8923 ( .A1(n7269), .A2(n9486), .ZN(n7258) );
  OAI21_X1 U8924 ( .B1(n9486), .B2(n7259), .A(n7258), .ZN(P1_U3528) );
  XNOR2_X1 U8925 ( .A(n7434), .B(n7435), .ZN(n7261) );
  NOR2_X1 U8926 ( .A1(n7261), .A2(n7260), .ZN(n7433) );
  AOI21_X1 U8927 ( .B1(n7261), .B2(n7260), .A(n7433), .ZN(n7268) );
  AOI22_X1 U8928 ( .A1(n9094), .A2(n9128), .B1(n9112), .B2(n9680), .ZN(n7267)
         );
  NOR2_X1 U8929 ( .A1(n9092), .A2(n7262), .ZN(n7263) );
  AOI211_X1 U8930 ( .C1(n7265), .C2(n9106), .A(n7264), .B(n7263), .ZN(n7266)
         );
  OAI211_X1 U8931 ( .C1(n7268), .C2(n9115), .A(n7267), .B(n7266), .ZN(P1_U3225) );
  INV_X1 U8932 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n7271) );
  NAND2_X1 U8933 ( .A1(n7269), .A2(n9722), .ZN(n7270) );
  OAI21_X1 U8934 ( .B1(n9722), .B2(n7271), .A(n7270), .ZN(P1_U3469) );
  INV_X1 U8935 ( .A(n7272), .ZN(n7273) );
  AND2_X2 U8936 ( .A1(n7274), .A2(n7273), .ZN(n9848) );
  XOR2_X1 U8937 ( .A(n7275), .B(n8239), .Z(n7339) );
  OAI21_X1 U8938 ( .B1(n8239), .B2(n7277), .A(n7276), .ZN(n7278) );
  AOI222_X1 U8939 ( .A1(n8813), .A2(n7278), .B1(n8377), .B2(n9744), .C1(n8378), 
        .C2(n9743), .ZN(n7328) );
  AOI21_X1 U8940 ( .B1(n8816), .B2(n7281), .A(n9825), .ZN(n7280) );
  AND2_X1 U8941 ( .A1(n7280), .A2(n7279), .ZN(n7330) );
  AOI21_X1 U8942 ( .B1(n9802), .B2(n7281), .A(n7330), .ZN(n7282) );
  OAI211_X1 U8943 ( .C1(n9797), .C2(n7339), .A(n7328), .B(n7282), .ZN(n7284)
         );
  NAND2_X1 U8944 ( .A1(n7284), .A2(n9848), .ZN(n7283) );
  OAI21_X1 U8945 ( .B1(n9848), .B2(n6871), .A(n7283), .ZN(P2_U3527) );
  INV_X1 U8946 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n7286) );
  NAND2_X1 U8947 ( .A1(n7284), .A2(n9833), .ZN(n7285) );
  OAI21_X1 U8948 ( .B1(n9833), .B2(n7286), .A(n7285), .ZN(P2_U3472) );
  INV_X1 U8949 ( .A(n7287), .ZN(n7935) );
  OAI222_X1 U8950 ( .A1(n7990), .A2(n7288), .B1(P2_U3152), .B2(n8343), .C1(
        n8967), .C2(n7935), .ZN(P2_U3338) );
  NAND2_X1 U8951 ( .A1(n7367), .A2(n7292), .ZN(n7293) );
  XNOR2_X1 U8952 ( .A(n7293), .B(n7302), .ZN(n7294) );
  OAI222_X1 U8953 ( .A1(n9331), .A2(n7300), .B1(n9333), .B2(n7295), .C1(n7294), 
        .C2(n9329), .ZN(n7412) );
  INV_X1 U8954 ( .A(n7412), .ZN(n7311) );
  NAND2_X1 U8955 ( .A1(n7297), .A2(n7296), .ZN(n7298) );
  NAND2_X1 U8956 ( .A1(n7388), .A2(n7387), .ZN(n7386) );
  NAND2_X1 U8957 ( .A1(n7300), .A2(n7469), .ZN(n7301) );
  OAI21_X1 U8958 ( .B1(n4388), .B2(n7302), .A(n7365), .ZN(n7303) );
  INV_X1 U8959 ( .A(n7303), .ZN(n7414) );
  AND2_X1 U8960 ( .A1(n7305), .A2(n7304), .ZN(n9679) );
  NAND2_X1 U8961 ( .A1(n9688), .A2(n9679), .ZN(n9411) );
  INV_X1 U8962 ( .A(n9411), .ZN(n7915) );
  NOR2_X1 U8963 ( .A1(n7390), .A2(n7487), .ZN(n7389) );
  NAND2_X1 U8964 ( .A1(n7389), .A2(n7411), .ZN(n7375) );
  OAI211_X1 U8965 ( .C1(n7389), .C2(n7411), .A(n9559), .B(n7375), .ZN(n7410)
         );
  AND2_X1 U8966 ( .A1(n9688), .A2(n9682), .ZN(n9335) );
  INV_X1 U8967 ( .A(n9335), .ZN(n7883) );
  INV_X1 U8968 ( .A(n7539), .ZN(n7306) );
  OAI22_X1 U8969 ( .A1(n9688), .A2(n6566), .B1(n7306), .B2(n9692), .ZN(n7307)
         );
  AOI21_X1 U8970 ( .B1(n9316), .B2(n7538), .A(n7307), .ZN(n7308) );
  OAI21_X1 U8971 ( .B1(n7410), .B2(n7883), .A(n7308), .ZN(n7309) );
  AOI21_X1 U8972 ( .B1(n7414), .B2(n7915), .A(n7309), .ZN(n7310) );
  OAI21_X1 U8973 ( .B1(n7311), .B2(n6638), .A(n7310), .ZN(P1_U3283) );
  NOR2_X1 U8974 ( .A1(n7318), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n7313) );
  NOR2_X1 U8975 ( .A1(n7313), .A2(n7312), .ZN(n7315) );
  INV_X1 U8976 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n8497) );
  AOI22_X1 U8977 ( .A1(n8493), .A2(n8497), .B1(P2_REG2_REG_14__SCAN_IN), .B2(
        n8498), .ZN(n7314) );
  NOR2_X1 U8978 ( .A1(n7315), .A2(n7314), .ZN(n8496) );
  AOI21_X1 U8979 ( .B1(n7315), .B2(n7314), .A(n8496), .ZN(n7327) );
  INV_X1 U8980 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n7316) );
  AOI22_X1 U8981 ( .A1(n8493), .A2(P2_REG1_REG_14__SCAN_IN), .B1(n7316), .B2(
        n8498), .ZN(n7320) );
  OAI21_X1 U8982 ( .B1(n7318), .B2(P2_REG1_REG_13__SCAN_IN), .A(n7317), .ZN(
        n7319) );
  NAND2_X1 U8983 ( .A1(n7320), .A2(n7319), .ZN(n8492) );
  OAI21_X1 U8984 ( .B1(n7320), .B2(n7319), .A(n8492), .ZN(n7321) );
  NAND2_X1 U8985 ( .A1(n7321), .A2(n9729), .ZN(n7326) );
  INV_X1 U8986 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7322) );
  NAND2_X1 U8987 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3152), .ZN(n7818) );
  OAI21_X1 U8988 ( .B1(n7323), .B2(n7322), .A(n7818), .ZN(n7324) );
  AOI21_X1 U8989 ( .B1(n9534), .B2(n8493), .A(n7324), .ZN(n7325) );
  OAI211_X1 U8990 ( .C1(n7327), .C2(n9732), .A(n7326), .B(n7325), .ZN(P2_U3259) );
  NOR2_X1 U8991 ( .A1(n7328), .A2(n8804), .ZN(n7337) );
  NOR2_X1 U8992 ( .A1(n8821), .A2(n7329), .ZN(n7336) );
  NOR2_X1 U8993 ( .A1(n8830), .A2(n6897), .ZN(n7335) );
  INV_X1 U8994 ( .A(n7330), .ZN(n7333) );
  INV_X1 U8995 ( .A(n7331), .ZN(n7332) );
  OAI22_X1 U8996 ( .A1(n7706), .A2(n7333), .B1(n7332), .B2(n7668), .ZN(n7334)
         );
  NOR4_X1 U8997 ( .A1(n7337), .A2(n7336), .A3(n7335), .A4(n7334), .ZN(n7338)
         );
  OAI21_X1 U8998 ( .B1(n8764), .B2(n7339), .A(n7338), .ZN(P2_U3289) );
  INV_X1 U8999 ( .A(n7340), .ZN(n7350) );
  OAI222_X1 U9000 ( .A1(n7342), .A2(P1_U3084), .B1(n9508), .B2(n7350), .C1(
        n7341), .C2(n9510), .ZN(P1_U3332) );
  XNOR2_X1 U9001 ( .A(n7344), .B(n7343), .ZN(n7349) );
  INV_X1 U9002 ( .A(n7634), .ZN(n9817) );
  OAI21_X1 U9003 ( .B1(n8146), .B2(n9817), .A(n7345), .ZN(n7347) );
  INV_X1 U9004 ( .A(n8374), .ZN(n7637) );
  OAI22_X1 U9005 ( .A1(n7456), .A2(n8160), .B1(n8159), .B2(n7637), .ZN(n7346)
         );
  AOI211_X1 U9006 ( .C1(n7460), .C2(n5616), .A(n7347), .B(n7346), .ZN(n7348)
         );
  OAI21_X1 U9007 ( .B1(n7349), .B2(n5614), .A(n7348), .ZN(P2_U3219) );
  OAI222_X1 U9008 ( .A1(n7990), .A2(n7351), .B1(P2_U3152), .B2(n8201), .C1(
        n8967), .C2(n7350), .ZN(P2_U3337) );
  OAI21_X1 U9009 ( .B1(n7352), .B2(n9776), .A(n9748), .ZN(n9777) );
  OAI21_X1 U9010 ( .B1(n7354), .B2(n8176), .A(n7353), .ZN(n9780) );
  AOI22_X1 U9011 ( .A1(n9754), .A2(n9780), .B1(n8827), .B2(n7355), .ZN(n7363)
         );
  INV_X1 U9012 ( .A(n9740), .ZN(n7356) );
  AOI21_X1 U9013 ( .B1(n8176), .B2(n7357), .A(n7356), .ZN(n7358) );
  OAI222_X1 U9014 ( .A1(n8754), .A2(n7359), .B1(n8756), .B2(n7025), .C1(n8751), 
        .C2(n7358), .ZN(n9778) );
  AOI22_X1 U9015 ( .A1(n9747), .A2(P2_REG3_REG_2__SCAN_IN), .B1(
        P2_REG2_REG_2__SCAN_IN), .B2(n8804), .ZN(n7360) );
  INV_X1 U9016 ( .A(n7360), .ZN(n7361) );
  AOI21_X1 U9017 ( .B1(n9778), .B2(n8830), .A(n7361), .ZN(n7362) );
  OAI211_X1 U9018 ( .C1(n8582), .C2(n9777), .A(n7363), .B(n7362), .ZN(P2_U3294) );
  NAND2_X1 U9019 ( .A1(n9126), .A2(n7538), .ZN(n7364) );
  XNOR2_X1 U9020 ( .A(n7496), .B(n7370), .ZN(n9718) );
  NAND2_X1 U9021 ( .A1(n7367), .A2(n7366), .ZN(n7369) );
  XNOR2_X1 U9022 ( .A(n7498), .B(n7370), .ZN(n7373) );
  OAI22_X1 U9023 ( .A1(n7620), .A2(n9333), .B1(n7480), .B2(n9331), .ZN(n7371)
         );
  INV_X1 U9024 ( .A(n7371), .ZN(n7372) );
  OAI21_X1 U9025 ( .B1(n7373), .B2(n9329), .A(n7372), .ZN(n7374) );
  AOI21_X1 U9026 ( .B1(n9718), .B2(n7625), .A(n7374), .ZN(n9720) );
  AOI21_X1 U9027 ( .B1(n7375), .B2(n7520), .A(n9707), .ZN(n7376) );
  NAND2_X1 U9028 ( .A1(n7376), .A2(n7505), .ZN(n9713) );
  INV_X1 U9029 ( .A(n7516), .ZN(n7377) );
  OAI22_X1 U9030 ( .A1(n9688), .A2(n6551), .B1(n7377), .B2(n9692), .ZN(n7378)
         );
  AOI21_X1 U9031 ( .B1(n9316), .B2(n7520), .A(n7378), .ZN(n7379) );
  OAI21_X1 U9032 ( .B1(n9713), .B2(n7883), .A(n7379), .ZN(n7380) );
  AOI21_X1 U9033 ( .B1(n9718), .B2(n7632), .A(n7380), .ZN(n7381) );
  OAI21_X1 U9034 ( .B1(n9720), .B2(n6638), .A(n7381), .ZN(P1_U3282) );
  NAND3_X1 U9035 ( .A1(n7383), .A2(n7382), .A3(n7387), .ZN(n7384) );
  NAND2_X1 U9036 ( .A1(n7367), .A2(n7384), .ZN(n7385) );
  AOI222_X1 U9037 ( .A1(n9406), .A2(n7385), .B1(n9128), .B2(n9401), .C1(n9126), 
        .C2(n9403), .ZN(n7468) );
  OAI21_X1 U9038 ( .B1(n7388), .B2(n7387), .A(n7386), .ZN(n7471) );
  INV_X1 U9039 ( .A(n7389), .ZN(n7392) );
  AOI21_X1 U9040 ( .B1(n7390), .B2(n7487), .A(n9707), .ZN(n7391) );
  NAND2_X1 U9041 ( .A1(n7392), .A2(n7391), .ZN(n7467) );
  NAND3_X1 U9042 ( .A1(n7394), .A2(n7393), .A3(n9682), .ZN(n7921) );
  AOI22_X1 U9043 ( .A1(n6638), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n7477), .B2(
        n9393), .ZN(n7396) );
  NAND2_X1 U9044 ( .A1(n9316), .A2(n7487), .ZN(n7395) );
  OAI211_X1 U9045 ( .C1(n7467), .C2(n7921), .A(n7396), .B(n7395), .ZN(n7397)
         );
  AOI21_X1 U9046 ( .B1(n7471), .B2(n7915), .A(n7397), .ZN(n7398) );
  OAI21_X1 U9047 ( .B1(n7468), .B2(n6638), .A(n7398), .ZN(P1_U3284) );
  XOR2_X1 U9048 ( .A(n7399), .B(n8180), .Z(n9798) );
  NOR2_X1 U9049 ( .A1(n8804), .A2(n8356), .ZN(n8762) );
  INV_X1 U9050 ( .A(n7400), .ZN(n7401) );
  AOI211_X1 U9051 ( .C1(n9794), .C2(n7401), .A(n9825), .B(n8814), .ZN(n9793)
         );
  OAI22_X1 U9052 ( .A1(n8821), .A2(n7403), .B1(n7668), .B2(n7402), .ZN(n7404)
         );
  AOI21_X1 U9053 ( .B1(n8762), .B2(n9793), .A(n7404), .ZN(n7409) );
  XNOR2_X1 U9054 ( .A(n7405), .B(n8180), .ZN(n7407) );
  AOI21_X1 U9055 ( .B1(n7407), .B2(n8813), .A(n7406), .ZN(n9796) );
  MUX2_X1 U9056 ( .A(n9796), .B(n6885), .S(n8804), .Z(n7408) );
  OAI211_X1 U9057 ( .C1(n9798), .C2(n8764), .A(n7409), .B(n7408), .ZN(P2_U3291) );
  INV_X1 U9058 ( .A(n9561), .ZN(n9578) );
  OAI21_X1 U9059 ( .B1(n7411), .B2(n9714), .A(n7410), .ZN(n7413) );
  AOI211_X1 U9060 ( .C1(n7414), .C2(n9578), .A(n7413), .B(n7412), .ZN(n7511)
         );
  NAND2_X1 U9061 ( .A1(n9725), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n7415) );
  OAI21_X1 U9062 ( .B1(n7511), .B2(n9725), .A(n7415), .ZN(P1_U3531) );
  NOR2_X1 U9063 ( .A1(n7422), .A2(n7416), .ZN(n7418) );
  NOR2_X1 U9064 ( .A1(n7418), .A2(n7417), .ZN(n7420) );
  NAND2_X1 U9065 ( .A1(n7588), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n7603) );
  OAI21_X1 U9066 ( .B1(n7588), .B2(P1_REG2_REG_16__SCAN_IN), .A(n7603), .ZN(
        n7419) );
  NOR2_X1 U9067 ( .A1(n7420), .A2(n7419), .ZN(n7601) );
  AOI211_X1 U9068 ( .C1(n7420), .C2(n7419), .A(n7601), .B(n9182), .ZN(n7432)
         );
  NOR2_X1 U9069 ( .A1(n7422), .A2(n7421), .ZN(n7424) );
  NOR2_X1 U9070 ( .A1(n7424), .A2(n7423), .ZN(n7427) );
  INV_X1 U9071 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9567) );
  NOR2_X1 U9072 ( .A1(n7588), .A2(n9567), .ZN(n7425) );
  AOI21_X1 U9073 ( .B1(n7588), .B2(n9567), .A(n7425), .ZN(n7426) );
  NOR2_X1 U9074 ( .A1(n7427), .A2(n7426), .ZN(n7589) );
  AOI211_X1 U9075 ( .C1(n7427), .C2(n7426), .A(n7589), .B(n9634), .ZN(n7431)
         );
  NAND2_X1 U9076 ( .A1(n9648), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n7428) );
  NAND2_X1 U9077 ( .A1(P1_U3084), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9024) );
  OAI211_X1 U9078 ( .C1(n7429), .C2(n9646), .A(n7428), .B(n9024), .ZN(n7430)
         );
  OR3_X1 U9079 ( .A1(n7432), .A2(n7431), .A3(n7430), .ZN(P1_U3257) );
  AOI21_X1 U9080 ( .B1(n7435), .B2(n7434), .A(n7433), .ZN(n7439) );
  XNOR2_X1 U9081 ( .A(n7437), .B(n7436), .ZN(n7438) );
  XNOR2_X1 U9082 ( .A(n7439), .B(n7438), .ZN(n7447) );
  AOI22_X1 U9083 ( .A1(n9094), .A2(n9127), .B1(n9112), .B2(n7440), .ZN(n7446)
         );
  NOR2_X1 U9084 ( .A1(n9092), .A2(n7441), .ZN(n7442) );
  AOI211_X1 U9085 ( .C1(n7444), .C2(n9106), .A(n7443), .B(n7442), .ZN(n7445)
         );
  OAI211_X1 U9086 ( .C1(n7447), .C2(n9115), .A(n7446), .B(n7445), .ZN(P1_U3237) );
  OR2_X1 U9087 ( .A1(n7772), .A2(n7456), .ZN(n8250) );
  NAND2_X1 U9088 ( .A1(n7772), .A2(n7456), .ZN(n8206) );
  INV_X1 U9089 ( .A(n8182), .ZN(n7449) );
  NAND2_X1 U9090 ( .A1(n7448), .A2(n8377), .ZN(n7657) );
  OR2_X1 U9091 ( .A1(n7772), .A2(n8376), .ZN(n7451) );
  AND2_X1 U9092 ( .A1(n7659), .A2(n7451), .ZN(n7453) );
  OR2_X1 U9093 ( .A1(n7634), .A2(n7655), .ZN(n8251) );
  NAND2_X1 U9094 ( .A1(n7634), .A2(n7655), .ZN(n8243) );
  NAND2_X1 U9095 ( .A1(n8251), .A2(n8243), .ZN(n8183) );
  AND2_X1 U9096 ( .A1(n8183), .A2(n7451), .ZN(n7452) );
  OAI21_X1 U9097 ( .B1(n7453), .B2(n8183), .A(n7636), .ZN(n9816) );
  INV_X1 U9098 ( .A(n8183), .ZN(n8203) );
  NAND2_X1 U9099 ( .A1(n7653), .A2(n8206), .ZN(n7455) );
  NAND2_X1 U9100 ( .A1(n7455), .A2(n8203), .ZN(n7640) );
  OAI21_X1 U9101 ( .B1(n8203), .B2(n7455), .A(n7640), .ZN(n7458) );
  OAI22_X1 U9102 ( .A1(n7456), .A2(n8756), .B1(n7637), .B2(n8754), .ZN(n7457)
         );
  AOI21_X1 U9103 ( .B1(n7458), .B2(n8813), .A(n7457), .ZN(n7459) );
  OAI21_X1 U9104 ( .B1(n9816), .B2(n8780), .A(n7459), .ZN(n9819) );
  NAND2_X1 U9105 ( .A1(n9819), .A2(n8830), .ZN(n7466) );
  INV_X1 U9106 ( .A(n7460), .ZN(n7461) );
  OAI22_X1 U9107 ( .A1(n8830), .A2(n6901), .B1(n7461), .B2(n7668), .ZN(n7464)
         );
  OR2_X1 U9108 ( .A1(n7665), .A2(n9817), .ZN(n7462) );
  NAND2_X1 U9109 ( .A1(n7804), .A2(n7462), .ZN(n9818) );
  NOR2_X1 U9110 ( .A1(n8582), .A2(n9818), .ZN(n7463) );
  AOI211_X1 U9111 ( .C1(n8827), .C2(n7634), .A(n7464), .B(n7463), .ZN(n7465)
         );
  OAI211_X1 U9112 ( .C1(n9816), .C2(n8790), .A(n7466), .B(n7465), .ZN(P2_U3286) );
  OAI211_X1 U9113 ( .C1(n7469), .C2(n9714), .A(n7468), .B(n7467), .ZN(n7470)
         );
  AOI21_X1 U9114 ( .B1(n9578), .B2(n7471), .A(n7470), .ZN(n7475) );
  NAND2_X1 U9115 ( .A1(n9725), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n7472) );
  OAI21_X1 U9116 ( .B1(n7475), .B2(n9725), .A(n7472), .ZN(P1_U3530) );
  INV_X1 U9117 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n7473) );
  OR2_X1 U9118 ( .A1(n9722), .A2(n7473), .ZN(n7474) );
  OAI21_X1 U9119 ( .B1(n7475), .B2(n9721), .A(n7474), .ZN(P1_U3475) );
  AOI21_X1 U9120 ( .B1(n9104), .B2(n9128), .A(n7476), .ZN(n7479) );
  NAND2_X1 U9121 ( .A1(n9106), .A2(n7477), .ZN(n7478) );
  OAI211_X1 U9122 ( .C1(n7480), .C2(n9109), .A(n7479), .B(n7478), .ZN(n7486)
         );
  INV_X1 U9123 ( .A(n7481), .ZN(n7482) );
  AOI211_X1 U9124 ( .C1(n7484), .C2(n7483), .A(n9115), .B(n7482), .ZN(n7485)
         );
  AOI211_X1 U9125 ( .C1(n7487), .C2(n9112), .A(n7486), .B(n7485), .ZN(n7488)
         );
  INV_X1 U9126 ( .A(n7488), .ZN(P1_U3211) );
  AOI22_X1 U9127 ( .A1(n9316), .A2(n6308), .B1(n9393), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n7489) );
  OAI21_X1 U9128 ( .B1(n9319), .B2(n7490), .A(n7489), .ZN(n7493) );
  MUX2_X1 U9129 ( .A(n7491), .B(P1_REG2_REG_2__SCAN_IN), .S(n6638), .Z(n7492)
         );
  AOI211_X1 U9130 ( .C1(n7632), .C2(n7494), .A(n7493), .B(n7492), .ZN(n7495)
         );
  INV_X1 U9131 ( .A(n7495), .ZN(P1_U3289) );
  XNOR2_X1 U9132 ( .A(n7612), .B(n7611), .ZN(n9544) );
  NAND2_X1 U9133 ( .A1(n7617), .A2(n7499), .ZN(n7500) );
  XNOR2_X1 U9134 ( .A(n7500), .B(n7611), .ZN(n7502) );
  AOI22_X1 U9135 ( .A1(n9401), .A2(n9125), .B1(n9123), .B2(n9403), .ZN(n7501)
         );
  OAI21_X1 U9136 ( .B1(n7502), .B2(n9329), .A(n7501), .ZN(n7503) );
  AOI21_X1 U9137 ( .B1(n9544), .B2(n7625), .A(n7503), .ZN(n9546) );
  NAND2_X1 U9138 ( .A1(n7505), .A2(n7685), .ZN(n7504) );
  NAND2_X1 U9139 ( .A1(n7504), .A2(n9559), .ZN(n7506) );
  OR2_X1 U9140 ( .A1(n7506), .A2(n7626), .ZN(n9541) );
  AOI22_X1 U9141 ( .A1(n6638), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n7688), .B2(
        n9393), .ZN(n7508) );
  NAND2_X1 U9142 ( .A1(n9316), .A2(n7685), .ZN(n7507) );
  OAI211_X1 U9143 ( .C1(n9541), .C2(n7921), .A(n7508), .B(n7507), .ZN(n7509)
         );
  AOI21_X1 U9144 ( .B1(n9544), .B2(n7632), .A(n7509), .ZN(n7510) );
  OAI21_X1 U9145 ( .B1(n9546), .B2(n6638), .A(n7510), .ZN(P1_U3281) );
  INV_X1 U9146 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n7513) );
  OR2_X1 U9147 ( .A1(n7511), .A2(n9721), .ZN(n7512) );
  OAI21_X1 U9148 ( .B1(n9722), .B2(n7513), .A(n7512), .ZN(P1_U3478) );
  XOR2_X1 U9149 ( .A(n7514), .B(n7515), .Z(n7522) );
  AND2_X1 U9150 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n9623) );
  AOI21_X1 U9151 ( .B1(n9104), .B2(n9126), .A(n9623), .ZN(n7518) );
  NAND2_X1 U9152 ( .A1(n9106), .A2(n7516), .ZN(n7517) );
  OAI211_X1 U9153 ( .C1(n7620), .C2(n9109), .A(n7518), .B(n7517), .ZN(n7519)
         );
  AOI21_X1 U9154 ( .B1(n7520), .B2(n9112), .A(n7519), .ZN(n7521) );
  OAI21_X1 U9155 ( .B1(n7522), .B2(n9115), .A(n7521), .ZN(P1_U3229) );
  INV_X1 U9156 ( .A(n7523), .ZN(n7528) );
  AOI21_X1 U9157 ( .B1(n7527), .B2(n7525), .A(n7524), .ZN(n7526) );
  AOI211_X1 U9158 ( .C1(n7528), .C2(n7527), .A(n5614), .B(n7526), .ZN(n7532)
         );
  INV_X1 U9159 ( .A(n8934), .ZN(n7807) );
  AOI22_X1 U9160 ( .A1(n5616), .A2(n7805), .B1(n8124), .B2(n8375), .ZN(n7530)
         );
  AOI22_X1 U9161 ( .A1(n8143), .A2(n8373), .B1(P2_REG3_REG_11__SCAN_IN), .B2(
        P2_U3152), .ZN(n7529) );
  OAI211_X1 U9162 ( .C1(n7807), .C2(n8146), .A(n7530), .B(n7529), .ZN(n7531)
         );
  OR2_X1 U9163 ( .A1(n7532), .A2(n7531), .ZN(P2_U3238) );
  NAND2_X1 U9164 ( .A1(n7534), .A2(n7533), .ZN(n7535) );
  XOR2_X1 U9165 ( .A(n7536), .B(n7535), .Z(n7545) );
  AOI21_X1 U9166 ( .B1(n9104), .B2(n9127), .A(n7537), .ZN(n7543) );
  NAND2_X1 U9167 ( .A1(n9112), .A2(n7538), .ZN(n7542) );
  NAND2_X1 U9168 ( .A1(n9106), .A2(n7539), .ZN(n7541) );
  NAND2_X1 U9169 ( .A1(n9094), .A2(n9125), .ZN(n7540) );
  NAND4_X1 U9170 ( .A1(n7543), .A2(n7542), .A3(n7541), .A4(n7540), .ZN(n7544)
         );
  AOI21_X1 U9171 ( .B1(n7545), .B2(n9087), .A(n7544), .ZN(n7546) );
  INV_X1 U9172 ( .A(n7546), .ZN(P1_U3219) );
  INV_X1 U9173 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10089) );
  NOR2_X1 U9174 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7547) );
  AOI21_X1 U9175 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n7547), .ZN(n9855) );
  NOR2_X1 U9176 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7548) );
  AOI21_X1 U9177 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n7548), .ZN(n9858) );
  NOR2_X1 U9178 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7549) );
  AOI21_X1 U9179 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n7549), .ZN(n9861) );
  NOR2_X1 U9180 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7550) );
  AOI21_X1 U9181 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n7550), .ZN(n9864) );
  NOR2_X1 U9182 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7551) );
  AOI21_X1 U9183 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n7551), .ZN(n9867) );
  NOR2_X1 U9184 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7557) );
  XNOR2_X1 U9185 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10097) );
  NAND2_X1 U9186 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7555) );
  XOR2_X1 U9187 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10095) );
  NAND2_X1 U9188 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n7553) );
  XOR2_X1 U9189 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(P1_ADDR_REG_2__SCAN_IN), .Z(
        n10092) );
  AOI21_X1 U9190 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9849) );
  INV_X1 U9191 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10021) );
  NAND3_X1 U9192 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n9851) );
  OAI21_X1 U9193 ( .B1(n9849), .B2(n10021), .A(n9851), .ZN(n10091) );
  NAND2_X1 U9194 ( .A1(n10092), .A2(n10091), .ZN(n7552) );
  NAND2_X1 U9195 ( .A1(n7553), .A2(n7552), .ZN(n10094) );
  NAND2_X1 U9196 ( .A1(n10095), .A2(n10094), .ZN(n7554) );
  NAND2_X1 U9197 ( .A1(n7555), .A2(n7554), .ZN(n10096) );
  NOR2_X1 U9198 ( .A1(n10097), .A2(n10096), .ZN(n7556) );
  NOR2_X1 U9199 ( .A1(n7557), .A2(n7556), .ZN(n7558) );
  NOR2_X1 U9200 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n7558), .ZN(n10085) );
  AND2_X1 U9201 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n7558), .ZN(n10084) );
  NOR2_X1 U9202 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10084), .ZN(n7559) );
  NOR2_X1 U9203 ( .A1(n10085), .A2(n7559), .ZN(n7560) );
  NAND2_X1 U9204 ( .A1(n7560), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n7562) );
  XOR2_X1 U9205 ( .A(n7560), .B(P1_ADDR_REG_6__SCAN_IN), .Z(n10083) );
  NAND2_X1 U9206 ( .A1(n10083), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n7561) );
  NAND2_X1 U9207 ( .A1(n7562), .A2(n7561), .ZN(n7563) );
  NAND2_X1 U9208 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n7563), .ZN(n7565) );
  XOR2_X1 U9209 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n7563), .Z(n10079) );
  NAND2_X1 U9210 ( .A1(n10079), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n7564) );
  NAND2_X1 U9211 ( .A1(n7565), .A2(n7564), .ZN(n7566) );
  NAND2_X1 U9212 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n7566), .ZN(n7569) );
  XNOR2_X1 U9213 ( .A(n7567), .B(n7566), .ZN(n10093) );
  NAND2_X1 U9214 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10093), .ZN(n7568) );
  NAND2_X1 U9215 ( .A1(n7569), .A2(n7568), .ZN(n7570) );
  AND2_X1 U9216 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n7570), .ZN(n7571) );
  XNOR2_X1 U9217 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n7570), .ZN(n10082) );
  INV_X1 U9218 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10081) );
  NOR2_X1 U9219 ( .A1(n10082), .A2(n10081), .ZN(n10080) );
  NAND2_X1 U9220 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n7572) );
  OAI21_X1 U9221 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n7572), .ZN(n9875) );
  AOI21_X1 U9222 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n9874), .ZN(n9873) );
  NAND2_X1 U9223 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n7573) );
  OAI21_X1 U9224 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n7573), .ZN(n9872) );
  NOR2_X1 U9225 ( .A1(n9873), .A2(n9872), .ZN(n9871) );
  AOI21_X1 U9226 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n9871), .ZN(n9870) );
  NOR2_X1 U9227 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7574) );
  AOI21_X1 U9228 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n7574), .ZN(n9869) );
  NAND2_X1 U9229 ( .A1(n9870), .A2(n9869), .ZN(n9868) );
  OAI21_X1 U9230 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n9868), .ZN(n9866) );
  NAND2_X1 U9231 ( .A1(n9867), .A2(n9866), .ZN(n9865) );
  OAI21_X1 U9232 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n9865), .ZN(n9863) );
  NAND2_X1 U9233 ( .A1(n9864), .A2(n9863), .ZN(n9862) );
  OAI21_X1 U9234 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n9862), .ZN(n9860) );
  NAND2_X1 U9235 ( .A1(n9861), .A2(n9860), .ZN(n9859) );
  OAI21_X1 U9236 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n9859), .ZN(n9857) );
  NAND2_X1 U9237 ( .A1(n9858), .A2(n9857), .ZN(n9856) );
  OAI21_X1 U9238 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n9856), .ZN(n9854) );
  NAND2_X1 U9239 ( .A1(n9855), .A2(n9854), .ZN(n9853) );
  OAI21_X1 U9240 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n9853), .ZN(n10088) );
  NOR2_X1 U9241 ( .A1(n10089), .A2(n10088), .ZN(n7575) );
  NAND2_X1 U9242 ( .A1(n10089), .A2(n10088), .ZN(n10087) );
  OAI21_X1 U9243 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n7575), .A(n10087), .ZN(
        n7579) );
  NOR2_X1 U9244 ( .A1(n7577), .A2(n7576), .ZN(n7578) );
  XNOR2_X1 U9245 ( .A(n7579), .B(n7578), .ZN(ADD_1071_U4) );
  NAND2_X1 U9246 ( .A1(n7581), .A2(n7580), .ZN(n7583) );
  XOR2_X1 U9247 ( .A(n7583), .B(n7582), .Z(n7587) );
  INV_X1 U9248 ( .A(n8372), .ZN(n7693) );
  AOI22_X1 U9249 ( .A1(n5616), .A2(n7647), .B1(n8124), .B2(n8374), .ZN(n7584)
         );
  NAND2_X1 U9250 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3152), .ZN(n8481) );
  OAI211_X1 U9251 ( .C1(n7693), .C2(n8159), .A(n7584), .B(n8481), .ZN(n7585)
         );
  AOI21_X1 U9252 ( .B1(n7691), .B2(n8166), .A(n7585), .ZN(n7586) );
  OAI21_X1 U9253 ( .B1(n7587), .B2(n5614), .A(n7586), .ZN(P2_U3226) );
  XNOR2_X1 U9254 ( .A(n9175), .B(P1_REG1_REG_18__SCAN_IN), .ZN(n7596) );
  NAND2_X1 U9255 ( .A1(n7588), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n7591) );
  INV_X1 U9256 ( .A(n7589), .ZN(n7590) );
  NAND2_X1 U9257 ( .A1(n7591), .A2(n7590), .ZN(n9169) );
  INV_X1 U9258 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n7592) );
  XNOR2_X1 U9259 ( .A(n9161), .B(n7592), .ZN(n9170) );
  NAND2_X1 U9260 ( .A1(n9169), .A2(n9170), .ZN(n9168) );
  NAND2_X1 U9261 ( .A1(n9161), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n7593) );
  NAND2_X1 U9262 ( .A1(n9168), .A2(n7593), .ZN(n7595) );
  OR2_X1 U9263 ( .A1(n7595), .A2(n7596), .ZN(n9177) );
  INV_X1 U9264 ( .A(n9177), .ZN(n7594) );
  AOI21_X1 U9265 ( .B1(n7596), .B2(n7595), .A(n7594), .ZN(n7610) );
  INV_X1 U9266 ( .A(n9175), .ZN(n7598) );
  NAND2_X1 U9267 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_U3084), .ZN(n7597) );
  OAI21_X1 U9268 ( .B1(n9646), .B2(n7598), .A(n7597), .ZN(n7599) );
  AOI21_X1 U9269 ( .B1(n9648), .B2(P1_ADDR_REG_18__SCAN_IN), .A(n7599), .ZN(
        n7609) );
  OR2_X1 U9270 ( .A1(n9175), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n7600) );
  NAND2_X1 U9271 ( .A1(n9175), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9179) );
  AND2_X1 U9272 ( .A1(n7600), .A2(n9179), .ZN(n7607) );
  INV_X1 U9273 ( .A(n7601), .ZN(n7602) );
  NAND2_X1 U9274 ( .A1(n7603), .A2(n7602), .ZN(n9166) );
  INV_X1 U9275 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n7604) );
  XNOR2_X1 U9276 ( .A(n9161), .B(n7604), .ZN(n9167) );
  NAND2_X1 U9277 ( .A1(n9166), .A2(n9167), .ZN(n9165) );
  NAND2_X1 U9278 ( .A1(n9161), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n7605) );
  NAND2_X1 U9279 ( .A1(n9165), .A2(n7605), .ZN(n7606) );
  NAND2_X1 U9280 ( .A1(n7606), .A2(n7607), .ZN(n9180) );
  OAI211_X1 U9281 ( .C1(n7607), .C2(n7606), .A(n9673), .B(n9180), .ZN(n7608)
         );
  OAI211_X1 U9282 ( .C1(n7610), .C2(n9634), .A(n7609), .B(n7608), .ZN(P1_U3259) );
  NAND2_X1 U9283 ( .A1(n7612), .A2(n7611), .ZN(n7614) );
  INV_X1 U9284 ( .A(n7620), .ZN(n9124) );
  OR2_X1 U9285 ( .A1(n7685), .A2(n9124), .ZN(n7613) );
  NAND2_X1 U9286 ( .A1(n7614), .A2(n7613), .ZN(n7755) );
  INV_X1 U9287 ( .A(n7619), .ZN(n7615) );
  XNOR2_X1 U9288 ( .A(n7755), .B(n7615), .ZN(n9584) );
  XNOR2_X1 U9289 ( .A(n7759), .B(n7619), .ZN(n7623) );
  OAI22_X1 U9290 ( .A1(n7620), .A2(n9331), .B1(n7787), .B2(n9333), .ZN(n7621)
         );
  INV_X1 U9291 ( .A(n7621), .ZN(n7622) );
  OAI21_X1 U9292 ( .B1(n7623), .B2(n9329), .A(n7622), .ZN(n7624) );
  AOI21_X1 U9293 ( .B1(n9584), .B2(n7625), .A(n7624), .ZN(n9586) );
  INV_X1 U9294 ( .A(n7629), .ZN(n9582) );
  NAND2_X1 U9295 ( .A1(n7626), .A2(n9582), .ZN(n7764) );
  OAI211_X1 U9296 ( .C1(n7626), .C2(n9582), .A(n9559), .B(n7764), .ZN(n9581)
         );
  INV_X1 U9297 ( .A(n7752), .ZN(n7627) );
  OAI22_X1 U9298 ( .A1(n9321), .A2(n9890), .B1(n7627), .B2(n9692), .ZN(n7628)
         );
  AOI21_X1 U9299 ( .B1(n7629), .B2(n9316), .A(n7628), .ZN(n7630) );
  OAI21_X1 U9300 ( .B1(n9581), .B2(n7883), .A(n7630), .ZN(n7631) );
  AOI21_X1 U9301 ( .B1(n9584), .B2(n7632), .A(n7631), .ZN(n7633) );
  OAI21_X1 U9302 ( .B1(n9586), .B2(n6638), .A(n7633), .ZN(P1_U3280) );
  NAND2_X1 U9303 ( .A1(n7634), .A2(n8375), .ZN(n7635) );
  OR2_X1 U9304 ( .A1(n8934), .A2(n7637), .ZN(n8259) );
  NAND2_X1 U9305 ( .A1(n8934), .A2(n7637), .ZN(n8244) );
  NAND2_X1 U9306 ( .A1(n8259), .A2(n8244), .ZN(n8184) );
  NAND2_X1 U9307 ( .A1(n7803), .A2(n8184), .ZN(n7639) );
  NAND2_X1 U9308 ( .A1(n8934), .A2(n8374), .ZN(n7638) );
  INV_X1 U9309 ( .A(n8373), .ZN(n7716) );
  OR2_X1 U9310 ( .A1(n7691), .A2(n7716), .ZN(n8263) );
  NAND2_X1 U9311 ( .A1(n7691), .A2(n7716), .ZN(n8261) );
  XNOR2_X1 U9312 ( .A(n7692), .B(n8187), .ZN(n9830) );
  INV_X1 U9313 ( .A(n9830), .ZN(n7652) );
  NAND2_X1 U9314 ( .A1(n7696), .A2(n8244), .ZN(n7641) );
  XNOR2_X1 U9315 ( .A(n7641), .B(n8187), .ZN(n7642) );
  NAND2_X1 U9316 ( .A1(n7642), .A2(n8813), .ZN(n7644) );
  AOI22_X1 U9317 ( .A1(n9743), .A2(n8374), .B1(n8372), .B2(n9744), .ZN(n7643)
         );
  NAND2_X1 U9318 ( .A1(n7644), .A2(n7643), .ZN(n9827) );
  INV_X1 U9319 ( .A(n7735), .ZN(n7646) );
  OAI21_X1 U9320 ( .B1(n4534), .B2(n4536), .A(n7646), .ZN(n9826) );
  AOI22_X1 U9321 ( .A1(n8804), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n7647), .B2(
        n9747), .ZN(n7649) );
  NAND2_X1 U9322 ( .A1(n8827), .A2(n7691), .ZN(n7648) );
  OAI211_X1 U9323 ( .C1(n9826), .C2(n8582), .A(n7649), .B(n7648), .ZN(n7650)
         );
  AOI21_X1 U9324 ( .B1(n9827), .B2(n8830), .A(n7650), .ZN(n7651) );
  OAI21_X1 U9325 ( .B1(n7652), .B2(n8764), .A(n7651), .ZN(P2_U3284) );
  OAI21_X1 U9326 ( .B1(n8182), .B2(n7654), .A(n7653), .ZN(n7664) );
  OAI22_X1 U9327 ( .A1(n7656), .A2(n8756), .B1(n7655), .B2(n8754), .ZN(n7663)
         );
  NAND2_X1 U9328 ( .A1(n7658), .A2(n7657), .ZN(n7661) );
  INV_X1 U9329 ( .A(n7659), .ZN(n7660) );
  AOI21_X1 U9330 ( .B1(n8182), .B2(n7661), .A(n7660), .ZN(n7776) );
  NOR2_X1 U9331 ( .A1(n7776), .A2(n8780), .ZN(n7662) );
  AOI211_X1 U9332 ( .C1(n8813), .C2(n7664), .A(n7663), .B(n7662), .ZN(n7775)
         );
  INV_X1 U9333 ( .A(n7776), .ZN(n7674) );
  INV_X1 U9334 ( .A(n8790), .ZN(n7743) );
  AOI21_X1 U9335 ( .B1(n7772), .B2(n7666), .A(n7665), .ZN(n7773) );
  INV_X1 U9336 ( .A(n7667), .ZN(n7669) );
  OAI22_X1 U9337 ( .A1(n8830), .A2(n6881), .B1(n7669), .B2(n7668), .ZN(n7670)
         );
  AOI21_X1 U9338 ( .B1(n7773), .B2(n7043), .A(n7670), .ZN(n7671) );
  OAI21_X1 U9339 ( .B1(n7672), .B2(n8821), .A(n7671), .ZN(n7673) );
  AOI21_X1 U9340 ( .B1(n7674), .B2(n7743), .A(n7673), .ZN(n7675) );
  OAI21_X1 U9341 ( .B1(n7775), .B2(n8804), .A(n7675), .ZN(P2_U3287) );
  INV_X1 U9342 ( .A(n7676), .ZN(n7988) );
  OAI222_X1 U9343 ( .A1(P1_U3084), .A2(n6241), .B1(n9508), .B2(n7988), .C1(
        n10076), .C2(n9510), .ZN(P1_U3331) );
  INV_X1 U9344 ( .A(n7677), .ZN(n7681) );
  NAND2_X1 U9345 ( .A1(n9506), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n7679) );
  OAI211_X1 U9346 ( .C1(n7681), .C2(n9508), .A(n7679), .B(n7678), .ZN(P1_U3330) );
  NAND2_X1 U9347 ( .A1(n8969), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n7680) );
  OAI211_X1 U9348 ( .C1(n7681), .C2(n8967), .A(n7680), .B(n8368), .ZN(P2_U3335) );
  XOR2_X1 U9349 ( .A(n7682), .B(n7683), .Z(n7690) );
  NAND2_X1 U9350 ( .A1(n9104), .A2(n9125), .ZN(n7684) );
  NAND2_X1 U9351 ( .A1(P1_U3084), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n9641) );
  OAI211_X1 U9352 ( .C1(n7763), .C2(n9109), .A(n7684), .B(n9641), .ZN(n7687)
         );
  INV_X1 U9353 ( .A(n7685), .ZN(n9542) );
  NOR2_X1 U9354 ( .A1(n9542), .A2(n9097), .ZN(n7686) );
  AOI211_X1 U9355 ( .C1(n7688), .C2(n9106), .A(n7687), .B(n7686), .ZN(n7689)
         );
  OAI21_X1 U9356 ( .B1(n7690), .B2(n9115), .A(n7689), .ZN(P1_U3215) );
  INV_X1 U9357 ( .A(n7722), .ZN(n7694) );
  OR2_X1 U9358 ( .A1(n7739), .A2(n7693), .ZN(n8267) );
  NAND2_X1 U9359 ( .A1(n7739), .A2(n7693), .ZN(n8266) );
  NAND2_X1 U9360 ( .A1(n7739), .A2(n8372), .ZN(n7695) );
  INV_X1 U9361 ( .A(n8802), .ZN(n8161) );
  NAND2_X1 U9362 ( .A1(n8925), .A2(n8161), .ZN(n8273) );
  INV_X1 U9363 ( .A(n8269), .ZN(n7699) );
  XNOR2_X1 U9364 ( .A(n7998), .B(n7699), .ZN(n8927) );
  AND2_X1 U9365 ( .A1(n8261), .A2(n8244), .ZN(n8262) );
  INV_X1 U9366 ( .A(n8188), .ZN(n8270) );
  INV_X1 U9367 ( .A(n8263), .ZN(n8260) );
  NOR2_X1 U9368 ( .A1(n8270), .A2(n8260), .ZN(n7697) );
  INV_X1 U9369 ( .A(n8266), .ZN(n7698) );
  NOR2_X1 U9370 ( .A1(n7699), .A2(n7698), .ZN(n7700) );
  NAND2_X1 U9371 ( .A1(n8023), .A2(n8813), .ZN(n7703) );
  AOI21_X1 U9372 ( .B1(n7726), .B2(n8266), .A(n8269), .ZN(n7702) );
  AOI22_X1 U9373 ( .A1(n9744), .A2(n8773), .B1(n8372), .B2(n9743), .ZN(n7701)
         );
  OAI21_X1 U9374 ( .B1(n7703), .B2(n7702), .A(n7701), .ZN(n8923) );
  INV_X1 U9375 ( .A(n8925), .ZN(n7710) );
  INV_X1 U9376 ( .A(n7739), .ZN(n8928) );
  INV_X1 U9377 ( .A(n7737), .ZN(n7705) );
  INV_X1 U9378 ( .A(n8796), .ZN(n7704) );
  AOI211_X1 U9379 ( .C1(n8925), .C2(n7705), .A(n9825), .B(n7704), .ZN(n8924)
         );
  INV_X1 U9380 ( .A(n7706), .ZN(n7707) );
  NAND2_X1 U9381 ( .A1(n8924), .A2(n7707), .ZN(n7709) );
  AOI22_X1 U9382 ( .A1(n8804), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n7817), .B2(
        n9747), .ZN(n7708) );
  OAI211_X1 U9383 ( .C1(n7710), .C2(n8821), .A(n7709), .B(n7708), .ZN(n7711)
         );
  AOI21_X1 U9384 ( .B1(n8923), .B2(n8830), .A(n7711), .ZN(n7712) );
  OAI21_X1 U9385 ( .B1(n8927), .B2(n8764), .A(n7712), .ZN(P2_U3282) );
  OAI211_X1 U9386 ( .C1(n7715), .C2(n7714), .A(n7713), .B(n4315), .ZN(n7720)
         );
  NOR2_X1 U9387 ( .A1(n8160), .A2(n7716), .ZN(n7718) );
  OAI22_X1 U9388 ( .A1(n8159), .A2(n8161), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7167), .ZN(n7717) );
  AOI211_X1 U9389 ( .C1(n5616), .C2(n7738), .A(n7718), .B(n7717), .ZN(n7719)
         );
  OAI211_X1 U9390 ( .C1(n8928), .C2(n8146), .A(n7720), .B(n7719), .ZN(P2_U3236) );
  NAND2_X1 U9391 ( .A1(n7722), .A2(n8188), .ZN(n7723) );
  NAND2_X1 U9392 ( .A1(n7721), .A2(n7723), .ZN(n7734) );
  OR2_X1 U9393 ( .A1(n7734), .A2(n8780), .ZN(n7733) );
  NAND2_X1 U9394 ( .A1(n7724), .A2(n8263), .ZN(n7725) );
  NAND2_X1 U9395 ( .A1(n7725), .A2(n8270), .ZN(n7727) );
  NAND2_X1 U9396 ( .A1(n7727), .A2(n7726), .ZN(n7731) );
  NAND2_X1 U9397 ( .A1(n8802), .A2(n9744), .ZN(n7729) );
  NAND2_X1 U9398 ( .A1(n8373), .A2(n9743), .ZN(n7728) );
  NAND2_X1 U9399 ( .A1(n7729), .A2(n7728), .ZN(n7730) );
  AOI21_X1 U9400 ( .B1(n7731), .B2(n8813), .A(n7730), .ZN(n7732) );
  INV_X1 U9401 ( .A(n7734), .ZN(n8931) );
  NOR2_X1 U9402 ( .A1(n7735), .A2(n8928), .ZN(n7736) );
  OR2_X1 U9403 ( .A1(n7737), .A2(n7736), .ZN(n8929) );
  AOI22_X1 U9404 ( .A1(n8804), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n7738), .B2(
        n9747), .ZN(n7741) );
  NAND2_X1 U9405 ( .A1(n8827), .A2(n7739), .ZN(n7740) );
  OAI211_X1 U9406 ( .C1(n8929), .C2(n8582), .A(n7741), .B(n7740), .ZN(n7742)
         );
  AOI21_X1 U9407 ( .B1(n8931), .B2(n7743), .A(n7742), .ZN(n7744) );
  OAI21_X1 U9408 ( .B1(n8933), .B2(n8804), .A(n7744), .ZN(P2_U3283) );
  AOI21_X1 U9409 ( .B1(n7745), .B2(n7746), .A(n9115), .ZN(n7748) );
  NAND2_X1 U9410 ( .A1(n7748), .A2(n7747), .ZN(n7754) );
  NAND2_X1 U9411 ( .A1(P1_U3084), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n9660) );
  INV_X1 U9412 ( .A(n9660), .ZN(n7749) );
  AOI21_X1 U9413 ( .B1(n9104), .B2(n9124), .A(n7749), .ZN(n7750) );
  OAI21_X1 U9414 ( .B1(n7787), .B2(n9109), .A(n7750), .ZN(n7751) );
  AOI21_X1 U9415 ( .B1(n7752), .B2(n9106), .A(n7751), .ZN(n7753) );
  OAI211_X1 U9416 ( .C1(n9582), .C2(n9097), .A(n7754), .B(n7753), .ZN(P1_U3234) );
  XNOR2_X1 U9417 ( .A(n7786), .B(n7785), .ZN(n9485) );
  NAND2_X1 U9418 ( .A1(n7779), .A2(n7760), .ZN(n7761) );
  XOR2_X1 U9419 ( .A(n7785), .B(n7761), .Z(n7762) );
  OAI222_X1 U9420 ( .A1(n9333), .A2(n7852), .B1(n9331), .B2(n7763), .C1(n9329), 
        .C2(n7762), .ZN(n9480) );
  INV_X1 U9421 ( .A(n9482), .ZN(n7857) );
  INV_X1 U9422 ( .A(n7792), .ZN(n7793) );
  AOI211_X1 U9423 ( .C1(n9482), .C2(n7764), .A(n9707), .B(n7793), .ZN(n9481)
         );
  INV_X1 U9424 ( .A(n7921), .ZN(n7846) );
  NAND2_X1 U9425 ( .A1(n9481), .A2(n7846), .ZN(n7766) );
  AOI22_X1 U9426 ( .A1(n6638), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n7854), .B2(
        n9393), .ZN(n7765) );
  OAI211_X1 U9427 ( .C1(n7857), .C2(n9396), .A(n7766), .B(n7765), .ZN(n7767)
         );
  AOI21_X1 U9428 ( .B1(n9480), .B2(n9688), .A(n7767), .ZN(n7768) );
  OAI21_X1 U9429 ( .B1(n9411), .B2(n9485), .A(n7768), .ZN(P1_U3279) );
  INV_X1 U9430 ( .A(n7769), .ZN(n7801) );
  NAND2_X1 U9431 ( .A1(n8969), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n7770) );
  OAI211_X1 U9432 ( .C1(n7801), .C2(n8967), .A(n7771), .B(n7770), .ZN(P2_U3334) );
  AOI22_X1 U9433 ( .A1(n7773), .A2(n9803), .B1(n9802), .B2(n7772), .ZN(n7774)
         );
  OAI211_X1 U9434 ( .C1(n7776), .C2(n9809), .A(n7775), .B(n7774), .ZN(n7798)
         );
  NAND2_X1 U9435 ( .A1(n7798), .A2(n9848), .ZN(n7777) );
  OAI21_X1 U9436 ( .B1(n9848), .B2(n6873), .A(n7777), .ZN(P2_U3529) );
  NAND2_X1 U9437 ( .A1(n7779), .A2(n7778), .ZN(n7781) );
  XNOR2_X1 U9438 ( .A(n7837), .B(n7836), .ZN(n7784) );
  NAND2_X1 U9439 ( .A1(n9120), .A2(n9403), .ZN(n7782) );
  OAI21_X1 U9440 ( .B1(n7787), .B2(n9331), .A(n7782), .ZN(n7783) );
  AOI21_X1 U9441 ( .B1(n7784), .B2(n9406), .A(n7783), .ZN(n9575) );
  INV_X1 U9442 ( .A(n7787), .ZN(n9122) );
  NAND2_X1 U9443 ( .A1(n9482), .A2(n9122), .ZN(n7788) );
  NAND2_X1 U9444 ( .A1(n7789), .A2(n7788), .ZN(n7831) );
  XNOR2_X1 U9445 ( .A(n7831), .B(n7836), .ZN(n9579) );
  NAND2_X1 U9446 ( .A1(n9579), .A2(n7915), .ZN(n7797) );
  INV_X1 U9447 ( .A(n7863), .ZN(n7790) );
  OAI22_X1 U9448 ( .A1(n9321), .A2(n7791), .B1(n7790), .B2(n9692), .ZN(n7795)
         );
  INV_X1 U9449 ( .A(n7868), .ZN(n9576) );
  NOR2_X2 U9450 ( .A1(n7792), .A2(n7868), .ZN(n7832) );
  INV_X1 U9451 ( .A(n7832), .ZN(n7833) );
  OAI211_X1 U9452 ( .C1(n9576), .C2(n7793), .A(n7833), .B(n9559), .ZN(n9574)
         );
  NOR2_X1 U9453 ( .A1(n9574), .A2(n7883), .ZN(n7794) );
  AOI211_X1 U9454 ( .C1(n9316), .C2(n7868), .A(n7795), .B(n7794), .ZN(n7796)
         );
  OAI211_X1 U9455 ( .C1(n6638), .C2(n9575), .A(n7797), .B(n7796), .ZN(P1_U3278) );
  INV_X1 U9456 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n7800) );
  NAND2_X1 U9457 ( .A1(n7798), .A2(n9833), .ZN(n7799) );
  OAI21_X1 U9458 ( .B1(n9833), .B2(n7800), .A(n7799), .ZN(P2_U3478) );
  OAI222_X1 U9459 ( .A1(n7802), .A2(P1_U3084), .B1(n9508), .B2(n7801), .C1(
        n10055), .C2(n9510), .ZN(P1_U3329) );
  XNOR2_X1 U9460 ( .A(n7803), .B(n8184), .ZN(n8938) );
  AOI21_X1 U9461 ( .B1(n8934), .B2(n7804), .A(n4536), .ZN(n8935) );
  AOI22_X1 U9462 ( .A1(n8804), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n7805), .B2(
        n9747), .ZN(n7806) );
  OAI21_X1 U9463 ( .B1(n7807), .B2(n8821), .A(n7806), .ZN(n7811) );
  XOR2_X1 U9464 ( .A(n8184), .B(n7808), .Z(n7809) );
  AOI222_X1 U9465 ( .A1(n8813), .A2(n7809), .B1(n8373), .B2(n9744), .C1(n8375), 
        .C2(n9743), .ZN(n8937) );
  NOR2_X1 U9466 ( .A1(n8937), .A2(n8804), .ZN(n7810) );
  AOI211_X1 U9467 ( .C1(n8935), .C2(n7043), .A(n7811), .B(n7810), .ZN(n7812)
         );
  OAI21_X1 U9468 ( .B1(n8764), .B2(n8938), .A(n7812), .ZN(P2_U3285) );
  INV_X1 U9469 ( .A(n7813), .ZN(n7814) );
  AOI21_X1 U9470 ( .B1(n7816), .B2(n7815), .A(n7814), .ZN(n7822) );
  INV_X1 U9471 ( .A(n8773), .ZN(n8001) );
  AOI22_X1 U9472 ( .A1(n5616), .A2(n7817), .B1(n8124), .B2(n8372), .ZN(n7819)
         );
  OAI211_X1 U9473 ( .C1(n8001), .C2(n8159), .A(n7819), .B(n7818), .ZN(n7820)
         );
  AOI21_X1 U9474 ( .B1(n8925), .B2(n8166), .A(n7820), .ZN(n7821) );
  OAI21_X1 U9475 ( .B1(n7822), .B2(n5614), .A(n7821), .ZN(P2_U3217) );
  INV_X1 U9476 ( .A(n7823), .ZN(n7827) );
  AOI22_X1 U9477 ( .A1(n7824), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_25__SCAN_IN), .B2(n8969), .ZN(n7825) );
  OAI21_X1 U9478 ( .B1(n7827), .B2(n8967), .A(n7825), .ZN(P2_U3333) );
  OAI222_X1 U9479 ( .A1(P1_U3084), .A2(n7828), .B1(n9508), .B2(n7827), .C1(
        n7826), .C2(n9510), .ZN(P1_U3328) );
  AND2_X1 U9480 ( .A1(n7868), .A2(n9121), .ZN(n7830) );
  XOR2_X1 U9481 ( .A(n7840), .B(n7879), .Z(n9479) );
  INV_X1 U9482 ( .A(n9476), .ZN(n7835) );
  AOI211_X1 U9483 ( .C1(n9476), .C2(n7833), .A(n9707), .B(n7882), .ZN(n9475)
         );
  AOI22_X1 U9484 ( .A1(n6638), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n7899), .B2(
        n9393), .ZN(n7834) );
  OAI21_X1 U9485 ( .B1(n7835), .B2(n9396), .A(n7834), .ZN(n7845) );
  NAND2_X1 U9486 ( .A1(n7837), .A2(n7836), .ZN(n7839) );
  NAND2_X1 U9487 ( .A1(n7839), .A2(n7838), .ZN(n7841) );
  AOI21_X1 U9488 ( .B1(n7841), .B2(n7840), .A(n9329), .ZN(n7843) );
  OAI22_X1 U9489 ( .A1(n7852), .A2(n9331), .B1(n7902), .B2(n9333), .ZN(n7842)
         );
  AOI21_X1 U9490 ( .B1(n7843), .B2(n7872), .A(n7842), .ZN(n9478) );
  NOR2_X1 U9491 ( .A1(n9478), .A2(n6638), .ZN(n7844) );
  AOI211_X1 U9492 ( .C1(n7846), .C2(n9475), .A(n7845), .B(n7844), .ZN(n7847)
         );
  OAI21_X1 U9493 ( .B1(n9479), .B2(n9411), .A(n7847), .ZN(P1_U3277) );
  OAI21_X1 U9494 ( .B1(n7849), .B2(n4384), .A(n7848), .ZN(n7850) );
  NAND2_X1 U9495 ( .A1(n7850), .A2(n9087), .ZN(n7856) );
  AOI22_X1 U9496 ( .A1(n9104), .A2(n9123), .B1(P1_REG3_REG_12__SCAN_IN), .B2(
        P1_U3084), .ZN(n7851) );
  OAI21_X1 U9497 ( .B1(n7852), .B2(n9109), .A(n7851), .ZN(n7853) );
  AOI21_X1 U9498 ( .B1(n7854), .B2(n9106), .A(n7853), .ZN(n7855) );
  OAI211_X1 U9499 ( .C1(n7857), .C2(n9097), .A(n7856), .B(n7855), .ZN(P1_U3222) );
  XNOR2_X1 U9500 ( .A(n7859), .B(n7858), .ZN(n7860) );
  XNOR2_X1 U9501 ( .A(n7861), .B(n7860), .ZN(n7870) );
  AOI21_X1 U9502 ( .B1(n9104), .B2(n9122), .A(n7862), .ZN(n7865) );
  NAND2_X1 U9503 ( .A1(n9106), .A2(n7863), .ZN(n7864) );
  OAI211_X1 U9504 ( .C1(n7866), .C2(n9109), .A(n7865), .B(n7864), .ZN(n7867)
         );
  AOI21_X1 U9505 ( .B1(n7868), .B2(n9112), .A(n7867), .ZN(n7869) );
  OAI21_X1 U9506 ( .B1(n7870), .B2(n9115), .A(n7869), .ZN(P1_U3232) );
  INV_X1 U9507 ( .A(n7880), .ZN(n7873) );
  XNOR2_X1 U9508 ( .A(n7907), .B(n7873), .ZN(n7876) );
  NAND2_X1 U9509 ( .A1(n9120), .A2(n9401), .ZN(n7874) );
  OAI21_X1 U9510 ( .B1(n9110), .B2(n9333), .A(n7874), .ZN(n7875) );
  AOI21_X1 U9511 ( .B1(n7876), .B2(n9406), .A(n7875), .ZN(n9569) );
  NOR2_X1 U9512 ( .A1(n9476), .A2(n9120), .ZN(n7878) );
  NAND2_X1 U9513 ( .A1(n9476), .A2(n9120), .ZN(n7877) );
  XNOR2_X1 U9514 ( .A(n7912), .B(n7880), .ZN(n9572) );
  NAND2_X1 U9515 ( .A1(n9572), .A2(n7915), .ZN(n7887) );
  INV_X1 U9516 ( .A(n9105), .ZN(n7881) );
  OAI22_X1 U9517 ( .A1(n9688), .A2(n9943), .B1(n7881), .B2(n9692), .ZN(n7885)
         );
  INV_X1 U9518 ( .A(n9113), .ZN(n9570) );
  OAI211_X1 U9519 ( .C1(n7882), .C2(n9570), .A(n9559), .B(n7919), .ZN(n9568)
         );
  NOR2_X1 U9520 ( .A1(n9568), .A2(n7883), .ZN(n7884) );
  AOI211_X1 U9521 ( .C1(n9316), .C2(n9113), .A(n7885), .B(n7884), .ZN(n7886)
         );
  OAI211_X1 U9522 ( .C1(n6638), .C2(n9569), .A(n7887), .B(n7886), .ZN(P1_U3276) );
  INV_X1 U9523 ( .A(n7888), .ZN(n7932) );
  OAI222_X1 U9524 ( .A1(P2_U3152), .A2(n7890), .B1(n8967), .B2(n7932), .C1(
        n7889), .C2(n7990), .ZN(P2_U3332) );
  INV_X1 U9525 ( .A(n7891), .ZN(n7927) );
  AOI21_X1 U9526 ( .B1(n9506), .B2(P2_DATAO_REG_27__SCAN_IN), .A(n7892), .ZN(
        n7893) );
  OAI21_X1 U9527 ( .B1(n7927), .B2(n9508), .A(n7893), .ZN(P1_U3326) );
  XNOR2_X1 U9528 ( .A(n7895), .B(n7894), .ZN(n7896) );
  XNOR2_X1 U9529 ( .A(n7897), .B(n7896), .ZN(n7905) );
  NOR2_X1 U9530 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7898), .ZN(n9662) );
  AOI21_X1 U9531 ( .B1(n9104), .B2(n9121), .A(n9662), .ZN(n7901) );
  NAND2_X1 U9532 ( .A1(n9106), .A2(n7899), .ZN(n7900) );
  OAI211_X1 U9533 ( .C1(n7902), .C2(n9109), .A(n7901), .B(n7900), .ZN(n7903)
         );
  AOI21_X1 U9534 ( .B1(n9476), .B2(n9112), .A(n7903), .ZN(n7904) );
  OAI21_X1 U9535 ( .B1(n7905), .B2(n9115), .A(n7904), .ZN(P1_U3213) );
  NAND2_X1 U9536 ( .A1(n7909), .A2(n7913), .ZN(n9398) );
  OAI21_X1 U9537 ( .B1(n7913), .B2(n7909), .A(n9398), .ZN(n7910) );
  AOI222_X1 U9538 ( .A1(n9406), .A2(n7910), .B1(n9384), .B2(n9403), .C1(n9119), 
        .C2(n9401), .ZN(n9564) );
  AND2_X1 U9539 ( .A1(n7914), .A2(n7913), .ZN(n9562) );
  INV_X1 U9540 ( .A(n9562), .ZN(n7916) );
  NAND3_X1 U9541 ( .A1(n7916), .A2(n7915), .A3(n7941), .ZN(n7925) );
  INV_X1 U9542 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n7918) );
  INV_X1 U9543 ( .A(n9029), .ZN(n7917) );
  OAI22_X1 U9544 ( .A1(n9688), .A2(n7918), .B1(n7917), .B2(n9692), .ZN(n7923)
         );
  INV_X1 U9545 ( .A(n7919), .ZN(n7920) );
  OAI211_X1 U9546 ( .C1(n7920), .C2(n4600), .A(n9559), .B(n9392), .ZN(n9563)
         );
  NOR2_X1 U9547 ( .A1(n9563), .A2(n7921), .ZN(n7922) );
  AOI211_X1 U9548 ( .C1(n9316), .C2(n7939), .A(n7923), .B(n7922), .ZN(n7924)
         );
  OAI211_X1 U9549 ( .C1(n6638), .C2(n9564), .A(n7925), .B(n7924), .ZN(P1_U3275) );
  INV_X1 U9550 ( .A(n7926), .ZN(n9512) );
  OAI222_X1 U9551 ( .A1(n8967), .A2(n9512), .B1(P2_U3152), .B2(n5620), .C1(
        n9988), .C2(n7990), .ZN(P2_U3330) );
  OAI222_X1 U9552 ( .A1(n7990), .A2(n7928), .B1(n8967), .B2(n7927), .C1(n8364), 
        .C2(P2_U3152), .ZN(P2_U3331) );
  INV_X1 U9553 ( .A(n8013), .ZN(n8972) );
  INV_X1 U9554 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n7929) );
  OAI222_X1 U9555 ( .A1(n9508), .A2(n8972), .B1(n7930), .B2(P1_U3084), .C1(
        n7929), .C2(n9510), .ZN(P1_U3324) );
  OAI222_X1 U9556 ( .A1(n7933), .A2(P1_U3084), .B1(n9508), .B2(n7932), .C1(
        n7931), .C2(n9510), .ZN(P1_U3327) );
  OAI222_X1 U9557 ( .A1(n7936), .A2(P1_U3084), .B1(n9508), .B2(n7935), .C1(
        n7934), .C2(n9510), .ZN(P1_U3333) );
  INV_X1 U9558 ( .A(n8172), .ZN(n8968) );
  OAI222_X1 U9559 ( .A1(n9510), .A2(n7938), .B1(n9508), .B2(n8968), .C1(
        P1_U3084), .C2(n7937), .ZN(P1_U3323) );
  INV_X1 U9560 ( .A(n9110), .ZN(n9402) );
  NAND2_X1 U9561 ( .A1(n7939), .A2(n9402), .ZN(n7940) );
  OR2_X1 U9562 ( .A1(n9470), .A2(n9384), .ZN(n7942) );
  NAND2_X1 U9563 ( .A1(n9389), .A2(n7942), .ZN(n7944) );
  NAND2_X1 U9564 ( .A1(n9470), .A2(n9384), .ZN(n7943) );
  INV_X1 U9565 ( .A(n9037), .ZN(n9404) );
  NAND2_X1 U9566 ( .A1(n9465), .A2(n9404), .ZN(n7945) );
  AND2_X1 U9567 ( .A1(n9460), .A2(n9383), .ZN(n7946) );
  NOR2_X1 U9568 ( .A1(n9455), .A2(n9369), .ZN(n7948) );
  NAND2_X1 U9569 ( .A1(n9455), .A2(n9369), .ZN(n7947) );
  NAND2_X1 U9570 ( .A1(n9325), .A2(n9324), .ZN(n7950) );
  INV_X1 U9571 ( .A(n9055), .ZN(n9352) );
  NAND2_X1 U9572 ( .A1(n9452), .A2(n9352), .ZN(n7949) );
  AND2_X1 U9573 ( .A1(n9317), .A2(n9118), .ZN(n7952) );
  OR2_X1 U9574 ( .A1(n9317), .A2(n9118), .ZN(n7951) );
  NOR2_X1 U9575 ( .A1(n9441), .A2(n9308), .ZN(n7954) );
  NAND2_X1 U9576 ( .A1(n9441), .A2(n9308), .ZN(n7953) );
  NAND2_X1 U9577 ( .A1(n9254), .A2(n9263), .ZN(n7956) );
  NAND2_X1 U9578 ( .A1(n7956), .A2(n7955), .ZN(n9238) );
  NOR2_X1 U9579 ( .A1(n9424), .A2(n9264), .ZN(n7958) );
  NAND2_X1 U9580 ( .A1(n9424), .A2(n9264), .ZN(n7957) );
  NAND2_X1 U9581 ( .A1(n9398), .A2(n7962), .ZN(n9380) );
  NAND2_X1 U9582 ( .A1(n9380), .A2(n7963), .ZN(n9366) );
  NAND2_X1 U9583 ( .A1(n9366), .A2(n9365), .ZN(n7965) );
  NAND2_X1 U9584 ( .A1(n7965), .A2(n7964), .ZN(n9368) );
  NAND2_X1 U9585 ( .A1(n9245), .A2(n7974), .ZN(n7976) );
  NOR2_X1 U9586 ( .A1(n7983), .A2(n7982), .ZN(n7984) );
  NOR2_X1 U9587 ( .A1(n9333), .A2(n7984), .ZN(n9194) );
  INV_X1 U9588 ( .A(n9460), .ZN(n9363) );
  NAND2_X1 U9589 ( .A1(n9375), .A2(n9363), .ZN(n9358) );
  OR2_X2 U9590 ( .A1(n9358), .A2(n9455), .ZN(n9344) );
  INV_X1 U9591 ( .A(n9317), .ZN(n9444) );
  INV_X1 U9592 ( .A(n9441), .ZN(n9298) );
  NOR2_X2 U9593 ( .A1(n9279), .A2(n9429), .ZN(n9255) );
  INV_X1 U9594 ( .A(n9424), .ZN(n9243) );
  AND2_X2 U9595 ( .A1(n9255), .A2(n9243), .ZN(n9239) );
  AOI22_X1 U9596 ( .A1(n7996), .A2(n9559), .B1(n9483), .B2(n7986), .ZN(n7987)
         );
  OAI211_X1 U9597 ( .C1(n7997), .C2(n9561), .A(n7994), .B(n7987), .ZN(n9487)
         );
  MUX2_X1 U9598 ( .A(n9487), .B(P1_REG1_REG_29__SCAN_IN), .S(n9725), .Z(
        P1_U3552) );
  OAI222_X1 U9599 ( .A1(n7990), .A2(n7989), .B1(n8967), .B2(n7988), .C1(n6820), 
        .C2(P2_U3152), .ZN(P2_U3336) );
  AOI22_X1 U9600 ( .A1(n7991), .A2(n9393), .B1(P1_REG2_REG_29__SCAN_IN), .B2(
        n6638), .ZN(n7992) );
  OAI21_X1 U9601 ( .B1(n7993), .B2(n9396), .A(n7992), .ZN(n7995) );
  INV_X1 U9602 ( .A(n8739), .ZN(n8026) );
  OR2_X1 U9603 ( .A1(n8925), .A2(n8802), .ZN(n7999) );
  NAND2_X1 U9604 ( .A1(n8000), .A2(n7999), .ZN(n8792) );
  NAND2_X1 U9605 ( .A1(n8918), .A2(n8001), .ZN(n8277) );
  NAND2_X1 U9606 ( .A1(n8278), .A2(n8277), .ZN(n8799) );
  OR2_X1 U9607 ( .A1(n8918), .A2(n8773), .ZN(n8002) );
  XNOR2_X1 U9608 ( .A(n8783), .B(n8801), .ZN(n8765) );
  INV_X1 U9609 ( .A(n8774), .ZN(n8283) );
  XNOR2_X1 U9610 ( .A(n8905), .B(n8283), .ZN(n8753) );
  NAND2_X1 U9611 ( .A1(n8750), .A2(n8283), .ZN(n8003) );
  NAND2_X1 U9612 ( .A1(n8899), .A2(n8371), .ZN(n8005) );
  INV_X1 U9613 ( .A(n8371), .ZN(n8755) );
  NAND2_X1 U9614 ( .A1(n8716), .A2(n8006), .ZN(n8007) );
  INV_X1 U9615 ( .A(n8698), .ZN(n8077) );
  NAND2_X1 U9616 ( .A1(n8889), .A2(n8077), .ZN(n8297) );
  NAND2_X1 U9617 ( .A1(n8301), .A2(n8297), .ZN(n8704) );
  NAND2_X1 U9618 ( .A1(n8884), .A2(n8711), .ZN(n8008) );
  INV_X1 U9619 ( .A(n8711), .ZN(n8681) );
  INV_X1 U9620 ( .A(n8884), .ZN(n8692) );
  INV_X1 U9621 ( .A(n8699), .ZN(n10075) );
  NAND2_X1 U9622 ( .A1(n8879), .A2(n10075), .ZN(n8306) );
  NAND2_X1 U9623 ( .A1(n8867), .A2(n8088), .ZN(n8312) );
  NAND2_X1 U9624 ( .A1(n8009), .A2(n8088), .ZN(n8010) );
  NAND2_X1 U9625 ( .A1(n8863), .A2(n8150), .ZN(n8315) );
  INV_X1 U9626 ( .A(n8863), .ZN(n8627) );
  NAND2_X1 U9627 ( .A1(n8858), .A2(n8087), .ZN(n8317) );
  NAND2_X1 U9628 ( .A1(n8852), .A2(n8149), .ZN(n8327) );
  INV_X1 U9629 ( .A(n8601), .ZN(n8048) );
  NAND2_X1 U9630 ( .A1(n8847), .A2(n8048), .ZN(n8329) );
  NAND2_X1 U9631 ( .A1(n8013), .A2(n8171), .ZN(n8016) );
  NAND2_X1 U9632 ( .A1(n8014), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n8015) );
  INV_X1 U9633 ( .A(n8590), .ZN(n8017) );
  NAND2_X1 U9634 ( .A1(n8842), .A2(n8017), .ZN(n8348) );
  INV_X1 U9635 ( .A(n8858), .ZN(n8612) );
  INV_X1 U9636 ( .A(n8905), .ZN(n8750) );
  INV_X1 U9637 ( .A(n8879), .ZN(n8674) );
  INV_X1 U9638 ( .A(n8873), .ZN(n8663) );
  AOI21_X1 U9639 ( .B1(n8842), .B2(n8584), .A(n8577), .ZN(n8843) );
  INV_X1 U9640 ( .A(n8842), .ZN(n8022) );
  INV_X1 U9641 ( .A(n8019), .ZN(n8020) );
  AOI22_X1 U9642 ( .A1(n8804), .A2(P2_REG2_REG_29__SCAN_IN), .B1(n8020), .B2(
        n9747), .ZN(n8021) );
  OAI21_X1 U9643 ( .B1(n8022), .B2(n8821), .A(n8021), .ZN(n8043) );
  INV_X1 U9644 ( .A(n8330), .ZN(n8034) );
  INV_X1 U9645 ( .A(n8799), .ZN(n8275) );
  INV_X1 U9646 ( .A(n8770), .ZN(n8024) );
  INV_X1 U9647 ( .A(n8765), .ZN(n8769) );
  INV_X1 U9648 ( .A(n8801), .ZN(n8757) );
  NAND2_X1 U9649 ( .A1(n8783), .A2(n8757), .ZN(n8285) );
  OR2_X1 U9650 ( .A1(n8899), .A2(n8755), .ZN(n8291) );
  NAND2_X1 U9651 ( .A1(n8899), .A2(n8755), .ZN(n8294) );
  NAND2_X1 U9652 ( .A1(n8291), .A2(n8294), .ZN(n8735) );
  NOR2_X1 U9653 ( .A1(n8905), .A2(n8283), .ZN(n8736) );
  NOR2_X1 U9654 ( .A1(n8735), .A2(n8736), .ZN(n8025) );
  NAND2_X1 U9655 ( .A1(n8737), .A2(n8294), .ZN(n8717) );
  OR2_X1 U9656 ( .A1(n8896), .A2(n8026), .ZN(n8299) );
  NAND2_X1 U9657 ( .A1(n8896), .A2(n8026), .ZN(n8295) );
  NAND2_X1 U9658 ( .A1(n8717), .A2(n8718), .ZN(n8027) );
  NAND2_X1 U9659 ( .A1(n8027), .A2(n8295), .ZN(n8710) );
  OR2_X1 U9660 ( .A1(n8884), .A2(n8681), .ZN(n8302) );
  NAND2_X1 U9661 ( .A1(n8884), .A2(n8681), .ZN(n8678) );
  NAND2_X1 U9662 ( .A1(n8302), .A2(n8678), .ZN(n8694) );
  INV_X1 U9663 ( .A(n8301), .ZN(n8695) );
  NOR2_X1 U9664 ( .A1(n8694), .A2(n8695), .ZN(n8029) );
  INV_X1 U9665 ( .A(n8678), .ZN(n8030) );
  NOR2_X1 U9666 ( .A1(n8667), .A2(n8030), .ZN(n8031) );
  INV_X1 U9667 ( .A(n8645), .ZN(n8682) );
  AND2_X1 U9668 ( .A1(n8873), .A2(n8682), .ZN(n8641) );
  NOR2_X1 U9669 ( .A1(n8640), .A2(n8641), .ZN(n8032) );
  NAND2_X1 U9670 ( .A1(n8643), .A2(n8311), .ZN(n8629) );
  INV_X1 U9671 ( .A(n8325), .ZN(n8331) );
  NAND2_X1 U9672 ( .A1(n4321), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8040) );
  NAND2_X1 U9673 ( .A1(n8036), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n8039) );
  NAND2_X1 U9674 ( .A1(n8037), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n8038) );
  NAND3_X1 U9675 ( .A1(n8040), .A2(n8039), .A3(n8038), .ZN(n8369) );
  INV_X1 U9676 ( .A(n8364), .ZN(n8041) );
  AOI21_X1 U9677 ( .B1(n8041), .B2(P2_B_REG_SCAN_IN), .A(n8754), .ZN(n8572) );
  NOR2_X1 U9678 ( .A1(n8845), .A2(n8804), .ZN(n8042) );
  AOI211_X1 U9679 ( .C1(n8843), .C2(n7043), .A(n8043), .B(n8042), .ZN(n8044)
         );
  OAI21_X1 U9680 ( .B1(n8846), .B2(n8764), .A(n8044), .ZN(P2_U3267) );
  XNOR2_X1 U9681 ( .A(n8045), .B(n8046), .ZN(n8053) );
  OAI22_X1 U9682 ( .A1(n8159), .A2(n8048), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8047), .ZN(n8051) );
  INV_X1 U9683 ( .A(n8597), .ZN(n8049) );
  OAI22_X1 U9684 ( .A1(n8163), .A2(n8049), .B1(n8087), .B2(n8160), .ZN(n8050)
         );
  AOI211_X1 U9685 ( .C1(n8852), .C2(n8166), .A(n8051), .B(n8050), .ZN(n8052)
         );
  OAI21_X1 U9686 ( .B1(n8053), .B2(n5614), .A(n8052), .ZN(P2_U3216) );
  INV_X1 U9687 ( .A(n8057), .ZN(n8054) );
  NOR2_X1 U9688 ( .A1(n8054), .A2(n8055), .ZN(n8112) );
  INV_X1 U9689 ( .A(n8055), .ZN(n8056) );
  OAI21_X1 U9690 ( .B1(n8057), .B2(n8056), .A(n4315), .ZN(n8062) );
  OAI22_X1 U9691 ( .A1(n8159), .A2(n8088), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8058), .ZN(n8060) );
  OAI22_X1 U9692 ( .A1(n8163), .A2(n8660), .B1(n10075), .B2(n8160), .ZN(n8059)
         );
  AOI211_X1 U9693 ( .C1(n8873), .C2(n8166), .A(n8060), .B(n8059), .ZN(n8061)
         );
  OAI21_X1 U9694 ( .B1(n8112), .B2(n8062), .A(n8061), .ZN(P2_U3218) );
  INV_X1 U9695 ( .A(n8063), .ZN(n8064) );
  AOI21_X1 U9696 ( .B1(n8066), .B2(n8065), .A(n8064), .ZN(n8072) );
  INV_X1 U9697 ( .A(n8067), .ZN(n8723) );
  AND2_X1 U9698 ( .A1(P2_U3152), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8571) );
  AOI22_X1 U9699 ( .A1(n8698), .A2(n9744), .B1(n9743), .B2(n8371), .ZN(n8719)
         );
  NOR2_X1 U9700 ( .A1(n8068), .A2(n8719), .ZN(n8069) );
  AOI211_X1 U9701 ( .C1(n5616), .C2(n8723), .A(n8571), .B(n8069), .ZN(n8071)
         );
  NAND2_X1 U9702 ( .A1(n8896), .A2(n8166), .ZN(n8070) );
  OAI211_X1 U9703 ( .C1(n8072), .C2(n5614), .A(n8071), .B(n8070), .ZN(P2_U3221) );
  OAI211_X1 U9704 ( .C1(n8075), .C2(n8074), .A(n8073), .B(n4315), .ZN(n8081)
         );
  OAI22_X1 U9705 ( .A1(n8159), .A2(n10075), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8076), .ZN(n8079) );
  OAI22_X1 U9706 ( .A1(n8163), .A2(n8689), .B1(n8077), .B2(n8160), .ZN(n8078)
         );
  AOI211_X1 U9707 ( .C1(n8884), .C2(n8166), .A(n8079), .B(n8078), .ZN(n8080)
         );
  NAND2_X1 U9708 ( .A1(n8081), .A2(n8080), .ZN(P2_U3225) );
  NOR2_X1 U9709 ( .A1(n4685), .A2(n8083), .ZN(n8084) );
  XNOR2_X1 U9710 ( .A(n8085), .B(n8084), .ZN(n8092) );
  OAI22_X1 U9711 ( .A1(n8159), .A2(n8087), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8086), .ZN(n8090) );
  OAI22_X1 U9712 ( .A1(n8163), .A2(n8624), .B1(n8088), .B2(n8160), .ZN(n8089)
         );
  AOI211_X1 U9713 ( .C1(n8863), .C2(n8166), .A(n8090), .B(n8089), .ZN(n8091)
         );
  OAI21_X1 U9714 ( .B1(n8092), .B2(n5614), .A(n8091), .ZN(P2_U3227) );
  XNOR2_X1 U9715 ( .A(n8093), .B(n8094), .ZN(n8157) );
  NOR2_X1 U9716 ( .A1(n8157), .A2(n8156), .ZN(n8155) );
  AOI21_X1 U9717 ( .B1(n8094), .B2(n8093), .A(n8155), .ZN(n8098) );
  XNOR2_X1 U9718 ( .A(n8096), .B(n8095), .ZN(n8097) );
  XNOR2_X1 U9719 ( .A(n8098), .B(n8097), .ZN(n8102) );
  AOI22_X1 U9720 ( .A1(n5616), .A2(n8784), .B1(n8124), .B2(n8773), .ZN(n8099)
         );
  NAND2_X1 U9721 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3152), .ZN(n8519) );
  OAI211_X1 U9722 ( .C1(n8283), .C2(n8159), .A(n8099), .B(n8519), .ZN(n8100)
         );
  AOI21_X1 U9723 ( .B1(n8783), .B2(n8166), .A(n8100), .ZN(n8101) );
  OAI21_X1 U9724 ( .B1(n8102), .B2(n5614), .A(n8101), .ZN(P2_U3228) );
  INV_X1 U9725 ( .A(n8103), .ZN(n8104) );
  AOI211_X1 U9726 ( .C1(n8106), .C2(n8105), .A(n5614), .B(n8104), .ZN(n8110)
         );
  AOI22_X1 U9727 ( .A1(n8143), .A2(n8371), .B1(P2_REG3_REG_17__SCAN_IN), .B2(
        P2_U3152), .ZN(n8108) );
  AOI22_X1 U9728 ( .A1(n5616), .A2(n8748), .B1(n8124), .B2(n8801), .ZN(n8107)
         );
  OAI211_X1 U9729 ( .C1(n8750), .C2(n8146), .A(n8108), .B(n8107), .ZN(n8109)
         );
  OR2_X1 U9730 ( .A1(n8110), .A2(n8109), .ZN(P2_U3230) );
  NOR2_X1 U9731 ( .A1(n8112), .A2(n8111), .ZN(n8114) );
  AOI22_X1 U9732 ( .A1(n8143), .A2(n8646), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3152), .ZN(n8118) );
  AOI22_X1 U9733 ( .A1(n5616), .A2(n8638), .B1(n8124), .B2(n8645), .ZN(n8117)
         );
  NAND2_X1 U9734 ( .A1(n8867), .A2(n8166), .ZN(n8116) );
  AOI21_X1 U9735 ( .B1(n8120), .B2(n8119), .A(n5614), .ZN(n8122) );
  NAND2_X1 U9736 ( .A1(n8122), .A2(n8121), .ZN(n8128) );
  AOI22_X1 U9737 ( .A1(n8143), .A2(n8711), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3152), .ZN(n8127) );
  INV_X1 U9738 ( .A(n8123), .ZN(n8708) );
  AOI22_X1 U9739 ( .A1(n5616), .A2(n8708), .B1(n8124), .B2(n8739), .ZN(n8126)
         );
  NAND2_X1 U9740 ( .A1(n8889), .A2(n8166), .ZN(n8125) );
  NAND4_X1 U9741 ( .A1(n8128), .A2(n8127), .A3(n8126), .A4(n8125), .ZN(
        P2_U3235) );
  XOR2_X1 U9742 ( .A(n8130), .B(n8129), .Z(n8136) );
  OAI22_X1 U9743 ( .A1(n8159), .A2(n8682), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8131), .ZN(n8134) );
  INV_X1 U9744 ( .A(n8672), .ZN(n8132) );
  OAI22_X1 U9745 ( .A1(n8163), .A2(n8132), .B1(n8681), .B2(n8160), .ZN(n8133)
         );
  AOI211_X1 U9746 ( .C1(n8879), .C2(n8166), .A(n8134), .B(n8133), .ZN(n8135)
         );
  OAI21_X1 U9747 ( .B1(n8136), .B2(n5614), .A(n8135), .ZN(P2_U3237) );
  OAI211_X1 U9748 ( .C1(n8140), .C2(n8139), .A(n8138), .B(n4315), .ZN(n8145)
         );
  AND2_X1 U9749 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8551) );
  INV_X1 U9750 ( .A(n8732), .ZN(n8141) );
  OAI22_X1 U9751 ( .A1(n8163), .A2(n8141), .B1(n8283), .B2(n8160), .ZN(n8142)
         );
  AOI211_X1 U9752 ( .C1(n8143), .C2(n8739), .A(n8551), .B(n8142), .ZN(n8144)
         );
  OAI211_X1 U9753 ( .C1(n8734), .C2(n8146), .A(n8145), .B(n8144), .ZN(P2_U3240) );
  XNOR2_X1 U9754 ( .A(n8147), .B(n8148), .ZN(n8154) );
  OAI22_X1 U9755 ( .A1(n8159), .A2(n8149), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9941), .ZN(n8152) );
  OAI22_X1 U9756 ( .A1(n8163), .A2(n8609), .B1(n8150), .B2(n8160), .ZN(n8151)
         );
  AOI211_X1 U9757 ( .C1(n8858), .C2(n8166), .A(n8152), .B(n8151), .ZN(n8153)
         );
  OAI21_X1 U9758 ( .B1(n8154), .B2(n5614), .A(n8153), .ZN(P2_U3242) );
  AOI21_X1 U9759 ( .B1(n8157), .B2(n8156), .A(n8155), .ZN(n8168) );
  OAI22_X1 U9760 ( .A1(n8159), .A2(n8757), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8158), .ZN(n8165) );
  INV_X1 U9761 ( .A(n8797), .ZN(n8162) );
  OAI22_X1 U9762 ( .A1(n8163), .A2(n8162), .B1(n8161), .B2(n8160), .ZN(n8164)
         );
  AOI211_X1 U9763 ( .C1(n8918), .C2(n8166), .A(n8165), .B(n8164), .ZN(n8167)
         );
  OAI21_X1 U9764 ( .B1(n8168), .B2(n5614), .A(n8167), .ZN(P2_U3243) );
  NOR2_X1 U9765 ( .A1(n8835), .A2(n8347), .ZN(n8341) );
  NAND2_X1 U9766 ( .A1(n8172), .A2(n8171), .ZN(n8174) );
  NAND2_X1 U9767 ( .A1(n8014), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n8173) );
  NOR2_X1 U9768 ( .A1(n8578), .A2(n8369), .ZN(n8332) );
  NOR2_X1 U9769 ( .A1(n8341), .A2(n8332), .ZN(n8354) );
  NAND2_X1 U9770 ( .A1(n8835), .A2(n8347), .ZN(n8352) );
  INV_X1 U9771 ( .A(n8369), .ZN(n8175) );
  NAND2_X1 U9772 ( .A1(n8352), .A2(n8351), .ZN(n8339) );
  INV_X1 U9773 ( .A(n8339), .ZN(n8196) );
  INV_X1 U9774 ( .A(n8589), .ZN(n8194) );
  INV_X1 U9775 ( .A(n8640), .ZN(n8310) );
  INV_X1 U9776 ( .A(n6818), .ZN(n8177) );
  NAND4_X1 U9777 ( .A1(n4855), .A2(n8220), .A3(n8199), .A4(n8177), .ZN(n8179)
         );
  NOR4_X1 U9778 ( .A1(n8180), .A2(n8179), .A3(n8178), .A4(n9769), .ZN(n8181)
         );
  NAND4_X1 U9779 ( .A1(n8247), .A2(n8239), .A3(n8819), .A4(n8181), .ZN(n8185)
         );
  NOR4_X1 U9780 ( .A1(n8185), .A2(n8184), .A3(n8183), .A4(n7449), .ZN(n8186)
         );
  NAND4_X1 U9781 ( .A1(n8269), .A2(n8188), .A3(n8187), .A4(n8186), .ZN(n8189)
         );
  NOR4_X1 U9782 ( .A1(n8735), .A2(n8769), .A3(n8799), .A4(n8189), .ZN(n8190)
         );
  INV_X1 U9783 ( .A(n8753), .ZN(n8282) );
  NAND4_X1 U9784 ( .A1(n8028), .A2(n8718), .A3(n8190), .A4(n8282), .ZN(n8191)
         );
  NOR4_X1 U9785 ( .A1(n4758), .A2(n8667), .A3(n8694), .A4(n8191), .ZN(n8192)
         );
  NAND4_X1 U9786 ( .A1(n8614), .A2(n8620), .A3(n8310), .A4(n8192), .ZN(n8193)
         );
  NOR4_X1 U9787 ( .A1(n8330), .A2(n8194), .A3(n8599), .A4(n8193), .ZN(n8195)
         );
  NAND3_X1 U9788 ( .A1(n8354), .A2(n8196), .A3(n8195), .ZN(n8197) );
  XNOR2_X1 U9789 ( .A(n8197), .B(n8569), .ZN(n8200) );
  OAI22_X1 U9790 ( .A1(n8200), .A2(n8346), .B1(n8199), .B2(n8198), .ZN(n8362)
         );
  NOR2_X1 U9791 ( .A1(n8201), .A2(n8569), .ZN(n8202) );
  NAND2_X1 U9792 ( .A1(n8251), .A2(n8250), .ZN(n8205) );
  NAND2_X1 U9793 ( .A1(n8203), .A2(n8206), .ZN(n8204) );
  MUX2_X1 U9794 ( .A(n8205), .B(n8204), .S(n8338), .Z(n8252) );
  INV_X1 U9795 ( .A(n8252), .ZN(n8258) );
  INV_X1 U9796 ( .A(n8206), .ZN(n8257) );
  INV_X1 U9797 ( .A(n8231), .ZN(n8210) );
  INV_X1 U9798 ( .A(n8237), .ZN(n8215) );
  NOR2_X1 U9799 ( .A1(n8216), .A2(n8322), .ZN(n8234) );
  AOI21_X1 U9800 ( .B1(n8346), .B2(n8225), .A(n8217), .ZN(n8219) );
  NAND2_X1 U9801 ( .A1(n8224), .A2(n8228), .ZN(n8218) );
  OAI211_X1 U9802 ( .C1(n8219), .C2(n8218), .A(n9739), .B(n8338), .ZN(n8221)
         );
  NAND2_X1 U9803 ( .A1(n8221), .A2(n8220), .ZN(n8222) );
  NOR2_X1 U9804 ( .A1(n8223), .A2(n8222), .ZN(n8233) );
  INV_X1 U9805 ( .A(n8224), .ZN(n8227) );
  INV_X1 U9806 ( .A(n8225), .ZN(n8226) );
  OAI211_X1 U9807 ( .C1(n8227), .C2(n8226), .A(n9739), .B(n7046), .ZN(n8229)
         );
  NAND3_X1 U9808 ( .A1(n8229), .A2(n8322), .A3(n8228), .ZN(n8230) );
  AND2_X1 U9809 ( .A1(n8231), .A2(n8230), .ZN(n8232) );
  OAI21_X1 U9810 ( .B1(n8234), .B2(n8233), .A(n8232), .ZN(n8235) );
  OAI211_X1 U9811 ( .C1(n8245), .C2(n8252), .A(n8244), .B(n8243), .ZN(n8255)
         );
  OAI211_X1 U9812 ( .C1(n8253), .C2(n8252), .A(n8259), .B(n8251), .ZN(n8254)
         );
  AOI21_X1 U9813 ( .B1(n8258), .B2(n8257), .A(n8256), .ZN(n8264) );
  OAI21_X1 U9814 ( .B1(n8264), .B2(n4409), .A(n8263), .ZN(n8265) );
  MUX2_X1 U9815 ( .A(n8267), .B(n8266), .S(n8338), .Z(n8268) );
  OAI211_X1 U9816 ( .C1(n8271), .C2(n8270), .A(n8269), .B(n8268), .ZN(n8276)
         );
  MUX2_X1 U9817 ( .A(n8273), .B(n8272), .S(n8338), .Z(n8274) );
  NAND3_X1 U9818 ( .A1(n8276), .A2(n8275), .A3(n8274), .ZN(n8280) );
  MUX2_X1 U9819 ( .A(n8278), .B(n8277), .S(n8338), .Z(n8279) );
  NAND4_X1 U9820 ( .A1(n8280), .A2(n8282), .A3(n8765), .A4(n8279), .ZN(n8290)
         );
  NOR2_X1 U9821 ( .A1(n8783), .A2(n8757), .ZN(n8281) );
  AOI21_X1 U9822 ( .B1(n8282), .B2(n8281), .A(n8736), .ZN(n8288) );
  NAND2_X1 U9823 ( .A1(n8905), .A2(n8283), .ZN(n8284) );
  OAI211_X1 U9824 ( .C1(n8753), .C2(n8285), .A(n8284), .B(n8294), .ZN(n8286)
         );
  INV_X1 U9825 ( .A(n8286), .ZN(n8287) );
  MUX2_X1 U9826 ( .A(n8288), .B(n8287), .S(n8322), .Z(n8289) );
  MUX2_X1 U9827 ( .A(n8322), .B(n8293), .S(n8292), .Z(n8307) );
  NAND3_X1 U9828 ( .A1(n8296), .A2(n8295), .A3(n8294), .ZN(n8300) );
  INV_X1 U9829 ( .A(n8297), .ZN(n8298) );
  AOI21_X1 U9830 ( .B1(n8300), .B2(n8299), .A(n8298), .ZN(n8304) );
  NAND2_X1 U9831 ( .A1(n8302), .A2(n8301), .ZN(n8303) );
  OAI211_X1 U9832 ( .C1(n8304), .C2(n8303), .A(n8306), .B(n8678), .ZN(n8305)
         );
  NAND3_X1 U9833 ( .A1(n8663), .A2(n8322), .A3(n8645), .ZN(n8309) );
  NAND3_X1 U9834 ( .A1(n8873), .A2(n8682), .A3(n8338), .ZN(n8308) );
  MUX2_X1 U9835 ( .A(n8312), .B(n8311), .S(n8338), .Z(n8313) );
  NAND2_X1 U9836 ( .A1(n8317), .A2(n8315), .ZN(n8316) );
  INV_X1 U9837 ( .A(n8321), .ZN(n8323) );
  NAND2_X1 U9838 ( .A1(n8329), .A2(n8327), .ZN(n8328) );
  INV_X1 U9839 ( .A(n8332), .ZN(n8335) );
  MUX2_X1 U9840 ( .A(n8333), .B(n8348), .S(n8338), .Z(n8334) );
  NAND3_X1 U9841 ( .A1(n8351), .A2(n8335), .A3(n8334), .ZN(n8336) );
  OAI22_X1 U9842 ( .A1(n8337), .A2(n8336), .B1(n8354), .B2(n8338), .ZN(n8340)
         );
  AOI22_X1 U9843 ( .A1(n8340), .A2(n8352), .B1(n8339), .B2(n8338), .ZN(n8345)
         );
  INV_X1 U9844 ( .A(n8341), .ZN(n8342) );
  NOR2_X1 U9845 ( .A1(n8342), .A2(n8322), .ZN(n8344) );
  NAND2_X1 U9846 ( .A1(n8347), .A2(n8346), .ZN(n8350) );
  INV_X1 U9847 ( .A(n8352), .ZN(n8353) );
  NOR2_X1 U9848 ( .A1(n8361), .A2(n8359), .ZN(n8360) );
  NOR4_X1 U9849 ( .A1(n9759), .A2(n8364), .A3(n8363), .A4(n8756), .ZN(n8367)
         );
  OAI21_X1 U9850 ( .B1(n8368), .B2(n8365), .A(P2_B_REG_SCAN_IN), .ZN(n8366) );
  MUX2_X1 U9851 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8369), .S(P2_U3966), .Z(
        P2_U3582) );
  MUX2_X1 U9852 ( .A(n8590), .B(P2_DATAO_REG_29__SCAN_IN), .S(n8370), .Z(
        P2_U3581) );
  MUX2_X1 U9853 ( .A(n8601), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8370), .Z(
        P2_U3580) );
  MUX2_X1 U9854 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8615), .S(P2_U3966), .Z(
        P2_U3579) );
  MUX2_X1 U9855 ( .A(n8630), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8370), .Z(
        P2_U3578) );
  MUX2_X1 U9856 ( .A(n8646), .B(P2_DATAO_REG_25__SCAN_IN), .S(n8370), .Z(
        P2_U3577) );
  MUX2_X1 U9857 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8653), .S(P2_U3966), .Z(
        P2_U3576) );
  MUX2_X1 U9858 ( .A(n8645), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8370), .Z(
        P2_U3575) );
  MUX2_X1 U9859 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8711), .S(P2_U3966), .Z(
        P2_U3573) );
  MUX2_X1 U9860 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8698), .S(P2_U3966), .Z(
        P2_U3572) );
  MUX2_X1 U9861 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8739), .S(P2_U3966), .Z(
        P2_U3571) );
  MUX2_X1 U9862 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8371), .S(P2_U3966), .Z(
        P2_U3570) );
  MUX2_X1 U9863 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8774), .S(P2_U3966), .Z(
        P2_U3569) );
  MUX2_X1 U9864 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8801), .S(P2_U3966), .Z(
        P2_U3568) );
  MUX2_X1 U9865 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8773), .S(P2_U3966), .Z(
        P2_U3567) );
  MUX2_X1 U9866 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8802), .S(P2_U3966), .Z(
        P2_U3566) );
  MUX2_X1 U9867 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n8372), .S(P2_U3966), .Z(
        P2_U3565) );
  MUX2_X1 U9868 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n8373), .S(P2_U3966), .Z(
        P2_U3564) );
  MUX2_X1 U9869 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n8374), .S(P2_U3966), .Z(
        P2_U3563) );
  MUX2_X1 U9870 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n8375), .S(P2_U3966), .Z(
        P2_U3562) );
  MUX2_X1 U9871 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n8376), .S(P2_U3966), .Z(
        P2_U3561) );
  MUX2_X1 U9872 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n8377), .S(P2_U3966), .Z(
        P2_U3560) );
  MUX2_X1 U9873 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n8811), .S(P2_U3966), .Z(
        P2_U3559) );
  MUX2_X1 U9874 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n8378), .S(P2_U3966), .Z(
        P2_U3558) );
  MUX2_X1 U9875 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n8810), .S(P2_U3966), .Z(
        P2_U3557) );
  MUX2_X1 U9876 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n9745), .S(P2_U3966), .Z(
        P2_U3556) );
  MUX2_X1 U9877 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n8379), .S(P2_U3966), .Z(
        P2_U3555) );
  MUX2_X1 U9878 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n7029), .S(P2_U3966), .Z(
        P2_U3554) );
  MUX2_X1 U9879 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n6817), .S(P2_U3966), .Z(
        P2_U3553) );
  MUX2_X1 U9880 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n8380), .S(P2_U3966), .Z(
        P2_U3552) );
  OAI211_X1 U9881 ( .C1(n8383), .C2(n8382), .A(n9728), .B(n8381), .ZN(n8393)
         );
  NOR2_X1 U9882 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5001), .ZN(n8384) );
  AOI21_X1 U9883 ( .B1(n9734), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n8384), .ZN(
        n8392) );
  NAND2_X1 U9884 ( .A1(n9534), .A2(n8385), .ZN(n8391) );
  AOI21_X1 U9885 ( .B1(n8388), .B2(n8387), .A(n8386), .ZN(n8389) );
  NAND2_X1 U9886 ( .A1(n9729), .A2(n8389), .ZN(n8390) );
  NAND4_X1 U9887 ( .A1(n8393), .A2(n8392), .A3(n8391), .A4(n8390), .ZN(
        P2_U3248) );
  OAI211_X1 U9888 ( .C1(n8396), .C2(n8395), .A(n9728), .B(n8394), .ZN(n8407)
         );
  INV_X1 U9889 ( .A(n8397), .ZN(n8398) );
  AOI21_X1 U9890 ( .B1(n9734), .B2(P2_ADDR_REG_4__SCAN_IN), .A(n8398), .ZN(
        n8406) );
  NAND2_X1 U9891 ( .A1(n9534), .A2(n8399), .ZN(n8405) );
  AOI21_X1 U9892 ( .B1(n8402), .B2(n8401), .A(n8400), .ZN(n8403) );
  NAND2_X1 U9893 ( .A1(n9729), .A2(n8403), .ZN(n8404) );
  NAND4_X1 U9894 ( .A1(n8407), .A2(n8406), .A3(n8405), .A4(n8404), .ZN(
        P2_U3249) );
  OAI211_X1 U9895 ( .C1(n8410), .C2(n8409), .A(n9728), .B(n8408), .ZN(n8421)
         );
  NOR2_X1 U9896 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8411), .ZN(n8412) );
  AOI21_X1 U9897 ( .B1(n9734), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n8412), .ZN(
        n8420) );
  NAND2_X1 U9898 ( .A1(n9534), .A2(n8413), .ZN(n8419) );
  AOI21_X1 U9899 ( .B1(n8416), .B2(n8415), .A(n8414), .ZN(n8417) );
  NAND2_X1 U9900 ( .A1(n9729), .A2(n8417), .ZN(n8418) );
  NAND4_X1 U9901 ( .A1(n8421), .A2(n8420), .A3(n8419), .A4(n8418), .ZN(
        P2_U3250) );
  OAI211_X1 U9902 ( .C1(n8424), .C2(n8423), .A(n9728), .B(n8422), .ZN(n8435)
         );
  INV_X1 U9903 ( .A(n8425), .ZN(n8426) );
  AOI21_X1 U9904 ( .B1(n9734), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n8426), .ZN(
        n8434) );
  NAND2_X1 U9905 ( .A1(n9534), .A2(n8427), .ZN(n8433) );
  AOI21_X1 U9906 ( .B1(n8430), .B2(n8429), .A(n8428), .ZN(n8431) );
  NAND2_X1 U9907 ( .A1(n9729), .A2(n8431), .ZN(n8432) );
  NAND4_X1 U9908 ( .A1(n8435), .A2(n8434), .A3(n8433), .A4(n8432), .ZN(
        P2_U3251) );
  OAI211_X1 U9909 ( .C1(n8438), .C2(n8437), .A(n9728), .B(n8436), .ZN(n8449)
         );
  NOR2_X1 U9910 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8439), .ZN(n8440) );
  AOI21_X1 U9911 ( .B1(n9734), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n8440), .ZN(
        n8448) );
  NAND2_X1 U9912 ( .A1(n9534), .A2(n8441), .ZN(n8447) );
  AOI21_X1 U9913 ( .B1(n8444), .B2(n8443), .A(n8442), .ZN(n8445) );
  NAND2_X1 U9914 ( .A1(n9729), .A2(n8445), .ZN(n8446) );
  NAND4_X1 U9915 ( .A1(n8449), .A2(n8448), .A3(n8447), .A4(n8446), .ZN(
        P2_U3252) );
  OAI211_X1 U9916 ( .C1(n8452), .C2(n8451), .A(n9728), .B(n8450), .ZN(n8463)
         );
  INV_X1 U9917 ( .A(n8453), .ZN(n8454) );
  AOI21_X1 U9918 ( .B1(n9734), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n8454), .ZN(
        n8462) );
  NAND2_X1 U9919 ( .A1(n9534), .A2(n8455), .ZN(n8461) );
  AOI21_X1 U9920 ( .B1(n8458), .B2(n8457), .A(n8456), .ZN(n8459) );
  NAND2_X1 U9921 ( .A1(n9729), .A2(n8459), .ZN(n8460) );
  NAND4_X1 U9922 ( .A1(n8463), .A2(n8462), .A3(n8461), .A4(n8460), .ZN(
        P2_U3253) );
  OAI211_X1 U9923 ( .C1(n8466), .C2(n8465), .A(n9728), .B(n8464), .ZN(n8477)
         );
  INV_X1 U9924 ( .A(n8467), .ZN(n8468) );
  AOI21_X1 U9925 ( .B1(n9734), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n8468), .ZN(
        n8476) );
  NAND2_X1 U9926 ( .A1(n9534), .A2(n8469), .ZN(n8475) );
  AOI21_X1 U9927 ( .B1(n8472), .B2(n8471), .A(n8470), .ZN(n8473) );
  NAND2_X1 U9928 ( .A1(n9729), .A2(n8473), .ZN(n8474) );
  NAND4_X1 U9929 ( .A1(n8477), .A2(n8476), .A3(n8475), .A4(n8474), .ZN(
        P2_U3254) );
  OAI211_X1 U9930 ( .C1(n8480), .C2(n8479), .A(n9728), .B(n8478), .ZN(n8491)
         );
  INV_X1 U9931 ( .A(n8481), .ZN(n8482) );
  AOI21_X1 U9932 ( .B1(n9734), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n8482), .ZN(
        n8490) );
  NAND2_X1 U9933 ( .A1(n9534), .A2(n8483), .ZN(n8489) );
  OAI21_X1 U9934 ( .B1(n8486), .B2(n8485), .A(n8484), .ZN(n8487) );
  NAND2_X1 U9935 ( .A1(n9729), .A2(n8487), .ZN(n8488) );
  NAND4_X1 U9936 ( .A1(n8491), .A2(n8490), .A3(n8489), .A4(n8488), .ZN(
        P2_U3257) );
  OAI21_X1 U9937 ( .B1(n8493), .B2(P2_REG1_REG_14__SCAN_IN), .A(n8492), .ZN(
        n8506) );
  XNOR2_X1 U9938 ( .A(n8506), .B(n8507), .ZN(n8495) );
  INV_X1 U9939 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8494) );
  NOR2_X1 U9940 ( .A1(n8494), .A2(n8495), .ZN(n8508) );
  AOI211_X1 U9941 ( .C1(n8495), .C2(n8494), .A(n8508), .B(n9528), .ZN(n8505)
         );
  AOI21_X1 U9942 ( .B1(n8498), .B2(n8497), .A(n8496), .ZN(n8512) );
  XNOR2_X1 U9943 ( .A(n8512), .B(n8513), .ZN(n8499) );
  NOR2_X1 U9944 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n8499), .ZN(n8514) );
  AOI21_X1 U9945 ( .B1(n8499), .B2(P2_REG2_REG_15__SCAN_IN), .A(n8514), .ZN(
        n8500) );
  NOR2_X1 U9946 ( .A1(n8500), .A2(n9732), .ZN(n8504) );
  AND2_X1 U9947 ( .A1(P2_U3152), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8501) );
  AOI21_X1 U9948 ( .B1(n9734), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n8501), .ZN(
        n8502) );
  OAI21_X1 U9949 ( .B1(n9730), .B2(n8507), .A(n8502), .ZN(n8503) );
  OR3_X1 U9950 ( .A1(n8505), .A2(n8504), .A3(n8503), .ZN(P2_U3260) );
  NOR2_X1 U9951 ( .A1(n8507), .A2(n8506), .ZN(n8509) );
  NOR2_X1 U9952 ( .A1(n8509), .A2(n8508), .ZN(n8511) );
  XNOR2_X1 U9953 ( .A(n8523), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n8510) );
  NAND2_X1 U9954 ( .A1(n8510), .A2(n8511), .ZN(n8534) );
  OAI21_X1 U9955 ( .B1(n8511), .B2(n8510), .A(n8534), .ZN(n8525) );
  NOR2_X1 U9956 ( .A1(n8513), .A2(n8512), .ZN(n8515) );
  NOR2_X1 U9957 ( .A1(n8515), .A2(n8514), .ZN(n8518) );
  INV_X1 U9958 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8516) );
  NOR2_X1 U9959 ( .A1(n8523), .A2(n8516), .ZN(n8527) );
  AOI21_X1 U9960 ( .B1(n8516), .B2(n8523), .A(n8527), .ZN(n8517) );
  NAND2_X1 U9961 ( .A1(n8517), .A2(n8518), .ZN(n8528) );
  OAI211_X1 U9962 ( .C1(n8518), .C2(n8517), .A(n9728), .B(n8528), .ZN(n8522)
         );
  INV_X1 U9963 ( .A(n8519), .ZN(n8520) );
  AOI21_X1 U9964 ( .B1(n9734), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n8520), .ZN(
        n8521) );
  OAI211_X1 U9965 ( .C1(n9730), .C2(n8523), .A(n8522), .B(n8521), .ZN(n8524)
         );
  AOI21_X1 U9966 ( .B1(n8525), .B2(n9729), .A(n8524), .ZN(n8526) );
  INV_X1 U9967 ( .A(n8526), .ZN(P2_U3261) );
  INV_X1 U9968 ( .A(n8527), .ZN(n8529) );
  NAND2_X1 U9969 ( .A1(n8529), .A2(n8528), .ZN(n8532) );
  OR2_X1 U9970 ( .A1(n8549), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8530) );
  NAND2_X1 U9971 ( .A1(n8549), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8544) );
  AND2_X1 U9972 ( .A1(n8530), .A2(n8544), .ZN(n8531) );
  NAND2_X1 U9973 ( .A1(n8531), .A2(n8532), .ZN(n8543) );
  OAI211_X1 U9974 ( .C1(n8532), .C2(n8531), .A(n9728), .B(n8543), .ZN(n8541)
         );
  NOR2_X1 U9975 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8533), .ZN(n8539) );
  XNOR2_X1 U9976 ( .A(n8549), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n8536) );
  AOI211_X1 U9977 ( .C1(n8537), .C2(n8536), .A(n8548), .B(n9528), .ZN(n8538)
         );
  AOI211_X1 U9978 ( .C1(P2_ADDR_REG_17__SCAN_IN), .C2(n9734), .A(n8539), .B(
        n8538), .ZN(n8540) );
  OAI211_X1 U9979 ( .C1(n9730), .C2(n8542), .A(n8541), .B(n8540), .ZN(P2_U3262) );
  NAND2_X1 U9980 ( .A1(n8544), .A2(n8543), .ZN(n8545) );
  NOR2_X1 U9981 ( .A1(n8545), .A2(n8560), .ZN(n8558) );
  AOI21_X1 U9982 ( .B1(n8545), .B2(n8560), .A(n8558), .ZN(n8546) );
  INV_X1 U9983 ( .A(n8546), .ZN(n8547) );
  NOR2_X1 U9984 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n8547), .ZN(n8557) );
  AOI21_X1 U9985 ( .B1(n8547), .B2(P2_REG2_REG_18__SCAN_IN), .A(n8557), .ZN(
        n8556) );
  INV_X1 U9986 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8550) );
  XNOR2_X1 U9987 ( .A(n8560), .B(n8550), .ZN(n8563) );
  XOR2_X1 U9988 ( .A(n8562), .B(n8563), .Z(n8553) );
  AOI21_X1 U9989 ( .B1(n9734), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n8551), .ZN(
        n8552) );
  OAI21_X1 U9990 ( .B1(n9528), .B2(n8553), .A(n8552), .ZN(n8554) );
  AOI21_X1 U9991 ( .B1(n8560), .B2(n9534), .A(n8554), .ZN(n8555) );
  OAI21_X1 U9992 ( .B1(n8556), .B2(n9732), .A(n8555), .ZN(P2_U3263) );
  NOR2_X1 U9993 ( .A1(n8558), .A2(n8557), .ZN(n8559) );
  XNOR2_X1 U9994 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n8559), .ZN(n8568) );
  INV_X1 U9995 ( .A(n8568), .ZN(n8566) );
  NOR2_X1 U9996 ( .A1(n8560), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8561) );
  XNOR2_X1 U9997 ( .A(n8564), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8567) );
  NAND2_X1 U9998 ( .A1(n9729), .A2(n8567), .ZN(n8565) );
  OAI22_X1 U9999 ( .A1(n8568), .A2(n9732), .B1(n8567), .B2(n9528), .ZN(n8570)
         );
  NAND2_X1 U10000 ( .A1(n8578), .A2(n8577), .ZN(n8576) );
  NAND2_X1 U10001 ( .A1(n8573), .A2(n8572), .ZN(n8840) );
  NOR2_X1 U10002 ( .A1(n8804), .A2(n8840), .ZN(n8580) );
  AOI21_X1 U10003 ( .B1(n8804), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8580), .ZN(
        n8575) );
  NAND2_X1 U10004 ( .A1(n8835), .A2(n8827), .ZN(n8574) );
  OAI211_X1 U10005 ( .C1(n8837), .C2(n8582), .A(n8575), .B(n8574), .ZN(
        P2_U3265) );
  OAI21_X1 U10006 ( .B1(n8578), .B2(n8577), .A(n8576), .ZN(n8841) );
  NOR2_X1 U10007 ( .A1(n8578), .A2(n8821), .ZN(n8579) );
  AOI211_X1 U10008 ( .C1(n8804), .C2(P2_REG2_REG_30__SCAN_IN), .A(n8580), .B(
        n8579), .ZN(n8581) );
  OAI21_X1 U10009 ( .B1(n8582), .B2(n8841), .A(n8581), .ZN(P2_U3266) );
  XOR2_X1 U10010 ( .A(n8589), .B(n8583), .Z(n8851) );
  INV_X1 U10011 ( .A(n8584), .ZN(n8585) );
  AOI21_X1 U10012 ( .B1(n8847), .B2(n8595), .A(n8585), .ZN(n8848) );
  AOI22_X1 U10013 ( .A1(n8804), .A2(P2_REG2_REG_28__SCAN_IN), .B1(n8586), .B2(
        n9747), .ZN(n8587) );
  OAI21_X1 U10014 ( .B1(n5613), .B2(n8821), .A(n8587), .ZN(n8592) );
  AOI211_X1 U10015 ( .C1(n7043), .C2(n8848), .A(n8592), .B(n8591), .ZN(n8593)
         );
  OAI21_X1 U10016 ( .B1(n8851), .B2(n8764), .A(n8593), .ZN(P2_U3268) );
  XNOR2_X1 U10017 ( .A(n8594), .B(n4779), .ZN(n8856) );
  INV_X1 U10018 ( .A(n8595), .ZN(n8596) );
  AOI21_X1 U10019 ( .B1(n8852), .B2(n8607), .A(n8596), .ZN(n8853) );
  AOI22_X1 U10020 ( .A1(n8804), .A2(P2_REG2_REG_27__SCAN_IN), .B1(n8597), .B2(
        n9747), .ZN(n8598) );
  OAI21_X1 U10021 ( .B1(n4529), .B2(n8821), .A(n8598), .ZN(n8604) );
  XNOR2_X1 U10022 ( .A(n8600), .B(n8599), .ZN(n8602) );
  AOI222_X1 U10023 ( .A1(n8813), .A2(n8602), .B1(n8630), .B2(n9743), .C1(n8601), .C2(n9744), .ZN(n8855) );
  NOR2_X1 U10024 ( .A1(n8855), .A2(n8804), .ZN(n8603) );
  AOI211_X1 U10025 ( .C1(n7043), .C2(n8853), .A(n8604), .B(n8603), .ZN(n8605)
         );
  OAI21_X1 U10026 ( .B1(n8856), .B2(n8764), .A(n8605), .ZN(P2_U3269) );
  XOR2_X1 U10027 ( .A(n8614), .B(n8606), .Z(n8861) );
  INV_X1 U10028 ( .A(n8607), .ZN(n8608) );
  AOI211_X1 U10029 ( .C1(n8858), .C2(n4533), .A(n9825), .B(n8608), .ZN(n8857)
         );
  INV_X1 U10030 ( .A(n8609), .ZN(n8610) );
  AOI22_X1 U10031 ( .A1(n8804), .A2(P2_REG2_REG_26__SCAN_IN), .B1(n8610), .B2(
        n9747), .ZN(n8611) );
  OAI21_X1 U10032 ( .B1(n8612), .B2(n8821), .A(n8611), .ZN(n8618) );
  XOR2_X1 U10033 ( .A(n8614), .B(n8613), .Z(n8616) );
  AOI222_X1 U10034 ( .A1(n8813), .A2(n8616), .B1(n8615), .B2(n9744), .C1(n8646), .C2(n9743), .ZN(n8860) );
  NOR2_X1 U10035 ( .A1(n8860), .A2(n8804), .ZN(n8617) );
  AOI211_X1 U10036 ( .C1(n8857), .C2(n8762), .A(n8618), .B(n8617), .ZN(n8619)
         );
  OAI21_X1 U10037 ( .B1(n8861), .B2(n8764), .A(n8619), .ZN(P2_U3270) );
  XNOR2_X1 U10038 ( .A(n8621), .B(n8620), .ZN(n8866) );
  AOI211_X1 U10039 ( .C1(n8863), .C2(n8623), .A(n9825), .B(n8622), .ZN(n8862)
         );
  INV_X1 U10040 ( .A(n8624), .ZN(n8625) );
  AOI22_X1 U10041 ( .A1(n8804), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n8625), .B2(
        n9747), .ZN(n8626) );
  OAI21_X1 U10042 ( .B1(n8627), .B2(n8821), .A(n8626), .ZN(n8633) );
  XNOR2_X1 U10043 ( .A(n8629), .B(n8628), .ZN(n8631) );
  AOI222_X1 U10044 ( .A1(n8813), .A2(n8631), .B1(n8630), .B2(n9744), .C1(n8653), .C2(n9743), .ZN(n8865) );
  NOR2_X1 U10045 ( .A1(n8865), .A2(n8804), .ZN(n8632) );
  AOI211_X1 U10046 ( .C1(n8762), .C2(n8862), .A(n8633), .B(n8632), .ZN(n8634)
         );
  OAI21_X1 U10047 ( .B1(n8866), .B2(n8764), .A(n8634), .ZN(P2_U3271) );
  OAI21_X1 U10048 ( .B1(n8636), .B2(n8640), .A(n8635), .ZN(n8637) );
  INV_X1 U10049 ( .A(n8637), .ZN(n8871) );
  XNOR2_X1 U10050 ( .A(n8658), .B(n8867), .ZN(n8868) );
  AOI22_X1 U10051 ( .A1(n8804), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n8638), .B2(
        n9747), .ZN(n8639) );
  OAI21_X1 U10052 ( .B1(n8009), .B2(n8821), .A(n8639), .ZN(n8650) );
  INV_X1 U10053 ( .A(n8652), .ZN(n8642) );
  OAI21_X1 U10054 ( .B1(n8642), .B2(n8641), .A(n8640), .ZN(n8644) );
  NAND3_X1 U10055 ( .A1(n8644), .A2(n8813), .A3(n8643), .ZN(n8648) );
  AOI22_X1 U10056 ( .A1(n8646), .A2(n9744), .B1(n9743), .B2(n8645), .ZN(n8647)
         );
  AND2_X1 U10057 ( .A1(n8648), .A2(n8647), .ZN(n8870) );
  NOR2_X1 U10058 ( .A1(n8870), .A2(n8804), .ZN(n8649) );
  AOI211_X1 U10059 ( .C1(n8868), .C2(n7043), .A(n8650), .B(n8649), .ZN(n8651)
         );
  OAI21_X1 U10060 ( .B1(n8871), .B2(n8764), .A(n8651), .ZN(P2_U3272) );
  OAI21_X1 U10061 ( .B1(n4894), .B2(n8655), .A(n8652), .ZN(n8654) );
  AOI222_X1 U10062 ( .A1(n8813), .A2(n8654), .B1(n8699), .B2(n9743), .C1(n8653), .C2(n9744), .ZN(n8876) );
  INV_X1 U10063 ( .A(n8878), .ZN(n8657) );
  NAND2_X1 U10064 ( .A1(n8656), .A2(n8655), .ZN(n8872) );
  NAND3_X1 U10065 ( .A1(n8657), .A2(n9754), .A3(n8872), .ZN(n8666) );
  INV_X1 U10066 ( .A(n8670), .ZN(n8659) );
  AOI21_X1 U10067 ( .B1(n8873), .B2(n8659), .A(n8658), .ZN(n8874) );
  INV_X1 U10068 ( .A(n8660), .ZN(n8661) );
  AOI22_X1 U10069 ( .A1(n8804), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n8661), .B2(
        n9747), .ZN(n8662) );
  OAI21_X1 U10070 ( .B1(n8663), .B2(n8821), .A(n8662), .ZN(n8664) );
  AOI21_X1 U10071 ( .B1(n8874), .B2(n7043), .A(n8664), .ZN(n8665) );
  OAI211_X1 U10072 ( .C1(n8804), .C2(n8876), .A(n8666), .B(n8665), .ZN(
        P2_U3273) );
  XNOR2_X1 U10073 ( .A(n8668), .B(n8667), .ZN(n8883) );
  INV_X1 U10074 ( .A(n8669), .ZN(n8671) );
  AOI21_X1 U10075 ( .B1(n8879), .B2(n8671), .A(n8670), .ZN(n8880) );
  AOI22_X1 U10076 ( .A1(n8804), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8672), .B2(
        n9747), .ZN(n8673) );
  OAI21_X1 U10077 ( .B1(n8674), .B2(n8821), .A(n8673), .ZN(n8686) );
  INV_X1 U10078 ( .A(n8675), .ZN(n8680) );
  AOI21_X1 U10079 ( .B1(n8676), .B2(n8678), .A(n8677), .ZN(n8679) );
  NOR3_X1 U10080 ( .A1(n8680), .A2(n8679), .A3(n8751), .ZN(n8684) );
  OAI22_X1 U10081 ( .A1(n8682), .A2(n8754), .B1(n8681), .B2(n8756), .ZN(n8683)
         );
  NOR2_X1 U10082 ( .A1(n8684), .A2(n8683), .ZN(n8882) );
  NOR2_X1 U10083 ( .A1(n8882), .A2(n8804), .ZN(n8685) );
  AOI211_X1 U10084 ( .C1(n8880), .C2(n7043), .A(n8686), .B(n8685), .ZN(n8687)
         );
  OAI21_X1 U10085 ( .B1(n8883), .B2(n8764), .A(n8687), .ZN(P2_U3274) );
  XOR2_X1 U10086 ( .A(n8694), .B(n4316), .Z(n8888) );
  XNOR2_X1 U10087 ( .A(n8706), .B(n8692), .ZN(n8885) );
  INV_X1 U10088 ( .A(n8689), .ZN(n8690) );
  AOI22_X1 U10089 ( .A1(n8804), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8690), .B2(
        n9747), .ZN(n8691) );
  OAI21_X1 U10090 ( .B1(n8692), .B2(n8821), .A(n8691), .ZN(n8702) );
  INV_X1 U10091 ( .A(n8693), .ZN(n8696) );
  OAI21_X1 U10092 ( .B1(n8696), .B2(n8695), .A(n8694), .ZN(n8697) );
  NAND2_X1 U10093 ( .A1(n8697), .A2(n8676), .ZN(n8700) );
  AOI222_X1 U10094 ( .A1(n8813), .A2(n8700), .B1(n8699), .B2(n9744), .C1(n8698), .C2(n9743), .ZN(n8887) );
  NOR2_X1 U10095 ( .A1(n8887), .A2(n8804), .ZN(n8701) );
  AOI211_X1 U10096 ( .C1(n8885), .C2(n7043), .A(n8702), .B(n8701), .ZN(n8703)
         );
  OAI21_X1 U10097 ( .B1(n8888), .B2(n8764), .A(n8703), .ZN(P2_U3275) );
  XNOR2_X1 U10098 ( .A(n8705), .B(n8704), .ZN(n8893) );
  INV_X1 U10099 ( .A(n8706), .ZN(n8707) );
  AOI21_X1 U10100 ( .B1(n8889), .B2(n8721), .A(n8707), .ZN(n8890) );
  AOI22_X1 U10101 ( .A1(n8804), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8708), .B2(
        n9747), .ZN(n8709) );
  OAI21_X1 U10102 ( .B1(n4526), .B2(n8821), .A(n8709), .ZN(n8714) );
  XNOR2_X1 U10103 ( .A(n8710), .B(n8028), .ZN(n8712) );
  AOI222_X1 U10104 ( .A1(n8813), .A2(n8712), .B1(n8739), .B2(n9743), .C1(n8711), .C2(n9744), .ZN(n8892) );
  NOR2_X1 U10105 ( .A1(n8892), .A2(n8804), .ZN(n8713) );
  AOI211_X1 U10106 ( .C1(n8890), .C2(n7043), .A(n8714), .B(n8713), .ZN(n8715)
         );
  OAI21_X1 U10107 ( .B1(n8893), .B2(n8764), .A(n8715), .ZN(P2_U3276) );
  XOR2_X1 U10108 ( .A(n8716), .B(n8718), .Z(n8898) );
  XOR2_X1 U10109 ( .A(n8718), .B(n8717), .Z(n8720) );
  OAI21_X1 U10110 ( .B1(n8720), .B2(n8751), .A(n8719), .ZN(n8894) );
  INV_X1 U10111 ( .A(n8721), .ZN(n8722) );
  AOI211_X1 U10112 ( .C1(n8896), .C2(n8729), .A(n9825), .B(n8722), .ZN(n8895)
         );
  NAND2_X1 U10113 ( .A1(n8895), .A2(n8762), .ZN(n8725) );
  AOI22_X1 U10114 ( .A1(n8804), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n8723), .B2(
        n9747), .ZN(n8724) );
  OAI211_X1 U10115 ( .C1(n4527), .C2(n8821), .A(n8725), .B(n8724), .ZN(n8726)
         );
  AOI21_X1 U10116 ( .B1(n8894), .B2(n8830), .A(n8726), .ZN(n8727) );
  OAI21_X1 U10117 ( .B1(n8898), .B2(n8764), .A(n8727), .ZN(P2_U3277) );
  XOR2_X1 U10118 ( .A(n8728), .B(n8735), .Z(n8903) );
  INV_X1 U10119 ( .A(n8746), .ZN(n8731) );
  INV_X1 U10120 ( .A(n8729), .ZN(n8730) );
  AOI21_X1 U10121 ( .B1(n8899), .B2(n8731), .A(n8730), .ZN(n8900) );
  AOI22_X1 U10122 ( .A1(n8804), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8732), .B2(
        n9747), .ZN(n8733) );
  OAI21_X1 U10123 ( .B1(n8734), .B2(n8821), .A(n8733), .ZN(n8742) );
  OAI21_X1 U10124 ( .B1(n4376), .B2(n8736), .A(n8735), .ZN(n8738) );
  NAND2_X1 U10125 ( .A1(n8738), .A2(n8737), .ZN(n8740) );
  AOI222_X1 U10126 ( .A1(n8813), .A2(n8740), .B1(n8739), .B2(n9744), .C1(n8774), .C2(n9743), .ZN(n8902) );
  NOR2_X1 U10127 ( .A1(n8902), .A2(n8804), .ZN(n8741) );
  AOI211_X1 U10128 ( .C1(n8900), .C2(n7043), .A(n8742), .B(n8741), .ZN(n8743)
         );
  OAI21_X1 U10129 ( .B1(n8903), .B2(n8764), .A(n8743), .ZN(P2_U3278) );
  OAI21_X1 U10130 ( .B1(n4383), .B2(n8753), .A(n8744), .ZN(n8745) );
  INV_X1 U10131 ( .A(n8745), .ZN(n8908) );
  INV_X1 U10132 ( .A(n8781), .ZN(n8747) );
  AOI211_X1 U10133 ( .C1(n8905), .C2(n8747), .A(n9825), .B(n8746), .ZN(n8904)
         );
  AOI22_X1 U10134 ( .A1(n8804), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n8748), .B2(
        n9747), .ZN(n8749) );
  OAI21_X1 U10135 ( .B1(n8750), .B2(n8821), .A(n8749), .ZN(n8761) );
  AOI211_X1 U10136 ( .C1(n8753), .C2(n8752), .A(n8751), .B(n4376), .ZN(n8759)
         );
  OAI22_X1 U10137 ( .A1(n8757), .A2(n8756), .B1(n8755), .B2(n8754), .ZN(n8758)
         );
  NOR2_X1 U10138 ( .A1(n8759), .A2(n8758), .ZN(n8907) );
  NOR2_X1 U10139 ( .A1(n8907), .A2(n8804), .ZN(n8760) );
  AOI211_X1 U10140 ( .C1(n8904), .C2(n8762), .A(n8761), .B(n8760), .ZN(n8763)
         );
  OAI21_X1 U10141 ( .B1(n8908), .B2(n8764), .A(n8763), .ZN(P2_U3279) );
  AND2_X1 U10142 ( .A1(n8766), .A2(n8765), .ZN(n8768) );
  OR2_X1 U10143 ( .A1(n8768), .A2(n8767), .ZN(n8913) );
  NAND2_X1 U10144 ( .A1(n8770), .A2(n8769), .ZN(n8771) );
  NAND2_X1 U10145 ( .A1(n8772), .A2(n8771), .ZN(n8778) );
  NAND2_X1 U10146 ( .A1(n8773), .A2(n9743), .ZN(n8776) );
  NAND2_X1 U10147 ( .A1(n8774), .A2(n9744), .ZN(n8775) );
  NAND2_X1 U10148 ( .A1(n8776), .A2(n8775), .ZN(n8777) );
  AOI21_X1 U10149 ( .B1(n8778), .B2(n8813), .A(n8777), .ZN(n8779) );
  OAI21_X1 U10150 ( .B1(n8913), .B2(n8780), .A(n8779), .ZN(n8915) );
  NAND2_X1 U10151 ( .A1(n8915), .A2(n8830), .ZN(n8789) );
  AND2_X1 U10152 ( .A1(n8794), .A2(n8783), .ZN(n8782) );
  OR2_X1 U10153 ( .A1(n8782), .A2(n8781), .ZN(n8910) );
  INV_X1 U10154 ( .A(n8910), .ZN(n8787) );
  INV_X1 U10155 ( .A(n8783), .ZN(n8909) );
  AOI22_X1 U10156 ( .A1(n8804), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n8784), .B2(
        n9747), .ZN(n8785) );
  OAI21_X1 U10157 ( .B1(n8909), .B2(n8821), .A(n8785), .ZN(n8786) );
  AOI21_X1 U10158 ( .B1(n8787), .B2(n7043), .A(n8786), .ZN(n8788) );
  OAI211_X1 U10159 ( .C1(n8913), .C2(n8790), .A(n8789), .B(n8788), .ZN(
        P2_U3280) );
  OAI21_X1 U10160 ( .B1(n8792), .B2(n8799), .A(n8791), .ZN(n8793) );
  INV_X1 U10161 ( .A(n8793), .ZN(n8922) );
  INV_X1 U10162 ( .A(n8794), .ZN(n8795) );
  AOI21_X1 U10163 ( .B1(n8918), .B2(n8796), .A(n8795), .ZN(n8919) );
  AOI22_X1 U10164 ( .A1(n8804), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n8797), .B2(
        n9747), .ZN(n8798) );
  OAI21_X1 U10165 ( .B1(n4538), .B2(n8821), .A(n8798), .ZN(n8806) );
  XNOR2_X1 U10166 ( .A(n8800), .B(n8799), .ZN(n8803) );
  AOI222_X1 U10167 ( .A1(n8813), .A2(n8803), .B1(n8802), .B2(n9743), .C1(n8801), .C2(n9744), .ZN(n8921) );
  NOR2_X1 U10168 ( .A1(n8921), .A2(n8804), .ZN(n8805) );
  AOI211_X1 U10169 ( .C1(n8919), .C2(n7043), .A(n8806), .B(n8805), .ZN(n8807)
         );
  OAI21_X1 U10170 ( .B1(n8922), .B2(n8764), .A(n8807), .ZN(P2_U3281) );
  OAI21_X1 U10171 ( .B1(n8819), .B2(n8809), .A(n8808), .ZN(n8812) );
  AOI222_X1 U10172 ( .A1(n8813), .A2(n8812), .B1(n8811), .B2(n9744), .C1(n8810), .C2(n9743), .ZN(n9806) );
  MUX2_X1 U10173 ( .A(n6883), .B(n9806), .S(n8830), .Z(n8825) );
  OR2_X1 U10174 ( .A1(n8814), .A2(n8820), .ZN(n8815) );
  AND2_X1 U10175 ( .A1(n8816), .A2(n8815), .ZN(n9804) );
  AOI22_X1 U10176 ( .A1(n7043), .A2(n9804), .B1(n8817), .B2(n9747), .ZN(n8824)
         );
  XOR2_X1 U10177 ( .A(n8818), .B(n8819), .Z(n9808) );
  NAND2_X1 U10178 ( .A1(n9808), .A2(n9754), .ZN(n8823) );
  OR2_X1 U10179 ( .A1(n8821), .A2(n8820), .ZN(n8822) );
  NAND4_X1 U10180 ( .A1(n8825), .A2(n8824), .A3(n8823), .A4(n8822), .ZN(
        P2_U3290) );
  AOI22_X1 U10181 ( .A1(n9754), .A2(n8828), .B1(n8827), .B2(n8826), .ZN(n8834)
         );
  AOI22_X1 U10182 ( .A1(n7043), .A2(n8829), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n9747), .ZN(n8833) );
  MUX2_X1 U10183 ( .A(n6890), .B(n8831), .S(n8830), .Z(n8832) );
  NAND3_X1 U10184 ( .A1(n8834), .A2(n8833), .A3(n8832), .ZN(P2_U3295) );
  NAND2_X1 U10185 ( .A1(n8835), .A2(n9802), .ZN(n8836) );
  OAI211_X1 U10186 ( .C1(n8837), .C2(n9825), .A(n8840), .B(n8836), .ZN(n8940)
         );
  MUX2_X1 U10187 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n8940), .S(n9848), .Z(
        P2_U3551) );
  NAND2_X1 U10188 ( .A1(n8838), .A2(n9802), .ZN(n8839) );
  OAI211_X1 U10189 ( .C1(n8841), .C2(n9825), .A(n8840), .B(n8839), .ZN(n8941)
         );
  MUX2_X1 U10190 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n8941), .S(n9848), .Z(
        P2_U3550) );
  AOI22_X1 U10191 ( .A1(n8843), .A2(n9803), .B1(n9802), .B2(n8842), .ZN(n8844)
         );
  MUX2_X1 U10192 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n8942), .S(n9848), .Z(
        P2_U3549) );
  AOI22_X1 U10193 ( .A1(n8848), .A2(n9803), .B1(n9802), .B2(n8847), .ZN(n8849)
         );
  OAI211_X1 U10194 ( .C1(n8851), .C2(n9797), .A(n8850), .B(n8849), .ZN(n8943)
         );
  MUX2_X1 U10195 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n8943), .S(n9848), .Z(
        P2_U3548) );
  AOI22_X1 U10196 ( .A1(n8853), .A2(n9803), .B1(n9802), .B2(n8852), .ZN(n8854)
         );
  OAI211_X1 U10197 ( .C1(n8856), .C2(n9797), .A(n8855), .B(n8854), .ZN(n8944)
         );
  MUX2_X1 U10198 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8944), .S(n9848), .Z(
        P2_U3547) );
  AOI21_X1 U10199 ( .B1(n9802), .B2(n8858), .A(n8857), .ZN(n8859) );
  OAI211_X1 U10200 ( .C1(n8861), .C2(n9797), .A(n8860), .B(n8859), .ZN(n8945)
         );
  MUX2_X1 U10201 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n8945), .S(n9848), .Z(
        P2_U3546) );
  AOI21_X1 U10202 ( .B1(n9802), .B2(n8863), .A(n8862), .ZN(n8864) );
  OAI211_X1 U10203 ( .C1(n8866), .C2(n9797), .A(n8865), .B(n8864), .ZN(n8946)
         );
  MUX2_X1 U10204 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8946), .S(n9848), .Z(
        P2_U3545) );
  AOI22_X1 U10205 ( .A1(n8868), .A2(n9803), .B1(n9802), .B2(n8867), .ZN(n8869)
         );
  OAI211_X1 U10206 ( .C1(n8871), .C2(n9797), .A(n8870), .B(n8869), .ZN(n8947)
         );
  MUX2_X1 U10207 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8947), .S(n9848), .Z(
        P2_U3544) );
  INV_X1 U10208 ( .A(n9797), .ZN(n9829) );
  NAND2_X1 U10209 ( .A1(n8872), .A2(n9829), .ZN(n8877) );
  AOI22_X1 U10210 ( .A1(n8874), .A2(n9803), .B1(n9802), .B2(n8873), .ZN(n8875)
         );
  OAI211_X1 U10211 ( .C1(n8878), .C2(n8877), .A(n8876), .B(n8875), .ZN(n8948)
         );
  MUX2_X1 U10212 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8948), .S(n9848), .Z(
        P2_U3543) );
  AOI22_X1 U10213 ( .A1(n8880), .A2(n9803), .B1(n9802), .B2(n8879), .ZN(n8881)
         );
  OAI211_X1 U10214 ( .C1(n8883), .C2(n9797), .A(n8882), .B(n8881), .ZN(n8949)
         );
  MUX2_X1 U10215 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n8949), .S(n9848), .Z(
        P2_U3542) );
  AOI22_X1 U10216 ( .A1(n8885), .A2(n9803), .B1(n9802), .B2(n8884), .ZN(n8886)
         );
  OAI211_X1 U10217 ( .C1(n8888), .C2(n9797), .A(n8887), .B(n8886), .ZN(n8950)
         );
  MUX2_X1 U10218 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n8950), .S(n9848), .Z(
        P2_U3541) );
  AOI22_X1 U10219 ( .A1(n8890), .A2(n9803), .B1(n9802), .B2(n8889), .ZN(n8891)
         );
  OAI211_X1 U10220 ( .C1(n8893), .C2(n9797), .A(n8892), .B(n8891), .ZN(n8951)
         );
  MUX2_X1 U10221 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n8951), .S(n9848), .Z(
        P2_U3540) );
  AOI211_X1 U10222 ( .C1(n9802), .C2(n8896), .A(n8895), .B(n8894), .ZN(n8897)
         );
  OAI21_X1 U10223 ( .B1(n8898), .B2(n9797), .A(n8897), .ZN(n8952) );
  MUX2_X1 U10224 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8952), .S(n9848), .Z(
        P2_U3539) );
  AOI22_X1 U10225 ( .A1(n8900), .A2(n9803), .B1(n9802), .B2(n8899), .ZN(n8901)
         );
  OAI211_X1 U10226 ( .C1(n8903), .C2(n9797), .A(n8902), .B(n8901), .ZN(n8953)
         );
  MUX2_X1 U10227 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n8953), .S(n9848), .Z(
        P2_U3538) );
  AOI21_X1 U10228 ( .B1(n9802), .B2(n8905), .A(n8904), .ZN(n8906) );
  OAI211_X1 U10229 ( .C1(n8908), .C2(n9797), .A(n8907), .B(n8906), .ZN(n8954)
         );
  MUX2_X1 U10230 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8954), .S(n9848), .Z(
        P2_U3537) );
  INV_X1 U10231 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8916) );
  INV_X1 U10232 ( .A(n9802), .ZN(n9824) );
  OAI22_X1 U10233 ( .A1(n8910), .A2(n9825), .B1(n8909), .B2(n9824), .ZN(n8911)
         );
  INV_X1 U10234 ( .A(n8911), .ZN(n8912) );
  OAI21_X1 U10235 ( .B1(n8913), .B2(n9809), .A(n8912), .ZN(n8914) );
  NOR2_X1 U10236 ( .A1(n8915), .A2(n8914), .ZN(n8955) );
  MUX2_X1 U10237 ( .A(n8916), .B(n8955), .S(n9848), .Z(n8917) );
  INV_X1 U10238 ( .A(n8917), .ZN(P2_U3536) );
  AOI22_X1 U10239 ( .A1(n8919), .A2(n9803), .B1(n9802), .B2(n8918), .ZN(n8920)
         );
  OAI211_X1 U10240 ( .C1(n8922), .C2(n9797), .A(n8921), .B(n8920), .ZN(n8958)
         );
  MUX2_X1 U10241 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n8958), .S(n9848), .Z(
        P2_U3535) );
  AOI211_X1 U10242 ( .C1(n9802), .C2(n8925), .A(n8924), .B(n8923), .ZN(n8926)
         );
  OAI21_X1 U10243 ( .B1(n9797), .B2(n8927), .A(n8926), .ZN(n8959) );
  MUX2_X1 U10244 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n8959), .S(n9848), .Z(
        P2_U3534) );
  INV_X1 U10245 ( .A(n9809), .ZN(n9822) );
  OAI22_X1 U10246 ( .A1(n8929), .A2(n9825), .B1(n8928), .B2(n9824), .ZN(n8930)
         );
  AOI21_X1 U10247 ( .B1(n8931), .B2(n9822), .A(n8930), .ZN(n8932) );
  NAND2_X1 U10248 ( .A1(n8933), .A2(n8932), .ZN(n8960) );
  MUX2_X1 U10249 ( .A(n8960), .B(P2_REG1_REG_13__SCAN_IN), .S(n9846), .Z(
        P2_U3533) );
  AOI22_X1 U10250 ( .A1(n8935), .A2(n9803), .B1(n9802), .B2(n8934), .ZN(n8936)
         );
  OAI211_X1 U10251 ( .C1(n9797), .C2(n8938), .A(n8937), .B(n8936), .ZN(n8961)
         );
  MUX2_X1 U10252 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n8961), .S(n9848), .Z(
        P2_U3531) );
  MUX2_X1 U10253 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n8939), .S(n9848), .Z(
        P2_U3521) );
  MUX2_X1 U10254 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n8940), .S(n9833), .Z(
        P2_U3519) );
  MUX2_X1 U10255 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n8941), .S(n9833), .Z(
        P2_U3518) );
  MUX2_X1 U10256 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n8942), .S(n9833), .Z(
        P2_U3517) );
  MUX2_X1 U10257 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n8943), .S(n9833), .Z(
        P2_U3516) );
  MUX2_X1 U10258 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8944), .S(n9833), .Z(
        P2_U3515) );
  MUX2_X1 U10259 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n8945), .S(n9833), .Z(
        P2_U3514) );
  MUX2_X1 U10260 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n8946), .S(n9833), .Z(
        P2_U3513) );
  MUX2_X1 U10261 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n8947), .S(n9833), .Z(
        P2_U3512) );
  MUX2_X1 U10262 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n8948), .S(n9833), .Z(
        P2_U3511) );
  MUX2_X1 U10263 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n8949), .S(n9833), .Z(
        P2_U3510) );
  MUX2_X1 U10264 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n8950), .S(n9833), .Z(
        P2_U3509) );
  MUX2_X1 U10265 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n8951), .S(n9833), .Z(
        P2_U3508) );
  MUX2_X1 U10266 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n8952), .S(n9833), .Z(
        P2_U3507) );
  MUX2_X1 U10267 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n8953), .S(n9833), .Z(
        P2_U3505) );
  MUX2_X1 U10268 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n8954), .S(n9833), .Z(
        P2_U3502) );
  INV_X1 U10269 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n8956) );
  MUX2_X1 U10270 ( .A(n8956), .B(n8955), .S(n9833), .Z(n8957) );
  INV_X1 U10271 ( .A(n8957), .ZN(P2_U3499) );
  MUX2_X1 U10272 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n8958), .S(n9833), .Z(
        P2_U3496) );
  MUX2_X1 U10273 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n8959), .S(n9833), .Z(
        P2_U3493) );
  MUX2_X1 U10274 ( .A(n8960), .B(P2_REG0_REG_13__SCAN_IN), .S(n9831), .Z(
        P2_U3490) );
  MUX2_X1 U10275 ( .A(P2_REG0_REG_11__SCAN_IN), .B(n8961), .S(n9833), .Z(
        P2_U3484) );
  NOR4_X1 U10276 ( .A1(n4324), .A2(P2_IR_REG_30__SCAN_IN), .A3(n8962), .A4(
        P2_U3152), .ZN(n8963) );
  AOI21_X1 U10277 ( .B1(n8969), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n8963), .ZN(
        n8964) );
  OAI21_X1 U10278 ( .B1(n9509), .B2(n8967), .A(n8964), .ZN(P2_U3327) );
  AOI22_X1 U10279 ( .A1(n8965), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n8969), .ZN(n8966) );
  OAI21_X1 U10280 ( .B1(n8968), .B2(n8967), .A(n8966), .ZN(P2_U3328) );
  AOI22_X1 U10281 ( .A1(n8970), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n8969), .ZN(n8971) );
  OAI21_X1 U10282 ( .B1(n8972), .B2(n8967), .A(n8971), .ZN(P2_U3329) );
  MUX2_X1 U10283 ( .A(n8973), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  XNOR2_X1 U10284 ( .A(n8975), .B(n8974), .ZN(n8976) );
  XNOR2_X1 U10285 ( .A(n8977), .B(n8976), .ZN(n8983) );
  OAI22_X1 U10286 ( .A1(n9230), .A2(n9092), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8978), .ZN(n8979) );
  AOI21_X1 U10287 ( .B1(n9226), .B2(n9106), .A(n8979), .ZN(n8980) );
  OAI21_X1 U10288 ( .B1(n9231), .B2(n9109), .A(n8980), .ZN(n8981) );
  AOI21_X1 U10289 ( .B1(n9420), .B2(n9112), .A(n8981), .ZN(n8982) );
  OAI21_X1 U10290 ( .B1(n8983), .B2(n9115), .A(n8982), .ZN(P1_U3212) );
  INV_X1 U10291 ( .A(n8984), .ZN(n8986) );
  NAND2_X1 U10292 ( .A1(n8986), .A2(n8985), .ZN(n8988) );
  XNOR2_X1 U10293 ( .A(n8988), .B(n8987), .ZN(n8994) );
  OAI22_X1 U10294 ( .A1(n9332), .A2(n9092), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8989), .ZN(n8990) );
  AOI21_X1 U10295 ( .B1(n9094), .B2(n9265), .A(n8990), .ZN(n8991) );
  OAI21_X1 U10296 ( .B1(n9071), .B2(n9294), .A(n8991), .ZN(n8992) );
  AOI21_X1 U10297 ( .B1(n9441), .B2(n9112), .A(n8992), .ZN(n8993) );
  OAI21_X1 U10298 ( .B1(n8994), .B2(n9115), .A(n8993), .ZN(P1_U3214) );
  NAND2_X1 U10299 ( .A1(n8996), .A2(n8995), .ZN(n8998) );
  XOR2_X1 U10300 ( .A(n8998), .B(n8997), .Z(n9003) );
  NAND2_X1 U10301 ( .A1(n9094), .A2(n9369), .ZN(n8999) );
  NAND2_X1 U10302 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9174) );
  OAI211_X1 U10303 ( .C1(n9037), .C2(n9092), .A(n8999), .B(n9174), .ZN(n9001)
         );
  NOR2_X1 U10304 ( .A1(n9363), .A2(n9097), .ZN(n9000) );
  AOI211_X1 U10305 ( .C1(n9361), .C2(n9106), .A(n9001), .B(n9000), .ZN(n9002)
         );
  OAI21_X1 U10306 ( .B1(n9003), .B2(n9115), .A(n9002), .ZN(P1_U3217) );
  NOR2_X1 U10307 ( .A1(n4377), .A2(n9005), .ZN(n9006) );
  XNOR2_X1 U10308 ( .A(n9004), .B(n9006), .ZN(n9011) );
  AOI22_X1 U10309 ( .A1(n9118), .A2(n9094), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3084), .ZN(n9008) );
  NAND2_X1 U10310 ( .A1(n9104), .A2(n9369), .ZN(n9007) );
  OAI211_X1 U10311 ( .C1(n9071), .C2(n9336), .A(n9008), .B(n9007), .ZN(n9009)
         );
  AOI21_X1 U10312 ( .B1(n9452), .B2(n9112), .A(n9009), .ZN(n9010) );
  OAI21_X1 U10313 ( .B1(n9011), .B2(n9115), .A(n9010), .ZN(P1_U3221) );
  XOR2_X1 U10314 ( .A(n9013), .B(n9012), .Z(n9018) );
  NAND2_X1 U10315 ( .A1(n9264), .A2(n9094), .ZN(n9015) );
  AOI22_X1 U10316 ( .A1(n9265), .A2(n9104), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3084), .ZN(n9014) );
  OAI211_X1 U10317 ( .C1(n9071), .C2(n9256), .A(n9015), .B(n9014), .ZN(n9016)
         );
  AOI21_X1 U10318 ( .B1(n9429), .B2(n9112), .A(n9016), .ZN(n9017) );
  OAI21_X1 U10319 ( .B1(n9018), .B2(n9115), .A(n9017), .ZN(P1_U3223) );
  INV_X1 U10320 ( .A(n9019), .ZN(n9023) );
  AOI21_X1 U10321 ( .B1(n9021), .B2(n9099), .A(n9020), .ZN(n9022) );
  OAI21_X1 U10322 ( .B1(n9023), .B2(n9022), .A(n9087), .ZN(n9031) );
  INV_X1 U10323 ( .A(n9024), .ZN(n9025) );
  AOI21_X1 U10324 ( .B1(n9104), .B2(n9119), .A(n9025), .ZN(n9026) );
  OAI21_X1 U10325 ( .B1(n9027), .B2(n9109), .A(n9026), .ZN(n9028) );
  AOI21_X1 U10326 ( .B1(n9029), .B2(n9106), .A(n9028), .ZN(n9030) );
  OAI211_X1 U10327 ( .C1(n4600), .C2(n9097), .A(n9031), .B(n9030), .ZN(
        P1_U3224) );
  OAI21_X1 U10328 ( .B1(n9034), .B2(n9032), .A(n9033), .ZN(n9035) );
  NAND2_X1 U10329 ( .A1(n9035), .A2(n9087), .ZN(n9040) );
  NAND2_X1 U10330 ( .A1(n9104), .A2(n9402), .ZN(n9036) );
  NAND2_X1 U10331 ( .A1(P1_U3084), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9162) );
  OAI211_X1 U10332 ( .C1(n9037), .C2(n9109), .A(n9036), .B(n9162), .ZN(n9038)
         );
  AOI21_X1 U10333 ( .B1(n9394), .B2(n9106), .A(n9038), .ZN(n9039) );
  OAI211_X1 U10334 ( .C1(n4599), .C2(n9097), .A(n9040), .B(n9039), .ZN(
        P1_U3226) );
  XOR2_X1 U10335 ( .A(n9042), .B(n9041), .Z(n9049) );
  NAND2_X1 U10336 ( .A1(n9308), .A2(n9104), .ZN(n9043) );
  OAI21_X1 U10337 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n9044), .A(n9043), .ZN(
        n9045) );
  AOI21_X1 U10338 ( .B1(n9280), .B2(n9106), .A(n9045), .ZN(n9046) );
  OAI21_X1 U10339 ( .B1(n9278), .B2(n9109), .A(n9046), .ZN(n9047) );
  AOI21_X1 U10340 ( .B1(n9436), .B2(n9112), .A(n9047), .ZN(n9048) );
  OAI21_X1 U10341 ( .B1(n9049), .B2(n9115), .A(n9048), .ZN(P1_U3227) );
  XNOR2_X1 U10342 ( .A(n9052), .B(n9051), .ZN(n9053) );
  XNOR2_X1 U10343 ( .A(n9050), .B(n9053), .ZN(n9060) );
  OAI22_X1 U10344 ( .A1(n9055), .A2(n9109), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9054), .ZN(n9056) );
  AOI21_X1 U10345 ( .B1(n9104), .B2(n9383), .A(n9056), .ZN(n9057) );
  OAI21_X1 U10346 ( .B1(n9071), .B2(n9346), .A(n9057), .ZN(n9058) );
  AOI21_X1 U10347 ( .B1(n9455), .B2(n9112), .A(n9058), .ZN(n9059) );
  OAI21_X1 U10348 ( .B1(n9060), .B2(n9115), .A(n9059), .ZN(P1_U3231) );
  INV_X1 U10349 ( .A(n9061), .ZN(n9063) );
  INV_X1 U10350 ( .A(n9065), .ZN(n9062) );
  OAI21_X1 U10351 ( .B1(n9066), .B2(n9063), .A(n9062), .ZN(n9068) );
  INV_X1 U10352 ( .A(n9064), .ZN(n9067) );
  AOI22_X1 U10353 ( .A1(n9068), .A2(n9067), .B1(n9066), .B2(n9065), .ZN(n9074)
         );
  AOI22_X1 U10354 ( .A1(n9308), .A2(n9094), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3084), .ZN(n9070) );
  NAND2_X1 U10355 ( .A1(n9352), .A2(n9104), .ZN(n9069) );
  OAI211_X1 U10356 ( .C1(n9071), .C2(n9314), .A(n9070), .B(n9069), .ZN(n9072)
         );
  AOI21_X1 U10357 ( .B1(n9317), .B2(n9112), .A(n9072), .ZN(n9073) );
  OAI21_X1 U10358 ( .B1(n9074), .B2(n9115), .A(n9073), .ZN(P1_U3233) );
  INV_X1 U10359 ( .A(n9465), .ZN(n9378) );
  INV_X1 U10360 ( .A(n9077), .ZN(n9081) );
  AOI21_X1 U10361 ( .B1(n9077), .B2(n9076), .A(n9075), .ZN(n9078) );
  NOR2_X1 U10362 ( .A1(n9078), .A2(n9115), .ZN(n9079) );
  OAI21_X1 U10363 ( .B1(n9081), .B2(n9080), .A(n9079), .ZN(n9086) );
  AOI22_X1 U10364 ( .A1(n9104), .A2(n9384), .B1(P1_REG3_REG_18__SCAN_IN), .B2(
        P1_U3084), .ZN(n9082) );
  OAI21_X1 U10365 ( .B1(n9083), .B2(n9109), .A(n9082), .ZN(n9084) );
  AOI21_X1 U10366 ( .B1(n9376), .B2(n9106), .A(n9084), .ZN(n9085) );
  OAI211_X1 U10367 ( .C1(n9378), .C2(n9097), .A(n9086), .B(n9085), .ZN(
        P1_U3236) );
  INV_X1 U10368 ( .A(n9090), .ZN(n9241) );
  AOI22_X1 U10369 ( .A1(n9241), .A2(n9106), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3084), .ZN(n9091) );
  OAI21_X1 U10370 ( .B1(n9278), .B2(n9092), .A(n9091), .ZN(n9093) );
  AOI21_X1 U10371 ( .B1(n9249), .B2(n9094), .A(n9093), .ZN(n9095) );
  OAI211_X1 U10372 ( .C1(n9243), .C2(n9097), .A(n9096), .B(n9095), .ZN(
        P1_U3238) );
  NAND2_X1 U10373 ( .A1(n9099), .A2(n9098), .ZN(n9100) );
  XOR2_X1 U10374 ( .A(n9101), .B(n9100), .Z(n9116) );
  INV_X1 U10375 ( .A(n9102), .ZN(n9103) );
  AOI21_X1 U10376 ( .B1(n9104), .B2(n9120), .A(n9103), .ZN(n9108) );
  NAND2_X1 U10377 ( .A1(n9106), .A2(n9105), .ZN(n9107) );
  OAI211_X1 U10378 ( .C1(n9110), .C2(n9109), .A(n9108), .B(n9107), .ZN(n9111)
         );
  AOI21_X1 U10379 ( .B1(n9113), .B2(n9112), .A(n9111), .ZN(n9114) );
  OAI21_X1 U10380 ( .B1(n9116), .B2(n9115), .A(n9114), .ZN(P1_U3239) );
  MUX2_X1 U10381 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n9195), .S(P1_U4006), .Z(
        P1_U3586) );
  MUX2_X1 U10382 ( .A(n9117), .B(P1_DATAO_REG_30__SCAN_IN), .S(n9134), .Z(
        P1_U3585) );
  MUX2_X1 U10383 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n7960), .S(P1_U4006), .Z(
        P1_U3583) );
  MUX2_X1 U10384 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9249), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U10385 ( .A(n9264), .B(P1_DATAO_REG_26__SCAN_IN), .S(n9134), .Z(
        P1_U3581) );
  MUX2_X1 U10386 ( .A(n9248), .B(P1_DATAO_REG_25__SCAN_IN), .S(n9134), .Z(
        P1_U3580) );
  MUX2_X1 U10387 ( .A(n9265), .B(P1_DATAO_REG_24__SCAN_IN), .S(n9134), .Z(
        P1_U3579) );
  MUX2_X1 U10388 ( .A(n9308), .B(P1_DATAO_REG_23__SCAN_IN), .S(n9134), .Z(
        P1_U3578) );
  MUX2_X1 U10389 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9118), .S(P1_U4006), .Z(
        P1_U3577) );
  MUX2_X1 U10390 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9352), .S(P1_U4006), .Z(
        P1_U3576) );
  MUX2_X1 U10391 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9369), .S(P1_U4006), .Z(
        P1_U3575) );
  MUX2_X1 U10392 ( .A(n9383), .B(P1_DATAO_REG_19__SCAN_IN), .S(n9134), .Z(
        P1_U3574) );
  MUX2_X1 U10393 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9404), .S(P1_U4006), .Z(
        P1_U3573) );
  MUX2_X1 U10394 ( .A(n9384), .B(P1_DATAO_REG_17__SCAN_IN), .S(n9134), .Z(
        P1_U3572) );
  MUX2_X1 U10395 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9402), .S(P1_U4006), .Z(
        P1_U3571) );
  MUX2_X1 U10396 ( .A(n9119), .B(P1_DATAO_REG_15__SCAN_IN), .S(n9134), .Z(
        P1_U3570) );
  MUX2_X1 U10397 ( .A(n9120), .B(P1_DATAO_REG_14__SCAN_IN), .S(n9134), .Z(
        P1_U3569) );
  MUX2_X1 U10398 ( .A(n9121), .B(P1_DATAO_REG_13__SCAN_IN), .S(n9134), .Z(
        P1_U3568) );
  MUX2_X1 U10399 ( .A(n9122), .B(P1_DATAO_REG_12__SCAN_IN), .S(n9134), .Z(
        P1_U3567) );
  MUX2_X1 U10400 ( .A(n9123), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9134), .Z(
        P1_U3566) );
  MUX2_X1 U10401 ( .A(n9124), .B(P1_DATAO_REG_10__SCAN_IN), .S(n9134), .Z(
        P1_U3565) );
  MUX2_X1 U10402 ( .A(n9125), .B(P1_DATAO_REG_9__SCAN_IN), .S(n9134), .Z(
        P1_U3564) );
  MUX2_X1 U10403 ( .A(n9126), .B(P1_DATAO_REG_8__SCAN_IN), .S(n9134), .Z(
        P1_U3563) );
  MUX2_X1 U10404 ( .A(n9127), .B(P1_DATAO_REG_7__SCAN_IN), .S(n9134), .Z(
        P1_U3562) );
  MUX2_X1 U10405 ( .A(n9128), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9134), .Z(
        P1_U3561) );
  MUX2_X1 U10406 ( .A(n9129), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9134), .Z(
        P1_U3560) );
  MUX2_X1 U10407 ( .A(n9130), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9134), .Z(
        P1_U3559) );
  MUX2_X1 U10408 ( .A(n9131), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9134), .Z(
        P1_U3558) );
  MUX2_X1 U10409 ( .A(n9132), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9134), .Z(
        P1_U3557) );
  MUX2_X1 U10410 ( .A(n9133), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9134), .Z(
        P1_U3556) );
  MUX2_X1 U10411 ( .A(n6306), .B(P1_DATAO_REG_0__SCAN_IN), .S(n9134), .Z(
        P1_U3555) );
  NAND2_X1 U10412 ( .A1(P1_REG3_REG_1__SCAN_IN), .A2(P1_U3084), .ZN(n9135) );
  OAI21_X1 U10413 ( .B1(n9646), .B2(n9136), .A(n9135), .ZN(n9137) );
  AOI21_X1 U10414 ( .B1(n9648), .B2(P1_ADDR_REG_1__SCAN_IN), .A(n9137), .ZN(
        n9146) );
  OAI211_X1 U10415 ( .C1(n9140), .C2(n9139), .A(n9672), .B(n9138), .ZN(n9145)
         );
  OAI211_X1 U10416 ( .C1(n9143), .C2(n9142), .A(n9673), .B(n9141), .ZN(n9144)
         );
  NAND3_X1 U10417 ( .A1(n9146), .A2(n9145), .A3(n9144), .ZN(P1_U3242) );
  OAI21_X1 U10418 ( .B1(n9646), .B2(n9148), .A(n9147), .ZN(n9149) );
  AOI21_X1 U10419 ( .B1(n9648), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n9149), .ZN(
        n9160) );
  MUX2_X1 U10420 ( .A(n6555), .B(P1_REG2_REG_3__SCAN_IN), .S(n9150), .Z(n9151)
         );
  NAND3_X1 U10421 ( .A1(n9612), .A2(n9152), .A3(n9151), .ZN(n9153) );
  NAND3_X1 U10422 ( .A1(n9673), .A2(n9154), .A3(n9153), .ZN(n9159) );
  OAI211_X1 U10423 ( .C1(n9157), .C2(n9156), .A(n9672), .B(n9155), .ZN(n9158)
         );
  NAND3_X1 U10424 ( .A1(n9160), .A2(n9159), .A3(n9158), .ZN(P1_U3244) );
  INV_X1 U10425 ( .A(n9161), .ZN(n9163) );
  OAI21_X1 U10426 ( .B1(n9646), .B2(n9163), .A(n9162), .ZN(n9164) );
  AOI21_X1 U10427 ( .B1(n9648), .B2(P1_ADDR_REG_17__SCAN_IN), .A(n9164), .ZN(
        n9173) );
  OAI211_X1 U10428 ( .C1(n9167), .C2(n9166), .A(n9673), .B(n9165), .ZN(n9172)
         );
  OAI211_X1 U10429 ( .C1(n9170), .C2(n9169), .A(n9672), .B(n9168), .ZN(n9171)
         );
  NAND3_X1 U10430 ( .A1(n9173), .A2(n9172), .A3(n9171), .ZN(P1_U3258) );
  INV_X1 U10431 ( .A(n9174), .ZN(n9190) );
  OR2_X1 U10432 ( .A1(n9175), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9176) );
  NAND2_X1 U10433 ( .A1(n9177), .A2(n9176), .ZN(n9178) );
  XNOR2_X1 U10434 ( .A(n9178), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n9186) );
  INV_X1 U10435 ( .A(n9186), .ZN(n9183) );
  NAND2_X1 U10436 ( .A1(n9180), .A2(n9179), .ZN(n9181) );
  XNOR2_X1 U10437 ( .A(n9181), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n9184) );
  OAI22_X1 U10438 ( .A1(n9634), .A2(n9183), .B1(n9182), .B2(n9184), .ZN(n9188)
         );
  NAND2_X1 U10439 ( .A1(n9643), .A2(n9184), .ZN(n9185) );
  OAI211_X1 U10440 ( .C1(n9634), .C2(n9186), .A(n9646), .B(n9185), .ZN(n9187)
         );
  MUX2_X1 U10441 ( .A(n9188), .B(n9187), .S(n9282), .Z(n9189) );
  AOI211_X1 U10442 ( .C1(P1_ADDR_REG_19__SCAN_IN), .C2(n9648), .A(n9190), .B(
        n9189), .ZN(n9191) );
  INV_X1 U10443 ( .A(n9191), .ZN(P1_U3260) );
  INV_X1 U10444 ( .A(n9193), .ZN(n9549) );
  NAND2_X1 U10445 ( .A1(n9556), .A2(n9199), .ZN(n9192) );
  XOR2_X1 U10446 ( .A(n9193), .B(n9192), .Z(n9551) );
  NAND2_X1 U10447 ( .A1(n9551), .A2(n9409), .ZN(n9197) );
  NAND2_X1 U10448 ( .A1(n9195), .A2(n9194), .ZN(n9555) );
  NOR2_X1 U10449 ( .A1(n6638), .A2(n9555), .ZN(n9200) );
  AOI21_X1 U10450 ( .B1(n6638), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9200), .ZN(
        n9196) );
  OAI211_X1 U10451 ( .C1(n9549), .C2(n9396), .A(n9197), .B(n9196), .ZN(
        P1_U3261) );
  XNOR2_X1 U10452 ( .A(n9199), .B(n9198), .ZN(n9558) );
  NAND2_X1 U10453 ( .A1(n9558), .A2(n9409), .ZN(n9202) );
  AOI21_X1 U10454 ( .B1(n6638), .B2(P1_REG2_REG_30__SCAN_IN), .A(n9200), .ZN(
        n9201) );
  OAI211_X1 U10455 ( .C1(n9556), .C2(n9396), .A(n9202), .B(n9201), .ZN(
        P1_U3262) );
  NAND2_X1 U10456 ( .A1(n9204), .A2(n9203), .ZN(n9205) );
  INV_X1 U10457 ( .A(n9416), .ZN(n9221) );
  AND2_X1 U10458 ( .A1(n9207), .A2(n4826), .ZN(n9208) );
  OAI21_X1 U10459 ( .B1(n4346), .B2(n9208), .A(n9406), .ZN(n9213) );
  OAI22_X1 U10460 ( .A1(n9210), .A2(n9331), .B1(n9209), .B2(n9333), .ZN(n9211)
         );
  INV_X1 U10461 ( .A(n9211), .ZN(n9212) );
  NAND2_X1 U10462 ( .A1(n9213), .A2(n9212), .ZN(n9414) );
  NAND2_X1 U10463 ( .A1(n9223), .A2(n9214), .ZN(n9215) );
  NAND2_X1 U10464 ( .A1(n4341), .A2(n9215), .ZN(n9412) );
  NOR2_X1 U10465 ( .A1(n9412), .A2(n9319), .ZN(n9219) );
  AOI22_X1 U10466 ( .A1(n9216), .A2(n9393), .B1(P1_REG2_REG_28__SCAN_IN), .B2(
        n6638), .ZN(n9217) );
  OAI21_X1 U10467 ( .B1(n4596), .B2(n9396), .A(n9217), .ZN(n9218) );
  AOI211_X1 U10468 ( .C1(n9414), .C2(n9688), .A(n9219), .B(n9218), .ZN(n9220)
         );
  OAI21_X1 U10469 ( .B1(n9221), .B2(n9411), .A(n9220), .ZN(P1_U3263) );
  XNOR2_X1 U10470 ( .A(n9222), .B(n9228), .ZN(n9423) );
  INV_X1 U10471 ( .A(n9239), .ZN(n9225) );
  INV_X1 U10472 ( .A(n9223), .ZN(n9224) );
  AOI211_X1 U10473 ( .C1(n9420), .C2(n9225), .A(n9707), .B(n9224), .ZN(n9419)
         );
  AOI22_X1 U10474 ( .A1(n9226), .A2(n9393), .B1(P1_REG2_REG_27__SCAN_IN), .B2(
        n6638), .ZN(n9227) );
  OAI21_X1 U10475 ( .B1(n4828), .B2(n9396), .A(n9227), .ZN(n9236) );
  AOI21_X1 U10476 ( .B1(n9229), .B2(n9228), .A(n9329), .ZN(n9234) );
  OAI22_X1 U10477 ( .A1(n9231), .A2(n9333), .B1(n9230), .B2(n9331), .ZN(n9232)
         );
  AOI21_X1 U10478 ( .B1(n9234), .B2(n9233), .A(n9232), .ZN(n9422) );
  NOR2_X1 U10479 ( .A1(n9422), .A2(n6638), .ZN(n9235) );
  AOI211_X1 U10480 ( .C1(n9419), .C2(n9335), .A(n9236), .B(n9235), .ZN(n9237)
         );
  OAI21_X1 U10481 ( .B1(n9423), .B2(n9411), .A(n9237), .ZN(P1_U3264) );
  XNOR2_X1 U10482 ( .A(n9238), .B(n9247), .ZN(n9428) );
  INV_X1 U10483 ( .A(n9255), .ZN(n9240) );
  AOI21_X1 U10484 ( .B1(n9424), .B2(n9240), .A(n9239), .ZN(n9425) );
  AOI22_X1 U10485 ( .A1(n9241), .A2(n9393), .B1(P1_REG2_REG_26__SCAN_IN), .B2(
        n6638), .ZN(n9242) );
  OAI21_X1 U10486 ( .B1(n9243), .B2(n9396), .A(n9242), .ZN(n9252) );
  NAND2_X1 U10487 ( .A1(n9245), .A2(n9244), .ZN(n9246) );
  XOR2_X1 U10488 ( .A(n9247), .B(n9246), .Z(n9250) );
  AOI222_X1 U10489 ( .A1(n9406), .A2(n9250), .B1(n9249), .B2(n9403), .C1(n9248), .C2(n9401), .ZN(n9427) );
  NOR2_X1 U10490 ( .A1(n9427), .A2(n6638), .ZN(n9251) );
  AOI211_X1 U10491 ( .C1(n9425), .C2(n9409), .A(n9252), .B(n9251), .ZN(n9253)
         );
  OAI21_X1 U10492 ( .B1(n9428), .B2(n9411), .A(n9253), .ZN(P1_U3265) );
  XOR2_X1 U10493 ( .A(n9254), .B(n9263), .Z(n9433) );
  AOI21_X1 U10494 ( .B1(n9429), .B2(n9279), .A(n9255), .ZN(n9430) );
  INV_X1 U10495 ( .A(n9429), .ZN(n9259) );
  INV_X1 U10496 ( .A(n9256), .ZN(n9257) );
  AOI22_X1 U10497 ( .A1(n9257), .A2(n9393), .B1(P1_REG2_REG_25__SCAN_IN), .B2(
        n6638), .ZN(n9258) );
  OAI21_X1 U10498 ( .B1(n9259), .B2(n9396), .A(n9258), .ZN(n9268) );
  NAND2_X1 U10499 ( .A1(n9261), .A2(n9260), .ZN(n9262) );
  XOR2_X1 U10500 ( .A(n9263), .B(n9262), .Z(n9266) );
  AOI222_X1 U10501 ( .A1(n9406), .A2(n9266), .B1(n9265), .B2(n9401), .C1(n9264), .C2(n9403), .ZN(n9432) );
  NOR2_X1 U10502 ( .A1(n9432), .A2(n6638), .ZN(n9267) );
  AOI211_X1 U10503 ( .C1(n9430), .C2(n9409), .A(n9268), .B(n9267), .ZN(n9269)
         );
  OAI21_X1 U10504 ( .B1(n9433), .B2(n9411), .A(n9269), .ZN(P1_U3266) );
  XNOR2_X1 U10505 ( .A(n9270), .B(n9271), .ZN(n9438) );
  AOI22_X1 U10506 ( .A1(n9436), .A2(n9316), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n6638), .ZN(n9286) );
  NAND2_X1 U10507 ( .A1(n9273), .A2(n9272), .ZN(n9275) );
  XNOR2_X1 U10508 ( .A(n9275), .B(n9274), .ZN(n9276) );
  OAI222_X1 U10509 ( .A1(n9333), .A2(n9278), .B1(n9331), .B2(n9277), .C1(n9329), .C2(n9276), .ZN(n9434) );
  AOI211_X1 U10510 ( .C1(n9436), .C2(n9292), .A(n9707), .B(n4607), .ZN(n9435)
         );
  INV_X1 U10511 ( .A(n9435), .ZN(n9283) );
  INV_X1 U10512 ( .A(n9280), .ZN(n9281) );
  OAI22_X1 U10513 ( .A1(n9283), .A2(n9282), .B1(n9692), .B2(n9281), .ZN(n9284)
         );
  OAI21_X1 U10514 ( .B1(n9434), .B2(n9284), .A(n9688), .ZN(n9285) );
  OAI211_X1 U10515 ( .C1(n9438), .C2(n9411), .A(n9286), .B(n9285), .ZN(
        P1_U3267) );
  XNOR2_X1 U10516 ( .A(n9287), .B(n9288), .ZN(n9443) );
  XNOR2_X1 U10517 ( .A(n9289), .B(n9288), .ZN(n9290) );
  OAI222_X1 U10518 ( .A1(n9333), .A2(n9291), .B1(n9331), .B2(n9332), .C1(n9290), .C2(n9329), .ZN(n9439) );
  INV_X1 U10519 ( .A(n9312), .ZN(n9293) );
  AOI211_X1 U10520 ( .C1(n9441), .C2(n9293), .A(n9707), .B(n4602), .ZN(n9440)
         );
  NAND2_X1 U10521 ( .A1(n9440), .A2(n9335), .ZN(n9297) );
  INV_X1 U10522 ( .A(n9294), .ZN(n9295) );
  AOI22_X1 U10523 ( .A1(n9295), .A2(n9393), .B1(P1_REG2_REG_23__SCAN_IN), .B2(
        n6638), .ZN(n9296) );
  OAI211_X1 U10524 ( .C1(n9298), .C2(n9396), .A(n9297), .B(n9296), .ZN(n9299)
         );
  AOI21_X1 U10525 ( .B1(n9439), .B2(n9688), .A(n9299), .ZN(n9300) );
  OAI21_X1 U10526 ( .B1(n9443), .B2(n9411), .A(n9300), .ZN(P1_U3268) );
  XNOR2_X1 U10527 ( .A(n9301), .B(n9305), .ZN(n9448) );
  INV_X1 U10528 ( .A(n9448), .ZN(n9323) );
  INV_X1 U10529 ( .A(n9302), .ZN(n9303) );
  AOI21_X1 U10530 ( .B1(n9327), .B2(n9304), .A(n9303), .ZN(n9306) );
  XNOR2_X1 U10531 ( .A(n9306), .B(n9305), .ZN(n9307) );
  NAND2_X1 U10532 ( .A1(n9307), .A2(n9406), .ZN(n9310) );
  AOI22_X1 U10533 ( .A1(n9403), .A2(n9308), .B1(n9352), .B2(n9401), .ZN(n9309)
         );
  NAND2_X1 U10534 ( .A1(n9310), .A2(n9309), .ZN(n9447) );
  NOR2_X1 U10535 ( .A1(n9334), .A2(n9444), .ZN(n9311) );
  OR2_X1 U10536 ( .A1(n9312), .A2(n9311), .ZN(n9445) );
  INV_X1 U10537 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n9313) );
  OAI22_X1 U10538 ( .A1(n9314), .A2(n9692), .B1(n9688), .B2(n9313), .ZN(n9315)
         );
  AOI21_X1 U10539 ( .B1(n9317), .B2(n9316), .A(n9315), .ZN(n9318) );
  OAI21_X1 U10540 ( .B1(n9445), .B2(n9319), .A(n9318), .ZN(n9320) );
  AOI21_X1 U10541 ( .B1(n9447), .B2(n9321), .A(n9320), .ZN(n9322) );
  OAI21_X1 U10542 ( .B1(n9323), .B2(n9411), .A(n9322), .ZN(P1_U3269) );
  XNOR2_X1 U10543 ( .A(n9325), .B(n9324), .ZN(n9454) );
  XNOR2_X1 U10544 ( .A(n9327), .B(n9326), .ZN(n9328) );
  OAI222_X1 U10545 ( .A1(n9333), .A2(n9332), .B1(n9331), .B2(n9330), .C1(n9329), .C2(n9328), .ZN(n9450) );
  INV_X1 U10546 ( .A(n9452), .ZN(n9340) );
  AOI211_X1 U10547 ( .C1(n9452), .C2(n9344), .A(n9707), .B(n9334), .ZN(n9451)
         );
  NAND2_X1 U10548 ( .A1(n9451), .A2(n9335), .ZN(n9339) );
  INV_X1 U10549 ( .A(n9336), .ZN(n9337) );
  AOI22_X1 U10550 ( .A1(n6638), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n9337), .B2(
        n9393), .ZN(n9338) );
  OAI211_X1 U10551 ( .C1(n9340), .C2(n9396), .A(n9339), .B(n9338), .ZN(n9341)
         );
  AOI21_X1 U10552 ( .B1(n9450), .B2(n9688), .A(n9341), .ZN(n9342) );
  OAI21_X1 U10553 ( .B1(n9454), .B2(n9411), .A(n9342), .ZN(P1_U3270) );
  XOR2_X1 U10554 ( .A(n9351), .B(n9343), .Z(n9459) );
  INV_X1 U10555 ( .A(n9344), .ZN(n9345) );
  AOI21_X1 U10556 ( .B1(n9455), .B2(n9358), .A(n9345), .ZN(n9456) );
  INV_X1 U10557 ( .A(n9455), .ZN(n9349) );
  INV_X1 U10558 ( .A(n9346), .ZN(n9347) );
  AOI22_X1 U10559 ( .A1(n6638), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9347), .B2(
        n9393), .ZN(n9348) );
  OAI21_X1 U10560 ( .B1(n9349), .B2(n9396), .A(n9348), .ZN(n9355) );
  XOR2_X1 U10561 ( .A(n9351), .B(n9350), .Z(n9353) );
  AOI222_X1 U10562 ( .A1(n9406), .A2(n9353), .B1(n9383), .B2(n9401), .C1(n9352), .C2(n9403), .ZN(n9458) );
  NOR2_X1 U10563 ( .A1(n9458), .A2(n6638), .ZN(n9354) );
  AOI211_X1 U10564 ( .C1(n9456), .C2(n9409), .A(n9355), .B(n9354), .ZN(n9356)
         );
  OAI21_X1 U10565 ( .B1(n9459), .B2(n9411), .A(n9356), .ZN(P1_U3271) );
  XNOR2_X1 U10566 ( .A(n9357), .B(n9364), .ZN(n9464) );
  INV_X1 U10567 ( .A(n9375), .ZN(n9360) );
  INV_X1 U10568 ( .A(n9358), .ZN(n9359) );
  AOI21_X1 U10569 ( .B1(n9460), .B2(n9360), .A(n9359), .ZN(n9461) );
  AOI22_X1 U10570 ( .A1(n6638), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9361), .B2(
        n9393), .ZN(n9362) );
  OAI21_X1 U10571 ( .B1(n9363), .B2(n9396), .A(n9362), .ZN(n9372) );
  NAND3_X1 U10572 ( .A1(n9366), .A2(n9365), .A3(n9364), .ZN(n9367) );
  NAND2_X1 U10573 ( .A1(n9368), .A2(n9367), .ZN(n9370) );
  AOI222_X1 U10574 ( .A1(n9406), .A2(n9370), .B1(n9404), .B2(n9401), .C1(n9369), .C2(n9403), .ZN(n9463) );
  NOR2_X1 U10575 ( .A1(n9463), .A2(n6638), .ZN(n9371) );
  AOI211_X1 U10576 ( .C1(n9461), .C2(n9409), .A(n9372), .B(n9371), .ZN(n9373)
         );
  OAI21_X1 U10577 ( .B1(n9411), .B2(n9464), .A(n9373), .ZN(P1_U3272) );
  XNOR2_X1 U10578 ( .A(n9374), .B(n9381), .ZN(n9469) );
  AOI21_X1 U10579 ( .B1(n9465), .B2(n9390), .A(n9375), .ZN(n9466) );
  AOI22_X1 U10580 ( .A1(n6638), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9376), .B2(
        n9393), .ZN(n9377) );
  OAI21_X1 U10581 ( .B1(n9378), .B2(n9396), .A(n9377), .ZN(n9387) );
  NAND2_X1 U10582 ( .A1(n9380), .A2(n9379), .ZN(n9382) );
  XNOR2_X1 U10583 ( .A(n9382), .B(n9381), .ZN(n9385) );
  AOI222_X1 U10584 ( .A1(n9406), .A2(n9385), .B1(n9384), .B2(n9401), .C1(n9383), .C2(n9403), .ZN(n9468) );
  NOR2_X1 U10585 ( .A1(n9468), .A2(n6638), .ZN(n9386) );
  AOI211_X1 U10586 ( .C1(n9466), .C2(n9409), .A(n9387), .B(n9386), .ZN(n9388)
         );
  OAI21_X1 U10587 ( .B1(n9411), .B2(n9469), .A(n9388), .ZN(P1_U3273) );
  XOR2_X1 U10588 ( .A(n9389), .B(n9399), .Z(n9474) );
  INV_X1 U10589 ( .A(n9390), .ZN(n9391) );
  AOI21_X1 U10590 ( .B1(n9470), .B2(n9392), .A(n9391), .ZN(n9471) );
  AOI22_X1 U10591 ( .A1(n6638), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9394), .B2(
        n9393), .ZN(n9395) );
  OAI21_X1 U10592 ( .B1(n4599), .B2(n9396), .A(n9395), .ZN(n9408) );
  NAND2_X1 U10593 ( .A1(n9398), .A2(n9397), .ZN(n9400) );
  XNOR2_X1 U10594 ( .A(n9400), .B(n9399), .ZN(n9405) );
  AOI222_X1 U10595 ( .A1(n9406), .A2(n9405), .B1(n9404), .B2(n9403), .C1(n9402), .C2(n9401), .ZN(n9473) );
  NOR2_X1 U10596 ( .A1(n9473), .A2(n6638), .ZN(n9407) );
  AOI211_X1 U10597 ( .C1(n9471), .C2(n9409), .A(n9408), .B(n9407), .ZN(n9410)
         );
  OAI21_X1 U10598 ( .B1(n9411), .B2(n9474), .A(n9410), .ZN(P1_U3274) );
  OAI22_X1 U10599 ( .A1(n9412), .A2(n9707), .B1(n4596), .B2(n9714), .ZN(n9413)
         );
  MUX2_X1 U10600 ( .A(n9417), .B(n9488), .S(n9486), .Z(n9418) );
  INV_X1 U10601 ( .A(n9418), .ZN(P1_U3551) );
  AOI21_X1 U10602 ( .B1(n9483), .B2(n9420), .A(n9419), .ZN(n9421) );
  OAI211_X1 U10603 ( .C1(n9423), .C2(n9561), .A(n9422), .B(n9421), .ZN(n9491)
         );
  MUX2_X1 U10604 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9491), .S(n9486), .Z(
        P1_U3550) );
  AOI22_X1 U10605 ( .A1(n9425), .A2(n9559), .B1(n9483), .B2(n9424), .ZN(n9426)
         );
  OAI211_X1 U10606 ( .C1(n9428), .C2(n9561), .A(n9427), .B(n9426), .ZN(n9492)
         );
  MUX2_X1 U10607 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9492), .S(n9486), .Z(
        P1_U3549) );
  AOI22_X1 U10608 ( .A1(n9430), .A2(n9559), .B1(n9483), .B2(n9429), .ZN(n9431)
         );
  OAI211_X1 U10609 ( .C1(n9433), .C2(n9561), .A(n9432), .B(n9431), .ZN(n9493)
         );
  MUX2_X1 U10610 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9493), .S(n9486), .Z(
        P1_U3548) );
  AOI211_X1 U10611 ( .C1(n9483), .C2(n9436), .A(n9435), .B(n9434), .ZN(n9437)
         );
  OAI21_X1 U10612 ( .B1(n9438), .B2(n9561), .A(n9437), .ZN(n9494) );
  MUX2_X1 U10613 ( .A(n9494), .B(P1_REG1_REG_24__SCAN_IN), .S(n9725), .Z(
        P1_U3547) );
  AOI211_X1 U10614 ( .C1(n9483), .C2(n9441), .A(n9440), .B(n9439), .ZN(n9442)
         );
  OAI21_X1 U10615 ( .B1(n9443), .B2(n9561), .A(n9442), .ZN(n9495) );
  MUX2_X1 U10616 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9495), .S(n9486), .Z(
        P1_U3546) );
  OAI22_X1 U10617 ( .A1(n9445), .A2(n9707), .B1(n9444), .B2(n9714), .ZN(n9446)
         );
  AOI211_X1 U10618 ( .C1(n9448), .C2(n9578), .A(n9447), .B(n9446), .ZN(n9449)
         );
  INV_X1 U10619 ( .A(n9449), .ZN(n9496) );
  MUX2_X1 U10620 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9496), .S(n9486), .Z(
        P1_U3545) );
  AOI211_X1 U10621 ( .C1(n9483), .C2(n9452), .A(n9451), .B(n9450), .ZN(n9453)
         );
  OAI21_X1 U10622 ( .B1(n9454), .B2(n9561), .A(n9453), .ZN(n9497) );
  MUX2_X1 U10623 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9497), .S(n9486), .Z(
        P1_U3544) );
  AOI22_X1 U10624 ( .A1(n9456), .A2(n9559), .B1(n9483), .B2(n9455), .ZN(n9457)
         );
  OAI211_X1 U10625 ( .C1(n9459), .C2(n9561), .A(n9458), .B(n9457), .ZN(n9498)
         );
  MUX2_X1 U10626 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9498), .S(n9486), .Z(
        P1_U3543) );
  AOI22_X1 U10627 ( .A1(n9461), .A2(n9559), .B1(n9483), .B2(n9460), .ZN(n9462)
         );
  OAI211_X1 U10628 ( .C1(n9464), .C2(n9561), .A(n9463), .B(n9462), .ZN(n9499)
         );
  MUX2_X1 U10629 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9499), .S(n9486), .Z(
        P1_U3542) );
  AOI22_X1 U10630 ( .A1(n9466), .A2(n9559), .B1(n9483), .B2(n9465), .ZN(n9467)
         );
  OAI211_X1 U10631 ( .C1(n9469), .C2(n9561), .A(n9468), .B(n9467), .ZN(n9500)
         );
  MUX2_X1 U10632 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9500), .S(n9486), .Z(
        P1_U3541) );
  AOI22_X1 U10633 ( .A1(n9471), .A2(n9559), .B1(n9483), .B2(n9470), .ZN(n9472)
         );
  OAI211_X1 U10634 ( .C1(n9474), .C2(n9561), .A(n9473), .B(n9472), .ZN(n9501)
         );
  MUX2_X1 U10635 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9501), .S(n9486), .Z(
        P1_U3540) );
  AOI21_X1 U10636 ( .B1(n9483), .B2(n9476), .A(n9475), .ZN(n9477) );
  OAI211_X1 U10637 ( .C1(n9479), .C2(n9561), .A(n9478), .B(n9477), .ZN(n9502)
         );
  MUX2_X1 U10638 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9502), .S(n9486), .Z(
        P1_U3537) );
  AOI211_X1 U10639 ( .C1(n9483), .C2(n9482), .A(n9481), .B(n9480), .ZN(n9484)
         );
  OAI21_X1 U10640 ( .B1(n9561), .B2(n9485), .A(n9484), .ZN(n9503) );
  MUX2_X1 U10641 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n9503), .S(n9486), .Z(
        P1_U3535) );
  MUX2_X1 U10642 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9487), .S(n9722), .Z(
        P1_U3520) );
  INV_X1 U10643 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n9489) );
  MUX2_X1 U10644 ( .A(n9489), .B(n9488), .S(n9722), .Z(n9490) );
  INV_X1 U10645 ( .A(n9490), .ZN(P1_U3519) );
  MUX2_X1 U10646 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9491), .S(n9722), .Z(
        P1_U3518) );
  MUX2_X1 U10647 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9492), .S(n9722), .Z(
        P1_U3517) );
  MUX2_X1 U10648 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9493), .S(n9722), .Z(
        P1_U3516) );
  MUX2_X1 U10649 ( .A(n9494), .B(P1_REG0_REG_24__SCAN_IN), .S(n9721), .Z(
        P1_U3515) );
  MUX2_X1 U10650 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9495), .S(n9722), .Z(
        P1_U3514) );
  MUX2_X1 U10651 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9496), .S(n9722), .Z(
        P1_U3513) );
  MUX2_X1 U10652 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9497), .S(n9722), .Z(
        P1_U3512) );
  MUX2_X1 U10653 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9498), .S(n9722), .Z(
        P1_U3511) );
  MUX2_X1 U10654 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9499), .S(n9722), .Z(
        P1_U3510) );
  MUX2_X1 U10655 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9500), .S(n9722), .Z(
        P1_U3508) );
  MUX2_X1 U10656 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9501), .S(n9722), .Z(
        P1_U3505) );
  MUX2_X1 U10657 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n9502), .S(n9722), .Z(
        P1_U3496) );
  MUX2_X1 U10658 ( .A(P1_REG0_REG_12__SCAN_IN), .B(n9503), .S(n9722), .Z(
        P1_U3490) );
  NOR4_X1 U10659 ( .A1(n5701), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3084), .A4(
        n9504), .ZN(n9505) );
  AOI21_X1 U10660 ( .B1(n9506), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9505), .ZN(
        n9507) );
  OAI21_X1 U10661 ( .B1(n9509), .B2(n9508), .A(n9507), .ZN(P1_U3322) );
  OAI222_X1 U10662 ( .A1(P1_U3084), .A2(n6249), .B1(n9508), .B2(n9512), .C1(
        n9511), .C2(n9510), .ZN(P1_U3325) );
  MUX2_X1 U10663 ( .A(n9513), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  AOI22_X1 U10664 ( .A1(n9734), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3152), .ZN(n9526) );
  OR2_X1 U10665 ( .A1(n9730), .A2(n4947), .ZN(n9520) );
  INV_X1 U10666 ( .A(n9514), .ZN(n9518) );
  NAND2_X1 U10667 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n9515) );
  NAND2_X1 U10668 ( .A1(n9516), .A2(n9515), .ZN(n9517) );
  NAND3_X1 U10669 ( .A1(n9729), .A2(n9518), .A3(n9517), .ZN(n9519) );
  AND2_X1 U10670 ( .A1(n9520), .A2(n9519), .ZN(n9525) );
  NOR2_X1 U10671 ( .A1(n9737), .A2(n9955), .ZN(n9523) );
  OAI211_X1 U10672 ( .C1(n9523), .C2(n9522), .A(n9728), .B(n9521), .ZN(n9524)
         );
  NAND3_X1 U10673 ( .A1(n9526), .A2(n9525), .A3(n9524), .ZN(P2_U3246) );
  AOI22_X1 U10674 ( .A1(n9734), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n9540) );
  AOI211_X1 U10675 ( .C1(n9531), .C2(n9530), .A(n9529), .B(n9528), .ZN(n9532)
         );
  AOI21_X1 U10676 ( .B1(n9534), .B2(n9533), .A(n9532), .ZN(n9539) );
  OAI211_X1 U10677 ( .C1(n9537), .C2(n9536), .A(n9728), .B(n9535), .ZN(n9538)
         );
  NAND3_X1 U10678 ( .A1(n9540), .A2(n9539), .A3(n9538), .ZN(P2_U3247) );
  OAI21_X1 U10679 ( .B1(n9542), .B2(n9714), .A(n9541), .ZN(n9543) );
  AOI21_X1 U10680 ( .B1(n9544), .B2(n9717), .A(n9543), .ZN(n9545) );
  AND2_X1 U10681 ( .A1(n9546), .A2(n9545), .ZN(n9548) );
  INV_X1 U10682 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n9547) );
  AOI22_X1 U10683 ( .A1(n9722), .A2(n9548), .B1(n9547), .B2(n9721), .ZN(
        P1_U3484) );
  AOI22_X1 U10684 ( .A1(n9486), .A2(n9548), .B1(n6598), .B2(n9725), .ZN(
        P1_U3533) );
  OAI21_X1 U10685 ( .B1(n9549), .B2(n9714), .A(n9555), .ZN(n9550) );
  AOI21_X1 U10686 ( .B1(n9551), .B2(n9559), .A(n9550), .ZN(n9554) );
  INV_X1 U10687 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9552) );
  AOI22_X1 U10688 ( .A1(n9486), .A2(n9554), .B1(n9552), .B2(n9725), .ZN(
        P1_U3554) );
  INV_X1 U10689 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n9553) );
  AOI22_X1 U10690 ( .A1(n9722), .A2(n9554), .B1(n9553), .B2(n9721), .ZN(
        P1_U3522) );
  OAI21_X1 U10691 ( .B1(n9556), .B2(n9714), .A(n9555), .ZN(n9557) );
  AOI21_X1 U10692 ( .B1(n9559), .B2(n9558), .A(n9557), .ZN(n9588) );
  INV_X1 U10693 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9560) );
  AOI22_X1 U10694 ( .A1(n9486), .A2(n9588), .B1(n9560), .B2(n9725), .ZN(
        P1_U3553) );
  NOR2_X1 U10695 ( .A1(n9562), .A2(n9561), .ZN(n9566) );
  OAI211_X1 U10696 ( .C1(n4600), .C2(n9714), .A(n9564), .B(n9563), .ZN(n9565)
         );
  AOI21_X1 U10697 ( .B1(n9566), .B2(n7941), .A(n9565), .ZN(n9590) );
  AOI22_X1 U10698 ( .A1(n9486), .A2(n9590), .B1(n9567), .B2(n9725), .ZN(
        P1_U3539) );
  OAI211_X1 U10699 ( .C1(n9570), .C2(n9714), .A(n9569), .B(n9568), .ZN(n9571)
         );
  AOI21_X1 U10700 ( .B1(n9572), .B2(n9578), .A(n9571), .ZN(n9592) );
  AOI22_X1 U10701 ( .A1(n9486), .A2(n9592), .B1(n9573), .B2(n9725), .ZN(
        P1_U3538) );
  OAI211_X1 U10702 ( .C1(n9576), .C2(n9714), .A(n9575), .B(n9574), .ZN(n9577)
         );
  AOI21_X1 U10703 ( .B1(n9579), .B2(n9578), .A(n9577), .ZN(n9594) );
  AOI22_X1 U10704 ( .A1(n9486), .A2(n9594), .B1(n9580), .B2(n9725), .ZN(
        P1_U3536) );
  OAI21_X1 U10705 ( .B1(n9582), .B2(n9714), .A(n9581), .ZN(n9583) );
  AOI21_X1 U10706 ( .B1(n9584), .B2(n9717), .A(n9583), .ZN(n9585) );
  AND2_X1 U10707 ( .A1(n9586), .A2(n9585), .ZN(n9596) );
  AOI22_X1 U10708 ( .A1(n9486), .A2(n9596), .B1(n6601), .B2(n9725), .ZN(
        P1_U3534) );
  INV_X1 U10709 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9587) );
  AOI22_X1 U10710 ( .A1(n9722), .A2(n9588), .B1(n9587), .B2(n9721), .ZN(
        P1_U3521) );
  INV_X1 U10711 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n9589) );
  AOI22_X1 U10712 ( .A1(n9722), .A2(n9590), .B1(n9589), .B2(n9721), .ZN(
        P1_U3502) );
  INV_X1 U10713 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n9591) );
  AOI22_X1 U10714 ( .A1(n9722), .A2(n9592), .B1(n9591), .B2(n9721), .ZN(
        P1_U3499) );
  INV_X1 U10715 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n9593) );
  AOI22_X1 U10716 ( .A1(n9722), .A2(n9594), .B1(n9593), .B2(n9721), .ZN(
        P1_U3493) );
  INV_X1 U10717 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n9595) );
  AOI22_X1 U10718 ( .A1(n9722), .A2(n9596), .B1(n9595), .B2(n9721), .ZN(
        P1_U3487) );
  XNOR2_X1 U10719 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  NOR2_X1 U10720 ( .A1(n9597), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n9600) );
  NOR2_X1 U10721 ( .A1(n9598), .A2(n6783), .ZN(n9599) );
  MUX2_X1 U10722 ( .A(n9600), .B(n9599), .S(P1_IR_REG_0__SCAN_IN), .Z(n9601)
         );
  OR2_X1 U10723 ( .A1(n9602), .A2(n9601), .ZN(n9605) );
  AOI22_X1 U10724 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(n9648), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3084), .ZN(n9603) );
  OAI21_X1 U10725 ( .B1(n9605), .B2(n9604), .A(n9603), .ZN(P1_U3241) );
  INV_X1 U10726 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n9617) );
  XOR2_X1 U10727 ( .A(n9607), .B(n9606), .Z(n9609) );
  OAI22_X1 U10728 ( .A1(n9634), .A2(n9609), .B1(n9646), .B2(n9608), .ZN(n9611)
         );
  AOI211_X1 U10729 ( .C1(n9648), .C2(P1_ADDR_REG_2__SCAN_IN), .A(n9611), .B(
        n9610), .ZN(n9616) );
  OAI211_X1 U10730 ( .C1(n9614), .C2(n9613), .A(n9673), .B(n9612), .ZN(n9615)
         );
  OAI211_X1 U10731 ( .C1(P1_STATE_REG_SCAN_IN), .C2(n9617), .A(n9616), .B(
        n9615), .ZN(P1_U3243) );
  AOI21_X1 U10732 ( .B1(n9620), .B2(n9619), .A(n9618), .ZN(n9621) );
  NOR2_X1 U10733 ( .A1(n9621), .A2(n9634), .ZN(n9622) );
  AOI211_X1 U10734 ( .C1(n9664), .C2(n9624), .A(n9623), .B(n9622), .ZN(n9629)
         );
  OAI211_X1 U10735 ( .C1(n9627), .C2(n9626), .A(n9673), .B(n9625), .ZN(n9628)
         );
  OAI211_X1 U10736 ( .C1(n10081), .C2(n9678), .A(n9629), .B(n9628), .ZN(
        P1_U3250) );
  AOI22_X1 U10737 ( .A1(n9648), .A2(P1_ADDR_REG_10__SCAN_IN), .B1(n9664), .B2(
        n9630), .ZN(n9642) );
  AOI21_X1 U10738 ( .B1(n9633), .B2(n9632), .A(n9631), .ZN(n9635) );
  OR2_X1 U10739 ( .A1(n9635), .A2(n9634), .ZN(n9640) );
  OAI211_X1 U10740 ( .C1(n9638), .C2(n9637), .A(n9673), .B(n9636), .ZN(n9639)
         );
  NAND4_X1 U10741 ( .A1(n9642), .A2(n9641), .A3(n9640), .A4(n9639), .ZN(
        P1_U3251) );
  NAND3_X1 U10742 ( .A1(n9657), .A2(P1_REG2_REG_11__SCAN_IN), .A3(n9643), .ZN(
        n9647) );
  INV_X1 U10743 ( .A(n9644), .ZN(n9653) );
  NAND3_X1 U10744 ( .A1(n9672), .A2(P1_REG1_REG_11__SCAN_IN), .A3(n9653), .ZN(
        n9645) );
  NAND3_X1 U10745 ( .A1(n9647), .A2(n9646), .A3(n9645), .ZN(n9649) );
  AOI22_X1 U10746 ( .A1(n9650), .A2(n9649), .B1(n9648), .B2(
        P1_ADDR_REG_11__SCAN_IN), .ZN(n9661) );
  OAI211_X1 U10747 ( .C1(n9653), .C2(n9652), .A(n9672), .B(n9651), .ZN(n9659)
         );
  NAND2_X1 U10748 ( .A1(n9654), .A2(n9890), .ZN(n9656) );
  OAI211_X1 U10749 ( .C1(n9657), .C2(n9656), .A(n9655), .B(n9673), .ZN(n9658)
         );
  NAND4_X1 U10750 ( .A1(n9661), .A2(n9660), .A3(n9659), .A4(n9658), .ZN(
        P1_U3252) );
  INV_X1 U10751 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n9677) );
  AOI21_X1 U10752 ( .B1(n9664), .B2(n9663), .A(n9662), .ZN(n9676) );
  OAI21_X1 U10753 ( .B1(n9667), .B2(n9666), .A(n9665), .ZN(n9674) );
  OAI21_X1 U10754 ( .B1(n9670), .B2(n9669), .A(n9668), .ZN(n9671) );
  AOI22_X1 U10755 ( .A1(n9674), .A2(n9673), .B1(n9672), .B2(n9671), .ZN(n9675)
         );
  OAI211_X1 U10756 ( .C1(n9678), .C2(n9677), .A(n9676), .B(n9675), .ZN(
        P1_U3255) );
  INV_X1 U10757 ( .A(n9679), .ZN(n9687) );
  AOI22_X1 U10758 ( .A1(n9683), .A2(n9682), .B1(n9681), .B2(n9680), .ZN(n9684)
         );
  OAI211_X1 U10759 ( .C1(n9687), .C2(n9686), .A(n9685), .B(n9684), .ZN(n9689)
         );
  AOI22_X1 U10760 ( .A1(n6638), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n9689), .B2(
        n9688), .ZN(n9690) );
  OAI21_X1 U10761 ( .B1(n9692), .B2(n9691), .A(n9690), .ZN(P1_U3286) );
  AND2_X1 U10762 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9694), .ZN(P1_U3292) );
  AND2_X1 U10763 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9694), .ZN(P1_U3293) );
  AND2_X1 U10764 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9694), .ZN(P1_U3294) );
  INV_X1 U10765 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n9894) );
  NOR2_X1 U10766 ( .A1(n9693), .A2(n9894), .ZN(P1_U3295) );
  AND2_X1 U10767 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9694), .ZN(P1_U3296) );
  AND2_X1 U10768 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9694), .ZN(P1_U3297) );
  AND2_X1 U10769 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9694), .ZN(P1_U3298) );
  AND2_X1 U10770 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9694), .ZN(P1_U3299) );
  AND2_X1 U10771 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9694), .ZN(P1_U3300) );
  AND2_X1 U10772 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9694), .ZN(P1_U3301) );
  AND2_X1 U10773 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9694), .ZN(P1_U3302) );
  AND2_X1 U10774 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9694), .ZN(P1_U3303) );
  AND2_X1 U10775 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9694), .ZN(P1_U3304) );
  INV_X1 U10776 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n10019) );
  NOR2_X1 U10777 ( .A1(n9693), .A2(n10019), .ZN(P1_U3305) );
  AND2_X1 U10778 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9694), .ZN(P1_U3306) );
  AND2_X1 U10779 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9694), .ZN(P1_U3307) );
  AND2_X1 U10780 ( .A1(n9694), .A2(P1_D_REG_15__SCAN_IN), .ZN(P1_U3308) );
  AND2_X1 U10781 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9694), .ZN(P1_U3309) );
  AND2_X1 U10782 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9694), .ZN(P1_U3310) );
  AND2_X1 U10783 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9694), .ZN(P1_U3311) );
  INV_X1 U10784 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n9965) );
  NOR2_X1 U10785 ( .A1(n9693), .A2(n9965), .ZN(P1_U3312) );
  AND2_X1 U10786 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9694), .ZN(P1_U3313) );
  INV_X1 U10787 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n10018) );
  NOR2_X1 U10788 ( .A1(n9693), .A2(n10018), .ZN(P1_U3314) );
  AND2_X1 U10789 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9694), .ZN(P1_U3315) );
  AND2_X1 U10790 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9694), .ZN(P1_U3316) );
  AND2_X1 U10791 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9694), .ZN(P1_U3317) );
  AND2_X1 U10792 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9694), .ZN(P1_U3318) );
  AND2_X1 U10793 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9694), .ZN(P1_U3319) );
  AND2_X1 U10794 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9694), .ZN(P1_U3320) );
  AND2_X1 U10795 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9694), .ZN(P1_U3321) );
  INV_X1 U10796 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n9696) );
  OAI21_X1 U10797 ( .B1(n9697), .B2(n9696), .A(n9695), .ZN(P1_U3440) );
  INV_X1 U10798 ( .A(n9698), .ZN(n9700) );
  OAI211_X1 U10799 ( .C1(n6618), .C2(n9714), .A(n9700), .B(n9699), .ZN(n9703)
         );
  INV_X1 U10800 ( .A(n9701), .ZN(n9702) );
  AOI211_X1 U10801 ( .C1(n9717), .C2(n9704), .A(n9703), .B(n9702), .ZN(n9723)
         );
  INV_X1 U10802 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9705) );
  AOI22_X1 U10803 ( .A1(n9722), .A2(n9723), .B1(n9705), .B2(n9721), .ZN(
        P1_U3457) );
  OAI22_X1 U10804 ( .A1(n9708), .A2(n9707), .B1(n9706), .B2(n9714), .ZN(n9710)
         );
  AOI211_X1 U10805 ( .C1(n9717), .C2(n9711), .A(n9710), .B(n9709), .ZN(n9724)
         );
  INV_X1 U10806 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n9712) );
  AOI22_X1 U10807 ( .A1(n9722), .A2(n9724), .B1(n9712), .B2(n9721), .ZN(
        P1_U3463) );
  OAI21_X1 U10808 ( .B1(n9715), .B2(n9714), .A(n9713), .ZN(n9716) );
  AOI21_X1 U10809 ( .B1(n9718), .B2(n9717), .A(n9716), .ZN(n9719) );
  AND2_X1 U10810 ( .A1(n9720), .A2(n9719), .ZN(n9727) );
  INV_X1 U10811 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9940) );
  AOI22_X1 U10812 ( .A1(n9722), .A2(n9727), .B1(n9940), .B2(n9721), .ZN(
        P1_U3481) );
  AOI22_X1 U10813 ( .A1(n9486), .A2(n9723), .B1(n6581), .B2(n9725), .ZN(
        P1_U3524) );
  AOI22_X1 U10814 ( .A1(n9486), .A2(n9724), .B1(n6586), .B2(n9725), .ZN(
        P1_U3526) );
  AOI22_X1 U10815 ( .A1(n9486), .A2(n9727), .B1(n9726), .B2(n9725), .ZN(
        P1_U3532) );
  AOI22_X1 U10816 ( .A1(n9728), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n9729), .ZN(n9738) );
  NAND2_X1 U10817 ( .A1(n9729), .A2(n9834), .ZN(n9731) );
  OAI211_X1 U10818 ( .C1(n9732), .C2(P2_REG2_REG_0__SCAN_IN), .A(n9731), .B(
        n9730), .ZN(n9733) );
  INV_X1 U10819 ( .A(n9733), .ZN(n9736) );
  AOI22_X1 U10820 ( .A1(n9734), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n9735) );
  OAI221_X1 U10821 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n9738), .C1(n9737), .C2(
        n9736), .A(n9735), .ZN(P2_U3245) );
  NAND3_X1 U10822 ( .A1(n9740), .A2(n9753), .A3(n9739), .ZN(n9741) );
  NAND2_X1 U10823 ( .A1(n9742), .A2(n9741), .ZN(n9746) );
  AOI222_X1 U10824 ( .A1(n8813), .A2(n9746), .B1(n9745), .B2(n9744), .C1(n7029), .C2(n9743), .ZN(n9782) );
  AOI22_X1 U10825 ( .A1(n9747), .A2(n5001), .B1(P2_REG2_REG_3__SCAN_IN), .B2(
        n8804), .ZN(n9757) );
  AND2_X1 U10826 ( .A1(n9748), .A2(n9803), .ZN(n9751) );
  OAI21_X1 U10827 ( .B1(n9748), .B2(n9825), .A(n9824), .ZN(n9750) );
  MUX2_X1 U10828 ( .A(n9751), .B(n9750), .S(n9749), .Z(n9784) );
  XNOR2_X1 U10829 ( .A(n9752), .B(n9753), .ZN(n9785) );
  AOI22_X1 U10830 ( .A1(n9755), .A2(n9784), .B1(n9754), .B2(n9785), .ZN(n9756)
         );
  OAI211_X1 U10831 ( .C1(n8804), .C2(n9782), .A(n9757), .B(n9756), .ZN(
        P2_U3293) );
  NOR2_X1 U10832 ( .A1(n9759), .A2(n9758), .ZN(n9761) );
  AND2_X1 U10833 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n9765), .ZN(P2_U3297) );
  AND2_X1 U10834 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n9765), .ZN(P2_U3298) );
  NOR2_X1 U10835 ( .A1(n9761), .A2(n10047), .ZN(P2_U3299) );
  AND2_X1 U10836 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n9765), .ZN(P2_U3300) );
  AND2_X1 U10837 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n9765), .ZN(P2_U3301) );
  AND2_X1 U10838 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n9765), .ZN(P2_U3302) );
  AND2_X1 U10839 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n9765), .ZN(P2_U3303) );
  AND2_X1 U10840 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n9765), .ZN(P2_U3304) );
  AND2_X1 U10841 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n9765), .ZN(P2_U3305) );
  AND2_X1 U10842 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n9765), .ZN(P2_U3306) );
  AND2_X1 U10843 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n9765), .ZN(P2_U3307) );
  AND2_X1 U10844 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n9765), .ZN(P2_U3308) );
  AND2_X1 U10845 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n9765), .ZN(P2_U3309) );
  AND2_X1 U10846 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n9765), .ZN(P2_U3310) );
  AND2_X1 U10847 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n9765), .ZN(P2_U3311) );
  AND2_X1 U10848 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n9765), .ZN(P2_U3312) );
  NOR2_X1 U10849 ( .A1(n9761), .A2(n10056), .ZN(P2_U3313) );
  NOR2_X1 U10850 ( .A1(n9761), .A2(n9760), .ZN(P2_U3314) );
  AND2_X1 U10851 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n9765), .ZN(P2_U3315) );
  AND2_X1 U10852 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n9765), .ZN(P2_U3316) );
  NOR2_X1 U10853 ( .A1(n9761), .A2(n10022), .ZN(P2_U3317) );
  AND2_X1 U10854 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n9765), .ZN(P2_U3318) );
  AND2_X1 U10855 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n9765), .ZN(P2_U3319) );
  AND2_X1 U10856 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n9765), .ZN(P2_U3320) );
  AND2_X1 U10857 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n9765), .ZN(P2_U3321) );
  INV_X1 U10858 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n10043) );
  NOR2_X1 U10859 ( .A1(n9761), .A2(n10043), .ZN(P2_U3322) );
  AND2_X1 U10860 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n9765), .ZN(P2_U3323) );
  AND2_X1 U10861 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n9765), .ZN(P2_U3324) );
  INV_X1 U10862 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n10044) );
  NOR2_X1 U10863 ( .A1(n9761), .A2(n10044), .ZN(P2_U3325) );
  AND2_X1 U10864 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n9765), .ZN(P2_U3326) );
  NOR2_X1 U10865 ( .A1(n9762), .A2(P2_U3152), .ZN(n9767) );
  AOI22_X1 U10866 ( .A1(n9764), .A2(n9767), .B1(n9763), .B2(n9765), .ZN(
        P2_U3437) );
  AOI22_X1 U10867 ( .A1(n9768), .A2(n9767), .B1(n9766), .B2(n9765), .ZN(
        P2_U3438) );
  NAND2_X1 U10868 ( .A1(n9769), .A2(n9829), .ZN(n9772) );
  NAND2_X1 U10869 ( .A1(n9770), .A2(n4702), .ZN(n9771) );
  NAND2_X1 U10870 ( .A1(n9772), .A2(n9771), .ZN(n9773) );
  NOR2_X1 U10871 ( .A1(n9774), .A2(n9773), .ZN(n9835) );
  INV_X1 U10872 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n9775) );
  AOI22_X1 U10873 ( .A1(n9833), .A2(n9835), .B1(n9775), .B2(n9831), .ZN(
        P2_U3451) );
  OAI22_X1 U10874 ( .A1(n9777), .A2(n9825), .B1(n9776), .B2(n9824), .ZN(n9779)
         );
  AOI211_X1 U10875 ( .C1(n9829), .C2(n9780), .A(n9779), .B(n9778), .ZN(n9837)
         );
  INV_X1 U10876 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n9781) );
  AOI22_X1 U10877 ( .A1(n9833), .A2(n9837), .B1(n9781), .B2(n9831), .ZN(
        P2_U3457) );
  INV_X1 U10878 ( .A(n9782), .ZN(n9783) );
  AOI211_X1 U10879 ( .C1(n9829), .C2(n9785), .A(n9784), .B(n9783), .ZN(n9838)
         );
  INV_X1 U10880 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n9786) );
  AOI22_X1 U10881 ( .A1(n9833), .A2(n9838), .B1(n9786), .B2(n9831), .ZN(
        P2_U3460) );
  INV_X1 U10882 ( .A(n9787), .ZN(n9789) );
  OAI22_X1 U10883 ( .A1(n9789), .A2(n9825), .B1(n9788), .B2(n9824), .ZN(n9791)
         );
  AOI211_X1 U10884 ( .C1(n9829), .C2(n9792), .A(n9791), .B(n9790), .ZN(n9840)
         );
  INV_X1 U10885 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n9930) );
  AOI22_X1 U10886 ( .A1(n9833), .A2(n9840), .B1(n9930), .B2(n9831), .ZN(
        P2_U3463) );
  AOI21_X1 U10887 ( .B1(n9802), .B2(n9794), .A(n9793), .ZN(n9795) );
  OAI211_X1 U10888 ( .C1(n9798), .C2(n9797), .A(n9796), .B(n9795), .ZN(n9799)
         );
  INV_X1 U10889 ( .A(n9799), .ZN(n9842) );
  INV_X1 U10890 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n9800) );
  AOI22_X1 U10891 ( .A1(n9833), .A2(n9842), .B1(n9800), .B2(n9831), .ZN(
        P2_U3466) );
  AOI22_X1 U10892 ( .A1(n9804), .A2(n9803), .B1(n9802), .B2(n9801), .ZN(n9805)
         );
  NAND2_X1 U10893 ( .A1(n9806), .A2(n9805), .ZN(n9807) );
  AOI21_X1 U10894 ( .B1(n9829), .B2(n9808), .A(n9807), .ZN(n9843) );
  INV_X1 U10895 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n9946) );
  AOI22_X1 U10896 ( .A1(n9833), .A2(n9843), .B1(n9946), .B2(n9831), .ZN(
        P2_U3469) );
  NOR2_X1 U10897 ( .A1(n9810), .A2(n9809), .ZN(n9813) );
  OAI22_X1 U10898 ( .A1(n9811), .A2(n9825), .B1(n4517), .B2(n9824), .ZN(n9812)
         );
  NOR3_X1 U10899 ( .A1(n9814), .A2(n9813), .A3(n9812), .ZN(n9844) );
  INV_X1 U10900 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n9815) );
  AOI22_X1 U10901 ( .A1(n9833), .A2(n9844), .B1(n9815), .B2(n9831), .ZN(
        P2_U3475) );
  INV_X1 U10902 ( .A(n9816), .ZN(n9821) );
  OAI22_X1 U10903 ( .A1(n9818), .A2(n9825), .B1(n9817), .B2(n9824), .ZN(n9820)
         );
  AOI211_X1 U10904 ( .C1(n9822), .C2(n9821), .A(n9820), .B(n9819), .ZN(n9845)
         );
  INV_X1 U10905 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n9823) );
  AOI22_X1 U10906 ( .A1(n9833), .A2(n9845), .B1(n9823), .B2(n9831), .ZN(
        P2_U3481) );
  OAI22_X1 U10907 ( .A1(n9826), .A2(n9825), .B1(n4534), .B2(n9824), .ZN(n9828)
         );
  AOI211_X1 U10908 ( .C1(n9830), .C2(n9829), .A(n9828), .B(n9827), .ZN(n9847)
         );
  INV_X1 U10909 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n9832) );
  AOI22_X1 U10910 ( .A1(n9833), .A2(n9847), .B1(n9832), .B2(n9831), .ZN(
        P2_U3487) );
  AOI22_X1 U10911 ( .A1(n9848), .A2(n9835), .B1(n9834), .B2(n9846), .ZN(
        P2_U3520) );
  INV_X1 U10912 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n9836) );
  AOI22_X1 U10913 ( .A1(n9848), .A2(n9837), .B1(n9836), .B2(n9846), .ZN(
        P2_U3522) );
  INV_X1 U10914 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n9964) );
  AOI22_X1 U10915 ( .A1(n9848), .A2(n9838), .B1(n9964), .B2(n9846), .ZN(
        P2_U3523) );
  INV_X1 U10916 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n9839) );
  AOI22_X1 U10917 ( .A1(n9848), .A2(n9840), .B1(n9839), .B2(n9846), .ZN(
        P2_U3524) );
  INV_X1 U10918 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n9841) );
  AOI22_X1 U10919 ( .A1(n9848), .A2(n9842), .B1(n9841), .B2(n9846), .ZN(
        P2_U3525) );
  INV_X1 U10920 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n9971) );
  AOI22_X1 U10921 ( .A1(n9848), .A2(n9843), .B1(n9971), .B2(n9846), .ZN(
        P2_U3526) );
  AOI22_X1 U10922 ( .A1(n9848), .A2(n9844), .B1(n6872), .B2(n9846), .ZN(
        P2_U3528) );
  AOI22_X1 U10923 ( .A1(n9848), .A2(n9845), .B1(n6874), .B2(n9846), .ZN(
        P2_U3530) );
  AOI22_X1 U10924 ( .A1(n9848), .A2(n9847), .B1(n7163), .B2(n9846), .ZN(
        P2_U3532) );
  INV_X1 U10925 ( .A(n9849), .ZN(n9850) );
  NAND2_X1 U10926 ( .A1(n9851), .A2(n9850), .ZN(n9852) );
  XOR2_X1 U10927 ( .A(n10021), .B(n9852), .Z(ADD_1071_U5) );
  XOR2_X1 U10928 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  OAI21_X1 U10929 ( .B1(n9855), .B2(n9854), .A(n9853), .ZN(ADD_1071_U56) );
  OAI21_X1 U10930 ( .B1(n9858), .B2(n9857), .A(n9856), .ZN(ADD_1071_U57) );
  OAI21_X1 U10931 ( .B1(n9861), .B2(n9860), .A(n9859), .ZN(ADD_1071_U58) );
  OAI21_X1 U10932 ( .B1(n9864), .B2(n9863), .A(n9862), .ZN(ADD_1071_U59) );
  OAI21_X1 U10933 ( .B1(n9867), .B2(n9866), .A(n9865), .ZN(ADD_1071_U60) );
  OAI21_X1 U10934 ( .B1(n9870), .B2(n9869), .A(n9868), .ZN(ADD_1071_U61) );
  AOI21_X1 U10935 ( .B1(n9873), .B2(n9872), .A(n9871), .ZN(ADD_1071_U62) );
  AOI21_X1 U10936 ( .B1(n9876), .B2(n9875), .A(n9874), .ZN(ADD_1071_U63) );
  AOI22_X1 U10937 ( .A1(n9947), .A2(keyinput1), .B1(keyinput59), .B2(n9878), 
        .ZN(n9877) );
  OAI221_X1 U10938 ( .B1(n9947), .B2(keyinput1), .C1(n9878), .C2(keyinput59), 
        .A(n9877), .ZN(n9887) );
  AOI22_X1 U10939 ( .A1(n10021), .A2(keyinput42), .B1(n9943), .B2(keyinput33), 
        .ZN(n9879) );
  OAI221_X1 U10940 ( .B1(n10021), .B2(keyinput42), .C1(n9943), .C2(keyinput33), 
        .A(n9879), .ZN(n9886) );
  AOI22_X1 U10941 ( .A1(n9946), .A2(keyinput34), .B1(n9881), .B2(keyinput16), 
        .ZN(n9880) );
  OAI221_X1 U10942 ( .B1(n9946), .B2(keyinput34), .C1(n9881), .C2(keyinput16), 
        .A(n9880), .ZN(n9885) );
  XNOR2_X1 U10943 ( .A(P2_IR_REG_19__SCAN_IN), .B(keyinput24), .ZN(n9883) );
  XNOR2_X1 U10944 ( .A(P1_IR_REG_22__SCAN_IN), .B(keyinput18), .ZN(n9882) );
  NAND2_X1 U10945 ( .A1(n9883), .A2(n9882), .ZN(n9884) );
  OR4_X1 U10946 ( .A1(n9887), .A2(n9886), .A3(n9885), .A4(n9884), .ZN(n10074)
         );
  INV_X1 U10947 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n9889) );
  OAI22_X1 U10948 ( .A1(n9890), .A2(keyinput53), .B1(n9889), .B2(keyinput45), 
        .ZN(n9888) );
  AOI221_X1 U10949 ( .B1(n9890), .B2(keyinput53), .C1(keyinput45), .C2(n9889), 
        .A(n9888), .ZN(n9901) );
  INV_X1 U10950 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n9985) );
  OAI22_X1 U10951 ( .A1(n5710), .A2(keyinput28), .B1(n9985), .B2(keyinput2), 
        .ZN(n9891) );
  AOI221_X1 U10952 ( .B1(n5710), .B2(keyinput28), .C1(keyinput2), .C2(n9985), 
        .A(n9891), .ZN(n9900) );
  OAI22_X1 U10953 ( .A1(n9894), .A2(keyinput7), .B1(n9893), .B2(keyinput50), 
        .ZN(n9892) );
  AOI221_X1 U10954 ( .B1(n9894), .B2(keyinput7), .C1(keyinput50), .C2(n9893), 
        .A(n9892), .ZN(n9899) );
  XNOR2_X1 U10955 ( .A(n9895), .B(keyinput26), .ZN(n9897) );
  XNOR2_X1 U10956 ( .A(keyinput13), .B(n9964), .ZN(n9896) );
  NOR2_X1 U10957 ( .A1(n9897), .A2(n9896), .ZN(n9898) );
  NAND4_X1 U10958 ( .A1(n9901), .A2(n9900), .A3(n9899), .A4(n9898), .ZN(n10073) );
  AOI22_X1 U10959 ( .A1(P2_REG2_REG_0__SCAN_IN), .A2(keyinput44), .B1(
        P2_REG1_REG_19__SCAN_IN), .B2(keyinput51), .ZN(n9902) );
  OAI221_X1 U10960 ( .B1(P2_REG2_REG_0__SCAN_IN), .B2(keyinput44), .C1(
        P2_REG1_REG_19__SCAN_IN), .C2(keyinput51), .A(n9902), .ZN(n9909) );
  AOI22_X1 U10961 ( .A1(P2_IR_REG_24__SCAN_IN), .A2(keyinput43), .B1(
        P1_REG2_REG_14__SCAN_IN), .B2(keyinput14), .ZN(n9903) );
  OAI221_X1 U10962 ( .B1(P2_IR_REG_24__SCAN_IN), .B2(keyinput43), .C1(
        P1_REG2_REG_14__SCAN_IN), .C2(keyinput14), .A(n9903), .ZN(n9908) );
  AOI22_X1 U10963 ( .A1(P2_D_REG_11__SCAN_IN), .A2(keyinput21), .B1(
        P1_D_REG_9__SCAN_IN), .B2(keyinput37), .ZN(n9904) );
  OAI221_X1 U10964 ( .B1(P2_D_REG_11__SCAN_IN), .B2(keyinput21), .C1(
        P1_D_REG_9__SCAN_IN), .C2(keyinput37), .A(n9904), .ZN(n9907) );
  AOI22_X1 U10965 ( .A1(P1_DATAO_REG_9__SCAN_IN), .A2(keyinput4), .B1(
        P1_IR_REG_25__SCAN_IN), .B2(keyinput9), .ZN(n9905) );
  OAI221_X1 U10966 ( .B1(P1_DATAO_REG_9__SCAN_IN), .B2(keyinput4), .C1(
        P1_IR_REG_25__SCAN_IN), .C2(keyinput9), .A(n9905), .ZN(n9906) );
  NOR4_X1 U10967 ( .A1(n9909), .A2(n9908), .A3(n9907), .A4(n9906), .ZN(n9938)
         );
  AOI22_X1 U10968 ( .A1(P1_REG0_REG_9__SCAN_IN), .A2(keyinput49), .B1(
        P1_REG3_REG_3__SCAN_IN), .B2(keyinput11), .ZN(n9910) );
  OAI221_X1 U10969 ( .B1(P1_REG0_REG_9__SCAN_IN), .B2(keyinput49), .C1(
        P1_REG3_REG_3__SCAN_IN), .C2(keyinput11), .A(n9910), .ZN(n9917) );
  AOI22_X1 U10970 ( .A1(P1_REG2_REG_19__SCAN_IN), .A2(keyinput23), .B1(SI_5_), 
        .B2(keyinput25), .ZN(n9911) );
  OAI221_X1 U10971 ( .B1(P1_REG2_REG_19__SCAN_IN), .B2(keyinput23), .C1(SI_5_), 
        .C2(keyinput25), .A(n9911), .ZN(n9916) );
  AOI22_X1 U10972 ( .A1(P2_D_REG_14__SCAN_IN), .A2(keyinput27), .B1(
        P1_REG3_REG_28__SCAN_IN), .B2(keyinput62), .ZN(n9912) );
  OAI221_X1 U10973 ( .B1(P2_D_REG_14__SCAN_IN), .B2(keyinput27), .C1(
        P1_REG3_REG_28__SCAN_IN), .C2(keyinput62), .A(n9912), .ZN(n9915) );
  AOI22_X1 U10974 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(keyinput12), .B1(
        P1_D_REG_15__SCAN_IN), .B2(keyinput5), .ZN(n9913) );
  OAI221_X1 U10975 ( .B1(P2_DATAO_REG_0__SCAN_IN), .B2(keyinput12), .C1(
        P1_D_REG_15__SCAN_IN), .C2(keyinput5), .A(n9913), .ZN(n9914) );
  NOR4_X1 U10976 ( .A1(n9917), .A2(n9916), .A3(n9915), .A4(n9914), .ZN(n9937)
         );
  AOI22_X1 U10977 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(keyinput0), .B1(
        P1_DATAO_REG_8__SCAN_IN), .B2(keyinput54), .ZN(n9918) );
  OAI221_X1 U10978 ( .B1(P2_REG1_REG_15__SCAN_IN), .B2(keyinput0), .C1(
        P1_DATAO_REG_8__SCAN_IN), .C2(keyinput54), .A(n9918), .ZN(n9925) );
  AOI22_X1 U10979 ( .A1(P1_REG0_REG_29__SCAN_IN), .A2(keyinput19), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(keyinput20), .ZN(n9919) );
  OAI221_X1 U10980 ( .B1(P1_REG0_REG_29__SCAN_IN), .B2(keyinput19), .C1(
        P2_DATAO_REG_5__SCAN_IN), .C2(keyinput20), .A(n9919), .ZN(n9924) );
  AOI22_X1 U10981 ( .A1(P2_REG1_REG_6__SCAN_IN), .A2(keyinput35), .B1(
        P1_REG0_REG_23__SCAN_IN), .B2(keyinput48), .ZN(n9920) );
  OAI221_X1 U10982 ( .B1(P2_REG1_REG_6__SCAN_IN), .B2(keyinput35), .C1(
        P1_REG0_REG_23__SCAN_IN), .C2(keyinput48), .A(n9920), .ZN(n9923) );
  AOI22_X1 U10983 ( .A1(P2_REG2_REG_26__SCAN_IN), .A2(keyinput3), .B1(
        P1_IR_REG_29__SCAN_IN), .B2(keyinput39), .ZN(n9921) );
  OAI221_X1 U10984 ( .B1(P2_REG2_REG_26__SCAN_IN), .B2(keyinput3), .C1(
        P1_IR_REG_29__SCAN_IN), .C2(keyinput39), .A(n9921), .ZN(n9922) );
  NOR4_X1 U10985 ( .A1(n9925), .A2(n9924), .A3(n9923), .A4(n9922), .ZN(n9936)
         );
  AOI22_X1 U10986 ( .A1(P2_REG2_REG_17__SCAN_IN), .A2(keyinput40), .B1(
        P1_RD_REG_SCAN_IN), .B2(keyinput57), .ZN(n9926) );
  OAI221_X1 U10987 ( .B1(P2_REG2_REG_17__SCAN_IN), .B2(keyinput40), .C1(
        P1_RD_REG_SCAN_IN), .C2(keyinput57), .A(n9926), .ZN(n9934) );
  AOI22_X1 U10988 ( .A1(P2_REG3_REG_26__SCAN_IN), .A2(keyinput41), .B1(
        P1_D_REG_11__SCAN_IN), .B2(keyinput30), .ZN(n9927) );
  OAI221_X1 U10989 ( .B1(P2_REG3_REG_26__SCAN_IN), .B2(keyinput41), .C1(
        P1_D_REG_11__SCAN_IN), .C2(keyinput30), .A(n9927), .ZN(n9933) );
  AOI22_X1 U10990 ( .A1(P1_REG0_REG_21__SCAN_IN), .A2(keyinput63), .B1(
        P1_D_REG_18__SCAN_IN), .B2(keyinput38), .ZN(n9928) );
  OAI221_X1 U10991 ( .B1(P1_REG0_REG_21__SCAN_IN), .B2(keyinput63), .C1(
        P1_D_REG_18__SCAN_IN), .C2(keyinput38), .A(n9928), .ZN(n9932) );
  AOI22_X1 U10992 ( .A1(n9930), .A2(keyinput32), .B1(keyinput46), .B2(n9983), 
        .ZN(n9929) );
  OAI221_X1 U10993 ( .B1(n9930), .B2(keyinput32), .C1(n9983), .C2(keyinput46), 
        .A(n9929), .ZN(n9931) );
  NOR4_X1 U10994 ( .A1(n9934), .A2(n9933), .A3(n9932), .A4(n9931), .ZN(n9935)
         );
  NAND4_X1 U10995 ( .A1(n9938), .A2(n9937), .A3(n9936), .A4(n9935), .ZN(n10072) );
  AOI22_X1 U10996 ( .A1(n9941), .A2(keyinput105), .B1(n9940), .B2(keyinput113), 
        .ZN(n9939) );
  OAI221_X1 U10997 ( .B1(n9941), .B2(keyinput105), .C1(n9940), .C2(keyinput113), .A(n9939), .ZN(n9953) );
  INV_X1 U10998 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n9944) );
  AOI22_X1 U10999 ( .A1(n9944), .A2(keyinput100), .B1(n9943), .B2(keyinput97), 
        .ZN(n9942) );
  OAI221_X1 U11000 ( .B1(n9944), .B2(keyinput100), .C1(n9943), .C2(keyinput97), 
        .A(n9942), .ZN(n9952) );
  AOI22_X1 U11001 ( .A1(n9946), .A2(keyinput98), .B1(n10055), .B2(keyinput120), 
        .ZN(n9945) );
  OAI221_X1 U11002 ( .B1(n9946), .B2(keyinput98), .C1(n10055), .C2(keyinput120), .A(n9945), .ZN(n9951) );
  XOR2_X1 U11003 ( .A(n9947), .B(keyinput65), .Z(n9949) );
  XNOR2_X1 U11004 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(keyinput76), .ZN(n9948) );
  NAND2_X1 U11005 ( .A1(n9949), .A2(n9948), .ZN(n9950) );
  NOR4_X1 U11006 ( .A1(n9953), .A2(n9952), .A3(n9951), .A4(n9950), .ZN(n9998)
         );
  AOI22_X1 U11007 ( .A1(n6202), .A2(keyinput126), .B1(keyinput108), .B2(n9955), 
        .ZN(n9954) );
  OAI221_X1 U11008 ( .B1(n6202), .B2(keyinput126), .C1(n9955), .C2(keyinput108), .A(n9954), .ZN(n9962) );
  AOI22_X1 U11009 ( .A1(n9958), .A2(keyinput83), .B1(n9957), .B2(keyinput84), 
        .ZN(n9956) );
  OAI221_X1 U11010 ( .B1(n9958), .B2(keyinput83), .C1(n9957), .C2(keyinput84), 
        .A(n9956), .ZN(n9961) );
  XNOR2_X1 U11011 ( .A(n9959), .B(keyinput95), .ZN(n9960) );
  OR3_X1 U11012 ( .A1(n9962), .A2(n9961), .A3(n9960), .ZN(n9968) );
  AOI22_X1 U11013 ( .A1(n9964), .A2(keyinput77), .B1(n5710), .B2(keyinput92), 
        .ZN(n9963) );
  OAI221_X1 U11014 ( .B1(n9964), .B2(keyinput77), .C1(n5710), .C2(keyinput92), 
        .A(n9963), .ZN(n9967) );
  XNOR2_X1 U11015 ( .A(n9965), .B(keyinput94), .ZN(n9966) );
  NOR3_X1 U11016 ( .A1(n9968), .A2(n9967), .A3(n9966), .ZN(n9997) );
  AOI22_X1 U11017 ( .A1(n5764), .A2(keyinput75), .B1(keyinput74), .B2(n10047), 
        .ZN(n9969) );
  OAI221_X1 U11018 ( .B1(n5764), .B2(keyinput75), .C1(n10047), .C2(keyinput74), 
        .A(n9969), .ZN(n9980) );
  AOI22_X1 U11019 ( .A1(n10044), .A2(keyinput70), .B1(keyinput99), .B2(n9971), 
        .ZN(n9970) );
  OAI221_X1 U11020 ( .B1(n10044), .B2(keyinput70), .C1(n9971), .C2(keyinput99), 
        .A(n9970), .ZN(n9979) );
  INV_X1 U11021 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n9974) );
  AOI22_X1 U11022 ( .A1(n9974), .A2(keyinput104), .B1(n9973), .B2(keyinput112), 
        .ZN(n9972) );
  OAI221_X1 U11023 ( .B1(n9974), .B2(keyinput104), .C1(n9973), .C2(keyinput112), .A(n9972), .ZN(n9978) );
  XNOR2_X1 U11024 ( .A(P1_REG0_REG_21__SCAN_IN), .B(keyinput127), .ZN(n9976)
         );
  XNOR2_X1 U11025 ( .A(P1_IR_REG_29__SCAN_IN), .B(keyinput103), .ZN(n9975) );
  NAND2_X1 U11026 ( .A1(n9976), .A2(n9975), .ZN(n9977) );
  NOR4_X1 U11027 ( .A1(n9980), .A2(n9979), .A3(n9978), .A4(n9977), .ZN(n9996)
         );
  INV_X1 U11028 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9982) );
  AOI22_X1 U11029 ( .A1(n9983), .A2(keyinput110), .B1(n9982), .B2(keyinput87), 
        .ZN(n9981) );
  OAI221_X1 U11030 ( .B1(n9983), .B2(keyinput110), .C1(n9982), .C2(keyinput87), 
        .A(n9981), .ZN(n9994) );
  AOI22_X1 U11031 ( .A1(n4906), .A2(keyinput107), .B1(keyinput66), .B2(n9985), 
        .ZN(n9984) );
  OAI221_X1 U11032 ( .B1(n4906), .B2(keyinput107), .C1(n9985), .C2(keyinput66), 
        .A(n9984), .ZN(n9993) );
  INV_X1 U11033 ( .A(P2_B_REG_SCAN_IN), .ZN(n9987) );
  AOI22_X1 U11034 ( .A1(n9988), .A2(keyinput81), .B1(keyinput116), .B2(n9987), 
        .ZN(n9986) );
  OAI221_X1 U11035 ( .B1(n9988), .B2(keyinput81), .C1(n9987), .C2(keyinput116), 
        .A(n9986), .ZN(n9992) );
  XNOR2_X1 U11036 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput125), .ZN(n9990) );
  XNOR2_X1 U11037 ( .A(P1_IR_REG_22__SCAN_IN), .B(keyinput82), .ZN(n9989) );
  NAND2_X1 U11038 ( .A1(n9990), .A2(n9989), .ZN(n9991) );
  NOR4_X1 U11039 ( .A1(n9994), .A2(n9993), .A3(n9992), .A4(n9991), .ZN(n9995)
         );
  NAND4_X1 U11040 ( .A1(n9998), .A2(n9997), .A3(n9996), .A4(n9995), .ZN(n10070) );
  AOI22_X1 U11041 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(keyinput122), .B1(SI_11_), .B2(keyinput86), .ZN(n9999) );
  OAI221_X1 U11042 ( .B1(P2_REG3_REG_14__SCAN_IN), .B2(keyinput122), .C1(
        SI_11_), .C2(keyinput86), .A(n9999), .ZN(n10006) );
  AOI22_X1 U11043 ( .A1(P2_REG0_REG_4__SCAN_IN), .A2(keyinput96), .B1(
        P2_IR_REG_19__SCAN_IN), .B2(keyinput88), .ZN(n10000) );
  OAI221_X1 U11044 ( .B1(P2_REG0_REG_4__SCAN_IN), .B2(keyinput96), .C1(
        P2_IR_REG_19__SCAN_IN), .C2(keyinput88), .A(n10000), .ZN(n10005) );
  AOI22_X1 U11045 ( .A1(P2_D_REG_14__SCAN_IN), .A2(keyinput91), .B1(
        P1_IR_REG_25__SCAN_IN), .B2(keyinput73), .ZN(n10001) );
  OAI221_X1 U11046 ( .B1(P2_D_REG_14__SCAN_IN), .B2(keyinput91), .C1(
        P1_IR_REG_25__SCAN_IN), .C2(keyinput73), .A(n10001), .ZN(n10004) );
  AOI22_X1 U11047 ( .A1(P2_REG2_REG_26__SCAN_IN), .A2(keyinput67), .B1(
        P1_D_REG_15__SCAN_IN), .B2(keyinput69), .ZN(n10002) );
  OAI221_X1 U11048 ( .B1(P2_REG2_REG_26__SCAN_IN), .B2(keyinput67), .C1(
        P1_D_REG_15__SCAN_IN), .C2(keyinput69), .A(n10002), .ZN(n10003) );
  NOR4_X1 U11049 ( .A1(n10006), .A2(n10005), .A3(n10004), .A4(n10003), .ZN(
        n10038) );
  AOI22_X1 U11050 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(keyinput114), .B1(
        P1_REG2_REG_14__SCAN_IN), .B2(keyinput78), .ZN(n10007) );
  OAI221_X1 U11051 ( .B1(P2_IR_REG_9__SCAN_IN), .B2(keyinput114), .C1(
        P1_REG2_REG_14__SCAN_IN), .C2(keyinput78), .A(n10007), .ZN(n10014) );
  AOI22_X1 U11052 ( .A1(P1_ADDR_REG_12__SCAN_IN), .A2(keyinput72), .B1(SI_5_), 
        .B2(keyinput89), .ZN(n10008) );
  OAI221_X1 U11053 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(keyinput72), .C1(SI_5_), 
        .C2(keyinput89), .A(n10008), .ZN(n10013) );
  AOI22_X1 U11054 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(keyinput64), .B1(
        P1_RD_REG_SCAN_IN), .B2(keyinput121), .ZN(n10009) );
  OAI221_X1 U11055 ( .B1(P2_REG1_REG_15__SCAN_IN), .B2(keyinput64), .C1(
        P1_RD_REG_SCAN_IN), .C2(keyinput121), .A(n10009), .ZN(n10012) );
  AOI22_X1 U11056 ( .A1(P2_D_REG_6__SCAN_IN), .A2(keyinput124), .B1(
        P1_D_REG_28__SCAN_IN), .B2(keyinput71), .ZN(n10010) );
  OAI221_X1 U11057 ( .B1(P2_D_REG_6__SCAN_IN), .B2(keyinput124), .C1(
        P1_D_REG_28__SCAN_IN), .C2(keyinput71), .A(n10010), .ZN(n10011) );
  NOR4_X1 U11058 ( .A1(n10014), .A2(n10013), .A3(n10012), .A4(n10011), .ZN(
        n10037) );
  AOI22_X1 U11059 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(keyinput80), .B1(
        P1_REG1_REG_4__SCAN_IN), .B2(keyinput93), .ZN(n10015) );
  OAI221_X1 U11060 ( .B1(P2_REG3_REG_11__SCAN_IN), .B2(keyinput80), .C1(
        P1_REG1_REG_4__SCAN_IN), .C2(keyinput93), .A(n10015), .ZN(n10026) );
  AOI22_X1 U11061 ( .A1(P1_REG1_REG_2__SCAN_IN), .A2(keyinput119), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(keyinput68), .ZN(n10016) );
  OAI221_X1 U11062 ( .B1(P1_REG1_REG_2__SCAN_IN), .B2(keyinput119), .C1(
        P1_DATAO_REG_9__SCAN_IN), .C2(keyinput68), .A(n10016), .ZN(n10025) );
  AOI22_X1 U11063 ( .A1(n10019), .A2(keyinput102), .B1(n10018), .B2(
        keyinput101), .ZN(n10017) );
  OAI221_X1 U11064 ( .B1(n10019), .B2(keyinput102), .C1(n10018), .C2(
        keyinput101), .A(n10017), .ZN(n10024) );
  AOI22_X1 U11065 ( .A1(n10022), .A2(keyinput85), .B1(keyinput106), .B2(n10021), .ZN(n10020) );
  OAI221_X1 U11066 ( .B1(n10022), .B2(keyinput85), .C1(n10021), .C2(
        keyinput106), .A(n10020), .ZN(n10023) );
  NOR4_X1 U11067 ( .A1(n10026), .A2(n10025), .A3(n10024), .A4(n10023), .ZN(
        n10036) );
  AOI22_X1 U11068 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(keyinput109), .B1(
        P2_D_REG_15__SCAN_IN), .B2(keyinput111), .ZN(n10027) );
  OAI221_X1 U11069 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(keyinput109), .C1(
        P2_D_REG_15__SCAN_IN), .C2(keyinput111), .A(n10027), .ZN(n10034) );
  AOI22_X1 U11070 ( .A1(P2_REG1_REG_19__SCAN_IN), .A2(keyinput115), .B1(
        P1_DATAO_REG_8__SCAN_IN), .B2(keyinput118), .ZN(n10028) );
  OAI221_X1 U11071 ( .B1(P2_REG1_REG_19__SCAN_IN), .B2(keyinput115), .C1(
        P1_DATAO_REG_8__SCAN_IN), .C2(keyinput118), .A(n10028), .ZN(n10033) );
  AOI22_X1 U11072 ( .A1(P2_REG2_REG_8__SCAN_IN), .A2(keyinput123), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(keyinput79), .ZN(n10029) );
  OAI221_X1 U11073 ( .B1(P2_REG2_REG_8__SCAN_IN), .B2(keyinput123), .C1(
        P2_DATAO_REG_6__SCAN_IN), .C2(keyinput79), .A(n10029), .ZN(n10032) );
  AOI22_X1 U11074 ( .A1(P1_REG2_REG_11__SCAN_IN), .A2(keyinput117), .B1(
        P1_IR_REG_2__SCAN_IN), .B2(keyinput90), .ZN(n10030) );
  OAI221_X1 U11075 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(keyinput117), .C1(
        P1_IR_REG_2__SCAN_IN), .C2(keyinput90), .A(n10030), .ZN(n10031) );
  NOR4_X1 U11076 ( .A1(n10034), .A2(n10033), .A3(n10032), .A4(n10031), .ZN(
        n10035) );
  NAND4_X1 U11077 ( .A1(n10038), .A2(n10037), .A3(n10036), .A4(n10035), .ZN(
        n10069) );
  AOI22_X1 U11078 ( .A1(n10041), .A2(keyinput15), .B1(keyinput29), .B2(n10040), 
        .ZN(n10039) );
  OAI221_X1 U11079 ( .B1(n10041), .B2(keyinput15), .C1(n10040), .C2(keyinput29), .A(n10039), .ZN(n10053) );
  AOI22_X1 U11080 ( .A1(n10044), .A2(keyinput6), .B1(keyinput60), .B2(n10043), 
        .ZN(n10042) );
  OAI221_X1 U11081 ( .B1(n10044), .B2(keyinput6), .C1(n10043), .C2(keyinput60), 
        .A(n10042), .ZN(n10052) );
  INV_X1 U11082 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n10046) );
  AOI22_X1 U11083 ( .A1(n10047), .A2(keyinput10), .B1(keyinput8), .B2(n10046), 
        .ZN(n10045) );
  OAI221_X1 U11084 ( .B1(n10047), .B2(keyinput10), .C1(n10046), .C2(keyinput8), 
        .A(n10045), .ZN(n10051) );
  XNOR2_X1 U11085 ( .A(P2_IR_REG_3__SCAN_IN), .B(keyinput36), .ZN(n10049) );
  XNOR2_X1 U11086 ( .A(P1_REG1_REG_2__SCAN_IN), .B(keyinput55), .ZN(n10048) );
  NAND2_X1 U11087 ( .A1(n10049), .A2(n10048), .ZN(n10050) );
  NOR4_X1 U11088 ( .A1(n10053), .A2(n10052), .A3(n10051), .A4(n10050), .ZN(
        n10068) );
  AOI22_X1 U11089 ( .A1(n10056), .A2(keyinput47), .B1(n10055), .B2(keyinput56), 
        .ZN(n10054) );
  OAI221_X1 U11090 ( .B1(n10056), .B2(keyinput47), .C1(n10055), .C2(keyinput56), .A(n10054), .ZN(n10066) );
  AOI22_X1 U11091 ( .A1(n10059), .A2(keyinput58), .B1(n10058), .B2(keyinput22), 
        .ZN(n10057) );
  OAI221_X1 U11092 ( .B1(n10059), .B2(keyinput58), .C1(n10058), .C2(keyinput22), .A(n10057), .ZN(n10065) );
  XNOR2_X1 U11093 ( .A(P2_B_REG_SCAN_IN), .B(keyinput52), .ZN(n10063) );
  XNOR2_X1 U11094 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput61), .ZN(n10062) );
  XNOR2_X1 U11095 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(keyinput17), .ZN(n10061)
         );
  XNOR2_X1 U11096 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput31), .ZN(n10060) );
  NAND4_X1 U11097 ( .A1(n10063), .A2(n10062), .A3(n10061), .A4(n10060), .ZN(
        n10064) );
  NOR3_X1 U11098 ( .A1(n10066), .A2(n10065), .A3(n10064), .ZN(n10067) );
  OAI211_X1 U11099 ( .C1(n10070), .C2(n10069), .A(n10068), .B(n10067), .ZN(
        n10071) );
  NOR4_X1 U11100 ( .A1(n10074), .A2(n10073), .A3(n10072), .A4(n10071), .ZN(
        n10078) );
  MUX2_X1 U11101 ( .A(n10076), .B(n10075), .S(P2_U3966), .Z(n10077) );
  XNOR2_X1 U11102 ( .A(n10078), .B(n10077), .ZN(P2_U3574) );
  XOR2_X1 U11103 ( .A(n10079), .B(P2_ADDR_REG_7__SCAN_IN), .Z(ADD_1071_U49) );
  AOI21_X1 U11104 ( .B1(n10082), .B2(n10081), .A(n10080), .ZN(ADD_1071_U47) );
  XOR2_X1 U11105 ( .A(n10083), .B(P2_ADDR_REG_6__SCAN_IN), .Z(ADD_1071_U50) );
  NOR2_X1 U11106 ( .A1(n10085), .A2(n10084), .ZN(n10086) );
  XOR2_X1 U11107 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n10086), .Z(ADD_1071_U51) );
  OAI21_X1 U11108 ( .B1(n10089), .B2(n10088), .A(n10087), .ZN(n10090) );
  XNOR2_X1 U11109 ( .A(n10090), .B(P1_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  XOR2_X1 U11110 ( .A(n10092), .B(n10091), .Z(ADD_1071_U54) );
  XOR2_X1 U11111 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n10093), .Z(ADD_1071_U48) );
  XOR2_X1 U11112 ( .A(n10095), .B(n10094), .Z(ADD_1071_U53) );
  XNOR2_X1 U11113 ( .A(n10097), .B(n10096), .ZN(ADD_1071_U52) );
  INV_X1 U4823 ( .A(n4987), .ZN(n8171) );
  INV_X2 U4853 ( .A(n4986), .ZN(n5115) );
  CLKBUF_X1 U4855 ( .A(n4973), .Z(n4318) );
  INV_X2 U4869 ( .A(n7304), .ZN(n6212) );
  AND2_X1 U4870 ( .A1(n4434), .A2(n4433), .ZN(n4432) );
  CLKBUF_X1 U4924 ( .A(n5213), .Z(n8037) );
  NAND2_X1 U5921 ( .A1(n6875), .A2(n5655), .ZN(n4987) );
  NAND2_X1 U6019 ( .A1(n7639), .A2(n7638), .ZN(n7692) );
endmodule

