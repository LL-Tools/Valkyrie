

module b21_C_gen_AntiSAT_k_256_9 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2, 
        keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7, 
        keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12, 
        keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17, 
        keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22, 
        keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27, 
        keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32, 
        keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37, 
        keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42, 
        keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47, 
        keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52, 
        keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57, 
        keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62, 
        keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66, keyinput_f67, 
        keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71, keyinput_f72, 
        keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76, keyinput_f77, 
        keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81, keyinput_f82, 
        keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86, keyinput_f87, 
        keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91, keyinput_f92, 
        keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96, keyinput_f97, 
        keyinput_f98, keyinput_f99, keyinput_f100, keyinput_f101, 
        keyinput_f102, keyinput_f103, keyinput_f104, keyinput_f105, 
        keyinput_f106, keyinput_f107, keyinput_f108, keyinput_f109, 
        keyinput_f110, keyinput_f111, keyinput_f112, keyinput_f113, 
        keyinput_f114, keyinput_f115, keyinput_f116, keyinput_f117, 
        keyinput_f118, keyinput_f119, keyinput_f120, keyinput_f121, 
        keyinput_f122, keyinput_f123, keyinput_f124, keyinput_f125, 
        keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, keyinput_g2, 
        keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, 
        keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, 
        keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, 
        keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, 
        keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, 
        keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, 
        keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, 
        keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, 
        keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, 
        keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, 
        keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, 
        keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, 
        keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, keyinput_g67, 
        keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, keyinput_g72, 
        keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, keyinput_g77, 
        keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, keyinput_g82, 
        keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, keyinput_g87, 
        keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, keyinput_g92, 
        keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, keyinput_g97, 
        keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101, 
        keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105, 
        keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109, 
        keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113, 
        keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117, 
        keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121, 
        keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125, 
        keyinput_g126, keyinput_g127, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, 
        ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, 
        ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, 
        ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, 
        ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, 
        P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, 
        P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, 
        P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, 
        P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, 
        P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, 
        P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, 
        P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, 
        P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, 
        P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, 
        P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, 
        P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, 
        P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, 
        P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, 
        P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, 
        P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, 
        P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, 
        P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, 
        P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, 
        P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, 
        P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, 
        P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, 
        P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, 
        P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, 
        P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, 
        P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, 
        P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, 
        P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, 
        P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, 
        P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, 
        P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, 
        P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, 
        P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, 
        P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, 
        P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, 
        P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, 
        P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, 
        P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, 
        P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, 
        P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, 
        P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, 
        P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, 
        P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, 
        P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, 
        P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3152, P2_U3151, P2_U3966 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66, keyinput_f67,
         keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71, keyinput_f72,
         keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76, keyinput_f77,
         keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81, keyinput_f82,
         keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86, keyinput_f87,
         keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91, keyinput_f92,
         keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96, keyinput_f97,
         keyinput_f98, keyinput_f99, keyinput_f100, keyinput_f101,
         keyinput_f102, keyinput_f103, keyinput_f104, keyinput_f105,
         keyinput_f106, keyinput_f107, keyinput_f108, keyinput_f109,
         keyinput_f110, keyinput_f111, keyinput_f112, keyinput_f113,
         keyinput_f114, keyinput_f115, keyinput_f116, keyinput_f117,
         keyinput_f118, keyinput_f119, keyinput_f120, keyinput_f121,
         keyinput_f122, keyinput_f123, keyinput_f124, keyinput_f125,
         keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, keyinput_g2,
         keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7,
         keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12,
         keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17,
         keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22,
         keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27,
         keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32,
         keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37,
         keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42,
         keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47,
         keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52,
         keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57,
         keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62,
         keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, keyinput_g67,
         keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, keyinput_g72,
         keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, keyinput_g77,
         keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, keyinput_g82,
         keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, keyinput_g87,
         keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, keyinput_g92,
         keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, keyinput_g97,
         keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101,
         keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105,
         keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109,
         keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113,
         keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117,
         keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121,
         keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125,
         keyinput_g126, keyinput_g127;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
         n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
         n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
         n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
         n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
         n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
         n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
         n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
         n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861,
         n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871,
         n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881,
         n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
         n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901,
         n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
         n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
         n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931,
         n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941,
         n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951,
         n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961,
         n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971,
         n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981,
         n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991,
         n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001,
         n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011,
         n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021,
         n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031,
         n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041,
         n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051,
         n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061,
         n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071,
         n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081,
         n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091,
         n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101,
         n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111,
         n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121,
         n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131,
         n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141,
         n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151,
         n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161,
         n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171,
         n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181,
         n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191,
         n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201,
         n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211,
         n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221,
         n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231,
         n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241,
         n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251,
         n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261,
         n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271,
         n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281,
         n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291,
         n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301,
         n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311,
         n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321,
         n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331,
         n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341,
         n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351,
         n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361,
         n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371,
         n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381,
         n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391,
         n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401,
         n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411,
         n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421,
         n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431,
         n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441,
         n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451,
         n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461,
         n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471,
         n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481,
         n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491,
         n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501,
         n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511,
         n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521,
         n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531,
         n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541,
         n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551,
         n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561,
         n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571,
         n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581,
         n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591,
         n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601,
         n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611,
         n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621,
         n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631,
         n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641,
         n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651,
         n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661,
         n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671,
         n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681,
         n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691,
         n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701,
         n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711,
         n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721,
         n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731,
         n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741,
         n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751,
         n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761,
         n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771,
         n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781,
         n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791,
         n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801,
         n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811,
         n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821,
         n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831,
         n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841,
         n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851,
         n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861,
         n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871,
         n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881,
         n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891,
         n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901,
         n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911,
         n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921,
         n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931,
         n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941,
         n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951,
         n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961,
         n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971,
         n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981,
         n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991,
         n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001,
         n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011,
         n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021,
         n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031,
         n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041,
         n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051,
         n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061,
         n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071,
         n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081,
         n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091,
         n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101,
         n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111,
         n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121,
         n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131,
         n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141,
         n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151,
         n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161,
         n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171,
         n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181,
         n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191,
         n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201,
         n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211,
         n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221,
         n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231,
         n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241,
         n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251,
         n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261,
         n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271,
         n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281,
         n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291,
         n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301,
         n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311,
         n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321,
         n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331,
         n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341,
         n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351,
         n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361,
         n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371,
         n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381,
         n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391,
         n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401,
         n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411,
         n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421,
         n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431,
         n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441,
         n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451,
         n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461,
         n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471,
         n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481,
         n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491,
         n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501,
         n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511,
         n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521,
         n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531,
         n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541,
         n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551,
         n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561,
         n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571,
         n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581,
         n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591,
         n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601,
         n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611,
         n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621,
         n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631,
         n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641,
         n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651,
         n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661,
         n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671,
         n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681,
         n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691,
         n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701,
         n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711,
         n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721,
         n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731,
         n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741,
         n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751,
         n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761,
         n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771,
         n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781,
         n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791,
         n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801,
         n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811,
         n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821,
         n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831,
         n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841,
         n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851,
         n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861,
         n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871,
         n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881,
         n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891,
         n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901,
         n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911,
         n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921,
         n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931,
         n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941,
         n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951,
         n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961,
         n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971,
         n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981,
         n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991,
         n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001,
         n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011,
         n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021,
         n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031,
         n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041,
         n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051,
         n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061,
         n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071,
         n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081,
         n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091,
         n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101,
         n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111,
         n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121,
         n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131,
         n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141,
         n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151,
         n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161,
         n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171,
         n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181,
         n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191,
         n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201,
         n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211,
         n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221,
         n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231,
         n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241,
         n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251,
         n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261,
         n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271,
         n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281,
         n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291,
         n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301,
         n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311,
         n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321,
         n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331,
         n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341,
         n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351,
         n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361,
         n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371,
         n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381,
         n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391,
         n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401,
         n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411,
         n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421,
         n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431,
         n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441,
         n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451,
         n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461,
         n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471,
         n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481,
         n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491,
         n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501,
         n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511,
         n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521,
         n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531,
         n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541,
         n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551,
         n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561,
         n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571,
         n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581,
         n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591,
         n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601,
         n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611,
         n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621,
         n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631,
         n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641,
         n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651,
         n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661,
         n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671,
         n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681,
         n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691,
         n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701,
         n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711,
         n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721,
         n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731,
         n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741,
         n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751,
         n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761,
         n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771,
         n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781,
         n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791,
         n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801,
         n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811,
         n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821,
         n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831,
         n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841,
         n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851,
         n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861,
         n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871,
         n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881,
         n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891,
         n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901,
         n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911,
         n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921,
         n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931,
         n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941,
         n7942, n7943, n7944, n7945, n7946, n7947, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073,
         n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083,
         n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093,
         n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103,
         n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113,
         n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123,
         n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133,
         n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143,
         n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153,
         n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163,
         n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173,
         n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183,
         n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193,
         n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203,
         n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213,
         n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223,
         n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233,
         n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243,
         n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253,
         n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263,
         n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273,
         n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283,
         n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293,
         n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303,
         n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313,
         n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323,
         n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333,
         n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343,
         n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353,
         n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363,
         n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373,
         n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383,
         n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393,
         n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403,
         n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413,
         n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423,
         n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433,
         n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443,
         n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453,
         n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463,
         n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473,
         n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483,
         n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493,
         n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503,
         n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513,
         n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523,
         n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533,
         n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543,
         n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553,
         n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563,
         n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573,
         n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583,
         n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593,
         n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603,
         n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613,
         n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623,
         n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633,
         n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643,
         n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653,
         n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663,
         n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673,
         n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683,
         n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693,
         n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703,
         n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713,
         n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723,
         n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733,
         n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743,
         n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753,
         n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763,
         n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773,
         n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783,
         n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793,
         n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803,
         n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813,
         n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823,
         n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833,
         n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843,
         n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853,
         n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863,
         n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873,
         n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883,
         n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893,
         n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903,
         n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913,
         n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923,
         n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933,
         n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943,
         n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953,
         n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963,
         n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973,
         n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983,
         n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993,
         n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003,
         n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013,
         n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023,
         n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033,
         n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043,
         n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053,
         n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063,
         n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073,
         n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083,
         n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093,
         n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103,
         n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113,
         n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123,
         n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133,
         n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143,
         n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153,
         n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163,
         n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173,
         n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183,
         n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193,
         n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203,
         n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213,
         n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223,
         n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233,
         n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243,
         n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253,
         n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263,
         n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273,
         n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283,
         n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293,
         n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303,
         n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313,
         n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323,
         n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333,
         n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343,
         n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353,
         n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363,
         n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373,
         n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383,
         n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393,
         n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403,
         n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413,
         n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423,
         n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433,
         n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443,
         n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453,
         n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463,
         n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473,
         n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483,
         n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493,
         n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503,
         n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513,
         n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523,
         n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533,
         n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543,
         n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553,
         n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563,
         n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573,
         n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583,
         n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593,
         n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603,
         n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613,
         n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623,
         n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633,
         n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643,
         n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653,
         n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663,
         n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673,
         n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683,
         n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693,
         n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703,
         n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713,
         n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723,
         n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733,
         n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743,
         n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753,
         n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763,
         n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773,
         n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783,
         n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793,
         n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803,
         n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813,
         n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823,
         n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833,
         n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843,
         n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853,
         n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863,
         n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873,
         n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883,
         n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893,
         n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903,
         n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913,
         n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923,
         n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933,
         n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943,
         n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953,
         n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963,
         n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973,
         n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983,
         n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993,
         n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002,
         n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010,
         n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018,
         n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026,
         n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034,
         n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042,
         n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050,
         n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058,
         n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066,
         n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074,
         n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082,
         n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090,
         n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098,
         n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106,
         n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114,
         n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122,
         n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130,
         n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138,
         n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146,
         n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154,
         n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162,
         n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170,
         n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178,
         n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186,
         n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194,
         n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202,
         n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210,
         n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218,
         n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226,
         n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234,
         n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242,
         n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250,
         n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258,
         n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266,
         n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274,
         n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282,
         n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290,
         n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298,
         n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306,
         n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314,
         n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322,
         n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330,
         n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338,
         n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346,
         n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354,
         n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362,
         n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370,
         n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378,
         n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386,
         n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394,
         n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402,
         n10403, n10404, n10405, n10406, n10407;

  INV_X1 U4987 ( .A(n7953), .ZN(n8156) );
  INV_X1 U4988 ( .A(n6062), .ZN(n6351) );
  NAND2_X2 U4989 ( .A1(n5111), .A2(n8873), .ZN(n5641) );
  CLKBUF_X2 U4990 ( .A(n6035), .Z(n6288) );
  OR2_X1 U4991 ( .A1(n7416), .A2(n8226), .ZN(n10245) );
  BUF_X1 U4992 ( .A(n10283), .Z(n4581) );
  INV_X1 U4993 ( .A(n7546), .ZN(n6712) );
  OAI21_X1 U4994 ( .B1(n5594), .B2(n5593), .A(n5592), .ZN(n5595) );
  INV_X1 U4996 ( .A(n8168), .ZN(n8243) );
  INV_X1 U4998 ( .A(n7338), .ZN(n7034) );
  AND2_X1 U4999 ( .A1(n5120), .A2(n5095), .ZN(n5163) );
  AND2_X2 U5000 ( .A1(n6788), .A2(n6537), .ZN(n6608) );
  INV_X1 U5002 ( .A(n9348), .ZN(n9349) );
  OR2_X1 U5003 ( .A1(n7804), .A2(n7812), .ZN(n7806) );
  NAND2_X1 U5004 ( .A1(n8965), .A2(n8969), .ZN(n8891) );
  AND4_X1 U5005 ( .A1(n6059), .A2(n6058), .A3(n6057), .A4(n6056), .ZN(n7539)
         );
  OAI21_X1 U5006 ( .B1(n9086), .B2(n9237), .A(n9088), .ZN(n9194) );
  NAND2_X1 U5007 ( .A1(n9483), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5926) );
  INV_X1 U5008 ( .A(n10138), .ZN(n9203) );
  AOI21_X1 U5009 ( .B1(n5391), .B2(n4991), .A(n4988), .ZN(n4987) );
  NOR2_X4 U5010 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n6020) );
  OR2_X2 U5011 ( .A1(n8153), .A2(n5954), .ZN(n6035) );
  XNOR2_X2 U5012 ( .A(n6371), .B(n6370), .ZN(n7577) );
  XNOR2_X2 U5013 ( .A(n5117), .B(n5116), .ZN(n7089) );
  OAI21_X2 U5014 ( .B1(n5881), .B2(n4506), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n5117) );
  BUF_X8 U5015 ( .A(n5159), .Z(n4483) );
  NAND2_X2 U5016 ( .A1(n4698), .A2(n4697), .ZN(n5159) );
  NAND2_X1 U5017 ( .A1(n5994), .A2(n5993), .ZN(n9452) );
  NAND2_X2 U5018 ( .A1(n10249), .A2(n5711), .ZN(n7444) );
  NAND2_X1 U5019 ( .A1(n6544), .A2(n7322), .ZN(n7245) );
  NAND2_X1 U5020 ( .A1(n5721), .A2(n5720), .ZN(n7367) );
  INV_X1 U5021 ( .A(n10259), .ZN(n10317) );
  CLKBUF_X1 U5022 ( .A(n6037), .Z(n4486) );
  INV_X1 U5023 ( .A(n7322), .ZN(n6542) );
  INV_X1 U5024 ( .A(n6047), .ZN(n6037) );
  INV_X1 U5025 ( .A(n10244), .ZN(n10308) );
  INV_X2 U5026 ( .A(n5657), .ZN(n5676) );
  INV_X4 U5027 ( .A(n6608), .ZN(n6727) );
  AOI21_X1 U5028 ( .B1(n8881), .B2(n8879), .A(n8878), .ZN(n6786) );
  AND2_X1 U5029 ( .A1(n4711), .A2(n4710), .ZN(n8881) );
  NAND2_X1 U5030 ( .A1(n4609), .A2(n4608), .ZN(n4711) );
  OAI22_X1 U5031 ( .A1(n9296), .A2(n9079), .B1(n9302), .B2(n9078), .ZN(n9281)
         );
  NAND2_X1 U5032 ( .A1(n9196), .A2(n9197), .ZN(n9195) );
  NAND2_X1 U5033 ( .A1(n5695), .A2(n5694), .ZN(n8744) );
  OAI21_X1 U5034 ( .B1(n8068), .B2(n4713), .A(n4712), .ZN(n8998) );
  NOR2_X1 U5035 ( .A1(n9233), .A2(n9232), .ZN(n9231) );
  NAND2_X1 U5036 ( .A1(n7938), .A2(n6623), .ZN(n8068) );
  NAND2_X1 U5037 ( .A1(n5047), .A2(n4521), .ZN(n7938) );
  NAND2_X1 U5038 ( .A1(n8031), .A2(n8030), .ZN(n9069) );
  AOI21_X1 U5039 ( .B1(n8662), .B2(n5017), .A(n5015), .ZN(n5014) );
  NAND2_X1 U5040 ( .A1(n7988), .A2(n7987), .ZN(n8031) );
  AOI21_X1 U5041 ( .B1(n9287), .B2(n9112), .A(n9111), .ZN(n9274) );
  NAND2_X2 U5042 ( .A1(n5634), .A2(n5633), .ZN(n8755) );
  AOI21_X1 U5043 ( .B1(n9311), .B2(n9108), .A(n9107), .ZN(n9303) );
  XNOR2_X1 U5044 ( .A(n5647), .B(n5646), .ZN(n8150) );
  NAND2_X1 U5045 ( .A1(n5632), .A2(n5631), .ZN(n5647) );
  NAND2_X1 U5046 ( .A1(n5016), .A2(n5084), .ZN(n5015) );
  NAND2_X1 U5047 ( .A1(n7627), .A2(n7626), .ZN(n10203) );
  AND2_X1 U5048 ( .A1(n4799), .A2(n4798), .ZN(n7627) );
  NAND2_X1 U5049 ( .A1(n7542), .A2(n6385), .ZN(n10179) );
  NAND2_X1 U5050 ( .A1(n6217), .A2(n6216), .ZN(n9925) );
  NAND2_X1 U5051 ( .A1(n5378), .A2(n5377), .ZN(n8111) );
  NAND2_X1 U5052 ( .A1(n6188), .A2(n6187), .ZN(n9932) );
  INV_X1 U5053 ( .A(n7239), .ZN(n10126) );
  INV_X2 U5054 ( .A(n10263), .ZN(n10266) );
  OR2_X1 U5055 ( .A1(n5325), .A2(n4975), .ZN(n4974) );
  NAND2_X2 U5056 ( .A1(n7229), .A2(n8620), .ZN(n10263) );
  NAND2_X2 U5057 ( .A1(n7534), .A2(n10151), .ZN(n10143) );
  NAND4_X1 U5058 ( .A1(n6041), .A2(n6040), .A3(n6039), .A4(n6038), .ZN(n9021)
         );
  INV_X2 U5059 ( .A(n4487), .ZN(n6358) );
  CLKBUF_X1 U5060 ( .A(n6037), .Z(n4487) );
  BUF_X2 U5061 ( .A(n6023), .Z(n6276) );
  NAND2_X1 U5062 ( .A1(n5842), .A2(n5843), .ZN(n7329) );
  NAND2_X1 U5063 ( .A1(n5955), .A2(n5954), .ZN(n6034) );
  OR2_X1 U5064 ( .A1(n6035), .A2(n6859), .ZN(n6016) );
  OR2_X1 U5065 ( .A1(n6032), .A2(n6014), .ZN(n6015) );
  INV_X1 U5066 ( .A(n7352), .ZN(n6538) );
  OAI211_X1 U5067 ( .C1(n6117), .C2(n6881), .A(n6055), .B(n6054), .ZN(n7322)
         );
  NAND3_X1 U5068 ( .A1(n5183), .A2(n5182), .A3(n4508), .ZN(n10244) );
  NAND2_X2 U5069 ( .A1(n7266), .A2(n6539), .ZN(n7546) );
  OAI211_X1 U5070 ( .C1(n5142), .C2(n7079), .A(n5133), .B(n5132), .ZN(n7338)
         );
  AND2_X2 U5071 ( .A1(n6788), .A2(n7266), .ZN(n6759) );
  NAND2_X1 U5072 ( .A1(n6478), .A2(n6737), .ZN(n6788) );
  NAND2_X1 U5074 ( .A1(n7247), .A2(n7524), .ZN(n7266) );
  NAND2_X2 U5075 ( .A1(n6480), .A2(n6481), .ZN(n6117) );
  XNOR2_X1 U5076 ( .A(n6477), .B(P1_IR_REG_26__SCAN_IN), .ZN(n6737) );
  XNOR2_X1 U5077 ( .A(n5928), .B(P1_IR_REG_29__SCAN_IN), .ZN(n5954) );
  XNOR2_X1 U5078 ( .A(n5914), .B(n5921), .ZN(n6480) );
  INV_X1 U5079 ( .A(n7577), .ZN(n7247) );
  XNOR2_X1 U5080 ( .A(n6475), .B(n6474), .ZN(n7952) );
  NAND2_X1 U5081 ( .A1(n6470), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6475) );
  AND2_X1 U5082 ( .A1(n5908), .A2(n5907), .ZN(n5910) );
  AND2_X1 U5083 ( .A1(n4792), .A2(n5908), .ZN(n4791) );
  AND2_X1 U5084 ( .A1(n5907), .A2(n6472), .ZN(n4792) );
  AND2_X1 U5085 ( .A1(n4494), .A2(n6468), .ZN(n5071) );
  NAND2_X1 U5086 ( .A1(n5141), .A2(n4783), .ZN(n7107) );
  NOR2_X1 U5087 ( .A1(n5906), .A2(n5905), .ZN(n5907) );
  AND4_X1 U5088 ( .A1(n5099), .A2(n5335), .A3(n5251), .A4(n5252), .ZN(n5044)
         );
  AND4_X1 U5089 ( .A1(n5097), .A2(n5098), .A3(n5100), .A4(n5096), .ZN(n5045)
         );
  AND4_X1 U5090 ( .A1(n5897), .A2(n5896), .A3(n5895), .A4(n6060), .ZN(n5900)
         );
  AND2_X1 U5091 ( .A1(n5909), .A2(n5073), .ZN(n5072) );
  INV_X1 U5092 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5990) );
  INV_X1 U5093 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5251) );
  INV_X2 U5094 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  NOR2_X1 U5095 ( .A1(P1_ADDR_REG_19__SCAN_IN), .A2(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n9889) );
  NOR2_X2 U5096 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5120) );
  INV_X4 U5097 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  INV_X1 U5098 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5252) );
  INV_X1 U5099 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5898) );
  NOR2_X1 U5100 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n5099) );
  NOR2_X1 U5101 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n5895) );
  NOR2_X1 U5102 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n5896) );
  NOR2_X1 U5103 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n5897) );
  NOR2_X1 U5104 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n5096) );
  NOR2_X1 U5105 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n5100) );
  NOR2_X1 U5106 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n5098) );
  INV_X1 U5107 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n5986) );
  INV_X1 U5108 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n6183) );
  INV_X1 U5109 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n9723) );
  NAND2_X1 U5110 ( .A1(n6117), .A2(n4483), .ZN(n4484) );
  NAND2_X1 U5111 ( .A1(n6117), .A2(n4483), .ZN(n6062) );
  XNOR2_X2 U5112 ( .A(n9021), .B(n6563), .ZN(n7393) );
  AND4_X4 U5113 ( .A1(n6051), .A2(n6050), .A3(n6049), .A4(n6048), .ZN(n6544)
         );
  OR2_X1 U5114 ( .A1(n6288), .A2(n6880), .ZN(n6049) );
  NAND2_X1 U5115 ( .A1(n5955), .A2(n5954), .ZN(n4485) );
  XNOR2_X2 U5116 ( .A(n6552), .B(n10160), .ZN(n7239) );
  XNOR2_X2 U5117 ( .A(n5926), .B(n5925), .ZN(n8153) );
  NAND2_X1 U5118 ( .A1(n5280), .A2(n5279), .ZN(n5295) );
  INV_X1 U5119 ( .A(n8873), .ZN(n5110) );
  NAND2_X1 U5120 ( .A1(n9186), .A2(n9092), .ZN(n4842) );
  NAND2_X1 U5121 ( .A1(n9416), .A2(n9092), .ZN(n6376) );
  OR2_X1 U5122 ( .A1(n9442), .A2(n9276), .ZN(n9081) );
  OR2_X1 U5123 ( .A1(n4809), .A2(n4807), .ZN(n4806) );
  NAND2_X1 U5124 ( .A1(n8153), .A2(n5954), .ZN(n6047) );
  NAND2_X1 U5125 ( .A1(n4678), .A2(n4679), .ZN(n4677) );
  INV_X1 U5126 ( .A(n5753), .ZN(n4679) );
  MUX2_X1 U5127 ( .A(n6012), .B(n9112), .S(n7351), .Z(n6245) );
  INV_X1 U5128 ( .A(n4796), .ZN(n4795) );
  OAI21_X1 U5129 ( .B1(n7857), .B2(n4797), .A(n7984), .ZN(n4796) );
  INV_X1 U5130 ( .A(SI_8_), .ZN(n9780) );
  AOI21_X1 U5131 ( .B1(n8096), .B2(n4851), .A(n4518), .ZN(n4850) );
  INV_X1 U5132 ( .A(n7963), .ZN(n4851) );
  INV_X1 U5133 ( .A(n8096), .ZN(n4852) );
  INV_X1 U5134 ( .A(n5169), .ZN(n5657) );
  OR2_X1 U5135 ( .A1(n8755), .A2(n8548), .ZN(n5816) );
  NAND2_X1 U5136 ( .A1(n8778), .A2(n8368), .ZN(n5797) );
  OR2_X1 U5137 ( .A1(n8778), .A2(n8368), .ZN(n5801) );
  NAND2_X1 U5138 ( .A1(n8654), .A2(n5543), .ZN(n8605) );
  OR2_X1 U5139 ( .A1(n8816), .A2(n8701), .ZN(n8499) );
  AOI21_X1 U5140 ( .B1(n4941), .B2(n4944), .A(n4526), .ZN(n4940) );
  OR2_X1 U5141 ( .A1(n8111), .A2(n8110), .ZN(n5761) );
  OR2_X1 U5142 ( .A1(n8009), .A2(n8008), .ZN(n5853) );
  OAI21_X1 U5143 ( .B1(n5056), .B2(n4598), .A(n4534), .ZN(n4597) );
  INV_X1 U5144 ( .A(n8911), .ZN(n4598) );
  NOR2_X1 U5145 ( .A1(n9400), .A2(n9405), .ZN(n4766) );
  NAND2_X1 U5146 ( .A1(n9272), .A2(n9080), .ZN(n4813) );
  AND2_X1 U5147 ( .A1(n6382), .A2(n9286), .ZN(n9112) );
  NOR2_X1 U5148 ( .A1(n4820), .A2(n4819), .ZN(n4818) );
  INV_X1 U5149 ( .A(n4826), .ZN(n4819) );
  INV_X1 U5150 ( .A(n4824), .ZN(n4820) );
  NAND2_X1 U5151 ( .A1(n9944), .A2(n4758), .ZN(n4761) );
  INV_X1 U5152 ( .A(n7881), .ZN(n4758) );
  OR2_X1 U5153 ( .A1(n7881), .A2(n7890), .ZN(n7886) );
  INV_X1 U5154 ( .A(n4483), .ZN(n5917) );
  NAND2_X1 U5155 ( .A1(n7246), .A2(n9203), .ZN(n6539) );
  OAI21_X1 U5156 ( .B1(n5552), .B2(n4998), .A(n4997), .ZN(n5594) );
  AOI21_X1 U5157 ( .B1(n4999), .B2(n5550), .A(n4564), .ZN(n4997) );
  INV_X1 U5158 ( .A(n4999), .ZN(n4998) );
  AND2_X1 U5159 ( .A1(n4982), .A2(n5488), .ZN(n4981) );
  AND2_X1 U5160 ( .A1(n5509), .A2(n5494), .ZN(n5507) );
  AND2_X1 U5161 ( .A1(n5435), .A2(n5413), .ZN(n5433) );
  AOI21_X1 U5162 ( .B1(n5371), .B2(n5370), .A(n4574), .ZN(n5391) );
  INV_X1 U5163 ( .A(n5372), .ZN(n4574) );
  NAND2_X1 U5164 ( .A1(n5330), .A2(n9644), .ZN(n5369) );
  NOR2_X1 U5165 ( .A1(n5278), .A2(n4667), .ZN(n4666) );
  INV_X1 U5166 ( .A(n5261), .ZN(n4667) );
  INV_X1 U5167 ( .A(n5276), .ZN(n5278) );
  AND2_X1 U5168 ( .A1(n5295), .A2(n5282), .ZN(n5293) );
  NAND2_X1 U5169 ( .A1(n5263), .A2(n9780), .ZN(n5277) );
  NAND2_X1 U5170 ( .A1(n7650), .A2(n4861), .ZN(n4611) );
  AOI21_X1 U5171 ( .B1(n4861), .B2(n4863), .A(n4859), .ZN(n4858) );
  INV_X1 U5172 ( .A(n7906), .ZN(n4859) );
  AND2_X1 U5173 ( .A1(n5109), .A2(n8873), .ZN(n5134) );
  NOR2_X1 U5174 ( .A1(n8467), .A2(n8466), .ZN(n8469) );
  OR2_X1 U5175 ( .A1(n8773), .A2(n8572), .ZN(n5803) );
  NAND2_X1 U5176 ( .A1(n8608), .A2(n4955), .ZN(n8594) );
  NOR2_X1 U5177 ( .A1(n8597), .A2(n4688), .ZN(n4955) );
  AND2_X1 U5178 ( .A1(n5799), .A2(n5798), .ZN(n8614) );
  OR2_X1 U5179 ( .A1(n8666), .A2(n8503), .ZN(n5085) );
  OR2_X1 U5180 ( .A1(n8495), .A2(n8494), .ZN(n8496) );
  OR2_X1 U5181 ( .A1(n8832), .A2(n8370), .ZN(n5089) );
  AOI21_X1 U5182 ( .B1(n7597), .B2(n5042), .A(n4530), .ZN(n5041) );
  INV_X1 U5183 ( .A(n5693), .ZN(n5669) );
  INV_X1 U5184 ( .A(n5142), .ZN(n6825) );
  OAI21_X1 U5185 ( .B1(n5242), .B2(n4959), .A(n4958), .ZN(n7683) );
  AOI21_X1 U5186 ( .B1(n4962), .B2(n7589), .A(n4532), .ZN(n4958) );
  INV_X1 U5187 ( .A(n4962), .ZN(n4959) );
  NAND2_X1 U5188 ( .A1(n8381), .A2(n10308), .ZN(n10249) );
  INV_X1 U5189 ( .A(n8702), .ZN(n8639) );
  OR2_X1 U5190 ( .A1(n10277), .A2(n5870), .ZN(n10336) );
  OR2_X1 U5191 ( .A1(n9405), .A2(n9095), .ZN(n9124) );
  AND2_X1 U5192 ( .A1(n6359), .A2(n6375), .ZN(n6466) );
  AND2_X1 U5193 ( .A1(n9388), .A2(n9061), .ZN(n6464) );
  AND2_X1 U5194 ( .A1(n5961), .A2(n5960), .ZN(n9092) );
  OR2_X1 U5195 ( .A1(n9183), .A2(n6235), .ZN(n5961) );
  NAND2_X1 U5196 ( .A1(n4836), .A2(n4841), .ZN(n4832) );
  NAND2_X1 U5197 ( .A1(n4831), .A2(n4841), .ZN(n4830) );
  INV_X1 U5198 ( .A(n4834), .ZN(n4831) );
  AOI21_X1 U5199 ( .B1(n4836), .B2(n4835), .A(n4535), .ZN(n4834) );
  AND3_X1 U5200 ( .A1(n6279), .A2(n6278), .A3(n6277), .ZN(n9235) );
  INV_X1 U5201 ( .A(n4802), .ZN(n9241) );
  AOI21_X1 U5202 ( .B1(n9281), .B2(n4504), .A(n4803), .ZN(n4802) );
  NAND2_X1 U5203 ( .A1(n4804), .A2(n5086), .ZN(n4803) );
  INV_X1 U5204 ( .A(n6352), .ZN(n6246) );
  AOI21_X1 U5205 ( .B1(n4934), .B2(n4933), .A(n4932), .ZN(n4931) );
  INV_X1 U5206 ( .A(n7527), .ZN(n4933) );
  NAND2_X1 U5207 ( .A1(n7388), .A2(n7241), .ZN(n7310) );
  OR2_X1 U5208 ( .A1(n7386), .A2(n7393), .ZN(n7388) );
  NAND2_X1 U5209 ( .A1(n4966), .A2(n5235), .ZN(n5258) );
  AND2_X1 U5210 ( .A1(n5628), .A2(n5627), .ZN(n8573) );
  OR2_X1 U5211 ( .A1(n7172), .A2(n7171), .ZN(n4786) );
  AOI21_X1 U5212 ( .B1(n4655), .B2(n10254), .A(n4652), .ZN(n8758) );
  NAND2_X1 U5213 ( .A1(n4654), .A2(n4653), .ZN(n4652) );
  XNOR2_X1 U5214 ( .A(n8526), .B(n8530), .ZN(n4655) );
  NAND2_X1 U5215 ( .A1(n8528), .A2(n8702), .ZN(n4653) );
  AND2_X1 U5216 ( .A1(n5740), .A2(n7597), .ZN(n4578) );
  NAND2_X1 U5217 ( .A1(n4676), .A2(n4675), .ZN(n4674) );
  NOR2_X1 U5218 ( .A1(n8051), .A2(n5759), .ZN(n4668) );
  AOI21_X1 U5219 ( .B1(n5778), .B2(n8667), .A(n5777), .ZN(n4577) );
  NAND2_X1 U5220 ( .A1(n4688), .A2(n4687), .ZN(n4686) );
  NAND2_X1 U5221 ( .A1(n5802), .A2(n4692), .ZN(n4682) );
  OR2_X1 U5222 ( .A1(n8075), .A2(n8082), .ZN(n6389) );
  OR2_X1 U5223 ( .A1(n7887), .A2(n4916), .ZN(n4915) );
  NAND2_X1 U5224 ( .A1(n7846), .A2(n7848), .ZN(n4916) );
  NAND2_X1 U5225 ( .A1(n5668), .A2(n5667), .ZN(n5686) );
  INV_X1 U5226 ( .A(n4664), .ZN(n4663) );
  OAI21_X1 U5227 ( .B1(n4666), .B2(n4665), .A(n5293), .ZN(n4664) );
  INV_X1 U5228 ( .A(n5277), .ZN(n4665) );
  INV_X1 U5229 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n4969) );
  INV_X1 U5230 ( .A(n4697), .ZN(n4695) );
  INV_X1 U5231 ( .A(n4866), .ZN(n4627) );
  OAI21_X1 U5232 ( .B1(n8318), .B2(n8317), .A(n5083), .ZN(n8185) );
  AND2_X1 U5233 ( .A1(n8744), .A2(n8485), .ZN(n5832) );
  NOR2_X1 U5234 ( .A1(n8194), .A2(n8755), .ZN(n4733) );
  NAND2_X1 U5235 ( .A1(n5860), .A2(n5767), .ZN(n4648) );
  NAND2_X1 U5236 ( .A1(n5461), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5482) );
  INV_X1 U5237 ( .A(n5462), .ZN(n5461) );
  NOR2_X1 U5238 ( .A1(n8111), .A2(n8369), .ZN(n5033) );
  NOR2_X1 U5239 ( .A1(n8112), .A2(n5035), .ZN(n5034) );
  INV_X1 U5240 ( .A(n5089), .ZN(n5035) );
  INV_X1 U5241 ( .A(n5039), .ZN(n5036) );
  NAND3_X1 U5242 ( .A1(n5144), .A2(n5143), .A3(n5093), .ZN(n10283) );
  NOR2_X1 U5243 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(n4951), .ZN(n4950) );
  NAND2_X1 U5244 ( .A1(n5102), .A2(n4952), .ZN(n4951) );
  INV_X1 U5245 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n4952) );
  NAND2_X1 U5246 ( .A1(n4949), .A2(n4950), .ZN(n5700) );
  NAND2_X1 U5247 ( .A1(n6729), .A2(n6728), .ZN(n6730) );
  OR2_X1 U5248 ( .A1(n9094), .A2(n6727), .ZN(n6729) );
  INV_X1 U5249 ( .A(n6630), .ZN(n5080) );
  AND2_X1 U5250 ( .A1(n4716), .A2(n4550), .ZN(n4714) );
  NAND2_X1 U5251 ( .A1(n4979), .A2(n6376), .ZN(n4978) );
  NAND2_X1 U5252 ( .A1(n6295), .A2(n6450), .ZN(n4979) );
  NAND2_X1 U5253 ( .A1(n6365), .A2(n5002), .ZN(n5001) );
  INV_X1 U5254 ( .A(n6462), .ZN(n5002) );
  NOR2_X1 U5255 ( .A1(n10049), .A2(n4569), .ZN(n9027) );
  NOR2_X1 U5256 ( .A1(n9134), .A2(n6775), .ZN(n6404) );
  AND2_X1 U5257 ( .A1(n9134), .A2(n6775), .ZN(n6459) );
  NOR2_X1 U5258 ( .A1(n4898), .A2(n4892), .ZN(n4891) );
  INV_X1 U5259 ( .A(n4832), .ZN(n4829) );
  NAND2_X1 U5260 ( .A1(n9411), .A2(n9165), .ZN(n4841) );
  AND2_X1 U5261 ( .A1(n9094), .A2(n9165), .ZN(n9123) );
  OR2_X1 U5262 ( .A1(n9421), .A2(n9089), .ZN(n6450) );
  NOR2_X1 U5263 ( .A1(n9426), .A2(n9432), .ZN(n4757) );
  NOR2_X1 U5264 ( .A1(n9115), .A2(n4929), .ZN(n4928) );
  INV_X1 U5265 ( .A(n9113), .ZN(n4929) );
  OR2_X1 U5266 ( .A1(n9439), .A2(n9235), .ZN(n6378) );
  AND2_X1 U5267 ( .A1(n9442), .A2(n9082), .ZN(n9115) );
  OR2_X1 U5268 ( .A1(n9452), .A2(n9011), .ZN(n6382) );
  NOR2_X1 U5269 ( .A1(n9323), .A2(n9458), .ZN(n4748) );
  NAND2_X1 U5270 ( .A1(n9925), .A2(n9313), .ZN(n4826) );
  NOR2_X1 U5271 ( .A1(n9075), .A2(n4825), .ZN(n4824) );
  INV_X1 U5272 ( .A(n9071), .ZN(n4825) );
  OR2_X1 U5273 ( .A1(n9463), .A2(n6198), .ZN(n9104) );
  NOR2_X1 U5274 ( .A1(n8075), .A2(n4761), .ZN(n4760) );
  INV_X1 U5275 ( .A(n7864), .ZN(n4759) );
  NAND2_X1 U5276 ( .A1(n4794), .A2(n4793), .ZN(n7989) );
  AOI21_X1 U5277 ( .B1(n4795), .B2(n4797), .A(n4531), .ZN(n4793) );
  AND2_X1 U5278 ( .A1(n7696), .A2(n7543), .ZN(n4801) );
  NAND2_X1 U5279 ( .A1(n5647), .A2(n5646), .ZN(n5664) );
  NAND2_X1 U5280 ( .A1(n5531), .A2(n5529), .ZN(n5545) );
  AOI21_X1 U5281 ( .B1(n5469), .B2(n4986), .A(n4563), .ZN(n4985) );
  INV_X1 U5282 ( .A(n5452), .ZN(n4986) );
  NAND2_X1 U5283 ( .A1(n4989), .A2(n5435), .ZN(n4988) );
  NAND2_X1 U5284 ( .A1(n4991), .A2(n4993), .ZN(n4989) );
  INV_X1 U5285 ( .A(n4992), .ZN(n4991) );
  NOR2_X1 U5286 ( .A1(n5408), .A2(n4996), .ZN(n4995) );
  INV_X1 U5287 ( .A(n5389), .ZN(n4996) );
  NAND2_X1 U5288 ( .A1(n4994), .A2(n5407), .ZN(n4993) );
  NAND2_X1 U5289 ( .A1(n4995), .A2(n5390), .ZN(n4994) );
  NAND2_X1 U5290 ( .A1(n5369), .A2(n5332), .ZN(n5349) );
  NAND2_X1 U5291 ( .A1(n5327), .A2(SI_11_), .ZN(n5328) );
  INV_X1 U5292 ( .A(n5324), .ZN(n4975) );
  OAI21_X1 U5293 ( .B1(n4482), .B2(n4632), .A(n4631), .ZN(n4630) );
  NAND2_X1 U5294 ( .A1(n4482), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n4631) );
  INV_X1 U5295 ( .A(n4873), .ZN(n4872) );
  OAI21_X1 U5296 ( .B1(n7293), .B2(n4628), .A(n4500), .ZN(n7513) );
  AOI21_X1 U5297 ( .B1(n4878), .B2(n4880), .A(n8180), .ZN(n4877) );
  INV_X1 U5298 ( .A(n4884), .ZN(n4878) );
  INV_X1 U5299 ( .A(n8254), .ZN(n4875) );
  NAND2_X1 U5300 ( .A1(n7962), .A2(n4850), .ZN(n4616) );
  INV_X1 U5301 ( .A(n8163), .ZN(n4849) );
  OR2_X1 U5302 ( .A1(n8165), .A2(n8278), .ZN(n4614) );
  NOR2_X1 U5303 ( .A1(n4881), .A2(n8312), .ZN(n4880) );
  INV_X1 U5304 ( .A(n4882), .ZN(n4881) );
  INV_X1 U5305 ( .A(n4862), .ZN(n4861) );
  OAI21_X1 U5306 ( .B1(n4863), .B2(n4503), .A(n7753), .ZN(n4862) );
  OR2_X1 U5307 ( .A1(n7754), .A2(n4864), .ZN(n4863) );
  AND2_X1 U5308 ( .A1(n4509), .A2(n7028), .ZN(n4847) );
  OR2_X1 U5309 ( .A1(n4549), .A2(n10277), .ZN(n8168) );
  AND2_X1 U5310 ( .A1(n5573), .A2(n5572), .ZN(n8368) );
  AND4_X1 U5311 ( .A1(n5487), .A2(n5486), .A3(n5485), .A4(n5484), .ZN(n8502)
         );
  NOR2_X1 U5312 ( .A1(n7483), .A2(n4775), .ZN(n8403) );
  AND2_X1 U5313 ( .A1(n7484), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n4775) );
  NAND2_X1 U5314 ( .A1(n8403), .A2(n8404), .ZN(n8402) );
  OAI21_X1 U5315 ( .B1(n7486), .B2(n4770), .A(n4768), .ZN(n7727) );
  AOI21_X1 U5316 ( .B1(n4773), .B2(n4769), .A(n7671), .ZN(n4768) );
  INV_X1 U5317 ( .A(n4773), .ZN(n4770) );
  INV_X1 U5318 ( .A(n7487), .ZN(n4769) );
  NAND2_X1 U5319 ( .A1(n5825), .A2(n5826), .ZN(n8515) );
  OAI21_X1 U5320 ( .B1(n8567), .B2(n4965), .A(n4963), .ZN(n5645) );
  INV_X1 U5321 ( .A(n4964), .ZN(n4963) );
  OAI21_X1 U5322 ( .B1(n4510), .B2(n4965), .A(n5865), .ZN(n4964) );
  NAND2_X1 U5323 ( .A1(n8585), .A2(n8599), .ZN(n8582) );
  AND2_X1 U5324 ( .A1(n8597), .A2(n4501), .ZN(n5023) );
  OAI22_X1 U5325 ( .A1(n8627), .A2(n8633), .B1(n8656), .B2(n8789), .ZN(n8613)
         );
  OR2_X1 U5326 ( .A1(n8613), .A2(n8614), .ZN(n5024) );
  NAND2_X1 U5327 ( .A1(n8605), .A2(n5560), .ZN(n8608) );
  NAND2_X1 U5328 ( .A1(n5789), .A2(n5787), .ZN(n8669) );
  NAND2_X1 U5329 ( .A1(n8662), .A2(n8669), .ZN(n8661) );
  INV_X1 U5330 ( .A(n5772), .ZN(n4646) );
  INV_X1 U5331 ( .A(n4648), .ZN(n4645) );
  NAND2_X1 U5332 ( .A1(n5027), .A2(n5025), .ZN(n8691) );
  AOI21_X1 U5333 ( .B1(n5028), .B2(n8728), .A(n5026), .ZN(n5025) );
  INV_X1 U5334 ( .A(n8499), .ZN(n5026) );
  NAND2_X1 U5335 ( .A1(n5431), .A2(n8728), .ZN(n5432) );
  AND2_X1 U5336 ( .A1(n8712), .A2(n4551), .ZN(n5028) );
  NAND2_X1 U5337 ( .A1(n9911), .A2(n4727), .ZN(n4726) );
  NOR2_X1 U5338 ( .A1(n4728), .A2(n8495), .ZN(n4727) );
  AND2_X1 U5339 ( .A1(n5768), .A2(n5767), .ZN(n8728) );
  OR2_X1 U5340 ( .A1(n8727), .A2(n8728), .ZN(n5029) );
  INV_X1 U5341 ( .A(n5386), .ZN(n4944) );
  INV_X1 U5342 ( .A(n5761), .ZN(n4942) );
  AND2_X1 U5343 ( .A1(n5761), .A2(n5760), .ZN(n8112) );
  OR2_X1 U5344 ( .A1(n5038), .A2(n4489), .ZN(n8048) );
  AND4_X1 U5345 ( .A1(n5404), .A2(n5403), .A3(n5402), .A4(n5401), .ZN(n8281)
         );
  INV_X1 U5346 ( .A(n4637), .ZN(n4636) );
  OAI21_X1 U5347 ( .B1(n5305), .B2(n4638), .A(n5854), .ZN(n4637) );
  INV_X1 U5348 ( .A(n5749), .ZN(n4638) );
  AND2_X1 U5349 ( .A1(n5853), .A2(n5852), .ZN(n8010) );
  AND4_X1 U5350 ( .A1(n5346), .A2(n5345), .A3(n5344), .A4(n5343), .ZN(n8008)
         );
  OR2_X1 U5351 ( .A1(n7823), .A2(n7768), .ZN(n5749) );
  AND4_X1 U5352 ( .A1(n5323), .A2(n5322), .A3(n5321), .A4(n5320), .ZN(n7926)
         );
  NAND2_X1 U5353 ( .A1(n7810), .A2(n5305), .ZN(n7811) );
  AND2_X1 U5354 ( .A1(n7809), .A2(n5850), .ZN(n7762) );
  OR2_X1 U5355 ( .A1(n7594), .A2(n7597), .ZN(n7682) );
  AND2_X1 U5356 ( .A1(n5267), .A2(n4513), .ZN(n4657) );
  INV_X1 U5357 ( .A(n7444), .ZN(n5184) );
  CLKBUF_X1 U5358 ( .A(n7410), .Z(n7411) );
  NAND2_X1 U5359 ( .A1(n5604), .A2(n5603), .ZN(n8768) );
  NAND2_X1 U5360 ( .A1(n5480), .A2(n5479), .ZN(n8805) );
  NAND2_X1 U5361 ( .A1(n5460), .A2(n5459), .ZN(n8809) );
  AND3_X1 U5362 ( .A1(n5168), .A2(n5167), .A3(n5166), .ZN(n10302) );
  NOR2_X1 U5363 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_26__SCAN_IN), .ZN(
        n5091) );
  INV_X1 U5364 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5118) );
  INV_X1 U5365 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5046) );
  INV_X1 U5366 ( .A(n5476), .ZN(n4949) );
  XNOR2_X1 U5367 ( .A(n5673), .B(P2_IR_REG_21__SCAN_IN), .ZN(n6987) );
  INV_X1 U5368 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5101) );
  AND2_X1 U5369 ( .A1(n5163), .A2(n5164), .ZN(n5455) );
  INV_X1 U5370 ( .A(n7553), .ZN(n6588) );
  AOI21_X1 U5371 ( .B1(n5078), .B2(n8069), .A(n4717), .ZN(n4716) );
  XNOR2_X1 U5372 ( .A(n6713), .B(n6712), .ZN(n8889) );
  OR2_X1 U5373 ( .A1(n6147), .A2(n6133), .ZN(n6158) );
  NAND2_X1 U5374 ( .A1(n6763), .A2(n8956), .ZN(n6781) );
  NOR2_X1 U5375 ( .A1(n6781), .A2(n8879), .ZN(n4707) );
  NAND2_X1 U5376 ( .A1(n6676), .A2(n8978), .ZN(n8901) );
  NAND2_X1 U5377 ( .A1(n5939), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n6081) );
  INV_X1 U5378 ( .A(n6067), .ZN(n5939) );
  XNOR2_X1 U5379 ( .A(n6540), .B(n6712), .ZN(n6577) );
  OAI22_X1 U5380 ( .A1(n7539), .A2(n6727), .B1(n6538), .B2(n6733), .ZN(n6540)
         );
  OAI22_X1 U5381 ( .A1(n7539), .A2(n6755), .B1(n6538), .B2(n6727), .ZN(n6578)
         );
  OR2_X1 U5382 ( .A1(n6545), .A2(n6574), .ZN(n7205) );
  AND2_X1 U5383 ( .A1(n4600), .A2(n5048), .ZN(n4599) );
  AND2_X1 U5384 ( .A1(n5049), .A2(n6606), .ZN(n5048) );
  NAND2_X1 U5385 ( .A1(n8901), .A2(n8903), .ZN(n8900) );
  OR2_X1 U5386 ( .A1(n6160), .A2(n8070), .ZN(n6191) );
  OR2_X1 U5387 ( .A1(n4597), .A2(n4541), .ZN(n4594) );
  NAND2_X1 U5388 ( .A1(n7830), .A2(n7828), .ZN(n5047) );
  NAND2_X1 U5389 ( .A1(n4507), .A2(n6947), .ZN(n8140) );
  NAND2_X1 U5390 ( .A1(n4592), .A2(n4591), .ZN(n7553) );
  INV_X1 U5391 ( .A(n6582), .ZN(n4591) );
  INV_X1 U5392 ( .A(n6583), .ZN(n4592) );
  NAND2_X1 U5393 ( .A1(n5061), .A2(n5060), .ZN(n8989) );
  AOI21_X1 U5394 ( .B1(n4491), .B2(n5065), .A(n4565), .ZN(n5060) );
  AND2_X1 U5395 ( .A1(n6320), .A2(n6319), .ZN(n9095) );
  AND2_X1 U5396 ( .A1(n6305), .A2(n6304), .ZN(n9093) );
  OR2_X1 U5397 ( .A1(n9177), .A2(n6235), .ZN(n6305) );
  INV_X1 U5398 ( .A(n6034), .ZN(n6346) );
  OR2_X1 U5399 ( .A1(n6101), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n6113) );
  NOR2_X1 U5400 ( .A1(n10010), .A2(n4743), .ZN(n6909) );
  AND2_X1 U5401 ( .A1(n10015), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n4743) );
  OR2_X1 U5402 ( .A1(n6909), .A2(n6908), .ZN(n4742) );
  OR2_X1 U5403 ( .A1(n10086), .A2(n10085), .ZN(n4740) );
  NAND2_X1 U5404 ( .A1(n4740), .A2(n4739), .ZN(n4738) );
  NAND2_X1 U5405 ( .A1(n10089), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n4739) );
  AND2_X1 U5406 ( .A1(n4738), .A2(n4737), .ZN(n10096) );
  INV_X1 U5407 ( .A(n10097), .ZN(n4737) );
  AND2_X1 U5408 ( .A1(n6333), .A2(n6341), .ZN(n9145) );
  NOR2_X1 U5409 ( .A1(n9182), .A2(n9411), .ZN(n9175) );
  OR2_X1 U5410 ( .A1(n6298), .A2(n8992), .ZN(n6332) );
  AND2_X1 U5411 ( .A1(n4842), .A2(n4843), .ZN(n4838) );
  INV_X1 U5412 ( .A(n4839), .ZN(n4837) );
  AOI21_X1 U5413 ( .B1(n4505), .B2(n4843), .A(n4840), .ZN(n4839) );
  INV_X1 U5414 ( .A(n9188), .ZN(n4840) );
  NOR2_X1 U5415 ( .A1(n9123), .A2(n6455), .ZN(n9172) );
  NAND2_X1 U5416 ( .A1(n9195), .A2(n9119), .ZN(n9187) );
  NAND2_X1 U5417 ( .A1(n9090), .A2(n9089), .ZN(n4843) );
  NAND2_X1 U5418 ( .A1(n4920), .A2(n4918), .ZN(n9233) );
  NAND2_X1 U5419 ( .A1(n4919), .A2(n6416), .ZN(n4918) );
  INV_X1 U5420 ( .A(n4923), .ZN(n4919) );
  OR2_X1 U5421 ( .A1(n9256), .A2(n9439), .ZN(n9247) );
  NOR2_X1 U5422 ( .A1(n9247), .A2(n9432), .ZN(n9225) );
  INV_X1 U5423 ( .A(n9432), .ZN(n9226) );
  NOR2_X1 U5424 ( .A1(n4924), .A2(n9244), .ZN(n4923) );
  INV_X1 U5425 ( .A(n4927), .ZN(n4924) );
  AOI21_X1 U5426 ( .B1(n4928), .B2(n9273), .A(n6380), .ZN(n4927) );
  NAND2_X1 U5427 ( .A1(n9274), .A2(n4928), .ZN(n4925) );
  NAND2_X1 U5428 ( .A1(n6378), .A2(n6416), .ZN(n9244) );
  AND2_X1 U5429 ( .A1(n9288), .A2(n4813), .ZN(n4809) );
  NOR2_X1 U5430 ( .A1(n4808), .A2(n4811), .ZN(n4807) );
  NOR2_X1 U5431 ( .A1(n4814), .A2(n4519), .ZN(n4811) );
  INV_X1 U5432 ( .A(n4813), .ZN(n4808) );
  AND2_X1 U5433 ( .A1(n9452), .A2(n9275), .ZN(n4814) );
  OR2_X1 U5434 ( .A1(n9925), .A2(n8932), .ZN(n9310) );
  NOR2_X1 U5435 ( .A1(n9330), .A2(n4822), .ZN(n4821) );
  INV_X1 U5436 ( .A(n9074), .ZN(n4822) );
  NAND2_X1 U5437 ( .A1(n9072), .A2(n4824), .ZN(n4823) );
  AND2_X1 U5438 ( .A1(n9310), .A2(n9105), .ZN(n9330) );
  NOR2_X1 U5439 ( .A1(n9357), .A2(n4908), .ZN(n4907) );
  INV_X1 U5440 ( .A(n9103), .ZN(n4908) );
  NAND2_X1 U5441 ( .A1(n9102), .A2(n9101), .ZN(n4909) );
  OR2_X1 U5442 ( .A1(n9350), .A2(n9463), .ZN(n9348) );
  OR2_X1 U5443 ( .A1(n7786), .A2(n7853), .ZN(n7864) );
  AND2_X1 U5444 ( .A1(n7886), .A2(n7885), .ZN(n7860) );
  NAND2_X1 U5445 ( .A1(n7858), .A2(n7857), .ZN(n7883) );
  NAND2_X1 U5446 ( .A1(n5942), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n6145) );
  INV_X1 U5447 ( .A(n6108), .ZN(n5942) );
  NAND2_X1 U5448 ( .A1(n4801), .A2(n10179), .ZN(n7695) );
  OR2_X1 U5449 ( .A1(n10124), .A2(n6563), .ZN(n7390) );
  NAND2_X1 U5450 ( .A1(n5917), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4887) );
  AND2_X1 U5451 ( .A1(n8151), .A2(n6790), .ZN(n9370) );
  NAND2_X1 U5452 ( .A1(n6329), .A2(n6328), .ZN(n9400) );
  NAND2_X1 U5453 ( .A1(n5938), .A2(n5937), .ZN(n9416) );
  NAND2_X1 U5454 ( .A1(n5630), .A2(n5629), .ZN(n5632) );
  XNOR2_X1 U5455 ( .A(n5936), .B(P1_IR_REG_22__SCAN_IN), .ZN(n7246) );
  NAND2_X1 U5456 ( .A1(n5510), .A2(n5509), .ZN(n5520) );
  OAI21_X1 U5457 ( .B1(n5391), .B2(n5390), .A(n5389), .ZN(n5409) );
  NAND2_X1 U5458 ( .A1(n4662), .A2(n5277), .ZN(n5294) );
  NAND2_X1 U5459 ( .A1(n5262), .A2(n4666), .ZN(n4662) );
  XNOR2_X1 U5460 ( .A(n5259), .B(SI_7_), .ZN(n5257) );
  NAND2_X1 U5461 ( .A1(n5217), .A2(n4582), .ZN(n5219) );
  INV_X1 U5462 ( .A(n5218), .ZN(n4582) );
  XNOR2_X1 U5463 ( .A(n5234), .B(n5221), .ZN(n5232) );
  XNOR2_X1 U5464 ( .A(n5197), .B(n5181), .ZN(n5195) );
  INV_X1 U5465 ( .A(SI_4_), .ZN(n5181) );
  OAI21_X1 U5466 ( .B1(n4483), .B2(n4580), .A(n4579), .ZN(n5139) );
  NAND2_X1 U5467 ( .A1(n4483), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4579) );
  XNOR2_X1 U5468 ( .A(n5128), .B(n5127), .ZN(n5140) );
  OAI21_X1 U5469 ( .B1(n8329), .B2(n8173), .A(n8328), .ZN(n8330) );
  NAND2_X1 U5470 ( .A1(n4500), .A2(n4628), .ZN(n4625) );
  AND4_X1 U5471 ( .A1(n5504), .A2(n5503), .A3(n5502), .A4(n5501), .ZN(n8503)
         );
  NAND2_X1 U5472 ( .A1(n5423), .A2(n5422), .ZN(n8820) );
  NAND2_X1 U5473 ( .A1(n7293), .A2(n7292), .ZN(n7345) );
  NOR2_X1 U5474 ( .A1(n8293), .A2(n8292), .ZN(n8329) );
  INV_X1 U5475 ( .A(n8670), .ZN(n8638) );
  INV_X1 U5476 ( .A(n8632), .ZN(n8789) );
  NAND2_X1 U5477 ( .A1(n5315), .A2(n5314), .ZN(n8840) );
  AND4_X1 U5478 ( .A1(n5367), .A2(n5366), .A3(n5365), .A4(n5364), .ZN(n8370)
         );
  AND2_X1 U5479 ( .A1(n7130), .A2(n4787), .ZN(n7172) );
  NAND2_X1 U5480 ( .A1(n7081), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n4787) );
  AND2_X1 U5481 ( .A1(n4786), .A2(n4785), .ZN(n7184) );
  NAND2_X1 U5482 ( .A1(n7083), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n4785) );
  XNOR2_X1 U5483 ( .A(n8465), .B(n8472), .ZN(n8450) );
  NAND2_X1 U5484 ( .A1(n8475), .A2(n8474), .ZN(n4782) );
  OAI22_X1 U5485 ( .A1(n8477), .A2(n10237), .B1(n8476), .B2(n10236), .ZN(n4779) );
  AOI21_X1 U5486 ( .B1(n8570), .B2(n8569), .A(n8568), .ZN(n8571) );
  NAND2_X1 U5487 ( .A1(n4633), .A2(n5803), .ZN(n8569) );
  OR2_X1 U5488 ( .A1(n8620), .A2(n9847), .ZN(n4855) );
  NAND2_X1 U5489 ( .A1(n4656), .A2(n8758), .ZN(n8845) );
  AND2_X1 U5490 ( .A1(n8759), .A2(n8757), .ZN(n4656) );
  NAND2_X1 U5491 ( .A1(n5104), .A2(n4956), .ZN(n8868) );
  AND2_X1 U5492 ( .A1(n4493), .A2(n4957), .ZN(n4956) );
  INV_X1 U5493 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n4957) );
  NAND2_X1 U5494 ( .A1(n7792), .A2(n6607), .ZN(n7830) );
  NAND2_X1 U5495 ( .A1(n6131), .A2(n6130), .ZN(n7881) );
  NAND2_X1 U5496 ( .A1(n4709), .A2(n4708), .ZN(n6764) );
  INV_X1 U5497 ( .A(n8881), .ZN(n4709) );
  AND4_X1 U5498 ( .A1(n6087), .A2(n6086), .A3(n6085), .A4(n6084), .ZN(n7544)
         );
  OAI211_X1 U5499 ( .C1(n6117), .C2(n6883), .A(n6076), .B(n6075), .ZN(n10176)
         );
  OR2_X1 U5500 ( .A1(n6034), .A2(n6033), .ZN(n6040) );
  NAND4_X2 U5501 ( .A1(n6025), .A2(n4499), .A3(n6024), .A4(n6026), .ZN(n6027)
         );
  OR2_X1 U5502 ( .A1(n6035), .A2(n6833), .ZN(n6025) );
  NAND2_X1 U5503 ( .A1(n4767), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5916) );
  INV_X1 U5504 ( .A(n5912), .ZN(n4885) );
  OR2_X1 U5505 ( .A1(n10002), .A2(n4546), .ZN(n6961) );
  NAND2_X1 U5506 ( .A1(n10103), .A2(n10104), .ZN(n10102) );
  AND2_X1 U5507 ( .A1(n5920), .A2(n5919), .ZN(n9388) );
  OR2_X1 U5508 ( .A1(n5910), .A2(n5913), .ZN(n4724) );
  AND2_X1 U5509 ( .A1(n5734), .A2(n4692), .ZN(n4586) );
  NAND2_X1 U5510 ( .A1(n4691), .A2(n4690), .ZN(n5747) );
  INV_X1 U5511 ( .A(n5852), .ZN(n4672) );
  NAND2_X1 U5512 ( .A1(n4677), .A2(n4515), .ZN(n4676) );
  AND2_X1 U5513 ( .A1(n4669), .A2(n4668), .ZN(n5766) );
  AND2_X1 U5514 ( .A1(n5788), .A2(n5781), .ZN(n4576) );
  NAND2_X1 U5515 ( .A1(n6494), .A2(n7351), .ZN(n4976) );
  AOI21_X1 U5516 ( .B1(n4978), .B2(n6366), .A(n4492), .ZN(n4977) );
  INV_X1 U5517 ( .A(n5800), .ZN(n4683) );
  NAND2_X1 U5518 ( .A1(n4682), .A2(n4681), .ZN(n4680) );
  INV_X1 U5519 ( .A(n5085), .ZN(n5019) );
  INV_X1 U5520 ( .A(n4606), .ZN(n4605) );
  NAND2_X1 U5521 ( .A1(n6349), .A2(n9394), .ZN(n5007) );
  NAND2_X1 U5522 ( .A1(n9120), .A2(n6450), .ZN(n6494) );
  INV_X1 U5523 ( .A(n7882), .ZN(n4797) );
  NOR2_X1 U5524 ( .A1(n5575), .A2(n5000), .ZN(n4999) );
  INV_X1 U5525 ( .A(n5561), .ZN(n5000) );
  INV_X1 U5526 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5901) );
  INV_X1 U5527 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5902) );
  INV_X1 U5528 ( .A(n5489), .ZN(n4984) );
  AND2_X1 U5529 ( .A1(n4985), .A2(n4984), .ZN(n4983) );
  OAI21_X1 U5530 ( .B1(n4993), .B2(n4995), .A(n5433), .ZN(n4992) );
  NAND2_X1 U5531 ( .A1(n5296), .A2(n9795), .ZN(n5308) );
  AOI21_X1 U5532 ( .B1(n4585), .B2(n4516), .A(n4495), .ZN(n5833) );
  NAND2_X1 U5533 ( .A1(n5830), .A2(n5829), .ZN(n4585) );
  INV_X1 U5534 ( .A(n5109), .ZN(n5111) );
  AND2_X1 U5535 ( .A1(n8748), .A2(n4733), .ZN(n4732) );
  OR2_X1 U5536 ( .A1(n8483), .A2(n8248), .ZN(n5825) );
  INV_X1 U5537 ( .A(n5814), .ZN(n4965) );
  OR2_X1 U5538 ( .A1(n8768), .A2(n8508), .ZN(n5807) );
  AND2_X1 U5539 ( .A1(n8618), .A2(n4722), .ZN(n4721) );
  NOR2_X1 U5540 ( .A1(n8789), .A2(n8794), .ZN(n4722) );
  INV_X1 U5541 ( .A(n5018), .ZN(n5017) );
  OAI21_X1 U5542 ( .B1(n8669), .B2(n5019), .A(n8504), .ZN(n5018) );
  OR2_X1 U5543 ( .A1(n8794), .A2(n8670), .ZN(n8504) );
  NAND2_X1 U5544 ( .A1(n5017), .A2(n5019), .ZN(n5016) );
  NAND2_X1 U5545 ( .A1(n5776), .A2(n4643), .ZN(n4642) );
  NAND2_X1 U5546 ( .A1(n5785), .A2(n4646), .ZN(n4643) );
  OR2_X1 U5547 ( .A1(n8805), .A2(n8502), .ZN(n5783) );
  OR2_X1 U5548 ( .A1(n8820), .A2(n8289), .ZN(n5768) );
  OR2_X1 U5549 ( .A1(n5399), .A2(n8358), .ZN(n5425) );
  NAND2_X1 U5550 ( .A1(n8832), .A2(n4729), .ZN(n4728) );
  NAND2_X1 U5551 ( .A1(n5360), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5380) );
  INV_X1 U5552 ( .A(n5362), .ZN(n5360) );
  NAND2_X1 U5553 ( .A1(n4636), .A2(n4638), .ZN(n4635) );
  NAND2_X1 U5554 ( .A1(n5316), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5341) );
  INV_X1 U5555 ( .A(n5318), .ZN(n5316) );
  OR2_X1 U5556 ( .A1(n5341), .A2(n9821), .ZN(n5362) );
  NAND2_X1 U5557 ( .A1(n5286), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5318) );
  INV_X1 U5558 ( .A(n5287), .ZN(n5286) );
  NOR2_X1 U5559 ( .A1(n7762), .A2(n5043), .ZN(n5042) );
  INV_X1 U5560 ( .A(n7681), .ZN(n5043) );
  OR2_X1 U5561 ( .A1(n5269), .A2(n5268), .ZN(n5287) );
  AND2_X1 U5562 ( .A1(n7597), .A2(n5243), .ZN(n4962) );
  NAND2_X1 U5563 ( .A1(n5202), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5226) );
  INV_X1 U5564 ( .A(n5203), .ZN(n5202) );
  AND2_X1 U5565 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5186) );
  NAND2_X1 U5566 ( .A1(n5186), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5203) );
  NOR2_X1 U5567 ( .A1(n10245), .A2(n7380), .ZN(n4700) );
  AND2_X1 U5568 ( .A1(n7444), .A2(n7371), .ZN(n5011) );
  INV_X1 U5569 ( .A(n7373), .ZN(n5012) );
  OR2_X1 U5570 ( .A1(n5641), .A2(n7228), .ZN(n5135) );
  XNOR2_X1 U5571 ( .A(n6543), .B(n6712), .ZN(n6575) );
  NAND2_X1 U5572 ( .A1(n5053), .A2(n5052), .ZN(n5049) );
  INV_X1 U5573 ( .A(n4604), .ZN(n4603) );
  OAI21_X1 U5574 ( .B1(n4607), .B2(n4605), .A(n5052), .ZN(n4604) );
  NAND2_X1 U5575 ( .A1(n4603), .A2(n4605), .ZN(n4600) );
  NAND2_X1 U5576 ( .A1(n8977), .A2(n8979), .ZN(n6676) );
  INV_X1 U5577 ( .A(n4597), .ZN(n4595) );
  INV_X1 U5578 ( .A(n8921), .ZN(n5062) );
  INV_X1 U5579 ( .A(n5077), .ZN(n5076) );
  OAI21_X1 U5580 ( .B1(n5078), .B2(n4717), .A(n6658), .ZN(n5077) );
  NAND2_X1 U5581 ( .A1(n5081), .A2(n5075), .ZN(n5074) );
  OR2_X1 U5582 ( .A1(n9064), .A2(n6401), .ZN(n6523) );
  OR2_X1 U5583 ( .A1(n9978), .A2(n6875), .ZN(n9980) );
  NOR2_X1 U5584 ( .A1(n10065), .A2(n9028), .ZN(n9030) );
  OR2_X1 U5585 ( .A1(n9400), .A2(n9096), .ZN(n6403) );
  INV_X1 U5586 ( .A(n4838), .ZN(n4835) );
  NAND2_X1 U5587 ( .A1(n4757), .A2(n9090), .ZN(n4756) );
  NOR2_X1 U5588 ( .A1(n9116), .A2(n4922), .ZN(n4921) );
  INV_X1 U5589 ( .A(n4928), .ZN(n4922) );
  NAND2_X1 U5590 ( .A1(n4504), .A2(n4807), .ZN(n4804) );
  AND2_X1 U5591 ( .A1(n6389), .A2(n7993), .ZN(n8032) );
  AOI21_X1 U5592 ( .B1(n4913), .B2(n4912), .A(n6201), .ZN(n4911) );
  INV_X1 U5593 ( .A(n4917), .ZN(n4912) );
  NOR2_X1 U5594 ( .A1(n7887), .A2(n6390), .ZN(n4917) );
  INV_X1 U5595 ( .A(n7545), .ZN(n4800) );
  AND2_X1 U5596 ( .A1(n6027), .A2(n7238), .ZN(n10128) );
  AND2_X1 U5597 ( .A1(n7698), .A2(n10192), .ZN(n7630) );
  XNOR2_X1 U5598 ( .A(n5686), .B(n5685), .ZN(n5683) );
  INV_X1 U5599 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5921) );
  NAND2_X1 U5600 ( .A1(n5595), .A2(n5601), .ZN(n5617) );
  INV_X1 U5601 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n6468) );
  INV_X1 U5602 ( .A(n5387), .ZN(n5390) );
  AOI21_X1 U5603 ( .B1(n4663), .B2(n4665), .A(n4661), .ZN(n4660) );
  INV_X1 U5604 ( .A(n5295), .ZN(n4661) );
  INV_X1 U5605 ( .A(SI_5_), .ZN(n9680) );
  NAND2_X1 U5606 ( .A1(n4630), .A2(SI_3_), .ZN(n5176) );
  OAI21_X1 U5607 ( .B1(n4483), .B2(n4584), .A(n4583), .ZN(n5158) );
  NAND2_X1 U5608 ( .A1(n4482), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n4583) );
  NAND2_X1 U5609 ( .A1(n4695), .A2(n4967), .ZN(n4694) );
  NOR2_X1 U5610 ( .A1(n4969), .A2(n4968), .ZN(n4967) );
  NAND2_X1 U5611 ( .A1(n9889), .A2(n5125), .ZN(n4698) );
  INV_X1 U5612 ( .A(P1_RD_REG_SCAN_IN), .ZN(n5125) );
  NAND2_X1 U5613 ( .A1(n9888), .A2(n5126), .ZN(n4697) );
  AND2_X1 U5614 ( .A1(n8241), .A2(n8199), .ZN(n8204) );
  INV_X1 U5615 ( .A(n7738), .ZN(n4865) );
  AND2_X1 U5616 ( .A1(n8233), .A2(n8175), .ZN(n4884) );
  INV_X1 U5617 ( .A(n7299), .ZN(n4628) );
  AND2_X1 U5618 ( .A1(n7502), .A2(n7496), .ZN(n4868) );
  NAND2_X1 U5619 ( .A1(n4627), .A2(n7299), .ZN(n4624) );
  NAND2_X1 U5620 ( .A1(n5224), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5244) );
  INV_X1 U5621 ( .A(n5226), .ZN(n5224) );
  OR2_X1 U5622 ( .A1(n5244), .A2(n7518), .ZN(n5269) );
  NAND2_X1 U5623 ( .A1(n4623), .A2(n4622), .ZN(n4621) );
  INV_X1 U5624 ( .A(n8212), .ZN(n4622) );
  NAND2_X1 U5625 ( .A1(n8299), .A2(n8368), .ZN(n4623) );
  INV_X1 U5626 ( .A(n6990), .ZN(n4846) );
  INV_X1 U5627 ( .A(n6991), .ZN(n4844) );
  INV_X1 U5628 ( .A(n5499), .ZN(n5497) );
  NAND2_X1 U5629 ( .A1(n8174), .A2(n4883), .ZN(n4882) );
  INV_X1 U5630 ( .A(n8176), .ZN(n4883) );
  AND2_X1 U5631 ( .A1(n8383), .A2(n8168), .ZN(n7030) );
  NOR2_X1 U5632 ( .A1(n7344), .A2(n4867), .ZN(n4866) );
  INV_X1 U5633 ( .A(n7292), .ZN(n4867) );
  OR2_X1 U5634 ( .A1(n8191), .A2(n8192), .ZN(n4873) );
  NAND2_X1 U5635 ( .A1(n4618), .A2(n4617), .ZN(n8266) );
  INV_X1 U5636 ( .A(n4620), .ZN(n4617) );
  NOR2_X1 U5637 ( .A1(n8189), .A2(n4619), .ZN(n4618) );
  INV_X1 U5638 ( .A(n8267), .ZN(n4619) );
  AND2_X1 U5639 ( .A1(n8266), .A2(n4561), .ZN(n8339) );
  OAI21_X1 U5640 ( .B1(n7962), .B2(n4852), .A(n4850), .ZN(n8275) );
  INV_X1 U5641 ( .A(n5644), .ZN(n5609) );
  AND4_X1 U5642 ( .A1(n5385), .A2(n5384), .A3(n5383), .A4(n5382), .ZN(n8110)
         );
  AND4_X1 U5643 ( .A1(n5173), .A2(n5172), .A3(n5171), .A4(n5170), .ZN(n7414)
         );
  AND2_X1 U5644 ( .A1(n5109), .A2(n5110), .ZN(n5169) );
  AND2_X1 U5645 ( .A1(n7102), .A2(n4789), .ZN(n9894) );
  NAND2_X1 U5646 ( .A1(n7080), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n4789) );
  NOR2_X1 U5647 ( .A1(n9894), .A2(n4788), .ZN(n9893) );
  NOR2_X1 U5648 ( .A1(n8386), .A2(n4776), .ZN(n7278) );
  AND2_X1 U5649 ( .A1(n8391), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n4776) );
  NOR2_X1 U5650 ( .A1(n7278), .A2(n7277), .ZN(n7483) );
  AND2_X1 U5651 ( .A1(n7676), .A2(n7673), .ZN(n4773) );
  NOR2_X1 U5652 ( .A1(n8447), .A2(n4572), .ZN(n8465) );
  AND2_X1 U5653 ( .A1(n8560), .A2(n4730), .ZN(n8489) );
  NOR2_X1 U5654 ( .A1(n4731), .A2(n8490), .ZN(n4730) );
  INV_X1 U5655 ( .A(n4732), .ZN(n4731) );
  AND2_X1 U5656 ( .A1(n5638), .A2(n5654), .ZN(n8533) );
  NAND2_X1 U5657 ( .A1(n8542), .A2(n5814), .ZN(n8526) );
  NAND2_X1 U5658 ( .A1(n8527), .A2(n8700), .ZN(n4654) );
  INV_X1 U5659 ( .A(n8540), .ZN(n8543) );
  NAND2_X1 U5660 ( .A1(n8768), .A2(n8508), .ZN(n5808) );
  XNOR2_X1 U5661 ( .A(n8194), .B(n8573), .ZN(n8540) );
  NAND2_X1 U5662 ( .A1(n4633), .A2(n4524), .ZN(n8567) );
  NAND2_X1 U5663 ( .A1(n8576), .A2(n4681), .ZN(n4633) );
  NAND2_X1 U5664 ( .A1(n5807), .A2(n5808), .ZN(n8570) );
  NAND2_X1 U5665 ( .A1(n5584), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n5607) );
  NAND2_X1 U5666 ( .A1(n5022), .A2(n5021), .ZN(n8581) );
  AOI21_X1 U5667 ( .B1(n5023), .B2(n8614), .A(n4533), .ZN(n5021) );
  NAND2_X1 U5668 ( .A1(n8594), .A2(n5801), .ZN(n8576) );
  AND2_X1 U5669 ( .A1(n8663), .A2(n4719), .ZN(n8599) );
  AND2_X1 U5670 ( .A1(n4721), .A2(n4720), .ZN(n4719) );
  NAND2_X1 U5671 ( .A1(n8663), .A2(n4721), .ZN(n8616) );
  AND2_X1 U5672 ( .A1(n5781), .A2(n5794), .ZN(n8633) );
  AOI21_X1 U5673 ( .B1(n8683), .B2(n5506), .A(n5777), .ZN(n8655) );
  NAND2_X1 U5674 ( .A1(n8655), .A2(n5519), .ZN(n8654) );
  NAND2_X1 U5675 ( .A1(n8663), .A2(n8652), .ZN(n8647) );
  NAND2_X1 U5676 ( .A1(n5432), .A2(n4647), .ZN(n4641) );
  NOR2_X1 U5677 ( .A1(n4648), .A2(n5840), .ZN(n4647) );
  INV_X1 U5678 ( .A(n4642), .ZN(n4639) );
  NAND2_X1 U5679 ( .A1(n4641), .A2(n4640), .ZN(n8683) );
  NOR2_X1 U5680 ( .A1(n8676), .A2(n4642), .ZN(n4640) );
  OR2_X1 U5681 ( .A1(n8692), .A2(n8805), .ZN(n8678) );
  AOI22_X1 U5682 ( .A1(n8691), .A2(n8501), .B1(n8500), .B2(n8697), .ZN(n8677)
         );
  AND2_X1 U5683 ( .A1(n8730), .A2(n8723), .ZN(n8717) );
  NAND2_X1 U5684 ( .A1(n5424), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5442) );
  INV_X1 U5685 ( .A(n5425), .ZN(n5424) );
  OR2_X1 U5686 ( .A1(n5442), .A2(n5441), .ZN(n5462) );
  INV_X1 U5687 ( .A(n8728), .ZN(n8735) );
  NOR2_X1 U5688 ( .A1(n4488), .A2(n8820), .ZN(n8730) );
  NAND2_X1 U5689 ( .A1(n5034), .A2(n5031), .ZN(n5030) );
  AOI21_X1 U5690 ( .B1(n5034), .B2(n4489), .A(n5033), .ZN(n5032) );
  INV_X1 U5691 ( .A(n8010), .ZN(n5031) );
  NOR2_X1 U5692 ( .A1(n7927), .A2(n4728), .ZN(n8054) );
  NAND2_X1 U5693 ( .A1(n8014), .A2(n8015), .ZN(n8050) );
  NOR2_X1 U5694 ( .A1(n7927), .A2(n8009), .ZN(n8021) );
  OR2_X1 U5695 ( .A1(n7820), .A2(n8840), .ZN(n7927) );
  NAND2_X1 U5696 ( .A1(n7806), .A2(n7764), .ZN(n7921) );
  AND2_X1 U5697 ( .A1(n5748), .A2(n5749), .ZN(n7812) );
  NAND2_X1 U5698 ( .A1(n4699), .A2(n10321), .ZN(n7685) );
  NOR2_X1 U5699 ( .A1(n4961), .A2(n4960), .ZN(n7598) );
  INV_X1 U5700 ( .A(n5243), .ZN(n4960) );
  INV_X1 U5701 ( .A(n7461), .ZN(n4961) );
  NAND2_X1 U5702 ( .A1(n7461), .A2(n4962), .ZN(n7596) );
  AND4_X1 U5703 ( .A1(n5208), .A2(n5207), .A3(n5206), .A4(n5205), .ZN(n7458)
         );
  AOI21_X1 U5704 ( .B1(n5846), .B2(n5713), .A(n5714), .ZN(n4947) );
  NAND2_X1 U5705 ( .A1(n5242), .A2(n5241), .ZN(n7461) );
  OAI21_X1 U5706 ( .B1(n10243), .B2(n7375), .A(n7374), .ZN(n7456) );
  AND2_X1 U5707 ( .A1(n4700), .A2(n7382), .ZN(n7463) );
  INV_X1 U5708 ( .A(n4700), .ZN(n10248) );
  OAI21_X1 U5709 ( .B1(n7332), .B2(n7367), .A(n5721), .ZN(n7412) );
  NAND2_X1 U5710 ( .A1(n7034), .A2(n4853), .ZN(n7416) );
  NAND2_X1 U5711 ( .A1(n5583), .A2(n5582), .ZN(n8773) );
  NAND2_X1 U5712 ( .A1(n5496), .A2(n5495), .ZN(n8799) );
  INV_X1 U5713 ( .A(n7823), .ZN(n10328) );
  AND2_X1 U5714 ( .A1(n6995), .A2(n6993), .ZN(n10267) );
  OR2_X1 U5715 ( .A1(n6249), .A2(n8906), .ZN(n6260) );
  INV_X1 U5716 ( .A(n6759), .ZN(n6733) );
  NAND2_X1 U5717 ( .A1(n7565), .A2(n7566), .ZN(n4606) );
  OR2_X1 U5718 ( .A1(n7565), .A2(n7566), .ZN(n4607) );
  AND2_X1 U5719 ( .A1(n5057), .A2(n6693), .ZN(n5056) );
  NAND2_X1 U5720 ( .A1(n8955), .A2(n5058), .ZN(n5057) );
  NOR2_X1 U5721 ( .A1(n5059), .A2(n5055), .ZN(n5054) );
  INV_X1 U5722 ( .A(n8903), .ZN(n5055) );
  INV_X1 U5723 ( .A(n8955), .ZN(n5059) );
  NAND2_X1 U5724 ( .A1(n5949), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n6274) );
  INV_X1 U5725 ( .A(n6260), .ZN(n5949) );
  NAND2_X1 U5726 ( .A1(n5944), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n6160) );
  INV_X1 U5727 ( .A(n6158), .ZN(n5944) );
  OR2_X1 U5728 ( .A1(n5067), .A2(n5088), .ZN(n5064) );
  AND2_X1 U5729 ( .A1(n8947), .A2(n5068), .ZN(n5067) );
  NAND2_X1 U5730 ( .A1(n6716), .A2(n6715), .ZN(n5068) );
  NAND2_X1 U5731 ( .A1(n5069), .A2(n6715), .ZN(n5065) );
  XNOR2_X1 U5732 ( .A(n6723), .B(n7546), .ZN(n6725) );
  OAI22_X1 U5733 ( .A1(n9186), .A2(n6727), .B1(n9092), .B2(n6755), .ZN(n6724)
         );
  NAND2_X1 U5734 ( .A1(n8937), .A2(n8939), .ZN(n8938) );
  OR2_X1 U5735 ( .A1(n7636), .A2(n7637), .ZN(n5052) );
  AND2_X1 U5736 ( .A1(n7636), .A2(n7637), .ZN(n5053) );
  NAND2_X1 U5737 ( .A1(n6608), .A2(n6027), .ZN(n6548) );
  AND2_X1 U5738 ( .A1(n6551), .A2(n6550), .ZN(n6949) );
  NAND2_X1 U5739 ( .A1(n5945), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n6193) );
  INV_X1 U5740 ( .A(n6191), .ZN(n5945) );
  INV_X1 U5741 ( .A(n8068), .ZN(n4718) );
  NAND2_X1 U5742 ( .A1(n5947), .A2(n5946), .ZN(n6007) );
  INV_X1 U5743 ( .A(n6234), .ZN(n5947) );
  NAND2_X1 U5744 ( .A1(n5948), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n6249) );
  INV_X1 U5745 ( .A(n6007), .ZN(n5948) );
  INV_X1 U5746 ( .A(n8989), .ZN(n4609) );
  AOI21_X1 U5747 ( .B1(n4714), .B2(n5079), .A(n4537), .ZN(n4712) );
  INV_X1 U5748 ( .A(n4714), .ZN(n4713) );
  INV_X1 U5749 ( .A(n6565), .ZN(n6755) );
  INV_X1 U5750 ( .A(n4978), .ZN(n6452) );
  AND2_X1 U5751 ( .A1(n6461), .A2(n6460), .ZN(n6522) );
  AND2_X1 U5752 ( .A1(n6367), .A2(n6366), .ZN(n6368) );
  AND4_X1 U5753 ( .A1(n6239), .A2(n6238), .A3(n6237), .A4(n6236), .ZN(n9012)
         );
  AND4_X1 U5754 ( .A1(n6225), .A2(n6224), .A3(n6223), .A4(n6222), .ZN(n8932)
         );
  AND4_X1 U5755 ( .A1(n6112), .A2(n6111), .A3(n6110), .A4(n6109), .ZN(n7557)
         );
  OR2_X1 U5756 ( .A1(n4485), .A2(n6013), .ZN(n6017) );
  OR2_X1 U5757 ( .A1(n6034), .A2(n6839), .ZN(n6026) );
  OR2_X1 U5758 ( .A1(n6929), .A2(n6928), .ZN(n6926) );
  OR2_X1 U5759 ( .A1(n6113), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n6102) );
  NAND2_X1 U5760 ( .A1(n9025), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4741) );
  NAND2_X1 U5761 ( .A1(n4511), .A2(n10028), .ZN(n10027) );
  XNOR2_X1 U5762 ( .A(n9027), .B(n9040), .ZN(n10066) );
  NOR2_X1 U5763 ( .A1(n10066), .A2(n6178), .ZN(n10065) );
  NOR2_X1 U5764 ( .A1(n10096), .A2(n4736), .ZN(n10112) );
  AND2_X1 U5765 ( .A1(n10101), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n4736) );
  NOR2_X1 U5766 ( .A1(n6404), .A2(n6459), .ZN(n9099) );
  NAND2_X1 U5767 ( .A1(n9400), .A2(n9096), .ZN(n9126) );
  AOI21_X1 U5768 ( .B1(n4897), .B2(n4896), .A(n4895), .ZN(n4894) );
  INV_X1 U5769 ( .A(n9124), .ZN(n4895) );
  NAND2_X1 U5770 ( .A1(n6403), .A2(n9126), .ZN(n9148) );
  AOI21_X1 U5771 ( .B1(n4827), .B2(n4517), .A(n4828), .ZN(n9142) );
  INV_X1 U5772 ( .A(n4901), .ZN(n4900) );
  OAI21_X1 U5773 ( .B1(n9123), .B2(n4902), .A(n9122), .ZN(n4901) );
  NAND2_X1 U5774 ( .A1(n9121), .A2(n9120), .ZN(n4902) );
  NAND2_X1 U5775 ( .A1(n4903), .A2(n4892), .ZN(n4893) );
  NAND2_X1 U5776 ( .A1(n5952), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n6298) );
  OR2_X1 U5777 ( .A1(n6285), .A2(n8896), .ZN(n5977) );
  NAND2_X1 U5778 ( .A1(n5951), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n5967) );
  INV_X1 U5779 ( .A(n5977), .ZN(n5951) );
  NOR2_X1 U5780 ( .A1(n9247), .A2(n4755), .ZN(n9219) );
  INV_X1 U5781 ( .A(n4757), .ZN(n4755) );
  OR2_X1 U5782 ( .A1(n6274), .A2(n8914), .ZN(n6283) );
  NAND2_X1 U5783 ( .A1(n5950), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n6285) );
  INV_X1 U5784 ( .A(n6283), .ZN(n5950) );
  AND2_X1 U5785 ( .A1(n9338), .A2(n4555), .ZN(n9269) );
  NAND2_X1 U5786 ( .A1(n9338), .A2(n4748), .ZN(n9297) );
  NOR2_X1 U5787 ( .A1(n9348), .A2(n9925), .ZN(n9338) );
  NAND2_X1 U5788 ( .A1(n9338), .A2(n9922), .ZN(n9319) );
  NAND2_X1 U5789 ( .A1(n4817), .A2(n4826), .ZN(n4816) );
  INV_X1 U5790 ( .A(n4821), .ZN(n4817) );
  OR2_X1 U5791 ( .A1(n6193), .A2(n6176), .ZN(n6219) );
  OR2_X1 U5792 ( .A1(n6219), .A2(n6218), .ZN(n6234) );
  AOI21_X1 U5793 ( .B1(n4907), .B2(n8036), .A(n4905), .ZN(n4904) );
  INV_X1 U5794 ( .A(n4907), .ZN(n4906) );
  INV_X1 U5795 ( .A(n9104), .ZN(n4905) );
  NAND2_X1 U5796 ( .A1(n4759), .A2(n4496), .ZN(n9350) );
  NAND2_X1 U5797 ( .A1(n4759), .A2(n4760), .ZN(n8041) );
  INV_X1 U5798 ( .A(n7994), .ZN(n7987) );
  NOR2_X1 U5799 ( .A1(n7864), .A2(n4761), .ZN(n8002) );
  NAND2_X1 U5800 ( .A1(n4910), .A2(n4913), .ZN(n7992) );
  NAND2_X1 U5801 ( .A1(n7847), .A2(n4917), .ZN(n4910) );
  NOR2_X1 U5802 ( .A1(n7864), .A2(n7881), .ZN(n7895) );
  NAND2_X1 U5803 ( .A1(n5943), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n6147) );
  INV_X1 U5804 ( .A(n6145), .ZN(n5943) );
  AND4_X1 U5805 ( .A1(n6100), .A2(n6099), .A3(n6098), .A4(n6097), .ZN(n7797)
         );
  AND4_X1 U5806 ( .A1(n6138), .A2(n6137), .A3(n6136), .A4(n6135), .ZN(n7890)
         );
  NAND2_X1 U5807 ( .A1(n5940), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n6106) );
  INV_X1 U5808 ( .A(n6081), .ZN(n5940) );
  NAND2_X1 U5809 ( .A1(n5941), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6108) );
  INV_X1 U5810 ( .A(n6106), .ZN(n5941) );
  NAND2_X1 U5811 ( .A1(n4930), .A2(n4934), .ZN(n7616) );
  NAND2_X1 U5812 ( .A1(n7704), .A2(n7527), .ZN(n4930) );
  NOR2_X1 U5813 ( .A1(n9374), .A2(n7701), .ZN(n7698) );
  OR2_X1 U5814 ( .A1(n9376), .A2(n10176), .ZN(n9374) );
  AND2_X1 U5815 ( .A1(n6503), .A2(n6426), .ZN(n9380) );
  NOR2_X1 U5816 ( .A1(n7390), .A2(n7322), .ZN(n7318) );
  NAND2_X1 U5817 ( .A1(n6538), .A2(n7318), .ZN(n9376) );
  NAND2_X1 U5818 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n6067) );
  AND4_X1 U5819 ( .A1(n6072), .A2(n6071), .A3(n6070), .A4(n6069), .ZN(n7558)
         );
  NAND2_X1 U5820 ( .A1(n5917), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n4751) );
  NAND2_X1 U5821 ( .A1(n6258), .A2(n6257), .ZN(n9442) );
  NAND2_X1 U5822 ( .A1(n6003), .A2(n6002), .ZN(n9458) );
  AND2_X1 U5823 ( .A1(n7260), .A2(n7524), .ZN(n10125) );
  XNOR2_X1 U5824 ( .A(n5691), .B(n5690), .ZN(n8863) );
  NAND2_X1 U5825 ( .A1(n5688), .A2(n5687), .ZN(n5691) );
  XNOR2_X1 U5826 ( .A(n5683), .B(SI_30_), .ZN(n8136) );
  XNOR2_X1 U5827 ( .A(n5651), .B(n5650), .ZN(n8872) );
  NAND2_X1 U5828 ( .A1(n5617), .A2(n5616), .ZN(n5630) );
  XNOR2_X1 U5829 ( .A(n5594), .B(n5593), .ZN(n7945) );
  NAND2_X1 U5830 ( .A1(n5562), .A2(n5561), .ZN(n5576) );
  NAND2_X1 U5831 ( .A1(n5545), .A2(n5544), .ZN(n5552) );
  NAND2_X1 U5832 ( .A1(n5910), .A2(n5072), .ZN(n6484) );
  OAI21_X1 U5833 ( .B1(n5453), .B2(n5468), .A(n4985), .ZN(n5490) );
  XNOR2_X1 U5834 ( .A(n5470), .B(n5468), .ZN(n7234) );
  INV_X1 U5835 ( .A(n4990), .ZN(n5434) );
  AOI21_X1 U5836 ( .B1(n5391), .B2(n4995), .A(n4993), .ZN(n4990) );
  NAND2_X1 U5837 ( .A1(n4974), .A2(n5328), .ZN(n5348) );
  AND2_X1 U5838 ( .A1(n5277), .A2(n5265), .ZN(n5276) );
  NAND2_X1 U5839 ( .A1(n5260), .A2(SI_7_), .ZN(n5261) );
  NAND2_X1 U5840 ( .A1(n5258), .A2(n5257), .ZN(n5262) );
  XNOR2_X1 U5841 ( .A(n5213), .B(n9680), .ZN(n5218) );
  XNOR2_X1 U5842 ( .A(n4630), .B(n5160), .ZN(n5177) );
  NAND2_X1 U5843 ( .A1(n7497), .A2(n7496), .ZN(n7505) );
  OAI21_X1 U5844 ( .B1(n8266), .B2(n4871), .A(n4869), .ZN(n8242) );
  INV_X1 U5845 ( .A(n4870), .ZN(n4869) );
  OAI21_X1 U5846 ( .B1(n4561), .B2(n4871), .A(n8204), .ZN(n4870) );
  INV_X1 U5847 ( .A(n8203), .ZN(n4871) );
  NAND2_X1 U5848 ( .A1(n8097), .A2(n8096), .ZN(n8160) );
  AND4_X1 U5849 ( .A1(n5274), .A2(n5273), .A3(n5272), .A4(n5271), .ZN(n7807)
         );
  NAND2_X1 U5850 ( .A1(n4860), .A2(n7742), .ZN(n7755) );
  NAND2_X1 U5851 ( .A1(n7650), .A2(n4503), .ZN(n4860) );
  INV_X1 U5852 ( .A(n10302), .ZN(n8226) );
  NAND2_X1 U5853 ( .A1(n8330), .A2(n4884), .ZN(n8231) );
  NAND2_X1 U5854 ( .A1(n8242), .A2(n8241), .ZN(n8247) );
  NAND2_X1 U5855 ( .A1(n8150), .A2(n5692), .ZN(n5634) );
  OAI21_X1 U5856 ( .B1(n8366), .B2(n4856), .A(n4854), .ZN(n7022) );
  OR2_X1 U5857 ( .A1(n7043), .A2(n9847), .ZN(n4854) );
  NAND2_X1 U5858 ( .A1(n4876), .A2(n4874), .ZN(n8258) );
  AOI21_X1 U5859 ( .B1(n4877), .B2(n4879), .A(n4875), .ZN(n4874) );
  INV_X1 U5860 ( .A(n4880), .ZN(n4879) );
  NAND2_X1 U5861 ( .A1(n4610), .A2(n7911), .ZN(n7959) );
  NAND2_X1 U5862 ( .A1(n4615), .A2(n4528), .ZN(n8293) );
  NAND2_X1 U5863 ( .A1(n4616), .A2(n4848), .ZN(n4615) );
  NAND2_X1 U5864 ( .A1(n5440), .A2(n5439), .ZN(n8816) );
  NAND2_X1 U5865 ( .A1(n7148), .A2(n7147), .ZN(n7293) );
  NAND2_X1 U5866 ( .A1(n7650), .A2(n7649), .ZN(n7743) );
  NAND2_X1 U5867 ( .A1(n5285), .A2(n5284), .ZN(n7839) );
  AND2_X1 U5868 ( .A1(n7151), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8344) );
  AND2_X1 U5869 ( .A1(n8231), .A2(n4880), .ZN(n8310) );
  NAND2_X1 U5870 ( .A1(n8231), .A2(n4882), .ZN(n8311) );
  NAND2_X1 U5871 ( .A1(n7962), .A2(n7963), .ZN(n8097) );
  XNOR2_X1 U5872 ( .A(n8183), .B(n4560), .ZN(n8318) );
  NAND2_X1 U5873 ( .A1(n4857), .A2(n4861), .ZN(n7907) );
  OR2_X1 U5874 ( .A1(n7650), .A2(n4863), .ZN(n4857) );
  NAND2_X1 U5875 ( .A1(n7293), .A2(n4866), .ZN(n7342) );
  NAND2_X1 U5876 ( .A1(n7342), .A2(n7299), .ZN(n7497) );
  INV_X1 U5877 ( .A(n8768), .ZN(n8562) );
  OR3_X1 U5878 ( .A1(n5872), .A2(n5838), .A3(n5837), .ZN(n5087) );
  AND2_X1 U5879 ( .A1(n5704), .A2(n5703), .ZN(n5880) );
  INV_X1 U5880 ( .A(P2_U3966), .ZN(n8384) );
  OR2_X1 U5881 ( .A1(n7114), .A2(n7113), .ZN(n7115) );
  NOR2_X1 U5882 ( .A1(n7182), .A2(n4562), .ZN(n7160) );
  NOR2_X1 U5883 ( .A1(n7160), .A2(n7159), .ZN(n7158) );
  NOR2_X1 U5884 ( .A1(n7158), .A2(n4774), .ZN(n7093) );
  AND2_X1 U5885 ( .A1(n7088), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n4774) );
  NOR2_X1 U5886 ( .A1(n7093), .A2(n7092), .ZN(n7272) );
  AND2_X1 U5887 ( .A1(n7485), .A2(n8402), .ZN(n7486) );
  NAND2_X1 U5888 ( .A1(n7486), .A2(n7487), .ZN(n7674) );
  NOR2_X1 U5889 ( .A1(n4772), .A2(n4771), .ZN(n7675) );
  INV_X1 U5890 ( .A(n7673), .ZN(n4771) );
  INV_X1 U5891 ( .A(n7674), .ZN(n4772) );
  NAND2_X1 U5892 ( .A1(n7674), .A2(n4773), .ZN(n7725) );
  NOR2_X1 U5893 ( .A1(n8450), .A2(n8449), .ZN(n8467) );
  AOI22_X1 U5894 ( .A1(n8136), .A2(n5692), .B1(P1_DATAO_REG_30__SCAN_IN), .B2(
        n5669), .ZN(n9906) );
  NAND2_X1 U5895 ( .A1(n5024), .A2(n5023), .ZN(n8596) );
  AND2_X1 U5896 ( .A1(n5024), .A2(n4501), .ZN(n8598) );
  NAND2_X1 U5897 ( .A1(n8608), .A2(n5798), .ZN(n8592) );
  AND2_X1 U5898 ( .A1(n5536), .A2(n5535), .ZN(n8632) );
  NAND2_X1 U5899 ( .A1(n8661), .A2(n5085), .ZN(n8646) );
  INV_X1 U5900 ( .A(n4644), .ZN(n8698) );
  AOI21_X1 U5901 ( .B1(n5432), .B2(n4645), .A(n4646), .ZN(n4644) );
  INV_X1 U5902 ( .A(n8809), .ZN(n8697) );
  NAND2_X1 U5903 ( .A1(n5432), .A2(n5767), .ZN(n8713) );
  NAND2_X1 U5904 ( .A1(n5029), .A2(n5028), .ZN(n8710) );
  NAND2_X1 U5905 ( .A1(n4939), .A2(n4941), .ZN(n8106) );
  OR2_X1 U5906 ( .A1(n8014), .A2(n4944), .ZN(n4939) );
  NAND2_X1 U5907 ( .A1(n5398), .A2(n5397), .ZN(n8495) );
  NAND2_X1 U5908 ( .A1(n8048), .A2(n5089), .ZN(n8113) );
  NAND2_X1 U5909 ( .A1(n4954), .A2(n5855), .ZN(n7924) );
  OAI21_X1 U5910 ( .B1(n7810), .B2(n4638), .A(n4636), .ZN(n4954) );
  NAND2_X1 U5911 ( .A1(n7811), .A2(n5749), .ZN(n7766) );
  NAND2_X1 U5912 ( .A1(n7682), .A2(n7681), .ZN(n7763) );
  AND3_X1 U5913 ( .A1(n5240), .A2(n5239), .A3(n5238), .ZN(n7591) );
  NAND2_X1 U5914 ( .A1(n10250), .A2(n5201), .ZN(n4948) );
  NAND2_X1 U5915 ( .A1(n5013), .A2(n7373), .ZN(n7442) );
  INV_X1 U5916 ( .A(n8733), .ZN(n8486) );
  NOR2_X1 U5917 ( .A1(n8751), .A2(n8750), .ZN(n8752) );
  AOI211_X1 U5918 ( .C1(n10284), .C2(n8768), .A(n8767), .B(n8766), .ZN(n8769)
         );
  XNOR2_X1 U5919 ( .A(n5106), .B(n8864), .ZN(n5109) );
  NAND2_X1 U5920 ( .A1(n8868), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5106) );
  NAND2_X1 U5921 ( .A1(n8868), .A2(n5108), .ZN(n8873) );
  MUX2_X1 U5922 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5107), .S(
        P2_IR_REG_29__SCAN_IN), .Z(n5108) );
  XNOR2_X1 U5923 ( .A(n5119), .B(n5118), .ZN(n8484) );
  NAND2_X1 U5924 ( .A1(n4703), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5119) );
  AND2_X1 U5925 ( .A1(n4949), .A2(n4545), .ZN(n4701) );
  INV_X1 U5926 ( .A(n6987), .ZN(n7578) );
  AND3_X1 U5927 ( .A1(n5045), .A2(n5044), .A3(n5101), .ZN(n5454) );
  INV_X1 U5928 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6812) );
  INV_X1 U5929 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6801) );
  AOI22_X1 U5930 ( .A1(n4538), .A2(P2_IR_REG_0__SCAN_IN), .B1(n4784), .B2(
        n5162), .ZN(n4783) );
  INV_X1 U5931 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n4784) );
  NAND2_X1 U5932 ( .A1(n6593), .A2(n7551), .ZN(n7568) );
  NAND2_X1 U5933 ( .A1(n4715), .A2(n4716), .ZN(n8125) );
  NAND2_X1 U5934 ( .A1(n8068), .A2(n5078), .ZN(n4715) );
  NAND2_X1 U5935 ( .A1(n4707), .A2(n6732), .ZN(n4705) );
  OR2_X1 U5936 ( .A1(n8989), .A2(n4706), .ZN(n4704) );
  NAND2_X1 U5937 ( .A1(n4707), .A2(n4608), .ZN(n4706) );
  INV_X1 U5938 ( .A(n6778), .ZN(n6779) );
  AOI211_X1 U5939 ( .C1(n9400), .C2(n9007), .A(n6777), .B(n6776), .ZN(n6778)
         );
  NAND2_X1 U5940 ( .A1(n4602), .A2(n4606), .ZN(n7639) );
  NAND2_X1 U5941 ( .A1(n7568), .A2(n4607), .ZN(n4602) );
  NAND2_X1 U5942 ( .A1(n4596), .A2(n5056), .ZN(n8912) );
  NAND2_X1 U5943 ( .A1(n8901), .A2(n5054), .ZN(n4596) );
  NAND2_X1 U5944 ( .A1(n5063), .A2(n5064), .ZN(n8920) );
  OR2_X1 U5945 ( .A1(n8891), .A2(n5065), .ZN(n5063) );
  NAND2_X1 U5946 ( .A1(n5066), .A2(n6715), .ZN(n8946) );
  NAND2_X1 U5947 ( .A1(n8891), .A2(n5070), .ZN(n5066) );
  AND2_X1 U5948 ( .A1(n7206), .A2(n7205), .ZN(n6576) );
  OR2_X1 U5949 ( .A1(n6062), .A2(n6805), .ZN(n6064) );
  NAND2_X1 U5950 ( .A1(n5051), .A2(n5050), .ZN(n7794) );
  INV_X1 U5951 ( .A(n5053), .ZN(n5050) );
  NAND2_X1 U5952 ( .A1(n7639), .A2(n5052), .ZN(n5051) );
  NAND2_X1 U5953 ( .A1(n8954), .A2(n8955), .ZN(n8953) );
  NAND2_X1 U5954 ( .A1(n8900), .A2(n8902), .ZN(n8954) );
  AND2_X1 U5955 ( .A1(n6765), .A2(n6754), .ZN(n8956) );
  NAND2_X1 U5956 ( .A1(n6709), .A2(n6708), .ZN(n8969) );
  NAND2_X1 U5957 ( .A1(n6281), .A2(n6280), .ZN(n9432) );
  AND4_X1 U5958 ( .A1(n6128), .A2(n6127), .A3(n6126), .A4(n6125), .ZN(n8082)
         );
  NAND2_X1 U5959 ( .A1(n5047), .A2(n7827), .ZN(n7937) );
  NAND2_X1 U5960 ( .A1(n6559), .A2(n4590), .ZN(n4589) );
  INV_X1 U5961 ( .A(n8956), .ZN(n9009) );
  INV_X1 U5962 ( .A(n7557), .ZN(n9018) );
  NAND2_X1 U5963 ( .A1(n6942), .A2(n6943), .ZN(n6941) );
  NAND2_X1 U5964 ( .A1(n6936), .A2(n4575), .ZN(n9975) );
  NAND2_X1 U5965 ( .A1(n6941), .A2(n4734), .ZN(n9968) );
  NAND2_X1 U5966 ( .A1(n4735), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n4734) );
  NAND2_X1 U5967 ( .A1(n6961), .A2(n4522), .ZN(n10016) );
  INV_X1 U5968 ( .A(n4742), .ZN(n9024) );
  INV_X1 U5969 ( .A(n4740), .ZN(n10084) );
  INV_X1 U5970 ( .A(n4738), .ZN(n10098) );
  NAND2_X1 U5971 ( .A1(n10090), .A2(n4570), .ZN(n10103) );
  NOR2_X1 U5972 ( .A1(n9064), .A2(n4765), .ZN(n4763) );
  OAI21_X1 U5973 ( .B1(n9194), .B2(n4832), .A(n4830), .ZN(n9156) );
  AOI21_X1 U5974 ( .B1(n9174), .B2(n10133), .A(n9173), .ZN(n9413) );
  OAI21_X1 U5975 ( .B1(n9187), .B2(n9121), .A(n9120), .ZN(n9171) );
  NAND2_X1 U5976 ( .A1(n4833), .A2(n4836), .ZN(n9170) );
  AOI21_X1 U5977 ( .B1(n9190), .B2(n10133), .A(n9189), .ZN(n9418) );
  OAI21_X1 U5978 ( .B1(n9194), .B2(n4505), .A(n4843), .ZN(n9181) );
  NAND2_X1 U5979 ( .A1(n6273), .A2(n6272), .ZN(n9439) );
  NAND2_X1 U5980 ( .A1(n4925), .A2(n4927), .ZN(n9243) );
  NAND2_X1 U5981 ( .A1(n4926), .A2(n9113), .ZN(n9262) );
  OR2_X1 U5982 ( .A1(n9274), .A2(n9273), .ZN(n4926) );
  INV_X1 U5983 ( .A(n4805), .ZN(n9255) );
  AOI21_X1 U5984 ( .B1(n9281), .B2(n4809), .A(n4807), .ZN(n4805) );
  INV_X1 U5985 ( .A(n4814), .ZN(n4810) );
  NAND2_X1 U5986 ( .A1(n9281), .A2(n9288), .ZN(n4812) );
  NAND2_X1 U5987 ( .A1(n4823), .A2(n9074), .ZN(n9328) );
  NAND2_X1 U5988 ( .A1(n4909), .A2(n4907), .ZN(n9360) );
  NAND2_X1 U5989 ( .A1(n4909), .A2(n9103), .ZN(n9358) );
  NAND2_X1 U5990 ( .A1(n6155), .A2(n6154), .ZN(n7986) );
  NAND2_X1 U5991 ( .A1(n7883), .A2(n7882), .ZN(n7985) );
  OAI21_X1 U5992 ( .B1(n7847), .B2(n7846), .A(n7848), .ZN(n7888) );
  NAND2_X1 U5993 ( .A1(n6144), .A2(n6143), .ZN(n7853) );
  NAND2_X1 U5994 ( .A1(n7695), .A2(n7545), .ZN(n7625) );
  AND2_X1 U5995 ( .A1(n10179), .A2(n7543), .ZN(n7697) );
  OAI21_X1 U5996 ( .B1(n6117), .B2(n4735), .A(n4886), .ZN(n4888) );
  NAND2_X1 U5997 ( .A1(n6117), .A2(n4887), .ZN(n4886) );
  OR2_X1 U5998 ( .A1(n6951), .A2(n6969), .ZN(n10151) );
  CLKBUF_X1 U5999 ( .A(n6480), .Z(n8151) );
  INV_X1 U6000 ( .A(n7246), .ZN(n7660) );
  INV_X1 U6001 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n9806) );
  XNOR2_X1 U6002 ( .A(n4629), .B(n5276), .ZN(n6811) );
  NAND2_X1 U6003 ( .A1(n5262), .A2(n5261), .ZN(n4629) );
  INV_X1 U6004 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n9833) );
  INV_X1 U6005 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n9657) );
  AND2_X1 U6006 ( .A1(n5220), .A2(n5219), .ZN(n5233) );
  XNOR2_X1 U6007 ( .A(n5196), .B(n5195), .ZN(n6805) );
  AND2_X1 U6008 ( .A1(n4658), .A2(n4502), .ZN(n5196) );
  NAND2_X1 U6009 ( .A1(n4483), .A2(SI_0_), .ZN(n6028) );
  AND2_X1 U6010 ( .A1(P2_ADDR_REG_19__SCAN_IN), .A2(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n9888) );
  AND2_X1 U6011 ( .A1(n7029), .A2(n7028), .ZN(n7033) );
  INV_X1 U6012 ( .A(n4786), .ZN(n7170) );
  INV_X1 U6013 ( .A(n8482), .ZN(n4777) );
  NAND2_X1 U6014 ( .A1(n4779), .A2(n8478), .ZN(n4778) );
  NAND2_X1 U6015 ( .A1(n4782), .A2(n4781), .ZN(n4780) );
  OAI21_X1 U6016 ( .B1(n8733), .B2(n4856), .A(n4855), .ZN(n7231) );
  OR2_X1 U6017 ( .A1(n10360), .A2(n4650), .ZN(n4649) );
  NAND2_X1 U6018 ( .A1(n8845), .A2(n10360), .ZN(n4651) );
  INV_X1 U6019 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n4650) );
  AOI21_X1 U6020 ( .B1(n10068), .B2(P1_ADDR_REG_19__SCAN_IN), .A(n9057), .ZN(
        n4744) );
  OR2_X1 U6021 ( .A1(n9051), .A2(n10138), .ZN(n4573) );
  OR2_X1 U6022 ( .A1(n7927), .A2(n4726), .ZN(n4488) );
  XNOR2_X1 U6023 ( .A(n7680), .B(n8377), .ZN(n7597) );
  NAND2_X1 U6024 ( .A1(n7301), .A2(n10259), .ZN(n5712) );
  OR2_X1 U6025 ( .A1(n8015), .A2(n5036), .ZN(n4489) );
  AND2_X1 U6026 ( .A1(n5103), .A2(n5046), .ZN(n4490) );
  AND2_X1 U6027 ( .A1(n5064), .A2(n5062), .ZN(n4491) );
  AND2_X1 U6028 ( .A1(n5984), .A2(n7351), .ZN(n4492) );
  AND2_X1 U6029 ( .A1(n4540), .A2(n5103), .ZN(n4493) );
  INV_X1 U6030 ( .A(n5798), .ZN(n4688) );
  NAND2_X1 U6031 ( .A1(n9421), .A2(n9089), .ZN(n9119) );
  INV_X1 U6032 ( .A(n9119), .ZN(n4892) );
  NAND2_X1 U6033 ( .A1(n5266), .A2(n4657), .ZN(n7680) );
  INV_X1 U6034 ( .A(n7589), .ZN(n5241) );
  NAND2_X1 U6035 ( .A1(n5964), .A2(n5963), .ZN(n9421) );
  INV_X1 U6036 ( .A(n9421), .ZN(n9090) );
  NAND2_X1 U6037 ( .A1(n6022), .A2(n6021), .ZN(n6939) );
  INV_X1 U6038 ( .A(n6939), .ZN(n4735) );
  NOR2_X1 U6039 ( .A1(n9123), .A2(n6321), .ZN(n4903) );
  INV_X1 U6040 ( .A(n4903), .ZN(n4896) );
  AND2_X1 U6041 ( .A1(n5072), .A2(n4525), .ZN(n4494) );
  AND2_X1 U6042 ( .A1(n5868), .A2(n4692), .ZN(n4495) );
  NAND2_X1 U6043 ( .A1(n5359), .A2(n5358), .ZN(n8024) );
  AND2_X1 U6044 ( .A1(n4760), .A2(n4762), .ZN(n4496) );
  NAND2_X1 U6045 ( .A1(n6354), .A2(n6353), .ZN(n9064) );
  OR2_X1 U6046 ( .A1(n5912), .A2(P1_IR_REG_27__SCAN_IN), .ZN(n4497) );
  AND2_X1 U6047 ( .A1(n4748), .A2(n4747), .ZN(n4498) );
  NAND2_X1 U6048 ( .A1(n9124), .A2(n6457), .ZN(n9164) );
  INV_X1 U6049 ( .A(n9164), .ZN(n4899) );
  OAI21_X1 U6050 ( .B1(n4830), .B2(n4899), .A(n4539), .ZN(n4828) );
  NAND2_X2 U6051 ( .A1(n6988), .A2(n7221), .ZN(n7953) );
  INV_X1 U6052 ( .A(n8069), .ZN(n5075) );
  NAND2_X1 U6053 ( .A1(n7402), .A2(n7404), .ZN(n7403) );
  AND4_X1 U6054 ( .A1(n5138), .A2(n5137), .A3(n5136), .A4(n5135), .ZN(n7361)
         );
  INV_X1 U6055 ( .A(n7361), .ZN(n5020) );
  INV_X1 U6056 ( .A(n6563), .ZN(n6046) );
  OR2_X1 U6057 ( .A1(n6047), .A2(n6836), .ZN(n4499) );
  AND2_X1 U6058 ( .A1(n4624), .A2(n4868), .ZN(n4500) );
  NAND2_X1 U6059 ( .A1(n8784), .A2(n8505), .ZN(n4501) );
  OR2_X1 U6060 ( .A1(n5178), .A2(n5177), .ZN(n4502) );
  OAI211_X1 U6061 ( .C1(n5142), .C2(n7191), .A(n5223), .B(n5222), .ZN(n7453)
         );
  INV_X1 U6062 ( .A(n5079), .ZN(n5078) );
  OR2_X1 U6063 ( .A1(n6635), .A2(n5080), .ZN(n5079) );
  AOI21_X1 U6064 ( .B1(n9426), .B2(n6608), .A(n6714), .ZN(n8888) );
  AND2_X1 U6065 ( .A1(n4865), .A2(n7649), .ZN(n4503) );
  AND2_X1 U6066 ( .A1(n4806), .A2(n9081), .ZN(n4504) );
  NOR2_X1 U6067 ( .A1(n9090), .A2(n9089), .ZN(n4505) );
  NAND2_X1 U6068 ( .A1(n5118), .A2(n4702), .ZN(n4506) );
  OR2_X1 U6069 ( .A1(n6948), .A2(n6712), .ZN(n4507) );
  OR2_X1 U6070 ( .A1(n5142), .A2(n7135), .ZN(n4508) );
  AND2_X1 U6071 ( .A1(n4613), .A2(n7140), .ZN(n4509) );
  AND2_X1 U6072 ( .A1(n8543), .A2(n5808), .ZN(n4510) );
  NAND2_X1 U6073 ( .A1(n5622), .A2(n5621), .ZN(n8194) );
  AND2_X1 U6074 ( .A1(n4742), .A2(n4741), .ZN(n4511) );
  XNOR2_X1 U6075 ( .A(n5630), .B(n5629), .ZN(n6312) );
  INV_X1 U6076 ( .A(n8879), .ZN(n4708) );
  AND2_X1 U6077 ( .A1(n9411), .A2(n7351), .ZN(n4512) );
  NAND2_X1 U6078 ( .A1(n6314), .A2(n6313), .ZN(n9405) );
  OR2_X1 U6079 ( .A1(n5142), .A2(n7281), .ZN(n4513) );
  OR3_X1 U6080 ( .A1(n5476), .A2(P2_IR_REG_19__SCAN_IN), .A3(
        P2_IR_REG_20__SCAN_IN), .ZN(n4514) );
  OR2_X1 U6081 ( .A1(n9416), .A2(n9092), .ZN(n9120) );
  NAND2_X1 U6082 ( .A1(n6231), .A2(n6230), .ZN(n9323) );
  NAND2_X1 U6083 ( .A1(n5803), .A2(n5804), .ZN(n8580) );
  INV_X1 U6084 ( .A(n8580), .ZN(n4681) );
  AND2_X1 U6085 ( .A1(n5852), .A2(n5854), .ZN(n4515) );
  NOR2_X1 U6086 ( .A1(n5831), .A2(n5828), .ZN(n4516) );
  AND2_X1 U6087 ( .A1(n6392), .A2(n9103), .ZN(n9101) );
  NAND2_X1 U6088 ( .A1(n5910), .A2(n5071), .ZN(n6471) );
  NAND2_X1 U6089 ( .A1(n5910), .A2(n5909), .ZN(n6482) );
  AND2_X1 U6090 ( .A1(n4829), .A2(n9164), .ZN(n4517) );
  AND2_X1 U6091 ( .A1(n8159), .A2(n8158), .ZN(n4518) );
  AND2_X1 U6092 ( .A1(n9447), .A2(n9290), .ZN(n4519) );
  AND2_X1 U6093 ( .A1(n5973), .A2(n5972), .ZN(n9089) );
  INV_X1 U6094 ( .A(n9426), .ZN(n9086) );
  NAND2_X1 U6095 ( .A1(n5975), .A2(n5974), .ZN(n9426) );
  INV_X1 U6096 ( .A(n8794), .ZN(n8652) );
  NAND2_X1 U6097 ( .A1(n5512), .A2(n5511), .ZN(n8794) );
  AND2_X1 U6098 ( .A1(n5219), .A2(n5232), .ZN(n4520) );
  NAND2_X1 U6099 ( .A1(n8663), .A2(n4722), .ZN(n4723) );
  AND2_X1 U6100 ( .A1(n6618), .A2(n7827), .ZN(n4521) );
  OR2_X1 U6101 ( .A1(n6964), .A2(n10226), .ZN(n4522) );
  AND2_X1 U6102 ( .A1(n4612), .A2(n7140), .ZN(n4523) );
  AND2_X1 U6103 ( .A1(n5615), .A2(n5803), .ZN(n4524) );
  AOI21_X1 U6104 ( .B1(n4850), .B2(n4852), .A(n4849), .ZN(n4848) );
  NOR2_X1 U6105 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n4525) );
  AND2_X1 U6106 ( .A1(n8495), .A2(n8281), .ZN(n4526) );
  AND2_X1 U6107 ( .A1(n6672), .A2(n6668), .ZN(n4527) );
  AND2_X1 U6108 ( .A1(n4614), .A2(n8164), .ZN(n4528) );
  OR2_X1 U6109 ( .A1(n8799), .A2(n8503), .ZN(n5789) );
  AND2_X1 U6110 ( .A1(n4925), .A2(n4923), .ZN(n4529) );
  NAND2_X1 U6111 ( .A1(n5801), .A2(n5797), .ZN(n8597) );
  AND2_X1 U6112 ( .A1(n7807), .A2(n7761), .ZN(n4530) );
  NOR2_X1 U6113 ( .A1(n7986), .A2(n9014), .ZN(n4531) );
  AND2_X1 U6114 ( .A1(n7459), .A2(n7680), .ZN(n4532) );
  INV_X1 U6115 ( .A(n4898), .ZN(n4897) );
  NAND2_X1 U6116 ( .A1(n4900), .A2(n4899), .ZN(n4898) );
  NOR2_X1 U6117 ( .A1(n8778), .A2(n8610), .ZN(n4533) );
  NAND2_X1 U6118 ( .A1(n6700), .A2(n6699), .ZN(n4534) );
  INV_X1 U6119 ( .A(n5081), .ZN(n4717) );
  AND2_X1 U6120 ( .A1(n9094), .A2(n9093), .ZN(n4535) );
  NAND2_X1 U6121 ( .A1(n5104), .A2(n4493), .ZN(n4536) );
  INV_X1 U6122 ( .A(n4765), .ZN(n4764) );
  NAND2_X1 U6123 ( .A1(n4766), .A2(n9394), .ZN(n4765) );
  NAND2_X1 U6124 ( .A1(n6659), .A2(n6658), .ZN(n4537) );
  AND2_X1 U6125 ( .A1(n8499), .A2(n5448), .ZN(n8712) );
  NAND2_X1 U6126 ( .A1(n6248), .A2(n6247), .ZN(n9447) );
  AND2_X1 U6127 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n4538) );
  NAND2_X1 U6128 ( .A1(n9162), .A2(n9095), .ZN(n4539) );
  NOR2_X1 U6129 ( .A1(n8889), .A2(n8888), .ZN(n6716) );
  AND2_X1 U6130 ( .A1(n5105), .A2(n5091), .ZN(n4540) );
  NAND2_X1 U6131 ( .A1(n4837), .A2(n4842), .ZN(n4836) );
  NAND2_X1 U6132 ( .A1(n6348), .A2(n6347), .ZN(n9134) );
  OR2_X1 U6133 ( .A1(n8080), .A2(n8079), .ZN(n5081) );
  OR2_X1 U6134 ( .A1(n9442), .A2(n9082), .ZN(n9114) );
  AND2_X1 U6135 ( .A1(n5054), .A2(n8911), .ZN(n4541) );
  OR2_X1 U6136 ( .A1(n5476), .A2(P2_IR_REG_19__SCAN_IN), .ZN(n4542) );
  AND2_X1 U6137 ( .A1(n5756), .A2(n8049), .ZN(n8015) );
  INV_X1 U6138 ( .A(n8015), .ZN(n4943) );
  AND3_X1 U6139 ( .A1(n5164), .A2(n5101), .A3(n5457), .ZN(n4543) );
  AND2_X1 U6140 ( .A1(n4812), .A2(n4810), .ZN(n4544) );
  AND4_X1 U6141 ( .A1(n5115), .A2(n5114), .A3(n5113), .A4(n5112), .ZN(n8223)
         );
  AND2_X1 U6142 ( .A1(n4950), .A2(n4702), .ZN(n4545) );
  OR2_X1 U6143 ( .A1(n6959), .A2(n6960), .ZN(n4546) );
  AND2_X1 U6144 ( .A1(n5853), .A2(n5855), .ZN(n4953) );
  AND2_X1 U6145 ( .A1(n7414), .A2(n10308), .ZN(n4547) );
  NOR2_X1 U6146 ( .A1(n6327), .A2(n4512), .ZN(n4548) );
  OR2_X1 U6147 ( .A1(n4781), .A2(n5870), .ZN(n4549) );
  NAND2_X1 U6148 ( .A1(n8123), .A2(n6645), .ZN(n4550) );
  AND4_X1 U6149 ( .A1(n5292), .A2(n5291), .A3(n5290), .A4(n5289), .ZN(n7768)
         );
  INV_X1 U6150 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n4702) );
  NAND2_X1 U6151 ( .A1(n8820), .A2(n8498), .ZN(n4551) );
  NAND2_X1 U6152 ( .A1(n6404), .A2(n6366), .ZN(n4552) );
  INV_X1 U6153 ( .A(n9094), .ZN(n9411) );
  AND2_X1 U6154 ( .A1(n6307), .A2(n6306), .ZN(n9094) );
  AND2_X1 U6155 ( .A1(n8543), .A2(n5809), .ZN(n4553) );
  AND2_X1 U6156 ( .A1(n5815), .A2(n5816), .ZN(n4554) );
  AND2_X1 U6157 ( .A1(n5555), .A2(n5554), .ZN(n8618) );
  INV_X1 U6158 ( .A(n8618), .ZN(n8784) );
  AND2_X1 U6159 ( .A1(n9272), .A2(n4498), .ZN(n4555) );
  AND2_X1 U6160 ( .A1(n4900), .A2(n4893), .ZN(n4556) );
  AND2_X1 U6161 ( .A1(n5350), .A2(n5328), .ZN(n4557) );
  INV_X1 U6162 ( .A(n5088), .ZN(n5069) );
  INV_X1 U6163 ( .A(n8483), .ZN(n8748) );
  NAND2_X1 U6164 ( .A1(n5653), .A2(n5652), .ZN(n8483) );
  AND2_X1 U6165 ( .A1(n4635), .A2(n4953), .ZN(n4558) );
  INV_X1 U6166 ( .A(n4935), .ZN(n4934) );
  NAND2_X1 U6167 ( .A1(n7529), .A2(n4936), .ZN(n4935) );
  INV_X1 U6168 ( .A(n4914), .ZN(n4913) );
  NAND2_X1 U6169 ( .A1(n4915), .A2(n7886), .ZN(n4914) );
  AND2_X1 U6170 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n4559) );
  XNOR2_X1 U6171 ( .A(n5326), .B(SI_11_), .ZN(n5324) );
  XOR2_X1 U6172 ( .A(n8632), .B(n7953), .Z(n4560) );
  NOR2_X1 U6173 ( .A1(n8011), .A2(n8010), .ZN(n5038) );
  INV_X1 U6174 ( .A(n8990), .ZN(n4608) );
  NAND2_X1 U6175 ( .A1(n5565), .A2(n5564), .ZN(n8778) );
  INV_X1 U6176 ( .A(n8778), .ZN(n4720) );
  INV_X1 U6177 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n4580) );
  INV_X1 U6178 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n4584) );
  INV_X1 U6179 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n4632) );
  NOR2_X1 U6180 ( .A1(n8342), .A2(n4872), .ZN(n4561) );
  NAND2_X1 U6181 ( .A1(n8066), .A2(n6630), .ZN(n8078) );
  INV_X1 U6182 ( .A(n8902), .ZN(n5058) );
  AND2_X1 U6183 ( .A1(n5029), .A2(n4551), .ZN(n8709) );
  NAND2_X1 U6184 ( .A1(n5104), .A2(n5103), .ZN(n5883) );
  NOR3_X1 U6185 ( .A1(n9247), .A2(n9416), .A3(n4756), .ZN(n4753) );
  INV_X1 U6186 ( .A(n7614), .ZN(n4932) );
  NAND2_X1 U6187 ( .A1(n8938), .A2(n4527), .ZN(n8977) );
  NAND2_X1 U6188 ( .A1(n9338), .A2(n4498), .ZN(n4749) );
  INV_X1 U6189 ( .A(n4754), .ZN(n9201) );
  NOR2_X1 U6190 ( .A1(n9247), .A2(n4756), .ZN(n4754) );
  INV_X1 U6191 ( .A(n4725), .ZN(n8117) );
  NOR3_X1 U6192 ( .A1(n7927), .A2(n8111), .A3(n4728), .ZN(n4725) );
  NAND2_X1 U6193 ( .A1(n8889), .A2(n8888), .ZN(n6715) );
  NAND2_X1 U6194 ( .A1(n4718), .A2(n5075), .ZN(n8066) );
  INV_X1 U6195 ( .A(n6732), .ZN(n4710) );
  AND2_X1 U6196 ( .A1(n6731), .A2(n6730), .ZN(n6732) );
  AND2_X1 U6197 ( .A1(n7086), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n4562) );
  INV_X1 U6198 ( .A(SI_0_), .ZN(n4968) );
  AND2_X1 U6199 ( .A1(n5471), .A2(SI_18_), .ZN(n4563) );
  AND2_X1 U6200 ( .A1(n5577), .A2(SI_24_), .ZN(n4564) );
  NOR2_X1 U6201 ( .A1(n6725), .A2(n6724), .ZN(n4565) );
  AND2_X1 U6202 ( .A1(n5521), .A2(n5509), .ZN(n4566) );
  AND2_X1 U6203 ( .A1(n4823), .A2(n4821), .ZN(n4567) );
  AND2_X1 U6204 ( .A1(n4641), .A2(n4639), .ZN(n4568) );
  NAND2_X1 U6205 ( .A1(n5340), .A2(n5339), .ZN(n8009) );
  INV_X1 U6206 ( .A(n8009), .ZN(n4729) );
  NAND2_X1 U6207 ( .A1(n4948), .A2(n5712), .ZN(n7376) );
  AND2_X1 U6208 ( .A1(n9039), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4569) );
  INV_X1 U6209 ( .A(n7742), .ZN(n4864) );
  INV_X1 U6210 ( .A(n9452), .ZN(n4747) );
  INV_X1 U6211 ( .A(n9932), .ZN(n4762) );
  NAND2_X1 U6212 ( .A1(n4601), .A2(n4599), .ZN(n7792) );
  NAND2_X1 U6213 ( .A1(n4945), .A2(n4947), .ZN(n7457) );
  AND2_X1 U6214 ( .A1(n5045), .A2(n5044), .ZN(n5420) );
  NAND2_X1 U6215 ( .A1(n7463), .A2(n7591), .ZN(n7606) );
  INV_X1 U6216 ( .A(n7606), .ZN(n4699) );
  AND2_X1 U6217 ( .A1(n6584), .A2(n7553), .ZN(n7402) );
  OR2_X1 U6218 ( .A1(n9043), .A2(n6232), .ZN(n4570) );
  NAND2_X1 U6219 ( .A1(n5910), .A2(n4494), .ZN(n4571) );
  AND2_X1 U6220 ( .A1(n8448), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n4572) );
  INV_X1 U6221 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n6060) );
  INV_X1 U6222 ( .A(n8478), .ZN(n4781) );
  INV_X1 U6223 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5073) );
  INV_X1 U6224 ( .A(n9892), .ZN(n4788) );
  INV_X1 U6225 ( .A(n4692), .ZN(n4687) );
  NOR2_X1 U6226 ( .A1(n4672), .A2(n5824), .ZN(n4671) );
  AND2_X1 U6227 ( .A1(n5853), .A2(n5824), .ZN(n4675) );
  NAND2_X1 U6228 ( .A1(n7809), .A2(n5824), .ZN(n4690) );
  INV_X1 U6229 ( .A(n5824), .ZN(n4692) );
  NAND3_X1 U6230 ( .A1(n4745), .A2(n4744), .A3(n4573), .ZN(P1_U3260) );
  NOR2_X1 U6231 ( .A1(n6877), .A2(n6876), .ZN(n6895) );
  NOR2_X1 U6232 ( .A1(n6898), .A2(n10018), .ZN(n6900) );
  AOI21_X1 U6233 ( .B1(n6156), .B2(n9037), .A(n10021), .ZN(n10036) );
  AOI21_X1 U6234 ( .B1(n6123), .B2(n9038), .A(n10034), .ZN(n10048) );
  AOI21_X1 U6235 ( .B1(n6189), .B2(n10053), .A(n10046), .ZN(n10061) );
  AOI21_X1 U6236 ( .B1(n9036), .B2(n6132), .A(n9035), .ZN(n10023) );
  OAI21_X1 U6237 ( .B1(n9056), .B2(n9055), .A(n9054), .ZN(n4746) );
  AOI21_X1 U6238 ( .B1(n9040), .B2(n6175), .A(n10059), .ZN(n9041) );
  AOI21_X1 U6239 ( .B1(n9047), .B2(n9046), .A(n10120), .ZN(n9049) );
  AOI21_X1 U6240 ( .B1(n6079), .B2(n6925), .A(n6922), .ZN(n10004) );
  NAND2_X1 U6241 ( .A1(n5220), .A2(n4520), .ZN(n4966) );
  AOI21_X1 U6242 ( .B1(n5386), .B2(n4943), .A(n4942), .ZN(n4941) );
  NAND2_X1 U6243 ( .A1(n9975), .A2(n9974), .ZN(n9973) );
  OR2_X1 U6244 ( .A1(n6939), .A2(n10218), .ZN(n4575) );
  NAND2_X1 U6245 ( .A1(n4746), .A2(n10138), .ZN(n4745) );
  AOI21_X1 U6246 ( .B1(n5820), .B2(n8548), .A(n8515), .ZN(n5823) );
  NAND2_X1 U6247 ( .A1(n5817), .A2(n4554), .ZN(n5820) );
  OAI21_X1 U6248 ( .B1(n4577), .B2(n5780), .A(n4576), .ZN(n5782) );
  OAI21_X1 U6249 ( .B1(n5742), .B2(n5741), .A(n4578), .ZN(n5746) );
  NAND2_X1 U6250 ( .A1(n4677), .A2(n4953), .ZN(n4673) );
  NAND2_X1 U6251 ( .A1(n5087), .A2(n5874), .ZN(n5879) );
  NAND2_X1 U6252 ( .A1(n5755), .A2(n5754), .ZN(n4678) );
  AOI21_X1 U6253 ( .B1(n4684), .B2(n4683), .A(n4680), .ZN(n5811) );
  AOI21_X1 U6254 ( .B1(n5711), .B2(n5710), .A(n5733), .ZN(n5715) );
  NAND2_X1 U6255 ( .A1(n7329), .A2(n7328), .ZN(n7331) );
  NAND2_X1 U6256 ( .A1(n4651), .A2(n4649), .ZN(P2_U3548) );
  NAND2_X1 U6257 ( .A1(n4974), .A2(n4557), .ZN(n5371) );
  NAND2_X1 U6258 ( .A1(n5216), .A2(n5215), .ZN(n5220) );
  MUX2_X1 U6259 ( .A(n6294), .B(n6293), .S(n7351), .Z(n6296) );
  NAND2_X1 U6260 ( .A1(n5005), .A2(n6362), .ZN(n5004) );
  NAND2_X1 U6261 ( .A1(n4973), .A2(n4548), .ZN(n4972) );
  NAND2_X1 U6262 ( .A1(n5003), .A2(n5001), .ZN(n6369) );
  NAND2_X1 U6263 ( .A1(n5180), .A2(n5179), .ZN(n4658) );
  NAND2_X1 U6264 ( .A1(n6350), .A2(n9134), .ZN(n5008) );
  MUX2_X2 U6265 ( .A(n6271), .B(n6270), .S(n7351), .Z(n6291) );
  NAND2_X1 U6266 ( .A1(n5004), .A2(n6462), .ZN(n5003) );
  NAND2_X1 U6267 ( .A1(n4970), .A2(n6340), .ZN(n6360) );
  NAND2_X1 U6268 ( .A1(n5006), .A2(n6466), .ZN(n5005) );
  NAND2_X1 U6269 ( .A1(n6326), .A2(n4972), .ZN(n4971) );
  NOR3_X1 U6270 ( .A1(n6369), .A2(n6464), .A3(n6368), .ZN(n6492) );
  NAND2_X1 U6271 ( .A1(n6308), .A2(n9094), .ZN(n4973) );
  OAI21_X1 U6272 ( .B1(n5811), .B2(n5810), .A(n4553), .ZN(n5817) );
  AOI21_X1 U6273 ( .B1(n5736), .B2(n5735), .A(n4586), .ZN(n5742) );
  NAND2_X1 U6274 ( .A1(n4673), .A2(n4671), .ZN(n4670) );
  NAND2_X1 U6275 ( .A1(n4685), .A2(n5801), .ZN(n4684) );
  OAI21_X1 U6276 ( .B1(n5880), .B2(n5879), .A(n5878), .ZN(n5894) );
  INV_X1 U6277 ( .A(n7049), .ZN(n6572) );
  NAND2_X1 U6278 ( .A1(n4589), .A2(n4587), .ZN(n7049) );
  NAND2_X1 U6279 ( .A1(n4588), .A2(n8141), .ZN(n4587) );
  NAND2_X1 U6280 ( .A1(n8143), .A2(n8140), .ZN(n4588) );
  INV_X1 U6281 ( .A(n8143), .ZN(n4590) );
  NAND2_X1 U6282 ( .A1(n4593), .A2(n4594), .ZN(n6706) );
  NAND3_X1 U6283 ( .A1(n6676), .A2(n4595), .A3(n8978), .ZN(n4593) );
  NAND2_X1 U6284 ( .A1(n7568), .A2(n4603), .ZN(n4601) );
  NAND2_X1 U6285 ( .A1(n7959), .A2(n7958), .ZN(n7961) );
  NAND2_X1 U6286 ( .A1(n4611), .A2(n4858), .ZN(n4610) );
  NAND3_X1 U6287 ( .A1(n4509), .A2(n7028), .A3(n4844), .ZN(n4612) );
  NAND2_X1 U6288 ( .A1(n7032), .A2(n8222), .ZN(n4613) );
  NOR2_X1 U6289 ( .A1(n4620), .A2(n8189), .ZN(n8268) );
  NOR2_X1 U6290 ( .A1(n8213), .A2(n4621), .ZN(n4620) );
  NAND2_X1 U6291 ( .A1(n7293), .A2(n4500), .ZN(n4626) );
  NAND3_X1 U6292 ( .A1(n4626), .A2(n7512), .A3(n4625), .ZN(n7515) );
  INV_X2 U6293 ( .A(n5700), .ZN(n5104) );
  NAND2_X1 U6294 ( .A1(n7810), .A2(n4636), .ZN(n4634) );
  NAND2_X1 U6295 ( .A1(n4558), .A2(n4634), .ZN(n5347) );
  NAND3_X1 U6296 ( .A1(n4658), .A2(n4502), .A3(n5195), .ZN(n5216) );
  NAND2_X1 U6297 ( .A1(n5262), .A2(n4663), .ZN(n4659) );
  NAND2_X1 U6298 ( .A1(n4659), .A2(n4660), .ZN(n5307) );
  NAND3_X1 U6299 ( .A1(n4674), .A2(n4670), .A3(n8015), .ZN(n4669) );
  NAND3_X1 U6300 ( .A1(n4689), .A2(n5797), .A3(n4686), .ZN(n4685) );
  NAND3_X1 U6301 ( .A1(n5795), .A2(n5796), .A3(n8614), .ZN(n4689) );
  NAND3_X1 U6302 ( .A1(n5850), .A2(n5749), .A3(n4692), .ZN(n4691) );
  INV_X1 U6303 ( .A(n4698), .ZN(n4693) );
  NAND2_X1 U6304 ( .A1(n4693), .A2(n4967), .ZN(n4696) );
  NAND3_X1 U6305 ( .A1(n5151), .A2(n4696), .A3(n4694), .ZN(n5128) );
  NAND3_X1 U6306 ( .A1(n4698), .A2(n4697), .A3(n4559), .ZN(n5151) );
  NAND2_X1 U6307 ( .A1(n4490), .A2(n5104), .ZN(n5881) );
  NAND2_X1 U6308 ( .A1(n4490), .A2(n4701), .ZN(n4703) );
  NAND2_X1 U6309 ( .A1(n4704), .A2(n4705), .ZN(n6780) );
  INV_X1 U6310 ( .A(n4711), .ZN(n8988) );
  INV_X1 U6311 ( .A(n4723), .ZN(n8628) );
  XNOR2_X2 U6312 ( .A(n4724), .B(P1_IR_REG_19__SCAN_IN), .ZN(n10138) );
  AND2_X1 U6313 ( .A1(n8560), .A2(n4733), .ZN(n8532) );
  NAND2_X1 U6314 ( .A1(n8560), .A2(n4732), .ZN(n8519) );
  NAND2_X1 U6315 ( .A1(n8560), .A2(n8760), .ZN(n8549) );
  MUX2_X1 U6316 ( .A(n6859), .B(P1_REG2_REG_1__SCAN_IN), .S(n6939), .Z(n6942)
         );
  INV_X1 U6317 ( .A(n4749), .ZN(n9282) );
  OAI211_X2 U6318 ( .C1(n6798), .C2(n6062), .A(n5092), .B(n4750), .ZN(n6563)
         );
  NAND2_X2 U6319 ( .A1(n6117), .A2(n5917), .ZN(n6352) );
  OR2_X1 U6320 ( .A1(n4752), .A2(n4751), .ZN(n4750) );
  INV_X2 U6321 ( .A(n6117), .ZN(n4752) );
  INV_X1 U6322 ( .A(n4753), .ZN(n9182) );
  AND2_X1 U6323 ( .A1(n9175), .A2(n4764), .ZN(n9133) );
  NAND2_X1 U6324 ( .A1(n9175), .A2(n4763), .ZN(n9058) );
  NAND2_X1 U6325 ( .A1(n9175), .A2(n4766), .ZN(n9143) );
  NAND2_X1 U6326 ( .A1(n9175), .A2(n9162), .ZN(n9157) );
  NAND4_X1 U6327 ( .A1(n5910), .A2(n5071), .A3(n4885), .A4(n6472), .ZN(n4767)
         );
  NAND3_X1 U6328 ( .A1(n4780), .A2(n4778), .A3(n4777), .ZN(P2_U3264) );
  MUX2_X1 U6329 ( .A(n7228), .B(P2_REG2_REG_1__SCAN_IN), .S(n7107), .Z(n7104)
         );
  NAND2_X1 U6330 ( .A1(n4790), .A2(n7240), .ZN(n7386) );
  OAI21_X1 U6331 ( .B1(n10129), .B2(n10128), .A(n4790), .ZN(n10139) );
  NAND2_X1 U6332 ( .A1(n10128), .A2(n7239), .ZN(n4790) );
  NAND2_X1 U6333 ( .A1(n6565), .A2(n6027), .ZN(n6551) );
  NAND2_X1 U6334 ( .A1(n4791), .A2(n5071), .ZN(n6470) );
  NOR2_X2 U6335 ( .A1(n6470), .A2(n4497), .ZN(n5922) );
  NAND2_X1 U6336 ( .A1(n7858), .A2(n4795), .ZN(n4794) );
  AOI21_X1 U6337 ( .B1(n7624), .B2(n4800), .A(n7623), .ZN(n4798) );
  NAND3_X1 U6338 ( .A1(n10179), .A2(n4801), .A3(n7624), .ZN(n4799) );
  NAND2_X1 U6339 ( .A1(n9072), .A2(n4818), .ZN(n4815) );
  NAND2_X1 U6340 ( .A1(n4815), .A2(n4816), .ZN(n9318) );
  NAND2_X1 U6341 ( .A1(n9072), .A2(n9071), .ZN(n9347) );
  INV_X1 U6342 ( .A(n9194), .ZN(n4827) );
  NAND2_X1 U6343 ( .A1(n9194), .A2(n4838), .ZN(n4833) );
  NAND2_X1 U6344 ( .A1(n5922), .A2(n5921), .ZN(n5927) );
  INV_X1 U6345 ( .A(n5927), .ZN(n5924) );
  NAND2_X1 U6346 ( .A1(n4845), .A2(n4523), .ZN(n7145) );
  NAND2_X1 U6347 ( .A1(n4846), .A2(n4847), .ZN(n4845) );
  NAND2_X1 U6348 ( .A1(n7029), .A2(n4847), .ZN(n8221) );
  NAND2_X1 U6349 ( .A1(n6990), .A2(n6991), .ZN(n7029) );
  OR2_X1 U6350 ( .A1(n7361), .A2(n10283), .ZN(n5842) );
  NAND2_X1 U6351 ( .A1(n10283), .A2(n7361), .ZN(n5843) );
  OR2_X1 U6352 ( .A1(n4581), .A2(n5020), .ZN(n7330) );
  NOR2_X1 U6353 ( .A1(n7363), .A2(n4581), .ZN(n4853) );
  INV_X1 U6354 ( .A(n4581), .ZN(n4856) );
  NAND2_X1 U6355 ( .A1(n8266), .A2(n4873), .ZN(n8341) );
  NAND2_X1 U6356 ( .A1(n8330), .A2(n4877), .ZN(n4876) );
  OR2_X1 U6357 ( .A1(n4484), .A2(n6797), .ZN(n4889) );
  INV_X2 U6358 ( .A(n6553), .ZN(n10160) );
  NAND2_X2 U6359 ( .A1(n4888), .A2(n4889), .ZN(n6553) );
  NAND2_X1 U6360 ( .A1(n9195), .A2(n4891), .ZN(n4890) );
  OAI21_X1 U6361 ( .B1(n9195), .B2(n4896), .A(n4556), .ZN(n9163) );
  NAND2_X1 U6362 ( .A1(n4890), .A2(n4894), .ZN(n9149) );
  OAI21_X1 U6363 ( .B1(n9102), .B2(n4906), .A(n4904), .ZN(n9332) );
  OAI21_X1 U6364 ( .B1(n7847), .B2(n4914), .A(n4911), .ZN(n8033) );
  NAND2_X1 U6365 ( .A1(n9274), .A2(n4921), .ZN(n4920) );
  OAI21_X1 U6366 ( .B1(n7704), .B2(n4935), .A(n4931), .ZN(n7780) );
  OAI21_X1 U6367 ( .B1(n7704), .B2(n7526), .A(n7527), .ZN(n7528) );
  NAND2_X1 U6368 ( .A1(n7526), .A2(n7527), .ZN(n4936) );
  INV_X1 U6369 ( .A(n7445), .ZN(n5185) );
  NAND2_X1 U6370 ( .A1(n4937), .A2(n5710), .ZN(n7445) );
  NAND2_X1 U6371 ( .A1(n7412), .A2(n7413), .ZN(n4937) );
  NAND2_X1 U6372 ( .A1(n4938), .A2(n4940), .ZN(n5406) );
  NAND2_X1 U6373 ( .A1(n8014), .A2(n4941), .ZN(n4938) );
  NAND2_X1 U6374 ( .A1(n10250), .A2(n4946), .ZN(n4945) );
  AND2_X1 U6375 ( .A1(n5201), .A2(n5846), .ZN(n4946) );
  NAND2_X1 U6376 ( .A1(n8567), .A2(n4510), .ZN(n8542) );
  AND2_X1 U6377 ( .A1(n8567), .A2(n5808), .ZN(n8544) );
  NAND2_X1 U6378 ( .A1(n5510), .A2(n4566), .ZN(n5531) );
  NAND3_X1 U6379 ( .A1(n4971), .A2(n6338), .A3(n6339), .ZN(n4970) );
  NAND3_X1 U6380 ( .A1(n6297), .A2(n4977), .A3(n4976), .ZN(n6325) );
  NAND2_X1 U6381 ( .A1(n5453), .A2(n4983), .ZN(n4980) );
  NAND2_X1 U6382 ( .A1(n4980), .A2(n4981), .ZN(n5508) );
  NAND2_X1 U6383 ( .A1(n5453), .A2(n5452), .ZN(n5470) );
  NAND3_X1 U6384 ( .A1(n4985), .A2(n5468), .A3(n4984), .ZN(n4982) );
  INV_X1 U6385 ( .A(n4987), .ZN(n5449) );
  NAND2_X1 U6386 ( .A1(n5552), .A2(n5551), .ZN(n5562) );
  NAND3_X1 U6387 ( .A1(n5008), .A2(n5007), .A3(n4552), .ZN(n5006) );
  NAND2_X1 U6388 ( .A1(n7411), .A2(n7371), .ZN(n5013) );
  NAND2_X1 U6389 ( .A1(n5010), .A2(n5009), .ZN(n10243) );
  AOI21_X1 U6390 ( .B1(n7444), .B2(n5012), .A(n4547), .ZN(n5009) );
  NAND2_X1 U6391 ( .A1(n7410), .A2(n5011), .ZN(n5010) );
  INV_X1 U6392 ( .A(n5014), .ZN(n8627) );
  NAND2_X1 U6393 ( .A1(n8613), .A2(n5023), .ZN(n5022) );
  INV_X1 U6394 ( .A(n5024), .ZN(n8612) );
  NAND2_X1 U6395 ( .A1(n8727), .A2(n5028), .ZN(n5027) );
  INV_X1 U6396 ( .A(n5029), .ZN(n8726) );
  OAI21_X2 U6397 ( .B1(n8011), .B2(n5030), .A(n5032), .ZN(n8115) );
  INV_X1 U6398 ( .A(n5038), .ZN(n5037) );
  NAND2_X1 U6399 ( .A1(n5037), .A2(n5039), .ZN(n8012) );
  OR2_X1 U6400 ( .A1(n8009), .A2(n8373), .ZN(n5039) );
  NAND2_X1 U6401 ( .A1(n7594), .A2(n5042), .ZN(n5040) );
  NAND2_X1 U6402 ( .A1(n5040), .A2(n5041), .ZN(n7804) );
  NAND4_X1 U6403 ( .A1(n5045), .A2(n5044), .A3(n5163), .A4(n4543), .ZN(n5476)
         );
  INV_X1 U6404 ( .A(n8153), .ZN(n5955) );
  NAND2_X1 U6405 ( .A1(n8153), .A2(n9490), .ZN(n6032) );
  NAND2_X1 U6406 ( .A1(n8938), .A2(n6668), .ZN(n6675) );
  NAND2_X1 U6407 ( .A1(n8891), .A2(n4491), .ZN(n5061) );
  INV_X1 U6408 ( .A(n6716), .ZN(n5070) );
  OAI21_X1 U6409 ( .B1(n8068), .B2(n5074), .A(n5076), .ZN(n6648) );
  NAND2_X1 U6410 ( .A1(n8579), .A2(n8507), .ZN(n8558) );
  NAND2_X1 U6411 ( .A1(n8581), .A2(n8580), .ZN(n8579) );
  NOR2_X1 U6412 ( .A1(n8514), .A2(n8515), .ZN(n8513) );
  NAND2_X1 U6413 ( .A1(n8497), .A2(n8496), .ZN(n8727) );
  OAI21_X1 U6414 ( .B1(n8182), .B2(n8181), .A(n8258), .ZN(n8183) );
  XNOR2_X1 U6415 ( .A(n8185), .B(n8184), .ZN(n8213) );
  INV_X1 U6416 ( .A(n5552), .ZN(n5549) );
  OR2_X1 U6417 ( .A1(n5922), .A2(n5913), .ZN(n5914) );
  NAND2_X1 U6418 ( .A1(n6553), .A2(n6759), .ZN(n6554) );
  NAND2_X1 U6419 ( .A1(n7392), .A2(n6499), .ZN(n7312) );
  NAND2_X1 U6420 ( .A1(n8539), .A2(n8510), .ZN(n8531) );
  INV_X1 U6421 ( .A(n9416), .ZN(n9186) );
  NAND2_X1 U6422 ( .A1(n7312), .A2(n7313), .ZN(n7311) );
  OR2_X1 U6423 ( .A1(n5693), .A2(n4580), .ZN(n5144) );
  NAND2_X1 U6424 ( .A1(n9120), .A2(n6376), .ZN(n9188) );
  NAND2_X1 U6425 ( .A1(n5508), .A2(n5507), .ZN(n5510) );
  NAND2_X1 U6426 ( .A1(n8115), .A2(n8114), .ZN(n8497) );
  NAND2_X2 U6427 ( .A1(n6078), .A2(n6426), .ZN(n7704) );
  OR2_X1 U6428 ( .A1(n5693), .A2(n4584), .ZN(n5133) );
  AOI211_X1 U6429 ( .C1(n10125), .C2(n9397), .A(n9396), .B(n9395), .ZN(n9398)
         );
  OAI21_X1 U6430 ( .B1(n9132), .B2(n9356), .A(n9131), .ZN(n9395) );
  NOR2_X1 U6431 ( .A1(n6492), .A2(n6374), .ZN(n6490) );
  NAND2_X1 U6432 ( .A1(n6555), .A2(n6554), .ZN(n6556) );
  NOR2_X1 U6433 ( .A1(n9211), .A2(n9118), .ZN(n9196) );
  OR2_X1 U6434 ( .A1(n5893), .A2(n5892), .ZN(n5082) );
  INV_X1 U6435 ( .A(n8653), .ZN(n5519) );
  NAND2_X1 U6436 ( .A1(n5983), .A2(n5982), .ZN(n9198) );
  OR2_X1 U6437 ( .A1(n8183), .A2(n4560), .ZN(n5083) );
  OR2_X1 U6438 ( .A1(n8638), .A2(n8652), .ZN(n5084) );
  OR2_X1 U6439 ( .A1(n9261), .A2(n9082), .ZN(n5086) );
  AND2_X1 U6440 ( .A1(n6720), .A2(n6719), .ZN(n5088) );
  OR2_X1 U6441 ( .A1(n8682), .A2(n8502), .ZN(n5090) );
  AOI21_X1 U6442 ( .B1(n9145), .B2(n6346), .A(n6337), .ZN(n9096) );
  INV_X1 U6443 ( .A(n7716), .ZN(n5878) );
  OR2_X1 U6444 ( .A1(n6117), .A2(n6860), .ZN(n5092) );
  OR2_X1 U6445 ( .A1(n5142), .A2(n7107), .ZN(n5093) );
  AND2_X1 U6446 ( .A1(n5591), .A2(n5590), .ZN(n8572) );
  INV_X1 U6447 ( .A(n5595), .ZN(n5599) );
  INV_X1 U6448 ( .A(n8570), .ZN(n5615) );
  OR2_X1 U6449 ( .A1(n6493), .A2(n9203), .ZN(n5094) );
  INV_X1 U6450 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5904) );
  NOR2_X1 U6451 ( .A1(n8744), .A2(n8485), .ZN(n5706) );
  INV_X1 U6452 ( .A(n5380), .ZN(n5379) );
  INV_X1 U6453 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5909) );
  INV_X1 U6454 ( .A(n5538), .ZN(n5537) );
  INV_X1 U6455 ( .A(n5585), .ZN(n5584) );
  NAND2_X1 U6456 ( .A1(n5379), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5399) );
  AND2_X1 U6457 ( .A1(n5116), .A2(n5118), .ZN(n5105) );
  INV_X1 U6458 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5335) );
  OAI22_X1 U6459 ( .A1(n6544), .A2(n6727), .B1(n6542), .B2(n6733), .ZN(n6543)
         );
  INV_X1 U6460 ( .A(n5967), .ZN(n5952) );
  INV_X1 U6461 ( .A(n9096), .ZN(n9097) );
  AND2_X1 U6462 ( .A1(n6389), .A2(n8034), .ZN(n7994) );
  INV_X1 U6463 ( .A(n6376), .ZN(n9121) );
  INV_X1 U6464 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5923) );
  AND2_X1 U6465 ( .A1(n5369), .A2(n5368), .ZN(n5370) );
  INV_X1 U6466 ( .A(n5349), .ZN(n5350) );
  INV_X1 U6467 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5126) );
  INV_X1 U6468 ( .A(n5607), .ZN(n5605) );
  INV_X1 U6469 ( .A(n7504), .ZN(n7502) );
  NAND2_X1 U6470 ( .A1(n5497), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5513) );
  OR2_X1 U6471 ( .A1(n7361), .A2(n8243), .ZN(n7027) );
  NAND2_X1 U6472 ( .A1(n5537), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5556) );
  NAND2_X1 U6473 ( .A1(n8755), .A2(n8548), .ZN(n5819) );
  OR2_X1 U6474 ( .A1(n5556), .A2(n8214), .ZN(n5566) );
  NAND2_X1 U6475 ( .A1(n5185), .A2(n5184), .ZN(n10250) );
  INV_X1 U6476 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5095) );
  OR2_X1 U6477 ( .A1(n6332), .A2(n6331), .ZN(n6341) );
  AND2_X1 U6478 ( .A1(n5528), .A2(n5530), .ZN(n5529) );
  NAND2_X1 U6479 ( .A1(n5605), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5637) );
  OR2_X1 U6480 ( .A1(n5513), .A2(n8260), .ZN(n5538) );
  XNOR2_X1 U6481 ( .A(n8778), .B(n8156), .ZN(n8299) );
  NAND2_X1 U6482 ( .A1(n5873), .A2(n5872), .ZN(n5874) );
  INV_X1 U6483 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n7518) );
  INV_X1 U6484 ( .A(n8805), .ZN(n8682) );
  OR2_X1 U6485 ( .A1(n8840), .A2(n7926), .ZN(n5855) );
  OR2_X1 U6486 ( .A1(n5890), .A2(n7872), .ZN(n7058) );
  NAND2_X1 U6487 ( .A1(n7050), .A2(n6573), .ZN(n7194) );
  XNOR2_X1 U6488 ( .A(n6556), .B(n6712), .ZN(n8143) );
  AOI22_X1 U6489 ( .A1(n9421), .A2(n6608), .B1(n6565), .B2(n9091), .ZN(n6719)
         );
  INV_X1 U6490 ( .A(n7936), .ZN(n6618) );
  INV_X1 U6491 ( .A(n9405), .ZN(n9162) );
  AND2_X1 U6492 ( .A1(n9323), .A2(n9076), .ZN(n9077) );
  AND2_X1 U6493 ( .A1(n6435), .A2(n9106), .ZN(n9317) );
  INV_X1 U6494 ( .A(n7777), .ZN(n10199) );
  XNOR2_X1 U6495 ( .A(n5388), .B(n9667), .ZN(n5387) );
  AND2_X1 U6496 ( .A1(n5308), .A2(n5298), .ZN(n5306) );
  AND2_X1 U6497 ( .A1(n5614), .A2(n5613), .ZN(n8508) );
  AND4_X1 U6498 ( .A1(n5430), .A2(n5429), .A3(n5428), .A4(n5427), .ZN(n8289)
         );
  NAND2_X1 U6499 ( .A1(n5783), .A2(n8667), .ZN(n8676) );
  NAND2_X1 U6500 ( .A1(n7331), .A2(n7330), .ZN(n7368) );
  AND2_X1 U6501 ( .A1(n7058), .A2(n10275), .ZN(n10268) );
  INV_X1 U6502 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5457) );
  INV_X1 U6503 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5164) );
  INV_X1 U6504 ( .A(n9370), .ZN(n9238) );
  AND4_X1 U6505 ( .A1(n6000), .A2(n5999), .A3(n5998), .A4(n5997), .ZN(n9011)
         );
  AND2_X1 U6506 ( .A1(n6837), .A2(n9965), .ZN(n10117) );
  AND2_X1 U6507 ( .A1(n6450), .A2(n9119), .ZN(n9197) );
  AND2_X1 U6508 ( .A1(n6857), .A2(n6790), .ZN(n9368) );
  INV_X1 U6509 ( .A(n10145), .ZN(n9343) );
  OR2_X1 U6510 ( .A1(n6977), .A2(n7259), .ZN(n10207) );
  INV_X1 U6511 ( .A(n8481), .ZN(n10234) );
  INV_X1 U6512 ( .A(n8194), .ZN(n8760) );
  INV_X1 U6513 ( .A(n8024), .ZN(n8832) );
  INV_X1 U6514 ( .A(n8324), .ZN(n8366) );
  INV_X1 U6515 ( .A(n8572), .ZN(n8506) );
  INV_X1 U6516 ( .A(n7768), .ZN(n8375) );
  INV_X1 U6517 ( .A(n9897), .ZN(n10235) );
  AND2_X1 U6518 ( .A1(n8019), .A2(n8018), .ZN(n8837) );
  INV_X1 U6519 ( .A(n10360), .ZN(n10357) );
  INV_X1 U6520 ( .A(n10344), .ZN(n10342) );
  AND2_X1 U6521 ( .A1(n7017), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10275) );
  NAND2_X1 U6522 ( .A1(n6786), .A2(n6782), .ZN(n6783) );
  INV_X1 U6523 ( .A(n8962), .ZN(n9005) );
  INV_X1 U6524 ( .A(n9442), .ZN(n9261) );
  INV_X1 U6525 ( .A(n9093), .ZN(n9165) );
  AND2_X1 U6526 ( .A1(n8000), .A2(n7999), .ZN(n9943) );
  INV_X1 U6527 ( .A(n10231), .ZN(n10228) );
  AND2_X1 U6528 ( .A1(n9943), .A2(n9942), .ZN(n9957) );
  INV_X1 U6529 ( .A(n10217), .ZN(n10215) );
  INV_X1 U6530 ( .A(n10158), .ZN(n10154) );
  INV_X1 U6531 ( .A(n5954), .ZN(n9490) );
  INV_X1 U6532 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n9669) );
  INV_X1 U6533 ( .A(n8372), .ZN(P2_U3966) );
  AOI21_X1 U6534 ( .B1(n6536), .B2(n5094), .A(n6535), .ZN(P1_U3240) );
  NOR2_X1 U6535 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n5097) );
  INV_X1 U6536 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5102) );
  NOR3_X1 U6537 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .A3(
        P2_IR_REG_24__SCAN_IN), .ZN(n5103) );
  INV_X1 U6538 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5116) );
  INV_X1 U6539 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n8864) );
  NAND2_X1 U6540 ( .A1(n4536), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5107) );
  NAND2_X1 U6541 ( .A1(n5134), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5115) );
  NAND2_X1 U6542 ( .A1(n5169), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5114) );
  AND2_X2 U6543 ( .A1(n5111), .A2(n5110), .ZN(n5644) );
  NAND2_X1 U6544 ( .A1(n5644), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5113) );
  NAND2_X1 U6545 ( .A1(n5677), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5112) );
  INV_X1 U6547 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5162) );
  NOR2_X1 U6548 ( .A1(n5120), .A2(n5162), .ZN(n5121) );
  MUX2_X1 U6549 ( .A(n5162), .B(n5121), .S(P2_IR_REG_2__SCAN_IN), .Z(n5122) );
  INV_X1 U6550 ( .A(n5122), .ZN(n5124) );
  INV_X1 U6551 ( .A(n5163), .ZN(n5123) );
  NAND2_X1 U6552 ( .A1(n5124), .A2(n5123), .ZN(n7079) );
  NAND2_X4 U6553 ( .A1(n5142), .A2(n4483), .ZN(n5693) );
  NAND2_X2 U6554 ( .A1(n5142), .A2(n5917), .ZN(n5283) );
  INV_X1 U6555 ( .A(SI_1_), .ZN(n5127) );
  NAND2_X1 U6556 ( .A1(n5140), .A2(n5139), .ZN(n5130) );
  NAND2_X1 U6557 ( .A1(n5128), .A2(SI_1_), .ZN(n5129) );
  NAND2_X1 U6558 ( .A1(n5130), .A2(n5129), .ZN(n5157) );
  INV_X1 U6559 ( .A(SI_2_), .ZN(n5131) );
  XNOR2_X1 U6560 ( .A(n5158), .B(n5131), .ZN(n5156) );
  XNOR2_X1 U6561 ( .A(n5156), .B(n5157), .ZN(n6798) );
  OR2_X1 U6562 ( .A1(n5283), .A2(n6798), .ZN(n5132) );
  NAND2_X1 U6563 ( .A1(n8223), .A2(n7338), .ZN(n5721) );
  INV_X1 U6564 ( .A(n8223), .ZN(n8383) );
  NAND2_X1 U6565 ( .A1(n8383), .A2(n7034), .ZN(n5720) );
  NAND2_X1 U6566 ( .A1(n5134), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5138) );
  NAND2_X1 U6567 ( .A1(n5169), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5137) );
  NAND2_X1 U6568 ( .A1(n5644), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n5136) );
  XNOR2_X1 U6569 ( .A(n5139), .B(n5140), .ZN(n6797) );
  OR2_X1 U6570 ( .A1(n5283), .A2(n6797), .ZN(n5143) );
  INV_X1 U6571 ( .A(n5120), .ZN(n5141) );
  NAND2_X1 U6572 ( .A1(n5134), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5148) );
  NAND2_X1 U6573 ( .A1(n5169), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5147) );
  NAND2_X1 U6574 ( .A1(n5644), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5146) );
  INV_X2 U6575 ( .A(n5641), .ZN(n5677) );
  NAND2_X1 U6576 ( .A1(n5677), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5145) );
  NAND4_X1 U6577 ( .A1(n5148), .A2(n5147), .A3(n5146), .A4(n5145), .ZN(n8385)
         );
  INV_X1 U6578 ( .A(n8385), .ZN(n7012) );
  INV_X1 U6579 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5149) );
  OAI21_X1 U6580 ( .B1(n4483), .B2(n4968), .A(n5149), .ZN(n5150) );
  AND2_X1 U6581 ( .A1(n5151), .A2(n5150), .ZN(n8877) );
  MUX2_X1 U6582 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8877), .S(n5142), .Z(n7363) );
  NAND2_X1 U6583 ( .A1(n7012), .A2(n7363), .ZN(n7223) );
  NAND2_X1 U6584 ( .A1(n5843), .A2(n7223), .ZN(n5719) );
  NAND2_X1 U6585 ( .A1(n5719), .A2(n5842), .ZN(n7332) );
  NAND2_X1 U6586 ( .A1(n5134), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5155) );
  NAND2_X1 U6587 ( .A1(n5169), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5154) );
  INV_X1 U6588 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n9820) );
  NAND2_X1 U6589 ( .A1(n5644), .A2(n9820), .ZN(n5153) );
  NAND2_X1 U6590 ( .A1(n5677), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5152) );
  NAND4_X1 U6591 ( .A1(n5155), .A2(n5154), .A3(n5153), .A4(n5152), .ZN(n8382)
         );
  OR2_X1 U6592 ( .A1(n5693), .A2(n4632), .ZN(n5168) );
  NAND2_X1 U6593 ( .A1(n5157), .A2(n5156), .ZN(n5180) );
  NAND2_X1 U6594 ( .A1(n5158), .A2(SI_2_), .ZN(n5175) );
  NAND2_X1 U6595 ( .A1(n5180), .A2(n5175), .ZN(n5161) );
  INV_X1 U6596 ( .A(SI_3_), .ZN(n5160) );
  XNOR2_X1 U6597 ( .A(n5161), .B(n5177), .ZN(n6799) );
  OR2_X1 U6598 ( .A1(n5283), .A2(n6799), .ZN(n5167) );
  OR2_X1 U6599 ( .A1(n5163), .A2(n5162), .ZN(n5165) );
  XNOR2_X1 U6600 ( .A(n5165), .B(n5164), .ZN(n7120) );
  OR2_X1 U6601 ( .A1(n5142), .A2(n7120), .ZN(n5166) );
  XNOR2_X1 U6602 ( .A(n8382), .B(n10302), .ZN(n7371) );
  INV_X1 U6603 ( .A(n7371), .ZN(n7413) );
  INV_X1 U6604 ( .A(n8382), .ZN(n7372) );
  NAND2_X1 U6605 ( .A1(n7372), .A2(n8226), .ZN(n5710) );
  NAND2_X1 U6606 ( .A1(n5134), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5173) );
  NAND2_X1 U6607 ( .A1(n5676), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5172) );
  INV_X2 U6608 ( .A(n5609), .ZN(n5660) );
  XNOR2_X1 U6609 ( .A(n9820), .B(P2_REG3_REG_4__SCAN_IN), .ZN(n7443) );
  NAND2_X1 U6610 ( .A1(n5660), .A2(n7443), .ZN(n5171) );
  NAND2_X1 U6611 ( .A1(n5677), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5170) );
  OR2_X1 U6612 ( .A1(n5455), .A2(n5162), .ZN(n5174) );
  INV_X1 U6613 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5194) );
  XNOR2_X1 U6614 ( .A(n5174), .B(n5194), .ZN(n7135) );
  INV_X1 U6615 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6802) );
  OR2_X1 U6616 ( .A1(n5693), .A2(n6802), .ZN(n5183) );
  AND2_X1 U6617 ( .A1(n5175), .A2(n5176), .ZN(n5179) );
  INV_X1 U6618 ( .A(n5176), .ZN(n5178) );
  MUX2_X1 U6619 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n4483), .Z(n5197) );
  OR2_X1 U6620 ( .A1(n5283), .A2(n6805), .ZN(n5182) );
  NAND2_X1 U6621 ( .A1(n7414), .A2(n10244), .ZN(n5711) );
  INV_X1 U6622 ( .A(n7414), .ZN(n8381) );
  NAND2_X1 U6623 ( .A1(n5134), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5193) );
  NAND2_X1 U6624 ( .A1(n5676), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5192) );
  INV_X1 U6625 ( .A(n5186), .ZN(n5188) );
  INV_X1 U6626 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5187) );
  NAND2_X1 U6627 ( .A1(n5188), .A2(n5187), .ZN(n5189) );
  AND2_X1 U6628 ( .A1(n5203), .A2(n5189), .ZN(n10256) );
  NAND2_X1 U6629 ( .A1(n5644), .A2(n10256), .ZN(n5191) );
  NAND2_X1 U6630 ( .A1(n5677), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5190) );
  NAND4_X1 U6631 ( .A1(n5193), .A2(n5192), .A3(n5191), .A4(n5190), .ZN(n8380)
         );
  INV_X1 U6632 ( .A(n8380), .ZN(n7301) );
  NAND2_X1 U6633 ( .A1(n5455), .A2(n5194), .ZN(n5254) );
  NAND2_X1 U6634 ( .A1(n5254), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5209) );
  XNOR2_X1 U6635 ( .A(n5209), .B(P2_IR_REG_5__SCAN_IN), .ZN(n7083) );
  INV_X1 U6636 ( .A(n7083), .ZN(n7179) );
  NAND2_X1 U6637 ( .A1(n5197), .A2(SI_4_), .ZN(n5214) );
  NAND2_X1 U6638 ( .A1(n5216), .A2(n5214), .ZN(n5198) );
  MUX2_X1 U6639 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n4482), .Z(n5213) );
  XNOR2_X1 U6640 ( .A(n5198), .B(n5218), .ZN(n6809) );
  OR2_X1 U6641 ( .A1(n5283), .A2(n6809), .ZN(n5200) );
  INV_X1 U6642 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6804) );
  OR2_X1 U6643 ( .A1(n5693), .A2(n6804), .ZN(n5199) );
  OAI211_X1 U6644 ( .C1(n5142), .C2(n7179), .A(n5200), .B(n5199), .ZN(n10259)
         );
  NAND2_X1 U6645 ( .A1(n8380), .A2(n10317), .ZN(n5731) );
  NAND2_X1 U6646 ( .A1(n5712), .A2(n5731), .ZN(n10251) );
  INV_X1 U6647 ( .A(n10249), .ZN(n5730) );
  NOR2_X1 U6648 ( .A1(n10251), .A2(n5730), .ZN(n5201) );
  NAND2_X1 U6649 ( .A1(n5134), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5208) );
  NAND2_X1 U6650 ( .A1(n5676), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5207) );
  INV_X1 U6651 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n9610) );
  NAND2_X1 U6652 ( .A1(n5203), .A2(n9610), .ZN(n5204) );
  AND2_X1 U6653 ( .A1(n5226), .A2(n5204), .ZN(n7303) );
  NAND2_X1 U6654 ( .A1(n5660), .A2(n7303), .ZN(n5206) );
  NAND2_X1 U6655 ( .A1(n5677), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5205) );
  NAND2_X1 U6656 ( .A1(n5209), .A2(n5251), .ZN(n5210) );
  NAND2_X1 U6657 ( .A1(n5210), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5211) );
  NAND2_X1 U6658 ( .A1(n5211), .A2(n5252), .ZN(n5236) );
  OR2_X1 U6659 ( .A1(n5211), .A2(n5252), .ZN(n5212) );
  NAND2_X1 U6660 ( .A1(n5236), .A2(n5212), .ZN(n7191) );
  NAND2_X1 U6661 ( .A1(n5213), .A2(SI_5_), .ZN(n5217) );
  AND2_X1 U6662 ( .A1(n5214), .A2(n5217), .ZN(n5215) );
  MUX2_X1 U6663 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n4483), .Z(n5234) );
  INV_X1 U6664 ( .A(SI_6_), .ZN(n5221) );
  XNOR2_X1 U6665 ( .A(n5233), .B(n5232), .ZN(n6807) );
  OR2_X1 U6666 ( .A1(n5283), .A2(n6807), .ZN(n5223) );
  INV_X1 U6667 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6803) );
  OR2_X1 U6668 ( .A1(n5693), .A2(n6803), .ZN(n5222) );
  NAND2_X1 U6669 ( .A1(n7458), .A2(n7453), .ZN(n5737) );
  INV_X1 U6670 ( .A(n7458), .ZN(n8379) );
  INV_X1 U6671 ( .A(n7453), .ZN(n7382) );
  NAND2_X1 U6672 ( .A1(n8379), .A2(n7382), .ZN(n5735) );
  NAND2_X1 U6673 ( .A1(n5737), .A2(n5735), .ZN(n7455) );
  INV_X1 U6674 ( .A(n7455), .ZN(n5846) );
  INV_X1 U6675 ( .A(n7457), .ZN(n5242) );
  NAND2_X1 U6676 ( .A1(n5675), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5231) );
  NAND2_X1 U6677 ( .A1(n5676), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5230) );
  INV_X1 U6678 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5225) );
  NAND2_X1 U6679 ( .A1(n5226), .A2(n5225), .ZN(n5227) );
  AND2_X1 U6680 ( .A1(n5244), .A2(n5227), .ZN(n7581) );
  NAND2_X1 U6681 ( .A1(n5660), .A2(n7581), .ZN(n5229) );
  NAND2_X1 U6682 ( .A1(n5677), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5228) );
  NAND4_X1 U6683 ( .A1(n5231), .A2(n5230), .A3(n5229), .A4(n5228), .ZN(n8378)
         );
  NAND2_X1 U6684 ( .A1(n5234), .A2(SI_6_), .ZN(n5235) );
  MUX2_X1 U6685 ( .A(n6801), .B(n9657), .S(n4483), .Z(n5259) );
  XNOR2_X1 U6686 ( .A(n5258), .B(n5257), .ZN(n6800) );
  OR2_X1 U6687 ( .A1(n5283), .A2(n6800), .ZN(n5240) );
  OR2_X1 U6688 ( .A1(n5693), .A2(n6801), .ZN(n5239) );
  NAND2_X1 U6689 ( .A1(n5236), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5237) );
  XNOR2_X1 U6690 ( .A(n5237), .B(P2_IR_REG_7__SCAN_IN), .ZN(n7088) );
  INV_X1 U6691 ( .A(n7088), .ZN(n7167) );
  OR2_X1 U6692 ( .A1(n5142), .A2(n7167), .ZN(n5238) );
  XNOR2_X1 U6693 ( .A(n8378), .B(n7591), .ZN(n7589) );
  NAND2_X1 U6694 ( .A1(n8378), .A2(n7591), .ZN(n5243) );
  NAND2_X1 U6695 ( .A1(n5675), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5249) );
  NAND2_X1 U6696 ( .A1(n5676), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5248) );
  NAND2_X1 U6697 ( .A1(n5244), .A2(n7518), .ZN(n5245) );
  AND2_X1 U6698 ( .A1(n5269), .A2(n5245), .ZN(n7608) );
  NAND2_X1 U6699 ( .A1(n5660), .A2(n7608), .ZN(n5247) );
  NAND2_X1 U6700 ( .A1(n5677), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5246) );
  NAND4_X1 U6701 ( .A1(n5249), .A2(n5248), .A3(n5247), .A4(n5246), .ZN(n8377)
         );
  INV_X1 U6702 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5250) );
  NAND3_X1 U6703 ( .A1(n5252), .A2(n5251), .A3(n5250), .ZN(n5253) );
  OR2_X1 U6704 ( .A1(n5254), .A2(n5253), .ZN(n5275) );
  NAND2_X1 U6705 ( .A1(n5275), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5256) );
  INV_X1 U6706 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5255) );
  XNOR2_X1 U6707 ( .A(n5256), .B(n5255), .ZN(n7281) );
  OR2_X1 U6708 ( .A1(n5693), .A2(n6812), .ZN(n5267) );
  INV_X1 U6709 ( .A(n5259), .ZN(n5260) );
  MUX2_X1 U6710 ( .A(n6812), .B(n9833), .S(n4483), .Z(n5263) );
  INV_X1 U6711 ( .A(n5263), .ZN(n5264) );
  NAND2_X1 U6712 ( .A1(n5264), .A2(SI_8_), .ZN(n5265) );
  OR2_X1 U6713 ( .A1(n5283), .A2(n6811), .ZN(n5266) );
  INV_X1 U6714 ( .A(n8377), .ZN(n7459) );
  NAND2_X1 U6715 ( .A1(n5676), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5274) );
  NAND2_X1 U6716 ( .A1(n5675), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5273) );
  INV_X1 U6717 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5268) );
  NAND2_X1 U6718 ( .A1(n5269), .A2(n5268), .ZN(n5270) );
  NAND2_X1 U6719 ( .A1(n5287), .A2(n5270), .ZN(n7688) );
  INV_X1 U6720 ( .A(n7688), .ZN(n7735) );
  NAND2_X1 U6721 ( .A1(n5660), .A2(n7735), .ZN(n5272) );
  NAND2_X1 U6722 ( .A1(n5677), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5271) );
  INV_X1 U6723 ( .A(n7807), .ZN(n8376) );
  NOR2_X1 U6724 ( .A1(n5275), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n5337) );
  OR2_X1 U6725 ( .A1(n5337), .A2(n5162), .ZN(n5299) );
  XNOR2_X1 U6726 ( .A(n5299), .B(P2_IR_REG_9__SCAN_IN), .ZN(n8391) );
  AOI22_X1 U6727 ( .A1(n5669), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6825), .B2(
        n8391), .ZN(n5285) );
  INV_X1 U6728 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6818) );
  MUX2_X1 U6729 ( .A(n6818), .B(n9806), .S(n4483), .Z(n5280) );
  INV_X1 U6730 ( .A(SI_9_), .ZN(n5279) );
  INV_X1 U6731 ( .A(n5280), .ZN(n5281) );
  NAND2_X1 U6732 ( .A1(n5281), .A2(SI_9_), .ZN(n5282) );
  XNOR2_X1 U6733 ( .A(n5294), .B(n5293), .ZN(n6817) );
  NAND2_X1 U6734 ( .A1(n6817), .A2(n5692), .ZN(n5284) );
  INV_X1 U6735 ( .A(n7839), .ZN(n7761) );
  NAND2_X1 U6736 ( .A1(n8376), .A2(n7761), .ZN(n5850) );
  NAND2_X1 U6737 ( .A1(n7683), .A2(n5850), .ZN(n7810) );
  NAND2_X1 U6738 ( .A1(n5675), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5292) );
  NAND2_X1 U6739 ( .A1(n5676), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5291) );
  INV_X1 U6740 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n7652) );
  NAND2_X1 U6741 ( .A1(n5287), .A2(n7652), .ZN(n5288) );
  AND2_X1 U6742 ( .A1(n5318), .A2(n5288), .ZN(n7653) );
  NAND2_X1 U6743 ( .A1(n5660), .A2(n7653), .ZN(n5290) );
  NAND2_X1 U6744 ( .A1(n5677), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5289) );
  INV_X1 U6745 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6823) );
  MUX2_X1 U6746 ( .A(n6823), .B(n9669), .S(n4483), .Z(n5296) );
  INV_X1 U6747 ( .A(SI_10_), .ZN(n9795) );
  INV_X1 U6748 ( .A(n5296), .ZN(n5297) );
  NAND2_X1 U6749 ( .A1(n5297), .A2(SI_10_), .ZN(n5298) );
  XNOR2_X1 U6750 ( .A(n5307), .B(n5306), .ZN(n6822) );
  NAND2_X1 U6751 ( .A1(n6822), .A2(n5692), .ZN(n5302) );
  NAND2_X1 U6752 ( .A1(n5299), .A2(n5335), .ZN(n5300) );
  NAND2_X1 U6753 ( .A1(n5300), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5311) );
  XNOR2_X1 U6754 ( .A(n5311), .B(P2_IR_REG_10__SCAN_IN), .ZN(n7484) );
  AOI22_X1 U6755 ( .A1(n5669), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6825), .B2(
        n7484), .ZN(n5301) );
  NAND2_X1 U6756 ( .A1(n5302), .A2(n5301), .ZN(n7823) );
  NAND2_X1 U6757 ( .A1(n7768), .A2(n7823), .ZN(n5748) );
  INV_X1 U6758 ( .A(n7812), .ZN(n5304) );
  NAND2_X1 U6759 ( .A1(n7807), .A2(n7839), .ZN(n7809) );
  INV_X1 U6760 ( .A(n7809), .ZN(n5303) );
  NOR2_X1 U6761 ( .A1(n5304), .A2(n5303), .ZN(n5305) );
  NAND2_X1 U6762 ( .A1(n5307), .A2(n5306), .ZN(n5309) );
  NAND2_X1 U6763 ( .A1(n5309), .A2(n5308), .ZN(n5325) );
  INV_X1 U6764 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n5310) );
  INV_X1 U6765 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6831) );
  MUX2_X1 U6766 ( .A(n5310), .B(n6831), .S(n4483), .Z(n5326) );
  XNOR2_X1 U6767 ( .A(n5325), .B(n5324), .ZN(n6820) );
  NAND2_X1 U6768 ( .A1(n6820), .A2(n5692), .ZN(n5315) );
  INV_X1 U6769 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5334) );
  NAND2_X1 U6770 ( .A1(n5311), .A2(n5334), .ZN(n5312) );
  NAND2_X1 U6771 ( .A1(n5312), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5313) );
  XNOR2_X1 U6772 ( .A(n5313), .B(P2_IR_REG_11__SCAN_IN), .ZN(n8407) );
  AOI22_X1 U6773 ( .A1(n5669), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6825), .B2(
        n8407), .ZN(n5314) );
  NAND2_X1 U6774 ( .A1(n5676), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5323) );
  NAND2_X1 U6775 ( .A1(n5677), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n5322) );
  INV_X1 U6776 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n5317) );
  NAND2_X1 U6777 ( .A1(n5318), .A2(n5317), .ZN(n5319) );
  AND2_X1 U6778 ( .A1(n5341), .A2(n5319), .ZN(n7756) );
  NAND2_X1 U6779 ( .A1(n5660), .A2(n7756), .ZN(n5321) );
  NAND2_X1 U6780 ( .A1(n5675), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5320) );
  NAND2_X1 U6781 ( .A1(n8840), .A2(n7926), .ZN(n5854) );
  INV_X1 U6782 ( .A(n5326), .ZN(n5327) );
  INV_X1 U6783 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n5329) );
  INV_X1 U6784 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6869) );
  MUX2_X1 U6785 ( .A(n5329), .B(n6869), .S(n4483), .Z(n5330) );
  INV_X1 U6786 ( .A(SI_12_), .ZN(n9644) );
  INV_X1 U6787 ( .A(n5330), .ZN(n5331) );
  NAND2_X1 U6788 ( .A1(n5331), .A2(SI_12_), .ZN(n5332) );
  XNOR2_X1 U6789 ( .A(n5348), .B(n5349), .ZN(n6844) );
  NAND2_X1 U6790 ( .A1(n6844), .A2(n5692), .ZN(n5340) );
  INV_X1 U6791 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5333) );
  AND3_X1 U6792 ( .A1(n5335), .A2(n5334), .A3(n5333), .ZN(n5336) );
  AND2_X1 U6793 ( .A1(n5337), .A2(n5336), .ZN(n5357) );
  OR2_X1 U6794 ( .A1(n5357), .A2(n5162), .ZN(n5338) );
  XNOR2_X1 U6795 ( .A(n5338), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7672) );
  AOI22_X1 U6796 ( .A1(n5669), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6825), .B2(
        n7672), .ZN(n5339) );
  NAND2_X1 U6797 ( .A1(n5675), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5346) );
  NAND2_X1 U6798 ( .A1(n5676), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5345) );
  INV_X1 U6799 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n9821) );
  NAND2_X1 U6800 ( .A1(n5341), .A2(n9821), .ZN(n5342) );
  AND2_X1 U6801 ( .A1(n5362), .A2(n5342), .ZN(n7930) );
  NAND2_X1 U6802 ( .A1(n5660), .A2(n7930), .ZN(n5344) );
  NAND2_X1 U6803 ( .A1(n5677), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5343) );
  NAND2_X1 U6804 ( .A1(n8009), .A2(n8008), .ZN(n5852) );
  NAND2_X1 U6805 ( .A1(n5347), .A2(n5852), .ZN(n8014) );
  NAND2_X1 U6806 ( .A1(n5371), .A2(n5369), .ZN(n5355) );
  INV_X1 U6807 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6894) );
  INV_X1 U6808 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n6892) );
  MUX2_X1 U6809 ( .A(n6894), .B(n6892), .S(n4483), .Z(n5352) );
  INV_X1 U6810 ( .A(SI_13_), .ZN(n5351) );
  NAND2_X1 U6811 ( .A1(n5352), .A2(n5351), .ZN(n5368) );
  INV_X1 U6812 ( .A(n5352), .ZN(n5353) );
  NAND2_X1 U6813 ( .A1(n5353), .A2(SI_13_), .ZN(n5372) );
  AND2_X1 U6814 ( .A1(n5368), .A2(n5372), .ZN(n5354) );
  XNOR2_X1 U6815 ( .A(n5355), .B(n5354), .ZN(n6891) );
  NAND2_X1 U6816 ( .A1(n6891), .A2(n5692), .ZN(n5359) );
  INV_X1 U6817 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5356) );
  NAND2_X1 U6818 ( .A1(n5357), .A2(n5356), .ZN(n5418) );
  NAND2_X1 U6819 ( .A1(n5418), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5373) );
  XNOR2_X1 U6820 ( .A(n5373), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7726) );
  AOI22_X1 U6821 ( .A1(n5669), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6825), .B2(
        n7726), .ZN(n5358) );
  NAND2_X1 U6822 ( .A1(n5134), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5367) );
  NAND2_X1 U6823 ( .A1(n5676), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n5366) );
  INV_X1 U6824 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5361) );
  NAND2_X1 U6825 ( .A1(n5362), .A2(n5361), .ZN(n5363) );
  AND2_X1 U6826 ( .A1(n5380), .A2(n5363), .ZN(n8023) );
  NAND2_X1 U6827 ( .A1(n5660), .A2(n8023), .ZN(n5365) );
  NAND2_X1 U6828 ( .A1(n5677), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5364) );
  OR2_X1 U6829 ( .A1(n8024), .A2(n8370), .ZN(n5756) );
  NAND2_X1 U6830 ( .A1(n8024), .A2(n8370), .ZN(n8049) );
  MUX2_X1 U6831 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n4483), .Z(n5388) );
  INV_X1 U6832 ( .A(SI_14_), .ZN(n9667) );
  XNOR2_X1 U6833 ( .A(n5391), .B(n5387), .ZN(n6916) );
  NAND2_X1 U6834 ( .A1(n6916), .A2(n5692), .ZN(n5378) );
  INV_X1 U6835 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5416) );
  NAND2_X1 U6836 ( .A1(n5373), .A2(n5416), .ZN(n5374) );
  NAND2_X1 U6837 ( .A1(n5374), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5375) );
  INV_X1 U6838 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5415) );
  NAND2_X1 U6839 ( .A1(n5375), .A2(n5415), .ZN(n5395) );
  OR2_X1 U6840 ( .A1(n5375), .A2(n5415), .ZN(n5376) );
  AND2_X1 U6841 ( .A1(n5395), .A2(n5376), .ZN(n7972) );
  AOI22_X1 U6842 ( .A1(n5669), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6825), .B2(
        n7972), .ZN(n5377) );
  NAND2_X1 U6843 ( .A1(n5675), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5385) );
  NAND2_X1 U6844 ( .A1(n5676), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n5384) );
  INV_X1 U6845 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n9839) );
  NAND2_X1 U6846 ( .A1(n5380), .A2(n9839), .ZN(n5381) );
  AND2_X1 U6847 ( .A1(n5399), .A2(n5381), .ZN(n8092) );
  NAND2_X1 U6848 ( .A1(n5660), .A2(n8092), .ZN(n5383) );
  NAND2_X1 U6849 ( .A1(n5677), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n5382) );
  NAND2_X1 U6850 ( .A1(n8111), .A2(n8110), .ZN(n5760) );
  INV_X1 U6851 ( .A(n8112), .ZN(n8051) );
  INV_X1 U6852 ( .A(n8049), .ZN(n5758) );
  NOR2_X1 U6853 ( .A1(n8051), .A2(n5758), .ZN(n5386) );
  NAND2_X1 U6854 ( .A1(n5388), .A2(SI_14_), .ZN(n5389) );
  INV_X1 U6855 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7041) );
  INV_X1 U6856 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n9584) );
  MUX2_X1 U6857 ( .A(n7041), .B(n9584), .S(n4483), .Z(n5392) );
  INV_X1 U6858 ( .A(SI_15_), .ZN(n9823) );
  NAND2_X1 U6859 ( .A1(n5392), .A2(n9823), .ZN(n5407) );
  INV_X1 U6860 ( .A(n5392), .ZN(n5393) );
  NAND2_X1 U6861 ( .A1(n5393), .A2(SI_15_), .ZN(n5394) );
  NAND2_X1 U6862 ( .A1(n5407), .A2(n5394), .ZN(n5408) );
  XNOR2_X1 U6863 ( .A(n5409), .B(n5408), .ZN(n7039) );
  NAND2_X1 U6864 ( .A1(n7039), .A2(n5692), .ZN(n5398) );
  NAND2_X1 U6865 ( .A1(n5395), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5396) );
  XNOR2_X1 U6866 ( .A(n5396), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8416) );
  AOI22_X1 U6867 ( .A1(n5669), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n6825), .B2(
        n8416), .ZN(n5397) );
  NAND2_X1 U6868 ( .A1(n5675), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5404) );
  NAND2_X1 U6869 ( .A1(n5676), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n5403) );
  INV_X1 U6870 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n8358) );
  NAND2_X1 U6871 ( .A1(n5399), .A2(n8358), .ZN(n5400) );
  AND2_X1 U6872 ( .A1(n5425), .A2(n5400), .ZN(n8116) );
  NAND2_X1 U6873 ( .A1(n5644), .A2(n8116), .ZN(n5402) );
  NAND2_X1 U6874 ( .A1(n5677), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n5401) );
  OR2_X1 U6875 ( .A1(n8495), .A2(n8281), .ZN(n5405) );
  NAND2_X1 U6876 ( .A1(n5406), .A2(n5405), .ZN(n8736) );
  INV_X1 U6877 ( .A(n8736), .ZN(n5431) );
  INV_X1 U6878 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n5410) );
  INV_X1 U6879 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n9849) );
  MUX2_X1 U6880 ( .A(n5410), .B(n9849), .S(n4483), .Z(n5411) );
  INV_X1 U6881 ( .A(SI_16_), .ZN(n9658) );
  NAND2_X1 U6882 ( .A1(n5411), .A2(n9658), .ZN(n5435) );
  INV_X1 U6883 ( .A(n5411), .ZN(n5412) );
  NAND2_X1 U6884 ( .A1(n5412), .A2(SI_16_), .ZN(n5413) );
  XNOR2_X1 U6885 ( .A(n5434), .B(n5433), .ZN(n7136) );
  NAND2_X1 U6886 ( .A1(n7136), .A2(n5692), .ZN(n5423) );
  INV_X1 U6887 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5414) );
  NAND3_X1 U6888 ( .A1(n5416), .A2(n5415), .A3(n5414), .ZN(n5417) );
  OAI21_X1 U6889 ( .B1(n5418), .B2(n5417), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n5419) );
  MUX2_X1 U6890 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5419), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n5421) );
  NAND2_X1 U6891 ( .A1(n5455), .A2(n5420), .ZN(n5437) );
  AND2_X1 U6892 ( .A1(n5421), .A2(n5437), .ZN(n8437) );
  AOI22_X1 U6893 ( .A1(n5669), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6825), .B2(
        n8437), .ZN(n5422) );
  NAND2_X1 U6894 ( .A1(n5675), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5430) );
  NAND2_X1 U6895 ( .A1(n5676), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n5429) );
  INV_X1 U6896 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n9860) );
  NAND2_X1 U6897 ( .A1(n5425), .A2(n9860), .ZN(n5426) );
  AND2_X1 U6898 ( .A1(n5442), .A2(n5426), .ZN(n8731) );
  NAND2_X1 U6899 ( .A1(n5660), .A2(n8731), .ZN(n5428) );
  NAND2_X1 U6900 ( .A1(n5677), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n5427) );
  NAND2_X1 U6901 ( .A1(n8820), .A2(n8289), .ZN(n5767) );
  MUX2_X1 U6902 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .S(n4483), .Z(n5451) );
  INV_X1 U6903 ( .A(SI_17_), .ZN(n5436) );
  XNOR2_X1 U6904 ( .A(n5451), .B(n5436), .ZN(n5450) );
  XNOR2_X1 U6905 ( .A(n5449), .B(n5450), .ZN(n7201) );
  NAND2_X1 U6906 ( .A1(n7201), .A2(n5692), .ZN(n5440) );
  NAND2_X1 U6907 ( .A1(n5437), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5438) );
  XNOR2_X1 U6908 ( .A(n5438), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8448) );
  AOI22_X1 U6909 ( .A1(n5669), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6825), .B2(
        n8448), .ZN(n5439) );
  NAND2_X1 U6910 ( .A1(n5675), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5447) );
  NAND2_X1 U6911 ( .A1(n5676), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n5446) );
  INV_X1 U6912 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n5441) );
  NAND2_X1 U6913 ( .A1(n5442), .A2(n5441), .ZN(n5443) );
  AND2_X1 U6914 ( .A1(n5462), .A2(n5443), .ZN(n8720) );
  NAND2_X1 U6915 ( .A1(n5660), .A2(n8720), .ZN(n5445) );
  NAND2_X1 U6916 ( .A1(n5677), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n5444) );
  NAND4_X1 U6917 ( .A1(n5447), .A2(n5446), .A3(n5445), .A4(n5444), .ZN(n8701)
         );
  NAND2_X1 U6918 ( .A1(n8816), .A2(n8701), .ZN(n5448) );
  INV_X1 U6919 ( .A(n8701), .ZN(n5771) );
  OR2_X1 U6920 ( .A1(n8816), .A2(n5771), .ZN(n5772) );
  NAND2_X1 U6921 ( .A1(n4987), .A2(n5450), .ZN(n5453) );
  NAND2_X1 U6922 ( .A1(n5451), .A2(SI_17_), .ZN(n5452) );
  MUX2_X1 U6923 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n4483), .Z(n5471) );
  XNOR2_X1 U6924 ( .A(n5471), .B(SI_18_), .ZN(n5468) );
  NAND2_X1 U6925 ( .A1(n7234), .A2(n5692), .ZN(n5460) );
  NAND2_X1 U6926 ( .A1(n5455), .A2(n5454), .ZN(n5456) );
  NAND2_X1 U6927 ( .A1(n5456), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5458) );
  XNOR2_X1 U6928 ( .A(n5458), .B(n5457), .ZN(n8472) );
  INV_X1 U6929 ( .A(n8472), .ZN(n8457) );
  AOI22_X1 U6930 ( .A1(n5669), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6825), .B2(
        n8457), .ZN(n5459) );
  NAND2_X1 U6931 ( .A1(n5675), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n5467) );
  NAND2_X1 U6932 ( .A1(n5676), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n5466) );
  INV_X1 U6933 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n9804) );
  NAND2_X1 U6934 ( .A1(n5462), .A2(n9804), .ZN(n5463) );
  AND2_X1 U6935 ( .A1(n5482), .A2(n5463), .ZN(n8695) );
  NAND2_X1 U6936 ( .A1(n5644), .A2(n8695), .ZN(n5465) );
  NAND2_X1 U6937 ( .A1(n5677), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n5464) );
  NAND4_X1 U6938 ( .A1(n5467), .A2(n5466), .A3(n5465), .A4(n5464), .ZN(n8685)
         );
  INV_X1 U6939 ( .A(n8685), .ZN(n8500) );
  NAND2_X1 U6940 ( .A1(n8809), .A2(n8500), .ZN(n5785) );
  AND2_X1 U6941 ( .A1(n8697), .A2(n8685), .ZN(n5841) );
  INV_X1 U6942 ( .A(n5468), .ZN(n5469) );
  INV_X1 U6943 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7327) );
  INV_X1 U6944 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n9796) );
  MUX2_X1 U6945 ( .A(n7327), .B(n9796), .S(n4483), .Z(n5473) );
  INV_X1 U6946 ( .A(SI_19_), .ZN(n5472) );
  NAND2_X1 U6947 ( .A1(n5473), .A2(n5472), .ZN(n5488) );
  INV_X1 U6948 ( .A(n5473), .ZN(n5474) );
  NAND2_X1 U6949 ( .A1(n5474), .A2(SI_19_), .ZN(n5475) );
  NAND2_X1 U6950 ( .A1(n5488), .A2(n5475), .ZN(n5489) );
  XNOR2_X1 U6951 ( .A(n5490), .B(n5489), .ZN(n7325) );
  NAND2_X1 U6952 ( .A1(n7325), .A2(n5692), .ZN(n5480) );
  NAND2_X1 U6953 ( .A1(n5476), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5478) );
  INV_X1 U6954 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5477) );
  XNOR2_X1 U6955 ( .A(n5478), .B(n5477), .ZN(n8478) );
  AOI22_X1 U6956 ( .A1(n5669), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n4781), .B2(
        n6825), .ZN(n5479) );
  NAND2_X1 U6957 ( .A1(n5675), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5487) );
  NAND2_X1 U6958 ( .A1(n5676), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n5486) );
  INV_X1 U6959 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n5481) );
  OR2_X2 U6960 ( .A1(n5482), .A2(n5481), .ZN(n5499) );
  NAND2_X1 U6961 ( .A1(n5482), .A2(n5481), .ZN(n5483) );
  AND2_X1 U6962 ( .A1(n5499), .A2(n5483), .ZN(n8680) );
  NAND2_X1 U6963 ( .A1(n5660), .A2(n8680), .ZN(n5485) );
  NAND2_X1 U6964 ( .A1(n5677), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n5484) );
  NAND2_X1 U6965 ( .A1(n8805), .A2(n8502), .ZN(n8667) );
  INV_X1 U6966 ( .A(n8676), .ZN(n8684) );
  INV_X1 U6967 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7492) );
  INV_X1 U6968 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n9793) );
  MUX2_X1 U6969 ( .A(n7492), .B(n9793), .S(n4483), .Z(n5492) );
  INV_X1 U6970 ( .A(SI_20_), .ZN(n5491) );
  NAND2_X1 U6971 ( .A1(n5492), .A2(n5491), .ZN(n5509) );
  INV_X1 U6972 ( .A(n5492), .ZN(n5493) );
  NAND2_X1 U6973 ( .A1(n5493), .A2(SI_20_), .ZN(n5494) );
  XNOR2_X1 U6974 ( .A(n5508), .B(n5507), .ZN(n7490) );
  NAND2_X1 U6975 ( .A1(n7490), .A2(n5692), .ZN(n5496) );
  OR2_X1 U6976 ( .A1(n5693), .A2(n7492), .ZN(n5495) );
  NAND2_X1 U6977 ( .A1(n5675), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n5504) );
  NAND2_X1 U6978 ( .A1(n5676), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n5503) );
  INV_X1 U6979 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n5498) );
  NAND2_X1 U6980 ( .A1(n5499), .A2(n5498), .ZN(n5500) );
  AND2_X1 U6981 ( .A1(n5513), .A2(n5500), .ZN(n8664) );
  NAND2_X1 U6982 ( .A1(n5644), .A2(n8664), .ZN(n5502) );
  NAND2_X1 U6983 ( .A1(n5677), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n5501) );
  NAND2_X1 U6984 ( .A1(n8799), .A2(n8503), .ZN(n5787) );
  INV_X1 U6985 ( .A(n8667), .ZN(n5505) );
  NOR2_X1 U6986 ( .A1(n8669), .A2(n5505), .ZN(n5506) );
  INV_X1 U6987 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7580) );
  INV_X1 U6988 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7576) );
  MUX2_X1 U6989 ( .A(n7580), .B(n7576), .S(n4483), .Z(n5526) );
  XNOR2_X1 U6990 ( .A(n5526), .B(SI_21_), .ZN(n5521) );
  XNOR2_X1 U6991 ( .A(n5520), .B(n5521), .ZN(n7575) );
  NAND2_X1 U6992 ( .A1(n7575), .A2(n5692), .ZN(n5512) );
  OR2_X1 U6993 ( .A1(n5693), .A2(n7580), .ZN(n5511) );
  INV_X1 U6994 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n8260) );
  NAND2_X1 U6995 ( .A1(n5513), .A2(n8260), .ZN(n5514) );
  AND2_X1 U6996 ( .A1(n5538), .A2(n5514), .ZN(n8650) );
  NAND2_X1 U6997 ( .A1(n8650), .A2(n5644), .ZN(n5518) );
  NAND2_X1 U6998 ( .A1(n5675), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n5517) );
  NAND2_X1 U6999 ( .A1(n5676), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n5516) );
  NAND2_X1 U7000 ( .A1(n5677), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n5515) );
  NAND4_X1 U7001 ( .A1(n5518), .A2(n5517), .A3(n5516), .A4(n5515), .ZN(n8670)
         );
  XNOR2_X1 U7002 ( .A(n8794), .B(n8638), .ZN(n8653) );
  INV_X1 U7003 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7663) );
  INV_X1 U7004 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7659) );
  MUX2_X1 U7005 ( .A(n7663), .B(n7659), .S(n4483), .Z(n5523) );
  INV_X1 U7006 ( .A(SI_22_), .ZN(n5522) );
  NAND2_X1 U7007 ( .A1(n5523), .A2(n5522), .ZN(n5544) );
  INV_X1 U7008 ( .A(n5523), .ZN(n5524) );
  NAND2_X1 U7009 ( .A1(n5524), .A2(SI_22_), .ZN(n5525) );
  NAND2_X1 U7010 ( .A1(n5544), .A2(n5525), .ZN(n5532) );
  INV_X1 U7011 ( .A(n5532), .ZN(n5528) );
  INV_X1 U7012 ( .A(n5526), .ZN(n5527) );
  NAND2_X1 U7013 ( .A1(n5527), .A2(SI_21_), .ZN(n5530) );
  NAND2_X1 U7014 ( .A1(n5531), .A2(n5530), .ZN(n5533) );
  NAND2_X1 U7015 ( .A1(n5533), .A2(n5532), .ZN(n5534) );
  NAND2_X1 U7016 ( .A1(n5545), .A2(n5534), .ZN(n7658) );
  NAND2_X1 U7017 ( .A1(n7658), .A2(n5692), .ZN(n5536) );
  OR2_X1 U7018 ( .A1(n5693), .A2(n7663), .ZN(n5535) );
  INV_X1 U7019 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n5542) );
  INV_X1 U7020 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n9792) );
  NAND2_X1 U7021 ( .A1(n5538), .A2(n9792), .ZN(n5539) );
  NAND2_X1 U7022 ( .A1(n5556), .A2(n5539), .ZN(n8629) );
  OR2_X1 U7023 ( .A1(n8629), .A2(n5609), .ZN(n5541) );
  AOI22_X1 U7024 ( .A1(n5675), .A2(P2_REG0_REG_22__SCAN_IN), .B1(n5676), .B2(
        P2_REG1_REG_22__SCAN_IN), .ZN(n5540) );
  OAI211_X1 U7025 ( .C1(n5641), .C2(n5542), .A(n5541), .B(n5540), .ZN(n8656)
         );
  NAND2_X1 U7026 ( .A1(n8632), .A2(n8656), .ZN(n5781) );
  INV_X1 U7027 ( .A(n8656), .ZN(n8261) );
  NAND2_X1 U7028 ( .A1(n8789), .A2(n8261), .ZN(n5794) );
  INV_X1 U7029 ( .A(n8633), .ZN(n8626) );
  AND2_X1 U7030 ( .A1(n8794), .A2(n8638), .ZN(n5779) );
  NOR2_X1 U7031 ( .A1(n8626), .A2(n5779), .ZN(n5543) );
  INV_X1 U7032 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7718) );
  INV_X1 U7033 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7714) );
  MUX2_X1 U7034 ( .A(n7718), .B(n7714), .S(n4483), .Z(n5546) );
  INV_X1 U7035 ( .A(SI_23_), .ZN(n9587) );
  NAND2_X1 U7036 ( .A1(n5546), .A2(n9587), .ZN(n5561) );
  INV_X1 U7037 ( .A(n5546), .ZN(n5547) );
  NAND2_X1 U7038 ( .A1(n5547), .A2(SI_23_), .ZN(n5548) );
  NAND2_X1 U7039 ( .A1(n5561), .A2(n5548), .ZN(n5550) );
  NAND2_X1 U7040 ( .A1(n5549), .A2(n5550), .ZN(n5553) );
  INV_X1 U7041 ( .A(n5550), .ZN(n5551) );
  NAND2_X1 U7042 ( .A1(n5553), .A2(n5562), .ZN(n7715) );
  NAND2_X1 U7043 ( .A1(n7715), .A2(n5692), .ZN(n5555) );
  OR2_X1 U7044 ( .A1(n5693), .A2(n7718), .ZN(n5554) );
  INV_X1 U7045 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8619) );
  INV_X1 U7046 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8214) );
  NAND2_X1 U7047 ( .A1(n5556), .A2(n8214), .ZN(n5557) );
  NAND2_X1 U7048 ( .A1(n5566), .A2(n5557), .ZN(n8621) );
  OR2_X1 U7049 ( .A1(n8621), .A2(n5609), .ZN(n5559) );
  AOI22_X1 U7050 ( .A1(n5675), .A2(P2_REG0_REG_23__SCAN_IN), .B1(n5676), .B2(
        P2_REG1_REG_23__SCAN_IN), .ZN(n5558) );
  OAI211_X1 U7051 ( .C1(n5641), .C2(n8619), .A(n5559), .B(n5558), .ZN(n8505)
         );
  NAND2_X1 U7052 ( .A1(n8618), .A2(n8505), .ZN(n5799) );
  INV_X1 U7053 ( .A(n8505), .ZN(n8640) );
  NAND2_X1 U7054 ( .A1(n8784), .A2(n8640), .ZN(n5798) );
  INV_X1 U7055 ( .A(n8614), .ZN(n8606) );
  INV_X1 U7056 ( .A(n5781), .ZN(n8607) );
  NOR2_X1 U7057 ( .A1(n8606), .A2(n8607), .ZN(n5560) );
  MUX2_X1 U7058 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(P2_DATAO_REG_24__SCAN_IN), 
        .S(n4483), .Z(n5577) );
  INV_X1 U7059 ( .A(SI_24_), .ZN(n5563) );
  XNOR2_X1 U7060 ( .A(n5577), .B(n5563), .ZN(n5574) );
  XNOR2_X1 U7061 ( .A(n5576), .B(n5574), .ZN(n5962) );
  NAND2_X1 U7062 ( .A1(n5962), .A2(n5692), .ZN(n5565) );
  INV_X1 U7063 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7871) );
  OR2_X1 U7064 ( .A1(n5693), .A2(n7871), .ZN(n5564) );
  INV_X1 U7065 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n8305) );
  OR2_X2 U7066 ( .A1(n5566), .A2(n8305), .ZN(n5585) );
  NAND2_X1 U7067 ( .A1(n5566), .A2(n8305), .ZN(n5567) );
  AND2_X1 U7068 ( .A1(n5585), .A2(n5567), .ZN(n8600) );
  NAND2_X1 U7069 ( .A1(n8600), .A2(n5644), .ZN(n5573) );
  INV_X1 U7070 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n5570) );
  NAND2_X1 U7071 ( .A1(n5675), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n5569) );
  NAND2_X1 U7072 ( .A1(n5676), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n5568) );
  OAI211_X1 U7073 ( .C1(n5570), .C2(n5641), .A(n5569), .B(n5568), .ZN(n5571)
         );
  INV_X1 U7074 ( .A(n5571), .ZN(n5572) );
  INV_X1 U7075 ( .A(n5574), .ZN(n5575) );
  INV_X1 U7076 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7949) );
  INV_X1 U7077 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7950) );
  MUX2_X1 U7078 ( .A(n7949), .B(n7950), .S(n4483), .Z(n5579) );
  INV_X1 U7079 ( .A(SI_25_), .ZN(n5578) );
  NAND2_X1 U7080 ( .A1(n5579), .A2(n5578), .ZN(n5592) );
  INV_X1 U7081 ( .A(n5579), .ZN(n5580) );
  NAND2_X1 U7082 ( .A1(n5580), .A2(SI_25_), .ZN(n5581) );
  NAND2_X1 U7083 ( .A1(n5592), .A2(n5581), .ZN(n5593) );
  NAND2_X1 U7084 ( .A1(n7945), .A2(n5692), .ZN(n5583) );
  OR2_X1 U7085 ( .A1(n5693), .A2(n7949), .ZN(n5582) );
  INV_X1 U7086 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8270) );
  NAND2_X1 U7087 ( .A1(n5585), .A2(n8270), .ZN(n5586) );
  NAND2_X1 U7088 ( .A1(n5607), .A2(n5586), .ZN(n8587) );
  OR2_X1 U7089 ( .A1(n8587), .A2(n5609), .ZN(n5591) );
  INV_X1 U7090 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n8586) );
  NAND2_X1 U7091 ( .A1(n5675), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n5588) );
  NAND2_X1 U7092 ( .A1(n5676), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n5587) );
  OAI211_X1 U7093 ( .C1(n8586), .C2(n5641), .A(n5588), .B(n5587), .ZN(n5589)
         );
  INV_X1 U7094 ( .A(n5589), .ZN(n5590) );
  NAND2_X1 U7095 ( .A1(n8773), .A2(n8572), .ZN(n5804) );
  INV_X1 U7096 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n8062) );
  INV_X1 U7097 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n9681) );
  MUX2_X1 U7098 ( .A(n8062), .B(n9681), .S(n4483), .Z(n5596) );
  INV_X1 U7099 ( .A(SI_26_), .ZN(n9836) );
  NAND2_X1 U7100 ( .A1(n5596), .A2(n9836), .ZN(n5616) );
  INV_X1 U7101 ( .A(n5596), .ZN(n5597) );
  NAND2_X1 U7102 ( .A1(n5597), .A2(SI_26_), .ZN(n5598) );
  NAND2_X1 U7103 ( .A1(n5616), .A2(n5598), .ZN(n5600) );
  NAND2_X1 U7104 ( .A1(n5599), .A2(n5600), .ZN(n5602) );
  INV_X1 U7105 ( .A(n5600), .ZN(n5601) );
  NAND2_X1 U7106 ( .A1(n5602), .A2(n5617), .ZN(n8060) );
  NAND2_X1 U7107 ( .A1(n8060), .A2(n5692), .ZN(n5604) );
  OR2_X1 U7108 ( .A1(n5693), .A2(n8062), .ZN(n5603) );
  INV_X1 U7109 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n5606) );
  NAND2_X1 U7110 ( .A1(n5607), .A2(n5606), .ZN(n5608) );
  NAND2_X1 U7111 ( .A1(n5637), .A2(n5608), .ZN(n8564) );
  OR2_X1 U7112 ( .A1(n8564), .A2(n5609), .ZN(n5614) );
  INV_X1 U7113 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8563) );
  NAND2_X1 U7114 ( .A1(n5675), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n5611) );
  NAND2_X1 U7115 ( .A1(n5676), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n5610) );
  OAI211_X1 U7116 ( .C1(n8563), .C2(n5641), .A(n5611), .B(n5610), .ZN(n5612)
         );
  INV_X1 U7117 ( .A(n5612), .ZN(n5613) );
  INV_X1 U7118 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n8139) );
  INV_X1 U7119 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n9863) );
  MUX2_X1 U7120 ( .A(n8139), .B(n9863), .S(n4483), .Z(n5618) );
  INV_X1 U7121 ( .A(SI_27_), .ZN(n9865) );
  NAND2_X1 U7122 ( .A1(n5618), .A2(n9865), .ZN(n5631) );
  INV_X1 U7123 ( .A(n5618), .ZN(n5619) );
  NAND2_X1 U7124 ( .A1(n5619), .A2(SI_27_), .ZN(n5620) );
  AND2_X1 U7125 ( .A1(n5631), .A2(n5620), .ZN(n5629) );
  NAND2_X1 U7126 ( .A1(n6312), .A2(n5692), .ZN(n5622) );
  OR2_X1 U7127 ( .A1(n5693), .A2(n8139), .ZN(n5621) );
  XNOR2_X1 U7128 ( .A(n5637), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n8551) );
  NAND2_X1 U7129 ( .A1(n8551), .A2(n5644), .ZN(n5628) );
  INV_X1 U7130 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n5625) );
  NAND2_X1 U7131 ( .A1(n5675), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n5624) );
  NAND2_X1 U7132 ( .A1(n5676), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n5623) );
  OAI211_X1 U7133 ( .C1(n5625), .C2(n5641), .A(n5624), .B(n5623), .ZN(n5626)
         );
  INV_X1 U7134 ( .A(n5626), .ZN(n5627) );
  OR2_X1 U7135 ( .A1(n8194), .A2(n8573), .ZN(n5814) );
  INV_X1 U7136 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8135) );
  INV_X1 U7137 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n9866) );
  MUX2_X1 U7138 ( .A(n8135), .B(n9866), .S(n4483), .Z(n5648) );
  XNOR2_X1 U7139 ( .A(n5648), .B(SI_28_), .ZN(n5646) );
  OR2_X1 U7140 ( .A1(n5693), .A2(n8135), .ZN(n5633) );
  INV_X1 U7141 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n8206) );
  INV_X1 U7142 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n5635) );
  OAI21_X1 U7143 ( .B1(n5637), .B2(n8206), .A(n5635), .ZN(n5638) );
  NAND2_X1 U7144 ( .A1(P2_REG3_REG_28__SCAN_IN), .A2(P2_REG3_REG_27__SCAN_IN), 
        .ZN(n5636) );
  OR2_X2 U7145 ( .A1(n5637), .A2(n5636), .ZN(n5654) );
  INV_X1 U7146 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n5642) );
  NAND2_X1 U7147 ( .A1(n5675), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n5640) );
  NAND2_X1 U7148 ( .A1(n5676), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n5639) );
  OAI211_X1 U7149 ( .C1(n5642), .C2(n5641), .A(n5640), .B(n5639), .ZN(n5643)
         );
  AOI21_X2 U7150 ( .B1(n8533), .B2(n5660), .A(n5643), .ZN(n8548) );
  NAND2_X1 U7151 ( .A1(n5816), .A2(n5819), .ZN(n8530) );
  INV_X1 U7152 ( .A(n8530), .ZN(n5865) );
  NAND2_X1 U7153 ( .A1(n5645), .A2(n5816), .ZN(n8514) );
  INV_X1 U7154 ( .A(SI_28_), .ZN(n9845) );
  NAND2_X1 U7155 ( .A1(n5648), .A2(n9845), .ZN(n5661) );
  NAND2_X1 U7156 ( .A1(n5664), .A2(n5661), .ZN(n5651) );
  MUX2_X1 U7157 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .S(n4483), .Z(n5666) );
  INV_X1 U7158 ( .A(SI_29_), .ZN(n5649) );
  XNOR2_X1 U7159 ( .A(n5666), .B(n5649), .ZN(n5650) );
  NAND2_X1 U7160 ( .A1(n8872), .A2(n5692), .ZN(n5653) );
  INV_X1 U7161 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8875) );
  OR2_X1 U7162 ( .A1(n5693), .A2(n8875), .ZN(n5652) );
  INV_X1 U7163 ( .A(n5654), .ZN(n8520) );
  INV_X1 U7164 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n5658) );
  NAND2_X1 U7165 ( .A1(n5675), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n5656) );
  NAND2_X1 U7166 ( .A1(n5677), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n5655) );
  OAI211_X1 U7167 ( .C1(n5658), .C2(n5657), .A(n5656), .B(n5655), .ZN(n5659)
         );
  AOI21_X1 U7168 ( .B1(n8520), .B2(n5660), .A(n5659), .ZN(n8248) );
  NAND2_X1 U7169 ( .A1(n8483), .A2(n8248), .ZN(n5826) );
  NOR2_X1 U7170 ( .A1(n5666), .A2(SI_29_), .ZN(n5663) );
  INV_X1 U7171 ( .A(n5661), .ZN(n5662) );
  NOR2_X1 U7172 ( .A1(n5663), .A2(n5662), .ZN(n5665) );
  NAND2_X1 U7173 ( .A1(n5665), .A2(n5664), .ZN(n5668) );
  NAND2_X1 U7174 ( .A1(n5666), .A2(SI_29_), .ZN(n5667) );
  MUX2_X1 U7175 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .S(n4483), .Z(n5685) );
  NAND2_X1 U7176 ( .A1(n5676), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n5672) );
  NAND2_X1 U7177 ( .A1(n5677), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n5671) );
  NAND2_X1 U7178 ( .A1(n5675), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n5670) );
  AND3_X1 U7179 ( .A1(n5672), .A2(n5671), .A3(n5670), .ZN(n8485) );
  NAND2_X1 U7180 ( .A1(n4514), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5673) );
  NAND2_X1 U7181 ( .A1(n8485), .A2(n6987), .ZN(n5674) );
  OAI21_X1 U7182 ( .B1(n9906), .B2(n5674), .A(n5826), .ZN(n5682) );
  INV_X1 U7183 ( .A(n5674), .ZN(n5681) );
  NAND2_X1 U7184 ( .A1(n5675), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n5680) );
  NAND2_X1 U7185 ( .A1(n5676), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n5679) );
  NAND2_X1 U7186 ( .A1(n5677), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n5678) );
  AND3_X1 U7187 ( .A1(n5680), .A2(n5679), .A3(n5678), .ZN(n8517) );
  INV_X1 U7188 ( .A(n8517), .ZN(n8367) );
  NAND2_X1 U7189 ( .A1(n9906), .A2(n8367), .ZN(n5827) );
  OAI22_X1 U7190 ( .A1(n8513), .A2(n5682), .B1(n5681), .B2(n5827), .ZN(n5696)
         );
  INV_X1 U7191 ( .A(n5683), .ZN(n5684) );
  NAND2_X1 U7192 ( .A1(n5684), .A2(SI_30_), .ZN(n5688) );
  NAND2_X1 U7193 ( .A1(n5686), .A2(n5685), .ZN(n5687) );
  MUX2_X1 U7194 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n4483), .Z(n5689) );
  XNOR2_X1 U7195 ( .A(n5689), .B(SI_31_), .ZN(n5690) );
  NAND2_X1 U7196 ( .A1(n8863), .A2(n5692), .ZN(n5695) );
  INV_X1 U7197 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n8866) );
  OR2_X1 U7198 ( .A1(n5693), .A2(n8866), .ZN(n5694) );
  NOR2_X1 U7199 ( .A1(n9906), .A2(n8367), .ZN(n5828) );
  NOR2_X1 U7200 ( .A1(n5706), .A2(n5828), .ZN(n5707) );
  NAND2_X1 U7201 ( .A1(n5696), .A2(n5707), .ZN(n5698) );
  INV_X1 U7202 ( .A(n5832), .ZN(n5697) );
  NAND2_X1 U7203 ( .A1(n5698), .A2(n5697), .ZN(n5699) );
  XNOR2_X1 U7204 ( .A(n5699), .B(n4781), .ZN(n5704) );
  NAND2_X1 U7205 ( .A1(n5700), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5876) );
  XNOR2_X1 U7206 ( .A(n5876), .B(P2_IR_REG_22__SCAN_IN), .ZN(n7219) );
  INV_X1 U7207 ( .A(n7219), .ZN(n7661) );
  NAND2_X1 U7208 ( .A1(n7661), .A2(n7578), .ZN(n10277) );
  NAND2_X1 U7209 ( .A1(n4542), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5701) );
  MUX2_X1 U7210 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5701), .S(
        P2_IR_REG_20__SCAN_IN), .Z(n5702) );
  NAND2_X1 U7211 ( .A1(n5702), .A2(n4514), .ZN(n7491) );
  INV_X1 U7212 ( .A(n7491), .ZN(n5870) );
  NAND2_X1 U7213 ( .A1(n6987), .A2(n5870), .ZN(n7224) );
  NAND2_X1 U7214 ( .A1(n8168), .A2(n7224), .ZN(n5703) );
  NAND2_X1 U7215 ( .A1(n6987), .A2(n4781), .ZN(n5705) );
  OR2_X1 U7216 ( .A1(n7219), .A2(n5705), .ZN(n5824) );
  INV_X1 U7217 ( .A(n5706), .ZN(n5835) );
  INV_X1 U7218 ( .A(n5707), .ZN(n5868) );
  INV_X1 U7219 ( .A(n5797), .ZN(n5802) );
  NAND2_X1 U7220 ( .A1(n10249), .A2(n5731), .ZN(n5709) );
  NAND2_X1 U7221 ( .A1(n5712), .A2(n5711), .ZN(n5708) );
  MUX2_X1 U7222 ( .A(n5709), .B(n5708), .S(n4692), .Z(n5733) );
  INV_X1 U7223 ( .A(n5737), .ZN(n5714) );
  INV_X1 U7224 ( .A(n5712), .ZN(n5713) );
  NOR3_X1 U7225 ( .A1(n5715), .A2(n5714), .A3(n5713), .ZN(n5729) );
  INV_X1 U7226 ( .A(n5842), .ZN(n5717) );
  INV_X1 U7227 ( .A(n7363), .ZN(n10276) );
  NAND2_X1 U7228 ( .A1(n8385), .A2(n10276), .ZN(n5844) );
  INV_X1 U7229 ( .A(n5844), .ZN(n5716) );
  OAI211_X1 U7230 ( .C1(n5717), .C2(n5716), .A(n5721), .B(n5843), .ZN(n5718)
         );
  NAND2_X1 U7231 ( .A1(n5718), .A2(n5720), .ZN(n5725) );
  AOI21_X1 U7232 ( .B1(n6987), .B2(n5844), .A(n5719), .ZN(n5723) );
  NAND2_X1 U7233 ( .A1(n5842), .A2(n5720), .ZN(n5722) );
  OAI21_X1 U7234 ( .B1(n5723), .B2(n5722), .A(n5721), .ZN(n5724) );
  MUX2_X1 U7235 ( .A(n5725), .B(n5724), .S(n5824), .Z(n5727) );
  INV_X1 U7236 ( .A(n5733), .ZN(n5726) );
  NAND3_X1 U7237 ( .A1(n5727), .A2(n5726), .A3(n7413), .ZN(n5728) );
  OAI21_X1 U7238 ( .B1(n5729), .B2(n4692), .A(n5728), .ZN(n5736) );
  AOI21_X1 U7239 ( .B1(n10302), .B2(n8382), .A(n5730), .ZN(n5732) );
  OAI211_X1 U7240 ( .C1(n5733), .C2(n5732), .A(n5735), .B(n5731), .ZN(n5734)
         );
  OAI21_X1 U7241 ( .B1(n5737), .B2(n5824), .A(n5241), .ZN(n5741) );
  INV_X1 U7242 ( .A(n8378), .ZN(n7599) );
  NAND2_X1 U7243 ( .A1(n7599), .A2(n5824), .ZN(n5739) );
  NAND2_X1 U7244 ( .A1(n8378), .A2(n4692), .ZN(n5738) );
  MUX2_X1 U7245 ( .A(n5739), .B(n5738), .S(n7591), .Z(n5740) );
  NAND2_X1 U7246 ( .A1(n7680), .A2(n4692), .ZN(n5744) );
  INV_X1 U7247 ( .A(n7680), .ZN(n10321) );
  NAND2_X1 U7248 ( .A1(n10321), .A2(n5824), .ZN(n5743) );
  MUX2_X1 U7249 ( .A(n5744), .B(n5743), .S(n8377), .Z(n5745) );
  NAND3_X1 U7250 ( .A1(n5746), .A2(n7809), .A3(n5745), .ZN(n5755) );
  NAND2_X1 U7251 ( .A1(n5747), .A2(n5748), .ZN(n5750) );
  INV_X1 U7252 ( .A(n5750), .ZN(n5754) );
  NAND2_X1 U7253 ( .A1(n5854), .A2(n5748), .ZN(n5752) );
  OAI211_X1 U7254 ( .C1(n5750), .C2(n5850), .A(n5855), .B(n5749), .ZN(n5751)
         );
  MUX2_X1 U7255 ( .A(n5752), .B(n5751), .S(n5824), .Z(n5753) );
  INV_X1 U7256 ( .A(n5756), .ZN(n5757) );
  MUX2_X1 U7257 ( .A(n5758), .B(n5757), .S(n5824), .Z(n5759) );
  XNOR2_X1 U7258 ( .A(n8495), .B(n8281), .ZN(n8114) );
  INV_X1 U7259 ( .A(n8114), .ZN(n5858) );
  MUX2_X1 U7260 ( .A(n5761), .B(n5760), .S(n5824), .Z(n5762) );
  NAND2_X1 U7261 ( .A1(n5858), .A2(n5762), .ZN(n5765) );
  INV_X1 U7262 ( .A(n8495), .ZN(n8826) );
  INV_X1 U7263 ( .A(n8281), .ZN(n8494) );
  MUX2_X1 U7264 ( .A(n8495), .B(n8494), .S(n5824), .Z(n5763) );
  OAI21_X1 U7265 ( .B1(n8826), .B2(n8281), .A(n5763), .ZN(n5764) );
  OAI211_X1 U7266 ( .C1(n5766), .C2(n5765), .A(n8728), .B(n5764), .ZN(n5770)
         );
  INV_X1 U7267 ( .A(n8712), .ZN(n5860) );
  MUX2_X1 U7268 ( .A(n5768), .B(n5767), .S(n5824), .Z(n5769) );
  NAND3_X1 U7269 ( .A1(n5770), .A2(n5860), .A3(n5769), .ZN(n5775) );
  INV_X1 U7270 ( .A(n5841), .ZN(n5776) );
  INV_X1 U7271 ( .A(n5785), .ZN(n5840) );
  AOI21_X1 U7272 ( .B1(n5771), .B2(n8816), .A(n5840), .ZN(n5773) );
  MUX2_X1 U7273 ( .A(n5773), .B(n5772), .S(n5824), .Z(n5774) );
  NAND3_X1 U7274 ( .A1(n5775), .A2(n5776), .A3(n5774), .ZN(n5786) );
  NAND3_X1 U7275 ( .A1(n5786), .A2(n5783), .A3(n5776), .ZN(n5778) );
  INV_X1 U7276 ( .A(n5789), .ZN(n5777) );
  INV_X1 U7277 ( .A(n5779), .ZN(n8634) );
  NAND2_X1 U7278 ( .A1(n8634), .A2(n5787), .ZN(n5780) );
  NAND2_X1 U7279 ( .A1(n8652), .A2(n8670), .ZN(n5788) );
  MUX2_X1 U7280 ( .A(n5782), .B(n5781), .S(n5824), .Z(n5796) );
  INV_X1 U7281 ( .A(n5783), .ZN(n5784) );
  AOI21_X1 U7282 ( .B1(n5786), .B2(n5785), .A(n5784), .ZN(n5791) );
  NAND2_X1 U7283 ( .A1(n5787), .A2(n8667), .ZN(n5790) );
  OAI211_X1 U7284 ( .C1(n5791), .C2(n5790), .A(n5789), .B(n5788), .ZN(n5792)
         );
  NAND3_X1 U7285 ( .A1(n5792), .A2(n5794), .A3(n8634), .ZN(n5793) );
  MUX2_X1 U7286 ( .A(n5794), .B(n5793), .S(n5824), .Z(n5795) );
  AOI21_X1 U7287 ( .B1(n5801), .B2(n5799), .A(n5824), .ZN(n5800) );
  NAND2_X1 U7288 ( .A1(n5807), .A2(n5803), .ZN(n5806) );
  NAND2_X1 U7289 ( .A1(n5615), .A2(n5804), .ZN(n5805) );
  MUX2_X1 U7290 ( .A(n5806), .B(n5805), .S(n5824), .Z(n5810) );
  MUX2_X1 U7291 ( .A(n5808), .B(n5807), .S(n5824), .Z(n5809) );
  INV_X1 U7292 ( .A(n5819), .ZN(n5812) );
  AOI21_X1 U7293 ( .B1(n8573), .B2(n8194), .A(n5812), .ZN(n5813) );
  MUX2_X1 U7294 ( .A(n5814), .B(n5813), .S(n5824), .Z(n5815) );
  INV_X1 U7295 ( .A(n5825), .ZN(n5818) );
  NOR2_X1 U7296 ( .A1(n5818), .A2(n5824), .ZN(n5822) );
  OAI211_X1 U7297 ( .C1(n4692), .C2(n8755), .A(n5820), .B(n5819), .ZN(n5821)
         );
  OAI21_X1 U7298 ( .B1(n5823), .B2(n5822), .A(n5821), .ZN(n5830) );
  MUX2_X1 U7299 ( .A(n5826), .B(n5825), .S(n4687), .Z(n5829) );
  INV_X1 U7300 ( .A(n5827), .ZN(n5831) );
  NOR2_X1 U7301 ( .A1(n5831), .A2(n5832), .ZN(n5839) );
  OAI22_X1 U7302 ( .A1(n5833), .A2(n5832), .B1(n5839), .B2(n4692), .ZN(n5834)
         );
  OAI21_X1 U7303 ( .B1(n4692), .B2(n5835), .A(n5834), .ZN(n5836) );
  NAND2_X1 U7304 ( .A1(n5836), .A2(n7491), .ZN(n5872) );
  NAND2_X1 U7305 ( .A1(n7219), .A2(n4781), .ZN(n7225) );
  INV_X1 U7306 ( .A(n7225), .ZN(n5838) );
  INV_X1 U7307 ( .A(n10277), .ZN(n5837) );
  INV_X1 U7308 ( .A(n5839), .ZN(n5867) );
  NOR2_X1 U7309 ( .A1(n5841), .A2(n5840), .ZN(n8699) );
  NOR2_X1 U7310 ( .A1(n7367), .A2(n7444), .ZN(n5848) );
  NOR2_X1 U7311 ( .A1(n10251), .A2(n7329), .ZN(n5847) );
  NAND2_X1 U7312 ( .A1(n7223), .A2(n5844), .ZN(n7362) );
  NOR2_X1 U7313 ( .A1(n7362), .A2(n7491), .ZN(n5845) );
  NAND4_X1 U7314 ( .A1(n5848), .A2(n5847), .A3(n5846), .A4(n5845), .ZN(n5849)
         );
  NOR2_X1 U7315 ( .A1(n5849), .A2(n7371), .ZN(n5851) );
  AND4_X1 U7316 ( .A1(n5851), .A2(n7762), .A3(n5241), .A4(n7597), .ZN(n5856)
         );
  NAND2_X1 U7317 ( .A1(n5855), .A2(n5854), .ZN(n7920) );
  INV_X1 U7318 ( .A(n7920), .ZN(n7765) );
  NAND4_X1 U7319 ( .A1(n5856), .A2(n8010), .A3(n7765), .A4(n7812), .ZN(n5857)
         );
  NOR4_X1 U7320 ( .A1(n8735), .A2(n8051), .A3(n4943), .A4(n5857), .ZN(n5859)
         );
  NAND4_X1 U7321 ( .A1(n5860), .A2(n8699), .A3(n5859), .A4(n5858), .ZN(n5861)
         );
  NOR4_X1 U7322 ( .A1(n8626), .A2(n8669), .A3(n8676), .A4(n5861), .ZN(n5862)
         );
  NAND2_X1 U7323 ( .A1(n8614), .A2(n5862), .ZN(n5863) );
  NOR4_X1 U7324 ( .A1(n8570), .A2(n8653), .A3(n8597), .A4(n5863), .ZN(n5864)
         );
  NAND4_X1 U7325 ( .A1(n5865), .A2(n4681), .A3(n5864), .A4(n8543), .ZN(n5866)
         );
  NOR4_X1 U7326 ( .A1(n5868), .A2(n5867), .A3(n8515), .A4(n5866), .ZN(n5869)
         );
  XNOR2_X1 U7327 ( .A(n5869), .B(n4781), .ZN(n5871) );
  OAI22_X1 U7328 ( .A1(n5871), .A2(n6987), .B1(n5870), .B2(n7225), .ZN(n5873)
         );
  INV_X1 U7329 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5875) );
  NAND2_X1 U7330 ( .A1(n5876), .A2(n5875), .ZN(n5877) );
  NAND2_X1 U7331 ( .A1(n5877), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5886) );
  INV_X1 U7332 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5885) );
  XNOR2_X1 U7333 ( .A(n5886), .B(n5885), .ZN(n7017) );
  OR2_X1 U7334 ( .A1(n7017), .A2(P2_U3152), .ZN(n7716) );
  NAND2_X1 U7335 ( .A1(n5881), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5882) );
  XNOR2_X1 U7336 ( .A(n5882), .B(P2_IR_REG_26__SCAN_IN), .ZN(n6995) );
  NAND2_X1 U7337 ( .A1(n5883), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5884) );
  XNOR2_X1 U7338 ( .A(n5884), .B(P2_IR_REG_25__SCAN_IN), .ZN(n7946) );
  NAND2_X1 U7339 ( .A1(n6995), .A2(n7946), .ZN(n5890) );
  NAND2_X1 U7340 ( .A1(n5886), .A2(n5885), .ZN(n5887) );
  NAND2_X1 U7341 ( .A1(n5887), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5889) );
  INV_X1 U7342 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5888) );
  XNOR2_X1 U7343 ( .A(n5889), .B(n5888), .ZN(n7872) );
  AND2_X1 U7344 ( .A1(n7491), .A2(n8478), .ZN(n7018) );
  NAND2_X1 U7345 ( .A1(n10268), .A2(n7018), .ZN(n7217) );
  INV_X1 U7346 ( .A(n7089), .ZN(n5891) );
  NAND2_X1 U7347 ( .A1(n7219), .A2(n6987), .ZN(n7057) );
  INV_X1 U7348 ( .A(n7057), .ZN(n7011) );
  NAND2_X1 U7349 ( .A1(n5891), .A2(n7011), .ZN(n8637) );
  NOR3_X1 U7350 ( .A1(n7217), .A2(n8484), .A3(n8637), .ZN(n5893) );
  OAI21_X1 U7351 ( .B1(n7716), .B2(n7219), .A(P2_B_REG_SCAN_IN), .ZN(n5892) );
  NAND2_X1 U7352 ( .A1(n5894), .A2(n5082), .ZN(P2_U3244) );
  NAND2_X1 U7353 ( .A1(n6020), .A2(n5898), .ZN(n6044) );
  INV_X1 U7354 ( .A(n6044), .ZN(n5899) );
  NAND2_X1 U7355 ( .A1(n5900), .A2(n5899), .ZN(n5985) );
  INV_X1 U7356 ( .A(n5985), .ZN(n5908) );
  NOR2_X1 U7357 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n5903) );
  NAND4_X1 U7358 ( .A1(n5903), .A2(n5990), .A3(n5902), .A4(n5901), .ZN(n5906)
         );
  NAND4_X1 U7359 ( .A1(n5904), .A2(n6183), .A3(n9723), .A4(n5986), .ZN(n5905)
         );
  INV_X1 U7360 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n6474) );
  INV_X1 U7361 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5911) );
  NAND2_X1 U7362 ( .A1(n6474), .A2(n5911), .ZN(n5912) );
  INV_X1 U7363 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5915) );
  INV_X1 U7364 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5913) );
  XNOR2_X2 U7365 ( .A(n5916), .B(n5915), .ZN(n6481) );
  NAND2_X1 U7366 ( .A1(n8863), .A2(n6351), .ZN(n5920) );
  INV_X1 U7367 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n5918) );
  OR2_X1 U7368 ( .A1(n6352), .A2(n5918), .ZN(n5919) );
  INV_X1 U7369 ( .A(n9388), .ZN(n5934) );
  NAND2_X1 U7370 ( .A1(n5924), .A2(n5923), .ZN(n9483) );
  INV_X1 U7371 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n5925) );
  NAND2_X1 U7372 ( .A1(n5927), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5928) );
  NAND2_X1 U7373 ( .A1(n4486), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n5933) );
  INV_X1 U7374 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n5929) );
  OR2_X1 U7375 ( .A1(n6035), .A2(n5929), .ZN(n5932) );
  INV_X1 U7376 ( .A(n6032), .ZN(n6023) );
  INV_X1 U7377 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n5930) );
  OR2_X1 U7378 ( .A1(n6032), .A2(n5930), .ZN(n5931) );
  AND3_X1 U7379 ( .A1(n5933), .A2(n5932), .A3(n5931), .ZN(n6363) );
  NAND2_X1 U7380 ( .A1(n5934), .A2(n6363), .ZN(n6375) );
  NAND2_X1 U7381 ( .A1(n6484), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6371) );
  INV_X1 U7382 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n6370) );
  NAND2_X1 U7383 ( .A1(n6371), .A2(n6370), .ZN(n5935) );
  NAND2_X1 U7384 ( .A1(n5935), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5936) );
  NAND2_X1 U7385 ( .A1(n7660), .A2(n10138), .ZN(n7351) );
  AND2_X1 U7386 ( .A1(n6375), .A2(n7351), .ZN(n6365) );
  NAND2_X1 U7387 ( .A1(n7945), .A2(n6351), .ZN(n5938) );
  OR2_X1 U7388 ( .A1(n6352), .A2(n7950), .ZN(n5937) );
  INV_X1 U7389 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n6133) );
  INV_X1 U7390 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n8070) );
  INV_X1 U7391 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n6176) );
  INV_X1 U7392 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n6218) );
  AND2_X1 U7393 ( .A1(P1_REG3_REG_17__SCAN_IN), .A2(P1_REG3_REG_16__SCAN_IN), 
        .ZN(n5946) );
  INV_X1 U7394 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n8906) );
  INV_X1 U7395 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n8914) );
  INV_X1 U7396 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n8896) );
  INV_X1 U7397 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n8922) );
  NAND2_X1 U7398 ( .A1(n5967), .A2(n8922), .ZN(n5953) );
  NAND2_X1 U7399 ( .A1(n6298), .A2(n5953), .ZN(n9183) );
  INV_X1 U7400 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n5958) );
  NAND2_X1 U7401 ( .A1(n6276), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5957) );
  NAND2_X1 U7402 ( .A1(n6036), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5956) );
  OAI211_X1 U7403 ( .C1(n6358), .C2(n5958), .A(n5957), .B(n5956), .ZN(n5959)
         );
  INV_X1 U7404 ( .A(n5959), .ZN(n5960) );
  NAND2_X1 U7405 ( .A1(n5962), .A2(n6351), .ZN(n5964) );
  INV_X1 U7406 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n9779) );
  OR2_X1 U7407 ( .A1(n6352), .A2(n9779), .ZN(n5963) );
  INV_X1 U7408 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n5965) );
  NAND2_X1 U7409 ( .A1(n5977), .A2(n5965), .ZN(n5966) );
  NAND2_X1 U7410 ( .A1(n5967), .A2(n5966), .ZN(n9205) );
  OR2_X1 U7411 ( .A1(n9205), .A2(n6235), .ZN(n5973) );
  INV_X1 U7412 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n5970) );
  NAND2_X1 U7413 ( .A1(n6036), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5969) );
  NAND2_X1 U7414 ( .A1(n6276), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5968) );
  OAI211_X1 U7415 ( .C1(n6358), .C2(n5970), .A(n5969), .B(n5968), .ZN(n5971)
         );
  INV_X1 U7416 ( .A(n5971), .ZN(n5972) );
  NAND2_X1 U7417 ( .A1(n7715), .A2(n6351), .ZN(n5975) );
  OR2_X1 U7418 ( .A1(n6352), .A2(n7714), .ZN(n5974) );
  NAND2_X1 U7419 ( .A1(n6285), .A2(n8896), .ZN(n5976) );
  AND2_X1 U7420 ( .A1(n5977), .A2(n5976), .ZN(n9210) );
  NAND2_X1 U7421 ( .A1(n9210), .A2(n6346), .ZN(n5983) );
  INV_X1 U7422 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n5980) );
  NAND2_X1 U7423 ( .A1(n6036), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n5979) );
  NAND2_X1 U7424 ( .A1(n6276), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5978) );
  OAI211_X1 U7425 ( .C1(n6358), .C2(n5980), .A(n5979), .B(n5978), .ZN(n5981)
         );
  INV_X1 U7426 ( .A(n5981), .ZN(n5982) );
  INV_X1 U7427 ( .A(n9198), .ZN(n9237) );
  NAND2_X1 U7428 ( .A1(n9426), .A2(n9237), .ZN(n6377) );
  NAND2_X1 U7429 ( .A1(n9119), .A2(n6377), .ZN(n6295) );
  NAND2_X1 U7430 ( .A1(n9086), .A2(n9198), .ZN(n6413) );
  INV_X1 U7431 ( .A(n6413), .ZN(n9118) );
  AND2_X1 U7432 ( .A1(n9119), .A2(n9118), .ZN(n5984) );
  NAND2_X1 U7433 ( .A1(n7234), .A2(n6351), .ZN(n5994) );
  NOR2_X1 U7434 ( .A1(n5985), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n6152) );
  AND2_X1 U7435 ( .A1(n6152), .A2(n5986), .ZN(n6120) );
  NOR2_X1 U7436 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n5987) );
  NAND2_X1 U7437 ( .A1(n6120), .A2(n5987), .ZN(n6171) );
  OR2_X1 U7438 ( .A1(n6171), .A2(P1_IR_REG_14__SCAN_IN), .ZN(n6214) );
  OAI21_X1 U7439 ( .B1(n6214), .B2(P1_IR_REG_15__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6229) );
  INV_X1 U7440 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5988) );
  NAND2_X1 U7441 ( .A1(n6229), .A2(n5988), .ZN(n5989) );
  NAND2_X1 U7442 ( .A1(n5989), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6001) );
  NAND2_X1 U7443 ( .A1(n6001), .A2(n5990), .ZN(n5991) );
  NAND2_X1 U7444 ( .A1(n5991), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5992) );
  XNOR2_X1 U7445 ( .A(n5992), .B(P1_IR_REG_18__SCAN_IN), .ZN(n10115) );
  AOI22_X1 U7446 ( .A1(n6246), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n4752), .B2(
        n10115), .ZN(n5993) );
  NAND2_X1 U7447 ( .A1(n6276), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n6000) );
  INV_X1 U7448 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9046) );
  OR2_X1 U7449 ( .A1(n6358), .A2(n9046), .ZN(n5999) );
  INV_X1 U7450 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n10108) );
  NAND2_X1 U7451 ( .A1(n6007), .A2(n10108), .ZN(n5995) );
  NAND2_X1 U7452 ( .A1(n6249), .A2(n5995), .ZN(n9283) );
  OR2_X1 U7453 ( .A1(n6235), .A2(n9283), .ZN(n5998) );
  INV_X1 U7454 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n5996) );
  OR2_X1 U7455 ( .A1(n6288), .A2(n5996), .ZN(n5997) );
  NAND2_X1 U7456 ( .A1(n9452), .A2(n9011), .ZN(n9110) );
  NAND2_X1 U7457 ( .A1(n7201), .A2(n6351), .ZN(n6003) );
  XNOR2_X1 U7458 ( .A(n6001), .B(P1_IR_REG_17__SCAN_IN), .ZN(n10101) );
  AOI22_X1 U7459 ( .A1(n6246), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n4752), .B2(
        n10101), .ZN(n6002) );
  NAND2_X1 U7460 ( .A1(n6276), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n6011) );
  INV_X1 U7461 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9044) );
  OR2_X1 U7462 ( .A1(n6358), .A2(n9044), .ZN(n6010) );
  INV_X1 U7463 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n6004) );
  OR2_X1 U7464 ( .A1(n6288), .A2(n6004), .ZN(n6009) );
  INV_X1 U7465 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n6233) );
  INV_X1 U7466 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n6005) );
  OAI21_X1 U7467 ( .B1(n6234), .B2(n6233), .A(n6005), .ZN(n6006) );
  NAND2_X1 U7468 ( .A1(n6007), .A2(n6006), .ZN(n9299) );
  OR2_X1 U7469 ( .A1(n6235), .A2(n9299), .ZN(n6008) );
  NAND4_X1 U7470 ( .A1(n6011), .A2(n6010), .A3(n6009), .A4(n6008), .ZN(n9314)
         );
  INV_X1 U7471 ( .A(n9314), .ZN(n9078) );
  NAND2_X1 U7472 ( .A1(n9458), .A2(n9078), .ZN(n9109) );
  AND2_X1 U7473 ( .A1(n9110), .A2(n9109), .ZN(n6012) );
  OR2_X1 U7474 ( .A1(n9458), .A2(n9078), .ZN(n9286) );
  NAND2_X1 U7475 ( .A1(n6037), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6018) );
  INV_X1 U7476 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n6013) );
  INV_X1 U7477 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6859) );
  INV_X1 U7478 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n6014) );
  NAND4_X4 U7479 ( .A1(n6018), .A2(n6017), .A3(n6016), .A4(n6015), .ZN(n6552)
         );
  INV_X1 U7480 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6793) );
  NAND2_X1 U7481 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n6019) );
  MUX2_X1 U7482 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6019), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n6022) );
  INV_X1 U7483 ( .A(n6020), .ZN(n6021) );
  INV_X1 U7484 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n6839) );
  INV_X1 U7485 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n6833) );
  NAND2_X1 U7486 ( .A1(n6023), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n6024) );
  INV_X1 U7487 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n6836) );
  XNOR2_X1 U7488 ( .A(n6028), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n9493) );
  MUX2_X1 U7489 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9493), .S(n6117), .Z(n7238) );
  INV_X1 U7490 ( .A(n7238), .ZN(n10144) );
  NOR2_X1 U7491 ( .A1(n6027), .A2(n10144), .ZN(n6384) );
  NAND2_X1 U7492 ( .A1(n10126), .A2(n6384), .ZN(n6030) );
  INV_X1 U7493 ( .A(n6552), .ZN(n7052) );
  NAND2_X1 U7494 ( .A1(n7052), .A2(n6553), .ZN(n6029) );
  NAND2_X1 U7495 ( .A1(n6030), .A2(n6029), .ZN(n7394) );
  INV_X1 U7496 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n6031) );
  OR2_X1 U7497 ( .A1(n6032), .A2(n6031), .ZN(n6041) );
  INV_X1 U7498 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n6033) );
  INV_X1 U7499 ( .A(n6035), .ZN(n6036) );
  NAND2_X1 U7500 ( .A1(n6036), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6039) );
  NAND2_X1 U7501 ( .A1(n4486), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6038) );
  INV_X1 U7502 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6795) );
  NOR2_X1 U7503 ( .A1(n6020), .A2(n5913), .ZN(n6042) );
  MUX2_X1 U7504 ( .A(n5913), .B(n6042), .S(P1_IR_REG_2__SCAN_IN), .Z(n6043) );
  INV_X1 U7505 ( .A(n6043), .ZN(n6045) );
  NAND2_X1 U7506 ( .A1(n6045), .A2(n6044), .ZN(n6860) );
  NAND2_X1 U7507 ( .A1(n7394), .A2(n7393), .ZN(n7392) );
  INV_X1 U7508 ( .A(n9021), .ZN(n7314) );
  NAND2_X1 U7509 ( .A1(n7314), .A2(n6563), .ZN(n6499) );
  NAND2_X1 U7510 ( .A1(n6023), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n6051) );
  INV_X1 U7511 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6871) );
  OR2_X1 U7512 ( .A1(n6047), .A2(n6871), .ZN(n6050) );
  INV_X1 U7513 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6880) );
  OR2_X1 U7514 ( .A1(n6034), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n6048) );
  NAND2_X1 U7515 ( .A1(n6044), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6053) );
  INV_X1 U7516 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n6052) );
  XNOR2_X1 U7517 ( .A(n6053), .B(n6052), .ZN(n6881) );
  OR2_X1 U7518 ( .A1(n6062), .A2(n6799), .ZN(n6055) );
  INV_X1 U7519 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6794) );
  OR2_X1 U7520 ( .A1(n6352), .A2(n6794), .ZN(n6054) );
  INV_X1 U7521 ( .A(n6544), .ZN(n9020) );
  NAND2_X1 U7522 ( .A1(n9020), .A2(n6542), .ZN(n6430) );
  NAND2_X1 U7523 ( .A1(n7245), .A2(n6430), .ZN(n7242) );
  INV_X1 U7524 ( .A(n7242), .ZN(n7313) );
  NAND2_X1 U7525 ( .A1(n7311), .A2(n7245), .ZN(n6066) );
  NAND2_X1 U7526 ( .A1(n4486), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6059) );
  INV_X1 U7527 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6882) );
  OR2_X1 U7528 ( .A1(n6288), .A2(n6882), .ZN(n6058) );
  OAI21_X1 U7529 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(n6067), .ZN(n7263) );
  OR2_X1 U7530 ( .A1(n6034), .A2(n7263), .ZN(n6057) );
  NAND2_X1 U7531 ( .A1(n6023), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n6056) );
  OR2_X1 U7532 ( .A1(n6044), .A2(P1_IR_REG_3__SCAN_IN), .ZN(n6073) );
  NAND2_X1 U7533 ( .A1(n6073), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6061) );
  XNOR2_X1 U7534 ( .A(n6061), .B(n6060), .ZN(n9979) );
  INV_X1 U7535 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6806) );
  OR2_X1 U7536 ( .A1(n6352), .A2(n6806), .ZN(n6063) );
  OAI211_X1 U7537 ( .C1(n6117), .C2(n9979), .A(n6064), .B(n6063), .ZN(n7352)
         );
  NAND2_X1 U7538 ( .A1(n7539), .A2(n7352), .ZN(n6504) );
  INV_X1 U7539 ( .A(n7539), .ZN(n9369) );
  NAND2_X1 U7540 ( .A1(n9369), .A2(n6538), .ZN(n6431) );
  NAND2_X1 U7541 ( .A1(n6504), .A2(n6431), .ZN(n7537) );
  INV_X1 U7542 ( .A(n7537), .ZN(n6065) );
  NAND2_X1 U7543 ( .A1(n6066), .A2(n6065), .ZN(n7251) );
  NAND2_X1 U7544 ( .A1(n7251), .A2(n6504), .ZN(n9367) );
  NAND2_X1 U7545 ( .A1(n6276), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n6072) );
  OR2_X1 U7546 ( .A1(n6358), .A2(n10222), .ZN(n6071) );
  INV_X1 U7547 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n9373) );
  OR2_X1 U7548 ( .A1(n6288), .A2(n9373), .ZN(n6070) );
  INV_X1 U7549 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n6870) );
  NAND2_X1 U7550 ( .A1(n6067), .A2(n6870), .ZN(n6068) );
  NAND2_X1 U7551 ( .A1(n6081), .A2(n6068), .ZN(n9377) );
  OR2_X1 U7552 ( .A1(n6034), .A2(n9377), .ZN(n6069) );
  NOR2_X1 U7553 ( .A1(n6073), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n6089) );
  OR2_X1 U7554 ( .A1(n6089), .A2(n5913), .ZN(n6074) );
  INV_X1 U7555 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n6088) );
  XNOR2_X1 U7556 ( .A(n6074), .B(n6088), .ZN(n6883) );
  OR2_X1 U7557 ( .A1(n6062), .A2(n6809), .ZN(n6076) );
  INV_X1 U7558 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6810) );
  OR2_X1 U7559 ( .A1(n6352), .A2(n6810), .ZN(n6075) );
  NAND2_X1 U7560 ( .A1(n7558), .A2(n10176), .ZN(n6503) );
  INV_X1 U7561 ( .A(n6503), .ZN(n6077) );
  OR2_X2 U7562 ( .A1(n9367), .A2(n6077), .ZN(n6078) );
  INV_X1 U7563 ( .A(n7558), .ZN(n9019) );
  INV_X1 U7564 ( .A(n10176), .ZN(n9378) );
  NAND2_X1 U7565 ( .A1(n9019), .A2(n9378), .ZN(n6426) );
  INV_X1 U7566 ( .A(n7351), .ZN(n6366) );
  XNOR2_X1 U7567 ( .A(n7704), .B(n6366), .ZN(n6094) );
  NAND2_X1 U7568 ( .A1(n6276), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n6087) );
  INV_X1 U7569 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6079) );
  OR2_X1 U7570 ( .A1(n6358), .A2(n6079), .ZN(n6086) );
  INV_X1 U7571 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6080) );
  NAND2_X1 U7572 ( .A1(n6081), .A2(n6080), .ZN(n6082) );
  NAND2_X1 U7573 ( .A1(n6106), .A2(n6082), .ZN(n7556) );
  OR2_X1 U7574 ( .A1(n6235), .A2(n7556), .ZN(n6085) );
  INV_X1 U7575 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6083) );
  OR2_X1 U7576 ( .A1(n6288), .A2(n6083), .ZN(n6084) );
  NAND2_X1 U7577 ( .A1(n6089), .A2(n6088), .ZN(n6101) );
  NAND2_X1 U7578 ( .A1(n6101), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6091) );
  INV_X1 U7579 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n6090) );
  XNOR2_X1 U7580 ( .A(n6091), .B(n6090), .ZN(n6925) );
  OR2_X1 U7581 ( .A1(n6062), .A2(n6807), .ZN(n6093) );
  INV_X1 U7582 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6808) );
  OR2_X1 U7583 ( .A1(n6352), .A2(n6808), .ZN(n6092) );
  OAI211_X1 U7584 ( .C1(n6117), .C2(n6925), .A(n6093), .B(n6092), .ZN(n7701)
         );
  NAND2_X1 U7585 ( .A1(n7544), .A2(n7701), .ZN(n7527) );
  INV_X1 U7586 ( .A(n7544), .ZN(n9371) );
  INV_X1 U7587 ( .A(n7701), .ZN(n10184) );
  NAND2_X1 U7588 ( .A1(n9371), .A2(n10184), .ZN(n7525) );
  NAND2_X1 U7589 ( .A1(n7527), .A2(n7525), .ZN(n7696) );
  INV_X1 U7590 ( .A(n7696), .ZN(n7703) );
  NAND2_X1 U7591 ( .A1(n6094), .A2(n7703), .ZN(n6206) );
  NAND2_X1 U7592 ( .A1(n6276), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n6100) );
  OR2_X1 U7593 ( .A1(n6358), .A2(n10226), .ZN(n6099) );
  INV_X1 U7594 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6095) );
  NAND2_X1 U7595 ( .A1(n6108), .A2(n6095), .ZN(n6096) );
  NAND2_X1 U7596 ( .A1(n6145), .A2(n6096), .ZN(n7642) );
  OR2_X1 U7597 ( .A1(n6235), .A2(n7642), .ZN(n6098) );
  INV_X1 U7598 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n7629) );
  OR2_X1 U7599 ( .A1(n6288), .A2(n7629), .ZN(n6097) );
  OR2_X1 U7600 ( .A1(n6811), .A2(n6062), .ZN(n6104) );
  NAND2_X1 U7601 ( .A1(n6102), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6140) );
  XNOR2_X1 U7602 ( .A(n6140), .B(P1_IR_REG_8__SCAN_IN), .ZN(n6956) );
  AOI22_X1 U7603 ( .A1(n6246), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n4752), .B2(
        n6956), .ZN(n6103) );
  NAND2_X1 U7604 ( .A1(n6104), .A2(n6103), .ZN(n7777) );
  NAND2_X1 U7605 ( .A1(n7797), .A2(n7777), .ZN(n6387) );
  NAND2_X1 U7606 ( .A1(n6276), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n6112) );
  INV_X1 U7607 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6896) );
  OR2_X1 U7608 ( .A1(n6358), .A2(n6896), .ZN(n6111) );
  INV_X1 U7609 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n6903) );
  OR2_X1 U7610 ( .A1(n6288), .A2(n6903), .ZN(n6110) );
  INV_X1 U7611 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n6105) );
  NAND2_X1 U7612 ( .A1(n6106), .A2(n6105), .ZN(n6107) );
  NAND2_X1 U7613 ( .A1(n6108), .A2(n6107), .ZN(n7571) );
  OR2_X1 U7614 ( .A1(n6034), .A2(n7571), .ZN(n6109) );
  NAND2_X1 U7615 ( .A1(n6113), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6114) );
  XNOR2_X1 U7616 ( .A(n6114), .B(P1_IR_REG_7__SCAN_IN), .ZN(n9997) );
  INV_X1 U7617 ( .A(n9997), .ZN(n6796) );
  OR2_X1 U7618 ( .A1(n6800), .A2(n6062), .ZN(n6116) );
  OR2_X1 U7619 ( .A1(n6352), .A2(n9657), .ZN(n6115) );
  OAI211_X1 U7620 ( .C1(n6117), .C2(n6796), .A(n6116), .B(n6115), .ZN(n7622)
         );
  NAND2_X1 U7621 ( .A1(n7557), .A2(n7622), .ZN(n7615) );
  AND2_X1 U7622 ( .A1(n6387), .A2(n7615), .ZN(n7614) );
  AND2_X1 U7623 ( .A1(n7614), .A2(n7527), .ZN(n6119) );
  INV_X1 U7624 ( .A(n7797), .ZN(n9017) );
  NAND2_X1 U7625 ( .A1(n9017), .A2(n10199), .ZN(n7779) );
  INV_X1 U7626 ( .A(n7622), .ZN(n10192) );
  NAND2_X1 U7627 ( .A1(n9018), .A2(n10192), .ZN(n6428) );
  NAND2_X1 U7628 ( .A1(n7779), .A2(n6428), .ZN(n6118) );
  AOI22_X1 U7629 ( .A1(n6206), .A2(n6119), .B1(n6387), .B2(n6118), .ZN(n6213)
         );
  NAND2_X1 U7630 ( .A1(n6844), .A2(n6351), .ZN(n6122) );
  OR2_X1 U7631 ( .A1(n6120), .A2(n5913), .ZN(n6184) );
  XNOR2_X1 U7632 ( .A(n6184), .B(P1_IR_REG_12__SCAN_IN), .ZN(n10038) );
  AOI22_X1 U7633 ( .A1(n6246), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n4752), .B2(
        n10038), .ZN(n6121) );
  NAND2_X2 U7634 ( .A1(n6122), .A2(n6121), .ZN(n8075) );
  NAND2_X1 U7635 ( .A1(n6276), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n6128) );
  INV_X1 U7636 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n6123) );
  OR2_X1 U7637 ( .A1(n6358), .A2(n6123), .ZN(n6127) );
  INV_X1 U7638 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n8003) );
  OR2_X1 U7639 ( .A1(n6288), .A2(n8003), .ZN(n6126) );
  NAND2_X1 U7640 ( .A1(n6160), .A2(n8070), .ZN(n6124) );
  NAND2_X1 U7641 ( .A1(n6191), .A2(n6124), .ZN(n8073) );
  OR2_X1 U7642 ( .A1(n6235), .A2(n8073), .ZN(n6125) );
  NAND2_X1 U7643 ( .A1(n8075), .A2(n8082), .ZN(n8034) );
  NAND2_X1 U7644 ( .A1(n6822), .A2(n6351), .ZN(n6131) );
  NAND2_X1 U7645 ( .A1(n5985), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6129) );
  XNOR2_X1 U7646 ( .A(n6129), .B(P1_IR_REG_10__SCAN_IN), .ZN(n9025) );
  AOI22_X1 U7647 ( .A1(n6246), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n4752), .B2(
        n9025), .ZN(n6130) );
  NAND2_X1 U7648 ( .A1(n6276), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n6138) );
  INV_X1 U7649 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6132) );
  OR2_X1 U7650 ( .A1(n6358), .A2(n6132), .ZN(n6137) );
  NAND2_X1 U7651 ( .A1(n6147), .A2(n6133), .ZN(n6134) );
  NAND2_X1 U7652 ( .A1(n6158), .A2(n6134), .ZN(n7861) );
  OR2_X1 U7653 ( .A1(n6235), .A2(n7861), .ZN(n6136) );
  INV_X1 U7654 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7862) );
  OR2_X1 U7655 ( .A1(n6288), .A2(n7862), .ZN(n6135) );
  NAND2_X1 U7656 ( .A1(n7881), .A2(n7890), .ZN(n7885) );
  NAND2_X1 U7657 ( .A1(n6817), .A2(n6351), .ZN(n6144) );
  INV_X1 U7658 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n6139) );
  NAND2_X1 U7659 ( .A1(n6140), .A2(n6139), .ZN(n6141) );
  NAND2_X1 U7660 ( .A1(n6141), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6142) );
  XNOR2_X1 U7661 ( .A(n6142), .B(P1_IR_REG_9__SCAN_IN), .ZN(n10015) );
  AOI22_X1 U7662 ( .A1(n6246), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n4752), .B2(
        n10015), .ZN(n6143) );
  NAND2_X1 U7663 ( .A1(n6276), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n6151) );
  OR2_X1 U7664 ( .A1(n6358), .A2(n10229), .ZN(n6150) );
  INV_X1 U7665 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n7796) );
  NAND2_X1 U7666 ( .A1(n6145), .A2(n7796), .ZN(n6146) );
  NAND2_X1 U7667 ( .A1(n6147), .A2(n6146), .ZN(n7800) );
  OR2_X1 U7668 ( .A1(n6235), .A2(n7800), .ZN(n6149) );
  INV_X1 U7669 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n7785) );
  OR2_X1 U7670 ( .A1(n6288), .A2(n7785), .ZN(n6148) );
  NAND4_X1 U7671 ( .A1(n6151), .A2(n6150), .A3(n6149), .A4(n6148), .ZN(n9016)
         );
  INV_X1 U7672 ( .A(n9016), .ZN(n7832) );
  NAND2_X1 U7673 ( .A1(n7853), .A2(n7832), .ZN(n7848) );
  NAND2_X1 U7674 ( .A1(n7885), .A2(n7848), .ZN(n6200) );
  INV_X1 U7675 ( .A(n6200), .ZN(n6165) );
  NAND2_X1 U7676 ( .A1(n6820), .A2(n6351), .ZN(n6155) );
  OR2_X1 U7677 ( .A1(n6152), .A2(n5913), .ZN(n6153) );
  XNOR2_X1 U7678 ( .A(n6153), .B(P1_IR_REG_11__SCAN_IN), .ZN(n10026) );
  AOI22_X1 U7679 ( .A1(n6246), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n4752), .B2(
        n10026), .ZN(n6154) );
  NAND2_X1 U7680 ( .A1(n6276), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n6164) );
  INV_X1 U7681 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n6156) );
  OR2_X1 U7682 ( .A1(n6358), .A2(n6156), .ZN(n6163) );
  INV_X1 U7683 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n6157) );
  NAND2_X1 U7684 ( .A1(n6158), .A2(n6157), .ZN(n6159) );
  NAND2_X1 U7685 ( .A1(n6160), .A2(n6159), .ZN(n7940) );
  OR2_X1 U7686 ( .A1(n6235), .A2(n7940), .ZN(n6162) );
  INV_X1 U7687 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7897) );
  OR2_X1 U7688 ( .A1(n6288), .A2(n7897), .ZN(n6161) );
  NAND4_X1 U7689 ( .A1(n6164), .A2(n6163), .A3(n6162), .A4(n6161), .ZN(n9014)
         );
  XNOR2_X1 U7690 ( .A(n7986), .B(n9014), .ZN(n7889) );
  NAND4_X1 U7691 ( .A1(n8034), .A2(n6165), .A3(n7889), .A4(n7351), .ZN(n6212)
         );
  INV_X1 U7692 ( .A(n9014), .ZN(n7831) );
  OR2_X1 U7693 ( .A1(n7986), .A2(n7831), .ZN(n7993) );
  INV_X1 U7694 ( .A(n7889), .ZN(n7884) );
  NAND3_X1 U7695 ( .A1(n8032), .A2(n7884), .A3(n7351), .ZN(n6170) );
  INV_X1 U7696 ( .A(n7853), .ZN(n10208) );
  AND2_X1 U7697 ( .A1(n10208), .A2(n9016), .ZN(n7846) );
  INV_X1 U7698 ( .A(n7846), .ZN(n6436) );
  NAND3_X1 U7699 ( .A1(n6436), .A2(n7886), .A3(n7351), .ZN(n6166) );
  OAI21_X1 U7700 ( .B1(n6366), .B2(n7885), .A(n6166), .ZN(n6167) );
  NAND2_X1 U7701 ( .A1(n8032), .A2(n6167), .ZN(n6169) );
  NAND3_X1 U7702 ( .A1(n8075), .A2(n8082), .A3(n7351), .ZN(n6168) );
  AND3_X1 U7703 ( .A1(n6170), .A2(n6169), .A3(n6168), .ZN(n6205) );
  NAND2_X1 U7704 ( .A1(n6916), .A2(n6351), .ZN(n6174) );
  NAND2_X1 U7705 ( .A1(n6171), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6172) );
  XNOR2_X1 U7706 ( .A(n6172), .B(P1_IR_REG_14__SCAN_IN), .ZN(n10064) );
  AOI22_X1 U7707 ( .A1(n6246), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n4752), .B2(
        n10064), .ZN(n6173) );
  NAND2_X2 U7708 ( .A1(n6174), .A2(n6173), .ZN(n9463) );
  NAND2_X1 U7709 ( .A1(n6276), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n6182) );
  INV_X1 U7710 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n6175) );
  OR2_X1 U7711 ( .A1(n6358), .A2(n6175), .ZN(n6181) );
  NAND2_X1 U7712 ( .A1(n6193), .A2(n6176), .ZN(n6177) );
  NAND2_X1 U7713 ( .A1(n6219), .A2(n6177), .ZN(n9351) );
  OR2_X1 U7714 ( .A1(n6235), .A2(n9351), .ZN(n6180) );
  INV_X1 U7715 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n6178) );
  OR2_X1 U7716 ( .A1(n6288), .A2(n6178), .ZN(n6179) );
  NAND4_X1 U7717 ( .A1(n6182), .A2(n6181), .A3(n6180), .A4(n6179), .ZN(n9073)
         );
  INV_X1 U7718 ( .A(n9073), .ZN(n6198) );
  NAND2_X1 U7719 ( .A1(n6891), .A2(n6351), .ZN(n6188) );
  NAND2_X1 U7720 ( .A1(n6184), .A2(n6183), .ZN(n6185) );
  NAND2_X1 U7721 ( .A1(n6185), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6186) );
  XNOR2_X1 U7722 ( .A(n6186), .B(P1_IR_REG_13__SCAN_IN), .ZN(n9039) );
  AOI22_X1 U7723 ( .A1(n6246), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n4752), .B2(
        n9039), .ZN(n6187) );
  NAND2_X1 U7724 ( .A1(n6276), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n6197) );
  INV_X1 U7725 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n6189) );
  OR2_X1 U7726 ( .A1(n6358), .A2(n6189), .ZN(n6196) );
  INV_X1 U7727 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n6190) );
  NAND2_X1 U7728 ( .A1(n6191), .A2(n6190), .ZN(n6192) );
  NAND2_X1 U7729 ( .A1(n6193), .A2(n6192), .ZN(n8085) );
  OR2_X1 U7730 ( .A1(n6235), .A2(n8085), .ZN(n6195) );
  INV_X1 U7731 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n8043) );
  OR2_X1 U7732 ( .A1(n6288), .A2(n8043), .ZN(n6194) );
  NAND4_X1 U7733 ( .A1(n6197), .A2(n6196), .A3(n6195), .A4(n6194), .ZN(n9070)
         );
  INV_X1 U7734 ( .A(n9070), .ZN(n6199) );
  OR2_X1 U7735 ( .A1(n9932), .A2(n6199), .ZN(n6392) );
  NAND2_X1 U7736 ( .A1(n9104), .A2(n6392), .ZN(n6442) );
  NAND2_X1 U7737 ( .A1(n9463), .A2(n6198), .ZN(n6383) );
  NAND2_X1 U7738 ( .A1(n9932), .A2(n6199), .ZN(n9103) );
  NAND2_X1 U7739 ( .A1(n6383), .A2(n9103), .ZN(n6418) );
  AND2_X1 U7740 ( .A1(n6200), .A2(n7886), .ZN(n6419) );
  NAND3_X1 U7741 ( .A1(n6389), .A2(n6419), .A3(n7889), .ZN(n6203) );
  NAND2_X1 U7742 ( .A1(n7986), .A2(n7831), .ZN(n7991) );
  INV_X1 U7743 ( .A(n7991), .ZN(n6201) );
  NAND2_X1 U7744 ( .A1(n6389), .A2(n6201), .ZN(n6202) );
  NAND4_X1 U7745 ( .A1(n6203), .A2(n6202), .A3(n6366), .A4(n8034), .ZN(n6204)
         );
  OAI22_X1 U7746 ( .A1(n6205), .A2(n6442), .B1(n6418), .B2(n6204), .ZN(n6211)
         );
  AND2_X1 U7747 ( .A1(n6428), .A2(n7525), .ZN(n6425) );
  NAND2_X1 U7748 ( .A1(n6206), .A2(n6425), .ZN(n6207) );
  NAND2_X1 U7749 ( .A1(n6207), .A2(n7614), .ZN(n6209) );
  AND4_X1 U7750 ( .A1(n6436), .A2(n7886), .A3(n6366), .A4(n7779), .ZN(n6208)
         );
  NAND4_X1 U7751 ( .A1(n6209), .A2(n6208), .A3(n7889), .A4(n6389), .ZN(n6210)
         );
  OAI211_X1 U7752 ( .C1(n6213), .C2(n6212), .A(n6211), .B(n6210), .ZN(n6228)
         );
  NAND2_X1 U7753 ( .A1(n7039), .A2(n6351), .ZN(n6217) );
  NAND2_X1 U7754 ( .A1(n6214), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6215) );
  XNOR2_X1 U7755 ( .A(n6215), .B(P1_IR_REG_15__SCAN_IN), .ZN(n10077) );
  AOI22_X1 U7756 ( .A1(n6246), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n4752), .B2(
        n10077), .ZN(n6216) );
  NAND2_X1 U7757 ( .A1(n6276), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n6225) );
  NAND2_X1 U7758 ( .A1(n6219), .A2(n6218), .ZN(n6220) );
  NAND2_X1 U7759 ( .A1(n6234), .A2(n6220), .ZN(n9336) );
  OR2_X1 U7760 ( .A1(n6235), .A2(n9336), .ZN(n6224) );
  INV_X1 U7761 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n6221) );
  OR2_X1 U7762 ( .A1(n6358), .A2(n6221), .ZN(n6223) );
  INV_X1 U7763 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9337) );
  OR2_X1 U7764 ( .A1(n6288), .A2(n9337), .ZN(n6222) );
  NAND2_X1 U7765 ( .A1(n9925), .A2(n8932), .ZN(n9105) );
  NAND2_X1 U7766 ( .A1(n6442), .A2(n6383), .ZN(n6226) );
  NAND2_X1 U7767 ( .A1(n6418), .A2(n9104), .ZN(n6440) );
  MUX2_X1 U7768 ( .A(n6226), .B(n6440), .S(n7351), .Z(n6227) );
  NAND3_X1 U7769 ( .A1(n6228), .A2(n9330), .A3(n6227), .ZN(n6241) );
  NAND2_X1 U7770 ( .A1(n7136), .A2(n6351), .ZN(n6231) );
  XNOR2_X1 U7771 ( .A(n6229), .B(P1_IR_REG_16__SCAN_IN), .ZN(n10089) );
  AOI22_X1 U7772 ( .A1(n6246), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n4752), .B2(
        n10089), .ZN(n6230) );
  NAND2_X1 U7773 ( .A1(n6276), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n6239) );
  INV_X1 U7774 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n6232) );
  OR2_X1 U7775 ( .A1(n6358), .A2(n6232), .ZN(n6238) );
  XNOR2_X1 U7776 ( .A(n6234), .B(n6233), .ZN(n9320) );
  OR2_X1 U7777 ( .A1(n6235), .A2(n9320), .ZN(n6237) );
  INV_X1 U7778 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n9321) );
  OR2_X1 U7779 ( .A1(n6288), .A2(n9321), .ZN(n6236) );
  OR2_X1 U7780 ( .A1(n9323), .A2(n9012), .ZN(n6435) );
  NAND2_X1 U7781 ( .A1(n9323), .A2(n9012), .ZN(n9106) );
  MUX2_X1 U7782 ( .A(n9310), .B(n9105), .S(n6366), .Z(n6240) );
  NAND3_X1 U7783 ( .A1(n6241), .A2(n9317), .A3(n6240), .ZN(n6243) );
  AND2_X1 U7784 ( .A1(n9286), .A2(n9109), .ZN(n9304) );
  MUX2_X1 U7785 ( .A(n6435), .B(n9106), .S(n7351), .Z(n6242) );
  NAND3_X1 U7786 ( .A1(n6243), .A2(n9304), .A3(n6242), .ZN(n6244) );
  NAND2_X1 U7787 ( .A1(n6245), .A2(n6244), .ZN(n6268) );
  NAND2_X1 U7788 ( .A1(n7325), .A2(n6351), .ZN(n6248) );
  AOI22_X1 U7789 ( .A1(n6246), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n10138), 
        .B2(n4752), .ZN(n6247) );
  NAND2_X1 U7790 ( .A1(n6249), .A2(n8906), .ZN(n6250) );
  AND2_X1 U7791 ( .A1(n6260), .A2(n6250), .ZN(n9270) );
  NAND2_X1 U7792 ( .A1(n6346), .A2(n9270), .ZN(n6256) );
  INV_X1 U7793 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n6251) );
  OR2_X1 U7794 ( .A1(n6032), .A2(n6251), .ZN(n6255) );
  INV_X1 U7795 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9048) );
  OR2_X1 U7796 ( .A1(n6358), .A2(n9048), .ZN(n6254) );
  INV_X1 U7797 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n6252) );
  OR2_X1 U7798 ( .A1(n6288), .A2(n6252), .ZN(n6253) );
  NAND4_X1 U7799 ( .A1(n6256), .A2(n6255), .A3(n6254), .A4(n6253), .ZN(n9290)
         );
  INV_X1 U7800 ( .A(n9290), .ZN(n9080) );
  OR2_X1 U7801 ( .A1(n9447), .A2(n9080), .ZN(n6381) );
  NAND3_X1 U7802 ( .A1(n6268), .A2(n6381), .A3(n6382), .ZN(n6267) );
  NAND2_X1 U7803 ( .A1(n7490), .A2(n6351), .ZN(n6258) );
  OR2_X1 U7804 ( .A1(n6352), .A2(n9793), .ZN(n6257) );
  INV_X1 U7805 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n6259) );
  NAND2_X1 U7806 ( .A1(n6260), .A2(n6259), .ZN(n6261) );
  NAND2_X1 U7807 ( .A1(n6274), .A2(n6261), .ZN(n8958) );
  OR2_X1 U7808 ( .A1(n8958), .A2(n6235), .ZN(n6265) );
  NAND2_X1 U7809 ( .A1(n4487), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n6264) );
  NAND2_X1 U7810 ( .A1(n6036), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n6263) );
  NAND2_X1 U7811 ( .A1(n6276), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n6262) );
  NAND4_X1 U7812 ( .A1(n6265), .A2(n6264), .A3(n6263), .A4(n6262), .ZN(n9276)
         );
  INV_X1 U7813 ( .A(n9276), .ZN(n9082) );
  INV_X1 U7814 ( .A(n9115), .ZN(n6266) );
  NAND2_X1 U7815 ( .A1(n9447), .A2(n9080), .ZN(n9113) );
  NAND3_X1 U7816 ( .A1(n6267), .A2(n6266), .A3(n9113), .ZN(n6271) );
  AND2_X1 U7817 ( .A1(n9114), .A2(n6381), .ZN(n6405) );
  AND2_X1 U7818 ( .A1(n9113), .A2(n9110), .ZN(n6406) );
  NAND2_X1 U7819 ( .A1(n6268), .A2(n6406), .ZN(n6269) );
  NAND2_X1 U7820 ( .A1(n6405), .A2(n6269), .ZN(n6270) );
  NAND2_X1 U7821 ( .A1(n7575), .A2(n6351), .ZN(n6273) );
  OR2_X1 U7822 ( .A1(n6352), .A2(n7576), .ZN(n6272) );
  NAND2_X1 U7823 ( .A1(n6274), .A2(n8914), .ZN(n6275) );
  AND2_X1 U7824 ( .A1(n6283), .A2(n6275), .ZN(n9249) );
  NAND2_X1 U7825 ( .A1(n9249), .A2(n6346), .ZN(n6279) );
  AOI22_X1 U7826 ( .A1(n4486), .A2(P1_REG1_REG_21__SCAN_IN), .B1(n6276), .B2(
        P1_REG0_REG_21__SCAN_IN), .ZN(n6278) );
  NAND2_X1 U7827 ( .A1(n6036), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n6277) );
  NAND2_X1 U7828 ( .A1(n9439), .A2(n9235), .ZN(n6416) );
  INV_X1 U7829 ( .A(n6416), .ZN(n9116) );
  AOI21_X1 U7830 ( .B1(n6291), .B2(n9114), .A(n9116), .ZN(n6289) );
  NAND2_X1 U7831 ( .A1(n7658), .A2(n6351), .ZN(n6281) );
  OR2_X1 U7832 ( .A1(n6352), .A2(n7659), .ZN(n6280) );
  INV_X1 U7833 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n9227) );
  INV_X1 U7834 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n6282) );
  NAND2_X1 U7835 ( .A1(n6283), .A2(n6282), .ZN(n6284) );
  NAND2_X1 U7836 ( .A1(n6285), .A2(n6284), .ZN(n9228) );
  OR2_X1 U7837 ( .A1(n9228), .A2(n6235), .ZN(n6287) );
  AOI22_X1 U7838 ( .A1(n4487), .A2(P1_REG1_REG_22__SCAN_IN), .B1(n6276), .B2(
        P1_REG0_REG_22__SCAN_IN), .ZN(n6286) );
  OAI211_X1 U7839 ( .C1(n6288), .C2(n9227), .A(n6287), .B(n6286), .ZN(n9083)
         );
  NAND2_X1 U7840 ( .A1(n9226), .A2(n9083), .ZN(n6379) );
  NAND2_X1 U7841 ( .A1(n6379), .A2(n6378), .ZN(n6412) );
  INV_X1 U7842 ( .A(n9083), .ZN(n9084) );
  NAND2_X1 U7843 ( .A1(n9432), .A2(n9084), .ZN(n9117) );
  OAI21_X1 U7844 ( .B1(n6289), .B2(n6412), .A(n9117), .ZN(n6294) );
  NAND2_X1 U7845 ( .A1(n6378), .A2(n9115), .ZN(n6415) );
  NAND3_X1 U7846 ( .A1(n9117), .A2(n6416), .A3(n6415), .ZN(n6290) );
  NAND2_X1 U7847 ( .A1(n6290), .A2(n6379), .ZN(n6410) );
  OAI21_X1 U7848 ( .B1(n6291), .B2(n6412), .A(n6410), .ZN(n6292) );
  INV_X1 U7849 ( .A(n6292), .ZN(n6293) );
  INV_X1 U7850 ( .A(n6295), .ZN(n6515) );
  NAND4_X1 U7851 ( .A1(n6296), .A2(n6515), .A3(n6450), .A4(n6413), .ZN(n6297)
         );
  INV_X1 U7852 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n8992) );
  NAND2_X1 U7853 ( .A1(n6298), .A2(n8992), .ZN(n6299) );
  NAND2_X1 U7854 ( .A1(n6332), .A2(n6299), .ZN(n9177) );
  INV_X1 U7855 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n6302) );
  NAND2_X1 U7856 ( .A1(n6023), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n6301) );
  NAND2_X1 U7857 ( .A1(n6036), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n6300) );
  OAI211_X1 U7858 ( .C1(n6358), .C2(n6302), .A(n6301), .B(n6300), .ZN(n6303)
         );
  INV_X1 U7859 ( .A(n6303), .ZN(n6304) );
  NOR2_X1 U7860 ( .A1(n6325), .A2(n9165), .ZN(n6308) );
  NAND2_X1 U7861 ( .A1(n8060), .A2(n6351), .ZN(n6307) );
  OR2_X1 U7862 ( .A1(n6352), .A2(n9681), .ZN(n6306) );
  OR2_X1 U7863 ( .A1(n6376), .A2(n9165), .ZN(n6309) );
  MUX2_X1 U7864 ( .A(n6309), .B(n9093), .S(n6366), .Z(n6311) );
  INV_X1 U7865 ( .A(n9120), .ZN(n6321) );
  NAND3_X1 U7866 ( .A1(n6321), .A2(n9094), .A3(n6366), .ZN(n6310) );
  NAND2_X1 U7867 ( .A1(n6311), .A2(n6310), .ZN(n6327) );
  NAND2_X1 U7868 ( .A1(n6312), .A2(n6351), .ZN(n6314) );
  OR2_X1 U7869 ( .A1(n6352), .A2(n9863), .ZN(n6313) );
  XNOR2_X1 U7870 ( .A(n6332), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n9160) );
  NAND2_X1 U7871 ( .A1(n9160), .A2(n6346), .ZN(n6320) );
  INV_X1 U7872 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n6317) );
  NAND2_X1 U7873 ( .A1(n6036), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n6316) );
  NAND2_X1 U7874 ( .A1(n6276), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6315) );
  OAI211_X1 U7875 ( .C1(n6358), .C2(n6317), .A(n6316), .B(n6315), .ZN(n6318)
         );
  INV_X1 U7876 ( .A(n6318), .ZN(n6319) );
  NAND2_X1 U7877 ( .A1(n9405), .A2(n9095), .ZN(n6457) );
  OAI21_X1 U7878 ( .B1(n6321), .B2(n9094), .A(n6457), .ZN(n6323) );
  OAI21_X1 U7879 ( .B1(n9121), .B2(n9093), .A(n9124), .ZN(n6322) );
  MUX2_X1 U7880 ( .A(n6323), .B(n6322), .S(n7351), .Z(n6324) );
  OAI21_X1 U7881 ( .B1(n6325), .B2(n9164), .A(n6324), .ZN(n6326) );
  NAND2_X1 U7882 ( .A1(n8150), .A2(n6351), .ZN(n6329) );
  OR2_X1 U7883 ( .A1(n6352), .A2(n9866), .ZN(n6328) );
  INV_X1 U7884 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n8882) );
  INV_X1 U7885 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n6330) );
  OAI21_X1 U7886 ( .B1(n6332), .B2(n8882), .A(n6330), .ZN(n6333) );
  NAND2_X1 U7887 ( .A1(P1_REG3_REG_28__SCAN_IN), .A2(P1_REG3_REG_27__SCAN_IN), 
        .ZN(n6331) );
  INV_X1 U7888 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n6336) );
  NAND2_X1 U7889 ( .A1(n6036), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n6335) );
  NAND2_X1 U7890 ( .A1(n6276), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6334) );
  OAI211_X1 U7891 ( .C1(n6358), .C2(n6336), .A(n6335), .B(n6334), .ZN(n6337)
         );
  INV_X1 U7892 ( .A(n9148), .ZN(n6339) );
  MUX2_X1 U7893 ( .A(n9124), .B(n6457), .S(n7351), .Z(n6338) );
  MUX2_X1 U7894 ( .A(n9126), .B(n6403), .S(n7351), .Z(n6340) );
  INV_X1 U7895 ( .A(n6341), .ZN(n9135) );
  INV_X1 U7896 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n6344) );
  NAND2_X1 U7897 ( .A1(n6276), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6343) );
  NAND2_X1 U7898 ( .A1(n6036), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6342) );
  OAI211_X1 U7899 ( .C1(n6358), .C2(n6344), .A(n6343), .B(n6342), .ZN(n6345)
         );
  AOI21_X1 U7900 ( .B1(n9135), .B2(n6346), .A(n6345), .ZN(n6775) );
  INV_X1 U7901 ( .A(n6775), .ZN(n9151) );
  AOI21_X1 U7902 ( .B1(n6360), .B2(n9151), .A(n6366), .ZN(n6350) );
  NOR2_X1 U7903 ( .A1(n6360), .A2(n9151), .ZN(n6349) );
  NAND2_X1 U7904 ( .A1(n8872), .A2(n6351), .ZN(n6348) );
  INV_X1 U7905 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n9598) );
  OR2_X1 U7906 ( .A1(n6352), .A2(n9598), .ZN(n6347) );
  INV_X1 U7907 ( .A(n9134), .ZN(n9394) );
  NAND2_X1 U7908 ( .A1(n8136), .A2(n6351), .ZN(n6354) );
  INV_X1 U7909 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n9807) );
  OR2_X1 U7910 ( .A1(n6352), .A2(n9807), .ZN(n6353) );
  INV_X1 U7911 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n6357) );
  NAND2_X1 U7912 ( .A1(n6036), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n6356) );
  NAND2_X1 U7913 ( .A1(n6276), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n6355) );
  OAI211_X1 U7914 ( .C1(n6358), .C2(n6357), .A(n6356), .B(n6355), .ZN(n9129)
         );
  INV_X1 U7915 ( .A(n9129), .ZN(n6401) );
  OR2_X1 U7916 ( .A1(n9388), .A2(n6523), .ZN(n6359) );
  INV_X1 U7917 ( .A(n6360), .ZN(n6361) );
  NAND3_X1 U7918 ( .A1(n6361), .A2(n6366), .A3(n9151), .ZN(n6362) );
  INV_X1 U7919 ( .A(n6363), .ZN(n9061) );
  NAND2_X1 U7920 ( .A1(n9129), .A2(n9061), .ZN(n6364) );
  NAND2_X1 U7921 ( .A1(n9064), .A2(n6364), .ZN(n6462) );
  INV_X1 U7922 ( .A(n6466), .ZN(n6367) );
  INV_X1 U7923 ( .A(n6464), .ZN(n6373) );
  NOR2_X1 U7924 ( .A1(n7246), .A2(n7577), .ZN(n6372) );
  NAND2_X1 U7925 ( .A1(n6373), .A2(n6372), .ZN(n6374) );
  INV_X1 U7926 ( .A(n6375), .ZN(n6526) );
  INV_X1 U7927 ( .A(n6523), .ZN(n6400) );
  INV_X1 U7928 ( .A(n9099), .ZN(n9127) );
  NAND2_X1 U7929 ( .A1(n9411), .A2(n9093), .ZN(n9122) );
  INV_X1 U7930 ( .A(n9122), .ZN(n6455) );
  NAND2_X1 U7931 ( .A1(n6413), .A2(n6377), .ZN(n9212) );
  NAND2_X1 U7932 ( .A1(n6379), .A2(n9117), .ZN(n9232) );
  INV_X1 U7933 ( .A(n9114), .ZN(n6380) );
  OR2_X1 U7934 ( .A1(n6380), .A2(n9115), .ZN(n9263) );
  NAND2_X1 U7935 ( .A1(n6381), .A2(n9113), .ZN(n9273) );
  NAND2_X1 U7936 ( .A1(n6382), .A2(n9110), .ZN(n9288) );
  NAND2_X1 U7937 ( .A1(n9104), .A2(n6383), .ZN(n9357) );
  INV_X1 U7938 ( .A(n9380), .ZN(n6385) );
  INV_X1 U7939 ( .A(n6384), .ZN(n10127) );
  NAND2_X1 U7940 ( .A1(n6027), .A2(n10144), .ZN(n6497) );
  NAND2_X1 U7941 ( .A1(n10127), .A2(n6497), .ZN(n6976) );
  NOR4_X1 U7942 ( .A1(n6385), .A2(n6976), .A3(n7537), .A4(n7242), .ZN(n6386)
         );
  NAND4_X1 U7943 ( .A1(n6386), .A2(n7703), .A3(n7393), .A4(n10126), .ZN(n6388)
         );
  NAND2_X1 U7944 ( .A1(n6387), .A2(n7779), .ZN(n7626) );
  NAND2_X1 U7945 ( .A1(n7615), .A2(n6428), .ZN(n7624) );
  NOR3_X1 U7946 ( .A1(n6388), .A2(n7626), .A3(n7624), .ZN(n6391) );
  INV_X1 U7947 ( .A(n7848), .ZN(n6390) );
  NOR2_X1 U7948 ( .A1(n7846), .A2(n6390), .ZN(n7781) );
  NAND4_X1 U7949 ( .A1(n6391), .A2(n7994), .A3(n7860), .A4(n7781), .ZN(n6393)
         );
  INV_X1 U7950 ( .A(n9101), .ZN(n8036) );
  NOR4_X1 U7951 ( .A1(n9357), .A2(n6393), .A3(n8036), .A4(n7884), .ZN(n6394)
         );
  NAND4_X1 U7952 ( .A1(n9304), .A2(n9317), .A3(n9330), .A4(n6394), .ZN(n6395)
         );
  OR4_X1 U7953 ( .A1(n9263), .A2(n9273), .A3(n9288), .A4(n6395), .ZN(n6396) );
  NOR4_X1 U7954 ( .A1(n9212), .A2(n9244), .A3(n9232), .A4(n6396), .ZN(n6397)
         );
  NAND3_X1 U7955 ( .A1(n9172), .A2(n9197), .A3(n6397), .ZN(n6398) );
  OR4_X1 U7956 ( .A1(n9148), .A2(n9164), .A3(n9188), .A4(n6398), .ZN(n6399) );
  NOR4_X1 U7957 ( .A1(n6526), .A2(n6400), .A3(n9127), .A4(n6399), .ZN(n6402)
         );
  AOI21_X1 U7958 ( .B1(n6401), .B2(n9064), .A(n6464), .ZN(n6528) );
  AOI21_X1 U7959 ( .B1(n6402), .B2(n6528), .A(n7247), .ZN(n6491) );
  INV_X1 U7960 ( .A(n6403), .ZN(n9125) );
  OR2_X1 U7961 ( .A1(n6404), .A2(n9125), .ZN(n6521) );
  INV_X1 U7962 ( .A(n9123), .ZN(n6454) );
  INV_X1 U7963 ( .A(n6405), .ZN(n6409) );
  INV_X1 U7964 ( .A(n6406), .ZN(n6407) );
  NOR2_X1 U7965 ( .A1(n6407), .A2(n9112), .ZN(n6408) );
  OR2_X1 U7966 ( .A1(n6409), .A2(n6408), .ZN(n6411) );
  OAI21_X1 U7967 ( .B1(n6412), .B2(n6411), .A(n6410), .ZN(n6414) );
  AND2_X1 U7968 ( .A1(n6414), .A2(n6413), .ZN(n6495) );
  NAND4_X1 U7969 ( .A1(n9117), .A2(n6416), .A3(n9113), .A4(n6415), .ZN(n6514)
         );
  INV_X1 U7970 ( .A(n6514), .ZN(n6448) );
  AND2_X1 U7971 ( .A1(n9109), .A2(n9106), .ZN(n6417) );
  NAND2_X1 U7972 ( .A1(n9110), .A2(n6417), .ZN(n6444) );
  OR2_X1 U7973 ( .A1(n6444), .A2(n6418), .ZN(n6512) );
  INV_X1 U7974 ( .A(n6419), .ZN(n6420) );
  AND2_X1 U7975 ( .A1(n6420), .A2(n7991), .ZN(n6421) );
  AND2_X1 U7976 ( .A1(n8034), .A2(n6421), .ZN(n6508) );
  NAND2_X1 U7977 ( .A1(n6504), .A2(n7245), .ZN(n6422) );
  NAND3_X1 U7978 ( .A1(n6422), .A2(n6431), .A3(n6426), .ZN(n6423) );
  NAND3_X1 U7979 ( .A1(n6423), .A2(n7527), .A3(n6503), .ZN(n6424) );
  AOI21_X1 U7980 ( .B1(n6425), .B2(n6424), .A(n4932), .ZN(n6434) );
  NAND2_X1 U7981 ( .A1(n7525), .A2(n6426), .ZN(n6427) );
  NAND2_X1 U7982 ( .A1(n7527), .A2(n6427), .ZN(n6429) );
  NAND2_X1 U7983 ( .A1(n6429), .A2(n6428), .ZN(n6509) );
  NAND2_X1 U7984 ( .A1(n6431), .A2(n6430), .ZN(n6502) );
  NOR2_X1 U7985 ( .A1(n6509), .A2(n6502), .ZN(n6432) );
  NAND2_X1 U7986 ( .A1(n7312), .A2(n6432), .ZN(n6433) );
  NAND4_X1 U7987 ( .A1(n9105), .A2(n6508), .A3(n6434), .A4(n6433), .ZN(n6446)
         );
  AND2_X1 U7988 ( .A1(n6435), .A2(n9310), .ZN(n9108) );
  INV_X1 U7989 ( .A(n8034), .ZN(n6439) );
  NAND3_X1 U7990 ( .A1(n6436), .A2(n7886), .A3(n7779), .ZN(n6437) );
  NAND2_X1 U7991 ( .A1(n6508), .A2(n6437), .ZN(n6438) );
  OAI21_X1 U7992 ( .B1(n8032), .B2(n6439), .A(n6438), .ZN(n6441) );
  OAI211_X1 U7993 ( .C1(n6442), .C2(n6441), .A(n6440), .B(n9105), .ZN(n6443)
         );
  AND2_X1 U7994 ( .A1(n9108), .A2(n6443), .ZN(n6445) );
  OR2_X1 U7995 ( .A1(n6445), .A2(n6444), .ZN(n6496) );
  OAI21_X1 U7996 ( .B1(n6512), .B2(n6446), .A(n6496), .ZN(n6447) );
  NAND2_X1 U7997 ( .A1(n6448), .A2(n6447), .ZN(n6449) );
  NAND3_X1 U7998 ( .A1(n6450), .A2(n6495), .A3(n6449), .ZN(n6451) );
  NAND2_X1 U7999 ( .A1(n6452), .A2(n6451), .ZN(n6453) );
  NAND4_X1 U8000 ( .A1(n9124), .A2(n9120), .A3(n6454), .A4(n6453), .ZN(n6463)
         );
  NAND2_X1 U8001 ( .A1(n9124), .A2(n6455), .ZN(n6456) );
  AND3_X1 U8002 ( .A1(n9126), .A2(n6457), .A3(n6456), .ZN(n6458) );
  OR2_X1 U8003 ( .A1(n6521), .A2(n6458), .ZN(n6461) );
  INV_X1 U8004 ( .A(n6459), .ZN(n6460) );
  OAI211_X1 U8005 ( .C1(n6521), .C2(n6463), .A(n6522), .B(n6462), .ZN(n6465)
         );
  AOI211_X1 U8006 ( .C1(n6466), .C2(n6465), .A(n7577), .B(n6464), .ZN(n6467)
         );
  NOR3_X1 U8007 ( .A1(n6491), .A2(n10138), .A3(n6467), .ZN(n6489) );
  NAND2_X1 U8008 ( .A1(n4571), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6469) );
  XNOR2_X1 U8009 ( .A(n6469), .B(n6468), .ZN(n6789) );
  OR2_X1 U8010 ( .A1(n6789), .A2(P1_U3084), .ZN(n7712) );
  INV_X1 U8011 ( .A(n7712), .ZN(n6488) );
  INV_X1 U8012 ( .A(P1_B_REG_SCAN_IN), .ZN(n6487) );
  NAND2_X1 U8013 ( .A1(n6471), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6473) );
  INV_X1 U8014 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n6472) );
  XNOR2_X1 U8015 ( .A(n6473), .B(n6472), .ZN(n7919) );
  NOR2_X1 U8016 ( .A1(n7952), .A2(n7919), .ZN(n6478) );
  NAND2_X1 U8017 ( .A1(n6475), .A2(n6474), .ZN(n6476) );
  NAND2_X1 U8018 ( .A1(n6476), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6477) );
  AND2_X1 U8019 ( .A1(n6789), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6479) );
  NAND2_X1 U8020 ( .A1(n6788), .A2(n6479), .ZN(n6951) );
  NAND2_X1 U8021 ( .A1(n6482), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6483) );
  MUX2_X1 U8022 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6483), .S(
        P1_IR_REG_20__SCAN_IN), .Z(n6485) );
  NAND2_X1 U8023 ( .A1(n6485), .A2(n6484), .ZN(n7524) );
  OR2_X1 U8024 ( .A1(n6539), .A2(n7266), .ZN(n7547) );
  NOR4_X1 U8025 ( .A1(n6951), .A2(n8151), .A3(n6481), .A4(n7547), .ZN(n6486)
         );
  AOI211_X1 U8026 ( .C1(n6488), .C2(n7660), .A(n6487), .B(n6486), .ZN(n6529)
         );
  NOR4_X1 U8027 ( .A1(n6490), .A2(n6489), .A3(n6529), .A4(n7524), .ZN(n6536)
         );
  AND2_X1 U8028 ( .A1(n7246), .A2(n7247), .ZN(n6790) );
  AOI21_X1 U8029 ( .B1(n6492), .B2(n6790), .A(n6491), .ZN(n6493) );
  INV_X1 U8030 ( .A(n6529), .ZN(n6531) );
  INV_X1 U8031 ( .A(n6494), .ZN(n6519) );
  OAI21_X1 U8032 ( .B1(n6514), .B2(n6496), .A(n6495), .ZN(n6517) );
  INV_X1 U8033 ( .A(n9105), .ZN(n6513) );
  AOI21_X1 U8034 ( .B1(n6552), .B2(n10160), .A(n7577), .ZN(n6498) );
  AOI21_X1 U8035 ( .B1(n6498), .B2(n6497), .A(n7394), .ZN(n6501) );
  NOR2_X1 U8036 ( .A1(n7314), .A2(n6563), .ZN(n6500) );
  OAI211_X1 U8037 ( .C1(n6501), .C2(n6500), .A(n7245), .B(n6499), .ZN(n6507)
         );
  INV_X1 U8038 ( .A(n6502), .ZN(n6506) );
  NAND3_X1 U8039 ( .A1(n7527), .A2(n6504), .A3(n6503), .ZN(n6505) );
  AOI21_X1 U8040 ( .B1(n6507), .B2(n6506), .A(n6505), .ZN(n6510) );
  OAI211_X1 U8041 ( .C1(n6510), .C2(n6509), .A(n6508), .B(n7614), .ZN(n6511)
         );
  NOR4_X1 U8042 ( .A1(n6514), .A2(n6513), .A3(n6512), .A4(n6511), .ZN(n6516)
         );
  OAI21_X1 U8043 ( .B1(n6517), .B2(n6516), .A(n6515), .ZN(n6518) );
  AOI21_X1 U8044 ( .B1(n6519), .B2(n6518), .A(n9121), .ZN(n6520) );
  NOR4_X1 U8045 ( .A1(n6521), .A2(n9123), .A3(n6520), .A4(n9164), .ZN(n6525)
         );
  INV_X1 U8046 ( .A(n6522), .ZN(n6524) );
  OAI21_X1 U8047 ( .B1(n6525), .B2(n6524), .A(n6523), .ZN(n6527) );
  AOI21_X1 U8048 ( .B1(n6528), .B2(n6527), .A(n6526), .ZN(n6532) );
  NAND2_X1 U8049 ( .A1(n7524), .A2(n9203), .ZN(n6768) );
  NOR3_X1 U8050 ( .A1(n6532), .A2(n6529), .A3(n6768), .ZN(n6530) );
  AOI21_X1 U8051 ( .B1(n7712), .B2(n6531), .A(n6530), .ZN(n6534) );
  NAND4_X1 U8052 ( .A1(n6532), .A2(n10138), .A3(n6531), .A4(n7524), .ZN(n6533)
         );
  NAND2_X1 U8053 ( .A1(n6534), .A2(n6533), .ZN(n6535) );
  INV_X1 U8054 ( .A(n7266), .ZN(n6537) );
  INV_X1 U8055 ( .A(n6768), .ZN(n7259) );
  NAND2_X1 U8056 ( .A1(n7660), .A2(n7259), .ZN(n6541) );
  AND2_X4 U8057 ( .A1(n6759), .A2(n6541), .ZN(n6565) );
  XNOR2_X1 U8058 ( .A(n6577), .B(n6578), .ZN(n7206) );
  INV_X1 U8059 ( .A(n6575), .ZN(n6545) );
  OAI22_X1 U8060 ( .A1(n6544), .A2(n6755), .B1(n6542), .B2(n6727), .ZN(n6574)
         );
  NOR2_X1 U8061 ( .A1(n6788), .A2(n6836), .ZN(n6546) );
  AOI21_X1 U8062 ( .B1(n7238), .B2(n6759), .A(n6546), .ZN(n6547) );
  NAND2_X1 U8063 ( .A1(n6548), .A2(n6547), .ZN(n6948) );
  INV_X1 U8064 ( .A(n6788), .ZN(n6549) );
  AOI22_X1 U8065 ( .A1(n7238), .A2(n6608), .B1(P1_IR_REG_0__SCAN_IN), .B2(
        n6549), .ZN(n6550) );
  NAND2_X1 U8066 ( .A1(n6949), .A2(n6948), .ZN(n6947) );
  NAND2_X1 U8067 ( .A1(n6552), .A2(n6608), .ZN(n6555) );
  NAND2_X1 U8068 ( .A1(n6552), .A2(n6565), .ZN(n6558) );
  NAND2_X1 U8069 ( .A1(n6553), .A2(n6608), .ZN(n6557) );
  NAND2_X1 U8070 ( .A1(n6558), .A2(n6557), .ZN(n8141) );
  INV_X1 U8071 ( .A(n8140), .ZN(n6559) );
  NAND2_X1 U8072 ( .A1(n9021), .A2(n6608), .ZN(n6561) );
  NAND2_X1 U8073 ( .A1(n6563), .A2(n6759), .ZN(n6560) );
  NAND2_X1 U8074 ( .A1(n6561), .A2(n6560), .ZN(n6562) );
  XNOR2_X1 U8075 ( .A(n6562), .B(n6712), .ZN(n6566) );
  AND2_X1 U8076 ( .A1(n6563), .A2(n6608), .ZN(n6564) );
  AOI21_X1 U8077 ( .B1(n9021), .B2(n6565), .A(n6564), .ZN(n6567) );
  NAND2_X1 U8078 ( .A1(n6566), .A2(n6567), .ZN(n6573) );
  INV_X1 U8079 ( .A(n6566), .ZN(n6569) );
  INV_X1 U8080 ( .A(n6567), .ZN(n6568) );
  NAND2_X1 U8081 ( .A1(n6569), .A2(n6568), .ZN(n6570) );
  NAND2_X1 U8082 ( .A1(n6573), .A2(n6570), .ZN(n7048) );
  INV_X1 U8083 ( .A(n7048), .ZN(n6571) );
  NAND2_X1 U8084 ( .A1(n6572), .A2(n6571), .ZN(n7050) );
  XNOR2_X1 U8085 ( .A(n6575), .B(n6574), .ZN(n7195) );
  NAND2_X1 U8086 ( .A1(n7194), .A2(n7195), .ZN(n7204) );
  NAND2_X1 U8087 ( .A1(n6576), .A2(n7204), .ZN(n7207) );
  INV_X1 U8088 ( .A(n6577), .ZN(n6579) );
  NAND2_X1 U8089 ( .A1(n6579), .A2(n6578), .ZN(n6580) );
  NAND2_X1 U8090 ( .A1(n7207), .A2(n6580), .ZN(n6583) );
  OAI22_X1 U8091 ( .A1(n7558), .A2(n6727), .B1(n9378), .B2(n6733), .ZN(n6581)
         );
  XNOR2_X1 U8092 ( .A(n6581), .B(n7546), .ZN(n6582) );
  NAND2_X1 U8093 ( .A1(n6583), .A2(n6582), .ZN(n6584) );
  OR2_X1 U8094 ( .A1(n7558), .A2(n6755), .ZN(n6586) );
  NAND2_X1 U8095 ( .A1(n10176), .A2(n6608), .ZN(n6585) );
  AND2_X1 U8096 ( .A1(n6586), .A2(n6585), .ZN(n7404) );
  OAI22_X1 U8097 ( .A1(n7544), .A2(n6727), .B1(n10184), .B2(n6733), .ZN(n6587)
         );
  XNOR2_X1 U8098 ( .A(n6587), .B(n7546), .ZN(n6592) );
  OAI22_X1 U8099 ( .A1(n7544), .A2(n6755), .B1(n10184), .B2(n6727), .ZN(n6591)
         );
  OR2_X1 U8100 ( .A1(n6592), .A2(n6591), .ZN(n7552) );
  INV_X1 U8101 ( .A(n7552), .ZN(n6589) );
  NOR2_X1 U8102 ( .A1(n6589), .A2(n6588), .ZN(n6590) );
  NAND2_X1 U8103 ( .A1(n7403), .A2(n6590), .ZN(n6593) );
  NAND2_X1 U8104 ( .A1(n6592), .A2(n6591), .ZN(n7551) );
  OR2_X1 U8105 ( .A1(n7557), .A2(n6755), .ZN(n6595) );
  NAND2_X1 U8106 ( .A1(n7622), .A2(n6608), .ZN(n6594) );
  NAND2_X1 U8107 ( .A1(n6595), .A2(n6594), .ZN(n7566) );
  OAI22_X1 U8108 ( .A1(n7557), .A2(n6727), .B1(n10192), .B2(n6733), .ZN(n6596)
         );
  XNOR2_X1 U8109 ( .A(n6596), .B(n7546), .ZN(n7565) );
  OR2_X1 U8110 ( .A1(n7797), .A2(n6755), .ZN(n6598) );
  NAND2_X1 U8111 ( .A1(n7777), .A2(n6608), .ZN(n6597) );
  NAND2_X1 U8112 ( .A1(n6598), .A2(n6597), .ZN(n7637) );
  OAI22_X1 U8113 ( .A1(n7797), .A2(n6727), .B1(n10199), .B2(n6733), .ZN(n6599)
         );
  XNOR2_X1 U8114 ( .A(n6599), .B(n7546), .ZN(n7636) );
  NAND2_X1 U8115 ( .A1(n7853), .A2(n6759), .ZN(n6601) );
  NAND2_X1 U8116 ( .A1(n9016), .A2(n6608), .ZN(n6600) );
  NAND2_X1 U8117 ( .A1(n6601), .A2(n6600), .ZN(n6602) );
  XNOR2_X1 U8118 ( .A(n6602), .B(n6712), .ZN(n6604) );
  AOI22_X1 U8119 ( .A1(n7853), .A2(n6608), .B1(n6565), .B2(n9016), .ZN(n6603)
         );
  NAND2_X1 U8120 ( .A1(n6604), .A2(n6603), .ZN(n6607) );
  OR2_X1 U8121 ( .A1(n6604), .A2(n6603), .ZN(n6605) );
  NAND2_X1 U8122 ( .A1(n6607), .A2(n6605), .ZN(n7795) );
  INV_X1 U8123 ( .A(n7795), .ZN(n6606) );
  NAND2_X1 U8124 ( .A1(n7881), .A2(n6759), .ZN(n6610) );
  OR2_X1 U8125 ( .A1(n7890), .A2(n6727), .ZN(n6609) );
  NAND2_X1 U8126 ( .A1(n6610), .A2(n6609), .ZN(n6611) );
  XNOR2_X1 U8127 ( .A(n6611), .B(n6712), .ZN(n6613) );
  INV_X1 U8128 ( .A(n7890), .ZN(n9015) );
  AOI22_X1 U8129 ( .A1(n7881), .A2(n6608), .B1(n6565), .B2(n9015), .ZN(n6612)
         );
  OR2_X1 U8130 ( .A1(n6613), .A2(n6612), .ZN(n7828) );
  NAND2_X1 U8131 ( .A1(n6613), .A2(n6612), .ZN(n7827) );
  NAND2_X1 U8132 ( .A1(n7986), .A2(n6759), .ZN(n6615) );
  NAND2_X1 U8133 ( .A1(n9014), .A2(n6608), .ZN(n6614) );
  NAND2_X1 U8134 ( .A1(n6615), .A2(n6614), .ZN(n6616) );
  XNOR2_X1 U8135 ( .A(n6616), .B(n6712), .ZN(n6619) );
  AND2_X1 U8136 ( .A1(n9014), .A2(n6565), .ZN(n6617) );
  AOI21_X1 U8137 ( .B1(n7986), .B2(n6608), .A(n6617), .ZN(n6620) );
  XNOR2_X1 U8138 ( .A(n6619), .B(n6620), .ZN(n7936) );
  INV_X1 U8139 ( .A(n6619), .ZN(n6622) );
  INV_X1 U8140 ( .A(n6620), .ZN(n6621) );
  NAND2_X1 U8141 ( .A1(n6622), .A2(n6621), .ZN(n6623) );
  NAND2_X1 U8142 ( .A1(n8075), .A2(n6759), .ZN(n6625) );
  OR2_X1 U8143 ( .A1(n8082), .A2(n6727), .ZN(n6624) );
  NAND2_X1 U8144 ( .A1(n6625), .A2(n6624), .ZN(n6626) );
  XNOR2_X1 U8145 ( .A(n6626), .B(n6712), .ZN(n6629) );
  NOR2_X1 U8146 ( .A1(n8082), .A2(n6755), .ZN(n6627) );
  AOI21_X1 U8147 ( .B1(n8075), .B2(n6608), .A(n6627), .ZN(n6628) );
  XNOR2_X1 U8148 ( .A(n6629), .B(n6628), .ZN(n8069) );
  NAND2_X1 U8149 ( .A1(n6629), .A2(n6628), .ZN(n6630) );
  NAND2_X1 U8150 ( .A1(n9932), .A2(n6759), .ZN(n6632) );
  NAND2_X1 U8151 ( .A1(n9070), .A2(n6608), .ZN(n6631) );
  NAND2_X1 U8152 ( .A1(n6632), .A2(n6631), .ZN(n6633) );
  XNOR2_X1 U8153 ( .A(n6633), .B(n6712), .ZN(n8080) );
  AND2_X1 U8154 ( .A1(n9070), .A2(n6565), .ZN(n6634) );
  AOI21_X1 U8155 ( .B1(n9932), .B2(n6608), .A(n6634), .ZN(n8079) );
  AND2_X1 U8156 ( .A1(n8080), .A2(n8079), .ZN(n6635) );
  NAND2_X1 U8157 ( .A1(n9463), .A2(n6759), .ZN(n6637) );
  NAND2_X1 U8158 ( .A1(n9073), .A2(n6608), .ZN(n6636) );
  NAND2_X1 U8159 ( .A1(n6637), .A2(n6636), .ZN(n6638) );
  XNOR2_X1 U8160 ( .A(n6638), .B(n7546), .ZN(n8123) );
  INV_X1 U8161 ( .A(n8123), .ZN(n6641) );
  NAND2_X1 U8162 ( .A1(n9463), .A2(n6608), .ZN(n6640) );
  NAND2_X1 U8163 ( .A1(n9073), .A2(n6565), .ZN(n6639) );
  NAND2_X1 U8164 ( .A1(n6640), .A2(n6639), .ZN(n6645) );
  INV_X1 U8165 ( .A(n6645), .ZN(n8122) );
  NAND2_X1 U8166 ( .A1(n6641), .A2(n8122), .ZN(n6658) );
  NAND2_X1 U8167 ( .A1(n9925), .A2(n6759), .ZN(n6643) );
  OR2_X1 U8168 ( .A1(n8932), .A2(n6727), .ZN(n6642) );
  NAND2_X1 U8169 ( .A1(n6643), .A2(n6642), .ZN(n6644) );
  XNOR2_X1 U8170 ( .A(n6644), .B(n7546), .ZN(n6659) );
  INV_X1 U8171 ( .A(n6659), .ZN(n6646) );
  AND2_X1 U8172 ( .A1(n6646), .A2(n4550), .ZN(n6647) );
  NAND2_X1 U8173 ( .A1(n6648), .A2(n6647), .ZN(n8997) );
  NAND2_X1 U8174 ( .A1(n9925), .A2(n6608), .ZN(n6650) );
  OR2_X1 U8175 ( .A1(n8932), .A2(n6755), .ZN(n6649) );
  NAND2_X1 U8176 ( .A1(n6650), .A2(n6649), .ZN(n9000) );
  NAND2_X1 U8177 ( .A1(n8997), .A2(n9000), .ZN(n8928) );
  NAND2_X1 U8178 ( .A1(n9323), .A2(n6759), .ZN(n6652) );
  OR2_X1 U8179 ( .A1(n9012), .A2(n6727), .ZN(n6651) );
  NAND2_X1 U8180 ( .A1(n6652), .A2(n6651), .ZN(n6653) );
  XNOR2_X1 U8181 ( .A(n6653), .B(n6712), .ZN(n6656) );
  NOR2_X1 U8182 ( .A1(n9012), .A2(n6755), .ZN(n6654) );
  AOI21_X1 U8183 ( .B1(n9323), .B2(n6608), .A(n6654), .ZN(n6655) );
  NAND2_X1 U8184 ( .A1(n6656), .A2(n6655), .ZN(n6660) );
  OR2_X1 U8185 ( .A1(n6656), .A2(n6655), .ZN(n6657) );
  AND2_X1 U8186 ( .A1(n6660), .A2(n6657), .ZN(n8929) );
  NAND3_X1 U8187 ( .A1(n8928), .A2(n8929), .A3(n8998), .ZN(n8927) );
  NAND2_X1 U8188 ( .A1(n8927), .A2(n6660), .ZN(n8937) );
  NAND2_X1 U8189 ( .A1(n9458), .A2(n6759), .ZN(n6662) );
  NAND2_X1 U8190 ( .A1(n9314), .A2(n6608), .ZN(n6661) );
  NAND2_X1 U8191 ( .A1(n6662), .A2(n6661), .ZN(n6663) );
  XNOR2_X1 U8192 ( .A(n6663), .B(n7546), .ZN(n6665) );
  AND2_X1 U8193 ( .A1(n9314), .A2(n6565), .ZN(n6664) );
  AOI21_X1 U8194 ( .B1(n9458), .B2(n6608), .A(n6664), .ZN(n6666) );
  XNOR2_X1 U8195 ( .A(n6665), .B(n6666), .ZN(n8939) );
  INV_X1 U8196 ( .A(n6665), .ZN(n6667) );
  NAND2_X1 U8197 ( .A1(n6667), .A2(n6666), .ZN(n6668) );
  NAND2_X1 U8198 ( .A1(n9452), .A2(n6759), .ZN(n6670) );
  OR2_X1 U8199 ( .A1(n9011), .A2(n6727), .ZN(n6669) );
  NAND2_X1 U8200 ( .A1(n6670), .A2(n6669), .ZN(n6671) );
  XNOR2_X1 U8201 ( .A(n6671), .B(n6712), .ZN(n6674) );
  INV_X1 U8202 ( .A(n6674), .ZN(n6672) );
  NOR2_X1 U8203 ( .A1(n9011), .A2(n6755), .ZN(n6673) );
  AOI21_X1 U8204 ( .B1(n9452), .B2(n6608), .A(n6673), .ZN(n8979) );
  NAND2_X1 U8205 ( .A1(n6675), .A2(n6674), .ZN(n8978) );
  NAND2_X1 U8206 ( .A1(n9447), .A2(n6759), .ZN(n6678) );
  NAND2_X1 U8207 ( .A1(n9290), .A2(n6608), .ZN(n6677) );
  NAND2_X1 U8208 ( .A1(n6678), .A2(n6677), .ZN(n6679) );
  XNOR2_X1 U8209 ( .A(n6679), .B(n7546), .ZN(n6682) );
  NAND2_X1 U8210 ( .A1(n9447), .A2(n6608), .ZN(n6681) );
  NAND2_X1 U8211 ( .A1(n9290), .A2(n6565), .ZN(n6680) );
  NAND2_X1 U8212 ( .A1(n6681), .A2(n6680), .ZN(n6683) );
  NAND2_X1 U8213 ( .A1(n6682), .A2(n6683), .ZN(n8903) );
  INV_X1 U8214 ( .A(n6682), .ZN(n6685) );
  INV_X1 U8215 ( .A(n6683), .ZN(n6684) );
  NAND2_X1 U8216 ( .A1(n6685), .A2(n6684), .ZN(n8902) );
  NAND2_X1 U8217 ( .A1(n9442), .A2(n6759), .ZN(n6687) );
  NAND2_X1 U8218 ( .A1(n9276), .A2(n6608), .ZN(n6686) );
  NAND2_X1 U8219 ( .A1(n6687), .A2(n6686), .ZN(n6688) );
  XNOR2_X1 U8220 ( .A(n6688), .B(n7546), .ZN(n6690) );
  AND2_X1 U8221 ( .A1(n9276), .A2(n6565), .ZN(n6689) );
  AOI21_X1 U8222 ( .B1(n9442), .B2(n6608), .A(n6689), .ZN(n6691) );
  XNOR2_X1 U8223 ( .A(n6690), .B(n6691), .ZN(n8955) );
  INV_X1 U8224 ( .A(n6690), .ZN(n6692) );
  NAND2_X1 U8225 ( .A1(n6692), .A2(n6691), .ZN(n6693) );
  NAND2_X1 U8226 ( .A1(n9439), .A2(n6759), .ZN(n6695) );
  INV_X1 U8227 ( .A(n9235), .ZN(n9264) );
  NAND2_X1 U8228 ( .A1(n9264), .A2(n6608), .ZN(n6694) );
  NAND2_X1 U8229 ( .A1(n6695), .A2(n6694), .ZN(n6696) );
  XNOR2_X1 U8230 ( .A(n6696), .B(n7546), .ZN(n6698) );
  NOR2_X1 U8231 ( .A1(n9235), .A2(n6755), .ZN(n6697) );
  AOI21_X1 U8232 ( .B1(n9439), .B2(n6608), .A(n6697), .ZN(n6699) );
  XNOR2_X1 U8233 ( .A(n6698), .B(n6699), .ZN(n8911) );
  INV_X1 U8234 ( .A(n6698), .ZN(n6700) );
  NAND2_X1 U8235 ( .A1(n9432), .A2(n6608), .ZN(n6702) );
  NAND2_X1 U8236 ( .A1(n9083), .A2(n6565), .ZN(n6701) );
  NAND2_X1 U8237 ( .A1(n6702), .A2(n6701), .ZN(n6707) );
  NAND2_X1 U8238 ( .A1(n6706), .A2(n6707), .ZN(n8967) );
  NAND2_X1 U8239 ( .A1(n9432), .A2(n6759), .ZN(n6704) );
  NAND2_X1 U8240 ( .A1(n9083), .A2(n6608), .ZN(n6703) );
  NAND2_X1 U8241 ( .A1(n6704), .A2(n6703), .ZN(n6705) );
  XNOR2_X1 U8242 ( .A(n6705), .B(n6712), .ZN(n8966) );
  NAND2_X1 U8243 ( .A1(n8967), .A2(n8966), .ZN(n8965) );
  INV_X1 U8244 ( .A(n6706), .ZN(n6709) );
  INV_X1 U8245 ( .A(n6707), .ZN(n6708) );
  NAND2_X1 U8246 ( .A1(n9426), .A2(n6759), .ZN(n6711) );
  NAND2_X1 U8247 ( .A1(n9198), .A2(n6608), .ZN(n6710) );
  NAND2_X1 U8248 ( .A1(n6711), .A2(n6710), .ZN(n6713) );
  AND2_X1 U8249 ( .A1(n9198), .A2(n6565), .ZN(n6714) );
  OAI22_X1 U8250 ( .A1(n9090), .A2(n6733), .B1(n9089), .B2(n6727), .ZN(n6717)
         );
  XNOR2_X1 U8251 ( .A(n6717), .B(n7546), .ZN(n6718) );
  INV_X1 U8252 ( .A(n9089), .ZN(n9091) );
  XNOR2_X1 U8253 ( .A(n6718), .B(n6719), .ZN(n8947) );
  INV_X1 U8254 ( .A(n6718), .ZN(n6720) );
  NAND2_X1 U8255 ( .A1(n9416), .A2(n6759), .ZN(n6722) );
  OR2_X1 U8256 ( .A1(n9092), .A2(n6727), .ZN(n6721) );
  NAND2_X1 U8257 ( .A1(n6722), .A2(n6721), .ZN(n6723) );
  XNOR2_X1 U8258 ( .A(n6725), .B(n6724), .ZN(n8921) );
  OAI22_X1 U8259 ( .A1(n9094), .A2(n6733), .B1(n9093), .B2(n6727), .ZN(n6726)
         );
  XNOR2_X1 U8260 ( .A(n6726), .B(n7546), .ZN(n6731) );
  NAND2_X1 U8261 ( .A1(n9165), .A2(n6565), .ZN(n6728) );
  XNOR2_X1 U8262 ( .A(n6731), .B(n6730), .ZN(n8990) );
  OAI22_X1 U8263 ( .A1(n9162), .A2(n6733), .B1(n9095), .B2(n6727), .ZN(n6734)
         );
  XOR2_X1 U8264 ( .A(n7546), .B(n6734), .Z(n8879) );
  NOR2_X1 U8265 ( .A1(n9095), .A2(n6755), .ZN(n6735) );
  AOI21_X1 U8266 ( .B1(n9405), .B2(n6608), .A(n6735), .ZN(n8878) );
  NAND3_X1 U8267 ( .A1(n7952), .A2(P1_B_REG_SCAN_IN), .A3(n7919), .ZN(n6736)
         );
  OAI211_X1 U8268 ( .C1(P1_B_REG_SCAN_IN), .C2(n7919), .A(n6737), .B(n6736), 
        .ZN(n10152) );
  OR2_X1 U8269 ( .A1(n10152), .A2(P1_D_REG_1__SCAN_IN), .ZN(n6739) );
  INV_X1 U8270 ( .A(n6737), .ZN(n8065) );
  NAND2_X1 U8271 ( .A1(n8065), .A2(n7952), .ZN(n6738) );
  NAND2_X1 U8272 ( .A1(n6739), .A2(n6738), .ZN(n6971) );
  INV_X1 U8273 ( .A(n6971), .ZN(n6813) );
  NOR4_X1 U8274 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n6743) );
  NOR4_X1 U8275 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n6742) );
  NOR4_X1 U8276 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n6741) );
  NOR4_X1 U8277 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n6740) );
  NAND4_X1 U8278 ( .A1(n6743), .A2(n6742), .A3(n6741), .A4(n6740), .ZN(n6749)
         );
  NOR2_X1 U8279 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .ZN(
        n6747) );
  NOR4_X1 U8280 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_2__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n6746) );
  NOR4_X1 U8281 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n6745) );
  NOR4_X1 U8282 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n6744) );
  NAND4_X1 U8283 ( .A1(n6747), .A2(n6746), .A3(n6745), .A4(n6744), .ZN(n6748)
         );
  NOR2_X1 U8284 ( .A1(n6749), .A2(n6748), .ZN(n6750) );
  OR2_X1 U8285 ( .A1(n10152), .A2(n6750), .ZN(n6970) );
  NAND2_X1 U8286 ( .A1(n6813), .A2(n6970), .ZN(n7254) );
  OR2_X1 U8287 ( .A1(n10152), .A2(P1_D_REG_0__SCAN_IN), .ZN(n6752) );
  NAND2_X1 U8288 ( .A1(n8065), .A2(n7919), .ZN(n6751) );
  NAND2_X1 U8289 ( .A1(n6752), .A2(n6751), .ZN(n6979) );
  OR2_X1 U8290 ( .A1(n7254), .A2(n6979), .ZN(n6772) );
  NOR2_X1 U8291 ( .A1(n6772), .A2(n6951), .ZN(n6765) );
  INV_X1 U8292 ( .A(n6790), .ZN(n6753) );
  AND2_X1 U8293 ( .A1(n7660), .A2(n7577), .ZN(n7260) );
  INV_X1 U8294 ( .A(n7260), .ZN(n6977) );
  AND2_X1 U8295 ( .A1(n6753), .A2(n10207), .ZN(n6754) );
  NAND2_X1 U8296 ( .A1(n9400), .A2(n6608), .ZN(n6757) );
  OR2_X1 U8297 ( .A1(n9096), .A2(n6755), .ZN(n6756) );
  NAND2_X1 U8298 ( .A1(n6757), .A2(n6756), .ZN(n6758) );
  XNOR2_X1 U8299 ( .A(n6758), .B(n7546), .ZN(n6761) );
  AOI22_X1 U8300 ( .A1(n9400), .A2(n6759), .B1(n6608), .B2(n9097), .ZN(n6760)
         );
  XNOR2_X1 U8301 ( .A(n6761), .B(n6760), .ZN(n6762) );
  NAND3_X1 U8302 ( .A1(n6764), .A2(n8956), .A3(n6762), .ZN(n6785) );
  INV_X1 U8303 ( .A(n6762), .ZN(n6763) );
  INV_X1 U8304 ( .A(n6765), .ZN(n6767) );
  INV_X1 U8305 ( .A(n7524), .ZN(n7350) );
  NAND2_X1 U8306 ( .A1(n7260), .A2(n7350), .ZN(n7262) );
  OR2_X1 U8307 ( .A1(n6767), .A2(n7262), .ZN(n6766) );
  NAND2_X1 U8308 ( .A1(n10125), .A2(n10138), .ZN(n6969) );
  NAND2_X1 U8309 ( .A1(n6766), .A2(n10151), .ZN(n9007) );
  OR2_X1 U8310 ( .A1(n6767), .A2(n6768), .ZN(n8915) );
  INV_X1 U8311 ( .A(n8151), .ZN(n6857) );
  INV_X1 U8312 ( .A(n9368), .ZN(n9236) );
  OR2_X1 U8313 ( .A1(n8915), .A2(n9236), .ZN(n8960) );
  NOR2_X1 U8314 ( .A1(n9095), .A2(n8960), .ZN(n6777) );
  OR2_X1 U8315 ( .A1(n8915), .A2(n9238), .ZN(n8981) );
  NAND2_X1 U8316 ( .A1(n6772), .A2(n10207), .ZN(n6952) );
  AND2_X1 U8317 ( .A1(n6790), .A2(n6768), .ZN(n6950) );
  INV_X1 U8318 ( .A(n6789), .ZN(n6787) );
  NOR2_X1 U8319 ( .A1(n6950), .A2(n6787), .ZN(n6769) );
  NAND3_X1 U8320 ( .A1(n6952), .A2(n6788), .A3(n6769), .ZN(n6770) );
  NAND2_X1 U8321 ( .A1(n6770), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6773) );
  NOR2_X1 U8322 ( .A1(n6951), .A2(n7262), .ZN(n6771) );
  NAND2_X1 U8323 ( .A1(n6772), .A2(n6771), .ZN(n6953) );
  NAND2_X1 U8324 ( .A1(n6773), .A2(n6953), .ZN(n8962) );
  AOI22_X1 U8325 ( .A1(n9145), .A2(n8962), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n6774) );
  OAI21_X1 U8326 ( .B1(n6775), .B2(n8981), .A(n6774), .ZN(n6776) );
  NOR2_X1 U8327 ( .A1(n6780), .A2(n6779), .ZN(n6784) );
  INV_X1 U8328 ( .A(n6781), .ZN(n6782) );
  OAI211_X1 U8329 ( .C1(n6786), .C2(n6785), .A(n6784), .B(n6783), .ZN(P1_U3218) );
  OR2_X1 U8330 ( .A1(n6788), .A2(n6787), .ZN(n6832) );
  NAND2_X1 U8331 ( .A1(n6790), .A2(n6789), .ZN(n6791) );
  NAND2_X1 U8332 ( .A1(n6832), .A2(n6791), .ZN(n6846) );
  OAI21_X1 U8333 ( .B1(n6846), .B2(n4752), .A(P1_STATE_REG_SCAN_IN), .ZN(
        P1_U3083) );
  NOR2_X2 U8334 ( .A1(n6832), .A2(P1_U3084), .ZN(P1_U4006) );
  INV_X1 U8335 ( .A(n7058), .ZN(n6792) );
  NAND2_X1 U8336 ( .A1(n6792), .A2(n10275), .ZN(n8372) );
  XNOR2_X1 U8337 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  NAND2_X1 U8338 ( .A1(n4483), .A2(P1_U3084), .ZN(n9487) );
  OR2_X1 U8339 ( .A1(n4483), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9489) );
  OAI222_X1 U8340 ( .A1(n6939), .A2(P1_U3084), .B1(n9487), .B2(n6797), .C1(
        n6793), .C2(n9489), .ZN(P1_U3352) );
  OAI222_X1 U8341 ( .A1(n6881), .A2(P1_U3084), .B1(n9487), .B2(n6799), .C1(
        n6794), .C2(n9489), .ZN(P1_U3350) );
  INV_X1 U8342 ( .A(n9487), .ZN(n8103) );
  INV_X1 U8343 ( .A(n8103), .ZN(n9492) );
  OAI222_X1 U8344 ( .A1(n6860), .A2(P1_U3084), .B1(n9492), .B2(n6798), .C1(
        n6795), .C2(n9489), .ZN(P1_U3351) );
  OAI222_X1 U8345 ( .A1(n9489), .A2(n9657), .B1(n9487), .B2(n6800), .C1(
        P1_U3084), .C2(n6796), .ZN(P1_U3346) );
  NAND2_X1 U8346 ( .A1(n4483), .A2(P2_U3152), .ZN(n8876) );
  INV_X1 U8347 ( .A(n8876), .ZN(n7137) );
  INV_X1 U8348 ( .A(n7137), .ZN(n8865) );
  OR2_X1 U8349 ( .A1(n4483), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8871) );
  INV_X1 U8350 ( .A(n8871), .ZN(n8132) );
  INV_X1 U8351 ( .A(n8132), .ZN(n8874) );
  OAI222_X1 U8352 ( .A1(n8865), .A2(n4580), .B1(n8874), .B2(n6797), .C1(
        P2_U3152), .C2(n7107), .ZN(P2_U3357) );
  OAI222_X1 U8353 ( .A1(n8865), .A2(n4584), .B1(n8871), .B2(n6798), .C1(
        P2_U3152), .C2(n7079), .ZN(P2_U3356) );
  OAI222_X1 U8354 ( .A1(n8865), .A2(n4632), .B1(n8874), .B2(n6799), .C1(
        P2_U3152), .C2(n7120), .ZN(P2_U3355) );
  OAI222_X1 U8355 ( .A1(n8865), .A2(n6801), .B1(n8874), .B2(n6800), .C1(
        P2_U3152), .C2(n7167), .ZN(P2_U3351) );
  OAI222_X1 U8356 ( .A1(n8865), .A2(n6802), .B1(n8871), .B2(n6805), .C1(
        P2_U3152), .C2(n7135), .ZN(P2_U3354) );
  OAI222_X1 U8357 ( .A1(n8865), .A2(n6803), .B1(n8874), .B2(n6807), .C1(
        P2_U3152), .C2(n7191), .ZN(P2_U3352) );
  OAI222_X1 U8358 ( .A1(n8865), .A2(n6804), .B1(n8874), .B2(n6809), .C1(
        P2_U3152), .C2(n7179), .ZN(P2_U3353) );
  INV_X1 U8359 ( .A(n9489), .ZN(n9485) );
  INV_X1 U8360 ( .A(n9485), .ZN(n8155) );
  OAI222_X1 U8361 ( .A1(n8155), .A2(n6806), .B1(n9492), .B2(n6805), .C1(
        P1_U3084), .C2(n9979), .ZN(P1_U3349) );
  OAI222_X1 U8362 ( .A1(n8155), .A2(n6808), .B1(n9487), .B2(n6807), .C1(
        P1_U3084), .C2(n6925), .ZN(P1_U3347) );
  OAI222_X1 U8363 ( .A1(n8155), .A2(n6810), .B1(n9487), .B2(n6809), .C1(
        P1_U3084), .C2(n6883), .ZN(P1_U3348) );
  INV_X1 U8364 ( .A(n6956), .ZN(n6964) );
  OAI222_X1 U8365 ( .A1(n8155), .A2(n9833), .B1(n9487), .B2(n6811), .C1(
        P1_U3084), .C2(n6964), .ZN(P1_U3345) );
  OAI222_X1 U8366 ( .A1(n8865), .A2(n6812), .B1(n8874), .B2(n6811), .C1(
        P2_U3152), .C2(n7281), .ZN(P2_U3350) );
  INV_X1 U8367 ( .A(n6951), .ZN(n10153) );
  INV_X1 U8368 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n9602) );
  NAND2_X1 U8369 ( .A1(n6813), .A2(n10153), .ZN(n6814) );
  OAI21_X1 U8370 ( .B1(n10153), .B2(n9602), .A(n6814), .ZN(P1_U3441) );
  INV_X1 U8371 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n9646) );
  INV_X1 U8372 ( .A(n6979), .ZN(n6815) );
  NAND2_X1 U8373 ( .A1(n6815), .A2(n10153), .ZN(n6816) );
  OAI21_X1 U8374 ( .B1(n10153), .B2(n9646), .A(n6816), .ZN(P1_U3440) );
  INV_X1 U8375 ( .A(n6817), .ZN(n6819) );
  INV_X1 U8376 ( .A(n8391), .ZN(n7283) );
  OAI222_X1 U8377 ( .A1(n8876), .A2(n6818), .B1(n8874), .B2(n6819), .C1(n7283), 
        .C2(P2_U3152), .ZN(P2_U3349) );
  INV_X1 U8378 ( .A(n10015), .ZN(n6897) );
  OAI222_X1 U8379 ( .A1(n8155), .A2(n9806), .B1(n9492), .B2(n6819), .C1(n6897), 
        .C2(P1_U3084), .ZN(P1_U3344) );
  INV_X1 U8380 ( .A(n6820), .ZN(n6830) );
  AOI22_X1 U8381 ( .A1(n8407), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n7137), .ZN(n6821) );
  OAI21_X1 U8382 ( .B1(n6830), .B2(n8871), .A(n6821), .ZN(P2_U3347) );
  INV_X1 U8383 ( .A(n6822), .ZN(n6824) );
  INV_X1 U8384 ( .A(n7484), .ZN(n7473) );
  OAI222_X1 U8385 ( .A1(n8876), .A2(n6823), .B1(n8874), .B2(n6824), .C1(n7473), 
        .C2(P2_U3152), .ZN(P2_U3348) );
  INV_X1 U8386 ( .A(n9025), .ZN(n9036) );
  OAI222_X1 U8387 ( .A1(n8155), .A2(n9669), .B1(n9492), .B2(n6824), .C1(n9036), 
        .C2(P1_U3084), .ZN(P1_U3343) );
  OAI21_X1 U8388 ( .B1(n10268), .B2(n5878), .A(n6825), .ZN(n6827) );
  NAND2_X1 U8389 ( .A1(n10268), .A2(n7011), .ZN(n6826) );
  AND2_X1 U8390 ( .A1(n6827), .A2(n6826), .ZN(n8481) );
  NOR2_X1 U8391 ( .A1(n10234), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U8392 ( .A(n8485), .ZN(n6828) );
  NAND2_X1 U8393 ( .A1(n6828), .A2(P2_U3966), .ZN(n6829) );
  OAI21_X1 U8394 ( .B1(n5918), .B2(P2_U3966), .A(n6829), .ZN(P2_U3583) );
  INV_X1 U8395 ( .A(n10026), .ZN(n9037) );
  OAI222_X1 U8396 ( .A1(n8155), .A2(n6831), .B1(n9492), .B2(n6830), .C1(n9037), 
        .C2(P1_U3084), .ZN(P1_U3342) );
  INV_X1 U8397 ( .A(n6832), .ZN(n9962) );
  OR2_X1 U8398 ( .A1(P1_U3083), .A2(n9962), .ZN(n10123) );
  INV_X1 U8399 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n6843) );
  INV_X1 U8400 ( .A(n6481), .ZN(n9059) );
  OR2_X1 U8401 ( .A1(n8151), .A2(n9059), .ZN(n9960) );
  OAI21_X1 U8402 ( .B1(n6833), .B2(n8151), .A(n9960), .ZN(n6834) );
  XNOR2_X1 U8403 ( .A(n6834), .B(P1_IR_REG_0__SCAN_IN), .ZN(n6835) );
  NOR2_X1 U8404 ( .A1(n6835), .A2(P1_U3084), .ZN(n9964) );
  AOI211_X1 U8405 ( .C1(n6481), .C2(n6836), .A(n4752), .B(n6846), .ZN(n6841)
         );
  INV_X1 U8406 ( .A(n6846), .ZN(n6837) );
  NOR2_X1 U8407 ( .A1(n9960), .A2(P1_U3084), .ZN(n9965) );
  NAND3_X1 U8408 ( .A1(n10117), .A2(P1_IR_REG_0__SCAN_IN), .A3(n6836), .ZN(
        n6838) );
  OAI21_X1 U8409 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n6839), .A(n6838), .ZN(n6840) );
  AOI21_X1 U8410 ( .B1(n9964), .B2(n6841), .A(n6840), .ZN(n6842) );
  OAI21_X1 U8411 ( .B1(n10123), .B2(n6843), .A(n6842), .ZN(P1_U3241) );
  INV_X1 U8412 ( .A(n6844), .ZN(n6868) );
  AOI22_X1 U8413 ( .A1(n7672), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_12__SCAN_IN), .B2(n7137), .ZN(n6845) );
  OAI21_X1 U8414 ( .B1(n6868), .B2(n8871), .A(n6845), .ZN(P2_U3346) );
  INV_X1 U8415 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n6867) );
  OR2_X1 U8416 ( .A1(n6481), .A2(P1_U3084), .ZN(n8104) );
  NOR2_X1 U8417 ( .A1(n6846), .A2(n8104), .ZN(n9052) );
  AND2_X1 U8418 ( .A1(n9052), .A2(n8151), .ZN(n10116) );
  INV_X1 U8419 ( .A(n6881), .ZN(n6856) );
  AND2_X1 U8420 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_U3084), .ZN(n7198) );
  INV_X1 U8421 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6847) );
  MUX2_X1 U8422 ( .A(n6847), .B(P1_REG1_REG_2__SCAN_IN), .S(n6860), .Z(n9974)
         );
  INV_X1 U8423 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10218) );
  MUX2_X1 U8424 ( .A(n10218), .B(P1_REG1_REG_1__SCAN_IN), .S(n6939), .Z(n6849)
         );
  AND2_X1 U8425 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n6848) );
  NAND2_X1 U8426 ( .A1(n6849), .A2(n6848), .ZN(n6936) );
  OR2_X1 U8427 ( .A1(n6860), .A2(n6847), .ZN(n6853) );
  NAND2_X1 U8428 ( .A1(n9973), .A2(n6853), .ZN(n6851) );
  MUX2_X1 U8429 ( .A(n6871), .B(P1_REG1_REG_3__SCAN_IN), .S(n6881), .Z(n6850)
         );
  NAND2_X1 U8430 ( .A1(n6851), .A2(n6850), .ZN(n6873) );
  MUX2_X1 U8431 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n6871), .S(n6881), .Z(n6852)
         );
  NAND3_X1 U8432 ( .A1(n9973), .A2(n6853), .A3(n6852), .ZN(n6854) );
  AND3_X1 U8433 ( .A1(n10117), .A2(n6873), .A3(n6854), .ZN(n6855) );
  AOI211_X1 U8434 ( .C1(n10116), .C2(n6856), .A(n7198), .B(n6855), .ZN(n6866)
         );
  AND2_X1 U8435 ( .A1(n9052), .A2(n6857), .ZN(n10030) );
  INV_X1 U8436 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6858) );
  MUX2_X1 U8437 ( .A(n6858), .B(P1_REG2_REG_2__SCAN_IN), .S(n6860), .Z(n9969)
         );
  AND2_X1 U8438 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n6943) );
  NAND2_X1 U8439 ( .A1(n9969), .A2(n9968), .ZN(n9967) );
  INV_X1 U8440 ( .A(n6860), .ZN(n9966) );
  NAND2_X1 U8441 ( .A1(n9966), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6863) );
  MUX2_X1 U8442 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n6880), .S(n6881), .Z(n6862)
         );
  AOI21_X1 U8443 ( .B1(n9967), .B2(n6863), .A(n6862), .ZN(n6861) );
  INV_X1 U8444 ( .A(n6861), .ZN(n6879) );
  NAND3_X1 U8445 ( .A1(n9967), .A2(n6863), .A3(n6862), .ZN(n6864) );
  NAND3_X1 U8446 ( .A1(n10030), .A2(n6879), .A3(n6864), .ZN(n6865) );
  OAI211_X1 U8447 ( .C1(n6867), .C2(n10123), .A(n6866), .B(n6865), .ZN(
        P1_U3244) );
  INV_X1 U8448 ( .A(n10038), .ZN(n9038) );
  OAI222_X1 U8449 ( .A1(n8155), .A2(n6869), .B1(n9487), .B2(n6868), .C1(
        P1_U3084), .C2(n9038), .ZN(P1_U3341) );
  INV_X1 U8450 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n6890) );
  INV_X1 U8451 ( .A(n6883), .ZN(n6902) );
  NOR2_X1 U8452 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6870), .ZN(n7407) );
  INV_X1 U8453 ( .A(n9979), .ZN(n9984) );
  OR2_X1 U8454 ( .A1(n6881), .A2(n6871), .ZN(n6872) );
  NAND2_X1 U8455 ( .A1(n6873), .A2(n6872), .ZN(n9978) );
  INV_X1 U8456 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6874) );
  MUX2_X1 U8457 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n6874), .S(n9979), .Z(n6875)
         );
  OAI21_X1 U8458 ( .B1(P1_REG1_REG_4__SCAN_IN), .B2(n9984), .A(n9980), .ZN(
        n6877) );
  INV_X1 U8459 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n10222) );
  MUX2_X1 U8460 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n10222), .S(n6883), .Z(n6876)
         );
  INV_X1 U8461 ( .A(n10117), .ZN(n10071) );
  AOI211_X1 U8462 ( .C1(n6877), .C2(n6876), .A(n6895), .B(n10071), .ZN(n6878)
         );
  AOI211_X1 U8463 ( .C1(n10116), .C2(n6902), .A(n7407), .B(n6878), .ZN(n6889)
         );
  OAI21_X1 U8464 ( .B1(n6881), .B2(n6880), .A(n6879), .ZN(n9990) );
  MUX2_X1 U8465 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n6882), .S(n9979), .Z(n9991)
         );
  NOR2_X1 U8466 ( .A1(n9990), .A2(n9991), .ZN(n9989) );
  NOR2_X1 U8467 ( .A1(n9984), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6884) );
  MUX2_X1 U8468 ( .A(n9373), .B(P1_REG2_REG_5__SCAN_IN), .S(n6883), .Z(n6885)
         );
  OAI21_X1 U8469 ( .B1(n9989), .B2(n6884), .A(n6885), .ZN(n6901) );
  INV_X1 U8470 ( .A(n6901), .ZN(n6887) );
  NOR3_X1 U8471 ( .A1(n9989), .A2(n6885), .A3(n6884), .ZN(n6886) );
  OAI21_X1 U8472 ( .B1(n6887), .B2(n6886), .A(n10030), .ZN(n6888) );
  OAI211_X1 U8473 ( .C1(n6890), .C2(n10123), .A(n6889), .B(n6888), .ZN(
        P1_U3246) );
  INV_X1 U8474 ( .A(n6891), .ZN(n6893) );
  INV_X1 U8475 ( .A(n9039), .ZN(n10053) );
  OAI222_X1 U8476 ( .A1(n9489), .A2(n6892), .B1(n9487), .B2(n6893), .C1(n10053), .C2(P1_U3084), .ZN(P1_U3340) );
  INV_X1 U8477 ( .A(n7726), .ZN(n7721) );
  OAI222_X1 U8478 ( .A1(n8876), .A2(n6894), .B1(n8874), .B2(n6893), .C1(n7721), 
        .C2(P2_U3152), .ZN(P2_U3345) );
  NOR2_X1 U8479 ( .A1(n10015), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6898) );
  AOI21_X1 U8480 ( .B1(n6902), .B2(P1_REG1_REG_5__SCAN_IN), .A(n6895), .ZN(
        n6920) );
  MUX2_X1 U8481 ( .A(n6079), .B(P1_REG1_REG_6__SCAN_IN), .S(n6925), .Z(n6919)
         );
  AND2_X1 U8482 ( .A1(n6920), .A2(n6919), .ZN(n6922) );
  MUX2_X1 U8483 ( .A(n6896), .B(P1_REG1_REG_7__SCAN_IN), .S(n9997), .Z(n10003)
         );
  NOR2_X1 U8484 ( .A1(n10004), .A2(n10003), .ZN(n10002) );
  NOR2_X1 U8485 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(n9997), .ZN(n6960) );
  INV_X1 U8486 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10226) );
  MUX2_X1 U8487 ( .A(n10226), .B(P1_REG1_REG_8__SCAN_IN), .S(n6956), .Z(n6959)
         );
  INV_X1 U8488 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10229) );
  AOI22_X1 U8489 ( .A1(n10015), .A2(n10229), .B1(P1_REG1_REG_9__SCAN_IN), .B2(
        n6897), .ZN(n10017) );
  NOR2_X1 U8490 ( .A1(n10016), .A2(n10017), .ZN(n10018) );
  AOI22_X1 U8491 ( .A1(n9025), .A2(n6132), .B1(P1_REG1_REG_10__SCAN_IN), .B2(
        n9036), .ZN(n6899) );
  NOR2_X1 U8492 ( .A1(n6900), .A2(n6899), .ZN(n9035) );
  AOI21_X1 U8493 ( .B1(n6900), .B2(n6899), .A(n9035), .ZN(n6915) );
  OAI21_X1 U8494 ( .B1(P1_REG2_REG_5__SCAN_IN), .B2(n6902), .A(n6901), .ZN(
        n6929) );
  MUX2_X1 U8495 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n6083), .S(n6925), .Z(n6928)
         );
  OAI21_X1 U8496 ( .B1(n6083), .B2(n6925), .A(n6926), .ZN(n9999) );
  MUX2_X1 U8497 ( .A(n6903), .B(P1_REG2_REG_7__SCAN_IN), .S(n9997), .Z(n10000)
         );
  NOR2_X1 U8498 ( .A1(n9999), .A2(n10000), .ZN(n9998) );
  NOR2_X1 U8499 ( .A1(P1_REG2_REG_7__SCAN_IN), .A2(n9997), .ZN(n6904) );
  NOR2_X1 U8500 ( .A1(n9998), .A2(n6904), .ZN(n6958) );
  NOR2_X1 U8501 ( .A1(n6964), .A2(n7629), .ZN(n6905) );
  OAI22_X1 U8502 ( .A1(n6958), .A2(n6905), .B1(n6956), .B2(
        P1_REG2_REG_8__SCAN_IN), .ZN(n10011) );
  NAND2_X1 U8503 ( .A1(n10015), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6906) );
  OAI21_X1 U8504 ( .B1(n10015), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6906), .ZN(
        n10012) );
  NOR2_X1 U8505 ( .A1(n10011), .A2(n10012), .ZN(n10010) );
  NAND2_X1 U8506 ( .A1(n9025), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6907) );
  OAI21_X1 U8507 ( .B1(n9025), .B2(P1_REG2_REG_10__SCAN_IN), .A(n6907), .ZN(
        n6908) );
  INV_X1 U8508 ( .A(n10030), .ZN(n10109) );
  AOI211_X1 U8509 ( .C1(n6909), .C2(n6908), .A(n9024), .B(n10109), .ZN(n6910)
         );
  INV_X1 U8510 ( .A(n6910), .ZN(n6914) );
  INV_X1 U8511 ( .A(n10123), .ZN(n10068) );
  AND2_X1 U8512 ( .A1(P1_U3084), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n6912) );
  INV_X1 U8513 ( .A(n10116), .ZN(n10054) );
  NOR2_X1 U8514 ( .A1(n10054), .A2(n9036), .ZN(n6911) );
  AOI211_X1 U8515 ( .C1(P1_ADDR_REG_10__SCAN_IN), .C2(n10068), .A(n6912), .B(
        n6911), .ZN(n6913) );
  OAI211_X1 U8516 ( .C1(n6915), .C2(n10071), .A(n6914), .B(n6913), .ZN(
        P1_U3251) );
  INV_X1 U8517 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n9824) );
  INV_X1 U8518 ( .A(n6916), .ZN(n6917) );
  INV_X1 U8519 ( .A(n10064), .ZN(n9040) );
  OAI222_X1 U8520 ( .A1(n9489), .A2(n9824), .B1(n9487), .B2(n6917), .C1(n9040), 
        .C2(P1_U3084), .ZN(P1_U3339) );
  INV_X1 U8521 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6918) );
  INV_X1 U8522 ( .A(n7972), .ZN(n7976) );
  OAI222_X1 U8523 ( .A1(n8876), .A2(n6918), .B1(n8874), .B2(n6917), .C1(n7976), 
        .C2(P2_U3152), .ZN(P2_U3344) );
  NAND2_X1 U8524 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3084), .ZN(n6924) );
  NOR2_X1 U8525 ( .A1(n6920), .A2(n6919), .ZN(n6921) );
  OAI21_X1 U8526 ( .B1(n6922), .B2(n6921), .A(n10117), .ZN(n6923) );
  OAI211_X1 U8527 ( .C1(n10054), .C2(n6925), .A(n6924), .B(n6923), .ZN(n6931)
         );
  INV_X1 U8528 ( .A(n6926), .ZN(n6927) );
  AOI211_X1 U8529 ( .C1(n6929), .C2(n6928), .A(n6927), .B(n10109), .ZN(n6930)
         );
  AOI211_X1 U8530 ( .C1(P1_ADDR_REG_6__SCAN_IN), .C2(n10068), .A(n6931), .B(
        n6930), .ZN(n6932) );
  INV_X1 U8531 ( .A(n6932), .ZN(P1_U3247) );
  INV_X1 U8532 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n6946) );
  NAND2_X1 U8533 ( .A1(P1_REG3_REG_1__SCAN_IN), .A2(P1_U3084), .ZN(n6938) );
  INV_X1 U8534 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n6934) );
  MUX2_X1 U8535 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n10218), .S(n6939), .Z(n6933)
         );
  OAI21_X1 U8536 ( .B1(n6836), .B2(n6934), .A(n6933), .ZN(n6935) );
  NAND3_X1 U8537 ( .A1(n10117), .A2(n6936), .A3(n6935), .ZN(n6937) );
  OAI211_X1 U8538 ( .C1(n10054), .C2(n6939), .A(n6938), .B(n6937), .ZN(n6940)
         );
  INV_X1 U8539 ( .A(n6940), .ZN(n6945) );
  OAI211_X1 U8540 ( .C1(n6943), .C2(n6942), .A(n10030), .B(n6941), .ZN(n6944)
         );
  OAI211_X1 U8541 ( .C1(n6946), .C2(n10123), .A(n6945), .B(n6944), .ZN(
        P1_U3242) );
  OAI21_X1 U8542 ( .B1(n6949), .B2(n6948), .A(n6947), .ZN(n9961) );
  NAND2_X1 U8543 ( .A1(n9961), .A2(n8956), .ZN(n6955) );
  OR2_X1 U8544 ( .A1(n6951), .A2(n6950), .ZN(n6972) );
  INV_X1 U8545 ( .A(n6972), .ZN(n6980) );
  NAND3_X1 U8546 ( .A1(n6953), .A2(n6952), .A3(n6980), .ZN(n8147) );
  AOI22_X1 U8547 ( .A1(n9007), .A2(n7238), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        n8147), .ZN(n6954) );
  OAI211_X1 U8548 ( .C1(n7052), .C2(n8981), .A(n6955), .B(n6954), .ZN(P1_U3230) );
  MUX2_X1 U8549 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n7629), .S(n6956), .Z(n6957)
         );
  XNOR2_X1 U8550 ( .A(n6958), .B(n6957), .ZN(n6968) );
  OAI21_X1 U8551 ( .B1(n10002), .B2(n6960), .A(n6959), .ZN(n6962) );
  NAND3_X1 U8552 ( .A1(n6962), .A2(n10117), .A3(n6961), .ZN(n6967) );
  NAND2_X1 U8553 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3084), .ZN(n6963) );
  OAI21_X1 U8554 ( .B1(n10054), .B2(n6964), .A(n6963), .ZN(n6965) );
  AOI21_X1 U8555 ( .B1(n10068), .B2(P1_ADDR_REG_8__SCAN_IN), .A(n6965), .ZN(
        n6966) );
  OAI211_X1 U8556 ( .C1(n6968), .C2(n10109), .A(n6967), .B(n6966), .ZN(
        P1_U3249) );
  AND3_X1 U8557 ( .A1(n6971), .A2(n6970), .A3(n6969), .ZN(n6981) );
  NOR2_X1 U8558 ( .A1(n6972), .A2(n6979), .ZN(n6973) );
  AND2_X2 U8559 ( .A1(n6981), .A2(n6973), .ZN(n10231) );
  INV_X1 U8560 ( .A(n7547), .ZN(n6974) );
  NOR2_X1 U8561 ( .A1(n6974), .A2(n7260), .ZN(n6975) );
  AOI22_X1 U8562 ( .A1(n6976), .A2(n6975), .B1(n9370), .B2(n6552), .ZN(n10147)
         );
  OAI21_X1 U8563 ( .B1(n10144), .B2(n6977), .A(n10147), .ZN(n6982) );
  NAND2_X1 U8564 ( .A1(n6982), .A2(n10231), .ZN(n6978) );
  OAI21_X1 U8565 ( .B1(n10231), .B2(n6836), .A(n6978), .ZN(P1_U3523) );
  AND2_X1 U8566 ( .A1(n6980), .A2(n6979), .ZN(n7255) );
  AND2_X2 U8567 ( .A1(n7255), .A2(n6981), .ZN(n10217) );
  INV_X1 U8568 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6984) );
  NAND2_X1 U8569 ( .A1(n6982), .A2(n10217), .ZN(n6983) );
  OAI21_X1 U8570 ( .B1(n10217), .B2(n6984), .A(n6983), .ZN(P1_U3454) );
  CLKBUF_X1 U8571 ( .A(P1_U4006), .Z(n9022) );
  NAND2_X1 U8572 ( .A1(n9061), .A2(n9022), .ZN(n6985) );
  OAI21_X1 U8573 ( .B1(n9022), .B2(n8866), .A(n6985), .ZN(P1_U3586) );
  NAND2_X1 U8574 ( .A1(n8505), .A2(P2_U3966), .ZN(n6986) );
  OAI21_X1 U8575 ( .B1(n7714), .B2(P2_U3966), .A(n6986), .ZN(P2_U3575) );
  NAND2_X1 U8576 ( .A1(n8385), .A2(n7363), .ZN(n7328) );
  INV_X1 U8577 ( .A(n7328), .ZN(n7214) );
  NAND2_X1 U8578 ( .A1(n7214), .A2(n8168), .ZN(n7042) );
  NAND3_X1 U8579 ( .A1(n7225), .A2(n10277), .A3(n7578), .ZN(n6988) );
  NAND2_X1 U8580 ( .A1(n6987), .A2(n7491), .ZN(n7221) );
  OR2_X1 U8581 ( .A1(n7363), .A2(n7953), .ZN(n6989) );
  AND2_X1 U8582 ( .A1(n7042), .A2(n6989), .ZN(n6991) );
  XNOR2_X1 U8583 ( .A(n4581), .B(n7953), .ZN(n7025) );
  XNOR2_X1 U8584 ( .A(n7027), .B(n7025), .ZN(n6990) );
  OAI21_X1 U8585 ( .B1(n6991), .B2(n6990), .A(n7029), .ZN(n7010) );
  XOR2_X1 U8586 ( .A(n7872), .B(P2_B_REG_SCAN_IN), .Z(n6992) );
  OR2_X1 U8587 ( .A1(n7946), .A2(n6992), .ZN(n6993) );
  INV_X1 U8588 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n10271) );
  AND2_X1 U8589 ( .A1(n10267), .A2(n10271), .ZN(n6994) );
  INV_X1 U8590 ( .A(n6995), .ZN(n8061) );
  AND2_X1 U8591 ( .A1(n8061), .A2(n7872), .ZN(n10270) );
  NOR2_X1 U8592 ( .A1(n6994), .A2(n10270), .ZN(n7437) );
  INV_X1 U8593 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n10273) );
  NOR2_X1 U8594 ( .A1(n7946), .A2(n6995), .ZN(n10274) );
  AOI21_X1 U8595 ( .B1(n10267), .B2(n10273), .A(n10274), .ZN(n7427) );
  NOR4_X1 U8596 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n6999) );
  NOR4_X1 U8597 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n6998) );
  NOR4_X1 U8598 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n6997) );
  NOR4_X1 U8599 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n6996) );
  NAND4_X1 U8600 ( .A1(n6999), .A2(n6998), .A3(n6997), .A4(n6996), .ZN(n7005)
         );
  NOR2_X1 U8601 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .ZN(
        n7003) );
  NOR4_X1 U8602 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n7002) );
  NOR4_X1 U8603 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n7001) );
  NOR4_X1 U8604 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n7000) );
  NAND4_X1 U8605 ( .A1(n7003), .A2(n7002), .A3(n7001), .A4(n7000), .ZN(n7004)
         );
  OAI21_X1 U8606 ( .B1(n7005), .B2(n7004), .A(n10267), .ZN(n7426) );
  NAND2_X1 U8607 ( .A1(n7427), .A2(n7426), .ZN(n7215) );
  INV_X1 U8608 ( .A(n7215), .ZN(n7006) );
  NAND2_X1 U8609 ( .A1(n7437), .A2(n7006), .ZN(n7016) );
  INV_X1 U8610 ( .A(n10268), .ZN(n7007) );
  OR2_X1 U8611 ( .A1(n7016), .A2(n7007), .ZN(n7015) );
  INV_X1 U8612 ( .A(n7015), .ZN(n7009) );
  OR2_X1 U8613 ( .A1(n10277), .A2(n7018), .ZN(n10335) );
  AND2_X1 U8614 ( .A1(n10335), .A2(n7057), .ZN(n7008) );
  NAND2_X1 U8615 ( .A1(n7009), .A2(n7008), .ZN(n8340) );
  INV_X1 U8616 ( .A(n8340), .ZN(n8353) );
  NAND2_X1 U8617 ( .A1(n7010), .A2(n8353), .ZN(n7024) );
  AND2_X1 U8618 ( .A1(n7089), .A2(n7011), .ZN(n8702) );
  OAI22_X1 U8619 ( .A1(n7012), .A2(n8637), .B1(n8223), .B2(n8639), .ZN(n7226)
         );
  OR2_X1 U8620 ( .A1(n7217), .A2(n7016), .ZN(n8291) );
  INV_X1 U8621 ( .A(n8291), .ZN(n8362) );
  NOR2_X1 U8622 ( .A1(n10277), .A2(n7491), .ZN(n10258) );
  INV_X1 U8623 ( .A(n10258), .ZN(n7014) );
  OR2_X1 U8624 ( .A1(n10336), .A2(n8478), .ZN(n7425) );
  INV_X1 U8625 ( .A(n7425), .ZN(n7013) );
  NAND2_X1 U8626 ( .A1(n10268), .A2(n7013), .ZN(n8620) );
  OAI21_X2 U8627 ( .B1(n7015), .B2(n7014), .A(n8620), .ZN(n8324) );
  NAND2_X1 U8628 ( .A1(n7016), .A2(n7425), .ZN(n7021) );
  OAI211_X1 U8629 ( .C1(n7018), .C2(n7057), .A(n7058), .B(n7017), .ZN(n7019)
         );
  INV_X1 U8630 ( .A(n7019), .ZN(n7020) );
  NAND2_X1 U8631 ( .A1(n7021), .A2(n7020), .ZN(n7151) );
  NOR2_X1 U8632 ( .A1(n7151), .A2(P2_U3152), .ZN(n7043) );
  INV_X1 U8633 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n9847) );
  AOI21_X1 U8634 ( .B1(n7226), .B2(n8362), .A(n7022), .ZN(n7023) );
  NAND2_X1 U8635 ( .A1(n7024), .A2(n7023), .ZN(P2_U3224) );
  INV_X1 U8636 ( .A(n7025), .ZN(n7026) );
  NAND2_X1 U8637 ( .A1(n7027), .A2(n7026), .ZN(n7028) );
  XNOR2_X1 U8638 ( .A(n7338), .B(n7953), .ZN(n7031) );
  NAND2_X1 U8639 ( .A1(n7030), .A2(n7031), .ZN(n7140) );
  INV_X1 U8640 ( .A(n7030), .ZN(n7032) );
  INV_X1 U8641 ( .A(n7031), .ZN(n8222) );
  OAI211_X1 U8642 ( .C1(n7033), .C2(n4509), .A(n8221), .B(n8353), .ZN(n7038)
         );
  INV_X1 U8643 ( .A(n8637), .ZN(n8700) );
  NAND2_X1 U8644 ( .A1(n8362), .A2(n8700), .ZN(n8347) );
  OAI22_X1 U8645 ( .A1(n7361), .A2(n8347), .B1(n8366), .B2(n7034), .ZN(n7036)
         );
  NOR2_X1 U8646 ( .A1(n8291), .A2(n8639), .ZN(n8349) );
  INV_X1 U8647 ( .A(n8349), .ZN(n8321) );
  OAI22_X1 U8648 ( .A1(n7372), .A2(n8321), .B1(n7043), .B2(n7336), .ZN(n7035)
         );
  NOR2_X1 U8649 ( .A1(n7036), .A2(n7035), .ZN(n7037) );
  NAND2_X1 U8650 ( .A1(n7038), .A2(n7037), .ZN(P2_U3239) );
  INV_X1 U8651 ( .A(n7039), .ZN(n7040) );
  INV_X1 U8652 ( .A(n10077), .ZN(n9029) );
  OAI222_X1 U8653 ( .A1(n9489), .A2(n9584), .B1(n9487), .B2(n7040), .C1(
        P1_U3084), .C2(n9029), .ZN(P1_U3338) );
  INV_X1 U8654 ( .A(n8416), .ZN(n8424) );
  OAI222_X1 U8655 ( .A1(n8865), .A2(n7041), .B1(n8874), .B2(n7040), .C1(
        P2_U3152), .C2(n8424), .ZN(P2_U3343) );
  INV_X1 U8656 ( .A(n7042), .ZN(n7047) );
  OR2_X1 U8657 ( .A1(n8340), .A2(n8243), .ZN(n8301) );
  INV_X1 U8658 ( .A(n8301), .ZN(n8352) );
  AOI22_X1 U8659 ( .A1(n8352), .A2(n8385), .B1(n7363), .B2(n8353), .ZN(n7046)
         );
  INV_X1 U8660 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n9599) );
  OAI22_X1 U8661 ( .A1(n7361), .A2(n8321), .B1(n7043), .B2(n9599), .ZN(n7044)
         );
  AOI21_X1 U8662 ( .B1(n7363), .B2(n8324), .A(n7044), .ZN(n7045) );
  OAI21_X1 U8663 ( .B1(n7047), .B2(n7046), .A(n7045), .ZN(P2_U3234) );
  INV_X1 U8664 ( .A(n7050), .ZN(n7051) );
  AOI21_X1 U8665 ( .B1(n7048), .B2(n7049), .A(n7051), .ZN(n7056) );
  INV_X1 U8666 ( .A(n9007), .ZN(n8996) );
  NOR2_X1 U8667 ( .A1(n8996), .A2(n6046), .ZN(n7054) );
  OAI22_X1 U8668 ( .A1(n6544), .A2(n8981), .B1(n8960), .B2(n7052), .ZN(n7053)
         );
  AOI211_X1 U8669 ( .C1(P1_REG3_REG_2__SCAN_IN), .C2(n8147), .A(n7054), .B(
        n7053), .ZN(n7055) );
  OAI21_X1 U8670 ( .B1(n7056), .B2(n9009), .A(n7055), .ZN(P1_U3235) );
  OR2_X1 U8671 ( .A1(n7089), .A2(P2_U3152), .ZN(n8133) );
  NAND2_X1 U8672 ( .A1(n10268), .A2(n7057), .ZN(n7216) );
  OAI211_X1 U8673 ( .C1(n8133), .C2(n7058), .A(n7216), .B(n7716), .ZN(n7074)
         );
  NAND2_X1 U8674 ( .A1(n7074), .A2(n5142), .ZN(n7059) );
  NAND2_X1 U8675 ( .A1(n7059), .A2(n8384), .ZN(n7091) );
  AND2_X1 U8676 ( .A1(n7091), .A2(n7089), .ZN(n9897) );
  NOR2_X1 U8677 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7518), .ZN(n7078) );
  NAND2_X1 U8678 ( .A1(n7088), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7072) );
  INV_X1 U8679 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n7060) );
  MUX2_X1 U8680 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n7060), .S(n7088), .Z(n7163)
         );
  INV_X1 U8681 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n7441) );
  MUX2_X1 U8682 ( .A(n7441), .B(P2_REG1_REG_6__SCAN_IN), .S(n7191), .Z(n7187)
         );
  NAND2_X1 U8683 ( .A1(n7083), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n7071) );
  INV_X1 U8684 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n7061) );
  MUX2_X1 U8685 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n7061), .S(n7083), .Z(n7175)
         );
  INV_X1 U8686 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n7122) );
  INV_X1 U8687 ( .A(n7107), .ZN(n7080) );
  INV_X1 U8688 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10346) );
  MUX2_X1 U8689 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n10346), .S(n7107), .Z(n7098)
         );
  INV_X1 U8690 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n7063) );
  INV_X1 U8691 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n7062) );
  NOR3_X1 U8692 ( .A1(n7098), .A2(n7063), .A3(n7062), .ZN(n7097) );
  AOI21_X1 U8693 ( .B1(n7080), .B2(P2_REG1_REG_1__SCAN_IN), .A(n7097), .ZN(
        n9900) );
  INV_X1 U8694 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10348) );
  MUX2_X1 U8695 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n10348), .S(n7079), .Z(n9899)
         );
  NOR2_X1 U8696 ( .A1(n9900), .A2(n9899), .ZN(n9898) );
  INV_X1 U8697 ( .A(n9898), .ZN(n7066) );
  NOR2_X1 U8698 ( .A1(n7079), .A2(n10348), .ZN(n7109) );
  INV_X1 U8699 ( .A(n7109), .ZN(n7065) );
  INV_X1 U8700 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10350) );
  MUX2_X1 U8701 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n10350), .S(n7120), .Z(n7064)
         );
  AOI21_X1 U8702 ( .B1(n7066), .B2(n7065), .A(n7064), .ZN(n7125) );
  INV_X1 U8703 ( .A(n7125), .ZN(n7069) );
  INV_X1 U8704 ( .A(n7120), .ZN(n7067) );
  NAND2_X1 U8705 ( .A1(n7067), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n7121) );
  MUX2_X1 U8706 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n7122), .S(n7135), .Z(n7068)
         );
  AOI21_X1 U8707 ( .B1(n7069), .B2(n7121), .A(n7068), .ZN(n7127) );
  INV_X1 U8708 ( .A(n7127), .ZN(n7070) );
  OAI21_X1 U8709 ( .B1(n7122), .B2(n7135), .A(n7070), .ZN(n7176) );
  NAND2_X1 U8710 ( .A1(n7175), .A2(n7176), .ZN(n7174) );
  NAND2_X1 U8711 ( .A1(n7071), .A2(n7174), .ZN(n7188) );
  NAND2_X1 U8712 ( .A1(n7187), .A2(n7188), .ZN(n7186) );
  OAI21_X1 U8713 ( .B1(n7191), .B2(n7441), .A(n7186), .ZN(n7164) );
  NAND2_X1 U8714 ( .A1(n7163), .A2(n7164), .ZN(n7162) );
  AND2_X1 U8715 ( .A1(n7072), .A2(n7162), .ZN(n7076) );
  INV_X1 U8716 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10354) );
  MUX2_X1 U8717 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n10354), .S(n7281), .Z(n7075)
         );
  AND2_X1 U8718 ( .A1(n5142), .A2(n8484), .ZN(n7073) );
  NAND2_X1 U8719 ( .A1(n7074), .A2(n7073), .ZN(n10236) );
  NOR2_X1 U8720 ( .A1(n7076), .A2(n7075), .ZN(n8398) );
  AOI211_X1 U8721 ( .C1(n7076), .C2(n7075), .A(n10236), .B(n8398), .ZN(n7077)
         );
  AOI211_X1 U8722 ( .C1(P2_ADDR_REG_8__SCAN_IN), .C2(n10234), .A(n7078), .B(
        n7077), .ZN(n7096) );
  INV_X1 U8723 ( .A(n7191), .ZN(n7086) );
  INV_X1 U8724 ( .A(n7135), .ZN(n7081) );
  INV_X1 U8725 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n7418) );
  INV_X1 U8726 ( .A(n7079), .ZN(n9896) );
  MUX2_X1 U8727 ( .A(n7334), .B(P2_REG2_REG_2__SCAN_IN), .S(n7079), .Z(n9892)
         );
  AND2_X1 U8728 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(
        n7103) );
  NAND2_X1 U8729 ( .A1(n7104), .A2(n7103), .ZN(n7102) );
  AOI21_X1 U8730 ( .B1(P2_REG2_REG_2__SCAN_IN), .B2(n9896), .A(n9893), .ZN(
        n7114) );
  XNOR2_X1 U8731 ( .A(n7120), .B(n7418), .ZN(n7113) );
  OAI21_X1 U8732 ( .B1(n7418), .B2(n7120), .A(n7115), .ZN(n7131) );
  XNOR2_X1 U8733 ( .A(n7135), .B(P2_REG2_REG_4__SCAN_IN), .ZN(n7132) );
  NAND2_X1 U8734 ( .A1(n7131), .A2(n7132), .ZN(n7130) );
  NAND2_X1 U8735 ( .A1(n7083), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n7082) );
  OAI21_X1 U8736 ( .B1(n7083), .B2(P2_REG2_REG_5__SCAN_IN), .A(n7082), .ZN(
        n7171) );
  INV_X1 U8737 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7084) );
  MUX2_X1 U8738 ( .A(n7084), .B(P2_REG2_REG_6__SCAN_IN), .S(n7191), .Z(n7085)
         );
  INV_X1 U8739 ( .A(n7085), .ZN(n7183) );
  NOR2_X1 U8740 ( .A1(n7184), .A2(n7183), .ZN(n7182) );
  NAND2_X1 U8741 ( .A1(n7088), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n7087) );
  OAI21_X1 U8742 ( .B1(n7088), .B2(P2_REG2_REG_7__SCAN_IN), .A(n7087), .ZN(
        n7159) );
  XOR2_X1 U8743 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n7281), .Z(n7092) );
  NOR2_X1 U8744 ( .A1(n7089), .A2(n8484), .ZN(n7090) );
  NAND2_X1 U8745 ( .A1(n7091), .A2(n7090), .ZN(n10237) );
  AOI211_X1 U8746 ( .C1(n7093), .C2(n7092), .A(n7272), .B(n10237), .ZN(n7094)
         );
  INV_X1 U8747 ( .A(n7094), .ZN(n7095) );
  OAI211_X1 U8748 ( .C1(n10235), .C2(n7281), .A(n7096), .B(n7095), .ZN(
        P2_U3253) );
  NAND2_X1 U8749 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n7099) );
  AOI211_X1 U8750 ( .C1(n7099), .C2(n7098), .A(n7097), .B(n10236), .ZN(n7101)
         );
  INV_X1 U8751 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n9499) );
  OAI22_X1 U8752 ( .A1(n8481), .A2(n9499), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9847), .ZN(n7100) );
  NOR2_X1 U8753 ( .A1(n7101), .A2(n7100), .ZN(n7106) );
  INV_X1 U8754 ( .A(n10237), .ZN(n10233) );
  OAI211_X1 U8755 ( .C1(n7104), .C2(n7103), .A(n10233), .B(n7102), .ZN(n7105)
         );
  OAI211_X1 U8756 ( .C1(n10235), .C2(n7107), .A(n7106), .B(n7105), .ZN(
        P2_U3246) );
  NOR2_X1 U8757 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9820), .ZN(n7112) );
  MUX2_X1 U8758 ( .A(n10350), .B(P2_REG1_REG_3__SCAN_IN), .S(n7120), .Z(n7108)
         );
  NOR3_X1 U8759 ( .A1(n9898), .A2(n7109), .A3(n7108), .ZN(n7110) );
  NOR3_X1 U8760 ( .A1(n10236), .A2(n7125), .A3(n7110), .ZN(n7111) );
  AOI211_X1 U8761 ( .C1(P2_ADDR_REG_3__SCAN_IN), .C2(n10234), .A(n7112), .B(
        n7111), .ZN(n7119) );
  INV_X1 U8762 ( .A(n7113), .ZN(n7117) );
  INV_X1 U8763 ( .A(n7114), .ZN(n7116) );
  OAI211_X1 U8764 ( .C1(n7117), .C2(n7116), .A(n10233), .B(n7115), .ZN(n7118)
         );
  OAI211_X1 U8765 ( .C1(n10235), .C2(n7120), .A(n7119), .B(n7118), .ZN(
        P2_U3248) );
  INV_X1 U8766 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n9621) );
  NOR2_X1 U8767 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9621), .ZN(n7129) );
  INV_X1 U8768 ( .A(n7121), .ZN(n7124) );
  MUX2_X1 U8769 ( .A(n7122), .B(P2_REG1_REG_4__SCAN_IN), .S(n7135), .Z(n7123)
         );
  NOR3_X1 U8770 ( .A1(n7125), .A2(n7124), .A3(n7123), .ZN(n7126) );
  NOR3_X1 U8771 ( .A1(n10236), .A2(n7127), .A3(n7126), .ZN(n7128) );
  AOI211_X1 U8772 ( .C1(P2_ADDR_REG_4__SCAN_IN), .C2(n10234), .A(n7129), .B(
        n7128), .ZN(n7134) );
  OAI211_X1 U8773 ( .C1(n7132), .C2(n7131), .A(n10233), .B(n7130), .ZN(n7133)
         );
  OAI211_X1 U8774 ( .C1(n10235), .C2(n7135), .A(n7134), .B(n7133), .ZN(
        P2_U3249) );
  INV_X1 U8775 ( .A(n7136), .ZN(n7139) );
  AOI22_X1 U8776 ( .A1(n8437), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n7137), .ZN(n7138) );
  OAI21_X1 U8777 ( .B1(n7139), .B2(n8871), .A(n7138), .ZN(P2_U3342) );
  INV_X1 U8778 ( .A(n10089), .ZN(n9043) );
  OAI222_X1 U8779 ( .A1(n9489), .A2(n9849), .B1(n9487), .B2(n7139), .C1(n9043), 
        .C2(P1_U3084), .ZN(P1_U3337) );
  OR2_X1 U8780 ( .A1(n7414), .A2(n8243), .ZN(n7291) );
  XNOR2_X1 U8781 ( .A(n10244), .B(n7953), .ZN(n7289) );
  XNOR2_X1 U8782 ( .A(n7291), .B(n7289), .ZN(n7150) );
  AND2_X1 U8783 ( .A1(n8382), .A2(n8168), .ZN(n7141) );
  XNOR2_X1 U8784 ( .A(n10302), .B(n8156), .ZN(n7142) );
  NAND2_X1 U8785 ( .A1(n7141), .A2(n7142), .ZN(n7146) );
  INV_X1 U8786 ( .A(n7141), .ZN(n7143) );
  INV_X1 U8787 ( .A(n7142), .ZN(n7149) );
  NAND2_X1 U8788 ( .A1(n7143), .A2(n7149), .ZN(n7144) );
  AND2_X1 U8789 ( .A1(n7146), .A2(n7144), .ZN(n8219) );
  NAND2_X1 U8790 ( .A1(n7145), .A2(n8219), .ZN(n7148) );
  AND2_X1 U8791 ( .A1(n7150), .A2(n7146), .ZN(n7147) );
  OAI21_X1 U8792 ( .B1(n7150), .B2(n7148), .A(n7293), .ZN(n7156) );
  NOR4_X1 U8793 ( .A1(n7150), .A2(n7372), .A3(n7149), .A4(n8301), .ZN(n7155)
         );
  OAI22_X1 U8794 ( .A1(n7372), .A2(n8637), .B1(n7301), .B2(n8639), .ZN(n7446)
         );
  NAND2_X1 U8795 ( .A1(n7446), .A2(n8362), .ZN(n7153) );
  AOI22_X1 U8796 ( .A1(n8344), .A2(n7443), .B1(P2_REG3_REG_4__SCAN_IN), .B2(
        P2_U3152), .ZN(n7152) );
  OAI211_X1 U8797 ( .C1(n10308), .C2(n8366), .A(n7153), .B(n7152), .ZN(n7154)
         );
  AOI211_X1 U8798 ( .C1(n7156), .C2(n8353), .A(n7155), .B(n7154), .ZN(n7157)
         );
  INV_X1 U8799 ( .A(n7157), .ZN(P2_U3232) );
  AOI211_X1 U8800 ( .C1(n7160), .C2(n7159), .A(n7158), .B(n10237), .ZN(n7169)
         );
  AND2_X1 U8801 ( .A1(P2_U3152), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7161) );
  AOI21_X1 U8802 ( .B1(n10234), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n7161), .ZN(
        n7166) );
  INV_X1 U8803 ( .A(n10236), .ZN(n10232) );
  OAI211_X1 U8804 ( .C1(n7164), .C2(n7163), .A(n10232), .B(n7162), .ZN(n7165)
         );
  OAI211_X1 U8805 ( .C1(n10235), .C2(n7167), .A(n7166), .B(n7165), .ZN(n7168)
         );
  OR2_X1 U8806 ( .A1(n7169), .A2(n7168), .ZN(P2_U3252) );
  AOI211_X1 U8807 ( .C1(n7172), .C2(n7171), .A(n7170), .B(n10237), .ZN(n7181)
         );
  NOR2_X1 U8808 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5187), .ZN(n7173) );
  AOI21_X1 U8809 ( .B1(n10234), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n7173), .ZN(
        n7178) );
  OAI211_X1 U8810 ( .C1(n7176), .C2(n7175), .A(n10232), .B(n7174), .ZN(n7177)
         );
  OAI211_X1 U8811 ( .C1(n10235), .C2(n7179), .A(n7178), .B(n7177), .ZN(n7180)
         );
  OR2_X1 U8812 ( .A1(n7181), .A2(n7180), .ZN(P2_U3250) );
  AOI211_X1 U8813 ( .C1(n7184), .C2(n7183), .A(n7182), .B(n10237), .ZN(n7193)
         );
  NOR2_X1 U8814 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9610), .ZN(n7185) );
  AOI21_X1 U8815 ( .B1(n10234), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n7185), .ZN(
        n7190) );
  OAI211_X1 U8816 ( .C1(n7188), .C2(n7187), .A(n10232), .B(n7186), .ZN(n7189)
         );
  OAI211_X1 U8817 ( .C1(n10235), .C2(n7191), .A(n7190), .B(n7189), .ZN(n7192)
         );
  OR2_X1 U8818 ( .A1(n7193), .A2(n7192), .ZN(P2_U3251) );
  OAI21_X1 U8819 ( .B1(n7195), .B2(n7194), .A(n7204), .ZN(n7196) );
  NAND2_X1 U8820 ( .A1(n7196), .A2(n8956), .ZN(n7200) );
  OAI22_X1 U8821 ( .A1(n7539), .A2(n8981), .B1(n8960), .B2(n7314), .ZN(n7197)
         );
  AOI211_X1 U8822 ( .C1(n7322), .C2(n9007), .A(n7198), .B(n7197), .ZN(n7199)
         );
  OAI211_X1 U8823 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n9005), .A(n7200), .B(
        n7199), .ZN(P1_U3216) );
  INV_X1 U8824 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n9790) );
  INV_X1 U8825 ( .A(n7201), .ZN(n7202) );
  INV_X1 U8826 ( .A(n10101), .ZN(n9045) );
  OAI222_X1 U8827 ( .A1(n9489), .A2(n9790), .B1(n9487), .B2(n7202), .C1(n9045), 
        .C2(P1_U3084), .ZN(P1_U3336) );
  INV_X1 U8828 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7203) );
  INV_X1 U8829 ( .A(n8448), .ZN(n8455) );
  OAI222_X1 U8830 ( .A1(n8865), .A2(n7203), .B1(n8874), .B2(n7202), .C1(n8455), 
        .C2(P2_U3152), .ZN(P2_U3341) );
  AND2_X1 U8831 ( .A1(n7205), .A2(n7204), .ZN(n7208) );
  OAI211_X1 U8832 ( .C1(n7208), .C2(n7206), .A(n8956), .B(n7207), .ZN(n7212)
         );
  NAND2_X1 U8833 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9995) );
  INV_X1 U8834 ( .A(n9995), .ZN(n7210) );
  OAI22_X1 U8835 ( .A1(n6544), .A2(n8960), .B1(n8981), .B2(n7558), .ZN(n7209)
         );
  AOI211_X1 U8836 ( .C1(n7352), .C2(n9007), .A(n7210), .B(n7209), .ZN(n7211)
         );
  OAI211_X1 U8837 ( .C1(n9005), .C2(n7263), .A(n7212), .B(n7211), .ZN(P1_U3228) );
  NAND2_X1 U8838 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(n8384), .ZN(n7213) );
  OAI21_X1 U8839 ( .B1(n8548), .B2(n8384), .A(n7213), .ZN(P2_U3580) );
  XNOR2_X1 U8840 ( .A(n7329), .B(n7214), .ZN(n10287) );
  NOR2_X1 U8841 ( .A1(n7437), .A2(n7215), .ZN(n7218) );
  NAND2_X1 U8842 ( .A1(n7217), .A2(n7216), .ZN(n7424) );
  NAND2_X1 U8843 ( .A1(n7218), .A2(n7424), .ZN(n7229) );
  XNOR2_X1 U8844 ( .A(n7219), .B(n7221), .ZN(n7220) );
  NAND2_X1 U8845 ( .A1(n7220), .A2(n8478), .ZN(n10298) );
  INV_X1 U8846 ( .A(n7221), .ZN(n7222) );
  NAND2_X1 U8847 ( .A1(n7222), .A2(n4781), .ZN(n7604) );
  NAND2_X1 U8848 ( .A1(n10298), .A2(n7604), .ZN(n10262) );
  NAND2_X1 U8849 ( .A1(n10263), .A2(n10262), .ZN(n8742) );
  INV_X1 U8850 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n7228) );
  XNOR2_X1 U8851 ( .A(n7223), .B(n7329), .ZN(n7227) );
  AND2_X1 U8852 ( .A1(n7225), .A2(n7224), .ZN(n8715) );
  INV_X1 U8853 ( .A(n8715), .ZN(n10254) );
  AOI21_X1 U8854 ( .B1(n7227), .B2(n10254), .A(n7226), .ZN(n10286) );
  MUX2_X1 U8855 ( .A(n7228), .B(n10286), .S(n10263), .Z(n7233) );
  OR2_X1 U8856 ( .A1(n7229), .A2(n4781), .ZN(n8561) );
  XNOR2_X1 U8857 ( .A(n4581), .B(n7363), .ZN(n7230) );
  NOR2_X1 U8858 ( .A1(n7230), .A2(n10336), .ZN(n10282) );
  NAND2_X1 U8859 ( .A1(n10263), .A2(n10258), .ZN(n8733) );
  AOI21_X1 U8860 ( .B1(n8719), .B2(n10282), .A(n7231), .ZN(n7232) );
  OAI211_X1 U8861 ( .C1(n10287), .C2(n8742), .A(n7233), .B(n7232), .ZN(
        P2_U3295) );
  INV_X1 U8862 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n7235) );
  INV_X1 U8863 ( .A(n7234), .ZN(n7236) );
  INV_X1 U8864 ( .A(n10115), .ZN(n9047) );
  OAI222_X1 U8865 ( .A1(n9489), .A2(n7235), .B1(n9492), .B2(n7236), .C1(
        P1_U3084), .C2(n9047), .ZN(P1_U3335) );
  INV_X1 U8866 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7237) );
  OAI222_X1 U8867 ( .A1(n8865), .A2(n7237), .B1(n8871), .B2(n7236), .C1(
        P2_U3152), .C2(n8472), .ZN(P2_U3340) );
  NAND3_X1 U8868 ( .A1(n7547), .A2(n7546), .A3(n9203), .ZN(n10130) );
  INV_X1 U8869 ( .A(n10130), .ZN(n8040) );
  NAND2_X1 U8870 ( .A1(n6552), .A2(n6553), .ZN(n7240) );
  NAND2_X1 U8871 ( .A1(n7314), .A2(n6046), .ZN(n7241) );
  NAND2_X1 U8872 ( .A1(n7310), .A2(n7242), .ZN(n7244) );
  NAND2_X1 U8873 ( .A1(n6544), .A2(n6542), .ZN(n7243) );
  NAND2_X1 U8874 ( .A1(n7244), .A2(n7243), .ZN(n7538) );
  XNOR2_X1 U8875 ( .A(n7538), .B(n7537), .ZN(n7349) );
  OAI22_X1 U8876 ( .A1(n6544), .A2(n9236), .B1(n7558), .B2(n9238), .ZN(n7253)
         );
  NAND3_X1 U8877 ( .A1(n7311), .A2(n7537), .A3(n7245), .ZN(n7250) );
  NAND2_X1 U8878 ( .A1(n7246), .A2(n10138), .ZN(n7249) );
  NAND2_X1 U8879 ( .A1(n7247), .A2(n7350), .ZN(n7248) );
  AND2_X1 U8880 ( .A1(n7249), .A2(n7248), .ZN(n9356) );
  AOI21_X1 U8881 ( .B1(n7251), .B2(n7250), .A(n9356), .ZN(n7252) );
  AOI211_X1 U8882 ( .C1(n8040), .C2(n7349), .A(n7253), .B(n7252), .ZN(n7355)
         );
  INV_X1 U8883 ( .A(n7254), .ZN(n7256) );
  NAND2_X1 U8884 ( .A1(n7256), .A2(n7255), .ZN(n7534) );
  INV_X1 U8885 ( .A(n10143), .ZN(n9353) );
  NAND2_X1 U8886 ( .A1(n10160), .A2(n10144), .ZN(n10124) );
  INV_X1 U8887 ( .A(n7318), .ZN(n7258) );
  INV_X1 U8888 ( .A(n9376), .ZN(n7257) );
  AOI21_X1 U8889 ( .B1(n7352), .B2(n7258), .A(n7257), .ZN(n7353) );
  AND2_X1 U8890 ( .A1(n7260), .A2(n7259), .ZN(n7261) );
  AND2_X1 U8891 ( .A1(n10143), .A2(n7261), .ZN(n9294) );
  INV_X1 U8892 ( .A(n7262), .ZN(n10136) );
  NAND2_X1 U8893 ( .A1(n10143), .A2(n10136), .ZN(n10145) );
  NOR2_X1 U8894 ( .A1(n10145), .A2(n6538), .ZN(n7265) );
  OAI22_X1 U8895 ( .A1(n10143), .A2(n6882), .B1(n7263), .B2(n10151), .ZN(n7264) );
  AOI211_X1 U8896 ( .C1(n7353), .C2(n9294), .A(n7265), .B(n7264), .ZN(n7269)
         );
  NOR2_X1 U8897 ( .A1(n7266), .A2(n9203), .ZN(n7267) );
  NAND2_X1 U8898 ( .A1(n10143), .A2(n7267), .ZN(n9346) );
  INV_X1 U8899 ( .A(n9346), .ZN(n10140) );
  NAND2_X1 U8900 ( .A1(n7349), .A2(n10140), .ZN(n7268) );
  OAI211_X1 U8901 ( .C1(n7355), .C2(n9353), .A(n7269), .B(n7268), .ZN(P1_U3287) );
  NOR2_X1 U8902 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7652), .ZN(n7270) );
  AOI21_X1 U8903 ( .B1(n10234), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n7270), .ZN(
        n7271) );
  INV_X1 U8904 ( .A(n7271), .ZN(n7280) );
  INV_X1 U8905 ( .A(n7281), .ZN(n7273) );
  AOI21_X1 U8906 ( .B1(n7273), .B2(P2_REG2_REG_8__SCAN_IN), .A(n7272), .ZN(
        n8388) );
  OR2_X1 U8907 ( .A1(n8391), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n7275) );
  NAND2_X1 U8908 ( .A1(n8391), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n7274) );
  NAND2_X1 U8909 ( .A1(n7275), .A2(n7274), .ZN(n8387) );
  NOR2_X1 U8910 ( .A1(n8388), .A2(n8387), .ZN(n8386) );
  NAND2_X1 U8911 ( .A1(n7484), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n7276) );
  OAI21_X1 U8912 ( .B1(n7484), .B2(P2_REG2_REG_10__SCAN_IN), .A(n7276), .ZN(
        n7277) );
  AOI211_X1 U8913 ( .C1(n7278), .C2(n7277), .A(n7483), .B(n10237), .ZN(n7279)
         );
  AOI211_X1 U8914 ( .C1(n9897), .C2(n7484), .A(n7280), .B(n7279), .ZN(n7288)
         );
  INV_X1 U8915 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n8392) );
  NOR2_X1 U8916 ( .A1(n7281), .A2(n10354), .ZN(n8393) );
  MUX2_X1 U8917 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n8392), .S(n8391), .Z(n7282)
         );
  OAI21_X1 U8918 ( .B1(n8398), .B2(n8393), .A(n7282), .ZN(n8396) );
  OAI21_X1 U8919 ( .B1(n8392), .B2(n7283), .A(n8396), .ZN(n7286) );
  INV_X1 U8920 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n7284) );
  MUX2_X1 U8921 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n7284), .S(n7484), .Z(n7285)
         );
  NAND2_X1 U8922 ( .A1(n7285), .A2(n7286), .ZN(n7472) );
  OAI211_X1 U8923 ( .C1(n7286), .C2(n7285), .A(n10232), .B(n7472), .ZN(n7287)
         );
  NAND2_X1 U8924 ( .A1(n7288), .A2(n7287), .ZN(P2_U3255) );
  OR2_X1 U8925 ( .A1(n7458), .A2(n8243), .ZN(n7495) );
  XNOR2_X1 U8926 ( .A(n7453), .B(n7953), .ZN(n7493) );
  XNOR2_X1 U8927 ( .A(n7495), .B(n7493), .ZN(n7302) );
  INV_X1 U8928 ( .A(n7289), .ZN(n7290) );
  NAND2_X1 U8929 ( .A1(n7291), .A2(n7290), .ZN(n7292) );
  AND2_X1 U8930 ( .A1(n8380), .A2(n8168), .ZN(n7294) );
  XNOR2_X1 U8931 ( .A(n10259), .B(n7953), .ZN(n7295) );
  NAND2_X1 U8932 ( .A1(n7294), .A2(n7295), .ZN(n7298) );
  INV_X1 U8933 ( .A(n7294), .ZN(n7296) );
  INV_X1 U8934 ( .A(n7295), .ZN(n7300) );
  NAND2_X1 U8935 ( .A1(n7296), .A2(n7300), .ZN(n7297) );
  NAND2_X1 U8936 ( .A1(n7298), .A2(n7297), .ZN(n7344) );
  AND2_X1 U8937 ( .A1(n7302), .A2(n7298), .ZN(n7299) );
  OAI21_X1 U8938 ( .B1(n7302), .B2(n7342), .A(n7497), .ZN(n7308) );
  NOR4_X1 U8939 ( .A1(n7302), .A2(n7301), .A3(n7300), .A4(n8301), .ZN(n7307)
         );
  AOI22_X1 U8940 ( .A1(n8700), .A2(n8380), .B1(n8378), .B2(n8702), .ZN(n7377)
         );
  INV_X1 U8941 ( .A(n8344), .ZN(n8360) );
  INV_X1 U8942 ( .A(n7303), .ZN(n7381) );
  OAI22_X1 U8943 ( .A1(n8360), .A2(n7381), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9610), .ZN(n7304) );
  AOI21_X1 U8944 ( .B1(n7453), .B2(n8324), .A(n7304), .ZN(n7305) );
  OAI21_X1 U8945 ( .B1(n7377), .B2(n8291), .A(n7305), .ZN(n7306) );
  AOI211_X1 U8946 ( .C1(n7308), .C2(n8353), .A(n7307), .B(n7306), .ZN(n7309)
         );
  INV_X1 U8947 ( .A(n7309), .ZN(P2_U3241) );
  XNOR2_X1 U8948 ( .A(n7310), .B(n7313), .ZN(n10169) );
  OAI21_X1 U8949 ( .B1(n7313), .B2(n7312), .A(n7311), .ZN(n7316) );
  INV_X1 U8950 ( .A(n9356), .ZN(n10133) );
  OAI22_X1 U8951 ( .A1(n7314), .A2(n9236), .B1(n7539), .B2(n9238), .ZN(n7315)
         );
  AOI21_X1 U8952 ( .B1(n7316), .B2(n10133), .A(n7315), .ZN(n7317) );
  OAI21_X1 U8953 ( .B1(n10169), .B2(n10130), .A(n7317), .ZN(n10171) );
  NAND2_X1 U8954 ( .A1(n10171), .A2(n10143), .ZN(n7324) );
  OAI22_X1 U8955 ( .A1(n10143), .A2(n6880), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n10151), .ZN(n7321) );
  AND2_X1 U8956 ( .A1(n7390), .A2(n7322), .ZN(n7319) );
  OR2_X1 U8957 ( .A1(n7319), .A2(n7318), .ZN(n10170) );
  INV_X1 U8958 ( .A(n9294), .ZN(n10146) );
  NOR2_X1 U8959 ( .A1(n10170), .A2(n10146), .ZN(n7320) );
  AOI211_X1 U8960 ( .C1(n9343), .C2(n7322), .A(n7321), .B(n7320), .ZN(n7323)
         );
  OAI211_X1 U8961 ( .C1(n10169), .C2(n9346), .A(n7324), .B(n7323), .ZN(
        P1_U3288) );
  INV_X1 U8962 ( .A(n7325), .ZN(n7326) );
  OAI222_X1 U8963 ( .A1(n9489), .A2(n9796), .B1(n9492), .B2(n7326), .C1(n9203), 
        .C2(P1_U3084), .ZN(P1_U3334) );
  OAI222_X1 U8964 ( .A1(n8865), .A2(n7327), .B1(n8871), .B2(n7326), .C1(
        P2_U3152), .C2(n8478), .ZN(P2_U3339) );
  XOR2_X1 U8965 ( .A(n7368), .B(n7367), .Z(n10291) );
  INV_X1 U8966 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n7334) );
  XNOR2_X1 U8967 ( .A(n7332), .B(n7367), .ZN(n7333) );
  AOI222_X1 U8968 ( .A1(n10254), .A2(n7333), .B1(n8382), .B2(n8702), .C1(n5020), .C2(n8700), .ZN(n10293) );
  MUX2_X1 U8969 ( .A(n7334), .B(n10293), .S(n10263), .Z(n7340) );
  INV_X1 U8970 ( .A(n10336), .ZN(n10246) );
  NAND2_X1 U8971 ( .A1(n8719), .A2(n10246), .ZN(n8550) );
  OAI21_X1 U8972 ( .B1(n4581), .B2(n7363), .A(n7338), .ZN(n7335) );
  NAND2_X1 U8973 ( .A1(n7416), .A2(n7335), .ZN(n10292) );
  INV_X1 U8974 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n7336) );
  OAI22_X1 U8975 ( .A1(n8550), .A2(n10292), .B1(n7336), .B2(n8620), .ZN(n7337)
         );
  AOI21_X1 U8976 ( .B1(n8486), .B2(n7338), .A(n7337), .ZN(n7339) );
  OAI211_X1 U8977 ( .C1(n10291), .C2(n8742), .A(n7340), .B(n7339), .ZN(
        P2_U3294) );
  OAI22_X1 U8978 ( .A1(n7414), .A2(n8637), .B1(n7458), .B2(n8639), .ZN(n10253)
         );
  AOI22_X1 U8979 ( .A1(n8344), .A2(n10256), .B1(P2_REG3_REG_5__SCAN_IN), .B2(
        P2_U3152), .ZN(n7341) );
  OAI21_X1 U8980 ( .B1(n8366), .B2(n10317), .A(n7341), .ZN(n7347) );
  INV_X1 U8981 ( .A(n7342), .ZN(n7343) );
  AOI211_X1 U8982 ( .C1(n7345), .C2(n7344), .A(n8340), .B(n7343), .ZN(n7346)
         );
  AOI211_X1 U8983 ( .C1(n8362), .C2(n10253), .A(n7347), .B(n7346), .ZN(n7348)
         );
  INV_X1 U8984 ( .A(n7348), .ZN(P2_U3229) );
  INV_X1 U8985 ( .A(n7349), .ZN(n7356) );
  OR2_X1 U8986 ( .A1(n7351), .A2(n7350), .ZN(n9931) );
  INV_X1 U8987 ( .A(n10207), .ZN(n10177) );
  AOI22_X1 U8988 ( .A1(n7353), .A2(n10125), .B1(n10177), .B2(n7352), .ZN(n7354) );
  OAI211_X1 U8989 ( .C1(n7356), .C2(n9931), .A(n7355), .B(n7354), .ZN(n7358)
         );
  NAND2_X1 U8990 ( .A1(n7358), .A2(n10231), .ZN(n7357) );
  OAI21_X1 U8991 ( .B1(n10231), .B2(n6874), .A(n7357), .ZN(P1_U3527) );
  INV_X1 U8992 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n7360) );
  NAND2_X1 U8993 ( .A1(n7358), .A2(n10217), .ZN(n7359) );
  OAI21_X1 U8994 ( .B1(n10217), .B2(n7360), .A(n7359), .ZN(P1_U3466) );
  INV_X1 U8995 ( .A(n8620), .ZN(n10257) );
  INV_X1 U8996 ( .A(n7362), .ZN(n10278) );
  OAI22_X1 U8997 ( .A1(n10278), .A2(n8715), .B1(n7361), .B2(n8639), .ZN(n10280) );
  AOI21_X1 U8998 ( .B1(n10257), .B2(P2_REG3_REG_0__SCAN_IN), .A(n10280), .ZN(
        n7366) );
  INV_X1 U8999 ( .A(n8742), .ZN(n8615) );
  AOI22_X1 U9000 ( .A1(n7362), .A2(n8615), .B1(P2_REG2_REG_0__SCAN_IN), .B2(
        n10266), .ZN(n7365) );
  INV_X1 U9001 ( .A(n8550), .ZN(n8707) );
  OAI21_X1 U9002 ( .B1(n8707), .B2(n8486), .A(n7363), .ZN(n7364) );
  OAI211_X1 U9003 ( .C1(n7366), .C2(n10266), .A(n7365), .B(n7364), .ZN(
        P2_U3296) );
  NAND2_X1 U9004 ( .A1(n7368), .A2(n7367), .ZN(n7370) );
  NAND2_X1 U9005 ( .A1(n8223), .A2(n7034), .ZN(n7369) );
  NAND2_X1 U9006 ( .A1(n7370), .A2(n7369), .ZN(n7410) );
  NAND2_X1 U9007 ( .A1(n7372), .A2(n10302), .ZN(n7373) );
  NOR2_X1 U9008 ( .A1(n8380), .A2(n10259), .ZN(n7375) );
  OR2_X1 U9009 ( .A1(n10251), .A2(n10317), .ZN(n7374) );
  XNOR2_X1 U9010 ( .A(n7456), .B(n7455), .ZN(n7434) );
  XNOR2_X1 U9011 ( .A(n7376), .B(n7455), .ZN(n7378) );
  OAI21_X1 U9012 ( .B1(n7378), .B2(n8715), .A(n7377), .ZN(n7431) );
  INV_X1 U9013 ( .A(n7431), .ZN(n7379) );
  MUX2_X1 U9014 ( .A(n7084), .B(n7379), .S(n10263), .Z(n7385) );
  OR2_X1 U9015 ( .A1(n10259), .A2(n10244), .ZN(n7380) );
  AOI211_X1 U9016 ( .C1(n7453), .C2(n10248), .A(n10336), .B(n7463), .ZN(n7432)
         );
  OAI22_X1 U9017 ( .A1(n8733), .A2(n7382), .B1(n8620), .B2(n7381), .ZN(n7383)
         );
  AOI21_X1 U9018 ( .B1(n7432), .B2(n8719), .A(n7383), .ZN(n7384) );
  OAI211_X1 U9019 ( .C1(n8742), .C2(n7434), .A(n7385), .B(n7384), .ZN(P2_U3290) );
  NAND2_X1 U9020 ( .A1(n7386), .A2(n7393), .ZN(n7387) );
  NAND2_X1 U9021 ( .A1(n7388), .A2(n7387), .ZN(n10168) );
  NAND2_X1 U9022 ( .A1(n10124), .A2(n6563), .ZN(n7389) );
  NAND2_X1 U9023 ( .A1(n7390), .A2(n7389), .ZN(n10165) );
  INV_X1 U9024 ( .A(n10151), .ZN(n10135) );
  AOI22_X1 U9025 ( .A1(n9343), .A2(n6563), .B1(n10135), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n7391) );
  OAI21_X1 U9026 ( .B1(n10146), .B2(n10165), .A(n7391), .ZN(n7400) );
  NAND2_X1 U9027 ( .A1(n10168), .A2(n8040), .ZN(n7398) );
  AOI22_X1 U9028 ( .A1(n9020), .A2(n9370), .B1(n9368), .B2(n6552), .ZN(n7397)
         );
  OAI21_X1 U9029 ( .B1(n7394), .B2(n7393), .A(n7392), .ZN(n7395) );
  NAND2_X1 U9030 ( .A1(n7395), .A2(n10133), .ZN(n7396) );
  NAND3_X1 U9031 ( .A1(n7398), .A2(n7397), .A3(n7396), .ZN(n10166) );
  MUX2_X1 U9032 ( .A(n10166), .B(P1_REG2_REG_2__SCAN_IN), .S(n9242), .Z(n7399)
         );
  AOI211_X1 U9033 ( .C1(n10140), .C2(n10168), .A(n7400), .B(n7399), .ZN(n7401)
         );
  INV_X1 U9034 ( .A(n7401), .ZN(P1_U3289) );
  OAI21_X1 U9035 ( .B1(n7404), .B2(n7402), .A(n7403), .ZN(n7405) );
  NAND2_X1 U9036 ( .A1(n7405), .A2(n8956), .ZN(n7409) );
  OAI22_X1 U9037 ( .A1(n7539), .A2(n8960), .B1(n8981), .B2(n7544), .ZN(n7406)
         );
  AOI211_X1 U9038 ( .C1(n10176), .C2(n9007), .A(n7407), .B(n7406), .ZN(n7408)
         );
  OAI211_X1 U9039 ( .C1(n9005), .C2(n9377), .A(n7409), .B(n7408), .ZN(P1_U3225) );
  XNOR2_X1 U9040 ( .A(n7411), .B(n7413), .ZN(n10299) );
  XNOR2_X1 U9041 ( .A(n7413), .B(n7412), .ZN(n7415) );
  OAI22_X1 U9042 ( .A1(n8223), .A2(n8637), .B1(n7414), .B2(n8639), .ZN(n8227)
         );
  AOI21_X1 U9043 ( .B1(n7415), .B2(n10254), .A(n8227), .ZN(n10301) );
  INV_X1 U9044 ( .A(n10301), .ZN(n7422) );
  AOI21_X1 U9045 ( .B1(n7416), .B2(n8226), .A(n10336), .ZN(n7417) );
  NAND2_X1 U9046 ( .A1(n7417), .A2(n10245), .ZN(n10300) );
  OAI22_X1 U9047 ( .A1(n10263), .A2(n7418), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n8620), .ZN(n7419) );
  AOI21_X1 U9048 ( .B1(n8486), .B2(n8226), .A(n7419), .ZN(n7420) );
  OAI21_X1 U9049 ( .B1(n10300), .B2(n8561), .A(n7420), .ZN(n7421) );
  AOI21_X1 U9050 ( .B1(n7422), .B2(n10263), .A(n7421), .ZN(n7423) );
  OAI21_X1 U9051 ( .B1(n8742), .B2(n10299), .A(n7423), .ZN(P2_U3293) );
  NAND3_X1 U9052 ( .A1(n7426), .A2(n7425), .A3(n7424), .ZN(n7428) );
  NOR2_X1 U9053 ( .A1(n7428), .A2(n7427), .ZN(n7438) );
  INV_X1 U9054 ( .A(n7437), .ZN(n7429) );
  AND2_X2 U9055 ( .A1(n7438), .A2(n7429), .ZN(n10344) );
  INV_X1 U9056 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n7436) );
  AND2_X1 U9057 ( .A1(n7491), .A2(n4781), .ZN(n7430) );
  NAND2_X1 U9058 ( .A1(n7661), .A2(n7430), .ZN(n8831) );
  NAND2_X1 U9059 ( .A1(n10298), .A2(n8831), .ZN(n10340) );
  INV_X1 U9060 ( .A(n10340), .ZN(n10288) );
  INV_X1 U9061 ( .A(n10335), .ZN(n10284) );
  AOI211_X1 U9062 ( .C1(n10284), .C2(n7453), .A(n7432), .B(n7431), .ZN(n7433)
         );
  OAI21_X1 U9063 ( .B1(n10288), .B2(n7434), .A(n7433), .ZN(n7439) );
  NAND2_X1 U9064 ( .A1(n7439), .A2(n10344), .ZN(n7435) );
  OAI21_X1 U9065 ( .B1(n10344), .B2(n7436), .A(n7435), .ZN(P2_U3469) );
  AND2_X2 U9066 ( .A1(n7438), .A2(n7437), .ZN(n10360) );
  NAND2_X1 U9067 ( .A1(n7439), .A2(n10360), .ZN(n7440) );
  OAI21_X1 U9068 ( .B1(n10360), .B2(n7441), .A(n7440), .ZN(P2_U3526) );
  XOR2_X1 U9069 ( .A(n7442), .B(n7444), .Z(n10307) );
  INV_X1 U9070 ( .A(n7443), .ZN(n7448) );
  AOI21_X1 U9071 ( .B1(n7445), .B2(n7444), .A(n8715), .ZN(n7447) );
  AOI21_X1 U9072 ( .B1(n7447), .B2(n10250), .A(n7446), .ZN(n10310) );
  OAI21_X1 U9073 ( .B1(n7448), .B2(n8620), .A(n10310), .ZN(n7451) );
  XNOR2_X1 U9074 ( .A(n10245), .B(n10244), .ZN(n10309) );
  AOI22_X1 U9075 ( .A1(n8486), .A2(n10244), .B1(n10266), .B2(
        P2_REG2_REG_4__SCAN_IN), .ZN(n7449) );
  OAI21_X1 U9076 ( .B1(n10309), .B2(n8550), .A(n7449), .ZN(n7450) );
  AOI21_X1 U9077 ( .B1(n7451), .B2(n10263), .A(n7450), .ZN(n7452) );
  OAI21_X1 U9078 ( .B1(n10307), .B2(n8742), .A(n7452), .ZN(P2_U3292) );
  INV_X1 U9079 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n7468) );
  AND2_X1 U9080 ( .A1(n8379), .A2(n7453), .ZN(n7454) );
  AOI21_X1 U9081 ( .B1(n7456), .B2(n7455), .A(n7454), .ZN(n7590) );
  XNOR2_X1 U9082 ( .A(n7590), .B(n5241), .ZN(n7588) );
  AOI21_X1 U9083 ( .B1(n7457), .B2(n7589), .A(n8715), .ZN(n7462) );
  OAI22_X1 U9084 ( .A1(n7459), .A2(n8639), .B1(n7458), .B2(n8637), .ZN(n7460)
         );
  AOI21_X1 U9085 ( .B1(n7462), .B2(n7461), .A(n7460), .ZN(n7583) );
  INV_X1 U9086 ( .A(n7591), .ZN(n7465) );
  INV_X1 U9087 ( .A(n7463), .ZN(n7464) );
  AOI21_X1 U9088 ( .B1(n7465), .B2(n7464), .A(n4699), .ZN(n7586) );
  AOI22_X1 U9089 ( .A1(n7586), .A2(n10246), .B1(n10284), .B2(n7465), .ZN(n7466) );
  OAI211_X1 U9090 ( .C1(n7588), .C2(n10288), .A(n7583), .B(n7466), .ZN(n7469)
         );
  NAND2_X1 U9091 ( .A1(n7469), .A2(n10344), .ZN(n7467) );
  OAI21_X1 U9092 ( .B1(n10344), .B2(n7468), .A(n7467), .ZN(P2_U3472) );
  NAND2_X1 U9093 ( .A1(n7469), .A2(n10360), .ZN(n7470) );
  OAI21_X1 U9094 ( .B1(n10360), .B2(n7060), .A(n7470), .ZN(P2_U3527) );
  INV_X1 U9095 ( .A(n7672), .ZN(n7665) );
  INV_X1 U9096 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n7471) );
  MUX2_X1 U9097 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n7471), .S(n8407), .Z(n8409)
         );
  OAI21_X1 U9098 ( .B1(n7473), .B2(n7284), .A(n7472), .ZN(n8410) );
  NAND2_X1 U9099 ( .A1(n8409), .A2(n8410), .ZN(n8408) );
  INV_X1 U9100 ( .A(n8408), .ZN(n7474) );
  AOI21_X1 U9101 ( .B1(n8407), .B2(P2_REG1_REG_11__SCAN_IN), .A(n7474), .ZN(
        n7477) );
  INV_X1 U9102 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n10358) );
  MUX2_X1 U9103 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n10358), .S(n7672), .Z(n7476) );
  AND2_X1 U9104 ( .A1(n7477), .A2(n7476), .ZN(n7664) );
  INV_X1 U9105 ( .A(n7664), .ZN(n7475) );
  OAI21_X1 U9106 ( .B1(n7477), .B2(n7476), .A(n7475), .ZN(n7481) );
  NAND2_X1 U9107 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3152), .ZN(n7913) );
  INV_X1 U9108 ( .A(n7913), .ZN(n7480) );
  INV_X1 U9109 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7478) );
  NOR2_X1 U9110 ( .A1(n8481), .A2(n7478), .ZN(n7479) );
  AOI211_X1 U9111 ( .C1(n10232), .C2(n7481), .A(n7480), .B(n7479), .ZN(n7489)
         );
  INV_X1 U9112 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7482) );
  XNOR2_X1 U9113 ( .A(n7672), .B(n7482), .ZN(n7487) );
  OR2_X1 U9114 ( .A1(n8407), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n7485) );
  INV_X1 U9115 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7771) );
  MUX2_X1 U9116 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n7771), .S(n8407), .Z(n8404)
         );
  OAI211_X1 U9117 ( .C1(n7487), .C2(n7486), .A(n10233), .B(n7674), .ZN(n7488)
         );
  OAI211_X1 U9118 ( .C1(n10235), .C2(n7665), .A(n7489), .B(n7488), .ZN(
        P2_U3257) );
  INV_X1 U9119 ( .A(n7490), .ZN(n7523) );
  OAI222_X1 U9120 ( .A1(n8876), .A2(n7492), .B1(n8871), .B2(n7523), .C1(n7491), 
        .C2(P2_U3152), .ZN(P2_U3338) );
  INV_X1 U9121 ( .A(n7493), .ZN(n7494) );
  NAND2_X1 U9122 ( .A1(n7495), .A2(n7494), .ZN(n7496) );
  AND2_X1 U9123 ( .A1(n8378), .A2(n8168), .ZN(n7498) );
  XNOR2_X1 U9124 ( .A(n7591), .B(n8156), .ZN(n7499) );
  NAND2_X1 U9125 ( .A1(n7498), .A2(n7499), .ZN(n7512) );
  INV_X1 U9126 ( .A(n7498), .ZN(n7500) );
  INV_X1 U9127 ( .A(n7499), .ZN(n7511) );
  NAND2_X1 U9128 ( .A1(n7500), .A2(n7511), .ZN(n7501) );
  NAND2_X1 U9129 ( .A1(n7512), .A2(n7501), .ZN(n7504) );
  INV_X1 U9130 ( .A(n7513), .ZN(n7503) );
  AOI211_X1 U9131 ( .C1(n7505), .C2(n7504), .A(n8340), .B(n7503), .ZN(n7509)
         );
  INV_X1 U9132 ( .A(n8347), .ZN(n8334) );
  AOI22_X1 U9133 ( .A1(n8379), .A2(n8334), .B1(n7581), .B2(n8344), .ZN(n7507)
         );
  AOI22_X1 U9134 ( .A1(n8377), .A2(n8349), .B1(P2_REG3_REG_7__SCAN_IN), .B2(
        P2_U3152), .ZN(n7506) );
  OAI211_X1 U9135 ( .C1(n7591), .C2(n8366), .A(n7507), .B(n7506), .ZN(n7508)
         );
  OR2_X1 U9136 ( .A1(n7509), .A2(n7508), .ZN(P2_U3215) );
  NAND2_X1 U9137 ( .A1(n8377), .A2(n8168), .ZN(n7646) );
  XNOR2_X1 U9138 ( .A(n7680), .B(n7953), .ZN(n7647) );
  XNOR2_X1 U9139 ( .A(n7646), .B(n7647), .ZN(n7514) );
  INV_X1 U9140 ( .A(n7514), .ZN(n7510) );
  AOI21_X1 U9141 ( .B1(n7513), .B2(n7510), .A(n8340), .ZN(n7517) );
  NOR3_X1 U9142 ( .A1(n7511), .A2(n7599), .A3(n8301), .ZN(n7516) );
  NAND2_X1 U9143 ( .A1(n7515), .A2(n7514), .ZN(n7650) );
  OAI21_X1 U9144 ( .B1(n7517), .B2(n7516), .A(n7650), .ZN(n7522) );
  NOR2_X1 U9145 ( .A1(n7599), .A2(n8347), .ZN(n7520) );
  OAI22_X1 U9146 ( .A1(n7807), .A2(n8321), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7518), .ZN(n7519) );
  AOI211_X1 U9147 ( .C1(n8344), .C2(n7608), .A(n7520), .B(n7519), .ZN(n7521)
         );
  OAI211_X1 U9148 ( .C1(n10321), .C2(n8366), .A(n7522), .B(n7521), .ZN(
        P2_U3223) );
  OAI222_X1 U9149 ( .A1(P1_U3084), .A2(n7524), .B1(n8155), .B2(n9793), .C1(
        n9492), .C2(n7523), .ZN(P1_U3333) );
  INV_X1 U9150 ( .A(n7624), .ZN(n7529) );
  INV_X1 U9151 ( .A(n7525), .ZN(n7526) );
  OAI21_X1 U9152 ( .B1(n7529), .B2(n7528), .A(n7616), .ZN(n7532) );
  OR2_X1 U9153 ( .A1(n7797), .A2(n9238), .ZN(n7531) );
  OR2_X1 U9154 ( .A1(n7544), .A2(n9236), .ZN(n7530) );
  NAND2_X1 U9155 ( .A1(n7531), .A2(n7530), .ZN(n7569) );
  AOI21_X1 U9156 ( .B1(n7532), .B2(n10133), .A(n7569), .ZN(n10191) );
  OAI22_X1 U9157 ( .A1(n10143), .A2(n6903), .B1(n7571), .B2(n10151), .ZN(n7536) );
  INV_X1 U9158 ( .A(n7630), .ZN(n7533) );
  OAI211_X1 U9159 ( .C1(n10192), .C2(n7698), .A(n7533), .B(n10125), .ZN(n10190) );
  OR2_X1 U9160 ( .A1(n7534), .A2(n10138), .ZN(n9325) );
  NOR2_X1 U9161 ( .A1(n10190), .A2(n9325), .ZN(n7535) );
  AOI211_X1 U9162 ( .C1(n9343), .C2(n7622), .A(n7536), .B(n7535), .ZN(n7550)
         );
  NAND2_X1 U9163 ( .A1(n7538), .A2(n7537), .ZN(n7541) );
  NAND2_X1 U9164 ( .A1(n7539), .A2(n6538), .ZN(n7540) );
  NAND2_X1 U9165 ( .A1(n7541), .A2(n7540), .ZN(n9381) );
  INV_X1 U9166 ( .A(n9381), .ZN(n7542) );
  NAND2_X1 U9167 ( .A1(n9019), .A2(n10176), .ZN(n7543) );
  NAND2_X1 U9168 ( .A1(n7544), .A2(n10184), .ZN(n7545) );
  XNOR2_X1 U9169 ( .A(n7625), .B(n7624), .ZN(n10194) );
  AND2_X1 U9170 ( .A1(n7547), .A2(n7546), .ZN(n7548) );
  NAND2_X1 U9171 ( .A1(n10143), .A2(n7548), .ZN(n9366) );
  INV_X1 U9172 ( .A(n9366), .ZN(n9382) );
  NAND2_X1 U9173 ( .A1(n10194), .A2(n9382), .ZN(n7549) );
  OAI211_X1 U9174 ( .C1(n10191), .C2(n9353), .A(n7550), .B(n7549), .ZN(
        P1_U3284) );
  NAND2_X1 U9175 ( .A1(n7552), .A2(n7551), .ZN(n7555) );
  AND2_X1 U9176 ( .A1(n7553), .A2(n7403), .ZN(n7554) );
  XOR2_X1 U9177 ( .A(n7555), .B(n7554), .Z(n7564) );
  INV_X1 U9178 ( .A(n7556), .ZN(n7700) );
  OR2_X1 U9179 ( .A1(n7557), .A2(n9238), .ZN(n7560) );
  OR2_X1 U9180 ( .A1(n7558), .A2(n9236), .ZN(n7559) );
  NAND2_X1 U9181 ( .A1(n7560), .A2(n7559), .ZN(n7705) );
  INV_X1 U9182 ( .A(n8915), .ZN(n9003) );
  AOI22_X1 U9183 ( .A1(n7705), .A2(n9003), .B1(P1_REG3_REG_6__SCAN_IN), .B2(
        P1_U3084), .ZN(n7561) );
  OAI21_X1 U9184 ( .B1(n10184), .B2(n8996), .A(n7561), .ZN(n7562) );
  AOI21_X1 U9185 ( .B1(n7700), .B2(n8962), .A(n7562), .ZN(n7563) );
  OAI21_X1 U9186 ( .B1(n7564), .B2(n9009), .A(n7563), .ZN(P1_U3237) );
  XOR2_X1 U9187 ( .A(n7566), .B(n7565), .Z(n7567) );
  XNOR2_X1 U9188 ( .A(n7568), .B(n7567), .ZN(n7574) );
  AOI22_X1 U9189 ( .A1(n7569), .A2(n9003), .B1(P1_REG3_REG_7__SCAN_IN), .B2(
        P1_U3084), .ZN(n7570) );
  OAI21_X1 U9190 ( .B1(n9005), .B2(n7571), .A(n7570), .ZN(n7572) );
  AOI21_X1 U9191 ( .B1(n7622), .B2(n9007), .A(n7572), .ZN(n7573) );
  OAI21_X1 U9192 ( .B1(n7574), .B2(n9009), .A(n7573), .ZN(P1_U3211) );
  INV_X1 U9193 ( .A(n7575), .ZN(n7579) );
  OAI222_X1 U9194 ( .A1(n9492), .A2(n7579), .B1(P1_U3084), .B2(n7577), .C1(
        n7576), .C2(n9489), .ZN(P1_U3332) );
  OAI222_X1 U9195 ( .A1(n8876), .A2(n7580), .B1(n8871), .B2(n7579), .C1(n7578), 
        .C2(P2_U3152), .ZN(P2_U3337) );
  AOI22_X1 U9196 ( .A1(n10266), .A2(P2_REG2_REG_7__SCAN_IN), .B1(n7581), .B2(
        n10257), .ZN(n7582) );
  OAI21_X1 U9197 ( .B1(n7591), .B2(n8733), .A(n7582), .ZN(n7585) );
  NOR2_X1 U9198 ( .A1(n7583), .A2(n10266), .ZN(n7584) );
  AOI211_X1 U9199 ( .C1(n7586), .C2(n8707), .A(n7585), .B(n7584), .ZN(n7587)
         );
  OAI21_X1 U9200 ( .B1(n7588), .B2(n8742), .A(n7587), .ZN(P2_U3289) );
  NAND2_X1 U9201 ( .A1(n7590), .A2(n7589), .ZN(n7593) );
  NAND2_X1 U9202 ( .A1(n7599), .A2(n7591), .ZN(n7592) );
  NAND2_X1 U9203 ( .A1(n7593), .A2(n7592), .ZN(n7594) );
  NAND2_X1 U9204 ( .A1(n7594), .A2(n7597), .ZN(n7595) );
  NAND2_X1 U9205 ( .A1(n7682), .A2(n7595), .ZN(n7603) );
  OAI21_X1 U9206 ( .B1(n7598), .B2(n7597), .A(n7596), .ZN(n7601) );
  OAI22_X1 U9207 ( .A1(n7599), .A2(n8637), .B1(n7807), .B2(n8639), .ZN(n7600)
         );
  AOI21_X1 U9208 ( .B1(n7601), .B2(n10254), .A(n7600), .ZN(n7602) );
  OAI21_X1 U9209 ( .B1(n7603), .B2(n10298), .A(n7602), .ZN(n10323) );
  INV_X1 U9210 ( .A(n10323), .ZN(n7613) );
  INV_X1 U9211 ( .A(n7603), .ZN(n10325) );
  INV_X1 U9212 ( .A(n7604), .ZN(n7605) );
  NAND2_X1 U9213 ( .A1(n10263), .A2(n7605), .ZN(n7826) );
  INV_X1 U9214 ( .A(n7826), .ZN(n8028) );
  NAND2_X1 U9215 ( .A1(n7606), .A2(n7680), .ZN(n7607) );
  NAND2_X1 U9216 ( .A1(n7685), .A2(n7607), .ZN(n10322) );
  AOI22_X1 U9217 ( .A1(n10266), .A2(P2_REG2_REG_8__SCAN_IN), .B1(n7608), .B2(
        n10257), .ZN(n7610) );
  NAND2_X1 U9218 ( .A1(n8486), .A2(n7680), .ZN(n7609) );
  OAI211_X1 U9219 ( .C1(n10322), .C2(n8550), .A(n7610), .B(n7609), .ZN(n7611)
         );
  AOI21_X1 U9220 ( .B1(n10325), .B2(n8028), .A(n7611), .ZN(n7612) );
  OAI21_X1 U9221 ( .B1(n7613), .B2(n10266), .A(n7612), .ZN(P2_U3288) );
  INV_X1 U9222 ( .A(n7779), .ZN(n7619) );
  NAND2_X1 U9223 ( .A1(n7616), .A2(n7615), .ZN(n7617) );
  NAND2_X1 U9224 ( .A1(n7617), .A2(n7626), .ZN(n7618) );
  OAI211_X1 U9225 ( .C1(n7780), .C2(n7619), .A(n7618), .B(n10133), .ZN(n7621)
         );
  AOI22_X1 U9226 ( .A1(n9018), .A2(n9368), .B1(n9370), .B2(n9016), .ZN(n7620)
         );
  NAND2_X1 U9227 ( .A1(n7621), .A2(n7620), .ZN(n10201) );
  INV_X1 U9228 ( .A(n10201), .ZN(n7635) );
  NOR2_X1 U9229 ( .A1(n9018), .A2(n7622), .ZN(n7623) );
  NOR2_X1 U9230 ( .A1(n7627), .A2(n7626), .ZN(n10198) );
  INV_X1 U9231 ( .A(n10198), .ZN(n7628) );
  NAND3_X1 U9232 ( .A1(n7628), .A2(n9382), .A3(n10203), .ZN(n7634) );
  OAI22_X1 U9233 ( .A1(n10143), .A2(n7629), .B1(n7642), .B2(n10151), .ZN(n7632) );
  NAND2_X1 U9234 ( .A1(n7630), .A2(n10199), .ZN(n7786) );
  OAI21_X1 U9235 ( .B1(n7630), .B2(n10199), .A(n7786), .ZN(n10200) );
  NOR2_X1 U9236 ( .A1(n10200), .A2(n10146), .ZN(n7631) );
  AOI211_X1 U9237 ( .C1(n9343), .C2(n7777), .A(n7632), .B(n7631), .ZN(n7633)
         );
  OAI211_X1 U9238 ( .C1(n9242), .C2(n7635), .A(n7634), .B(n7633), .ZN(P1_U3283) );
  XOR2_X1 U9239 ( .A(n7637), .B(n7636), .Z(n7638) );
  XNOR2_X1 U9240 ( .A(n7639), .B(n7638), .ZN(n7645) );
  INV_X1 U9241 ( .A(n8960), .ZN(n8983) );
  AOI22_X1 U9242 ( .A1(n8983), .A2(n9018), .B1(P1_REG3_REG_8__SCAN_IN), .B2(
        P1_U3084), .ZN(n7641) );
  INV_X1 U9243 ( .A(n8981), .ZN(n8971) );
  NAND2_X1 U9244 ( .A1(n8971), .A2(n9016), .ZN(n7640) );
  OAI211_X1 U9245 ( .C1(n9005), .C2(n7642), .A(n7641), .B(n7640), .ZN(n7643)
         );
  AOI21_X1 U9246 ( .B1(n7777), .B2(n9007), .A(n7643), .ZN(n7644) );
  OAI21_X1 U9247 ( .B1(n7645), .B2(n9009), .A(n7644), .ZN(P1_U3219) );
  INV_X1 U9248 ( .A(n7646), .ZN(n7648) );
  NAND2_X1 U9249 ( .A1(n7648), .A2(n7647), .ZN(n7649) );
  OR2_X1 U9250 ( .A1(n7807), .A2(n8243), .ZN(n7651) );
  XNOR2_X1 U9251 ( .A(n7839), .B(n8156), .ZN(n7739) );
  NOR2_X1 U9252 ( .A1(n7651), .A2(n7739), .ZN(n7738) );
  NAND2_X1 U9253 ( .A1(n7651), .A2(n7739), .ZN(n7742) );
  XNOR2_X1 U9254 ( .A(n7823), .B(n8156), .ZN(n7750) );
  OR2_X1 U9255 ( .A1(n7768), .A2(n8243), .ZN(n7749) );
  XNOR2_X1 U9256 ( .A(n7750), .B(n7749), .ZN(n7754) );
  XNOR2_X1 U9257 ( .A(n7755), .B(n7754), .ZN(n7657) );
  OAI22_X1 U9258 ( .A1(n7926), .A2(n8321), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7652), .ZN(n7655) );
  INV_X1 U9259 ( .A(n7653), .ZN(n7816) );
  OAI22_X1 U9260 ( .A1(n7807), .A2(n8347), .B1(n8360), .B2(n7816), .ZN(n7654)
         );
  AOI211_X1 U9261 ( .C1(n7823), .C2(n8324), .A(n7655), .B(n7654), .ZN(n7656)
         );
  OAI21_X1 U9262 ( .B1(n7657), .B2(n8340), .A(n7656), .ZN(P2_U3219) );
  INV_X1 U9263 ( .A(n7658), .ZN(n7662) );
  OAI222_X1 U9264 ( .A1(n7660), .A2(P1_U3084), .B1(n9492), .B2(n7662), .C1(
        n7659), .C2(n8155), .ZN(P1_U3331) );
  OAI222_X1 U9265 ( .A1(n8876), .A2(n7663), .B1(n8871), .B2(n7662), .C1(
        P2_U3152), .C2(n7661), .ZN(P2_U3336) );
  NAND2_X1 U9266 ( .A1(P2_U3152), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n7966) );
  INV_X1 U9267 ( .A(n7966), .ZN(n7670) );
  AOI21_X1 U9268 ( .B1(n10358), .B2(n7665), .A(n7664), .ZN(n7667) );
  INV_X1 U9269 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n7720) );
  AOI22_X1 U9270 ( .A1(n7726), .A2(n7720), .B1(P2_REG1_REG_13__SCAN_IN), .B2(
        n7721), .ZN(n7666) );
  NOR2_X1 U9271 ( .A1(n7667), .A2(n7666), .ZN(n7719) );
  AOI21_X1 U9272 ( .B1(n7667), .B2(n7666), .A(n7719), .ZN(n7668) );
  NOR2_X1 U9273 ( .A1(n10236), .A2(n7668), .ZN(n7669) );
  AOI211_X1 U9274 ( .C1(P2_ADDR_REG_13__SCAN_IN), .C2(n10234), .A(n7670), .B(
        n7669), .ZN(n7679) );
  NOR2_X1 U9275 ( .A1(n7726), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n7671) );
  AOI21_X1 U9276 ( .B1(P2_REG2_REG_13__SCAN_IN), .B2(n7726), .A(n7671), .ZN(
        n7676) );
  NAND2_X1 U9277 ( .A1(n7672), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n7673) );
  OAI21_X1 U9278 ( .B1(n7676), .B2(n7675), .A(n7725), .ZN(n7677) );
  NAND2_X1 U9279 ( .A1(n10233), .A2(n7677), .ZN(n7678) );
  OAI211_X1 U9280 ( .C1(n10235), .C2(n7721), .A(n7679), .B(n7678), .ZN(
        P2_U3258) );
  NAND2_X1 U9281 ( .A1(n8377), .A2(n7680), .ZN(n7681) );
  XOR2_X1 U9282 ( .A(n7762), .B(n7763), .Z(n7841) );
  XOR2_X1 U9283 ( .A(n7683), .B(n7762), .Z(n7684) );
  AOI22_X1 U9284 ( .A1(n8375), .A2(n8702), .B1(n8700), .B2(n8377), .ZN(n7737)
         );
  OAI21_X1 U9285 ( .B1(n7684), .B2(n8715), .A(n7737), .ZN(n7837) );
  NOR2_X2 U9286 ( .A1(n7685), .A2(n7839), .ZN(n7818) );
  NAND2_X1 U9287 ( .A1(n7685), .A2(n7839), .ZN(n7686) );
  NAND2_X1 U9288 ( .A1(n7686), .A2(n10246), .ZN(n7687) );
  NOR2_X1 U9289 ( .A1(n7818), .A2(n7687), .ZN(n7838) );
  NAND2_X1 U9290 ( .A1(n7838), .A2(n8719), .ZN(n7692) );
  INV_X1 U9291 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7689) );
  OAI22_X1 U9292 ( .A1(n10263), .A2(n7689), .B1(n7688), .B2(n8620), .ZN(n7690)
         );
  AOI21_X1 U9293 ( .B1(n8486), .B2(n7839), .A(n7690), .ZN(n7691) );
  NAND2_X1 U9294 ( .A1(n7692), .A2(n7691), .ZN(n7693) );
  AOI21_X1 U9295 ( .B1(n7837), .B2(n10263), .A(n7693), .ZN(n7694) );
  OAI21_X1 U9296 ( .B1(n8742), .B2(n7841), .A(n7694), .ZN(P2_U3287) );
  OAI21_X1 U9297 ( .B1(n7697), .B2(n7696), .A(n7695), .ZN(n10188) );
  AND2_X1 U9298 ( .A1(n9374), .A2(n7701), .ZN(n7699) );
  OR2_X1 U9299 ( .A1(n7699), .A2(n7698), .ZN(n10185) );
  AOI22_X1 U9300 ( .A1(n9343), .A2(n7701), .B1(n7700), .B2(n10135), .ZN(n7702)
         );
  OAI21_X1 U9301 ( .B1(n10185), .B2(n10146), .A(n7702), .ZN(n7710) );
  XNOR2_X1 U9302 ( .A(n7704), .B(n7703), .ZN(n7708) );
  NAND2_X1 U9303 ( .A1(n10188), .A2(n8040), .ZN(n7707) );
  INV_X1 U9304 ( .A(n7705), .ZN(n7706) );
  OAI211_X1 U9305 ( .C1(n9356), .C2(n7708), .A(n7707), .B(n7706), .ZN(n10186)
         );
  MUX2_X1 U9306 ( .A(n10186), .B(P1_REG2_REG_6__SCAN_IN), .S(n9242), .Z(n7709)
         );
  AOI211_X1 U9307 ( .C1(n10140), .C2(n10188), .A(n7710), .B(n7709), .ZN(n7711)
         );
  INV_X1 U9308 ( .A(n7711), .ZN(P1_U3285) );
  NAND2_X1 U9309 ( .A1(n7715), .A2(n8103), .ZN(n7713) );
  OAI211_X1 U9310 ( .C1(n7714), .C2(n8155), .A(n7713), .B(n7712), .ZN(P1_U3330) );
  NAND2_X1 U9311 ( .A1(n7715), .A2(n8132), .ZN(n7717) );
  OAI211_X1 U9312 ( .C1(n7718), .C2(n8865), .A(n7717), .B(n7716), .ZN(P2_U3335) );
  AOI21_X1 U9313 ( .B1(n7721), .B2(n7720), .A(n7719), .ZN(n7723) );
  INV_X1 U9314 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n9915) );
  AOI22_X1 U9315 ( .A1(n7972), .A2(n9915), .B1(P2_REG1_REG_14__SCAN_IN), .B2(
        n7976), .ZN(n7722) );
  NOR2_X1 U9316 ( .A1(n7723), .A2(n7722), .ZN(n7975) );
  AOI21_X1 U9317 ( .B1(n7723), .B2(n7722), .A(n7975), .ZN(n7734) );
  INV_X1 U9318 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n7724) );
  AOI22_X1 U9319 ( .A1(n7972), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n7724), .B2(
        n7976), .ZN(n7728) );
  NAND2_X1 U9320 ( .A1(n7728), .A2(n7727), .ZN(n7971) );
  OAI21_X1 U9321 ( .B1(n7728), .B2(n7727), .A(n7971), .ZN(n7732) );
  INV_X1 U9322 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7730) );
  NAND2_X1 U9323 ( .A1(n9897), .A2(n7972), .ZN(n7729) );
  NAND2_X1 U9324 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3152), .ZN(n8093) );
  OAI211_X1 U9325 ( .C1(n8481), .C2(n7730), .A(n7729), .B(n8093), .ZN(n7731)
         );
  AOI21_X1 U9326 ( .B1(n7732), .B2(n10233), .A(n7731), .ZN(n7733) );
  OAI21_X1 U9327 ( .B1(n7734), .B2(n10236), .A(n7733), .ZN(P2_U3259) );
  AOI22_X1 U9328 ( .A1(n8344), .A2(n7735), .B1(P2_REG3_REG_9__SCAN_IN), .B2(
        P2_U3152), .ZN(n7736) );
  OAI21_X1 U9329 ( .B1(n7737), .B2(n8291), .A(n7736), .ZN(n7747) );
  NOR3_X1 U9330 ( .A1(n7738), .A2(n4864), .A3(n8340), .ZN(n7745) );
  INV_X1 U9331 ( .A(n7739), .ZN(n7740) );
  NAND3_X1 U9332 ( .A1(n8376), .A2(n7740), .A3(n8352), .ZN(n7741) );
  OAI21_X1 U9333 ( .B1(n7742), .B2(n8340), .A(n7741), .ZN(n7744) );
  MUX2_X1 U9334 ( .A(n7745), .B(n7744), .S(n7743), .Z(n7746) );
  AOI211_X1 U9335 ( .C1(n7839), .C2(n8324), .A(n7747), .B(n7746), .ZN(n7748)
         );
  INV_X1 U9336 ( .A(n7748), .ZN(P2_U3233) );
  INV_X1 U9337 ( .A(n7749), .ZN(n7752) );
  INV_X1 U9338 ( .A(n7750), .ZN(n7751) );
  NAND2_X1 U9339 ( .A1(n7752), .A2(n7751), .ZN(n7753) );
  XNOR2_X1 U9340 ( .A(n8840), .B(n8156), .ZN(n7908) );
  NOR2_X1 U9341 ( .A1(n7926), .A2(n8243), .ZN(n7909) );
  XNOR2_X1 U9342 ( .A(n7908), .B(n7909), .ZN(n7906) );
  XNOR2_X1 U9343 ( .A(n7907), .B(n7906), .ZN(n7760) );
  OAI22_X1 U9344 ( .A1(n8008), .A2(n8321), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5317), .ZN(n7758) );
  INV_X1 U9345 ( .A(n7756), .ZN(n7770) );
  OAI22_X1 U9346 ( .A1(n7768), .A2(n8347), .B1(n8360), .B2(n7770), .ZN(n7757)
         );
  AOI211_X1 U9347 ( .C1(n8840), .C2(n8324), .A(n7758), .B(n7757), .ZN(n7759)
         );
  OAI21_X1 U9348 ( .B1(n7760), .B2(n8340), .A(n7759), .ZN(P2_U3238) );
  NAND2_X1 U9349 ( .A1(n8375), .A2(n7823), .ZN(n7764) );
  XNOR2_X1 U9350 ( .A(n7921), .B(n7920), .ZN(n8842) );
  XNOR2_X1 U9351 ( .A(n7766), .B(n7765), .ZN(n7767) );
  OAI222_X1 U9352 ( .A1(n8639), .A2(n8008), .B1(n8637), .B2(n7768), .C1(n8715), 
        .C2(n7767), .ZN(n8838) );
  NAND2_X1 U9353 ( .A1(n7818), .A2(n10328), .ZN(n7820) );
  AOI21_X1 U9354 ( .B1(n7820), .B2(n8840), .A(n10336), .ZN(n7769) );
  AND2_X1 U9355 ( .A1(n7769), .A2(n7927), .ZN(n8839) );
  NAND2_X1 U9356 ( .A1(n8839), .A2(n8719), .ZN(n7774) );
  OAI22_X1 U9357 ( .A1(n10263), .A2(n7771), .B1(n7770), .B2(n8620), .ZN(n7772)
         );
  AOI21_X1 U9358 ( .B1(n8840), .B2(n8486), .A(n7772), .ZN(n7773) );
  NAND2_X1 U9359 ( .A1(n7774), .A2(n7773), .ZN(n7775) );
  AOI21_X1 U9360 ( .B1(n8838), .B2(n10263), .A(n7775), .ZN(n7776) );
  OAI21_X1 U9361 ( .B1(n8742), .B2(n8842), .A(n7776), .ZN(P2_U3285) );
  NAND2_X1 U9362 ( .A1(n9017), .A2(n7777), .ZN(n7778) );
  NAND2_X1 U9363 ( .A1(n10203), .A2(n7778), .ZN(n7852) );
  XOR2_X1 U9364 ( .A(n7852), .B(n7781), .Z(n10206) );
  NAND2_X1 U9365 ( .A1(n7780), .A2(n7779), .ZN(n7847) );
  XOR2_X1 U9366 ( .A(n7781), .B(n7847), .Z(n7783) );
  OAI22_X1 U9367 ( .A1(n7797), .A2(n9236), .B1(n7890), .B2(n9238), .ZN(n7782)
         );
  AOI21_X1 U9368 ( .B1(n7783), .B2(n10133), .A(n7782), .ZN(n7784) );
  OAI21_X1 U9369 ( .B1(n10206), .B2(n10130), .A(n7784), .ZN(n10211) );
  NAND2_X1 U9370 ( .A1(n10211), .A2(n10143), .ZN(n7791) );
  OAI22_X1 U9371 ( .A1(n10143), .A2(n7785), .B1(n7800), .B2(n10151), .ZN(n7789) );
  NAND2_X1 U9372 ( .A1(n7786), .A2(n7853), .ZN(n7787) );
  NAND2_X1 U9373 ( .A1(n7864), .A2(n7787), .ZN(n10210) );
  NOR2_X1 U9374 ( .A1(n10210), .A2(n10146), .ZN(n7788) );
  AOI211_X1 U9375 ( .C1(n9343), .C2(n7853), .A(n7789), .B(n7788), .ZN(n7790)
         );
  OAI211_X1 U9376 ( .C1(n10206), .C2(n9346), .A(n7791), .B(n7790), .ZN(
        P1_U3282) );
  INV_X1 U9377 ( .A(n7792), .ZN(n7793) );
  AOI21_X1 U9378 ( .B1(n7795), .B2(n7794), .A(n7793), .ZN(n7803) );
  NOR2_X1 U9379 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7796), .ZN(n10014) );
  NOR2_X1 U9380 ( .A1(n8960), .A2(n7797), .ZN(n7798) );
  AOI211_X1 U9381 ( .C1(n8971), .C2(n9015), .A(n10014), .B(n7798), .ZN(n7799)
         );
  OAI21_X1 U9382 ( .B1(n9005), .B2(n7800), .A(n7799), .ZN(n7801) );
  AOI21_X1 U9383 ( .B1(n7853), .B2(n9007), .A(n7801), .ZN(n7802) );
  OAI21_X1 U9384 ( .B1(n7803), .B2(n9009), .A(n7802), .ZN(P1_U3229) );
  NAND2_X1 U9385 ( .A1(n7804), .A2(n7812), .ZN(n7805) );
  NAND2_X1 U9386 ( .A1(n7806), .A2(n7805), .ZN(n10327) );
  OAI22_X1 U9387 ( .A1(n7807), .A2(n8637), .B1(n7926), .B2(n8639), .ZN(n7808)
         );
  INV_X1 U9388 ( .A(n7808), .ZN(n7815) );
  AND2_X1 U9389 ( .A1(n7810), .A2(n7809), .ZN(n7813) );
  OAI211_X1 U9390 ( .C1(n7813), .C2(n7812), .A(n7811), .B(n10254), .ZN(n7814)
         );
  OAI211_X1 U9391 ( .C1(n10327), .C2(n10298), .A(n7815), .B(n7814), .ZN(n10330) );
  NAND2_X1 U9392 ( .A1(n10330), .A2(n10263), .ZN(n7825) );
  INV_X1 U9393 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7817) );
  OAI22_X1 U9394 ( .A1(n10263), .A2(n7817), .B1(n7816), .B2(n8620), .ZN(n7822)
         );
  OR2_X1 U9395 ( .A1(n7818), .A2(n10328), .ZN(n7819) );
  NAND2_X1 U9396 ( .A1(n7820), .A2(n7819), .ZN(n10329) );
  NOR2_X1 U9397 ( .A1(n10329), .A2(n8550), .ZN(n7821) );
  AOI211_X1 U9398 ( .C1(n8486), .C2(n7823), .A(n7822), .B(n7821), .ZN(n7824)
         );
  OAI211_X1 U9399 ( .C1(n10327), .C2(n7826), .A(n7825), .B(n7824), .ZN(
        P2_U3286) );
  NAND2_X1 U9400 ( .A1(n7828), .A2(n7827), .ZN(n7829) );
  XNOR2_X1 U9401 ( .A(n7830), .B(n7829), .ZN(n7836) );
  OAI22_X1 U9402 ( .A1(n7832), .A2(n9236), .B1(n7831), .B2(n9238), .ZN(n7849)
         );
  AOI22_X1 U9403 ( .A1(n7849), .A2(n9003), .B1(P1_REG3_REG_10__SCAN_IN), .B2(
        P1_U3084), .ZN(n7833) );
  OAI21_X1 U9404 ( .B1(n9005), .B2(n7861), .A(n7833), .ZN(n7834) );
  AOI21_X1 U9405 ( .B1(n7881), .B2(n9007), .A(n7834), .ZN(n7835) );
  OAI21_X1 U9406 ( .B1(n7836), .B2(n9009), .A(n7835), .ZN(P1_U3215) );
  INV_X1 U9407 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n7843) );
  AOI211_X1 U9408 ( .C1(n10284), .C2(n7839), .A(n7838), .B(n7837), .ZN(n7840)
         );
  OAI21_X1 U9409 ( .B1(n10288), .B2(n7841), .A(n7840), .ZN(n7844) );
  NAND2_X1 U9410 ( .A1(n7844), .A2(n10344), .ZN(n7842) );
  OAI21_X1 U9411 ( .B1(n10344), .B2(n7843), .A(n7842), .ZN(P2_U3478) );
  NAND2_X1 U9412 ( .A1(n7844), .A2(n10360), .ZN(n7845) );
  OAI21_X1 U9413 ( .B1(n10360), .B2(n8392), .A(n7845), .ZN(P2_U3529) );
  XNOR2_X1 U9414 ( .A(n7888), .B(n7860), .ZN(n7850) );
  AOI21_X1 U9415 ( .B1(n7850), .B2(n10133), .A(n7849), .ZN(n7875) );
  OR2_X1 U9416 ( .A1(n9016), .A2(n7853), .ZN(n7851) );
  NAND2_X1 U9417 ( .A1(n7852), .A2(n7851), .ZN(n7855) );
  NAND2_X1 U9418 ( .A1(n7853), .A2(n9016), .ZN(n7854) );
  NAND2_X1 U9419 ( .A1(n7855), .A2(n7854), .ZN(n7856) );
  INV_X1 U9420 ( .A(n7856), .ZN(n7858) );
  INV_X1 U9421 ( .A(n7860), .ZN(n7857) );
  INV_X1 U9422 ( .A(n7883), .ZN(n7859) );
  AOI21_X1 U9423 ( .B1(n7860), .B2(n7856), .A(n7859), .ZN(n7876) );
  OAI22_X1 U9424 ( .A1(n10143), .A2(n7862), .B1(n7861), .B2(n10151), .ZN(n7863) );
  AOI21_X1 U9425 ( .B1(n7881), .B2(n9343), .A(n7863), .ZN(n7868) );
  NAND2_X1 U9426 ( .A1(n7864), .A2(n7881), .ZN(n7865) );
  NAND2_X1 U9427 ( .A1(n7865), .A2(n10125), .ZN(n7866) );
  NOR2_X1 U9428 ( .A1(n7895), .A2(n7866), .ZN(n7873) );
  INV_X1 U9429 ( .A(n9325), .ZN(n9364) );
  NAND2_X1 U9430 ( .A1(n7873), .A2(n9364), .ZN(n7867) );
  OAI211_X1 U9431 ( .C1(n7876), .C2(n9366), .A(n7868), .B(n7867), .ZN(n7869)
         );
  INV_X1 U9432 ( .A(n7869), .ZN(n7870) );
  OAI21_X1 U9433 ( .B1(n9353), .B2(n7875), .A(n7870), .ZN(P1_U3281) );
  INV_X1 U9434 ( .A(n5962), .ZN(n7918) );
  OAI222_X1 U9435 ( .A1(P2_U3152), .A2(n7872), .B1(n8871), .B2(n7918), .C1(
        n7871), .C2(n8865), .ZN(P2_U3334) );
  INV_X1 U9436 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n7878) );
  NAND2_X1 U9437 ( .A1(n10130), .A2(n9931), .ZN(n10195) );
  INV_X1 U9438 ( .A(n10195), .ZN(n10197) );
  AOI21_X1 U9439 ( .B1(n10177), .B2(n7881), .A(n7873), .ZN(n7874) );
  OAI211_X1 U9440 ( .C1(n7876), .C2(n10197), .A(n7875), .B(n7874), .ZN(n7879)
         );
  NAND2_X1 U9441 ( .A1(n7879), .A2(n10217), .ZN(n7877) );
  OAI21_X1 U9442 ( .B1(n10217), .B2(n7878), .A(n7877), .ZN(P1_U3484) );
  NAND2_X1 U9443 ( .A1(n7879), .A2(n10231), .ZN(n7880) );
  OAI21_X1 U9444 ( .B1(n10231), .B2(n6132), .A(n7880), .ZN(P1_U3533) );
  OR2_X1 U9445 ( .A1(n7881), .A2(n9015), .ZN(n7882) );
  XNOR2_X1 U9446 ( .A(n7985), .B(n7884), .ZN(n9947) );
  INV_X1 U9447 ( .A(n7885), .ZN(n7887) );
  XNOR2_X1 U9448 ( .A(n7992), .B(n7889), .ZN(n7893) );
  OAI22_X1 U9449 ( .A1(n7890), .A2(n9236), .B1(n8082), .B2(n9238), .ZN(n7891)
         );
  INV_X1 U9450 ( .A(n7891), .ZN(n7892) );
  OAI21_X1 U9451 ( .B1(n7893), .B2(n9356), .A(n7892), .ZN(n7894) );
  AOI21_X1 U9452 ( .B1(n9947), .B2(n8040), .A(n7894), .ZN(n9949) );
  INV_X1 U9453 ( .A(n10143), .ZN(n9242) );
  INV_X1 U9454 ( .A(n7986), .ZN(n9944) );
  NOR2_X1 U9455 ( .A1(n7895), .A2(n9944), .ZN(n7896) );
  OR2_X1 U9456 ( .A1(n8002), .A2(n7896), .ZN(n9945) );
  OAI22_X1 U9457 ( .A1(n10143), .A2(n7897), .B1(n7940), .B2(n10151), .ZN(n7898) );
  AOI21_X1 U9458 ( .B1(n7986), .B2(n9343), .A(n7898), .ZN(n7899) );
  OAI21_X1 U9459 ( .B1(n9945), .B2(n10146), .A(n7899), .ZN(n7900) );
  AOI21_X1 U9460 ( .B1(n9947), .B2(n10140), .A(n7900), .ZN(n7901) );
  OAI21_X1 U9461 ( .B1(n9949), .B2(n9242), .A(n7901), .ZN(P1_U3280) );
  XNOR2_X1 U9462 ( .A(n8009), .B(n8156), .ZN(n7905) );
  INV_X1 U9463 ( .A(n7905), .ZN(n7903) );
  OR2_X1 U9464 ( .A1(n8008), .A2(n8243), .ZN(n7904) );
  INV_X1 U9465 ( .A(n7904), .ZN(n7902) );
  NAND2_X1 U9466 ( .A1(n7903), .A2(n7902), .ZN(n7960) );
  NAND2_X1 U9467 ( .A1(n7905), .A2(n7904), .ZN(n7958) );
  NAND2_X1 U9468 ( .A1(n7960), .A2(n7958), .ZN(n7912) );
  INV_X1 U9469 ( .A(n7908), .ZN(n7910) );
  NAND2_X1 U9470 ( .A1(n7910), .A2(n7909), .ZN(n7911) );
  XOR2_X1 U9471 ( .A(n7912), .B(n7959), .Z(n7917) );
  INV_X1 U9472 ( .A(n7926), .ZN(n8374) );
  AOI22_X1 U9473 ( .A1(n8374), .A2(n8334), .B1(n7930), .B2(n8344), .ZN(n7914)
         );
  OAI211_X1 U9474 ( .C1(n8370), .C2(n8321), .A(n7914), .B(n7913), .ZN(n7915)
         );
  AOI21_X1 U9475 ( .B1(n8009), .B2(n8324), .A(n7915), .ZN(n7916) );
  OAI21_X1 U9476 ( .B1(n7917), .B2(n8340), .A(n7916), .ZN(P2_U3226) );
  OAI222_X1 U9477 ( .A1(P1_U3084), .A2(n7919), .B1(n8155), .B2(n9779), .C1(
        n9492), .C2(n7918), .ZN(P1_U3329) );
  NAND2_X1 U9478 ( .A1(n7921), .A2(n7920), .ZN(n7923) );
  NAND2_X1 U9479 ( .A1(n8840), .A2(n8374), .ZN(n7922) );
  NAND2_X1 U9480 ( .A1(n7923), .A2(n7922), .ZN(n8011) );
  XNOR2_X1 U9481 ( .A(n8011), .B(n8010), .ZN(n10341) );
  INV_X1 U9482 ( .A(n10341), .ZN(n7935) );
  XNOR2_X1 U9483 ( .A(n7924), .B(n8010), .ZN(n7925) );
  OAI222_X1 U9484 ( .A1(n8639), .A2(n8370), .B1(n8637), .B2(n7926), .C1(n8715), 
        .C2(n7925), .ZN(n10338) );
  INV_X1 U9485 ( .A(n7927), .ZN(n7929) );
  INV_X1 U9486 ( .A(n8021), .ZN(n7928) );
  OAI21_X1 U9487 ( .B1(n4729), .B2(n7929), .A(n7928), .ZN(n10337) );
  AOI22_X1 U9488 ( .A1(n10266), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n7930), .B2(
        n10257), .ZN(n7932) );
  NAND2_X1 U9489 ( .A1(n8009), .A2(n8486), .ZN(n7931) );
  OAI211_X1 U9490 ( .C1(n10337), .C2(n8550), .A(n7932), .B(n7931), .ZN(n7933)
         );
  AOI21_X1 U9491 ( .B1(n10338), .B2(n10263), .A(n7933), .ZN(n7934) );
  OAI21_X1 U9492 ( .B1(n8742), .B2(n7935), .A(n7934), .ZN(P2_U3284) );
  AOI21_X1 U9493 ( .B1(n7937), .B2(n7936), .A(n9009), .ZN(n7939) );
  NAND2_X1 U9494 ( .A1(n7939), .A2(n7938), .ZN(n7944) );
  NAND2_X1 U9495 ( .A1(P1_U3084), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n10024) );
  OAI21_X1 U9496 ( .B1(n8981), .B2(n8082), .A(n10024), .ZN(n7942) );
  NOR2_X1 U9497 ( .A1(n9005), .A2(n7940), .ZN(n7941) );
  AOI211_X1 U9498 ( .C1(n8983), .C2(n9015), .A(n7942), .B(n7941), .ZN(n7943)
         );
  OAI211_X1 U9499 ( .C1(n9944), .C2(n8996), .A(n7944), .B(n7943), .ZN(P1_U3234) );
  INV_X1 U9500 ( .A(n7945), .ZN(n7951) );
  INV_X1 U9501 ( .A(n7946), .ZN(n7947) );
  OAI222_X1 U9502 ( .A1(n8876), .A2(n7949), .B1(n8871), .B2(n7951), .C1(
        P2_U3152), .C2(n7947), .ZN(P2_U3333) );
  OAI222_X1 U9503 ( .A1(n7952), .A2(P1_U3084), .B1(n9492), .B2(n7951), .C1(
        n7950), .C2(n8155), .ZN(P1_U3328) );
  XNOR2_X1 U9504 ( .A(n8024), .B(n7953), .ZN(n7954) );
  NOR2_X1 U9505 ( .A1(n8370), .A2(n8243), .ZN(n7955) );
  NAND2_X1 U9506 ( .A1(n7954), .A2(n7955), .ZN(n8095) );
  INV_X1 U9507 ( .A(n7954), .ZN(n8089) );
  INV_X1 U9508 ( .A(n7955), .ZN(n7956) );
  NAND2_X1 U9509 ( .A1(n8089), .A2(n7956), .ZN(n7957) );
  AND2_X1 U9510 ( .A1(n8095), .A2(n7957), .ZN(n7963) );
  NAND2_X1 U9511 ( .A1(n7961), .A2(n7960), .ZN(n7962) );
  OAI211_X1 U9512 ( .C1(n7963), .C2(n7962), .A(n8097), .B(n8353), .ZN(n7970)
         );
  OR2_X1 U9513 ( .A1(n8008), .A2(n8637), .ZN(n7965) );
  OR2_X1 U9514 ( .A1(n8110), .A2(n8639), .ZN(n7964) );
  NAND2_X1 U9515 ( .A1(n7965), .A2(n7964), .ZN(n8016) );
  INV_X1 U9516 ( .A(n8023), .ZN(n7967) );
  OAI21_X1 U9517 ( .B1(n8360), .B2(n7967), .A(n7966), .ZN(n7968) );
  AOI21_X1 U9518 ( .B1(n8016), .B2(n8362), .A(n7968), .ZN(n7969) );
  OAI211_X1 U9519 ( .C1(n8832), .C2(n8366), .A(n7970), .B(n7969), .ZN(P2_U3236) );
  OAI21_X1 U9520 ( .B1(n7972), .B2(P2_REG2_REG_14__SCAN_IN), .A(n7971), .ZN(
        n8423) );
  XNOR2_X1 U9521 ( .A(n8423), .B(n8416), .ZN(n7974) );
  INV_X1 U9522 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n7973) );
  NAND2_X1 U9523 ( .A1(n7974), .A2(n7973), .ZN(n8425) );
  OAI21_X1 U9524 ( .B1(n7974), .B2(n7973), .A(n8425), .ZN(n7982) );
  AOI21_X1 U9525 ( .B1(n7976), .B2(n9915), .A(n7975), .ZN(n8415) );
  XNOR2_X1 U9526 ( .A(n8415), .B(n8424), .ZN(n7977) );
  NAND2_X1 U9527 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n7977), .ZN(n8417) );
  OAI211_X1 U9528 ( .C1(n7977), .C2(P2_REG1_REG_15__SCAN_IN), .A(n10232), .B(
        n8417), .ZN(n7980) );
  NOR2_X1 U9529 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8358), .ZN(n7978) );
  AOI21_X1 U9530 ( .B1(n10234), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n7978), .ZN(
        n7979) );
  OAI211_X1 U9531 ( .C1(n10235), .C2(n8424), .A(n7980), .B(n7979), .ZN(n7981)
         );
  AOI21_X1 U9532 ( .B1(n10233), .B2(n7982), .A(n7981), .ZN(n7983) );
  INV_X1 U9533 ( .A(n7983), .ZN(P2_U3260) );
  NAND2_X1 U9534 ( .A1(n7986), .A2(n9014), .ZN(n7984) );
  INV_X1 U9535 ( .A(n7989), .ZN(n7988) );
  NAND2_X1 U9536 ( .A1(n7989), .A2(n7994), .ZN(n7990) );
  NAND2_X1 U9537 ( .A1(n8031), .A2(n7990), .ZN(n8001) );
  OR2_X1 U9538 ( .A1(n8001), .A2(n10130), .ZN(n8000) );
  NAND2_X1 U9539 ( .A1(n8033), .A2(n7993), .ZN(n7995) );
  XNOR2_X1 U9540 ( .A(n7995), .B(n7987), .ZN(n7998) );
  NAND2_X1 U9541 ( .A1(n9070), .A2(n9370), .ZN(n7997) );
  NAND2_X1 U9542 ( .A1(n9014), .A2(n9368), .ZN(n7996) );
  NAND2_X1 U9543 ( .A1(n7997), .A2(n7996), .ZN(n8071) );
  AOI21_X1 U9544 ( .B1(n7998), .B2(n10133), .A(n8071), .ZN(n7999) );
  INV_X1 U9545 ( .A(n8001), .ZN(n9941) );
  INV_X1 U9546 ( .A(n8075), .ZN(n9939) );
  OAI211_X1 U9547 ( .C1(n8002), .C2(n9939), .A(n10125), .B(n8041), .ZN(n9938)
         );
  OAI22_X1 U9548 ( .A1(n10143), .A2(n8003), .B1(n8073), .B2(n10151), .ZN(n8004) );
  AOI21_X1 U9549 ( .B1(n8075), .B2(n9343), .A(n8004), .ZN(n8005) );
  OAI21_X1 U9550 ( .B1(n9938), .B2(n9325), .A(n8005), .ZN(n8006) );
  AOI21_X1 U9551 ( .B1(n9941), .B2(n10140), .A(n8006), .ZN(n8007) );
  OAI21_X1 U9552 ( .B1(n9943), .B2(n9242), .A(n8007), .ZN(P1_U3279) );
  INV_X1 U9553 ( .A(n8008), .ZN(n8373) );
  NAND2_X1 U9554 ( .A1(n8012), .A2(n8015), .ZN(n8013) );
  NAND2_X1 U9555 ( .A1(n8048), .A2(n8013), .ZN(n8020) );
  OR2_X1 U9556 ( .A1(n8020), .A2(n10298), .ZN(n8019) );
  OAI21_X1 U9557 ( .B1(n8015), .B2(n8014), .A(n8050), .ZN(n8017) );
  AOI21_X1 U9558 ( .B1(n8017), .B2(n10254), .A(n8016), .ZN(n8018) );
  INV_X1 U9559 ( .A(n8020), .ZN(n8835) );
  NOR2_X1 U9560 ( .A1(n8021), .A2(n8832), .ZN(n8022) );
  OR2_X1 U9561 ( .A1(n8054), .A2(n8022), .ZN(n8833) );
  AOI22_X1 U9562 ( .A1(n10266), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n8023), .B2(
        n10257), .ZN(n8026) );
  NAND2_X1 U9563 ( .A1(n8024), .A2(n8486), .ZN(n8025) );
  OAI211_X1 U9564 ( .C1(n8833), .C2(n8550), .A(n8026), .B(n8025), .ZN(n8027)
         );
  AOI21_X1 U9565 ( .B1(n8835), .B2(n8028), .A(n8027), .ZN(n8029) );
  OAI21_X1 U9566 ( .B1(n8837), .B2(n10266), .A(n8029), .ZN(P2_U3283) );
  INV_X1 U9567 ( .A(n8082), .ZN(n9013) );
  NAND2_X1 U9568 ( .A1(n8075), .A2(n9013), .ZN(n8030) );
  XNOR2_X1 U9569 ( .A(n9069), .B(n9101), .ZN(n9935) );
  NAND2_X1 U9570 ( .A1(n8033), .A2(n8032), .ZN(n8035) );
  NAND2_X1 U9571 ( .A1(n8035), .A2(n8034), .ZN(n9102) );
  XNOR2_X1 U9572 ( .A(n9102), .B(n8036), .ZN(n8038) );
  AOI22_X1 U9573 ( .A1(n9013), .A2(n9368), .B1(n9370), .B2(n9073), .ZN(n8037)
         );
  OAI21_X1 U9574 ( .B1(n8038), .B2(n9356), .A(n8037), .ZN(n8039) );
  AOI21_X1 U9575 ( .B1(n9935), .B2(n8040), .A(n8039), .ZN(n9937) );
  NAND2_X1 U9576 ( .A1(n8041), .A2(n9932), .ZN(n8042) );
  NAND2_X1 U9577 ( .A1(n9350), .A2(n8042), .ZN(n9933) );
  OAI22_X1 U9578 ( .A1(n10143), .A2(n8043), .B1(n8085), .B2(n10151), .ZN(n8044) );
  AOI21_X1 U9579 ( .B1(n9932), .B2(n9343), .A(n8044), .ZN(n8045) );
  OAI21_X1 U9580 ( .B1(n9933), .B2(n10146), .A(n8045), .ZN(n8046) );
  AOI21_X1 U9581 ( .B1(n9935), .B2(n10140), .A(n8046), .ZN(n8047) );
  OAI21_X1 U9582 ( .B1(n9937), .B2(n9242), .A(n8047), .ZN(P1_U3278) );
  XNOR2_X1 U9583 ( .A(n8113), .B(n8112), .ZN(n9914) );
  INV_X1 U9584 ( .A(n9914), .ZN(n8059) );
  NAND2_X1 U9585 ( .A1(n8050), .A2(n8049), .ZN(n8052) );
  XNOR2_X1 U9586 ( .A(n8052), .B(n8051), .ZN(n8053) );
  OAI222_X1 U9587 ( .A1(n8639), .A2(n8281), .B1(n8637), .B2(n8370), .C1(n8053), 
        .C2(n8715), .ZN(n9912) );
  INV_X1 U9588 ( .A(n8111), .ZN(n9911) );
  OAI211_X1 U9589 ( .C1(n8054), .C2(n9911), .A(n10246), .B(n8117), .ZN(n9910)
         );
  AOI22_X1 U9590 ( .A1(n10266), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n8092), .B2(
        n10257), .ZN(n8056) );
  NAND2_X1 U9591 ( .A1(n8111), .A2(n8486), .ZN(n8055) );
  OAI211_X1 U9592 ( .C1(n9910), .C2(n8561), .A(n8056), .B(n8055), .ZN(n8057)
         );
  AOI21_X1 U9593 ( .B1(n9912), .B2(n10263), .A(n8057), .ZN(n8058) );
  OAI21_X1 U9594 ( .B1(n8059), .B2(n8742), .A(n8058), .ZN(P2_U3282) );
  INV_X1 U9595 ( .A(n8060), .ZN(n8063) );
  OAI222_X1 U9596 ( .A1(n8876), .A2(n8062), .B1(n8871), .B2(n8063), .C1(
        P2_U3152), .C2(n8061), .ZN(P2_U3332) );
  OAI222_X1 U9597 ( .A1(n8065), .A2(P1_U3084), .B1(n9492), .B2(n8063), .C1(
        n9681), .C2(n9489), .ZN(P1_U3327) );
  INV_X1 U9598 ( .A(n8066), .ZN(n8067) );
  AOI21_X1 U9599 ( .B1(n8069), .B2(n8068), .A(n8067), .ZN(n8077) );
  NOR2_X1 U9600 ( .A1(n8070), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10037) );
  AOI21_X1 U9601 ( .B1(n9003), .B2(n8071), .A(n10037), .ZN(n8072) );
  OAI21_X1 U9602 ( .B1(n9005), .B2(n8073), .A(n8072), .ZN(n8074) );
  AOI21_X1 U9603 ( .B1(n8075), .B2(n9007), .A(n8074), .ZN(n8076) );
  OAI21_X1 U9604 ( .B1(n8077), .B2(n9009), .A(n8076), .ZN(P1_U3222) );
  XNOR2_X1 U9605 ( .A(n8080), .B(n8079), .ZN(n8081) );
  XNOR2_X1 U9606 ( .A(n8078), .B(n8081), .ZN(n8088) );
  NAND2_X1 U9607 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n10052) );
  OAI21_X1 U9608 ( .B1(n8960), .B2(n8082), .A(n10052), .ZN(n8083) );
  AOI21_X1 U9609 ( .B1(n8971), .B2(n9073), .A(n8083), .ZN(n8084) );
  OAI21_X1 U9610 ( .B1(n9005), .B2(n8085), .A(n8084), .ZN(n8086) );
  AOI21_X1 U9611 ( .B1(n9932), .B2(n9007), .A(n8086), .ZN(n8087) );
  OAI21_X1 U9612 ( .B1(n8088), .B2(n9009), .A(n8087), .ZN(P1_U3232) );
  INV_X1 U9613 ( .A(n8097), .ZN(n8091) );
  NOR3_X1 U9614 ( .A1(n8089), .A2(n8370), .A3(n8301), .ZN(n8090) );
  AOI21_X1 U9615 ( .B1(n8091), .B2(n8353), .A(n8090), .ZN(n8102) );
  XNOR2_X1 U9616 ( .A(n8111), .B(n8156), .ZN(n8159) );
  NOR2_X1 U9617 ( .A1(n8110), .A2(n8243), .ZN(n8157) );
  XNOR2_X1 U9618 ( .A(n8159), .B(n8157), .ZN(n8101) );
  AOI22_X1 U9619 ( .A1(n8494), .A2(n8349), .B1(n8344), .B2(n8092), .ZN(n8094)
         );
  OAI211_X1 U9620 ( .C1(n8370), .C2(n8347), .A(n8094), .B(n8093), .ZN(n8099)
         );
  AND2_X1 U9621 ( .A1(n8101), .A2(n8095), .ZN(n8096) );
  NOR2_X1 U9622 ( .A1(n8160), .A2(n8340), .ZN(n8098) );
  AOI211_X1 U9623 ( .C1(n8111), .C2(n8324), .A(n8099), .B(n8098), .ZN(n8100)
         );
  OAI21_X1 U9624 ( .B1(n8102), .B2(n8101), .A(n8100), .ZN(P2_U3217) );
  NAND2_X1 U9625 ( .A1(n6312), .A2(n8103), .ZN(n8105) );
  OAI211_X1 U9626 ( .C1(n8155), .C2(n9863), .A(n8105), .B(n8104), .ZN(P1_U3326) );
  XNOR2_X1 U9627 ( .A(n8106), .B(n8114), .ZN(n8109) );
  OR2_X1 U9628 ( .A1(n8289), .A2(n8639), .ZN(n8108) );
  OR2_X1 U9629 ( .A1(n8110), .A2(n8637), .ZN(n8107) );
  NAND2_X1 U9630 ( .A1(n8108), .A2(n8107), .ZN(n8363) );
  AOI21_X1 U9631 ( .B1(n8109), .B2(n10254), .A(n8363), .ZN(n8825) );
  INV_X1 U9632 ( .A(n8110), .ZN(n8369) );
  OAI21_X1 U9633 ( .B1(n8115), .B2(n8114), .A(n8497), .ZN(n8828) );
  NAND2_X1 U9634 ( .A1(n8828), .A2(n8615), .ZN(n8121) );
  INV_X1 U9635 ( .A(n8116), .ZN(n8359) );
  OAI22_X1 U9636 ( .A1(n10263), .A2(n7973), .B1(n8359), .B2(n8620), .ZN(n8119)
         );
  OAI211_X1 U9637 ( .C1(n4725), .C2(n8826), .A(n10246), .B(n4488), .ZN(n8824)
         );
  NOR2_X1 U9638 ( .A1(n8824), .A2(n8561), .ZN(n8118) );
  AOI211_X1 U9639 ( .C1(n8486), .C2(n8495), .A(n8119), .B(n8118), .ZN(n8120)
         );
  OAI211_X1 U9640 ( .C1(n10266), .C2(n8825), .A(n8121), .B(n8120), .ZN(
        P2_U3281) );
  XNOR2_X1 U9641 ( .A(n8123), .B(n8122), .ZN(n8124) );
  XNOR2_X1 U9642 ( .A(n8125), .B(n8124), .ZN(n8131) );
  NAND2_X1 U9643 ( .A1(P1_U3084), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n10062) );
  OR2_X1 U9644 ( .A1(n8932), .A2(n9238), .ZN(n8127) );
  NAND2_X1 U9645 ( .A1(n9070), .A2(n9368), .ZN(n8126) );
  NAND2_X1 U9646 ( .A1(n8127), .A2(n8126), .ZN(n9359) );
  NAND2_X1 U9647 ( .A1(n9359), .A2(n9003), .ZN(n8128) );
  OAI211_X1 U9648 ( .C1(n9005), .C2(n9351), .A(n10062), .B(n8128), .ZN(n8129)
         );
  AOI21_X1 U9649 ( .B1(n9463), .B2(n9007), .A(n8129), .ZN(n8130) );
  OAI21_X1 U9650 ( .B1(n8131), .B2(n9009), .A(n8130), .ZN(P1_U3213) );
  NAND2_X1 U9651 ( .A1(n8150), .A2(n8132), .ZN(n8134) );
  OAI211_X1 U9652 ( .C1(n8876), .C2(n8135), .A(n8134), .B(n8133), .ZN(P2_U3330) );
  INV_X1 U9653 ( .A(n8136), .ZN(n8154) );
  INV_X1 U9654 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8137) );
  OAI222_X1 U9655 ( .A1(P2_U3152), .A2(n5109), .B1(n8871), .B2(n8154), .C1(
        n8137), .C2(n8865), .ZN(P2_U3328) );
  INV_X1 U9656 ( .A(n6312), .ZN(n8138) );
  OAI222_X1 U9657 ( .A1(n8876), .A2(n8139), .B1(n8874), .B2(n8138), .C1(n8484), 
        .C2(P2_U3152), .ZN(P2_U3331) );
  XNOR2_X1 U9658 ( .A(n8141), .B(n8140), .ZN(n8142) );
  XNOR2_X1 U9659 ( .A(n8143), .B(n8142), .ZN(n8144) );
  NAND2_X1 U9660 ( .A1(n8144), .A2(n8956), .ZN(n8149) );
  NAND2_X1 U9661 ( .A1(n9021), .A2(n9370), .ZN(n8146) );
  NAND2_X1 U9662 ( .A1(n6027), .A2(n9368), .ZN(n8145) );
  NAND2_X1 U9663 ( .A1(n8146), .A2(n8145), .ZN(n10132) );
  AOI22_X1 U9664 ( .A1(n9003), .A2(n10132), .B1(P1_REG3_REG_1__SCAN_IN), .B2(
        n8147), .ZN(n8148) );
  OAI211_X1 U9665 ( .C1(n10160), .C2(n8996), .A(n8149), .B(n8148), .ZN(
        P1_U3220) );
  INV_X1 U9666 ( .A(n8150), .ZN(n8152) );
  OAI222_X1 U9667 ( .A1(n9492), .A2(n8152), .B1(P1_U3084), .B2(n8151), .C1(
        n9866), .C2(n9489), .ZN(P1_U3325) );
  OAI222_X1 U9668 ( .A1(n8155), .A2(n9807), .B1(n9487), .B2(n8154), .C1(n8153), 
        .C2(P1_U3084), .ZN(P1_U3323) );
  NAND2_X1 U9669 ( .A1(n8506), .A2(n8168), .ZN(n8190) );
  INV_X1 U9670 ( .A(n8190), .ZN(n8192) );
  XNOR2_X1 U9671 ( .A(n8773), .B(n7953), .ZN(n8191) );
  NAND2_X1 U9672 ( .A1(n8505), .A2(n8168), .ZN(n8212) );
  XNOR2_X1 U9673 ( .A(n8794), .B(n7953), .ZN(n8179) );
  INV_X1 U9674 ( .A(n8179), .ZN(n8182) );
  NAND2_X1 U9675 ( .A1(n8670), .A2(n8168), .ZN(n8181) );
  NOR2_X1 U9676 ( .A1(n8502), .A2(n8243), .ZN(n8176) );
  XNOR2_X1 U9677 ( .A(n8682), .B(n7953), .ZN(n8174) );
  XNOR2_X1 U9678 ( .A(n8495), .B(n7953), .ZN(n8274) );
  INV_X1 U9679 ( .A(n8274), .ZN(n8276) );
  NOR2_X1 U9680 ( .A1(n8281), .A2(n8243), .ZN(n8161) );
  INV_X1 U9681 ( .A(n8161), .ZN(n8354) );
  NOR2_X1 U9682 ( .A1(n8289), .A2(n8243), .ZN(n8162) );
  INV_X1 U9683 ( .A(n8162), .ZN(n8277) );
  AOI21_X1 U9684 ( .B1(n8276), .B2(n8354), .A(n8277), .ZN(n8165) );
  XNOR2_X1 U9685 ( .A(n8820), .B(n7953), .ZN(n8278) );
  INV_X1 U9686 ( .A(n8157), .ZN(n8158) );
  AOI22_X1 U9687 ( .A1(n8278), .A2(n8162), .B1(n8161), .B2(n8274), .ZN(n8163)
         );
  NAND3_X1 U9688 ( .A1(n8276), .A2(n8354), .A3(n8277), .ZN(n8164) );
  XNOR2_X1 U9689 ( .A(n8816), .B(n7953), .ZN(n8327) );
  AND2_X1 U9690 ( .A1(n8701), .A2(n8168), .ZN(n8166) );
  NAND2_X1 U9691 ( .A1(n8327), .A2(n8166), .ZN(n8167) );
  OAI21_X1 U9692 ( .B1(n8327), .B2(n8166), .A(n8167), .ZN(n8292) );
  INV_X1 U9693 ( .A(n8167), .ZN(n8173) );
  XNOR2_X1 U9694 ( .A(n8809), .B(n7953), .ZN(n8169) );
  AND2_X1 U9695 ( .A1(n8685), .A2(n8168), .ZN(n8170) );
  NAND2_X1 U9696 ( .A1(n8169), .A2(n8170), .ZN(n8175) );
  INV_X1 U9697 ( .A(n8169), .ZN(n8232) );
  INV_X1 U9698 ( .A(n8170), .ZN(n8171) );
  NAND2_X1 U9699 ( .A1(n8232), .A2(n8171), .ZN(n8172) );
  AND2_X1 U9700 ( .A1(n8175), .A2(n8172), .ZN(n8328) );
  XNOR2_X1 U9701 ( .A(n8174), .B(n8176), .ZN(n8233) );
  XNOR2_X1 U9702 ( .A(n8799), .B(n7953), .ZN(n8255) );
  NOR2_X1 U9703 ( .A1(n8503), .A2(n8243), .ZN(n8177) );
  NAND2_X1 U9704 ( .A1(n8255), .A2(n8177), .ZN(n8178) );
  OAI21_X1 U9705 ( .B1(n8255), .B2(n8177), .A(n8178), .ZN(n8312) );
  INV_X1 U9706 ( .A(n8178), .ZN(n8180) );
  XNOR2_X1 U9707 ( .A(n8179), .B(n8181), .ZN(n8254) );
  NOR2_X1 U9708 ( .A1(n8261), .A2(n8243), .ZN(n8317) );
  XNOR2_X1 U9709 ( .A(n8618), .B(n7953), .ZN(n8184) );
  NOR2_X1 U9710 ( .A1(n8368), .A2(n8243), .ZN(n8187) );
  INV_X1 U9711 ( .A(n8187), .ZN(n8303) );
  INV_X1 U9712 ( .A(n8299), .ZN(n8186) );
  NOR2_X1 U9713 ( .A1(n8185), .A2(n8184), .ZN(n8297) );
  OAI21_X1 U9714 ( .B1(n8187), .B2(n8186), .A(n8297), .ZN(n8188) );
  OAI21_X1 U9715 ( .B1(n8299), .B2(n8303), .A(n8188), .ZN(n8189) );
  XNOR2_X1 U9716 ( .A(n8191), .B(n8190), .ZN(n8267) );
  XNOR2_X1 U9717 ( .A(n8768), .B(n7953), .ZN(n8200) );
  NOR2_X1 U9718 ( .A1(n8508), .A2(n8243), .ZN(n8193) );
  NAND2_X1 U9719 ( .A1(n8200), .A2(n8193), .ZN(n8203) );
  OAI21_X1 U9720 ( .B1(n8200), .B2(n8193), .A(n8203), .ZN(n8342) );
  XNOR2_X1 U9721 ( .A(n8194), .B(n7953), .ZN(n8195) );
  NOR2_X1 U9722 ( .A1(n8573), .A2(n8243), .ZN(n8196) );
  NAND2_X1 U9723 ( .A1(n8195), .A2(n8196), .ZN(n8241) );
  INV_X1 U9724 ( .A(n8195), .ZN(n8198) );
  INV_X1 U9725 ( .A(n8196), .ZN(n8197) );
  NAND2_X1 U9726 ( .A1(n8198), .A2(n8197), .ZN(n8199) );
  NOR2_X1 U9727 ( .A1(n8339), .A2(n8204), .ZN(n8202) );
  INV_X1 U9728 ( .A(n8508), .ZN(n8545) );
  NAND3_X1 U9729 ( .A1(n8200), .A2(n8352), .A3(n8545), .ZN(n8201) );
  OAI21_X1 U9730 ( .B1(n8202), .B2(n8340), .A(n8201), .ZN(n8205) );
  NAND2_X1 U9731 ( .A1(n8205), .A2(n8242), .ZN(n8210) );
  OAI22_X1 U9732 ( .A1(n8508), .A2(n8347), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8206), .ZN(n8208) );
  NOR2_X1 U9733 ( .A1(n8548), .A2(n8321), .ZN(n8207) );
  AOI211_X1 U9734 ( .C1(n8344), .C2(n8551), .A(n8208), .B(n8207), .ZN(n8209)
         );
  OAI211_X1 U9735 ( .C1(n8760), .C2(n8366), .A(n8210), .B(n8209), .ZN(P2_U3216) );
  INV_X1 U9736 ( .A(n8213), .ZN(n8211) );
  AOI22_X1 U9737 ( .A1(n8211), .A2(n8353), .B1(n8352), .B2(n8505), .ZN(n8218)
         );
  NOR2_X1 U9738 ( .A1(n8213), .A2(n8212), .ZN(n8298) );
  OAI22_X1 U9739 ( .A1(n8261), .A2(n8347), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8214), .ZN(n8216) );
  OAI22_X1 U9740 ( .A1(n8368), .A2(n8321), .B1(n8360), .B2(n8621), .ZN(n8215)
         );
  AOI211_X1 U9741 ( .C1(n8784), .C2(n8324), .A(n8216), .B(n8215), .ZN(n8217)
         );
  OAI21_X1 U9742 ( .B1(n8218), .B2(n8298), .A(n8217), .ZN(P2_U3218) );
  INV_X1 U9743 ( .A(n8219), .ZN(n8220) );
  AOI21_X1 U9744 ( .B1(n8221), .B2(n8220), .A(n8340), .ZN(n8225) );
  NOR3_X1 U9745 ( .A1(n8223), .A2(n8222), .A3(n8301), .ZN(n8224) );
  OAI21_X1 U9746 ( .B1(n8225), .B2(n8224), .A(n7148), .ZN(n8230) );
  AOI22_X1 U9747 ( .A1(n8227), .A2(n8362), .B1(n8226), .B2(n8324), .ZN(n8229)
         );
  MUX2_X1 U9748 ( .A(P2_STATE_REG_SCAN_IN), .B(n8360), .S(n9820), .Z(n8228) );
  NAND3_X1 U9749 ( .A1(n8230), .A2(n8229), .A3(n8228), .ZN(P2_U3220) );
  OAI21_X1 U9750 ( .B1(n8233), .B2(n8330), .A(n8231), .ZN(n8239) );
  NOR3_X1 U9751 ( .A1(n8233), .A2(n8232), .A3(n8301), .ZN(n8234) );
  OAI21_X1 U9752 ( .B1(n8234), .B2(n8334), .A(n8685), .ZN(n8237) );
  NAND2_X1 U9753 ( .A1(P2_U3152), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8479) );
  OAI21_X1 U9754 ( .B1(n8503), .B2(n8321), .A(n8479), .ZN(n8235) );
  AOI21_X1 U9755 ( .B1(n8680), .B2(n8344), .A(n8235), .ZN(n8236) );
  OAI211_X1 U9756 ( .C1(n8682), .C2(n8366), .A(n8237), .B(n8236), .ZN(n8238)
         );
  AOI21_X1 U9757 ( .B1(n8239), .B2(n8353), .A(n8238), .ZN(n8240) );
  INV_X1 U9758 ( .A(n8240), .ZN(P2_U3221) );
  NOR2_X1 U9759 ( .A1(n8548), .A2(n8243), .ZN(n8244) );
  XOR2_X1 U9760 ( .A(n7953), .B(n8244), .Z(n8245) );
  XNOR2_X1 U9761 ( .A(n8755), .B(n8245), .ZN(n8246) );
  XNOR2_X1 U9762 ( .A(n8247), .B(n8246), .ZN(n8253) );
  INV_X1 U9763 ( .A(n8248), .ZN(n8528) );
  NAND2_X1 U9764 ( .A1(n8528), .A2(n8349), .ZN(n8250) );
  AOI22_X1 U9765 ( .A1(n8533), .A2(n8344), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3152), .ZN(n8249) );
  OAI211_X1 U9766 ( .C1(n8573), .C2(n8347), .A(n8250), .B(n8249), .ZN(n8251)
         );
  AOI21_X1 U9767 ( .B1(n8755), .B2(n8324), .A(n8251), .ZN(n8252) );
  OAI21_X1 U9768 ( .B1(n8253), .B2(n8340), .A(n8252), .ZN(P2_U3222) );
  OAI21_X1 U9769 ( .B1(n8310), .B2(n8254), .A(n8353), .ZN(n8257) );
  INV_X1 U9770 ( .A(n8503), .ZN(n8686) );
  NAND3_X1 U9771 ( .A1(n8255), .A2(n8352), .A3(n8686), .ZN(n8256) );
  NAND2_X1 U9772 ( .A1(n8257), .A2(n8256), .ZN(n8259) );
  NAND2_X1 U9773 ( .A1(n8259), .A2(n8258), .ZN(n8265) );
  NOR2_X1 U9774 ( .A1(n8503), .A2(n8347), .ZN(n8263) );
  OAI22_X1 U9775 ( .A1(n8261), .A2(n8321), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8260), .ZN(n8262) );
  AOI211_X1 U9776 ( .C1(n8344), .C2(n8650), .A(n8263), .B(n8262), .ZN(n8264)
         );
  OAI211_X1 U9777 ( .C1(n8652), .C2(n8366), .A(n8265), .B(n8264), .ZN(P2_U3225) );
  INV_X1 U9778 ( .A(n8773), .ZN(n8585) );
  OAI21_X1 U9779 ( .B1(n8268), .B2(n8267), .A(n8266), .ZN(n8269) );
  NAND2_X1 U9780 ( .A1(n8269), .A2(n8353), .ZN(n8273) );
  OAI22_X1 U9781 ( .A1(n8508), .A2(n8639), .B1(n8368), .B2(n8637), .ZN(n8577)
         );
  OAI22_X1 U9782 ( .A1(n8587), .A2(n8360), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8270), .ZN(n8271) );
  AOI21_X1 U9783 ( .B1(n8577), .B2(n8362), .A(n8271), .ZN(n8272) );
  OAI211_X1 U9784 ( .C1(n8585), .C2(n8366), .A(n8273), .B(n8272), .ZN(P2_U3227) );
  XNOR2_X1 U9785 ( .A(n8275), .B(n8274), .ZN(n8355) );
  AOI22_X1 U9786 ( .A1(n8355), .A2(n8354), .B1(n8276), .B2(n8275), .ZN(n8280)
         );
  XNOR2_X1 U9787 ( .A(n8278), .B(n8277), .ZN(n8279) );
  XNOR2_X1 U9788 ( .A(n8280), .B(n8279), .ZN(n8288) );
  OR2_X1 U9789 ( .A1(n8281), .A2(n8637), .ZN(n8283) );
  NAND2_X1 U9790 ( .A1(n8701), .A2(n8702), .ZN(n8282) );
  NAND2_X1 U9791 ( .A1(n8283), .A2(n8282), .ZN(n8737) );
  INV_X1 U9792 ( .A(n8731), .ZN(n8284) );
  OAI22_X1 U9793 ( .A1(n8360), .A2(n8284), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9860), .ZN(n8285) );
  AOI21_X1 U9794 ( .B1(n8737), .B2(n8362), .A(n8285), .ZN(n8287) );
  NAND2_X1 U9795 ( .A1(n8820), .A2(n8324), .ZN(n8286) );
  OAI211_X1 U9796 ( .C1(n8288), .C2(n8340), .A(n8287), .B(n8286), .ZN(P2_U3228) );
  INV_X1 U9797 ( .A(n8289), .ZN(n8498) );
  AOI22_X1 U9798 ( .A1(n8498), .A2(n8700), .B1(n8702), .B2(n8685), .ZN(n8714)
         );
  AOI22_X1 U9799 ( .A1(n8344), .A2(n8720), .B1(P2_REG3_REG_17__SCAN_IN), .B2(
        P2_U3152), .ZN(n8290) );
  OAI21_X1 U9800 ( .B1(n8714), .B2(n8291), .A(n8290), .ZN(n8295) );
  AOI211_X1 U9801 ( .C1(n8293), .C2(n8292), .A(n8340), .B(n8329), .ZN(n8294)
         );
  AOI211_X1 U9802 ( .C1(n8816), .C2(n8324), .A(n8295), .B(n8294), .ZN(n8296)
         );
  INV_X1 U9803 ( .A(n8296), .ZN(P2_U3230) );
  NOR2_X1 U9804 ( .A1(n8298), .A2(n8297), .ZN(n8300) );
  XNOR2_X1 U9805 ( .A(n8300), .B(n8299), .ZN(n8304) );
  OAI22_X1 U9806 ( .A1(n8304), .A2(n8340), .B1(n8368), .B2(n8301), .ZN(n8302)
         );
  OAI21_X1 U9807 ( .B1(n8304), .B2(n8303), .A(n8302), .ZN(n8309) );
  OAI22_X1 U9808 ( .A1(n8572), .A2(n8639), .B1(n8640), .B2(n8637), .ZN(n8593)
         );
  INV_X1 U9809 ( .A(n8600), .ZN(n8306) );
  OAI22_X1 U9810 ( .A1(n8306), .A2(n8360), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8305), .ZN(n8307) );
  AOI21_X1 U9811 ( .B1(n8593), .B2(n8362), .A(n8307), .ZN(n8308) );
  OAI211_X1 U9812 ( .C1(n4720), .C2(n8366), .A(n8309), .B(n8308), .ZN(P2_U3231) );
  AOI211_X1 U9813 ( .C1(n8312), .C2(n8311), .A(n8340), .B(n8310), .ZN(n8316)
         );
  INV_X1 U9814 ( .A(n8799), .ZN(n8666) );
  AOI22_X1 U9815 ( .A1(n8670), .A2(n8349), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3152), .ZN(n8314) );
  INV_X1 U9816 ( .A(n8502), .ZN(n8703) );
  AOI22_X1 U9817 ( .A1(n8703), .A2(n8334), .B1(n8664), .B2(n8344), .ZN(n8313)
         );
  OAI211_X1 U9818 ( .C1(n8666), .C2(n8366), .A(n8314), .B(n8313), .ZN(n8315)
         );
  OR2_X1 U9819 ( .A1(n8316), .A2(n8315), .ZN(P2_U3235) );
  OR2_X1 U9820 ( .A1(n8317), .A2(n8340), .ZN(n8320) );
  NAND2_X1 U9821 ( .A1(n8656), .A2(n8352), .ZN(n8319) );
  MUX2_X1 U9822 ( .A(n8320), .B(n8319), .S(n8318), .Z(n8326) );
  OAI22_X1 U9823 ( .A1(n8638), .A2(n8347), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9792), .ZN(n8323) );
  OAI22_X1 U9824 ( .A1(n8640), .A2(n8321), .B1(n8360), .B2(n8629), .ZN(n8322)
         );
  AOI211_X1 U9825 ( .C1(n8789), .C2(n8324), .A(n8323), .B(n8322), .ZN(n8325)
         );
  NAND2_X1 U9826 ( .A1(n8326), .A2(n8325), .ZN(P2_U3237) );
  NAND3_X1 U9827 ( .A1(n8327), .A2(n8352), .A3(n8701), .ZN(n8333) );
  OAI21_X1 U9828 ( .B1(n8329), .B2(n8328), .A(n8353), .ZN(n8332) );
  INV_X1 U9829 ( .A(n8330), .ZN(n8331) );
  AOI21_X1 U9830 ( .B1(n8333), .B2(n8332), .A(n8331), .ZN(n8338) );
  AOI22_X1 U9831 ( .A1(n8703), .A2(n8349), .B1(P2_REG3_REG_18__SCAN_IN), .B2(
        P2_U3152), .ZN(n8336) );
  AOI22_X1 U9832 ( .A1(n8334), .A2(n8701), .B1(n8344), .B2(n8695), .ZN(n8335)
         );
  OAI211_X1 U9833 ( .C1(n8697), .C2(n8366), .A(n8336), .B(n8335), .ZN(n8337)
         );
  OR2_X1 U9834 ( .A1(n8338), .A2(n8337), .ZN(P2_U3240) );
  AOI211_X1 U9835 ( .C1(n8342), .C2(n8341), .A(n8340), .B(n8339), .ZN(n8343)
         );
  INV_X1 U9836 ( .A(n8343), .ZN(n8351) );
  INV_X1 U9837 ( .A(n8573), .ZN(n8527) );
  INV_X1 U9838 ( .A(n8564), .ZN(n8345) );
  AOI22_X1 U9839 ( .A1(n8345), .A2(n8344), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3152), .ZN(n8346) );
  OAI21_X1 U9840 ( .B1(n8572), .B2(n8347), .A(n8346), .ZN(n8348) );
  AOI21_X1 U9841 ( .B1(n8527), .B2(n8349), .A(n8348), .ZN(n8350) );
  OAI211_X1 U9842 ( .C1(n8562), .C2(n8366), .A(n8351), .B(n8350), .ZN(P2_U3242) );
  NAND2_X1 U9843 ( .A1(n8494), .A2(n8352), .ZN(n8357) );
  NAND2_X1 U9844 ( .A1(n8354), .A2(n8353), .ZN(n8356) );
  MUX2_X1 U9845 ( .A(n8357), .B(n8356), .S(n8355), .Z(n8365) );
  OAI22_X1 U9846 ( .A1(n8360), .A2(n8359), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8358), .ZN(n8361) );
  AOI21_X1 U9847 ( .B1(n8363), .B2(n8362), .A(n8361), .ZN(n8364) );
  OAI211_X1 U9848 ( .C1(n8826), .C2(n8366), .A(n8365), .B(n8364), .ZN(P2_U3243) );
  MUX2_X1 U9849 ( .A(n8367), .B(P2_DATAO_REG_30__SCAN_IN), .S(n8384), .Z(
        P2_U3582) );
  MUX2_X1 U9850 ( .A(n8528), .B(P2_DATAO_REG_29__SCAN_IN), .S(n8384), .Z(
        P2_U3581) );
  MUX2_X1 U9851 ( .A(n8527), .B(P2_DATAO_REG_27__SCAN_IN), .S(n8384), .Z(
        P2_U3579) );
  MUX2_X1 U9852 ( .A(n8545), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8372), .Z(
        P2_U3578) );
  MUX2_X1 U9853 ( .A(n8506), .B(P2_DATAO_REG_25__SCAN_IN), .S(n8372), .Z(
        P2_U3577) );
  INV_X1 U9854 ( .A(n8368), .ZN(n8610) );
  MUX2_X1 U9855 ( .A(n8610), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8372), .Z(
        P2_U3576) );
  MUX2_X1 U9856 ( .A(n8656), .B(P2_DATAO_REG_22__SCAN_IN), .S(n8372), .Z(
        P2_U3574) );
  MUX2_X1 U9857 ( .A(n8670), .B(P2_DATAO_REG_21__SCAN_IN), .S(n8372), .Z(
        P2_U3573) );
  MUX2_X1 U9858 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8686), .S(P2_U3966), .Z(
        P2_U3572) );
  MUX2_X1 U9859 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8703), .S(P2_U3966), .Z(
        P2_U3571) );
  MUX2_X1 U9860 ( .A(n8685), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8372), .Z(
        P2_U3570) );
  MUX2_X1 U9861 ( .A(n8701), .B(P2_DATAO_REG_17__SCAN_IN), .S(n8372), .Z(
        P2_U3569) );
  MUX2_X1 U9862 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8498), .S(P2_U3966), .Z(
        P2_U3568) );
  MUX2_X1 U9863 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8494), .S(P2_U3966), .Z(
        P2_U3567) );
  MUX2_X1 U9864 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8369), .S(P2_U3966), .Z(
        P2_U3566) );
  INV_X1 U9865 ( .A(n8370), .ZN(n8371) );
  MUX2_X1 U9866 ( .A(n8371), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8372), .Z(
        P2_U3565) );
  MUX2_X1 U9867 ( .A(n8373), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8372), .Z(
        P2_U3564) );
  MUX2_X1 U9868 ( .A(n8374), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8384), .Z(
        P2_U3563) );
  MUX2_X1 U9869 ( .A(n8375), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8384), .Z(
        P2_U3562) );
  MUX2_X1 U9870 ( .A(n8376), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8384), .Z(
        P2_U3561) );
  MUX2_X1 U9871 ( .A(n8377), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8384), .Z(
        P2_U3560) );
  MUX2_X1 U9872 ( .A(n8378), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8384), .Z(
        P2_U3559) );
  MUX2_X1 U9873 ( .A(n8379), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8384), .Z(
        P2_U3558) );
  MUX2_X1 U9874 ( .A(n8380), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8384), .Z(
        P2_U3557) );
  MUX2_X1 U9875 ( .A(n8381), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8384), .Z(
        P2_U3556) );
  MUX2_X1 U9876 ( .A(n8382), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8384), .Z(
        P2_U3555) );
  MUX2_X1 U9877 ( .A(n8383), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8384), .Z(
        P2_U3554) );
  MUX2_X1 U9878 ( .A(n5020), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8384), .Z(
        P2_U3553) );
  MUX2_X1 U9879 ( .A(n8385), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8384), .Z(
        P2_U3552) );
  AOI211_X1 U9880 ( .C1(n8388), .C2(n8387), .A(n8386), .B(n10237), .ZN(n8389)
         );
  AOI21_X1 U9881 ( .B1(n9897), .B2(n8391), .A(n8389), .ZN(n8401) );
  NOR2_X1 U9882 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5268), .ZN(n8390) );
  AOI21_X1 U9883 ( .B1(n10234), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n8390), .ZN(
        n8400) );
  MUX2_X1 U9884 ( .A(n8392), .B(P2_REG1_REG_9__SCAN_IN), .S(n8391), .Z(n8395)
         );
  INV_X1 U9885 ( .A(n8393), .ZN(n8394) );
  NAND2_X1 U9886 ( .A1(n8395), .A2(n8394), .ZN(n8397) );
  OAI211_X1 U9887 ( .C1(n8398), .C2(n8397), .A(n8396), .B(n10232), .ZN(n8399)
         );
  NAND3_X1 U9888 ( .A1(n8401), .A2(n8400), .A3(n8399), .ZN(P2_U3254) );
  OAI21_X1 U9889 ( .B1(n8404), .B2(n8403), .A(n8402), .ZN(n8405) );
  NAND2_X1 U9890 ( .A1(n10233), .A2(n8405), .ZN(n8414) );
  NOR2_X1 U9891 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5317), .ZN(n8406) );
  AOI21_X1 U9892 ( .B1(n10234), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n8406), .ZN(
        n8413) );
  NAND2_X1 U9893 ( .A1(n9897), .A2(n8407), .ZN(n8412) );
  OAI211_X1 U9894 ( .C1(n8410), .C2(n8409), .A(n10232), .B(n8408), .ZN(n8411)
         );
  NAND4_X1 U9895 ( .A1(n8414), .A2(n8413), .A3(n8412), .A4(n8411), .ZN(
        P2_U3256) );
  NAND2_X1 U9896 ( .A1(n8416), .A2(n8415), .ZN(n8418) );
  NAND2_X1 U9897 ( .A1(n8418), .A2(n8417), .ZN(n8420) );
  XNOR2_X1 U9898 ( .A(n8437), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n8419) );
  NOR2_X1 U9899 ( .A1(n8420), .A2(n8419), .ZN(n8440) );
  AOI21_X1 U9900 ( .B1(n8420), .B2(n8419), .A(n8440), .ZN(n8432) );
  NOR2_X1 U9901 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9860), .ZN(n8421) );
  AOI21_X1 U9902 ( .B1(n10234), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n8421), .ZN(
        n8422) );
  INV_X1 U9903 ( .A(n8422), .ZN(n8430) );
  NAND2_X1 U9904 ( .A1(n8424), .A2(n8423), .ZN(n8426) );
  NAND2_X1 U9905 ( .A1(n8426), .A2(n8425), .ZN(n8428) );
  XNOR2_X1 U9906 ( .A(n8437), .B(P2_REG2_REG_16__SCAN_IN), .ZN(n8427) );
  NOR2_X1 U9907 ( .A1(n8428), .A2(n8427), .ZN(n8433) );
  AOI211_X1 U9908 ( .C1(n8428), .C2(n8427), .A(n10237), .B(n8433), .ZN(n8429)
         );
  AOI211_X1 U9909 ( .C1(n9897), .C2(n8437), .A(n8430), .B(n8429), .ZN(n8431)
         );
  OAI21_X1 U9910 ( .B1(n8432), .B2(n10236), .A(n8431), .ZN(P2_U3261) );
  AOI21_X1 U9911 ( .B1(P2_REG2_REG_16__SCAN_IN), .B2(n8437), .A(n8433), .ZN(
        n8436) );
  NAND2_X1 U9912 ( .A1(n8448), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8434) );
  OAI21_X1 U9913 ( .B1(n8448), .B2(P2_REG2_REG_17__SCAN_IN), .A(n8434), .ZN(
        n8435) );
  NOR2_X1 U9914 ( .A1(n8436), .A2(n8435), .ZN(n8447) );
  AOI211_X1 U9915 ( .C1(n8436), .C2(n8435), .A(n10237), .B(n8447), .ZN(n8446)
         );
  NOR2_X1 U9916 ( .A1(n8437), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n8439) );
  XNOR2_X1 U9917 ( .A(n8448), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n8438) );
  OAI21_X1 U9918 ( .B1(n8440), .B2(n8439), .A(n8438), .ZN(n8441) );
  OR3_X1 U9919 ( .A1(n8440), .A2(n8439), .A3(n8438), .ZN(n8454) );
  NAND3_X1 U9920 ( .A1(n8441), .A2(n10232), .A3(n8454), .ZN(n8444) );
  NOR2_X1 U9921 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5441), .ZN(n8442) );
  AOI21_X1 U9922 ( .B1(n10234), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n8442), .ZN(
        n8443) );
  OAI211_X1 U9923 ( .C1(n10235), .C2(n8455), .A(n8444), .B(n8443), .ZN(n8445)
         );
  OR2_X1 U9924 ( .A1(n8446), .A2(n8445), .ZN(P2_U3262) );
  INV_X1 U9925 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8449) );
  AOI21_X1 U9926 ( .B1(n8450), .B2(n8449), .A(n8467), .ZN(n8463) );
  NAND2_X1 U9927 ( .A1(n9897), .A2(n8457), .ZN(n8453) );
  NOR2_X1 U9928 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9804), .ZN(n8451) );
  AOI21_X1 U9929 ( .B1(n10234), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n8451), .ZN(
        n8452) );
  NAND2_X1 U9930 ( .A1(n8453), .A2(n8452), .ZN(n8462) );
  INV_X1 U9931 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8456) );
  OAI21_X1 U9932 ( .B1(n8456), .B2(n8455), .A(n8454), .ZN(n8459) );
  XNOR2_X1 U9933 ( .A(n8457), .B(P2_REG1_REG_18__SCAN_IN), .ZN(n8458) );
  NOR2_X1 U9934 ( .A1(n8459), .A2(n8458), .ZN(n8470) );
  AOI21_X1 U9935 ( .B1(n8459), .B2(n8458), .A(n8470), .ZN(n8460) );
  NOR2_X1 U9936 ( .A1(n8460), .A2(n10236), .ZN(n8461) );
  AOI211_X1 U9937 ( .C1(n10233), .C2(n8463), .A(n8462), .B(n8461), .ZN(n8464)
         );
  INV_X1 U9938 ( .A(n8464), .ZN(P2_U3263) );
  NOR2_X1 U9939 ( .A1(n8465), .A2(n8472), .ZN(n8466) );
  INV_X1 U9940 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8468) );
  XNOR2_X1 U9941 ( .A(n8469), .B(n8468), .ZN(n8477) );
  NAND2_X1 U9942 ( .A1(n8477), .A2(n10233), .ZN(n8475) );
  INV_X1 U9943 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8471) );
  AOI21_X1 U9944 ( .B1(n8472), .B2(n8471), .A(n8470), .ZN(n8473) );
  XNOR2_X1 U9945 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8473), .ZN(n8476) );
  AOI21_X1 U9946 ( .B1(n8476), .B2(n10232), .A(n9897), .ZN(n8474) );
  INV_X1 U9947 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n8480) );
  OAI21_X1 U9948 ( .B1(n8481), .B2(n8480), .A(n8479), .ZN(n8482) );
  INV_X1 U9949 ( .A(n9906), .ZN(n8490) );
  INV_X1 U9950 ( .A(n8816), .ZN(n8723) );
  NAND2_X1 U9951 ( .A1(n8717), .A2(n8697), .ZN(n8692) );
  NOR2_X2 U9952 ( .A1(n8678), .A2(n8799), .ZN(n8663) );
  NOR2_X2 U9953 ( .A1(n8582), .A2(n8768), .ZN(n8560) );
  XOR2_X1 U9954 ( .A(n8744), .B(n8489), .Z(n8746) );
  INV_X1 U9955 ( .A(P2_B_REG_SCAN_IN), .ZN(n9655) );
  OAI21_X1 U9956 ( .B1(n8484), .B2(n9655), .A(n8702), .ZN(n8518) );
  NOR2_X1 U9957 ( .A1(n8485), .A2(n8518), .ZN(n8743) );
  INV_X1 U9958 ( .A(n8743), .ZN(n9905) );
  NOR2_X1 U9959 ( .A1(n9905), .A2(n10266), .ZN(n8491) );
  AOI21_X1 U9960 ( .B1(n10266), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8491), .ZN(
        n8488) );
  NAND2_X1 U9961 ( .A1(n8744), .A2(n8486), .ZN(n8487) );
  OAI211_X1 U9962 ( .C1(n8746), .C2(n8550), .A(n8488), .B(n8487), .ZN(P2_U3265) );
  AOI21_X1 U9963 ( .B1(n8519), .B2(n8490), .A(n8489), .ZN(n9908) );
  NAND2_X1 U9964 ( .A1(n9908), .A2(n8707), .ZN(n8493) );
  AOI21_X1 U9965 ( .B1(n10266), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8491), .ZN(
        n8492) );
  OAI211_X1 U9966 ( .C1(n9906), .C2(n8733), .A(n8493), .B(n8492), .ZN(P2_U3266) );
  NAND2_X1 U9967 ( .A1(n8809), .A2(n8685), .ZN(n8501) );
  NAND2_X1 U9968 ( .A1(n8677), .A2(n8676), .ZN(n8675) );
  NAND2_X1 U9969 ( .A1(n8675), .A2(n5090), .ZN(n8662) );
  NAND2_X1 U9970 ( .A1(n8585), .A2(n8572), .ZN(n8507) );
  NAND2_X1 U9971 ( .A1(n8558), .A2(n8570), .ZN(n8557) );
  NAND2_X1 U9972 ( .A1(n8562), .A2(n8508), .ZN(n8509) );
  NAND2_X1 U9973 ( .A1(n8557), .A2(n8509), .ZN(n8541) );
  NAND2_X1 U9974 ( .A1(n8541), .A2(n8540), .ZN(n8539) );
  NAND2_X1 U9975 ( .A1(n8760), .A2(n8573), .ZN(n8510) );
  NAND2_X1 U9976 ( .A1(n8531), .A2(n8530), .ZN(n8529) );
  INV_X1 U9977 ( .A(n8755), .ZN(n8535) );
  NAND2_X1 U9978 ( .A1(n8535), .A2(n8548), .ZN(n8511) );
  NAND2_X1 U9979 ( .A1(n8529), .A2(n8511), .ZN(n8512) );
  XNOR2_X1 U9980 ( .A(n8512), .B(n8515), .ZN(n8747) );
  INV_X1 U9981 ( .A(n8747), .ZN(n8525) );
  AOI21_X1 U9982 ( .B1(n8515), .B2(n8514), .A(n8513), .ZN(n8516) );
  OAI222_X1 U9983 ( .A1(n8637), .A2(n8548), .B1(n8518), .B2(n8517), .C1(n8516), 
        .C2(n8715), .ZN(n8751) );
  OAI21_X1 U9984 ( .B1(n8532), .B2(n8748), .A(n8519), .ZN(n8749) );
  NOR2_X1 U9985 ( .A1(n8749), .A2(n8550), .ZN(n8523) );
  AOI22_X1 U9986 ( .A1(n8520), .A2(n10257), .B1(P2_REG2_REG_29__SCAN_IN), .B2(
        n10266), .ZN(n8521) );
  OAI21_X1 U9987 ( .B1(n8748), .B2(n8733), .A(n8521), .ZN(n8522) );
  AOI211_X1 U9988 ( .C1(n8751), .C2(n10263), .A(n8523), .B(n8522), .ZN(n8524)
         );
  OAI21_X1 U9989 ( .B1(n8525), .B2(n8742), .A(n8524), .ZN(P2_U3267) );
  OAI21_X1 U9990 ( .B1(n8531), .B2(n8530), .A(n8529), .ZN(n8754) );
  NAND2_X1 U9991 ( .A1(n8754), .A2(n8615), .ZN(n8538) );
  AOI21_X1 U9992 ( .B1(n8755), .B2(n8549), .A(n8532), .ZN(n8756) );
  AOI22_X1 U9993 ( .A1(n8533), .A2(n10257), .B1(P2_REG2_REG_28__SCAN_IN), .B2(
        n10266), .ZN(n8534) );
  OAI21_X1 U9994 ( .B1(n8535), .B2(n8733), .A(n8534), .ZN(n8536) );
  AOI21_X1 U9995 ( .B1(n8756), .B2(n8707), .A(n8536), .ZN(n8537) );
  OAI211_X1 U9996 ( .C1(n10266), .C2(n8758), .A(n8538), .B(n8537), .ZN(
        P2_U3268) );
  OAI21_X1 U9997 ( .B1(n8541), .B2(n8540), .A(n8539), .ZN(n8764) );
  INV_X1 U9998 ( .A(n8764), .ZN(n8556) );
  OAI211_X1 U9999 ( .C1(n8544), .C2(n8543), .A(n8542), .B(n10254), .ZN(n8547)
         );
  NAND2_X1 U10000 ( .A1(n8545), .A2(n8700), .ZN(n8546) );
  OAI211_X1 U10001 ( .C1(n8548), .C2(n8639), .A(n8547), .B(n8546), .ZN(n8763)
         );
  OAI21_X1 U10002 ( .B1(n8560), .B2(n8760), .A(n8549), .ZN(n8761) );
  NOR2_X1 U10003 ( .A1(n8761), .A2(n8550), .ZN(n8554) );
  AOI22_X1 U10004 ( .A1(n8551), .A2(n10257), .B1(P2_REG2_REG_27__SCAN_IN), 
        .B2(n10266), .ZN(n8552) );
  OAI21_X1 U10005 ( .B1(n8760), .B2(n8733), .A(n8552), .ZN(n8553) );
  AOI211_X1 U10006 ( .C1(n8763), .C2(n10263), .A(n8554), .B(n8553), .ZN(n8555)
         );
  OAI21_X1 U10007 ( .B1(n8556), .B2(n8742), .A(n8555), .ZN(P2_U3269) );
  OAI21_X1 U10008 ( .B1(n8558), .B2(n8570), .A(n8557), .ZN(n8559) );
  INV_X1 U10009 ( .A(n8559), .ZN(n8770) );
  AOI211_X1 U10010 ( .C1(n8768), .C2(n8582), .A(n10336), .B(n8560), .ZN(n8767)
         );
  INV_X1 U10011 ( .A(n8561), .ZN(n8719) );
  NOR2_X1 U10012 ( .A1(n8562), .A2(n8733), .ZN(n8566) );
  OAI22_X1 U10013 ( .A1(n8564), .A2(n8620), .B1(n8563), .B2(n10263), .ZN(n8565) );
  AOI211_X1 U10014 ( .C1(n8767), .C2(n8719), .A(n8566), .B(n8565), .ZN(n8575)
         );
  INV_X1 U10015 ( .A(n8567), .ZN(n8568) );
  OAI222_X1 U10016 ( .A1(n8639), .A2(n8573), .B1(n8637), .B2(n8572), .C1(n8715), .C2(n8571), .ZN(n8766) );
  NAND2_X1 U10017 ( .A1(n8766), .A2(n10263), .ZN(n8574) );
  OAI211_X1 U10018 ( .C1(n8770), .C2(n8742), .A(n8575), .B(n8574), .ZN(
        P2_U3270) );
  XNOR2_X1 U10019 ( .A(n8576), .B(n8580), .ZN(n8578) );
  AOI21_X1 U10020 ( .B1(n8578), .B2(n10254), .A(n8577), .ZN(n8775) );
  OAI21_X1 U10021 ( .B1(n8581), .B2(n8580), .A(n8579), .ZN(n8771) );
  NAND2_X1 U10022 ( .A1(n8771), .A2(n8615), .ZN(n8591) );
  INV_X1 U10023 ( .A(n8599), .ZN(n8584) );
  INV_X1 U10024 ( .A(n8582), .ZN(n8583) );
  AOI211_X1 U10025 ( .C1(n8773), .C2(n8584), .A(n10336), .B(n8583), .ZN(n8772)
         );
  NOR2_X1 U10026 ( .A1(n8585), .A2(n8733), .ZN(n8589) );
  OAI22_X1 U10027 ( .A1(n8587), .A2(n8620), .B1(n8586), .B2(n10263), .ZN(n8588) );
  AOI211_X1 U10028 ( .C1(n8772), .C2(n8719), .A(n8589), .B(n8588), .ZN(n8590)
         );
  OAI211_X1 U10029 ( .C1(n10266), .C2(n8775), .A(n8591), .B(n8590), .ZN(
        P2_U3271) );
  AOI21_X1 U10030 ( .B1(n8592), .B2(n8597), .A(n8715), .ZN(n8595) );
  AOI21_X1 U10031 ( .B1(n8595), .B2(n8594), .A(n8593), .ZN(n8781) );
  OAI21_X1 U10032 ( .B1(n8598), .B2(n8597), .A(n8596), .ZN(n8777) );
  NAND2_X1 U10033 ( .A1(n8777), .A2(n8615), .ZN(n8604) );
  AOI21_X1 U10034 ( .B1(n8778), .B2(n8616), .A(n8599), .ZN(n8779) );
  AOI22_X1 U10035 ( .A1(n8600), .A2(n10257), .B1(P2_REG2_REG_24__SCAN_IN), 
        .B2(n10266), .ZN(n8601) );
  OAI21_X1 U10036 ( .B1(n4720), .B2(n8733), .A(n8601), .ZN(n8602) );
  AOI21_X1 U10037 ( .B1(n8779), .B2(n8707), .A(n8602), .ZN(n8603) );
  OAI211_X1 U10038 ( .C1(n10266), .C2(n8781), .A(n8604), .B(n8603), .ZN(
        P2_U3272) );
  INV_X1 U10039 ( .A(n8605), .ZN(n8636) );
  OAI21_X1 U10040 ( .B1(n8636), .B2(n8607), .A(n8606), .ZN(n8609) );
  NAND2_X1 U10041 ( .A1(n8609), .A2(n8608), .ZN(n8611) );
  AOI222_X1 U10042 ( .A1(n10254), .A2(n8611), .B1(n8610), .B2(n8702), .C1(
        n8656), .C2(n8700), .ZN(n8787) );
  AOI21_X1 U10043 ( .B1(n8614), .B2(n8613), .A(n8612), .ZN(n8783) );
  NAND2_X1 U10044 ( .A1(n8783), .A2(n8615), .ZN(n8625) );
  INV_X1 U10045 ( .A(n8616), .ZN(n8617) );
  AOI21_X1 U10046 ( .B1(n8784), .B2(n4723), .A(n8617), .ZN(n8785) );
  NOR2_X1 U10047 ( .A1(n8618), .A2(n8733), .ZN(n8623) );
  OAI22_X1 U10048 ( .A1(n8621), .A2(n8620), .B1(n8619), .B2(n10263), .ZN(n8622) );
  AOI211_X1 U10049 ( .C1(n8785), .C2(n8707), .A(n8623), .B(n8622), .ZN(n8624)
         );
  OAI211_X1 U10050 ( .C1(n10266), .C2(n8787), .A(n8625), .B(n8624), .ZN(
        P2_U3273) );
  XNOR2_X1 U10051 ( .A(n8627), .B(n8626), .ZN(n8793) );
  AOI21_X1 U10052 ( .B1(n8789), .B2(n8647), .A(n8628), .ZN(n8790) );
  INV_X1 U10053 ( .A(n8629), .ZN(n8630) );
  AOI22_X1 U10054 ( .A1(n8630), .A2(n10257), .B1(n10266), .B2(
        P2_REG2_REG_22__SCAN_IN), .ZN(n8631) );
  OAI21_X1 U10055 ( .B1(n8632), .B2(n8733), .A(n8631), .ZN(n8644) );
  AOI21_X1 U10056 ( .B1(n8654), .B2(n8634), .A(n8633), .ZN(n8635) );
  NOR3_X1 U10057 ( .A1(n8636), .A2(n8635), .A3(n8715), .ZN(n8642) );
  OAI22_X1 U10058 ( .A1(n8640), .A2(n8639), .B1(n8638), .B2(n8637), .ZN(n8641)
         );
  NOR2_X1 U10059 ( .A1(n8642), .A2(n8641), .ZN(n8792) );
  NOR2_X1 U10060 ( .A1(n8792), .A2(n10266), .ZN(n8643) );
  AOI211_X1 U10061 ( .C1(n8790), .C2(n8707), .A(n8644), .B(n8643), .ZN(n8645)
         );
  OAI21_X1 U10062 ( .B1(n8793), .B2(n8742), .A(n8645), .ZN(P2_U3274) );
  XNOR2_X1 U10063 ( .A(n8646), .B(n8653), .ZN(n8798) );
  INV_X1 U10064 ( .A(n8663), .ZN(n8649) );
  INV_X1 U10065 ( .A(n8647), .ZN(n8648) );
  AOI21_X1 U10066 ( .B1(n8794), .B2(n8649), .A(n8648), .ZN(n8795) );
  AOI22_X1 U10067 ( .A1(n10266), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8650), 
        .B2(n10257), .ZN(n8651) );
  OAI21_X1 U10068 ( .B1(n8652), .B2(n8733), .A(n8651), .ZN(n8659) );
  OAI21_X1 U10069 ( .B1(n8655), .B2(n5519), .A(n8654), .ZN(n8657) );
  AOI222_X1 U10070 ( .A1(n10254), .A2(n8657), .B1(n8656), .B2(n8702), .C1(
        n8686), .C2(n8700), .ZN(n8797) );
  NOR2_X1 U10071 ( .A1(n8797), .A2(n10266), .ZN(n8658) );
  AOI211_X1 U10072 ( .C1(n8795), .C2(n8707), .A(n8659), .B(n8658), .ZN(n8660)
         );
  OAI21_X1 U10073 ( .B1(n8798), .B2(n8742), .A(n8660), .ZN(P2_U3275) );
  OAI21_X1 U10074 ( .B1(n8662), .B2(n8669), .A(n8661), .ZN(n8803) );
  AOI21_X1 U10075 ( .B1(n8799), .B2(n8678), .A(n8663), .ZN(n8800) );
  AOI22_X1 U10076 ( .A1(n10266), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8664), 
        .B2(n10257), .ZN(n8665) );
  OAI21_X1 U10077 ( .B1(n8666), .B2(n8733), .A(n8665), .ZN(n8673) );
  NAND2_X1 U10078 ( .A1(n8683), .A2(n8667), .ZN(n8668) );
  XOR2_X1 U10079 ( .A(n8669), .B(n8668), .Z(n8671) );
  AOI222_X1 U10080 ( .A1(n10254), .A2(n8671), .B1(n8703), .B2(n8700), .C1(
        n8670), .C2(n8702), .ZN(n8802) );
  NOR2_X1 U10081 ( .A1(n8802), .A2(n10266), .ZN(n8672) );
  AOI211_X1 U10082 ( .C1(n8800), .C2(n8707), .A(n8673), .B(n8672), .ZN(n8674)
         );
  OAI21_X1 U10083 ( .B1(n8742), .B2(n8803), .A(n8674), .ZN(P2_U3276) );
  OAI21_X1 U10084 ( .B1(n8677), .B2(n8676), .A(n8675), .ZN(n8808) );
  INV_X1 U10085 ( .A(n8678), .ZN(n8679) );
  AOI211_X1 U10086 ( .C1(n8805), .C2(n8692), .A(n10336), .B(n8679), .ZN(n8804)
         );
  AOI22_X1 U10087 ( .A1(n10266), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n8680), 
        .B2(n10257), .ZN(n8681) );
  OAI21_X1 U10088 ( .B1(n8682), .B2(n8733), .A(n8681), .ZN(n8689) );
  OAI21_X1 U10089 ( .B1(n8684), .B2(n4568), .A(n8683), .ZN(n8687) );
  AOI222_X1 U10090 ( .A1(n10254), .A2(n8687), .B1(n8686), .B2(n8702), .C1(
        n8685), .C2(n8700), .ZN(n8807) );
  NOR2_X1 U10091 ( .A1(n8807), .A2(n10266), .ZN(n8688) );
  AOI211_X1 U10092 ( .C1(n8804), .C2(n8719), .A(n8689), .B(n8688), .ZN(n8690)
         );
  OAI21_X1 U10093 ( .B1(n8742), .B2(n8808), .A(n8690), .ZN(P2_U3277) );
  XNOR2_X1 U10094 ( .A(n8691), .B(n8699), .ZN(n8813) );
  INV_X1 U10095 ( .A(n8717), .ZN(n8694) );
  INV_X1 U10096 ( .A(n8692), .ZN(n8693) );
  AOI21_X1 U10097 ( .B1(n8809), .B2(n8694), .A(n8693), .ZN(n8810) );
  AOI22_X1 U10098 ( .A1(n10266), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8695), 
        .B2(n10257), .ZN(n8696) );
  OAI21_X1 U10099 ( .B1(n8697), .B2(n8733), .A(n8696), .ZN(n8706) );
  XOR2_X1 U10100 ( .A(n8699), .B(n8698), .Z(n8704) );
  AOI222_X1 U10101 ( .A1(n10254), .A2(n8704), .B1(n8703), .B2(n8702), .C1(
        n8701), .C2(n8700), .ZN(n8812) );
  NOR2_X1 U10102 ( .A1(n8812), .A2(n10266), .ZN(n8705) );
  AOI211_X1 U10103 ( .C1(n8810), .C2(n8707), .A(n8706), .B(n8705), .ZN(n8708)
         );
  OAI21_X1 U10104 ( .B1(n8813), .B2(n8742), .A(n8708), .ZN(P2_U3278) );
  OAI21_X1 U10105 ( .B1(n8709), .B2(n8712), .A(n8710), .ZN(n8711) );
  INV_X1 U10106 ( .A(n8711), .ZN(n8818) );
  XNOR2_X1 U10107 ( .A(n8713), .B(n8712), .ZN(n8716) );
  OAI21_X1 U10108 ( .B1(n8716), .B2(n8715), .A(n8714), .ZN(n8814) );
  INV_X1 U10109 ( .A(n8730), .ZN(n8718) );
  AOI211_X1 U10110 ( .C1(n8816), .C2(n8718), .A(n10336), .B(n8717), .ZN(n8815)
         );
  NAND2_X1 U10111 ( .A1(n8815), .A2(n8719), .ZN(n8722) );
  AOI22_X1 U10112 ( .A1(n10266), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n8720), 
        .B2(n10257), .ZN(n8721) );
  OAI211_X1 U10113 ( .C1(n8723), .C2(n8733), .A(n8722), .B(n8721), .ZN(n8724)
         );
  AOI21_X1 U10114 ( .B1(n8814), .B2(n10263), .A(n8724), .ZN(n8725) );
  OAI21_X1 U10115 ( .B1(n8818), .B2(n8742), .A(n8725), .ZN(P2_U3279) );
  AOI21_X1 U10116 ( .B1(n8728), .B2(n8727), .A(n8726), .ZN(n8729) );
  INV_X1 U10117 ( .A(n8729), .ZN(n8823) );
  AOI211_X1 U10118 ( .C1(n8820), .C2(n4488), .A(n10336), .B(n8730), .ZN(n8819)
         );
  INV_X1 U10119 ( .A(n8820), .ZN(n8734) );
  AOI22_X1 U10120 ( .A1(n10266), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n8731), 
        .B2(n10257), .ZN(n8732) );
  OAI21_X1 U10121 ( .B1(n8734), .B2(n8733), .A(n8732), .ZN(n8740) );
  XNOR2_X1 U10122 ( .A(n8736), .B(n8735), .ZN(n8738) );
  AOI21_X1 U10123 ( .B1(n8738), .B2(n10254), .A(n8737), .ZN(n8822) );
  NOR2_X1 U10124 ( .A1(n8822), .A2(n10266), .ZN(n8739) );
  AOI211_X1 U10125 ( .C1(n8819), .C2(n8719), .A(n8740), .B(n8739), .ZN(n8741)
         );
  OAI21_X1 U10126 ( .B1(n8823), .B2(n8742), .A(n8741), .ZN(P2_U3280) );
  AOI21_X1 U10127 ( .B1(n8744), .B2(n10284), .A(n8743), .ZN(n8745) );
  OAI21_X1 U10128 ( .B1(n8746), .B2(n10336), .A(n8745), .ZN(n8843) );
  MUX2_X1 U10129 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n8843), .S(n10360), .Z(
        P2_U3551) );
  NAND2_X1 U10130 ( .A1(n8747), .A2(n10340), .ZN(n8753) );
  OAI22_X1 U10131 ( .A1(n8749), .A2(n10336), .B1(n8748), .B2(n10335), .ZN(
        n8750) );
  NAND2_X1 U10132 ( .A1(n8753), .A2(n8752), .ZN(n8844) );
  MUX2_X1 U10133 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n8844), .S(n10360), .Z(
        P2_U3549) );
  NAND2_X1 U10134 ( .A1(n8754), .A2(n10340), .ZN(n8759) );
  AOI22_X1 U10135 ( .A1(n8756), .A2(n10246), .B1(n10284), .B2(n8755), .ZN(
        n8757) );
  OAI22_X1 U10136 ( .A1(n8761), .A2(n10336), .B1(n8760), .B2(n10335), .ZN(
        n8762) );
  AOI211_X1 U10137 ( .C1(n8764), .C2(n10340), .A(n8763), .B(n8762), .ZN(n8765)
         );
  INV_X1 U10138 ( .A(n8765), .ZN(n8846) );
  MUX2_X1 U10139 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8846), .S(n10360), .Z(
        P2_U3547) );
  OAI21_X1 U10140 ( .B1(n8770), .B2(n10288), .A(n8769), .ZN(n8847) );
  MUX2_X1 U10141 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n8847), .S(n10360), .Z(
        P2_U3546) );
  INV_X1 U10142 ( .A(n8771), .ZN(n8776) );
  AOI21_X1 U10143 ( .B1(n10284), .B2(n8773), .A(n8772), .ZN(n8774) );
  OAI211_X1 U10144 ( .C1(n8776), .C2(n10288), .A(n8775), .B(n8774), .ZN(n8848)
         );
  MUX2_X1 U10145 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8848), .S(n10360), .Z(
        P2_U3545) );
  INV_X1 U10146 ( .A(n8777), .ZN(n8782) );
  AOI22_X1 U10147 ( .A1(n8779), .A2(n10246), .B1(n10284), .B2(n8778), .ZN(
        n8780) );
  OAI211_X1 U10148 ( .C1(n8782), .C2(n10288), .A(n8781), .B(n8780), .ZN(n8849)
         );
  MUX2_X1 U10149 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8849), .S(n10360), .Z(
        P2_U3544) );
  INV_X1 U10150 ( .A(n8783), .ZN(n8788) );
  AOI22_X1 U10151 ( .A1(n8785), .A2(n10246), .B1(n10284), .B2(n8784), .ZN(
        n8786) );
  OAI211_X1 U10152 ( .C1(n8788), .C2(n10288), .A(n8787), .B(n8786), .ZN(n8850)
         );
  MUX2_X1 U10153 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8850), .S(n10360), .Z(
        P2_U3543) );
  AOI22_X1 U10154 ( .A1(n8790), .A2(n10246), .B1(n10284), .B2(n8789), .ZN(
        n8791) );
  OAI211_X1 U10155 ( .C1(n8793), .C2(n10288), .A(n8792), .B(n8791), .ZN(n8851)
         );
  MUX2_X1 U10156 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n8851), .S(n10360), .Z(
        P2_U3542) );
  AOI22_X1 U10157 ( .A1(n8795), .A2(n10246), .B1(n10284), .B2(n8794), .ZN(
        n8796) );
  OAI211_X1 U10158 ( .C1(n8798), .C2(n10288), .A(n8797), .B(n8796), .ZN(n8852)
         );
  MUX2_X1 U10159 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n8852), .S(n10360), .Z(
        P2_U3541) );
  AOI22_X1 U10160 ( .A1(n8800), .A2(n10246), .B1(n10284), .B2(n8799), .ZN(
        n8801) );
  OAI211_X1 U10161 ( .C1(n8803), .C2(n10288), .A(n8802), .B(n8801), .ZN(n8853)
         );
  MUX2_X1 U10162 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n8853), .S(n10360), .Z(
        P2_U3540) );
  AOI21_X1 U10163 ( .B1(n10284), .B2(n8805), .A(n8804), .ZN(n8806) );
  OAI211_X1 U10164 ( .C1(n8808), .C2(n10288), .A(n8807), .B(n8806), .ZN(n8854)
         );
  MUX2_X1 U10165 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8854), .S(n10360), .Z(
        P2_U3539) );
  AOI22_X1 U10166 ( .A1(n8810), .A2(n10246), .B1(n10284), .B2(n8809), .ZN(
        n8811) );
  OAI211_X1 U10167 ( .C1(n8813), .C2(n10288), .A(n8812), .B(n8811), .ZN(n8855)
         );
  MUX2_X1 U10168 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n8855), .S(n10360), .Z(
        P2_U3538) );
  AOI211_X1 U10169 ( .C1(n10284), .C2(n8816), .A(n8815), .B(n8814), .ZN(n8817)
         );
  OAI21_X1 U10170 ( .B1(n8818), .B2(n10288), .A(n8817), .ZN(n8856) );
  MUX2_X1 U10171 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8856), .S(n10360), .Z(
        P2_U3537) );
  AOI21_X1 U10172 ( .B1(n10284), .B2(n8820), .A(n8819), .ZN(n8821) );
  OAI211_X1 U10173 ( .C1(n8823), .C2(n10288), .A(n8822), .B(n8821), .ZN(n8857)
         );
  MUX2_X1 U10174 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8857), .S(n10360), .Z(
        P2_U3536) );
  INV_X1 U10175 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8829) );
  OAI211_X1 U10176 ( .C1(n8826), .C2(n10335), .A(n8825), .B(n8824), .ZN(n8827)
         );
  AOI21_X1 U10177 ( .B1(n8828), .B2(n10340), .A(n8827), .ZN(n8858) );
  MUX2_X1 U10178 ( .A(n8829), .B(n8858), .S(n10360), .Z(n8830) );
  INV_X1 U10179 ( .A(n8830), .ZN(P2_U3535) );
  INV_X1 U10180 ( .A(n8831), .ZN(n10333) );
  OAI22_X1 U10181 ( .A1(n8833), .A2(n10336), .B1(n8832), .B2(n10335), .ZN(
        n8834) );
  AOI21_X1 U10182 ( .B1(n8835), .B2(n10333), .A(n8834), .ZN(n8836) );
  NAND2_X1 U10183 ( .A1(n8837), .A2(n8836), .ZN(n8861) );
  MUX2_X1 U10184 ( .A(n8861), .B(P2_REG1_REG_13__SCAN_IN), .S(n10357), .Z(
        P2_U3533) );
  AOI211_X1 U10185 ( .C1(n10284), .C2(n8840), .A(n8839), .B(n8838), .ZN(n8841)
         );
  OAI21_X1 U10186 ( .B1(n10288), .B2(n8842), .A(n8841), .ZN(n8862) );
  MUX2_X1 U10187 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n8862), .S(n10360), .Z(
        P2_U3531) );
  MUX2_X1 U10188 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n8843), .S(n10344), .Z(
        P2_U3519) );
  MUX2_X1 U10189 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n8844), .S(n10344), .Z(
        P2_U3517) );
  MUX2_X1 U10190 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n8845), .S(n10344), .Z(
        P2_U3516) );
  MUX2_X1 U10191 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8846), .S(n10344), .Z(
        P2_U3515) );
  MUX2_X1 U10192 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n8847), .S(n10344), .Z(
        P2_U3514) );
  MUX2_X1 U10193 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n8848), .S(n10344), .Z(
        P2_U3513) );
  MUX2_X1 U10194 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n8849), .S(n10344), .Z(
        P2_U3512) );
  MUX2_X1 U10195 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n8850), .S(n10344), .Z(
        P2_U3511) );
  MUX2_X1 U10196 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n8851), .S(n10344), .Z(
        P2_U3510) );
  MUX2_X1 U10197 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n8852), .S(n10344), .Z(
        P2_U3509) );
  MUX2_X1 U10198 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n8853), .S(n10344), .Z(
        P2_U3508) );
  MUX2_X1 U10199 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n8854), .S(n10344), .Z(
        P2_U3507) );
  MUX2_X1 U10200 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n8855), .S(n10344), .Z(
        P2_U3505) );
  MUX2_X1 U10201 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n8856), .S(n10344), .Z(
        P2_U3502) );
  MUX2_X1 U10202 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n8857), .S(n10344), .Z(
        P2_U3499) );
  INV_X1 U10203 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n8859) );
  MUX2_X1 U10204 ( .A(n8859), .B(n8858), .S(n10344), .Z(n8860) );
  INV_X1 U10205 ( .A(n8860), .ZN(P2_U3496) );
  MUX2_X1 U10206 ( .A(P2_REG0_REG_13__SCAN_IN), .B(n8861), .S(n10344), .Z(
        P2_U3490) );
  MUX2_X1 U10207 ( .A(P2_REG0_REG_11__SCAN_IN), .B(n8862), .S(n10344), .Z(
        P2_U3484) );
  INV_X1 U10208 ( .A(n8863), .ZN(n9488) );
  NAND3_X1 U10209 ( .A1(n8864), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n8867) );
  OAI22_X1 U10210 ( .A1(n8868), .A2(n8867), .B1(n8866), .B2(n8865), .ZN(n8869)
         );
  INV_X1 U10211 ( .A(n8869), .ZN(n8870) );
  OAI21_X1 U10212 ( .B1(n9488), .B2(n8871), .A(n8870), .ZN(P2_U3327) );
  INV_X1 U10213 ( .A(n8872), .ZN(n9491) );
  OAI222_X1 U10214 ( .A1(n8876), .A2(n8875), .B1(n8874), .B2(n9491), .C1(n8873), .C2(P2_U3152), .ZN(P2_U3329) );
  MUX2_X1 U10215 ( .A(n8877), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  XNOR2_X1 U10216 ( .A(n8879), .B(n8878), .ZN(n8880) );
  XNOR2_X1 U10217 ( .A(n8881), .B(n8880), .ZN(n8887) );
  OAI22_X1 U10218 ( .A1(n9093), .A2(n8960), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8882), .ZN(n8883) );
  AOI21_X1 U10219 ( .B1(n9160), .B2(n8962), .A(n8883), .ZN(n8884) );
  OAI21_X1 U10220 ( .B1(n9096), .B2(n8981), .A(n8884), .ZN(n8885) );
  AOI21_X1 U10221 ( .B1(n9405), .B2(n9007), .A(n8885), .ZN(n8886) );
  OAI21_X1 U10222 ( .B1(n8887), .B2(n9009), .A(n8886), .ZN(P1_U3212) );
  XNOR2_X1 U10223 ( .A(n8889), .B(n8888), .ZN(n8890) );
  XNOR2_X1 U10224 ( .A(n8891), .B(n8890), .ZN(n8899) );
  OR2_X1 U10225 ( .A1(n9089), .A2(n9238), .ZN(n8893) );
  NAND2_X1 U10226 ( .A1(n9083), .A2(n9368), .ZN(n8892) );
  NAND2_X1 U10227 ( .A1(n8893), .A2(n8892), .ZN(n9214) );
  NAND2_X1 U10228 ( .A1(n9214), .A2(n9003), .ZN(n8895) );
  NAND2_X1 U10229 ( .A1(n8962), .A2(n9210), .ZN(n8894) );
  OAI211_X1 U10230 ( .C1(P1_STATE_REG_SCAN_IN), .C2(n8896), .A(n8895), .B(
        n8894), .ZN(n8897) );
  AOI21_X1 U10231 ( .B1(n9426), .B2(n9007), .A(n8897), .ZN(n8898) );
  OAI21_X1 U10232 ( .B1(n8899), .B2(n9009), .A(n8898), .ZN(P1_U3214) );
  INV_X1 U10233 ( .A(n9447), .ZN(n9272) );
  NOR2_X1 U10234 ( .A1(n8900), .A2(n5058), .ZN(n8905) );
  AOI21_X1 U10235 ( .B1(n8903), .B2(n8902), .A(n8901), .ZN(n8904) );
  OAI21_X1 U10236 ( .B1(n8905), .B2(n8904), .A(n8956), .ZN(n8910) );
  NOR2_X1 U10237 ( .A1(n8906), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9057) );
  AOI21_X1 U10238 ( .B1(n8971), .B2(n9276), .A(n9057), .ZN(n8907) );
  OAI21_X1 U10239 ( .B1(n9011), .B2(n8960), .A(n8907), .ZN(n8908) );
  AOI21_X1 U10240 ( .B1(n9270), .B2(n8962), .A(n8908), .ZN(n8909) );
  OAI211_X1 U10241 ( .C1(n9272), .C2(n8996), .A(n8910), .B(n8909), .ZN(
        P1_U3217) );
  XOR2_X1 U10242 ( .A(n8912), .B(n8911), .Z(n8919) );
  AND2_X1 U10243 ( .A1(n9276), .A2(n9368), .ZN(n8913) );
  AOI21_X1 U10244 ( .B1(n9083), .B2(n9370), .A(n8913), .ZN(n9245) );
  OAI22_X1 U10245 ( .A1(n9245), .A2(n8915), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8914), .ZN(n8916) );
  AOI21_X1 U10246 ( .B1(n9249), .B2(n8962), .A(n8916), .ZN(n8918) );
  NAND2_X1 U10247 ( .A1(n9439), .A2(n9007), .ZN(n8917) );
  OAI211_X1 U10248 ( .C1(n8919), .C2(n9009), .A(n8918), .B(n8917), .ZN(
        P1_U3221) );
  XOR2_X1 U10249 ( .A(n8921), .B(n8920), .Z(n8926) );
  OAI22_X1 U10250 ( .A1(n9093), .A2(n9238), .B1(n9089), .B2(n9236), .ZN(n9189)
         );
  OAI22_X1 U10251 ( .A1(n9183), .A2(n9005), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8922), .ZN(n8924) );
  NOR2_X1 U10252 ( .A1(n9186), .A2(n8996), .ZN(n8923) );
  AOI211_X1 U10253 ( .C1(n9003), .C2(n9189), .A(n8924), .B(n8923), .ZN(n8925)
         );
  OAI21_X1 U10254 ( .B1(n8926), .B2(n9009), .A(n8925), .ZN(P1_U3223) );
  INV_X1 U10255 ( .A(n9323), .ZN(n9922) );
  INV_X1 U10256 ( .A(n8927), .ZN(n8931) );
  AOI21_X1 U10257 ( .B1(n8928), .B2(n8998), .A(n8929), .ZN(n8930) );
  OAI21_X1 U10258 ( .B1(n8931), .B2(n8930), .A(n8956), .ZN(n8936) );
  INV_X1 U10259 ( .A(n8932), .ZN(n9313) );
  NAND2_X1 U10260 ( .A1(P1_REG3_REG_16__SCAN_IN), .A2(P1_U3084), .ZN(n10083)
         );
  OAI21_X1 U10261 ( .B1(n8981), .B2(n9078), .A(n10083), .ZN(n8934) );
  NOR2_X1 U10262 ( .A1(n9005), .A2(n9320), .ZN(n8933) );
  AOI211_X1 U10263 ( .C1(n8983), .C2(n9313), .A(n8934), .B(n8933), .ZN(n8935)
         );
  OAI211_X1 U10264 ( .C1(n9922), .C2(n8996), .A(n8936), .B(n8935), .ZN(
        P1_U3224) );
  INV_X1 U10265 ( .A(n9458), .ZN(n9302) );
  OAI21_X1 U10266 ( .B1(n8939), .B2(n8937), .A(n8938), .ZN(n8940) );
  NAND2_X1 U10267 ( .A1(n8940), .A2(n8956), .ZN(n8945) );
  OR2_X1 U10268 ( .A1(n9011), .A2(n9238), .ZN(n8942) );
  OR2_X1 U10269 ( .A1(n9012), .A2(n9236), .ZN(n8941) );
  NAND2_X1 U10270 ( .A1(n8942), .A2(n8941), .ZN(n9305) );
  AND2_X1 U10271 ( .A1(P1_U3084), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n10100) );
  NOR2_X1 U10272 ( .A1(n9005), .A2(n9299), .ZN(n8943) );
  AOI211_X1 U10273 ( .C1(n9003), .C2(n9305), .A(n10100), .B(n8943), .ZN(n8944)
         );
  OAI211_X1 U10274 ( .C1(n9302), .C2(n8996), .A(n8945), .B(n8944), .ZN(
        P1_U3226) );
  XOR2_X1 U10275 ( .A(n8947), .B(n8946), .Z(n8952) );
  NOR2_X1 U10276 ( .A1(n9205), .A2(n9005), .ZN(n8950) );
  AOI22_X1 U10277 ( .A1(n9198), .A2(n8983), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3084), .ZN(n8948) );
  OAI21_X1 U10278 ( .B1(n9092), .B2(n8981), .A(n8948), .ZN(n8949) );
  AOI211_X1 U10279 ( .C1(n9421), .C2(n9007), .A(n8950), .B(n8949), .ZN(n8951)
         );
  OAI21_X1 U10280 ( .B1(n8952), .B2(n9009), .A(n8951), .ZN(P1_U3227) );
  OAI21_X1 U10281 ( .B1(n8955), .B2(n8954), .A(n8953), .ZN(n8957) );
  NAND2_X1 U10282 ( .A1(n8957), .A2(n8956), .ZN(n8964) );
  INV_X1 U10283 ( .A(n8958), .ZN(n9259) );
  AOI22_X1 U10284 ( .A1(n9264), .A2(n8971), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3084), .ZN(n8959) );
  OAI21_X1 U10285 ( .B1(n9080), .B2(n8960), .A(n8959), .ZN(n8961) );
  AOI21_X1 U10286 ( .B1(n9259), .B2(n8962), .A(n8961), .ZN(n8963) );
  OAI211_X1 U10287 ( .C1(n9261), .C2(n8996), .A(n8964), .B(n8963), .ZN(
        P1_U3231) );
  INV_X1 U10288 ( .A(n8965), .ZN(n8970) );
  AOI21_X1 U10289 ( .B1(n8967), .B2(n8969), .A(n8966), .ZN(n8968) );
  AOI21_X1 U10290 ( .B1(n8970), .B2(n8969), .A(n8968), .ZN(n8976) );
  AOI22_X1 U10291 ( .A1(n9198), .A2(n8971), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3084), .ZN(n8973) );
  NAND2_X1 U10292 ( .A1(n9264), .A2(n8983), .ZN(n8972) );
  OAI211_X1 U10293 ( .C1(n9005), .C2(n9228), .A(n8973), .B(n8972), .ZN(n8974)
         );
  AOI21_X1 U10294 ( .B1(n9432), .B2(n9007), .A(n8974), .ZN(n8975) );
  OAI21_X1 U10295 ( .B1(n8976), .B2(n9009), .A(n8975), .ZN(P1_U3233) );
  NAND2_X1 U10296 ( .A1(n8977), .A2(n8978), .ZN(n8980) );
  XNOR2_X1 U10297 ( .A(n8980), .B(n8979), .ZN(n8987) );
  OAI22_X1 U10298 ( .A1(n8981), .A2(n9080), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10108), .ZN(n8982) );
  AOI21_X1 U10299 ( .B1(n8983), .B2(n9314), .A(n8982), .ZN(n8984) );
  OAI21_X1 U10300 ( .B1(n9005), .B2(n9283), .A(n8984), .ZN(n8985) );
  AOI21_X1 U10301 ( .B1(n9452), .B2(n9007), .A(n8985), .ZN(n8986) );
  OAI21_X1 U10302 ( .B1(n8987), .B2(n9009), .A(n8986), .ZN(P1_U3236) );
  AOI211_X1 U10303 ( .C1(n8990), .C2(n8989), .A(n9009), .B(n8988), .ZN(n8991)
         );
  INV_X1 U10304 ( .A(n8991), .ZN(n8995) );
  OAI22_X1 U10305 ( .A1(n9095), .A2(n9238), .B1(n9092), .B2(n9236), .ZN(n9173)
         );
  OAI22_X1 U10306 ( .A1(n9177), .A2(n9005), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8992), .ZN(n8993) );
  AOI21_X1 U10307 ( .B1(n9173), .B2(n9003), .A(n8993), .ZN(n8994) );
  OAI211_X1 U10308 ( .C1(n9094), .C2(n8996), .A(n8995), .B(n8994), .ZN(
        P1_U3238) );
  NAND2_X1 U10309 ( .A1(n8998), .A2(n8997), .ZN(n8999) );
  XOR2_X1 U10310 ( .A(n9000), .B(n8999), .Z(n9010) );
  OR2_X1 U10311 ( .A1(n9012), .A2(n9238), .ZN(n9002) );
  NAND2_X1 U10312 ( .A1(n9073), .A2(n9368), .ZN(n9001) );
  NAND2_X1 U10313 ( .A1(n9002), .A2(n9001), .ZN(n9333) );
  AOI22_X1 U10314 ( .A1(n9333), .A2(n9003), .B1(P1_REG3_REG_15__SCAN_IN), .B2(
        P1_U3084), .ZN(n9004) );
  OAI21_X1 U10315 ( .B1(n9005), .B2(n9336), .A(n9004), .ZN(n9006) );
  AOI21_X1 U10316 ( .B1(n9925), .B2(n9007), .A(n9006), .ZN(n9008) );
  OAI21_X1 U10317 ( .B1(n9010), .B2(n9009), .A(n9008), .ZN(P1_U3239) );
  MUX2_X1 U10318 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9129), .S(n9022), .Z(
        P1_U3585) );
  MUX2_X1 U10319 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9151), .S(n9022), .Z(
        P1_U3584) );
  MUX2_X1 U10320 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9097), .S(n9022), .Z(
        P1_U3583) );
  INV_X1 U10321 ( .A(n9095), .ZN(n9150) );
  MUX2_X1 U10322 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9150), .S(n9022), .Z(
        P1_U3582) );
  MUX2_X1 U10323 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9165), .S(n9022), .Z(
        P1_U3581) );
  INV_X1 U10324 ( .A(n9092), .ZN(n9199) );
  MUX2_X1 U10325 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9199), .S(n9022), .Z(
        P1_U3580) );
  MUX2_X1 U10326 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9091), .S(n9022), .Z(
        P1_U3579) );
  MUX2_X1 U10327 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9198), .S(n9022), .Z(
        P1_U3578) );
  MUX2_X1 U10328 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9083), .S(n9022), .Z(
        P1_U3577) );
  MUX2_X1 U10329 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9264), .S(n9022), .Z(
        P1_U3576) );
  MUX2_X1 U10330 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9276), .S(n9022), .Z(
        P1_U3575) );
  MUX2_X1 U10331 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9290), .S(n9022), .Z(
        P1_U3574) );
  INV_X1 U10332 ( .A(n9011), .ZN(n9275) );
  MUX2_X1 U10333 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9275), .S(n9022), .Z(
        P1_U3573) );
  MUX2_X1 U10334 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9314), .S(n9022), .Z(
        P1_U3572) );
  INV_X1 U10335 ( .A(n9012), .ZN(n9076) );
  MUX2_X1 U10336 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9076), .S(n9022), .Z(
        P1_U3571) );
  MUX2_X1 U10337 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9313), .S(P1_U4006), .Z(
        P1_U3570) );
  MUX2_X1 U10338 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9073), .S(P1_U4006), .Z(
        P1_U3569) );
  MUX2_X1 U10339 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9070), .S(P1_U4006), .Z(
        P1_U3568) );
  MUX2_X1 U10340 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9013), .S(P1_U4006), .Z(
        P1_U3567) );
  MUX2_X1 U10341 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9014), .S(P1_U4006), .Z(
        P1_U3566) );
  MUX2_X1 U10342 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9015), .S(P1_U4006), .Z(
        P1_U3565) );
  MUX2_X1 U10343 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9016), .S(P1_U4006), .Z(
        P1_U3564) );
  MUX2_X1 U10344 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9017), .S(P1_U4006), .Z(
        P1_U3563) );
  MUX2_X1 U10345 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9018), .S(P1_U4006), .Z(
        P1_U3562) );
  MUX2_X1 U10346 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9371), .S(P1_U4006), .Z(
        P1_U3561) );
  MUX2_X1 U10347 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9019), .S(P1_U4006), .Z(
        P1_U3560) );
  MUX2_X1 U10348 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9369), .S(P1_U4006), .Z(
        P1_U3559) );
  MUX2_X1 U10349 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9020), .S(P1_U4006), .Z(
        P1_U3558) );
  MUX2_X1 U10350 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n9021), .S(P1_U4006), .Z(
        P1_U3557) );
  MUX2_X1 U10351 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n6552), .S(P1_U4006), .Z(
        P1_U3556) );
  MUX2_X1 U10352 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n6027), .S(n9022), .Z(
        P1_U3555) );
  NAND2_X1 U10353 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n10038), .ZN(n9023) );
  OAI21_X1 U10354 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n10038), .A(n9023), .ZN(
        n10041) );
  AOI22_X1 U10355 ( .A1(P1_REG2_REG_11__SCAN_IN), .A2(n10026), .B1(n9037), 
        .B2(n7897), .ZN(n10028) );
  OAI21_X1 U10356 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n10026), .A(n10027), 
        .ZN(n10040) );
  NOR2_X1 U10357 ( .A1(n10041), .A2(n10040), .ZN(n10039) );
  AOI21_X1 U10358 ( .B1(n10038), .B2(P1_REG2_REG_12__SCAN_IN), .A(n10039), 
        .ZN(n10051) );
  NAND2_X1 U10359 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n9039), .ZN(n9026) );
  OAI21_X1 U10360 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n9039), .A(n9026), .ZN(
        n10050) );
  NOR2_X1 U10361 ( .A1(n10051), .A2(n10050), .ZN(n10049) );
  NOR2_X1 U10362 ( .A1(n9027), .A2(n9040), .ZN(n9028) );
  NOR2_X1 U10363 ( .A1(n9030), .A2(n9029), .ZN(n9031) );
  XOR2_X1 U10364 ( .A(n10077), .B(n9030), .Z(n10074) );
  NOR2_X1 U10365 ( .A1(n9337), .A2(n10074), .ZN(n10073) );
  NOR2_X1 U10366 ( .A1(n9031), .A2(n10073), .ZN(n10086) );
  NAND2_X1 U10367 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n10089), .ZN(n9032) );
  OAI21_X1 U10368 ( .B1(P1_REG2_REG_16__SCAN_IN), .B2(n10089), .A(n9032), .ZN(
        n10085) );
  NAND2_X1 U10369 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(n10101), .ZN(n9033) );
  OAI21_X1 U10370 ( .B1(P1_REG2_REG_17__SCAN_IN), .B2(n10101), .A(n9033), .ZN(
        n10097) );
  AOI22_X1 U10371 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n9047), .B1(n10115), 
        .B2(n5996), .ZN(n10111) );
  NOR2_X1 U10372 ( .A1(n10112), .A2(n10111), .ZN(n10110) );
  AOI21_X1 U10373 ( .B1(n10115), .B2(P1_REG2_REG_18__SCAN_IN), .A(n10110), 
        .ZN(n9034) );
  XNOR2_X1 U10374 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n9034), .ZN(n9056) );
  AOI22_X1 U10375 ( .A1(P1_REG1_REG_18__SCAN_IN), .A2(n9047), .B1(n10115), 
        .B2(n9046), .ZN(n10118) );
  AOI22_X1 U10376 ( .A1(P1_REG1_REG_17__SCAN_IN), .A2(n10101), .B1(n9045), 
        .B2(n9044), .ZN(n10104) );
  AOI22_X1 U10377 ( .A1(P1_REG1_REG_16__SCAN_IN), .A2(n10089), .B1(n9043), 
        .B2(n6232), .ZN(n10092) );
  AOI22_X1 U10378 ( .A1(P1_REG1_REG_11__SCAN_IN), .A2(n9037), .B1(n10026), 
        .B2(n6156), .ZN(n10022) );
  NOR2_X1 U10379 ( .A1(n10023), .A2(n10022), .ZN(n10021) );
  AOI22_X1 U10380 ( .A1(P1_REG1_REG_12__SCAN_IN), .A2(n9038), .B1(n10038), 
        .B2(n6123), .ZN(n10035) );
  NOR2_X1 U10381 ( .A1(n10036), .A2(n10035), .ZN(n10034) );
  AOI22_X1 U10382 ( .A1(P1_REG1_REG_13__SCAN_IN), .A2(n10053), .B1(n9039), 
        .B2(n6189), .ZN(n10047) );
  NOR2_X1 U10383 ( .A1(n10048), .A2(n10047), .ZN(n10046) );
  AOI22_X1 U10384 ( .A1(n10064), .A2(n6175), .B1(P1_REG1_REG_14__SCAN_IN), 
        .B2(n9040), .ZN(n10060) );
  NOR2_X1 U10385 ( .A1(n10061), .A2(n10060), .ZN(n10059) );
  NAND2_X1 U10386 ( .A1(n10077), .A2(n9041), .ZN(n9042) );
  XOR2_X1 U10387 ( .A(n10077), .B(n9041), .Z(n10079) );
  NAND2_X1 U10388 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n10079), .ZN(n10078) );
  NAND2_X1 U10389 ( .A1(n9042), .A2(n10078), .ZN(n10091) );
  NAND2_X1 U10390 ( .A1(n10092), .A2(n10091), .ZN(n10090) );
  OAI21_X1 U10391 ( .B1(n9045), .B2(n9044), .A(n10102), .ZN(n10119) );
  NOR2_X1 U10392 ( .A1(n10118), .A2(n10119), .ZN(n10120) );
  XOR2_X1 U10393 ( .A(n9049), .B(n9048), .Z(n9053) );
  INV_X1 U10394 ( .A(n9053), .ZN(n9050) );
  AOI22_X1 U10395 ( .A1(n9056), .A2(n10030), .B1(n10117), .B2(n9050), .ZN(
        n9051) );
  INV_X1 U10396 ( .A(n9052), .ZN(n9055) );
  AOI21_X1 U10397 ( .B1(n9053), .B2(n10117), .A(n10116), .ZN(n9054) );
  INV_X1 U10398 ( .A(n9064), .ZN(n9392) );
  NAND2_X1 U10399 ( .A1(n9269), .A2(n9261), .ZN(n9256) );
  XNOR2_X1 U10400 ( .A(n9388), .B(n9058), .ZN(n9386) );
  NAND2_X1 U10401 ( .A1(n9386), .A2(n9294), .ZN(n9063) );
  NAND2_X1 U10402 ( .A1(n9059), .A2(P1_B_REG_SCAN_IN), .ZN(n9060) );
  AND2_X1 U10403 ( .A1(n9370), .A2(n9060), .ZN(n9130) );
  NAND2_X1 U10404 ( .A1(n9061), .A2(n9130), .ZN(n9390) );
  NOR2_X1 U10405 ( .A1(n9390), .A2(n9353), .ZN(n9065) );
  AOI21_X1 U10406 ( .B1(n9242), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9065), .ZN(
        n9062) );
  OAI211_X1 U10407 ( .C1(n9388), .C2(n10145), .A(n9063), .B(n9062), .ZN(
        P1_U3261) );
  XNOR2_X1 U10408 ( .A(n9064), .B(n9133), .ZN(n9389) );
  NAND2_X1 U10409 ( .A1(n9389), .A2(n9294), .ZN(n9067) );
  AOI21_X1 U10410 ( .B1(n9353), .B2(P1_REG2_REG_30__SCAN_IN), .A(n9065), .ZN(
        n9066) );
  OAI211_X1 U10411 ( .C1(n9392), .C2(n10145), .A(n9067), .B(n9066), .ZN(
        P1_U3262) );
  OR2_X1 U10412 ( .A1(n9932), .A2(n9070), .ZN(n9068) );
  NAND2_X1 U10413 ( .A1(n9069), .A2(n9068), .ZN(n9072) );
  NAND2_X1 U10414 ( .A1(n9932), .A2(n9070), .ZN(n9071) );
  AND2_X1 U10415 ( .A1(n9463), .A2(n9073), .ZN(n9075) );
  OR2_X1 U10416 ( .A1(n9463), .A2(n9073), .ZN(n9074) );
  NOR2_X1 U10417 ( .A1(n9318), .A2(n9317), .ZN(n9316) );
  NOR2_X1 U10418 ( .A1(n9316), .A2(n9077), .ZN(n9296) );
  NOR2_X1 U10419 ( .A1(n9458), .A2(n9314), .ZN(n9079) );
  AOI22_X2 U10420 ( .A1(n9241), .A2(n9244), .B1(n9439), .B2(n9264), .ZN(n9224)
         );
  NAND2_X1 U10421 ( .A1(n9432), .A2(n9083), .ZN(n9085) );
  AOI22_X2 U10422 ( .A1(n9224), .A2(n9085), .B1(n9226), .B2(n9084), .ZN(n9209)
         );
  NAND2_X1 U10423 ( .A1(n9086), .A2(n9237), .ZN(n9087) );
  NAND2_X1 U10424 ( .A1(n9209), .A2(n9087), .ZN(n9088) );
  NAND2_X1 U10425 ( .A1(n9142), .A2(n9148), .ZN(n9141) );
  INV_X1 U10426 ( .A(n9400), .ZN(n9147) );
  NAND2_X1 U10427 ( .A1(n9400), .A2(n9097), .ZN(n9098) );
  NAND2_X1 U10428 ( .A1(n9141), .A2(n9098), .ZN(n9100) );
  XNOR2_X1 U10429 ( .A(n9100), .B(n9099), .ZN(n9393) );
  INV_X1 U10430 ( .A(n9393), .ZN(n9140) );
  NAND2_X1 U10431 ( .A1(n9332), .A2(n9105), .ZN(n9311) );
  INV_X1 U10432 ( .A(n9106), .ZN(n9107) );
  NAND2_X1 U10433 ( .A1(n9303), .A2(n9109), .ZN(n9287) );
  INV_X1 U10434 ( .A(n9110), .ZN(n9111) );
  INV_X1 U10435 ( .A(n9117), .ZN(n9213) );
  NOR3_X2 U10436 ( .A1(n9231), .A2(n9213), .A3(n9212), .ZN(n9211) );
  AOI21_X1 U10437 ( .B1(n9149), .B2(n9126), .A(n9125), .ZN(n9128) );
  XNOR2_X1 U10438 ( .A(n9128), .B(n9127), .ZN(n9132) );
  AOI22_X1 U10439 ( .A1(n9097), .A2(n9368), .B1(n9130), .B2(n9129), .ZN(n9131)
         );
  AOI21_X1 U10440 ( .B1(n9134), .B2(n9143), .A(n9133), .ZN(n9397) );
  NAND2_X1 U10441 ( .A1(n9397), .A2(n9294), .ZN(n9137) );
  AOI22_X1 U10442 ( .A1(n9135), .A2(n10135), .B1(P1_REG2_REG_29__SCAN_IN), 
        .B2(n9242), .ZN(n9136) );
  OAI211_X1 U10443 ( .C1(n9394), .C2(n10145), .A(n9137), .B(n9136), .ZN(n9138)
         );
  AOI21_X1 U10444 ( .B1(n9395), .B2(n10143), .A(n9138), .ZN(n9139) );
  OAI21_X1 U10445 ( .B1(n9140), .B2(n9366), .A(n9139), .ZN(P1_U3355) );
  OAI21_X1 U10446 ( .B1(n9142), .B2(n9148), .A(n9141), .ZN(n9404) );
  INV_X1 U10447 ( .A(n9143), .ZN(n9144) );
  AOI21_X1 U10448 ( .B1(n9400), .B2(n9157), .A(n9144), .ZN(n9401) );
  AOI22_X1 U10449 ( .A1(n9145), .A2(n10135), .B1(P1_REG2_REG_28__SCAN_IN), 
        .B2(n9242), .ZN(n9146) );
  OAI21_X1 U10450 ( .B1(n9147), .B2(n10145), .A(n9146), .ZN(n9154) );
  XNOR2_X1 U10451 ( .A(n9149), .B(n9148), .ZN(n9152) );
  AOI222_X1 U10452 ( .A1(n10133), .A2(n9152), .B1(n9151), .B2(n9370), .C1(
        n9150), .C2(n9368), .ZN(n9403) );
  NOR2_X1 U10453 ( .A1(n9403), .A2(n9242), .ZN(n9153) );
  AOI211_X1 U10454 ( .C1(n9401), .C2(n9294), .A(n9154), .B(n9153), .ZN(n9155)
         );
  OAI21_X1 U10455 ( .B1(n9366), .B2(n9404), .A(n9155), .ZN(P1_U3263) );
  XOR2_X1 U10456 ( .A(n9164), .B(n9156), .Z(n9409) );
  INV_X1 U10457 ( .A(n9175), .ZN(n9159) );
  INV_X1 U10458 ( .A(n9157), .ZN(n9158) );
  AOI21_X1 U10459 ( .B1(n9405), .B2(n9159), .A(n9158), .ZN(n9406) );
  AOI22_X1 U10460 ( .A1(n9160), .A2(n10135), .B1(P1_REG2_REG_27__SCAN_IN), 
        .B2(n9242), .ZN(n9161) );
  OAI21_X1 U10461 ( .B1(n9162), .B2(n10145), .A(n9161), .ZN(n9168) );
  XOR2_X1 U10462 ( .A(n9164), .B(n9163), .Z(n9166) );
  AOI222_X1 U10463 ( .A1(n10133), .A2(n9166), .B1(n9097), .B2(n9370), .C1(
        n9165), .C2(n9368), .ZN(n9408) );
  NOR2_X1 U10464 ( .A1(n9408), .A2(n9242), .ZN(n9167) );
  AOI211_X1 U10465 ( .C1(n9294), .C2(n9406), .A(n9168), .B(n9167), .ZN(n9169)
         );
  OAI21_X1 U10466 ( .B1(n9409), .B2(n9366), .A(n9169), .ZN(P1_U3264) );
  XOR2_X1 U10467 ( .A(n9172), .B(n9170), .Z(n9414) );
  AOI22_X1 U10468 ( .A1(n9411), .A2(n9343), .B1(n9353), .B2(
        P1_REG2_REG_26__SCAN_IN), .ZN(n9180) );
  XOR2_X1 U10469 ( .A(n9172), .B(n9171), .Z(n9174) );
  INV_X1 U10470 ( .A(n10125), .ZN(n10209) );
  AOI211_X1 U10471 ( .C1(n9411), .C2(n9182), .A(n10209), .B(n9175), .ZN(n9410)
         );
  NAND2_X1 U10472 ( .A1(n9410), .A2(n9203), .ZN(n9176) );
  OAI211_X1 U10473 ( .C1(n10151), .C2(n9177), .A(n9413), .B(n9176), .ZN(n9178)
         );
  NAND2_X1 U10474 ( .A1(n9178), .A2(n10143), .ZN(n9179) );
  OAI211_X1 U10475 ( .C1(n9414), .C2(n9366), .A(n9180), .B(n9179), .ZN(
        P1_U3265) );
  XOR2_X1 U10476 ( .A(n9188), .B(n9181), .Z(n9419) );
  AOI211_X1 U10477 ( .C1(n9416), .C2(n9201), .A(n10209), .B(n4753), .ZN(n9415)
         );
  INV_X1 U10478 ( .A(n9183), .ZN(n9184) );
  AOI22_X1 U10479 ( .A1(n9184), .A2(n10135), .B1(P1_REG2_REG_25__SCAN_IN), 
        .B2(n9242), .ZN(n9185) );
  OAI21_X1 U10480 ( .B1(n9186), .B2(n10145), .A(n9185), .ZN(n9192) );
  XOR2_X1 U10481 ( .A(n9188), .B(n9187), .Z(n9190) );
  NOR2_X1 U10482 ( .A1(n9418), .A2(n9242), .ZN(n9191) );
  AOI211_X1 U10483 ( .C1(n9415), .C2(n9364), .A(n9192), .B(n9191), .ZN(n9193)
         );
  OAI21_X1 U10484 ( .B1(n9419), .B2(n9366), .A(n9193), .ZN(P1_U3266) );
  XOR2_X1 U10485 ( .A(n9197), .B(n9194), .Z(n9424) );
  AOI22_X1 U10486 ( .A1(n9421), .A2(n9343), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n9242), .ZN(n9208) );
  OAI21_X1 U10487 ( .B1(n9197), .B2(n9196), .A(n9195), .ZN(n9200) );
  AOI222_X1 U10488 ( .A1(n10133), .A2(n9200), .B1(n9199), .B2(n9370), .C1(
        n9198), .C2(n9368), .ZN(n9423) );
  INV_X1 U10489 ( .A(n9219), .ZN(n9202) );
  AOI211_X1 U10490 ( .C1(n9421), .C2(n9202), .A(n10209), .B(n4754), .ZN(n9420)
         );
  NAND2_X1 U10491 ( .A1(n9420), .A2(n9203), .ZN(n9204) );
  OAI211_X1 U10492 ( .C1(n10151), .C2(n9205), .A(n9423), .B(n9204), .ZN(n9206)
         );
  NAND2_X1 U10493 ( .A1(n9206), .A2(n10143), .ZN(n9207) );
  OAI211_X1 U10494 ( .C1(n9424), .C2(n9366), .A(n9208), .B(n9207), .ZN(
        P1_U3267) );
  XNOR2_X1 U10495 ( .A(n9209), .B(n9212), .ZN(n9430) );
  INV_X1 U10496 ( .A(n9210), .ZN(n9217) );
  NOR2_X1 U10497 ( .A1(n9211), .A2(n9356), .ZN(n9216) );
  OAI21_X1 U10498 ( .B1(n9231), .B2(n9213), .A(n9212), .ZN(n9215) );
  AOI21_X1 U10499 ( .B1(n9216), .B2(n9215), .A(n9214), .ZN(n9429) );
  OAI21_X1 U10500 ( .B1(n9217), .B2(n10151), .A(n9429), .ZN(n9222) );
  NOR2_X1 U10501 ( .A1(n9225), .A2(n9086), .ZN(n9218) );
  OR2_X1 U10502 ( .A1(n9219), .A2(n9218), .ZN(n9425) );
  AOI22_X1 U10503 ( .A1(n9426), .A2(n9343), .B1(n9353), .B2(
        P1_REG2_REG_23__SCAN_IN), .ZN(n9220) );
  OAI21_X1 U10504 ( .B1(n9425), .B2(n10146), .A(n9220), .ZN(n9221) );
  AOI21_X1 U10505 ( .B1(n9222), .B2(n10143), .A(n9221), .ZN(n9223) );
  OAI21_X1 U10506 ( .B1(n9430), .B2(n9366), .A(n9223), .ZN(P1_U3268) );
  XOR2_X1 U10507 ( .A(n9232), .B(n9224), .Z(n9436) );
  AOI21_X1 U10508 ( .B1(n9432), .B2(n9247), .A(n9225), .ZN(n9433) );
  NOR2_X1 U10509 ( .A1(n9226), .A2(n10145), .ZN(n9230) );
  OAI22_X1 U10510 ( .A1(n9228), .A2(n10151), .B1(n10143), .B2(n9227), .ZN(
        n9229) );
  AOI211_X1 U10511 ( .C1(n9433), .C2(n9294), .A(n9230), .B(n9229), .ZN(n9240)
         );
  AOI21_X1 U10512 ( .B1(n9233), .B2(n9232), .A(n9231), .ZN(n9234) );
  OAI222_X1 U10513 ( .A1(n9238), .A2(n9237), .B1(n9236), .B2(n9235), .C1(n9356), .C2(n9234), .ZN(n9431) );
  NAND2_X1 U10514 ( .A1(n9431), .A2(n10143), .ZN(n9239) );
  OAI211_X1 U10515 ( .C1(n9436), .C2(n9366), .A(n9240), .B(n9239), .ZN(
        P1_U3269) );
  XNOR2_X1 U10516 ( .A(n9241), .B(n9244), .ZN(n9441) );
  AOI22_X1 U10517 ( .A1(n9439), .A2(n9343), .B1(P1_REG2_REG_21__SCAN_IN), .B2(
        n9242), .ZN(n9254) );
  AOI21_X1 U10518 ( .B1(n9244), .B2(n9243), .A(n4529), .ZN(n9246) );
  OAI21_X1 U10519 ( .B1(n9246), .B2(n9356), .A(n9245), .ZN(n9437) );
  INV_X1 U10520 ( .A(n9247), .ZN(n9248) );
  AOI211_X1 U10521 ( .C1(n9439), .C2(n9256), .A(n10209), .B(n9248), .ZN(n9438)
         );
  INV_X1 U10522 ( .A(n9438), .ZN(n9251) );
  INV_X1 U10523 ( .A(n9249), .ZN(n9250) );
  OAI22_X1 U10524 ( .A1(n9251), .A2(n10138), .B1(n10151), .B2(n9250), .ZN(
        n9252) );
  OAI21_X1 U10525 ( .B1(n9437), .B2(n9252), .A(n10143), .ZN(n9253) );
  OAI211_X1 U10526 ( .C1(n9441), .C2(n9366), .A(n9254), .B(n9253), .ZN(
        P1_U3270) );
  XNOR2_X1 U10527 ( .A(n9255), .B(n9263), .ZN(n9446) );
  INV_X1 U10528 ( .A(n9269), .ZN(n9258) );
  INV_X1 U10529 ( .A(n9256), .ZN(n9257) );
  AOI21_X1 U10530 ( .B1(n9442), .B2(n9258), .A(n9257), .ZN(n9443) );
  AOI22_X1 U10531 ( .A1(n9353), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9259), .B2(
        n10135), .ZN(n9260) );
  OAI21_X1 U10532 ( .B1(n9261), .B2(n10145), .A(n9260), .ZN(n9267) );
  XOR2_X1 U10533 ( .A(n9263), .B(n9262), .Z(n9265) );
  AOI222_X1 U10534 ( .A1(n10133), .A2(n9265), .B1(n9264), .B2(n9370), .C1(
        n9290), .C2(n9368), .ZN(n9445) );
  NOR2_X1 U10535 ( .A1(n9445), .A2(n9242), .ZN(n9266) );
  AOI211_X1 U10536 ( .C1(n9443), .C2(n9294), .A(n9267), .B(n9266), .ZN(n9268)
         );
  OAI21_X1 U10537 ( .B1(n9446), .B2(n9366), .A(n9268), .ZN(P1_U3271) );
  XOR2_X1 U10538 ( .A(n4544), .B(n9273), .Z(n9451) );
  AOI21_X1 U10539 ( .B1(n9447), .B2(n4749), .A(n9269), .ZN(n9448) );
  AOI22_X1 U10540 ( .A1(n9353), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9270), .B2(
        n10135), .ZN(n9271) );
  OAI21_X1 U10541 ( .B1(n9272), .B2(n10145), .A(n9271), .ZN(n9279) );
  XNOR2_X1 U10542 ( .A(n9274), .B(n9273), .ZN(n9277) );
  AOI222_X1 U10543 ( .A1(n10133), .A2(n9277), .B1(n9276), .B2(n9370), .C1(
        n9275), .C2(n9368), .ZN(n9450) );
  NOR2_X1 U10544 ( .A1(n9450), .A2(n9242), .ZN(n9278) );
  AOI211_X1 U10545 ( .C1(n9448), .C2(n9294), .A(n9279), .B(n9278), .ZN(n9280)
         );
  OAI21_X1 U10546 ( .B1(n9451), .B2(n9366), .A(n9280), .ZN(P1_U3272) );
  XNOR2_X1 U10547 ( .A(n9281), .B(n9288), .ZN(n9456) );
  AOI21_X1 U10548 ( .B1(n9452), .B2(n9297), .A(n9282), .ZN(n9453) );
  INV_X1 U10549 ( .A(n9283), .ZN(n9284) );
  AOI22_X1 U10550 ( .A1(n9353), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9284), .B2(
        n10135), .ZN(n9285) );
  OAI21_X1 U10551 ( .B1(n4747), .B2(n10145), .A(n9285), .ZN(n9293) );
  NAND2_X1 U10552 ( .A1(n9287), .A2(n9286), .ZN(n9289) );
  XNOR2_X1 U10553 ( .A(n9289), .B(n9288), .ZN(n9291) );
  AOI222_X1 U10554 ( .A1(n10133), .A2(n9291), .B1(n9290), .B2(n9370), .C1(
        n9314), .C2(n9368), .ZN(n9455) );
  NOR2_X1 U10555 ( .A1(n9455), .A2(n9242), .ZN(n9292) );
  AOI211_X1 U10556 ( .C1(n9453), .C2(n9294), .A(n9293), .B(n9292), .ZN(n9295)
         );
  OAI21_X1 U10557 ( .B1(n9456), .B2(n9366), .A(n9295), .ZN(P1_U3273) );
  XNOR2_X1 U10558 ( .A(n9296), .B(n9304), .ZN(n9461) );
  INV_X1 U10559 ( .A(n9297), .ZN(n9298) );
  AOI211_X1 U10560 ( .C1(n9458), .C2(n9319), .A(n10209), .B(n9298), .ZN(n9457)
         );
  INV_X1 U10561 ( .A(n9299), .ZN(n9300) );
  AOI22_X1 U10562 ( .A1(n9353), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9300), .B2(
        n10135), .ZN(n9301) );
  OAI21_X1 U10563 ( .B1(n9302), .B2(n10145), .A(n9301), .ZN(n9308) );
  XOR2_X1 U10564 ( .A(n9304), .B(n9303), .Z(n9306) );
  AOI21_X1 U10565 ( .B1(n9306), .B2(n10133), .A(n9305), .ZN(n9460) );
  NOR2_X1 U10566 ( .A1(n9460), .A2(n9242), .ZN(n9307) );
  AOI211_X1 U10567 ( .C1(n9457), .C2(n9364), .A(n9308), .B(n9307), .ZN(n9309)
         );
  OAI21_X1 U10568 ( .B1(n9461), .B2(n9366), .A(n9309), .ZN(P1_U3274) );
  NAND2_X1 U10569 ( .A1(n9311), .A2(n9310), .ZN(n9312) );
  XOR2_X1 U10570 ( .A(n9317), .B(n9312), .Z(n9315) );
  AOI222_X1 U10571 ( .A1(n10133), .A2(n9315), .B1(n9314), .B2(n9370), .C1(
        n9313), .C2(n9368), .ZN(n9921) );
  AOI21_X1 U10572 ( .B1(n9318), .B2(n9317), .A(n9316), .ZN(n9924) );
  OAI211_X1 U10573 ( .C1(n9338), .C2(n9922), .A(n10125), .B(n9319), .ZN(n9920)
         );
  OAI22_X1 U10574 ( .A1(n10143), .A2(n9321), .B1(n9320), .B2(n10151), .ZN(
        n9322) );
  AOI21_X1 U10575 ( .B1(n9323), .B2(n9343), .A(n9322), .ZN(n9324) );
  OAI21_X1 U10576 ( .B1(n9920), .B2(n9325), .A(n9324), .ZN(n9326) );
  AOI21_X1 U10577 ( .B1(n9924), .B2(n9382), .A(n9326), .ZN(n9327) );
  OAI21_X1 U10578 ( .B1(n9242), .B2(n9921), .A(n9327), .ZN(P1_U3275) );
  AND2_X1 U10579 ( .A1(n9328), .A2(n9330), .ZN(n9329) );
  OR2_X1 U10580 ( .A1(n9329), .A2(n4567), .ZN(n9928) );
  INV_X1 U10581 ( .A(n9330), .ZN(n9331) );
  XNOR2_X1 U10582 ( .A(n9332), .B(n9331), .ZN(n9334) );
  AOI21_X1 U10583 ( .B1(n9334), .B2(n10133), .A(n9333), .ZN(n9335) );
  OAI21_X1 U10584 ( .B1(n9928), .B2(n10130), .A(n9335), .ZN(n9930) );
  NAND2_X1 U10585 ( .A1(n9930), .A2(n10143), .ZN(n9345) );
  OAI22_X1 U10586 ( .A1(n10143), .A2(n9337), .B1(n9336), .B2(n10151), .ZN(
        n9342) );
  INV_X1 U10587 ( .A(n9338), .ZN(n9340) );
  AOI21_X1 U10588 ( .B1(n9348), .B2(n9925), .A(n10209), .ZN(n9339) );
  NAND2_X1 U10589 ( .A1(n9340), .A2(n9339), .ZN(n9927) );
  NOR2_X1 U10590 ( .A1(n9927), .A2(n9325), .ZN(n9341) );
  AOI211_X1 U10591 ( .C1(n9343), .C2(n9925), .A(n9342), .B(n9341), .ZN(n9344)
         );
  OAI211_X1 U10592 ( .C1(n9928), .C2(n9346), .A(n9345), .B(n9344), .ZN(
        P1_U3276) );
  XNOR2_X1 U10593 ( .A(n9347), .B(n9357), .ZN(n9466) );
  AOI211_X1 U10594 ( .C1(n9463), .C2(n9350), .A(n10209), .B(n9349), .ZN(n9462)
         );
  INV_X1 U10595 ( .A(n9463), .ZN(n9355) );
  INV_X1 U10596 ( .A(n9351), .ZN(n9352) );
  AOI22_X1 U10597 ( .A1(n9353), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n9352), .B2(
        n10135), .ZN(n9354) );
  OAI21_X1 U10598 ( .B1(n9355), .B2(n10145), .A(n9354), .ZN(n9363) );
  AOI21_X1 U10599 ( .B1(n9358), .B2(n9357), .A(n9356), .ZN(n9361) );
  AOI21_X1 U10600 ( .B1(n9361), .B2(n9360), .A(n9359), .ZN(n9465) );
  NOR2_X1 U10601 ( .A1(n9465), .A2(n9242), .ZN(n9362) );
  AOI211_X1 U10602 ( .C1(n9364), .C2(n9462), .A(n9363), .B(n9362), .ZN(n9365)
         );
  OAI21_X1 U10603 ( .B1(n9366), .B2(n9466), .A(n9365), .ZN(P1_U3277) );
  XNOR2_X1 U10604 ( .A(n9367), .B(n9380), .ZN(n9372) );
  AOI222_X1 U10605 ( .A1(n10133), .A2(n9372), .B1(n9371), .B2(n9370), .C1(
        n9369), .C2(n9368), .ZN(n10182) );
  MUX2_X1 U10606 ( .A(n9373), .B(n10182), .S(n10143), .Z(n9385) );
  INV_X1 U10607 ( .A(n9374), .ZN(n9375) );
  AOI211_X1 U10608 ( .C1(n10176), .C2(n9376), .A(n10209), .B(n9375), .ZN(
        n10175) );
  OAI22_X1 U10609 ( .A1(n10145), .A2(n9378), .B1(n9377), .B2(n10151), .ZN(
        n9379) );
  AOI21_X1 U10610 ( .B1(n10175), .B2(n9364), .A(n9379), .ZN(n9384) );
  NAND2_X1 U10611 ( .A1(n9381), .A2(n9380), .ZN(n10178) );
  NAND3_X1 U10612 ( .A1(n10179), .A2(n10178), .A3(n9382), .ZN(n9383) );
  NAND3_X1 U10613 ( .A1(n9385), .A2(n9384), .A3(n9383), .ZN(P1_U3286) );
  NAND2_X1 U10614 ( .A1(n9386), .A2(n10125), .ZN(n9387) );
  OAI211_X1 U10615 ( .C1(n9388), .C2(n10207), .A(n9387), .B(n9390), .ZN(n9467)
         );
  MUX2_X1 U10616 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9467), .S(n10231), .Z(
        P1_U3554) );
  NAND2_X1 U10617 ( .A1(n9389), .A2(n10125), .ZN(n9391) );
  OAI211_X1 U10618 ( .C1(n9392), .C2(n10207), .A(n9391), .B(n9390), .ZN(n9468)
         );
  MUX2_X1 U10619 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n9468), .S(n10231), .Z(
        P1_U3553) );
  NAND2_X1 U10620 ( .A1(n9393), .A2(n10195), .ZN(n9399) );
  NOR2_X1 U10621 ( .A1(n9394), .A2(n10207), .ZN(n9396) );
  NAND2_X1 U10622 ( .A1(n9399), .A2(n9398), .ZN(n9469) );
  MUX2_X1 U10623 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9469), .S(n10231), .Z(
        P1_U3552) );
  AOI22_X1 U10624 ( .A1(n9401), .A2(n10125), .B1(n10177), .B2(n9400), .ZN(
        n9402) );
  OAI211_X1 U10625 ( .C1(n9404), .C2(n10197), .A(n9403), .B(n9402), .ZN(n9470)
         );
  MUX2_X1 U10626 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9470), .S(n10231), .Z(
        P1_U3551) );
  AOI22_X1 U10627 ( .A1(n9406), .A2(n10125), .B1(n10177), .B2(n9405), .ZN(
        n9407) );
  OAI211_X1 U10628 ( .C1(n9409), .C2(n10197), .A(n9408), .B(n9407), .ZN(n9471)
         );
  MUX2_X1 U10629 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9471), .S(n10231), .Z(
        P1_U3550) );
  AOI21_X1 U10630 ( .B1(n10177), .B2(n9411), .A(n9410), .ZN(n9412) );
  OAI211_X1 U10631 ( .C1(n9414), .C2(n10197), .A(n9413), .B(n9412), .ZN(n9472)
         );
  MUX2_X1 U10632 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9472), .S(n10231), .Z(
        P1_U3549) );
  AOI21_X1 U10633 ( .B1(n10177), .B2(n9416), .A(n9415), .ZN(n9417) );
  OAI211_X1 U10634 ( .C1(n9419), .C2(n10197), .A(n9418), .B(n9417), .ZN(n9473)
         );
  MUX2_X1 U10635 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9473), .S(n10231), .Z(
        P1_U3548) );
  AOI21_X1 U10636 ( .B1(n10177), .B2(n9421), .A(n9420), .ZN(n9422) );
  OAI211_X1 U10637 ( .C1(n9424), .C2(n10197), .A(n9423), .B(n9422), .ZN(n9474)
         );
  MUX2_X1 U10638 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9474), .S(n10231), .Z(
        P1_U3547) );
  INV_X1 U10639 ( .A(n9425), .ZN(n9427) );
  AOI22_X1 U10640 ( .A1(n9427), .A2(n10125), .B1(n10177), .B2(n9426), .ZN(
        n9428) );
  OAI211_X1 U10641 ( .C1(n9430), .C2(n10197), .A(n9429), .B(n9428), .ZN(n9475)
         );
  MUX2_X1 U10642 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9475), .S(n10231), .Z(
        P1_U3546) );
  INV_X1 U10643 ( .A(n9431), .ZN(n9435) );
  AOI22_X1 U10644 ( .A1(n9433), .A2(n10125), .B1(n10177), .B2(n9432), .ZN(
        n9434) );
  OAI211_X1 U10645 ( .C1(n9436), .C2(n10197), .A(n9435), .B(n9434), .ZN(n9476)
         );
  MUX2_X1 U10646 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9476), .S(n10231), .Z(
        P1_U3545) );
  AOI211_X1 U10647 ( .C1(n10177), .C2(n9439), .A(n9438), .B(n9437), .ZN(n9440)
         );
  OAI21_X1 U10648 ( .B1(n9441), .B2(n10197), .A(n9440), .ZN(n9477) );
  MUX2_X1 U10649 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9477), .S(n10231), .Z(
        P1_U3544) );
  AOI22_X1 U10650 ( .A1(n9443), .A2(n10125), .B1(n10177), .B2(n9442), .ZN(
        n9444) );
  OAI211_X1 U10651 ( .C1(n9446), .C2(n10197), .A(n9445), .B(n9444), .ZN(n9478)
         );
  MUX2_X1 U10652 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9478), .S(n10231), .Z(
        P1_U3543) );
  AOI22_X1 U10653 ( .A1(n9448), .A2(n10125), .B1(n10177), .B2(n9447), .ZN(
        n9449) );
  OAI211_X1 U10654 ( .C1(n9451), .C2(n10197), .A(n9450), .B(n9449), .ZN(n9479)
         );
  MUX2_X1 U10655 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9479), .S(n10231), .Z(
        P1_U3542) );
  AOI22_X1 U10656 ( .A1(n9453), .A2(n10125), .B1(n10177), .B2(n9452), .ZN(
        n9454) );
  OAI211_X1 U10657 ( .C1(n9456), .C2(n10197), .A(n9455), .B(n9454), .ZN(n9480)
         );
  MUX2_X1 U10658 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9480), .S(n10231), .Z(
        P1_U3541) );
  AOI21_X1 U10659 ( .B1(n10177), .B2(n9458), .A(n9457), .ZN(n9459) );
  OAI211_X1 U10660 ( .C1(n9461), .C2(n10197), .A(n9460), .B(n9459), .ZN(n9481)
         );
  MUX2_X1 U10661 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9481), .S(n10231), .Z(
        P1_U3540) );
  AOI21_X1 U10662 ( .B1(n10177), .B2(n9463), .A(n9462), .ZN(n9464) );
  OAI211_X1 U10663 ( .C1(n9466), .C2(n10197), .A(n9465), .B(n9464), .ZN(n9482)
         );
  MUX2_X1 U10664 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9482), .S(n10231), .Z(
        P1_U3537) );
  MUX2_X1 U10665 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9467), .S(n10217), .Z(
        P1_U3522) );
  MUX2_X1 U10666 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n9468), .S(n10217), .Z(
        P1_U3521) );
  MUX2_X1 U10667 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9469), .S(n10217), .Z(
        P1_U3520) );
  MUX2_X1 U10668 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9470), .S(n10217), .Z(
        P1_U3519) );
  MUX2_X1 U10669 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9471), .S(n10217), .Z(
        P1_U3518) );
  MUX2_X1 U10670 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9472), .S(n10217), .Z(
        P1_U3517) );
  MUX2_X1 U10671 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9473), .S(n10217), .Z(
        P1_U3516) );
  MUX2_X1 U10672 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9474), .S(n10217), .Z(
        P1_U3515) );
  MUX2_X1 U10673 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9475), .S(n10217), .Z(
        P1_U3514) );
  MUX2_X1 U10674 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9476), .S(n10217), .Z(
        P1_U3513) );
  MUX2_X1 U10675 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9477), .S(n10217), .Z(
        P1_U3512) );
  MUX2_X1 U10676 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9478), .S(n10217), .Z(
        P1_U3511) );
  MUX2_X1 U10677 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9479), .S(n10217), .Z(
        P1_U3510) );
  MUX2_X1 U10678 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9480), .S(n10217), .Z(
        P1_U3508) );
  MUX2_X1 U10679 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9481), .S(n10217), .Z(
        P1_U3505) );
  MUX2_X1 U10680 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n9482), .S(n10217), .Z(
        P1_U3496) );
  NOR4_X1 U10681 ( .A1(n9483), .A2(P1_IR_REG_30__SCAN_IN), .A3(n5913), .A4(
        P1_U3084), .ZN(n9484) );
  AOI21_X1 U10682 ( .B1(n9485), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9484), .ZN(
        n9486) );
  OAI21_X1 U10683 ( .B1(n9488), .B2(n9487), .A(n9486), .ZN(P1_U3322) );
  OAI222_X1 U10684 ( .A1(n9492), .A2(n9491), .B1(P1_U3084), .B2(n9490), .C1(
        n9598), .C2(n9489), .ZN(P1_U3324) );
  MUX2_X1 U10685 ( .A(n9493), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  INV_X1 U10686 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10400) );
  NOR2_X1 U10687 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n9494) );
  AOI21_X1 U10688 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n9494), .ZN(n10367) );
  NOR2_X1 U10689 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n9495) );
  AOI21_X1 U10690 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n9495), .ZN(n10370) );
  NOR2_X1 U10691 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n9496) );
  AOI21_X1 U10692 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n9496), .ZN(n10373) );
  NOR2_X1 U10693 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n9497) );
  AOI21_X1 U10694 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n9497), .ZN(n10376) );
  NOR2_X1 U10695 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n9498) );
  AOI21_X1 U10696 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n9498), .ZN(n10379) );
  NOR2_X1 U10697 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n9505) );
  XNOR2_X1 U10698 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10407) );
  NAND2_X1 U10699 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n9503) );
  XOR2_X1 U10700 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10405) );
  NAND2_X1 U10701 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n9501) );
  XOR2_X1 U10702 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(P1_ADDR_REG_2__SCAN_IN), .Z(
        n10394) );
  AOI21_X1 U10703 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10361) );
  NAND3_X1 U10704 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n10363) );
  OAI21_X1 U10705 ( .B1(n10361), .B2(n9499), .A(n10363), .ZN(n10393) );
  NAND2_X1 U10706 ( .A1(n10394), .A2(n10393), .ZN(n9500) );
  NAND2_X1 U10707 ( .A1(n9501), .A2(n9500), .ZN(n10404) );
  NAND2_X1 U10708 ( .A1(n10405), .A2(n10404), .ZN(n9502) );
  NAND2_X1 U10709 ( .A1(n9503), .A2(n9502), .ZN(n10406) );
  NOR2_X1 U10710 ( .A1(n10407), .A2(n10406), .ZN(n9504) );
  NOR2_X1 U10711 ( .A1(n9505), .A2(n9504), .ZN(n9506) );
  NOR2_X1 U10712 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n9506), .ZN(n10396) );
  AND2_X1 U10713 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n9506), .ZN(n10395) );
  NOR2_X1 U10714 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10395), .ZN(n9507) );
  NOR2_X1 U10715 ( .A1(n10396), .A2(n9507), .ZN(n9508) );
  NAND2_X1 U10716 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(n9508), .ZN(n9510) );
  XOR2_X1 U10717 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(n9508), .Z(n10403) );
  NAND2_X1 U10718 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(n10403), .ZN(n9509) );
  NAND2_X1 U10719 ( .A1(n9510), .A2(n9509), .ZN(n9511) );
  NAND2_X1 U10720 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n9511), .ZN(n9513) );
  XOR2_X1 U10721 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n9511), .Z(n10392) );
  NAND2_X1 U10722 ( .A1(n10392), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n9512) );
  NAND2_X1 U10723 ( .A1(n9513), .A2(n9512), .ZN(n9514) );
  NAND2_X1 U10724 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n9514), .ZN(n9516) );
  XOR2_X1 U10725 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n9514), .Z(n10402) );
  NAND2_X1 U10726 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10402), .ZN(n9515) );
  NAND2_X1 U10727 ( .A1(n9516), .A2(n9515), .ZN(n9517) );
  AND2_X1 U10728 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n9517), .ZN(n9518) );
  XNOR2_X1 U10729 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n9517), .ZN(n10391) );
  INV_X1 U10730 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10390) );
  NOR2_X1 U10731 ( .A1(n10391), .A2(n10390), .ZN(n10389) );
  NOR2_X1 U10732 ( .A1(n9518), .A2(n10389), .ZN(n10388) );
  NAND2_X1 U10733 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n9519) );
  OAI21_X1 U10734 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n9519), .ZN(n10387) );
  NOR2_X1 U10735 ( .A1(n10388), .A2(n10387), .ZN(n10386) );
  AOI21_X1 U10736 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10386), .ZN(n10385) );
  NAND2_X1 U10737 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n9520) );
  OAI21_X1 U10738 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n9520), .ZN(n10384) );
  NOR2_X1 U10739 ( .A1(n10385), .A2(n10384), .ZN(n10383) );
  AOI21_X1 U10740 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10383), .ZN(n10382) );
  NOR2_X1 U10741 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n9521) );
  AOI21_X1 U10742 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n9521), .ZN(n10381) );
  NAND2_X1 U10743 ( .A1(n10382), .A2(n10381), .ZN(n10380) );
  OAI21_X1 U10744 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10380), .ZN(n10378) );
  NAND2_X1 U10745 ( .A1(n10379), .A2(n10378), .ZN(n10377) );
  OAI21_X1 U10746 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10377), .ZN(n10375) );
  NAND2_X1 U10747 ( .A1(n10376), .A2(n10375), .ZN(n10374) );
  OAI21_X1 U10748 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10374), .ZN(n10372) );
  NAND2_X1 U10749 ( .A1(n10373), .A2(n10372), .ZN(n10371) );
  OAI21_X1 U10750 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10371), .ZN(n10369) );
  NAND2_X1 U10751 ( .A1(n10370), .A2(n10369), .ZN(n10368) );
  OAI21_X1 U10752 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10368), .ZN(n10366) );
  NAND2_X1 U10753 ( .A1(n10367), .A2(n10366), .ZN(n10365) );
  OAI21_X1 U10754 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10365), .ZN(n10399) );
  NOR2_X1 U10755 ( .A1(n10400), .A2(n10399), .ZN(n9522) );
  NAND2_X1 U10756 ( .A1(n10400), .A2(n10399), .ZN(n10398) );
  OAI21_X1 U10757 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n9522), .A(n10398), .ZN(
        n9887) );
  INV_X1 U10758 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n9885) );
  XOR2_X1 U10759 ( .A(SI_20_), .B(keyinput_g12), .Z(n9529) );
  AOI22_X1 U10760 ( .A1(SI_17_), .A2(keyinput_g15), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(keyinput_g75), .ZN(n9523) );
  OAI221_X1 U10761 ( .B1(SI_17_), .B2(keyinput_g15), .C1(
        P2_DATAO_REG_21__SCAN_IN), .C2(keyinput_g75), .A(n9523), .ZN(n9528) );
  AOI22_X1 U10762 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(keyinput_g60), .B1(
        P1_IR_REG_9__SCAN_IN), .B2(keyinput_g100), .ZN(n9524) );
  OAI221_X1 U10763 ( .B1(P2_REG3_REG_18__SCAN_IN), .B2(keyinput_g60), .C1(
        P1_IR_REG_9__SCAN_IN), .C2(keyinput_g100), .A(n9524), .ZN(n9527) );
  AOI22_X1 U10764 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(keyinput_g68), .B1(
        P1_IR_REG_14__SCAN_IN), .B2(keyinput_g105), .ZN(n9525) );
  OAI221_X1 U10765 ( .B1(P2_DATAO_REG_28__SCAN_IN), .B2(keyinput_g68), .C1(
        P1_IR_REG_14__SCAN_IN), .C2(keyinput_g105), .A(n9525), .ZN(n9526) );
  NOR4_X1 U10766 ( .A1(n9529), .A2(n9528), .A3(n9527), .A4(n9526), .ZN(n9557)
         );
  AOI22_X1 U10767 ( .A1(SI_31_), .A2(keyinput_g1), .B1(P1_D_REG_4__SCAN_IN), 
        .B2(keyinput_g127), .ZN(n9530) );
  OAI221_X1 U10768 ( .B1(SI_31_), .B2(keyinput_g1), .C1(P1_D_REG_4__SCAN_IN), 
        .C2(keyinput_g127), .A(n9530), .ZN(n9537) );
  AOI22_X1 U10769 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(keyinput_g49), .B1(
        P1_IR_REG_17__SCAN_IN), .B2(keyinput_g108), .ZN(n9531) );
  OAI221_X1 U10770 ( .B1(P2_REG3_REG_5__SCAN_IN), .B2(keyinput_g49), .C1(
        P1_IR_REG_17__SCAN_IN), .C2(keyinput_g108), .A(n9531), .ZN(n9536) );
  AOI22_X1 U10771 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(keyinput_g35), .B1(SI_15_), .B2(keyinput_g17), .ZN(n9532) );
  OAI221_X1 U10772 ( .B1(P2_REG3_REG_7__SCAN_IN), .B2(keyinput_g35), .C1(
        SI_15_), .C2(keyinput_g17), .A(n9532), .ZN(n9535) );
  AOI22_X1 U10773 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(keyinput_g40), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(keyinput_g74), .ZN(n9533) );
  OAI221_X1 U10774 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(keyinput_g40), .C1(
        P2_DATAO_REG_22__SCAN_IN), .C2(keyinput_g74), .A(n9533), .ZN(n9534) );
  NOR4_X1 U10775 ( .A1(n9537), .A2(n9536), .A3(n9535), .A4(n9534), .ZN(n9556)
         );
  AOI22_X1 U10776 ( .A1(P1_D_REG_3__SCAN_IN), .A2(keyinput_g126), .B1(
        P1_IR_REG_25__SCAN_IN), .B2(keyinput_g116), .ZN(n9538) );
  OAI221_X1 U10777 ( .B1(P1_D_REG_3__SCAN_IN), .B2(keyinput_g126), .C1(
        P1_IR_REG_25__SCAN_IN), .C2(keyinput_g116), .A(n9538), .ZN(n9545) );
  AOI22_X1 U10778 ( .A1(P2_REG3_REG_20__SCAN_IN), .A2(keyinput_g55), .B1(
        P1_IR_REG_21__SCAN_IN), .B2(keyinput_g112), .ZN(n9539) );
  OAI221_X1 U10779 ( .B1(P2_REG3_REG_20__SCAN_IN), .B2(keyinput_g55), .C1(
        P1_IR_REG_21__SCAN_IN), .C2(keyinput_g112), .A(n9539), .ZN(n9544) );
  AOI22_X1 U10780 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(keyinput_g80), .B1(
        SI_22_), .B2(keyinput_g10), .ZN(n9540) );
  OAI221_X1 U10781 ( .B1(P2_DATAO_REG_16__SCAN_IN), .B2(keyinput_g80), .C1(
        SI_22_), .C2(keyinput_g10), .A(n9540), .ZN(n9543) );
  AOI22_X1 U10782 ( .A1(SI_30_), .A2(keyinput_g2), .B1(SI_19_), .B2(
        keyinput_g13), .ZN(n9541) );
  OAI221_X1 U10783 ( .B1(SI_30_), .B2(keyinput_g2), .C1(SI_19_), .C2(
        keyinput_g13), .A(n9541), .ZN(n9542) );
  NOR4_X1 U10784 ( .A1(n9545), .A2(n9544), .A3(n9543), .A4(n9542), .ZN(n9555)
         );
  AOI22_X1 U10785 ( .A1(SI_21_), .A2(keyinput_g11), .B1(P1_IR_REG_19__SCAN_IN), 
        .B2(keyinput_g110), .ZN(n9546) );
  OAI221_X1 U10786 ( .B1(SI_21_), .B2(keyinput_g11), .C1(P1_IR_REG_19__SCAN_IN), .C2(keyinput_g110), .A(n9546), .ZN(n9553) );
  AOI22_X1 U10787 ( .A1(SI_6_), .A2(keyinput_g26), .B1(P1_IR_REG_13__SCAN_IN), 
        .B2(keyinput_g104), .ZN(n9547) );
  OAI221_X1 U10788 ( .B1(SI_6_), .B2(keyinput_g26), .C1(P1_IR_REG_13__SCAN_IN), 
        .C2(keyinput_g104), .A(n9547), .ZN(n9552) );
  AOI22_X1 U10789 ( .A1(P2_REG3_REG_1__SCAN_IN), .A2(keyinput_g44), .B1(
        P1_IR_REG_31__SCAN_IN), .B2(keyinput_g122), .ZN(n9548) );
  OAI221_X1 U10790 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(keyinput_g44), .C1(
        P1_IR_REG_31__SCAN_IN), .C2(keyinput_g122), .A(n9548), .ZN(n9551) );
  AOI22_X1 U10791 ( .A1(P2_DATAO_REG_9__SCAN_IN), .A2(keyinput_g87), .B1(
        P1_IR_REG_24__SCAN_IN), .B2(keyinput_g115), .ZN(n9549) );
  OAI221_X1 U10792 ( .B1(P2_DATAO_REG_9__SCAN_IN), .B2(keyinput_g87), .C1(
        P1_IR_REG_24__SCAN_IN), .C2(keyinput_g115), .A(n9549), .ZN(n9550) );
  NOR4_X1 U10793 ( .A1(n9553), .A2(n9552), .A3(n9551), .A4(n9550), .ZN(n9554)
         );
  NAND4_X1 U10794 ( .A1(n9557), .A2(n9556), .A3(n9555), .A4(n9554), .ZN(n9695)
         );
  AOI22_X1 U10795 ( .A1(SI_29_), .A2(keyinput_g3), .B1(SI_3_), .B2(
        keyinput_g29), .ZN(n9558) );
  OAI221_X1 U10796 ( .B1(SI_29_), .B2(keyinput_g3), .C1(SI_3_), .C2(
        keyinput_g29), .A(n9558), .ZN(n9565) );
  AOI22_X1 U10797 ( .A1(SI_10_), .A2(keyinput_g22), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(keyinput_g85), .ZN(n9559) );
  OAI221_X1 U10798 ( .B1(SI_10_), .B2(keyinput_g22), .C1(
        P2_DATAO_REG_11__SCAN_IN), .C2(keyinput_g85), .A(n9559), .ZN(n9564) );
  AOI22_X1 U10799 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(keyinput_g39), .B1(
        P1_IR_REG_3__SCAN_IN), .B2(keyinput_g94), .ZN(n9560) );
  OAI221_X1 U10800 ( .B1(P2_REG3_REG_10__SCAN_IN), .B2(keyinput_g39), .C1(
        P1_IR_REG_3__SCAN_IN), .C2(keyinput_g94), .A(n9560), .ZN(n9563) );
  AOI22_X1 U10801 ( .A1(P2_DATAO_REG_13__SCAN_IN), .A2(keyinput_g83), .B1(
        P1_IR_REG_12__SCAN_IN), .B2(keyinput_g103), .ZN(n9561) );
  OAI221_X1 U10802 ( .B1(P2_DATAO_REG_13__SCAN_IN), .B2(keyinput_g83), .C1(
        P1_IR_REG_12__SCAN_IN), .C2(keyinput_g103), .A(n9561), .ZN(n9562) );
  NOR4_X1 U10803 ( .A1(n9565), .A2(n9564), .A3(n9563), .A4(n9562), .ZN(n9595)
         );
  AOI22_X1 U10804 ( .A1(P2_REG3_REG_21__SCAN_IN), .A2(keyinput_g45), .B1(
        P1_IR_REG_23__SCAN_IN), .B2(keyinput_g114), .ZN(n9566) );
  OAI221_X1 U10805 ( .B1(P2_REG3_REG_21__SCAN_IN), .B2(keyinput_g45), .C1(
        P1_IR_REG_23__SCAN_IN), .C2(keyinput_g114), .A(n9566), .ZN(n9573) );
  AOI22_X1 U10806 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(keyinput_g43), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(keyinput_g71), .ZN(n9567) );
  OAI221_X1 U10807 ( .B1(P2_REG3_REG_8__SCAN_IN), .B2(keyinput_g43), .C1(
        P2_DATAO_REG_25__SCAN_IN), .C2(keyinput_g71), .A(n9567), .ZN(n9572) );
  AOI22_X1 U10808 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(keyinput_g58), .B1(
        SI_13_), .B2(keyinput_g19), .ZN(n9568) );
  OAI221_X1 U10809 ( .B1(P2_REG3_REG_11__SCAN_IN), .B2(keyinput_g58), .C1(
        SI_13_), .C2(keyinput_g19), .A(n9568), .ZN(n9571) );
  AOI22_X1 U10810 ( .A1(P1_IR_REG_30__SCAN_IN), .A2(keyinput_g121), .B1(SI_25_), .B2(keyinput_g7), .ZN(n9569) );
  OAI221_X1 U10811 ( .B1(P1_IR_REG_30__SCAN_IN), .B2(keyinput_g121), .C1(
        SI_25_), .C2(keyinput_g7), .A(n9569), .ZN(n9570) );
  NOR4_X1 U10812 ( .A1(n9573), .A2(n9572), .A3(n9571), .A4(n9570), .ZN(n9594)
         );
  AOI22_X1 U10813 ( .A1(P2_REG3_REG_28__SCAN_IN), .A2(keyinput_g42), .B1(
        P1_IR_REG_8__SCAN_IN), .B2(keyinput_g99), .ZN(n9574) );
  OAI221_X1 U10814 ( .B1(P2_REG3_REG_28__SCAN_IN), .B2(keyinput_g42), .C1(
        P1_IR_REG_8__SCAN_IN), .C2(keyinput_g99), .A(n9574), .ZN(n9581) );
  AOI22_X1 U10815 ( .A1(P2_REG3_REG_2__SCAN_IN), .A2(keyinput_g59), .B1(SI_9_), 
        .B2(keyinput_g23), .ZN(n9575) );
  OAI221_X1 U10816 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(keyinput_g59), .C1(SI_9_), .C2(keyinput_g23), .A(n9575), .ZN(n9580) );
  AOI22_X1 U10817 ( .A1(SI_26_), .A2(keyinput_g6), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(keyinput_g69), .ZN(n9576) );
  OAI221_X1 U10818 ( .B1(SI_26_), .B2(keyinput_g6), .C1(
        P2_DATAO_REG_27__SCAN_IN), .C2(keyinput_g69), .A(n9576), .ZN(n9579) );
  AOI22_X1 U10819 ( .A1(SI_4_), .A2(keyinput_g28), .B1(P1_IR_REG_18__SCAN_IN), 
        .B2(keyinput_g109), .ZN(n9577) );
  OAI221_X1 U10820 ( .B1(SI_4_), .B2(keyinput_g28), .C1(P1_IR_REG_18__SCAN_IN), 
        .C2(keyinput_g109), .A(n9577), .ZN(n9578) );
  NOR4_X1 U10821 ( .A1(n9581), .A2(n9580), .A3(n9579), .A4(n9578), .ZN(n9593)
         );
  AOI22_X1 U10822 ( .A1(P2_RD_REG_SCAN_IN), .A2(keyinput_g33), .B1(
        P1_D_REG_2__SCAN_IN), .B2(keyinput_g125), .ZN(n9582) );
  OAI221_X1 U10823 ( .B1(P2_RD_REG_SCAN_IN), .B2(keyinput_g33), .C1(
        P1_D_REG_2__SCAN_IN), .C2(keyinput_g125), .A(n9582), .ZN(n9591) );
  AOI22_X1 U10824 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(keyinput_g50), .B1(n9584), .B2(keyinput_g81), .ZN(n9583) );
  OAI221_X1 U10825 ( .B1(P2_REG3_REG_17__SCAN_IN), .B2(keyinput_g50), .C1(
        n9584), .C2(keyinput_g81), .A(n9583), .ZN(n9590) );
  AOI22_X1 U10826 ( .A1(n9824), .A2(keyinput_g82), .B1(keyinput_g65), .B2(
        n5918), .ZN(n9585) );
  OAI221_X1 U10827 ( .B1(n9824), .B2(keyinput_g82), .C1(n5918), .C2(
        keyinput_g65), .A(n9585), .ZN(n9589) );
  AOI22_X1 U10828 ( .A1(n9792), .A2(keyinput_g57), .B1(n9587), .B2(keyinput_g9), .ZN(n9586) );
  OAI221_X1 U10829 ( .B1(n9792), .B2(keyinput_g57), .C1(n9587), .C2(
        keyinput_g9), .A(n9586), .ZN(n9588) );
  NOR4_X1 U10830 ( .A1(n9591), .A2(n9590), .A3(n9589), .A4(n9588), .ZN(n9592)
         );
  NAND4_X1 U10831 ( .A1(n9595), .A2(n9594), .A3(n9593), .A4(n9592), .ZN(n9694)
         );
  AOI22_X1 U10832 ( .A1(n5268), .A2(keyinput_g53), .B1(n9845), .B2(keyinput_g4), .ZN(n9596) );
  OAI221_X1 U10833 ( .B1(n5268), .B2(keyinput_g53), .C1(n9845), .C2(
        keyinput_g4), .A(n9596), .ZN(n9608) );
  AOI22_X1 U10834 ( .A1(n9599), .A2(keyinput_g54), .B1(keyinput_g67), .B2(
        n9598), .ZN(n9597) );
  OAI221_X1 U10835 ( .B1(n9599), .B2(keyinput_g54), .C1(n9598), .C2(
        keyinput_g67), .A(n9597), .ZN(n9607) );
  INV_X1 U10836 ( .A(SI_11_), .ZN(n9601) );
  AOI22_X1 U10837 ( .A1(n9601), .A2(keyinput_g21), .B1(keyinput_g48), .B2(
        n9860), .ZN(n9600) );
  OAI221_X1 U10838 ( .B1(n9601), .B2(keyinput_g21), .C1(n9860), .C2(
        keyinput_g48), .A(n9600), .ZN(n9606) );
  XOR2_X1 U10839 ( .A(n9602), .B(keyinput_g124), .Z(n9604) );
  XNOR2_X1 U10840 ( .A(P1_IR_REG_0__SCAN_IN), .B(keyinput_g91), .ZN(n9603) );
  NAND2_X1 U10841 ( .A1(n9604), .A2(n9603), .ZN(n9605) );
  NOR4_X1 U10842 ( .A1(n9608), .A2(n9607), .A3(n9606), .A4(n9605), .ZN(n9641)
         );
  AOI22_X1 U10843 ( .A1(n9610), .A2(keyinput_g61), .B1(n6090), .B2(
        keyinput_g97), .ZN(n9609) );
  OAI221_X1 U10844 ( .B1(n9610), .B2(keyinput_g61), .C1(n6090), .C2(
        keyinput_g97), .A(n9609), .ZN(n9618) );
  INV_X1 U10845 ( .A(SI_18_), .ZN(n9858) );
  AOI22_X1 U10846 ( .A1(n8270), .A2(keyinput_g47), .B1(n9858), .B2(
        keyinput_g14), .ZN(n9611) );
  OAI221_X1 U10847 ( .B1(n8270), .B2(keyinput_g47), .C1(n9858), .C2(
        keyinput_g14), .A(n9611), .ZN(n9617) );
  AOI22_X1 U10848 ( .A1(P2_U3152), .A2(keyinput_g34), .B1(n9779), .B2(
        keyinput_g72), .ZN(n9612) );
  OAI221_X1 U10849 ( .B1(P2_U3152), .B2(keyinput_g34), .C1(n9779), .C2(
        keyinput_g72), .A(n9612), .ZN(n9616) );
  XNOR2_X1 U10850 ( .A(P1_IR_REG_10__SCAN_IN), .B(keyinput_g101), .ZN(n9614)
         );
  XNOR2_X1 U10851 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(keyinput_g77), .ZN(n9613)
         );
  NAND2_X1 U10852 ( .A1(n9614), .A2(n9613), .ZN(n9615) );
  NOR4_X1 U10853 ( .A1(n9618), .A2(n9617), .A3(n9616), .A4(n9615), .ZN(n9640)
         );
  AOI22_X1 U10854 ( .A1(n8206), .A2(keyinput_g36), .B1(keyinput_g63), .B2(
        n8358), .ZN(n9619) );
  OAI221_X1 U10855 ( .B1(n8206), .B2(keyinput_g36), .C1(n8358), .C2(
        keyinput_g63), .A(n9619), .ZN(n9628) );
  AOI22_X1 U10856 ( .A1(n9621), .A2(keyinput_g52), .B1(n5915), .B2(
        keyinput_g118), .ZN(n9620) );
  OAI221_X1 U10857 ( .B1(n9621), .B2(keyinput_g52), .C1(n5915), .C2(
        keyinput_g118), .A(n9620), .ZN(n9627) );
  INV_X1 U10858 ( .A(P2_WR_REG_SCAN_IN), .ZN(n9770) );
  AOI22_X1 U10859 ( .A1(n9770), .A2(keyinput_g0), .B1(n9833), .B2(keyinput_g88), .ZN(n9622) );
  OAI221_X1 U10860 ( .B1(n9770), .B2(keyinput_g0), .C1(n9833), .C2(
        keyinput_g88), .A(n9622), .ZN(n9626) );
  XNOR2_X1 U10861 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput_g98), .ZN(n9624) );
  XNOR2_X1 U10862 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(keyinput_g78), .ZN(n9623)
         );
  NAND2_X1 U10863 ( .A1(n9624), .A2(n9623), .ZN(n9625) );
  NOR4_X1 U10864 ( .A1(n9628), .A2(n9627), .A3(n9626), .A4(n9625), .ZN(n9639)
         );
  AOI22_X1 U10865 ( .A1(n9839), .A2(keyinput_g37), .B1(n8214), .B2(
        keyinput_g38), .ZN(n9629) );
  OAI221_X1 U10866 ( .B1(n9839), .B2(keyinput_g37), .C1(n8214), .C2(
        keyinput_g38), .A(n9629), .ZN(n9637) );
  AOI22_X1 U10867 ( .A1(n7714), .A2(keyinput_g73), .B1(keyinput_g24), .B2(
        n9780), .ZN(n9630) );
  OAI221_X1 U10868 ( .B1(n7714), .B2(keyinput_g73), .C1(n9780), .C2(
        keyinput_g24), .A(n9630), .ZN(n9636) );
  XOR2_X1 U10869 ( .A(n5073), .B(keyinput_g111), .Z(n9634) );
  XNOR2_X1 U10870 ( .A(SI_2_), .B(keyinput_g30), .ZN(n9633) );
  XNOR2_X1 U10871 ( .A(P2_REG3_REG_24__SCAN_IN), .B(keyinput_g51), .ZN(n9632)
         );
  XNOR2_X1 U10872 ( .A(SI_1_), .B(keyinput_g31), .ZN(n9631) );
  NAND4_X1 U10873 ( .A1(n9634), .A2(n9633), .A3(n9632), .A4(n9631), .ZN(n9635)
         );
  NOR3_X1 U10874 ( .A1(n9637), .A2(n9636), .A3(n9635), .ZN(n9638) );
  NAND4_X1 U10875 ( .A1(n9641), .A2(n9640), .A3(n9639), .A4(n9638), .ZN(n9693)
         );
  AOI22_X1 U10876 ( .A1(n9865), .A2(keyinput_g5), .B1(keyinput_g76), .B2(n9793), .ZN(n9642) );
  OAI221_X1 U10877 ( .B1(n9865), .B2(keyinput_g5), .C1(n9793), .C2(
        keyinput_g76), .A(n9642), .ZN(n9653) );
  INV_X1 U10878 ( .A(SI_7_), .ZN(n9645) );
  AOI22_X1 U10879 ( .A1(n9645), .A2(keyinput_g25), .B1(n9644), .B2(
        keyinput_g20), .ZN(n9643) );
  OAI221_X1 U10880 ( .B1(n9645), .B2(keyinput_g25), .C1(n9644), .C2(
        keyinput_g20), .A(n9643), .ZN(n9652) );
  XOR2_X1 U10881 ( .A(n9646), .B(keyinput_g123), .Z(n9650) );
  XNOR2_X1 U10882 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput_g119), .ZN(n9649)
         );
  XNOR2_X1 U10883 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(keyinput_g84), .ZN(n9648)
         );
  XNOR2_X1 U10884 ( .A(P1_IR_REG_11__SCAN_IN), .B(keyinput_g102), .ZN(n9647)
         );
  NAND4_X1 U10885 ( .A1(n9650), .A2(n9649), .A3(n9648), .A4(n9647), .ZN(n9651)
         );
  NOR3_X1 U10886 ( .A1(n9653), .A2(n9652), .A3(n9651), .ZN(n9691) );
  AOI22_X1 U10887 ( .A1(n9655), .A2(keyinput_g64), .B1(keyinput_g66), .B2(
        n9807), .ZN(n9654) );
  OAI221_X1 U10888 ( .B1(n9655), .B2(keyinput_g64), .C1(n9807), .C2(
        keyinput_g66), .A(n9654), .ZN(n9665) );
  AOI22_X1 U10889 ( .A1(n9658), .A2(keyinput_g16), .B1(keyinput_g89), .B2(
        n9657), .ZN(n9656) );
  OAI221_X1 U10890 ( .B1(n9658), .B2(keyinput_g16), .C1(n9657), .C2(
        keyinput_g89), .A(n9656), .ZN(n9664) );
  XOR2_X1 U10891 ( .A(n5923), .B(keyinput_g120), .Z(n9662) );
  XOR2_X1 U10892 ( .A(n5563), .B(keyinput_g8), .Z(n9661) );
  XNOR2_X1 U10893 ( .A(P1_IR_REG_26__SCAN_IN), .B(keyinput_g117), .ZN(n9660)
         );
  XNOR2_X1 U10894 ( .A(P1_IR_REG_15__SCAN_IN), .B(keyinput_g106), .ZN(n9659)
         );
  NAND4_X1 U10895 ( .A1(n9662), .A2(n9661), .A3(n9660), .A4(n9659), .ZN(n9663)
         );
  NOR3_X1 U10896 ( .A1(n9665), .A2(n9664), .A3(n9663), .ZN(n9690) );
  AOI22_X1 U10897 ( .A1(n9667), .A2(keyinput_g18), .B1(n5898), .B2(
        keyinput_g93), .ZN(n9666) );
  OAI221_X1 U10898 ( .B1(n9667), .B2(keyinput_g18), .C1(n5898), .C2(
        keyinput_g93), .A(n9666), .ZN(n9676) );
  AOI22_X1 U10899 ( .A1(n5988), .A2(keyinput_g107), .B1(keyinput_g86), .B2(
        n9669), .ZN(n9668) );
  OAI221_X1 U10900 ( .B1(n5988), .B2(keyinput_g107), .C1(n9669), .C2(
        keyinput_g86), .A(n9668), .ZN(n9675) );
  XNOR2_X1 U10901 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(keyinput_g79), .ZN(n9673)
         );
  XNOR2_X1 U10902 ( .A(P1_IR_REG_22__SCAN_IN), .B(keyinput_g113), .ZN(n9672)
         );
  XNOR2_X1 U10903 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(keyinput_g90), .ZN(n9671)
         );
  XNOR2_X1 U10904 ( .A(SI_0_), .B(keyinput_g32), .ZN(n9670) );
  NAND4_X1 U10905 ( .A1(n9673), .A2(n9672), .A3(n9671), .A4(n9670), .ZN(n9674)
         );
  NOR3_X1 U10906 ( .A1(n9676), .A2(n9675), .A3(n9674), .ZN(n9689) );
  AOI22_X1 U10907 ( .A1(n5361), .A2(keyinput_g56), .B1(n5481), .B2(
        keyinput_g41), .ZN(n9677) );
  OAI221_X1 U10908 ( .B1(n5361), .B2(keyinput_g56), .C1(n5481), .C2(
        keyinput_g41), .A(n9677), .ZN(n9687) );
  AOI22_X1 U10909 ( .A1(n9821), .A2(keyinput_g46), .B1(n6060), .B2(
        keyinput_g95), .ZN(n9678) );
  OAI221_X1 U10910 ( .B1(n9821), .B2(keyinput_g46), .C1(n6060), .C2(
        keyinput_g95), .A(n9678), .ZN(n9686) );
  AOI22_X1 U10911 ( .A1(n9681), .A2(keyinput_g70), .B1(keyinput_g27), .B2(
        n9680), .ZN(n9679) );
  OAI221_X1 U10912 ( .B1(n9681), .B2(keyinput_g70), .C1(n9680), .C2(
        keyinput_g27), .A(n9679), .ZN(n9685) );
  XNOR2_X1 U10913 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput_g96), .ZN(n9683) );
  XNOR2_X1 U10914 ( .A(P2_REG3_REG_26__SCAN_IN), .B(keyinput_g62), .ZN(n9682)
         );
  NAND2_X1 U10915 ( .A1(n9683), .A2(n9682), .ZN(n9684) );
  NOR4_X1 U10916 ( .A1(n9687), .A2(n9686), .A3(n9685), .A4(n9684), .ZN(n9688)
         );
  NAND4_X1 U10917 ( .A1(n9691), .A2(n9690), .A3(n9689), .A4(n9688), .ZN(n9692)
         );
  NOR4_X1 U10918 ( .A1(n9695), .A2(n9694), .A3(n9693), .A4(n9692), .ZN(n9884)
         );
  OAI22_X1 U10919 ( .A1(SI_2_), .A2(keyinput_f30), .B1(keyinput_f1), .B2(
        SI_31_), .ZN(n9696) );
  AOI221_X1 U10920 ( .B1(SI_2_), .B2(keyinput_f30), .C1(SI_31_), .C2(
        keyinput_f1), .A(n9696), .ZN(n9703) );
  OAI22_X1 U10921 ( .A1(P2_RD_REG_SCAN_IN), .A2(keyinput_f33), .B1(
        keyinput_f64), .B2(P2_B_REG_SCAN_IN), .ZN(n9697) );
  AOI221_X1 U10922 ( .B1(P2_RD_REG_SCAN_IN), .B2(keyinput_f33), .C1(
        P2_B_REG_SCAN_IN), .C2(keyinput_f64), .A(n9697), .ZN(n9702) );
  OAI22_X1 U10923 ( .A1(SI_17_), .A2(keyinput_f15), .B1(keyinput_f81), .B2(
        P2_DATAO_REG_15__SCAN_IN), .ZN(n9698) );
  AOI221_X1 U10924 ( .B1(SI_17_), .B2(keyinput_f15), .C1(
        P2_DATAO_REG_15__SCAN_IN), .C2(keyinput_f81), .A(n9698), .ZN(n9701) );
  OAI22_X1 U10925 ( .A1(P2_STATE_REG_SCAN_IN), .A2(keyinput_f34), .B1(
        P2_REG3_REG_21__SCAN_IN), .B2(keyinput_f45), .ZN(n9699) );
  AOI221_X1 U10926 ( .B1(P2_STATE_REG_SCAN_IN), .B2(keyinput_f34), .C1(
        keyinput_f45), .C2(P2_REG3_REG_21__SCAN_IN), .A(n9699), .ZN(n9700) );
  NAND4_X1 U10927 ( .A1(n9703), .A2(n9702), .A3(n9701), .A4(n9700), .ZN(n9733)
         );
  OAI22_X1 U10928 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(keyinput_f103), .B1(
        keyinput_f32), .B2(SI_0_), .ZN(n9704) );
  AOI221_X1 U10929 ( .B1(P1_IR_REG_12__SCAN_IN), .B2(keyinput_f103), .C1(SI_0_), .C2(keyinput_f32), .A(n9704), .ZN(n9711) );
  OAI22_X1 U10930 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(keyinput_f96), .B1(
        keyinput_f51), .B2(P2_REG3_REG_24__SCAN_IN), .ZN(n9705) );
  AOI221_X1 U10931 ( .B1(P1_IR_REG_5__SCAN_IN), .B2(keyinput_f96), .C1(
        P2_REG3_REG_24__SCAN_IN), .C2(keyinput_f51), .A(n9705), .ZN(n9710) );
  OAI22_X1 U10932 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(keyinput_f108), .B1(SI_9_), 
        .B2(keyinput_f23), .ZN(n9706) );
  AOI221_X1 U10933 ( .B1(P1_IR_REG_17__SCAN_IN), .B2(keyinput_f108), .C1(
        keyinput_f23), .C2(SI_9_), .A(n9706), .ZN(n9709) );
  OAI22_X1 U10934 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(keyinput_f101), .B1(
        keyinput_f67), .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n9707) );
  AOI221_X1 U10935 ( .B1(P1_IR_REG_10__SCAN_IN), .B2(keyinput_f101), .C1(
        P2_DATAO_REG_29__SCAN_IN), .C2(keyinput_f67), .A(n9707), .ZN(n9708) );
  NAND4_X1 U10936 ( .A1(n9711), .A2(n9710), .A3(n9709), .A4(n9708), .ZN(n9732)
         );
  OAI22_X1 U10937 ( .A1(SI_14_), .A2(keyinput_f18), .B1(keyinput_f29), .B2(
        SI_3_), .ZN(n9712) );
  AOI221_X1 U10938 ( .B1(SI_14_), .B2(keyinput_f18), .C1(SI_3_), .C2(
        keyinput_f29), .A(n9712), .ZN(n9719) );
  OAI22_X1 U10939 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(keyinput_f104), .B1(
        keyinput_f95), .B2(P1_IR_REG_4__SCAN_IN), .ZN(n9713) );
  AOI221_X1 U10940 ( .B1(P1_IR_REG_13__SCAN_IN), .B2(keyinput_f104), .C1(
        P1_IR_REG_4__SCAN_IN), .C2(keyinput_f95), .A(n9713), .ZN(n9718) );
  OAI22_X1 U10941 ( .A1(SI_6_), .A2(keyinput_f26), .B1(keyinput_f90), .B2(
        P2_DATAO_REG_6__SCAN_IN), .ZN(n9714) );
  AOI221_X1 U10942 ( .B1(SI_6_), .B2(keyinput_f26), .C1(
        P2_DATAO_REG_6__SCAN_IN), .C2(keyinput_f90), .A(n9714), .ZN(n9717) );
  OAI22_X1 U10943 ( .A1(SI_23_), .A2(keyinput_f9), .B1(SI_20_), .B2(
        keyinput_f12), .ZN(n9715) );
  AOI221_X1 U10944 ( .B1(SI_23_), .B2(keyinput_f9), .C1(keyinput_f12), .C2(
        SI_20_), .A(n9715), .ZN(n9716) );
  NAND4_X1 U10945 ( .A1(n9719), .A2(n9718), .A3(n9717), .A4(n9716), .ZN(n9731)
         );
  OAI22_X1 U10946 ( .A1(P2_DATAO_REG_7__SCAN_IN), .A2(keyinput_f89), .B1(
        keyinput_f43), .B2(P2_REG3_REG_8__SCAN_IN), .ZN(n9720) );
  AOI221_X1 U10947 ( .B1(P2_DATAO_REG_7__SCAN_IN), .B2(keyinput_f89), .C1(
        P2_REG3_REG_8__SCAN_IN), .C2(keyinput_f43), .A(n9720), .ZN(n9729) );
  OAI22_X1 U10948 ( .A1(P1_IR_REG_25__SCAN_IN), .A2(keyinput_f116), .B1(
        keyinput_f3), .B2(SI_29_), .ZN(n9721) );
  AOI221_X1 U10949 ( .B1(P1_IR_REG_25__SCAN_IN), .B2(keyinput_f116), .C1(
        SI_29_), .C2(keyinput_f3), .A(n9721), .ZN(n9728) );
  OAI22_X1 U10950 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(keyinput_f74), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(keyinput_f59), .ZN(n9722) );
  AOI221_X1 U10951 ( .B1(P2_DATAO_REG_22__SCAN_IN), .B2(keyinput_f74), .C1(
        keyinput_f59), .C2(P2_REG3_REG_2__SCAN_IN), .A(n9722), .ZN(n9727) );
  XNOR2_X1 U10952 ( .A(n9723), .B(keyinput_f106), .ZN(n9725) );
  XNOR2_X1 U10953 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(keyinput_f65), .ZN(n9724)
         );
  NOR2_X1 U10954 ( .A1(n9725), .A2(n9724), .ZN(n9726) );
  NAND4_X1 U10955 ( .A1(n9729), .A2(n9728), .A3(n9727), .A4(n9726), .ZN(n9730)
         );
  NOR4_X1 U10956 ( .A1(n9733), .A2(n9732), .A3(n9731), .A4(n9730), .ZN(n9880)
         );
  OAI22_X1 U10957 ( .A1(P1_IR_REG_29__SCAN_IN), .A2(keyinput_f120), .B1(
        P2_REG3_REG_4__SCAN_IN), .B2(keyinput_f52), .ZN(n9734) );
  AOI221_X1 U10958 ( .B1(P1_IR_REG_29__SCAN_IN), .B2(keyinput_f120), .C1(
        keyinput_f52), .C2(P2_REG3_REG_4__SCAN_IN), .A(n9734), .ZN(n9741) );
  OAI22_X1 U10959 ( .A1(SI_13_), .A2(keyinput_f19), .B1(keyinput_f35), .B2(
        P2_REG3_REG_7__SCAN_IN), .ZN(n9735) );
  AOI221_X1 U10960 ( .B1(SI_13_), .B2(keyinput_f19), .C1(
        P2_REG3_REG_7__SCAN_IN), .C2(keyinput_f35), .A(n9735), .ZN(n9740) );
  OAI22_X1 U10961 ( .A1(P2_DATAO_REG_13__SCAN_IN), .A2(keyinput_f83), .B1(
        SI_5_), .B2(keyinput_f27), .ZN(n9736) );
  AOI221_X1 U10962 ( .B1(P2_DATAO_REG_13__SCAN_IN), .B2(keyinput_f83), .C1(
        keyinput_f27), .C2(SI_5_), .A(n9736), .ZN(n9739) );
  OAI22_X1 U10963 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(keyinput_f71), .B1(
        keyinput_f13), .B2(SI_19_), .ZN(n9737) );
  AOI221_X1 U10964 ( .B1(P2_DATAO_REG_25__SCAN_IN), .B2(keyinput_f71), .C1(
        SI_19_), .C2(keyinput_f13), .A(n9737), .ZN(n9738) );
  NAND4_X1 U10965 ( .A1(n9741), .A2(n9740), .A3(n9739), .A4(n9738), .ZN(n9878)
         );
  OAI22_X1 U10966 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(keyinput_f114), .B1(
        P2_REG3_REG_13__SCAN_IN), .B2(keyinput_f56), .ZN(n9742) );
  AOI221_X1 U10967 ( .B1(P1_IR_REG_23__SCAN_IN), .B2(keyinput_f114), .C1(
        keyinput_f56), .C2(P2_REG3_REG_13__SCAN_IN), .A(n9742), .ZN(n9767) );
  OAI22_X1 U10968 ( .A1(SI_22_), .A2(keyinput_f10), .B1(keyinput_f75), .B2(
        P2_DATAO_REG_21__SCAN_IN), .ZN(n9743) );
  AOI221_X1 U10969 ( .B1(SI_22_), .B2(keyinput_f10), .C1(
        P2_DATAO_REG_21__SCAN_IN), .C2(keyinput_f75), .A(n9743), .ZN(n9746) );
  OAI22_X1 U10970 ( .A1(SI_11_), .A2(keyinput_f21), .B1(keyinput_f62), .B2(
        P2_REG3_REG_26__SCAN_IN), .ZN(n9744) );
  AOI221_X1 U10971 ( .B1(SI_11_), .B2(keyinput_f21), .C1(
        P2_REG3_REG_26__SCAN_IN), .C2(keyinput_f62), .A(n9744), .ZN(n9745) );
  OAI211_X1 U10972 ( .C1(n8206), .C2(keyinput_f36), .A(n9746), .B(n9745), .ZN(
        n9747) );
  AOI21_X1 U10973 ( .B1(n8206), .B2(keyinput_f36), .A(n9747), .ZN(n9766) );
  AOI22_X1 U10974 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(keyinput_f61), .B1(
        P1_IR_REG_19__SCAN_IN), .B2(keyinput_f110), .ZN(n9748) );
  OAI221_X1 U10975 ( .B1(P2_REG3_REG_6__SCAN_IN), .B2(keyinput_f61), .C1(
        P1_IR_REG_19__SCAN_IN), .C2(keyinput_f110), .A(n9748), .ZN(n9755) );
  AOI22_X1 U10976 ( .A1(P2_REG3_REG_0__SCAN_IN), .A2(keyinput_f54), .B1(
        P1_IR_REG_31__SCAN_IN), .B2(keyinput_f122), .ZN(n9749) );
  OAI221_X1 U10977 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(keyinput_f54), .C1(
        P1_IR_REG_31__SCAN_IN), .C2(keyinput_f122), .A(n9749), .ZN(n9754) );
  AOI22_X1 U10978 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(keyinput_f58), .B1(
        SI_25_), .B2(keyinput_f7), .ZN(n9750) );
  OAI221_X1 U10979 ( .B1(P2_REG3_REG_11__SCAN_IN), .B2(keyinput_f58), .C1(
        SI_25_), .C2(keyinput_f7), .A(n9750), .ZN(n9753) );
  AOI22_X1 U10980 ( .A1(P2_DATAO_REG_11__SCAN_IN), .A2(keyinput_f85), .B1(
        P1_IR_REG_20__SCAN_IN), .B2(keyinput_f111), .ZN(n9751) );
  OAI221_X1 U10981 ( .B1(P2_DATAO_REG_11__SCAN_IN), .B2(keyinput_f85), .C1(
        P1_IR_REG_20__SCAN_IN), .C2(keyinput_f111), .A(n9751), .ZN(n9752) );
  NOR4_X1 U10982 ( .A1(n9755), .A2(n9754), .A3(n9753), .A4(n9752), .ZN(n9765)
         );
  AOI22_X1 U10983 ( .A1(P1_D_REG_1__SCAN_IN), .A2(keyinput_f124), .B1(
        P1_D_REG_0__SCAN_IN), .B2(keyinput_f123), .ZN(n9756) );
  OAI221_X1 U10984 ( .B1(P1_D_REG_1__SCAN_IN), .B2(keyinput_f124), .C1(
        P1_D_REG_0__SCAN_IN), .C2(keyinput_f123), .A(n9756), .ZN(n9763) );
  AOI22_X1 U10985 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(keyinput_f39), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(keyinput_f70), .ZN(n9757) );
  OAI221_X1 U10986 ( .B1(P2_REG3_REG_10__SCAN_IN), .B2(keyinput_f39), .C1(
        P2_DATAO_REG_26__SCAN_IN), .C2(keyinput_f70), .A(n9757), .ZN(n9762) );
  AOI22_X1 U10987 ( .A1(SI_16_), .A2(keyinput_f16), .B1(P1_IR_REG_18__SCAN_IN), 
        .B2(keyinput_f109), .ZN(n9758) );
  OAI221_X1 U10988 ( .B1(SI_16_), .B2(keyinput_f16), .C1(P1_IR_REG_18__SCAN_IN), .C2(keyinput_f109), .A(n9758), .ZN(n9761) );
  AOI22_X1 U10989 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(keyinput_f53), .B1(SI_12_), .B2(keyinput_f20), .ZN(n9759) );
  OAI221_X1 U10990 ( .B1(P2_REG3_REG_9__SCAN_IN), .B2(keyinput_f53), .C1(
        SI_12_), .C2(keyinput_f20), .A(n9759), .ZN(n9760) );
  NOR4_X1 U10991 ( .A1(n9763), .A2(n9762), .A3(n9761), .A4(n9760), .ZN(n9764)
         );
  NAND4_X1 U10992 ( .A1(n9767), .A2(n9766), .A3(n9765), .A4(n9764), .ZN(n9877)
         );
  AOI22_X1 U10993 ( .A1(n5563), .A2(keyinput_f8), .B1(keyinput_f38), .B2(n8214), .ZN(n9768) );
  OAI221_X1 U10994 ( .B1(n5563), .B2(keyinput_f8), .C1(n8214), .C2(
        keyinput_f38), .A(n9768), .ZN(n9777) );
  AOI22_X1 U10995 ( .A1(n5635), .A2(keyinput_f42), .B1(keyinput_f0), .B2(n9770), .ZN(n9769) );
  OAI221_X1 U10996 ( .B1(n5635), .B2(keyinput_f42), .C1(n9770), .C2(
        keyinput_f0), .A(n9769), .ZN(n9776) );
  XOR2_X1 U10997 ( .A(n5187), .B(keyinput_f49), .Z(n9774) );
  XNOR2_X1 U10998 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(keyinput_f84), .ZN(n9773)
         );
  XNOR2_X1 U10999 ( .A(P1_IR_REG_26__SCAN_IN), .B(keyinput_f117), .ZN(n9772)
         );
  XNOR2_X1 U11000 ( .A(P1_IR_REG_11__SCAN_IN), .B(keyinput_f102), .ZN(n9771)
         );
  NAND4_X1 U11001 ( .A1(n9774), .A2(n9773), .A3(n9772), .A4(n9771), .ZN(n9775)
         );
  NOR3_X1 U11002 ( .A1(n9777), .A2(n9776), .A3(n9775), .ZN(n9818) );
  AOI22_X1 U11003 ( .A1(n9780), .A2(keyinput_f24), .B1(n9779), .B2(
        keyinput_f72), .ZN(n9778) );
  OAI221_X1 U11004 ( .B1(n9780), .B2(keyinput_f24), .C1(n9779), .C2(
        keyinput_f72), .A(n9778), .ZN(n9788) );
  XOR2_X1 U11005 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput_f98), .Z(n9787) );
  XNOR2_X1 U11006 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(keyinput_f86), .ZN(n9784)
         );
  XNOR2_X1 U11007 ( .A(P1_IR_REG_0__SCAN_IN), .B(keyinput_f91), .ZN(n9783) );
  XNOR2_X1 U11008 ( .A(SI_7_), .B(keyinput_f25), .ZN(n9782) );
  XNOR2_X1 U11009 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput_f94), .ZN(n9781) );
  NAND4_X1 U11010 ( .A1(n9784), .A2(n9783), .A3(n9782), .A4(n9781), .ZN(n9786)
         );
  XNOR2_X1 U11011 ( .A(keyinput_f107), .B(n5988), .ZN(n9785) );
  NOR4_X1 U11012 ( .A1(n9788), .A2(n9787), .A3(n9786), .A4(n9785), .ZN(n9817)
         );
  AOI22_X1 U11013 ( .A1(n8358), .A2(keyinput_f63), .B1(n9790), .B2(
        keyinput_f79), .ZN(n9789) );
  OAI221_X1 U11014 ( .B1(n8358), .B2(keyinput_f63), .C1(n9790), .C2(
        keyinput_f79), .A(n9789), .ZN(n9802) );
  AOI22_X1 U11015 ( .A1(n9793), .A2(keyinput_f76), .B1(keyinput_f57), .B2(
        n9792), .ZN(n9791) );
  OAI221_X1 U11016 ( .B1(n9793), .B2(keyinput_f76), .C1(n9792), .C2(
        keyinput_f57), .A(n9791), .ZN(n9801) );
  AOI22_X1 U11017 ( .A1(n9796), .A2(keyinput_f77), .B1(keyinput_f22), .B2(
        n9795), .ZN(n9794) );
  OAI221_X1 U11018 ( .B1(n9796), .B2(keyinput_f77), .C1(n9795), .C2(
        keyinput_f22), .A(n9794), .ZN(n9800) );
  XOR2_X1 U11019 ( .A(n7714), .B(keyinput_f73), .Z(n9798) );
  XNOR2_X1 U11020 ( .A(P1_IR_REG_21__SCAN_IN), .B(keyinput_f112), .ZN(n9797)
         );
  NAND2_X1 U11021 ( .A1(n9798), .A2(n9797), .ZN(n9799) );
  NOR4_X1 U11022 ( .A1(n9802), .A2(n9801), .A3(n9800), .A4(n9799), .ZN(n9816)
         );
  INV_X1 U11023 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n10155) );
  AOI22_X1 U11024 ( .A1(n9804), .A2(keyinput_f60), .B1(n10155), .B2(
        keyinput_f127), .ZN(n9803) );
  OAI221_X1 U11025 ( .B1(n9804), .B2(keyinput_f60), .C1(n10155), .C2(
        keyinput_f127), .A(n9803), .ZN(n9814) );
  AOI22_X1 U11026 ( .A1(n9807), .A2(keyinput_f66), .B1(n9806), .B2(
        keyinput_f87), .ZN(n9805) );
  OAI221_X1 U11027 ( .B1(n9807), .B2(keyinput_f66), .C1(n9806), .C2(
        keyinput_f87), .A(n9805), .ZN(n9813) );
  XOR2_X1 U11028 ( .A(n6090), .B(keyinput_f97), .Z(n9811) );
  XOR2_X1 U11029 ( .A(n5915), .B(keyinput_f118), .Z(n9810) );
  XNOR2_X1 U11030 ( .A(SI_1_), .B(keyinput_f31), .ZN(n9809) );
  XNOR2_X1 U11031 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput_f119), .ZN(n9808)
         );
  NAND4_X1 U11032 ( .A1(n9811), .A2(n9810), .A3(n9809), .A4(n9808), .ZN(n9812)
         );
  NOR3_X1 U11033 ( .A1(n9814), .A2(n9813), .A3(n9812), .ZN(n9815) );
  NAND4_X1 U11034 ( .A1(n9818), .A2(n9817), .A3(n9816), .A4(n9815), .ZN(n9876)
         );
  AOI22_X1 U11035 ( .A1(n9821), .A2(keyinput_f46), .B1(keyinput_f40), .B2(
        n9820), .ZN(n9819) );
  OAI221_X1 U11036 ( .B1(n9821), .B2(keyinput_f46), .C1(n9820), .C2(
        keyinput_f40), .A(n9819), .ZN(n9831) );
  AOI22_X1 U11037 ( .A1(n9824), .A2(keyinput_f82), .B1(n9823), .B2(
        keyinput_f17), .ZN(n9822) );
  OAI221_X1 U11038 ( .B1(n9824), .B2(keyinput_f82), .C1(n9823), .C2(
        keyinput_f17), .A(n9822), .ZN(n9830) );
  XNOR2_X1 U11039 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(keyinput_f78), .ZN(n9828)
         );
  XNOR2_X1 U11040 ( .A(P1_IR_REG_14__SCAN_IN), .B(keyinput_f105), .ZN(n9827)
         );
  XNOR2_X1 U11041 ( .A(P2_REG3_REG_20__SCAN_IN), .B(keyinput_f55), .ZN(n9826)
         );
  XNOR2_X1 U11042 ( .A(SI_4_), .B(keyinput_f28), .ZN(n9825) );
  NAND4_X1 U11043 ( .A1(n9828), .A2(n9827), .A3(n9826), .A4(n9825), .ZN(n9829)
         );
  NOR3_X1 U11044 ( .A1(n9831), .A2(n9830), .A3(n9829), .ZN(n9874) );
  INV_X1 U11045 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n10156) );
  AOI22_X1 U11046 ( .A1(n10156), .A2(keyinput_f126), .B1(keyinput_f88), .B2(
        n9833), .ZN(n9832) );
  OAI221_X1 U11047 ( .B1(n10156), .B2(keyinput_f126), .C1(n9833), .C2(
        keyinput_f88), .A(n9832), .ZN(n9843) );
  AOI22_X1 U11048 ( .A1(n6139), .A2(keyinput_f99), .B1(keyinput_f121), .B2(
        n5925), .ZN(n9834) );
  OAI221_X1 U11049 ( .B1(n6139), .B2(keyinput_f99), .C1(n5925), .C2(
        keyinput_f121), .A(n9834), .ZN(n9842) );
  INV_X1 U11050 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n10157) );
  AOI22_X1 U11051 ( .A1(n10157), .A2(keyinput_f125), .B1(keyinput_f6), .B2(
        n9836), .ZN(n9835) );
  OAI221_X1 U11052 ( .B1(n10157), .B2(keyinput_f125), .C1(n9836), .C2(
        keyinput_f6), .A(n9835), .ZN(n9841) );
  INV_X1 U11053 ( .A(SI_21_), .ZN(n9838) );
  AOI22_X1 U11054 ( .A1(n9839), .A2(keyinput_f37), .B1(n9838), .B2(
        keyinput_f11), .ZN(n9837) );
  OAI221_X1 U11055 ( .B1(n9839), .B2(keyinput_f37), .C1(n9838), .C2(
        keyinput_f11), .A(n9837), .ZN(n9840) );
  NOR4_X1 U11056 ( .A1(n9843), .A2(n9842), .A3(n9841), .A4(n9840), .ZN(n9873)
         );
  AOI22_X1 U11057 ( .A1(n9845), .A2(keyinput_f4), .B1(keyinput_f50), .B2(n5441), .ZN(n9844) );
  OAI221_X1 U11058 ( .B1(n9845), .B2(keyinput_f4), .C1(n5441), .C2(
        keyinput_f50), .A(n9844), .ZN(n9856) );
  AOI22_X1 U11059 ( .A1(n9847), .A2(keyinput_f44), .B1(n6472), .B2(
        keyinput_f115), .ZN(n9846) );
  OAI221_X1 U11060 ( .B1(n9847), .B2(keyinput_f44), .C1(n6472), .C2(
        keyinput_f115), .A(n9846), .ZN(n9855) );
  AOI22_X1 U11061 ( .A1(n8270), .A2(keyinput_f47), .B1(n9849), .B2(
        keyinput_f80), .ZN(n9848) );
  OAI221_X1 U11062 ( .B1(n8270), .B2(keyinput_f47), .C1(n9849), .C2(
        keyinput_f80), .A(n9848), .ZN(n9854) );
  INV_X1 U11063 ( .A(SI_30_), .ZN(n9850) );
  XOR2_X1 U11064 ( .A(n9850), .B(keyinput_f2), .Z(n9852) );
  XNOR2_X1 U11065 ( .A(P1_IR_REG_22__SCAN_IN), .B(keyinput_f113), .ZN(n9851)
         );
  NAND2_X1 U11066 ( .A1(n9852), .A2(n9851), .ZN(n9853) );
  NOR4_X1 U11067 ( .A1(n9856), .A2(n9855), .A3(n9854), .A4(n9853), .ZN(n9872)
         );
  AOI22_X1 U11068 ( .A1(n9858), .A2(keyinput_f14), .B1(keyinput_f41), .B2(
        n5481), .ZN(n9857) );
  OAI221_X1 U11069 ( .B1(n9858), .B2(keyinput_f14), .C1(n5481), .C2(
        keyinput_f41), .A(n9857), .ZN(n9870) );
  AOI22_X1 U11070 ( .A1(n9860), .A2(keyinput_f48), .B1(n5898), .B2(
        keyinput_f93), .ZN(n9859) );
  OAI221_X1 U11071 ( .B1(n9860), .B2(keyinput_f48), .C1(n5898), .C2(
        keyinput_f93), .A(n9859), .ZN(n9869) );
  INV_X1 U11072 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n9862) );
  AOI22_X1 U11073 ( .A1(n9863), .A2(keyinput_f69), .B1(n9862), .B2(
        keyinput_f100), .ZN(n9861) );
  OAI221_X1 U11074 ( .B1(n9863), .B2(keyinput_f69), .C1(n9862), .C2(
        keyinput_f100), .A(n9861), .ZN(n9868) );
  AOI22_X1 U11075 ( .A1(n9866), .A2(keyinput_f68), .B1(n9865), .B2(keyinput_f5), .ZN(n9864) );
  OAI221_X1 U11076 ( .B1(n9866), .B2(keyinput_f68), .C1(n9865), .C2(
        keyinput_f5), .A(n9864), .ZN(n9867) );
  NOR4_X1 U11077 ( .A1(n9870), .A2(n9869), .A3(n9868), .A4(n9867), .ZN(n9871)
         );
  NAND4_X1 U11078 ( .A1(n9874), .A2(n9873), .A3(n9872), .A4(n9871), .ZN(n9875)
         );
  NOR4_X1 U11079 ( .A1(n9878), .A2(n9877), .A3(n9876), .A4(n9875), .ZN(n9879)
         );
  AOI22_X1 U11080 ( .A1(n9880), .A2(n9879), .B1(keyinput_f92), .B2(
        P1_IR_REG_1__SCAN_IN), .ZN(n9881) );
  OAI21_X1 U11081 ( .B1(keyinput_f92), .B2(P1_IR_REG_1__SCAN_IN), .A(n9881), 
        .ZN(n9882) );
  OAI21_X1 U11082 ( .B1(n9885), .B2(keyinput_g92), .A(n9882), .ZN(n9883) );
  AOI211_X1 U11083 ( .C1(n9885), .C2(keyinput_g92), .A(n9884), .B(n9883), .ZN(
        n9886) );
  XNOR2_X1 U11084 ( .A(n9887), .B(n9886), .ZN(n9891) );
  NOR2_X1 U11085 ( .A1(n9889), .A2(n9888), .ZN(n9890) );
  XOR2_X1 U11086 ( .A(n9891), .B(n9890), .Z(ADD_1071_U4) );
  AOI22_X1 U11087 ( .A1(n10234), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n9904) );
  AOI211_X1 U11088 ( .C1(n9894), .C2(n4788), .A(n9893), .B(n10237), .ZN(n9895)
         );
  AOI21_X1 U11089 ( .B1(n9897), .B2(n9896), .A(n9895), .ZN(n9903) );
  AOI211_X1 U11090 ( .C1(n9900), .C2(n9899), .A(n9898), .B(n10236), .ZN(n9901)
         );
  INV_X1 U11091 ( .A(n9901), .ZN(n9902) );
  NAND3_X1 U11092 ( .A1(n9904), .A2(n9903), .A3(n9902), .ZN(P2_U3247) );
  OAI21_X1 U11093 ( .B1(n9906), .B2(n10335), .A(n9905), .ZN(n9907) );
  AOI21_X1 U11094 ( .B1(n9908), .B2(n10246), .A(n9907), .ZN(n9917) );
  INV_X1 U11095 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n9909) );
  AOI22_X1 U11096 ( .A1(n10360), .A2(n9917), .B1(n9909), .B2(n10357), .ZN(
        P2_U3550) );
  OAI21_X1 U11097 ( .B1(n9911), .B2(n10335), .A(n9910), .ZN(n9913) );
  AOI211_X1 U11098 ( .C1(n9914), .C2(n10340), .A(n9913), .B(n9912), .ZN(n9919)
         );
  AOI22_X1 U11099 ( .A1(n10360), .A2(n9919), .B1(n9915), .B2(n10357), .ZN(
        P2_U3534) );
  INV_X1 U11100 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n9916) );
  AOI22_X1 U11101 ( .A1(n10344), .A2(n9917), .B1(n9916), .B2(n10342), .ZN(
        P2_U3518) );
  INV_X1 U11102 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n9918) );
  AOI22_X1 U11103 ( .A1(n10344), .A2(n9919), .B1(n9918), .B2(n10342), .ZN(
        P2_U3493) );
  OAI211_X1 U11104 ( .C1(n9922), .C2(n10207), .A(n9921), .B(n9920), .ZN(n9923)
         );
  AOI21_X1 U11105 ( .B1(n9924), .B2(n10195), .A(n9923), .ZN(n9951) );
  AOI22_X1 U11106 ( .A1(n10231), .A2(n9951), .B1(n6232), .B2(n10228), .ZN(
        P1_U3539) );
  NAND2_X1 U11107 ( .A1(n9925), .A2(n10177), .ZN(n9926) );
  OAI211_X1 U11108 ( .C1(n9928), .C2(n9931), .A(n9927), .B(n9926), .ZN(n9929)
         );
  NOR2_X1 U11109 ( .A1(n9930), .A2(n9929), .ZN(n9953) );
  AOI22_X1 U11110 ( .A1(n10231), .A2(n9953), .B1(n6221), .B2(n10228), .ZN(
        P1_U3538) );
  INV_X1 U11111 ( .A(n9931), .ZN(n10214) );
  OAI22_X1 U11112 ( .A1(n9933), .A2(n10209), .B1(n4762), .B2(n10207), .ZN(
        n9934) );
  AOI21_X1 U11113 ( .B1(n9935), .B2(n10214), .A(n9934), .ZN(n9936) );
  AND2_X1 U11114 ( .A1(n9937), .A2(n9936), .ZN(n9955) );
  AOI22_X1 U11115 ( .A1(n10231), .A2(n9955), .B1(n6189), .B2(n10228), .ZN(
        P1_U3536) );
  OAI21_X1 U11116 ( .B1(n9939), .B2(n10207), .A(n9938), .ZN(n9940) );
  AOI21_X1 U11117 ( .B1(n9941), .B2(n10214), .A(n9940), .ZN(n9942) );
  AOI22_X1 U11118 ( .A1(n10231), .A2(n9957), .B1(n6123), .B2(n10228), .ZN(
        P1_U3535) );
  OAI22_X1 U11119 ( .A1(n9945), .A2(n10209), .B1(n9944), .B2(n10207), .ZN(
        n9946) );
  AOI21_X1 U11120 ( .B1(n9947), .B2(n10214), .A(n9946), .ZN(n9948) );
  AND2_X1 U11121 ( .A1(n9949), .A2(n9948), .ZN(n9959) );
  AOI22_X1 U11122 ( .A1(n10231), .A2(n9959), .B1(n6156), .B2(n10228), .ZN(
        P1_U3534) );
  INV_X1 U11123 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n9950) );
  AOI22_X1 U11124 ( .A1(n10217), .A2(n9951), .B1(n9950), .B2(n10215), .ZN(
        P1_U3502) );
  INV_X1 U11125 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n9952) );
  AOI22_X1 U11126 ( .A1(n10217), .A2(n9953), .B1(n9952), .B2(n10215), .ZN(
        P1_U3499) );
  INV_X1 U11127 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n9954) );
  AOI22_X1 U11128 ( .A1(n10217), .A2(n9955), .B1(n9954), .B2(n10215), .ZN(
        P1_U3493) );
  INV_X1 U11129 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n9956) );
  AOI22_X1 U11130 ( .A1(n10217), .A2(n9957), .B1(n9956), .B2(n10215), .ZN(
        P1_U3490) );
  INV_X1 U11131 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n9958) );
  AOI22_X1 U11132 ( .A1(n10217), .A2(n9959), .B1(n9958), .B2(n10215), .ZN(
        P1_U3487) );
  XNOR2_X1 U11133 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  OR2_X1 U11134 ( .A1(n9961), .A2(n9960), .ZN(n9963) );
  OAI211_X1 U11135 ( .C1(n9965), .C2(n9964), .A(n9963), .B(n9962), .ZN(n9994)
         );
  NAND2_X1 U11136 ( .A1(n10068), .A2(P1_ADDR_REG_2__SCAN_IN), .ZN(n9972) );
  NAND2_X1 U11137 ( .A1(n10116), .A2(n9966), .ZN(n9971) );
  OAI211_X1 U11138 ( .C1(n9969), .C2(n9968), .A(n10030), .B(n9967), .ZN(n9970)
         );
  AND4_X1 U11139 ( .A1(n9994), .A2(n9972), .A3(n9971), .A4(n9970), .ZN(n9977)
         );
  OAI211_X1 U11140 ( .C1(n9975), .C2(n9974), .A(n10117), .B(n9973), .ZN(n9976)
         );
  OAI211_X1 U11141 ( .C1(P1_STATE_REG_SCAN_IN), .C2(n6033), .A(n9977), .B(
        n9976), .ZN(P1_U3243) );
  INV_X1 U11142 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9987) );
  INV_X1 U11143 ( .A(n9978), .ZN(n9982) );
  MUX2_X1 U11144 ( .A(n6874), .B(P1_REG1_REG_4__SCAN_IN), .S(n9979), .Z(n9981)
         );
  OAI21_X1 U11145 ( .B1(n9982), .B2(n9981), .A(n9980), .ZN(n9983) );
  NAND2_X1 U11146 ( .A1(n10117), .A2(n9983), .ZN(n9986) );
  NAND2_X1 U11147 ( .A1(n10116), .A2(n9984), .ZN(n9985) );
  OAI211_X1 U11148 ( .C1(n10123), .C2(n9987), .A(n9986), .B(n9985), .ZN(n9988)
         );
  INV_X1 U11149 ( .A(n9988), .ZN(n9996) );
  AOI21_X1 U11150 ( .B1(n9991), .B2(n9990), .A(n9989), .ZN(n9992) );
  OR2_X1 U11151 ( .A1(n10109), .A2(n9992), .ZN(n9993) );
  NAND4_X1 U11152 ( .A1(n9996), .A2(n9995), .A3(n9994), .A4(n9993), .ZN(
        P1_U3245) );
  AOI22_X1 U11153 ( .A1(n10068), .A2(P1_ADDR_REG_7__SCAN_IN), .B1(n9997), .B2(
        n10116), .ZN(n10009) );
  NAND2_X1 U11154 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3084), .ZN(n10008) );
  AOI21_X1 U11155 ( .B1(n10000), .B2(n9999), .A(n9998), .ZN(n10001) );
  OR2_X1 U11156 ( .A1(n10001), .A2(n10109), .ZN(n10007) );
  AOI21_X1 U11157 ( .B1(n10004), .B2(n10003), .A(n10002), .ZN(n10005) );
  OR2_X1 U11158 ( .A1(n10005), .A2(n10071), .ZN(n10006) );
  NAND4_X1 U11159 ( .A1(n10009), .A2(n10008), .A3(n10007), .A4(n10006), .ZN(
        P1_U3248) );
  AOI211_X1 U11160 ( .C1(n10012), .C2(n10011), .A(n10109), .B(n10010), .ZN(
        n10013) );
  AOI211_X1 U11161 ( .C1(n10116), .C2(n10015), .A(n10014), .B(n10013), .ZN(
        n10020) );
  OAI221_X1 U11162 ( .B1(n10018), .B2(n10017), .C1(n10018), .C2(n10016), .A(
        n10117), .ZN(n10019) );
  OAI211_X1 U11163 ( .C1(n10390), .C2(n10123), .A(n10020), .B(n10019), .ZN(
        P1_U3250) );
  AOI21_X1 U11164 ( .B1(n10023), .B2(n10022), .A(n10021), .ZN(n10033) );
  INV_X1 U11165 ( .A(n10024), .ZN(n10025) );
  AOI21_X1 U11166 ( .B1(n10116), .B2(n10026), .A(n10025), .ZN(n10032) );
  OAI21_X1 U11167 ( .B1(n10028), .B2(n4511), .A(n10027), .ZN(n10029) );
  AOI22_X1 U11168 ( .A1(n10030), .A2(n10029), .B1(n10068), .B2(
        P1_ADDR_REG_11__SCAN_IN), .ZN(n10031) );
  OAI211_X1 U11169 ( .C1(n10033), .C2(n10071), .A(n10032), .B(n10031), .ZN(
        P1_U3252) );
  AOI21_X1 U11170 ( .B1(n10036), .B2(n10035), .A(n10034), .ZN(n10045) );
  AOI21_X1 U11171 ( .B1(n10116), .B2(n10038), .A(n10037), .ZN(n10044) );
  AOI211_X1 U11172 ( .C1(n10041), .C2(n10040), .A(n10039), .B(n10109), .ZN(
        n10042) );
  AOI21_X1 U11173 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(n10068), .A(n10042), 
        .ZN(n10043) );
  OAI211_X1 U11174 ( .C1(n10045), .C2(n10071), .A(n10044), .B(n10043), .ZN(
        P1_U3253) );
  AOI21_X1 U11175 ( .B1(n10048), .B2(n10047), .A(n10046), .ZN(n10058) );
  AOI211_X1 U11176 ( .C1(n10051), .C2(n10050), .A(n10049), .B(n10109), .ZN(
        n10056) );
  OAI21_X1 U11177 ( .B1(n10054), .B2(n10053), .A(n10052), .ZN(n10055) );
  AOI211_X1 U11178 ( .C1(P1_ADDR_REG_13__SCAN_IN), .C2(n10068), .A(n10056), 
        .B(n10055), .ZN(n10057) );
  OAI21_X1 U11179 ( .B1(n10058), .B2(n10071), .A(n10057), .ZN(P1_U3254) );
  AOI21_X1 U11180 ( .B1(n10061), .B2(n10060), .A(n10059), .ZN(n10072) );
  INV_X1 U11181 ( .A(n10062), .ZN(n10063) );
  AOI21_X1 U11182 ( .B1(n10116), .B2(n10064), .A(n10063), .ZN(n10070) );
  AOI211_X1 U11183 ( .C1(n6178), .C2(n10066), .A(n10065), .B(n10109), .ZN(
        n10067) );
  AOI21_X1 U11184 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(n10068), .A(n10067), 
        .ZN(n10069) );
  OAI211_X1 U11185 ( .C1(n10072), .C2(n10071), .A(n10070), .B(n10069), .ZN(
        P1_U3255) );
  INV_X1 U11186 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n10082) );
  AND2_X1 U11187 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n10076) );
  AOI211_X1 U11188 ( .C1(n10074), .C2(n9337), .A(n10073), .B(n10109), .ZN(
        n10075) );
  AOI211_X1 U11189 ( .C1(n10116), .C2(n10077), .A(n10076), .B(n10075), .ZN(
        n10081) );
  OAI211_X1 U11190 ( .C1(P1_REG1_REG_15__SCAN_IN), .C2(n10079), .A(n10117), 
        .B(n10078), .ZN(n10080) );
  OAI211_X1 U11191 ( .C1(n10082), .C2(n10123), .A(n10081), .B(n10080), .ZN(
        P1_U3256) );
  INV_X1 U11192 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n10095) );
  INV_X1 U11193 ( .A(n10083), .ZN(n10088) );
  AOI211_X1 U11194 ( .C1(n10086), .C2(n10085), .A(n10084), .B(n10109), .ZN(
        n10087) );
  AOI211_X1 U11195 ( .C1(n10116), .C2(n10089), .A(n10088), .B(n10087), .ZN(
        n10094) );
  OAI211_X1 U11196 ( .C1(n10092), .C2(n10091), .A(n10117), .B(n10090), .ZN(
        n10093) );
  OAI211_X1 U11197 ( .C1(n10095), .C2(n10123), .A(n10094), .B(n10093), .ZN(
        P1_U3257) );
  INV_X1 U11198 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n10107) );
  AOI211_X1 U11199 ( .C1(n10098), .C2(n10097), .A(n10096), .B(n10109), .ZN(
        n10099) );
  AOI211_X1 U11200 ( .C1(n10116), .C2(n10101), .A(n10100), .B(n10099), .ZN(
        n10106) );
  OAI211_X1 U11201 ( .C1(n10104), .C2(n10103), .A(n10117), .B(n10102), .ZN(
        n10105) );
  OAI211_X1 U11202 ( .C1(n10107), .C2(n10123), .A(n10106), .B(n10105), .ZN(
        P1_U3258) );
  NOR2_X1 U11203 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10108), .ZN(n10114) );
  AOI211_X1 U11204 ( .C1(n10112), .C2(n10111), .A(n10110), .B(n10109), .ZN(
        n10113) );
  AOI211_X1 U11205 ( .C1(n10116), .C2(n10115), .A(n10114), .B(n10113), .ZN(
        n10122) );
  OAI221_X1 U11206 ( .B1(n10120), .B2(n10119), .C1(n10120), .C2(n10118), .A(
        n10117), .ZN(n10121) );
  OAI211_X1 U11207 ( .C1(n10400), .C2(n10123), .A(n10122), .B(n10121), .ZN(
        P1_U3259) );
  OAI211_X1 U11208 ( .C1(n10144), .C2(n10160), .A(n10125), .B(n10124), .ZN(
        n10159) );
  INV_X1 U11209 ( .A(n10126), .ZN(n10129) );
  XNOR2_X1 U11210 ( .A(n10127), .B(n10129), .ZN(n10134) );
  NOR2_X1 U11211 ( .A1(n10139), .A2(n10130), .ZN(n10131) );
  AOI211_X1 U11212 ( .C1(n10134), .C2(n10133), .A(n10132), .B(n10131), .ZN(
        n10161) );
  AOI22_X1 U11213 ( .A1(n6553), .A2(n10136), .B1(P1_REG3_REG_1__SCAN_IN), .B2(
        n10135), .ZN(n10137) );
  OAI211_X1 U11214 ( .C1(n10138), .C2(n10159), .A(n10161), .B(n10137), .ZN(
        n10141) );
  INV_X1 U11215 ( .A(n10139), .ZN(n10164) );
  AOI22_X1 U11216 ( .A1(n10141), .A2(n10143), .B1(n10164), .B2(n10140), .ZN(
        n10142) );
  OAI21_X1 U11217 ( .B1(n6859), .B2(n10143), .A(n10142), .ZN(P1_U3290) );
  AOI21_X1 U11218 ( .B1(n10146), .B2(n10145), .A(n10144), .ZN(n10149) );
  NOR2_X1 U11219 ( .A1(n10147), .A2(n9242), .ZN(n10148) );
  AOI211_X1 U11220 ( .C1(n9242), .C2(P1_REG2_REG_0__SCAN_IN), .A(n10149), .B(
        n10148), .ZN(n10150) );
  OAI21_X1 U11221 ( .B1(n10151), .B2(n6839), .A(n10150), .ZN(P1_U3291) );
  AND2_X1 U11222 ( .A1(n10153), .A2(n10152), .ZN(n10158) );
  AND2_X1 U11223 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n10154), .ZN(P1_U3292) );
  AND2_X1 U11224 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n10154), .ZN(P1_U3293) );
  AND2_X1 U11225 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n10154), .ZN(P1_U3294) );
  AND2_X1 U11226 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n10154), .ZN(P1_U3295) );
  AND2_X1 U11227 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n10154), .ZN(P1_U3296) );
  AND2_X1 U11228 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10154), .ZN(P1_U3297) );
  AND2_X1 U11229 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10154), .ZN(P1_U3298) );
  AND2_X1 U11230 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n10154), .ZN(P1_U3299) );
  AND2_X1 U11231 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n10154), .ZN(P1_U3300) );
  AND2_X1 U11232 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n10154), .ZN(P1_U3301) );
  AND2_X1 U11233 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n10154), .ZN(P1_U3302) );
  AND2_X1 U11234 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n10154), .ZN(P1_U3303) );
  AND2_X1 U11235 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n10154), .ZN(P1_U3304) );
  AND2_X1 U11236 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n10154), .ZN(P1_U3305) );
  AND2_X1 U11237 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n10154), .ZN(P1_U3306) );
  AND2_X1 U11238 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n10154), .ZN(P1_U3307) );
  AND2_X1 U11239 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n10154), .ZN(P1_U3308) );
  AND2_X1 U11240 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n10154), .ZN(P1_U3309) );
  AND2_X1 U11241 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n10154), .ZN(P1_U3310) );
  AND2_X1 U11242 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n10154), .ZN(P1_U3311) );
  AND2_X1 U11243 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n10154), .ZN(P1_U3312) );
  AND2_X1 U11244 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n10154), .ZN(P1_U3313) );
  AND2_X1 U11245 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10154), .ZN(P1_U3314) );
  AND2_X1 U11246 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n10154), .ZN(P1_U3315) );
  AND2_X1 U11247 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n10154), .ZN(P1_U3316) );
  AND2_X1 U11248 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n10154), .ZN(P1_U3317) );
  AND2_X1 U11249 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n10154), .ZN(P1_U3318) );
  NOR2_X1 U11250 ( .A1(n10158), .A2(n10155), .ZN(P1_U3319) );
  NOR2_X1 U11251 ( .A1(n10158), .A2(n10156), .ZN(P1_U3320) );
  NOR2_X1 U11252 ( .A1(n10158), .A2(n10157), .ZN(P1_U3321) );
  OAI21_X1 U11253 ( .B1(n10160), .B2(n10207), .A(n10159), .ZN(n10163) );
  INV_X1 U11254 ( .A(n10161), .ZN(n10162) );
  AOI211_X1 U11255 ( .C1(n10214), .C2(n10164), .A(n10163), .B(n10162), .ZN(
        n10219) );
  AOI22_X1 U11256 ( .A1(n10217), .A2(n10219), .B1(n6014), .B2(n10215), .ZN(
        P1_U3457) );
  OAI22_X1 U11257 ( .A1(n10165), .A2(n10209), .B1(n6046), .B2(n10207), .ZN(
        n10167) );
  AOI211_X1 U11258 ( .C1(n10214), .C2(n10168), .A(n10167), .B(n10166), .ZN(
        n10220) );
  AOI22_X1 U11259 ( .A1(n10217), .A2(n10220), .B1(n6031), .B2(n10215), .ZN(
        P1_U3460) );
  INV_X1 U11260 ( .A(n10169), .ZN(n10173) );
  OAI22_X1 U11261 ( .A1(n10170), .A2(n10209), .B1(n6542), .B2(n10207), .ZN(
        n10172) );
  AOI211_X1 U11262 ( .C1(n10214), .C2(n10173), .A(n10172), .B(n10171), .ZN(
        n10221) );
  INV_X1 U11263 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n10174) );
  AOI22_X1 U11264 ( .A1(n10217), .A2(n10221), .B1(n10174), .B2(n10215), .ZN(
        P1_U3463) );
  AOI21_X1 U11265 ( .B1(n10177), .B2(n10176), .A(n10175), .ZN(n10181) );
  NAND3_X1 U11266 ( .A1(n10179), .A2(n10178), .A3(n10195), .ZN(n10180) );
  AND3_X1 U11267 ( .A1(n10182), .A2(n10181), .A3(n10180), .ZN(n10223) );
  INV_X1 U11268 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n10183) );
  AOI22_X1 U11269 ( .A1(n10217), .A2(n10223), .B1(n10183), .B2(n10215), .ZN(
        P1_U3469) );
  OAI22_X1 U11270 ( .A1(n10185), .A2(n10209), .B1(n10184), .B2(n10207), .ZN(
        n10187) );
  AOI211_X1 U11271 ( .C1(n10214), .C2(n10188), .A(n10187), .B(n10186), .ZN(
        n10224) );
  INV_X1 U11272 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10189) );
  AOI22_X1 U11273 ( .A1(n10217), .A2(n10224), .B1(n10189), .B2(n10215), .ZN(
        P1_U3472) );
  OAI211_X1 U11274 ( .C1(n10192), .C2(n10207), .A(n10191), .B(n10190), .ZN(
        n10193) );
  AOI21_X1 U11275 ( .B1(n10195), .B2(n10194), .A(n10193), .ZN(n10225) );
  INV_X1 U11276 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n10196) );
  AOI22_X1 U11277 ( .A1(n10217), .A2(n10225), .B1(n10196), .B2(n10215), .ZN(
        P1_U3475) );
  NOR2_X1 U11278 ( .A1(n10198), .A2(n10197), .ZN(n10204) );
  OAI22_X1 U11279 ( .A1(n10200), .A2(n10209), .B1(n10199), .B2(n10207), .ZN(
        n10202) );
  AOI211_X1 U11280 ( .C1(n10204), .C2(n10203), .A(n10202), .B(n10201), .ZN(
        n10227) );
  INV_X1 U11281 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n10205) );
  AOI22_X1 U11282 ( .A1(n10217), .A2(n10227), .B1(n10205), .B2(n10215), .ZN(
        P1_U3478) );
  INV_X1 U11283 ( .A(n10206), .ZN(n10213) );
  OAI22_X1 U11284 ( .A1(n10210), .A2(n10209), .B1(n10208), .B2(n10207), .ZN(
        n10212) );
  AOI211_X1 U11285 ( .C1(n10214), .C2(n10213), .A(n10212), .B(n10211), .ZN(
        n10230) );
  INV_X1 U11286 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10216) );
  AOI22_X1 U11287 ( .A1(n10217), .A2(n10230), .B1(n10216), .B2(n10215), .ZN(
        P1_U3481) );
  AOI22_X1 U11288 ( .A1(n10231), .A2(n10219), .B1(n10218), .B2(n10228), .ZN(
        P1_U3524) );
  AOI22_X1 U11289 ( .A1(n10231), .A2(n10220), .B1(n6847), .B2(n10228), .ZN(
        P1_U3525) );
  AOI22_X1 U11290 ( .A1(n10231), .A2(n10221), .B1(n6871), .B2(n10228), .ZN(
        P1_U3526) );
  AOI22_X1 U11291 ( .A1(n10231), .A2(n10223), .B1(n10222), .B2(n10228), .ZN(
        P1_U3528) );
  AOI22_X1 U11292 ( .A1(n10231), .A2(n10224), .B1(n6079), .B2(n10228), .ZN(
        P1_U3529) );
  AOI22_X1 U11293 ( .A1(n10231), .A2(n10225), .B1(n6896), .B2(n10228), .ZN(
        P1_U3530) );
  AOI22_X1 U11294 ( .A1(n10231), .A2(n10227), .B1(n10226), .B2(n10228), .ZN(
        P1_U3531) );
  AOI22_X1 U11295 ( .A1(n10231), .A2(n10230), .B1(n10229), .B2(n10228), .ZN(
        P1_U3532) );
  AOI22_X1 U11296 ( .A1(n10233), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n10232), .ZN(n10242) );
  AOI22_X1 U11297 ( .A1(n10234), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n10241) );
  OAI21_X1 U11298 ( .B1(P2_REG1_REG_0__SCAN_IN), .B2(n10236), .A(n10235), .ZN(
        n10239) );
  NOR2_X1 U11299 ( .A1(n10237), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n10238) );
  OAI21_X1 U11300 ( .B1(n10239), .B2(n10238), .A(P2_IR_REG_0__SCAN_IN), .ZN(
        n10240) );
  OAI211_X1 U11301 ( .C1(P2_IR_REG_0__SCAN_IN), .C2(n10242), .A(n10241), .B(
        n10240), .ZN(P2_U3245) );
  INV_X1 U11302 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n10265) );
  XNOR2_X1 U11303 ( .A(n10243), .B(n10251), .ZN(n10319) );
  OAI21_X1 U11304 ( .B1(n10245), .B2(n10244), .A(n10259), .ZN(n10247) );
  NAND3_X1 U11305 ( .A1(n10248), .A2(n10247), .A3(n10246), .ZN(n10315) );
  NAND2_X1 U11306 ( .A1(n10250), .A2(n10249), .ZN(n10252) );
  XNOR2_X1 U11307 ( .A(n10252), .B(n10251), .ZN(n10255) );
  AOI21_X1 U11308 ( .B1(n10255), .B2(n10254), .A(n10253), .ZN(n10316) );
  AOI22_X1 U11309 ( .A1(n10259), .A2(n10258), .B1(n10257), .B2(n10256), .ZN(
        n10260) );
  OAI211_X1 U11310 ( .C1(n4781), .C2(n10315), .A(n10316), .B(n10260), .ZN(
        n10261) );
  AOI21_X1 U11311 ( .B1(n10262), .B2(n10319), .A(n10261), .ZN(n10264) );
  AOI22_X1 U11312 ( .A1(n10266), .A2(n10265), .B1(n10264), .B2(n10263), .ZN(
        P2_U3291) );
  INV_X1 U11313 ( .A(n10267), .ZN(n10269) );
  NAND2_X1 U11314 ( .A1(n10269), .A2(n10268), .ZN(n10272) );
  AND2_X1 U11315 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n10272), .ZN(P2_U3297) );
  AND2_X1 U11316 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n10272), .ZN(P2_U3298) );
  AND2_X1 U11317 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n10272), .ZN(P2_U3299) );
  AND2_X1 U11318 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n10272), .ZN(P2_U3300) );
  AND2_X1 U11319 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n10272), .ZN(P2_U3301) );
  AND2_X1 U11320 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n10272), .ZN(P2_U3302) );
  AND2_X1 U11321 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n10272), .ZN(P2_U3303) );
  AND2_X1 U11322 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n10272), .ZN(P2_U3304) );
  AND2_X1 U11323 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n10272), .ZN(P2_U3305) );
  AND2_X1 U11324 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n10272), .ZN(P2_U3306) );
  AND2_X1 U11325 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n10272), .ZN(P2_U3307) );
  AND2_X1 U11326 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n10272), .ZN(P2_U3308) );
  AND2_X1 U11327 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n10272), .ZN(P2_U3309) );
  AND2_X1 U11328 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n10272), .ZN(P2_U3310) );
  AND2_X1 U11329 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n10272), .ZN(P2_U3311) );
  AND2_X1 U11330 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n10272), .ZN(P2_U3312) );
  AND2_X1 U11331 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n10272), .ZN(P2_U3313) );
  AND2_X1 U11332 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n10272), .ZN(P2_U3314) );
  AND2_X1 U11333 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n10272), .ZN(P2_U3315) );
  AND2_X1 U11334 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n10272), .ZN(P2_U3316) );
  AND2_X1 U11335 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n10272), .ZN(P2_U3317) );
  AND2_X1 U11336 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n10272), .ZN(P2_U3318) );
  AND2_X1 U11337 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n10272), .ZN(P2_U3319) );
  AND2_X1 U11338 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n10272), .ZN(P2_U3320) );
  AND2_X1 U11339 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n10272), .ZN(P2_U3321) );
  AND2_X1 U11340 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n10272), .ZN(P2_U3322) );
  AND2_X1 U11341 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n10272), .ZN(P2_U3323) );
  AND2_X1 U11342 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n10272), .ZN(P2_U3324) );
  AND2_X1 U11343 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n10272), .ZN(P2_U3325) );
  AND2_X1 U11344 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n10272), .ZN(P2_U3326) );
  AOI22_X1 U11345 ( .A1(n10271), .A2(n10272), .B1(n10275), .B2(n10270), .ZN(
        P2_U3437) );
  AOI22_X1 U11346 ( .A1(n10275), .A2(n10274), .B1(n10273), .B2(n10272), .ZN(
        P2_U3438) );
  OAI22_X1 U11347 ( .A1(n10278), .A2(n10288), .B1(n10277), .B2(n10276), .ZN(
        n10279) );
  NOR2_X1 U11348 ( .A1(n10280), .A2(n10279), .ZN(n10345) );
  INV_X1 U11349 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n10281) );
  AOI22_X1 U11350 ( .A1(n10344), .A2(n10345), .B1(n10281), .B2(n10342), .ZN(
        P2_U3451) );
  AOI21_X1 U11351 ( .B1(n10284), .B2(n4581), .A(n10282), .ZN(n10285) );
  OAI211_X1 U11352 ( .C1(n10288), .C2(n10287), .A(n10286), .B(n10285), .ZN(
        n10289) );
  INV_X1 U11353 ( .A(n10289), .ZN(n10347) );
  INV_X1 U11354 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10290) );
  AOI22_X1 U11355 ( .A1(n10344), .A2(n10347), .B1(n10290), .B2(n10342), .ZN(
        P2_U3454) );
  INV_X1 U11356 ( .A(n10291), .ZN(n10296) );
  OAI22_X1 U11357 ( .A1(n10292), .A2(n10336), .B1(n7034), .B2(n10335), .ZN(
        n10295) );
  INV_X1 U11358 ( .A(n10293), .ZN(n10294) );
  AOI211_X1 U11359 ( .C1(n10340), .C2(n10296), .A(n10295), .B(n10294), .ZN(
        n10349) );
  INV_X1 U11360 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10297) );
  AOI22_X1 U11361 ( .A1(n10344), .A2(n10349), .B1(n10297), .B2(n10342), .ZN(
        P2_U3457) );
  INV_X1 U11362 ( .A(n10299), .ZN(n10305) );
  NOR2_X1 U11363 ( .A1(n10299), .A2(n10298), .ZN(n10304) );
  OAI211_X1 U11364 ( .C1(n10302), .C2(n10335), .A(n10301), .B(n10300), .ZN(
        n10303) );
  AOI211_X1 U11365 ( .C1(n10305), .C2(n10333), .A(n10304), .B(n10303), .ZN(
        n10351) );
  INV_X1 U11366 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10306) );
  AOI22_X1 U11367 ( .A1(n10344), .A2(n10351), .B1(n10306), .B2(n10342), .ZN(
        P2_U3460) );
  INV_X1 U11368 ( .A(n10307), .ZN(n10313) );
  OAI22_X1 U11369 ( .A1(n10309), .A2(n10336), .B1(n10308), .B2(n10335), .ZN(
        n10312) );
  INV_X1 U11370 ( .A(n10310), .ZN(n10311) );
  AOI211_X1 U11371 ( .C1(n10340), .C2(n10313), .A(n10312), .B(n10311), .ZN(
        n10352) );
  INV_X1 U11372 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10314) );
  AOI22_X1 U11373 ( .A1(n10344), .A2(n10352), .B1(n10314), .B2(n10342), .ZN(
        P2_U3463) );
  OAI211_X1 U11374 ( .C1(n10317), .C2(n10335), .A(n10316), .B(n10315), .ZN(
        n10318) );
  AOI21_X1 U11375 ( .B1(n10340), .B2(n10319), .A(n10318), .ZN(n10353) );
  INV_X1 U11376 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10320) );
  AOI22_X1 U11377 ( .A1(n10344), .A2(n10353), .B1(n10320), .B2(n10342), .ZN(
        P2_U3466) );
  OAI22_X1 U11378 ( .A1(n10322), .A2(n10336), .B1(n10321), .B2(n10335), .ZN(
        n10324) );
  AOI211_X1 U11379 ( .C1(n10333), .C2(n10325), .A(n10324), .B(n10323), .ZN(
        n10355) );
  INV_X1 U11380 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10326) );
  AOI22_X1 U11381 ( .A1(n10344), .A2(n10355), .B1(n10326), .B2(n10342), .ZN(
        P2_U3475) );
  INV_X1 U11382 ( .A(n10327), .ZN(n10332) );
  OAI22_X1 U11383 ( .A1(n10329), .A2(n10336), .B1(n10328), .B2(n10335), .ZN(
        n10331) );
  AOI211_X1 U11384 ( .C1(n10333), .C2(n10332), .A(n10331), .B(n10330), .ZN(
        n10356) );
  INV_X1 U11385 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10334) );
  AOI22_X1 U11386 ( .A1(n10344), .A2(n10356), .B1(n10334), .B2(n10342), .ZN(
        P2_U3481) );
  OAI22_X1 U11387 ( .A1(n10337), .A2(n10336), .B1(n4729), .B2(n10335), .ZN(
        n10339) );
  AOI211_X1 U11388 ( .C1(n10341), .C2(n10340), .A(n10339), .B(n10338), .ZN(
        n10359) );
  INV_X1 U11389 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10343) );
  AOI22_X1 U11390 ( .A1(n10344), .A2(n10359), .B1(n10343), .B2(n10342), .ZN(
        P2_U3487) );
  AOI22_X1 U11391 ( .A1(n10360), .A2(n10345), .B1(n7062), .B2(n10357), .ZN(
        P2_U3520) );
  AOI22_X1 U11392 ( .A1(n10360), .A2(n10347), .B1(n10346), .B2(n10357), .ZN(
        P2_U3521) );
  AOI22_X1 U11393 ( .A1(n10360), .A2(n10349), .B1(n10348), .B2(n10357), .ZN(
        P2_U3522) );
  AOI22_X1 U11394 ( .A1(n10360), .A2(n10351), .B1(n10350), .B2(n10357), .ZN(
        P2_U3523) );
  AOI22_X1 U11395 ( .A1(n10360), .A2(n10352), .B1(n7122), .B2(n10357), .ZN(
        P2_U3524) );
  AOI22_X1 U11396 ( .A1(n10360), .A2(n10353), .B1(n7061), .B2(n10357), .ZN(
        P2_U3525) );
  AOI22_X1 U11397 ( .A1(n10360), .A2(n10355), .B1(n10354), .B2(n10357), .ZN(
        P2_U3528) );
  AOI22_X1 U11398 ( .A1(n10360), .A2(n10356), .B1(n7284), .B2(n10357), .ZN(
        P2_U3530) );
  AOI22_X1 U11399 ( .A1(n10360), .A2(n10359), .B1(n10358), .B2(n10357), .ZN(
        P2_U3532) );
  INV_X1 U11400 ( .A(n10361), .ZN(n10362) );
  NAND2_X1 U11401 ( .A1(n10363), .A2(n10362), .ZN(n10364) );
  XNOR2_X1 U11402 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n10364), .ZN(ADD_1071_U5)
         );
  XOR2_X1 U11403 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  OAI21_X1 U11404 ( .B1(n10367), .B2(n10366), .A(n10365), .ZN(ADD_1071_U56) );
  OAI21_X1 U11405 ( .B1(n10370), .B2(n10369), .A(n10368), .ZN(ADD_1071_U57) );
  OAI21_X1 U11406 ( .B1(n10373), .B2(n10372), .A(n10371), .ZN(ADD_1071_U58) );
  OAI21_X1 U11407 ( .B1(n10376), .B2(n10375), .A(n10374), .ZN(ADD_1071_U59) );
  OAI21_X1 U11408 ( .B1(n10379), .B2(n10378), .A(n10377), .ZN(ADD_1071_U60) );
  OAI21_X1 U11409 ( .B1(n10382), .B2(n10381), .A(n10380), .ZN(ADD_1071_U61) );
  AOI21_X1 U11410 ( .B1(n10385), .B2(n10384), .A(n10383), .ZN(ADD_1071_U62) );
  AOI21_X1 U11411 ( .B1(n10388), .B2(n10387), .A(n10386), .ZN(ADD_1071_U63) );
  AOI21_X1 U11412 ( .B1(n10391), .B2(n10390), .A(n10389), .ZN(ADD_1071_U47) );
  XOR2_X1 U11413 ( .A(n10392), .B(P2_ADDR_REG_7__SCAN_IN), .Z(ADD_1071_U49) );
  XOR2_X1 U11414 ( .A(n10394), .B(n10393), .Z(ADD_1071_U54) );
  NOR2_X1 U11415 ( .A1(n10396), .A2(n10395), .ZN(n10397) );
  XOR2_X1 U11416 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n10397), .Z(ADD_1071_U51) );
  OAI21_X1 U11417 ( .B1(n10400), .B2(n10399), .A(n10398), .ZN(n10401) );
  XNOR2_X1 U11418 ( .A(n10401), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  XOR2_X1 U11419 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n10402), .Z(ADD_1071_U48) );
  XOR2_X1 U11420 ( .A(P2_ADDR_REG_6__SCAN_IN), .B(n10403), .Z(ADD_1071_U50) );
  XOR2_X1 U11421 ( .A(n10405), .B(n10404), .Z(ADD_1071_U53) );
  XNOR2_X1 U11422 ( .A(n10407), .B(n10406), .ZN(ADD_1071_U52) );
  INV_X1 U5073 ( .A(n5283), .ZN(n5692) );
  CLKBUF_X1 U4995 ( .A(n5159), .Z(n4482) );
  CLKBUF_X1 U4997 ( .A(n5134), .Z(n5675) );
  NAND2_X2 U5001 ( .A1(n7089), .A2(n8484), .ZN(n5142) );
  CLKBUF_X1 U6546 ( .A(n6034), .Z(n6235) );
endmodule

