

module b15_C_gen_AntiSAT_k_256_10 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput_f0, keyinput_f1, 
        keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, 
        keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, 
        keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, 
        keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, 
        keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, 
        keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, 
        keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, 
        keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, 
        keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, 
        keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, 
        keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, 
        keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, 
        keyinput_f62, keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66, 
        keyinput_f67, keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71, 
        keyinput_f72, keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76, 
        keyinput_f77, keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81, 
        keyinput_f82, keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86, 
        keyinput_f87, keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91, 
        keyinput_f92, keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96, 
        keyinput_f97, keyinput_f98, keyinput_f99, keyinput_f100, keyinput_f101, 
        keyinput_f102, keyinput_f103, keyinput_f104, keyinput_f105, 
        keyinput_f106, keyinput_f107, keyinput_f108, keyinput_f109, 
        keyinput_f110, keyinput_f111, keyinput_f112, keyinput_f113, 
        keyinput_f114, keyinput_f115, keyinput_f116, keyinput_f117, 
        keyinput_f118, keyinput_f119, keyinput_f120, keyinput_f121, 
        keyinput_f122, keyinput_f123, keyinput_f124, keyinput_f125, 
        keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, keyinput_g2, 
        keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, 
        keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, 
        keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, 
        keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, 
        keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, 
        keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, 
        keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, 
        keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, 
        keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, 
        keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, 
        keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, 
        keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, 
        keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, keyinput_g67, 
        keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, keyinput_g72, 
        keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, keyinput_g77, 
        keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, keyinput_g82, 
        keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, keyinput_g87, 
        keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, keyinput_g92, 
        keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, keyinput_g97, 
        keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101, 
        keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105, 
        keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109, 
        keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113, 
        keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117, 
        keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121, 
        keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125, 
        keyinput_g126, keyinput_g127, U3445, U3446, U3447, U3448, U3213, U3212, 
        U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, U3203, U3202, 
        U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, U3193, U3192, 
        U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, U3183, U3182, 
        U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, U3175, U3174, 
        U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, U3165, U3164, 
        U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, U3155, U3154, 
        U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, U3146, U3145, 
        U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, U3136, U3135, 
        U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, U3126, U3125, 
        U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, U3116, U3115, 
        U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, U3106, U3105, 
        U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, U3096, U3095, 
        U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, U3086, U3085, 
        U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, U3076, U3075, 
        U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, U3066, U3065, 
        U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, U3056, U3055, 
        U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, U3046, U3045, 
        U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, U3036, U3035, 
        U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, U3026, U3025, 
        U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, U3460, U3461, 
        U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, U3015, U3014, 
        U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, U3005, U3004, 
        U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, U2995, U2994, 
        U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, U2985, U2984, 
        U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, U2975, U2974, 
        U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, U2965, U2964, 
        U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, U2955, U2954, 
        U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, U2945, U2944, 
        U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, U2935, U2934, 
        U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, U2925, U2924, 
        U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, U2915, U2914, 
        U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, U2905, U2904, 
        U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, U2895, U2894, 
        U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, U2885, U2884, 
        U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, U2875, U2874, 
        U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, U2865, U2864, 
        U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, U2855, U2854, 
        U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, U2845, U2844, 
        U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, U2835, U2834, 
        U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, U2825, U2824, 
        U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, U2815, U2814, 
        U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, U2805, U2804, 
        U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, U2795, U3468, 
        U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, U3473, U2790, 
        U2789, U3474, U2788 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput_f0, keyinput_f1,
         keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6,
         keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11,
         keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16,
         keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21,
         keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26,
         keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31,
         keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36,
         keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41,
         keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46,
         keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51,
         keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56,
         keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61,
         keyinput_f62, keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66,
         keyinput_f67, keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71,
         keyinput_f72, keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76,
         keyinput_f77, keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81,
         keyinput_f82, keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86,
         keyinput_f87, keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91,
         keyinput_f92, keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96,
         keyinput_f97, keyinput_f98, keyinput_f99, keyinput_f100,
         keyinput_f101, keyinput_f102, keyinput_f103, keyinput_f104,
         keyinput_f105, keyinput_f106, keyinput_f107, keyinput_f108,
         keyinput_f109, keyinput_f110, keyinput_f111, keyinput_f112,
         keyinput_f113, keyinput_f114, keyinput_f115, keyinput_f116,
         keyinput_f117, keyinput_f118, keyinput_f119, keyinput_f120,
         keyinput_f121, keyinput_f122, keyinput_f123, keyinput_f124,
         keyinput_f125, keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1,
         keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6,
         keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11,
         keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16,
         keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21,
         keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26,
         keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31,
         keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36,
         keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41,
         keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46,
         keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51,
         keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56,
         keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61,
         keyinput_g62, keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66,
         keyinput_g67, keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71,
         keyinput_g72, keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76,
         keyinput_g77, keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81,
         keyinput_g82, keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86,
         keyinput_g87, keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91,
         keyinput_g92, keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96,
         keyinput_g97, keyinput_g98, keyinput_g99, keyinput_g100,
         keyinput_g101, keyinput_g102, keyinput_g103, keyinput_g104,
         keyinput_g105, keyinput_g106, keyinput_g107, keyinput_g108,
         keyinput_g109, keyinput_g110, keyinput_g111, keyinput_g112,
         keyinput_g113, keyinput_g114, keyinput_g115, keyinput_g116,
         keyinput_g117, keyinput_g118, keyinput_g119, keyinput_g120,
         keyinput_g121, keyinput_g122, keyinput_g123, keyinput_g124,
         keyinput_g125, keyinput_g126, keyinput_g127;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
         n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
         n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
         n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
         n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
         n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
         n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
         n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
         n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
         n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
         n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
         n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
         n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
         n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
         n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
         n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
         n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
         n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
         n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
         n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
         n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
         n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424,
         n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
         n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
         n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
         n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
         n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
         n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
         n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
         n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
         n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
         n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
         n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
         n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
         n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
         n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
         n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
         n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
         n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
         n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
         n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
         n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
         n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
         n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644,
         n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
         n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664,
         n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674,
         n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684,
         n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
         n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
         n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
         n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
         n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
         n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744,
         n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
         n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764,
         n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
         n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
         n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
         n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
         n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
         n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
         n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
         n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
         n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854,
         n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864,
         n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874,
         n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884,
         n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894,
         n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904,
         n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914,
         n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924,
         n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
         n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
         n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
         n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
         n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
         n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
         n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
         n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004,
         n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014,
         n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024,
         n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034,
         n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044,
         n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
         n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
         n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
         n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084,
         n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094,
         n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104,
         n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114,
         n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124,
         n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134,
         n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144,
         n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
         n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164,
         n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
         n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184,
         n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194,
         n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204,
         n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214,
         n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224,
         n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234,
         n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244,
         n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254,
         n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264,
         n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
         n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
         n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
         n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
         n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
         n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
         n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
         n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
         n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
         n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
         n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
         n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
         n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
         n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
         n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
         n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
         n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
         n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294,
         n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304,
         n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314,
         n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324,
         n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334,
         n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344,
         n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354,
         n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364,
         n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374,
         n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384,
         n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394,
         n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404,
         n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414,
         n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424,
         n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434,
         n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444,
         n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454,
         n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464,
         n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474,
         n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484,
         n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494,
         n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504,
         n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514,
         n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524,
         n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534,
         n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544,
         n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554,
         n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564,
         n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574,
         n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584,
         n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594,
         n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604,
         n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614,
         n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624,
         n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634,
         n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644,
         n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654,
         n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664,
         n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674,
         n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684,
         n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694,
         n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704,
         n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714,
         n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724,
         n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734,
         n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744,
         n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754,
         n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764,
         n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774,
         n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784,
         n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794,
         n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804,
         n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814,
         n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824,
         n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834,
         n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844,
         n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854,
         n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864,
         n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874,
         n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884,
         n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894,
         n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904,
         n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914,
         n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924,
         n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934,
         n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944,
         n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954,
         n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964,
         n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974,
         n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984,
         n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994,
         n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004,
         n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014,
         n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024,
         n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034,
         n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044,
         n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054,
         n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064,
         n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074,
         n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084,
         n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094,
         n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104,
         n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114,
         n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124,
         n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134,
         n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144,
         n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154,
         n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164,
         n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174,
         n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184,
         n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194,
         n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204,
         n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214,
         n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224,
         n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234,
         n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244,
         n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254,
         n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264,
         n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274,
         n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284,
         n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294,
         n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304,
         n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314,
         n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324,
         n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334,
         n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344,
         n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354,
         n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364,
         n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
         n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
         n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
         n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
         n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414,
         n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
         n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434,
         n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444,
         n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454,
         n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
         n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
         n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484,
         n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494,
         n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504,
         n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514,
         n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
         n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
         n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
         n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
         n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
         n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
         n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
         n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
         n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
         n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
         n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624,
         n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634,
         n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644,
         n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654,
         n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664,
         n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674,
         n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684,
         n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694,
         n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704,
         n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714,
         n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724,
         n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734,
         n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744,
         n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754,
         n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764,
         n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774,
         n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784,
         n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794,
         n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804,
         n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814,
         n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824,
         n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834,
         n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844,
         n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854,
         n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864,
         n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874,
         n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884,
         n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894,
         n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904,
         n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914,
         n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924,
         n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934,
         n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944,
         n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954,
         n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964,
         n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974,
         n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984,
         n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994,
         n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004,
         n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014,
         n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024,
         n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034,
         n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044,
         n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054,
         n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064,
         n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074,
         n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084,
         n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094,
         n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104,
         n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114,
         n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124,
         n7125;

  NAND2_X1 U3603 ( .A1(n3575), .A2(n3574), .ZN(n3675) );
  INV_X2 U3604 ( .A(n5665), .ZN(n5344) );
  CLKBUF_X2 U3605 ( .A(n3414), .Z(n3545) );
  CLKBUF_X2 U3606 ( .A(n3536), .Z(n4149) );
  CLKBUF_X2 U3607 ( .A(n3521), .Z(n4151) );
  CLKBUF_X2 U3608 ( .A(n3519), .Z(n4140) );
  BUF_X1 U3609 ( .A(n3474), .Z(n4324) );
  CLKBUF_X2 U3610 ( .A(n3537), .Z(n3158) );
  INV_X1 U3611 ( .A(n3482), .ZN(n4498) );
  CLKBUF_X2 U3612 ( .A(n3547), .Z(n4150) );
  CLKBUF_X2 U3613 ( .A(n3415), .Z(n4148) );
  CLKBUF_X2 U3614 ( .A(n3413), .Z(n4098) );
  CLKBUF_X2 U3615 ( .A(n3518), .Z(n4143) );
  BUF_X1 U3616 ( .A(n3427), .Z(n3421) );
  INV_X1 U3617 ( .A(n3498), .ZN(n4503) );
  INV_X1 U3618 ( .A(n3423), .ZN(n3428) );
  CLKBUF_X1 U3619 ( .A(n6705), .Z(n3155) );
  NOR2_X1 U3620 ( .A1(n7123), .A2(n6093), .ZN(n6705) );
  XNOR2_X1 U3621 ( .A(n3698), .B(n3707), .ZN(n4517) );
  AND4_X1 U3622 ( .A1(n3195), .A2(n3194), .A3(n3193), .A4(n3192), .ZN(n3211)
         );
  NAND4_X2 U3623 ( .A1(n3211), .A2(n3210), .A3(n3209), .A4(n3208), .ZN(n3482)
         );
  AND2_X2 U3624 ( .A1(n3451), .A2(n3482), .ZN(n6240) );
  OR3_X1 U3625 ( .A1(n6721), .A2(n6639), .A3(n3438), .ZN(n5267) );
  AND2_X2 U3626 ( .A1(n5517), .A2(n5504), .ZN(n5506) );
  NAND2_X1 U3627 ( .A1(n5609), .A2(n5610), .ZN(n5678) );
  OR2_X1 U3628 ( .A1(n4225), .A2(n4224), .ZN(n4227) );
  NOR2_X1 U3629 ( .A1(n5725), .A2(n5419), .ZN(n5421) );
  NAND2_X1 U3630 ( .A1(n5287), .A2(n5286), .ZN(n5389) );
  AOI21_X1 U3631 ( .B1(n5499), .B2(n7100), .A(n5498), .ZN(n5500) );
  INV_X1 U3632 ( .A(n6193), .ZN(n6186) );
  AND2_X1 U3633 ( .A1(n5794), .A2(n5411), .ZN(n3156) );
  NOR2_X2 U3634 ( .A1(n5543), .A2(n5545), .ZN(n5529) );
  AOI21_X2 U3635 ( .B1(n5730), .B2(n6354), .A(n5729), .ZN(n5731) );
  NOR2_X2 U3636 ( .A1(n5741), .A2(n5761), .ZN(n5754) );
  OAI21_X2 U3637 ( .B1(n5389), .B2(n5392), .A(n5390), .ZN(n5361) );
  XNOR2_X2 U3638 ( .A(n3573), .B(n3571), .ZN(n3619) );
  NAND2_X1 U3639 ( .A1(n3405), .A2(n3463), .ZN(n3461) );
  XNOR2_X1 U3640 ( .A(n5421), .B(n5420), .ZN(n5456) );
  OR2_X1 U3641 ( .A1(n5822), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5823)
         );
  OAI21_X1 U3642 ( .B1(n5445), .B2(n6391), .A(n5450), .ZN(n5446) );
  NAND2_X1 U3643 ( .A1(n5568), .A2(n5570), .ZN(n5569) );
  NAND2_X1 U3644 ( .A1(n5114), .A2(n5143), .ZN(n5145) );
  NOR2_X1 U3645 ( .A1(n5655), .A2(n5654), .ZN(n3287) );
  AND2_X1 U3646 ( .A1(n4545), .A2(n4544), .ZN(n3726) );
  NAND2_X1 U3647 ( .A1(n3731), .A2(n3730), .ZN(n4796) );
  NAND2_X2 U3648 ( .A1(n5698), .A2(n4325), .ZN(n6024) );
  XNOR2_X1 U3649 ( .A(n3603), .B(n3602), .ZN(n3651) );
  NAND2_X1 U3650 ( .A1(n3599), .A2(n3598), .ZN(n3603) );
  CLKBUF_X1 U3651 ( .A(n4367), .Z(n6189) );
  NOR2_X1 U3652 ( .A1(n4266), .A2(n3509), .ZN(n3529) );
  CLKBUF_X1 U3653 ( .A(n3480), .Z(n5480) );
  NOR2_X1 U3654 ( .A1(n4200), .A2(n4498), .ZN(n3480) );
  AND2_X1 U3655 ( .A1(n3234), .A2(n3233), .ZN(n4401) );
  CLKBUF_X1 U3656 ( .A(n4200), .Z(n4352) );
  INV_X1 U3657 ( .A(n3734), .ZN(n3709) );
  OAI21_X1 U3658 ( .B1(n3473), .B2(n3472), .A(n4498), .ZN(n3476) );
  NAND2_X1 U3659 ( .A1(n3226), .A2(n3225), .ZN(n3230) );
  AOI21_X1 U3660 ( .B1(n3838), .B2(n3461), .A(n4503), .ZN(n3473) );
  INV_X1 U3661 ( .A(n3236), .ZN(n3157) );
  NAND2_X1 U3662 ( .A1(n4306), .A2(n5665), .ZN(n3301) );
  OR2_X1 U3663 ( .A1(n3543), .A2(n3542), .ZN(n4800) );
  NAND2_X1 U3664 ( .A1(n3174), .A2(n3341), .ZN(n3427) );
  AND4_X1 U3665 ( .A1(n3203), .A2(n3202), .A3(n3201), .A4(n3200), .ZN(n3209)
         );
  AND4_X1 U3666 ( .A1(n3207), .A2(n3206), .A3(n3205), .A4(n3204), .ZN(n3208)
         );
  AND4_X1 U3667 ( .A1(n3340), .A2(n3339), .A3(n3338), .A4(n3337), .ZN(n3341)
         );
  AND4_X1 U3668 ( .A1(n3215), .A2(n3214), .A3(n3213), .A4(n3212), .ZN(n3221)
         );
  AND4_X1 U3669 ( .A1(n3312), .A2(n3311), .A3(n3310), .A4(n3309), .ZN(n3318)
         );
  BUF_X1 U3670 ( .A(n3772), .Z(n3773) );
  AND4_X1 U3671 ( .A1(n3316), .A2(n3315), .A3(n3314), .A4(n3313), .ZN(n3317)
         );
  NAND2_X2 U3672 ( .A1(STATE_REG_2__SCAN_IN), .A2(n7123), .ZN(n6696) );
  BUF_X2 U3673 ( .A(n3544), .Z(n4139) );
  AND2_X2 U3674 ( .A1(n6644), .A2(n4474), .ZN(n4333) );
  BUF_X2 U3675 ( .A(n3408), .Z(n4142) );
  NAND2_X1 U3676 ( .A1(n4249), .A2(n4294), .ZN(n3462) );
  INV_X2 U3677 ( .A(n4294), .ZN(n4508) );
  AND4_X2 U3678 ( .A1(n3190), .A2(n3189), .A3(n3188), .A4(n3187), .ZN(n3191)
         );
  NAND2_X1 U3679 ( .A1(n5794), .A2(n5411), .ZN(n3159) );
  CLKBUF_X1 U3680 ( .A(n6327), .Z(n3160) );
  NAND2_X1 U3681 ( .A1(n6343), .A2(n3164), .ZN(n3161) );
  OAI21_X1 U3683 ( .B1(n3467), .B2(n3426), .A(n5696), .ZN(n3163) );
  XNOR2_X1 U3684 ( .A(n4431), .B(n6417), .ZN(n3164) );
  NAND2_X1 U3685 ( .A1(n5794), .A2(n5411), .ZN(n5822) );
  OAI21_X1 U3686 ( .B1(n3467), .B2(n3426), .A(n5696), .ZN(n3472) );
  AND2_X1 U3687 ( .A1(n3428), .A2(n3464), .ZN(n3426) );
  AND2_X2 U3688 ( .A1(n5340), .A2(n3981), .ZN(n5568) );
  NAND3_X1 U3689 ( .A1(n3675), .A2(n4482), .A3(n3674), .ZN(n3705) );
  AND2_X2 U3691 ( .A1(n3186), .A2(n4357), .ZN(n3414) );
  AND2_X4 U3692 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4368) );
  NOR3_X2 U3693 ( .A1(n5678), .A2(n5677), .A3(n5676), .ZN(n3275) );
  AND2_X1 U3694 ( .A1(n3186), .A2(n4357), .ZN(n3165) );
  AND2_X2 U3695 ( .A1(n5081), .A2(n5115), .ZN(n5114) );
  NOR2_X4 U3696 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4369) );
  INV_X2 U3697 ( .A(n4249), .ZN(n3451) );
  OR2_X2 U3698 ( .A1(n6039), .A2(n5408), .ZN(n5794) );
  NOR2_X2 U3699 ( .A1(n5069), .A2(n5070), .ZN(n5093) );
  OR2_X2 U3700 ( .A1(n4770), .A2(n4703), .ZN(n5069) );
  BUF_X4 U3701 ( .A(n3462), .Z(n5665) );
  AND2_X1 U3702 ( .A1(n5696), .A2(n4294), .ZN(n3465) );
  OR2_X1 U3703 ( .A1(n3474), .A2(n3464), .ZN(n3466) );
  INV_X1 U3704 ( .A(n3729), .ZN(n3730) );
  INV_X1 U3705 ( .A(n3728), .ZN(n3731) );
  NAND2_X1 U3706 ( .A1(n3319), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3734) );
  INV_X1 U3707 ( .A(n3332), .ZN(n3319) );
  NOR2_X1 U3708 ( .A1(n3464), .A2(n6644), .ZN(n4797) );
  AND2_X2 U3709 ( .A1(n4463), .A2(n4368), .ZN(n3537) );
  NAND2_X1 U3710 ( .A1(n3482), .A2(n3464), .ZN(n3332) );
  AND2_X2 U3711 ( .A1(n3186), .A2(n4368), .ZN(n3520) );
  AND2_X1 U3712 ( .A1(n5479), .A2(n6641), .ZN(n6238) );
  NAND2_X1 U3713 ( .A1(n3173), .A2(n3470), .ZN(n3471) );
  AOI22_X1 U3714 ( .A1(n3544), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3414), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3338) );
  OR2_X1 U3715 ( .A1(n3344), .A2(n3345), .ZN(n3322) );
  CLKBUF_X1 U3716 ( .A(n3512), .Z(n3772) );
  NAND2_X1 U3717 ( .A1(n3500), .A2(n3499), .ZN(n4266) );
  OR2_X1 U3718 ( .A1(n3734), .A2(n4290), .ZN(n3372) );
  AND2_X1 U3719 ( .A1(n3331), .A2(n3330), .ZN(n3434) );
  NAND2_X1 U3720 ( .A1(n3586), .A2(n3585), .ZN(n3631) );
  AND2_X1 U3722 ( .A1(n3979), .A2(n5342), .ZN(n5649) );
  XNOR2_X1 U3724 ( .A(n4796), .B(n3735), .ZN(n4783) );
  INV_X1 U3725 ( .A(n5348), .ZN(n4269) );
  NAND2_X1 U3726 ( .A1(n3636), .A2(n3635), .ZN(n4922) );
  INV_X1 U3727 ( .A(n3372), .ZN(n3380) );
  AND2_X1 U3728 ( .A1(n4268), .A2(n3484), .ZN(n4350) );
  INV_X1 U3729 ( .A(n3820), .ZN(n4039) );
  OR2_X1 U3730 ( .A1(n4116), .A2(n5746), .ZN(n4117) );
  OR2_X1 U3731 ( .A1(n4117), .A2(n5494), .ZN(n4171) );
  NOR2_X1 U3732 ( .A1(n3736), .A2(n5260), .ZN(n3737) );
  AND2_X1 U3733 ( .A1(n4248), .A2(n6641), .ZN(n4276) );
  INV_X1 U3734 ( .A(n3617), .ZN(n3618) );
  AND2_X2 U3735 ( .A1(n3318), .A2(n3317), .ZN(n4582) );
  AND2_X1 U3736 ( .A1(n5267), .A2(n4185), .ZN(n6193) );
  AND2_X1 U3737 ( .A1(n5728), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4185) );
  AND2_X1 U3738 ( .A1(n5698), .A2(n5697), .ZN(n6214) );
  INV_X1 U3739 ( .A(n5698), .ZN(n6213) );
  NAND2_X1 U3740 ( .A1(n6096), .A2(n4233), .ZN(n6047) );
  AOI22_X1 U3741 ( .A1(n3415), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3536), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3337) );
  AND2_X1 U3742 ( .A1(n3324), .A2(n3323), .ZN(n3361) );
  INV_X1 U3743 ( .A(n3705), .ZN(n3708) );
  AND2_X1 U3744 ( .A1(n3722), .A2(n3721), .ZN(n3729) );
  OR2_X1 U3745 ( .A1(n3696), .A2(n3695), .ZN(n4564) );
  OR2_X1 U3746 ( .A1(n3662), .A2(n3661), .ZN(n4565) );
  NAND2_X1 U3747 ( .A1(n3709), .A2(n4324), .ZN(n3478) );
  AOI22_X1 U3748 ( .A1(n3413), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3537), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3216) );
  AND2_X1 U3749 ( .A1(n3980), .A2(n5649), .ZN(n3981) );
  AND2_X1 U3750 ( .A1(n5811), .A2(n5812), .ZN(n5781) );
  OR2_X1 U3751 ( .A1(n3560), .A2(n3559), .ZN(n4292) );
  AND2_X1 U3752 ( .A1(n3607), .A2(n3606), .ZN(n3566) );
  OR2_X1 U3753 ( .A1(n3647), .A2(n3646), .ZN(n4434) );
  XNOR2_X1 U3754 ( .A(n3630), .B(n3587), .ZN(n4450) );
  XNOR2_X1 U3755 ( .A(n4384), .B(n4922), .ZN(n4367) );
  OR3_X1 U3756 ( .A1(n4347), .A2(n4346), .A3(n4345), .ZN(n6614) );
  AND2_X1 U3757 ( .A1(n3633), .A2(n4911), .ZN(n5020) );
  AND4_X1 U3758 ( .A1(n3199), .A2(n3198), .A3(n3197), .A4(n3196), .ZN(n3210)
         );
  INV_X1 U3759 ( .A(n6637), .ZN(n4472) );
  INV_X1 U3760 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4681) );
  INV_X1 U3761 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6620) );
  AND2_X2 U3762 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4463) );
  OR2_X1 U3763 ( .A1(n5481), .A2(n6648), .ZN(n4205) );
  OR2_X1 U3764 ( .A1(n3436), .A2(n3435), .ZN(n5469) );
  CLKBUF_X1 U3765 ( .A(n3481), .Z(n5476) );
  INV_X1 U3766 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n5260) );
  NAND2_X1 U3767 ( .A1(n3630), .A2(n3631), .ZN(n4384) );
  INV_X1 U3768 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n5166) );
  CLKBUF_X1 U3769 ( .A(n3482), .Z(n3348) );
  AND2_X1 U3770 ( .A1(n6238), .A2(n4202), .ZN(n6217) );
  NOR2_X1 U3771 ( .A1(n4078), .A2(n5765), .ZN(n4079) );
  BUF_X1 U3772 ( .A(n5514), .Z(n5530) );
  OR2_X1 U3773 ( .A1(n4044), .A2(n5553), .ZN(n4078) );
  CLKBUF_X1 U3774 ( .A(n5529), .Z(n5544) );
  CLKBUF_X1 U3776 ( .A(n5568), .Z(n5652) );
  AND2_X1 U3777 ( .A1(PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n3855), .ZN(n3893)
         );
  NAND2_X1 U3778 ( .A1(n3893), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3892)
         );
  NAND2_X1 U3779 ( .A1(n3958), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n3957)
         );
  NOR2_X1 U3780 ( .A1(n3926), .A2(n3927), .ZN(n3912) );
  OR2_X1 U3781 ( .A1(n5622), .A2(n5381), .ZN(n5673) );
  OR2_X1 U3782 ( .A1(n5849), .A2(n5848), .ZN(n5365) );
  AND2_X1 U3783 ( .A1(n5849), .A2(n5848), .ZN(n5366) );
  NAND2_X1 U3784 ( .A1(n3972), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3926)
         );
  NAND2_X1 U3785 ( .A1(n5650), .A2(n5620), .ZN(n5622) );
  NAND2_X1 U3786 ( .A1(n3819), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3854)
         );
  NOR2_X1 U3787 ( .A1(n3805), .A2(n3804), .ZN(n3819) );
  NOR2_X1 U3788 ( .A1(n3771), .A2(n5240), .ZN(n3788) );
  NAND2_X1 U3790 ( .A1(n3755), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3771)
         );
  INV_X1 U3791 ( .A(n3741), .ZN(n3755) );
  AOI21_X1 U3792 ( .B1(n4783), .B2(n3961), .A(n3740), .ZN(n4707) );
  CLKBUF_X1 U3793 ( .A(n4699), .Z(n4705) );
  NAND2_X1 U3794 ( .A1(n3699), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3736)
         );
  AND2_X1 U3795 ( .A1(n4406), .A2(n4479), .ZN(n3685) );
  NOR2_X1 U3796 ( .A1(n3677), .A2(n5166), .ZN(n3699) );
  INV_X1 U3797 ( .A(n3667), .ZN(n3678) );
  NAND2_X1 U3798 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3667) );
  AND2_X2 U3799 ( .A1(n5506), .A2(n5488), .ZN(n4180) );
  NOR2_X2 U3800 ( .A1(n5657), .A2(n5571), .ZN(n5923) );
  INV_X1 U3801 ( .A(n5781), .ZN(n5810) );
  AND2_X1 U3802 ( .A1(n5626), .A2(n5625), .ZN(n5609) );
  AND2_X1 U3803 ( .A1(n4276), .A2(n4271), .ZN(n6070) );
  NOR2_X2 U3804 ( .A1(n5274), .A2(n5275), .ZN(n5626) );
  OAI21_X1 U3805 ( .B1(n5158), .B2(n5284), .A(n5283), .ZN(n5285) );
  AND2_X1 U3806 ( .A1(n3261), .A2(n3260), .ZN(n5118) );
  AND2_X1 U3807 ( .A1(n5093), .A2(n5092), .ZN(n5091) );
  CLKBUF_X1 U3808 ( .A(n5156), .Z(n5074) );
  NAND2_X1 U3809 ( .A1(n3251), .A2(n3250), .ZN(n4770) );
  INV_X1 U3810 ( .A(n4767), .ZN(n3250) );
  INV_X1 U3811 ( .A(n4768), .ZN(n3251) );
  NAND2_X1 U3812 ( .A1(n4549), .A2(n4548), .ZN(n4768) );
  NAND2_X1 U3813 ( .A1(n3243), .A2(n3242), .ZN(n4537) );
  INV_X1 U3814 ( .A(n4408), .ZN(n3242) );
  NAND2_X1 U3815 ( .A1(n5194), .A2(n4306), .ZN(n4311) );
  INV_X1 U3816 ( .A(n6426), .ZN(n6399) );
  OR2_X1 U3817 ( .A1(n6073), .A2(n6070), .ZN(n4534) );
  INV_X1 U3818 ( .A(n3651), .ZN(n3674) );
  AND2_X2 U3819 ( .A1(n3177), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4358)
         );
  INV_X1 U3820 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4360) );
  CLKBUF_X1 U3821 ( .A(n4450), .Z(n5134) );
  INV_X1 U3822 ( .A(n6614), .ZN(n4467) );
  OR2_X1 U3823 ( .A1(n5986), .A2(n5978), .ZN(n4977) );
  INV_X1 U3824 ( .A(n4920), .ZN(n4976) );
  NAND2_X1 U3825 ( .A1(n6644), .A2(n4492), .ZN(n4646) );
  AND2_X1 U3826 ( .A1(n5981), .A2(n4591), .ZN(n4598) );
  AOI21_X1 U3827 ( .B1(n3384), .B2(n3383), .A(n3382), .ZN(n5479) );
  NOR2_X1 U3828 ( .A1(n3381), .A2(n3733), .ZN(n3382) );
  NAND2_X1 U3829 ( .A1(n4196), .A2(n4195), .ZN(n4197) );
  AND2_X1 U3830 ( .A1(REIP_REG_18__SCAN_IN), .A2(n5582), .ZN(n6012) );
  INV_X1 U3831 ( .A(n6123), .ZN(n6191) );
  OR2_X1 U3832 ( .A1(n5127), .A2(n3439), .ZN(n6198) );
  INV_X1 U3833 ( .A(n6044), .ZN(n6207) );
  NAND2_X1 U3834 ( .A1(n4323), .A2(n6272), .ZN(n5698) );
  INV_X1 U3835 ( .A(n5720), .ZN(n5291) );
  BUF_X1 U3836 ( .A(n6234), .Z(n6229) );
  CLKBUF_X2 U3837 ( .A(n6317), .Z(n6321) );
  XNOR2_X1 U3838 ( .A(n4172), .B(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5728)
         );
  AOI21_X1 U3839 ( .B1(n5662), .B2(n5661), .A(n5660), .ZN(n6032) );
  OAI21_X1 U3840 ( .B1(n5588), .B2(n5343), .A(n5661), .ZN(n6035) );
  BUF_X1 U3841 ( .A(n5847), .Z(n5851) );
  NAND2_X1 U3842 ( .A1(n6047), .A2(n4300), .ZN(n6360) );
  INV_X1 U3843 ( .A(n6047), .ZN(n6350) );
  INV_X1 U3844 ( .A(n5898), .ZN(n5914) );
  NOR2_X1 U3845 ( .A1(n5439), .A2(n6057), .ZN(n6052) );
  AND2_X1 U3846 ( .A1(n4276), .A2(n4273), .ZN(n6424) );
  NOR2_X1 U3847 ( .A1(n4534), .A2(n6399), .ZN(n5438) );
  AND2_X1 U3848 ( .A1(n4276), .A2(n5355), .ZN(n6073) );
  INV_X1 U3849 ( .A(n6424), .ZN(n6391) );
  AND2_X1 U3850 ( .A1(n4276), .A2(n4256), .ZN(n6429) );
  CLKBUF_X1 U3851 ( .A(n4481), .Z(n5978) );
  CLKBUF_X1 U3852 ( .A(n4348), .Z(n4349) );
  CLKBUF_X1 U3853 ( .A(n4483), .Z(n5981) );
  AND2_X1 U3854 ( .A1(n5978), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6438) );
  INV_X1 U3855 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n5467) );
  NOR2_X1 U3856 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_1__SCAN_IN), .ZN(
        n5463) );
  OR2_X1 U3857 ( .A1(n5203), .A2(n5292), .ZN(n6476) );
  OR2_X1 U3858 ( .A1(n5986), .A2(n4921), .ZN(n6525) );
  OR3_X1 U3859 ( .A1(n6532), .A2(n4920), .A3(n5978), .ZN(n4874) );
  INV_X1 U3860 ( .A(n5060), .ZN(n5032) );
  OR2_X1 U3861 ( .A1(n6532), .A2(n5292), .ZN(n6592) );
  AND2_X1 U3862 ( .A1(n5479), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6637) );
  INV_X1 U3863 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n6645) );
  AND2_X1 U3864 ( .A1(n6635), .A2(n6634), .ZN(n6706) );
  CLKBUF_X1 U3865 ( .A(n6700), .Z(n6697) );
  INV_X1 U3866 ( .A(n5701), .ZN(n5454) );
  INV_X1 U3867 ( .A(n3227), .ZN(n3236) );
  INV_X2 U3868 ( .A(n3535), .ZN(n3546) );
  NOR2_X1 U3869 ( .A1(n3463), .A2(n3462), .ZN(n3166) );
  AND2_X2 U3870 ( .A1(n4369), .A2(n4368), .ZN(n3553) );
  NAND2_X1 U3872 ( .A1(n3580), .A2(n3579), .ZN(n3630) );
  INV_X1 U3873 ( .A(n3224), .ZN(n4306) );
  INV_X1 U3874 ( .A(n4554), .ZN(n3243) );
  AND3_X1 U3875 ( .A1(n5791), .A2(n5954), .A3(n5443), .ZN(n3167) );
  INV_X1 U3876 ( .A(n5158), .ZN(n5277) );
  AND2_X1 U3877 ( .A1(n3506), .A2(n3505), .ZN(n3168) );
  INV_X2 U3878 ( .A(n5277), .ZN(n5849) );
  NAND2_X1 U3879 ( .A1(n4796), .A2(n4798), .ZN(n5158) );
  AND2_X1 U3880 ( .A1(n3707), .A2(n3706), .ZN(n3169) );
  AND3_X1 U3881 ( .A1(n4929), .A2(n4928), .A3(n4927), .ZN(n3170) );
  INV_X1 U3882 ( .A(n6157), .ZN(n6171) );
  INV_X1 U3883 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4447) );
  OR2_X1 U3884 ( .A1(n3491), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3171)
         );
  NAND2_X1 U3885 ( .A1(n5921), .A2(n5561), .ZN(n5549) );
  AND2_X2 U3886 ( .A1(n3179), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4357)
         );
  AND4_X1 U3887 ( .A1(n3184), .A2(n3183), .A3(n3182), .A4(n3181), .ZN(n3172)
         );
  OR2_X1 U3888 ( .A1(n4249), .A2(n3469), .ZN(n3173) );
  INV_X1 U3889 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5420) );
  AND4_X1 U3890 ( .A1(n3336), .A2(n3335), .A3(n3334), .A4(n3333), .ZN(n3174)
         );
  AND4_X1 U3891 ( .A1(n3412), .A2(n3411), .A3(n3410), .A4(n3409), .ZN(n3175)
         );
  AND2_X2 U3892 ( .A1(n4699), .A2(n4698), .ZN(n3176) );
  NAND2_X1 U3893 ( .A1(n5692), .A2(n6023), .ZN(n5689) );
  INV_X1 U3894 ( .A(n5068), .ZN(n3770) );
  AOI21_X1 U3895 ( .B1(n4220), .B2(n4324), .A(n4203), .ZN(n3475) );
  NAND2_X1 U3896 ( .A1(n4797), .A2(n4415), .ZN(n3598) );
  OR2_X1 U3897 ( .A1(n3719), .A2(n3718), .ZN(n4785) );
  INV_X1 U3898 ( .A(n3427), .ZN(n3424) );
  OR2_X1 U3899 ( .A1(n3527), .A2(n3526), .ZN(n4291) );
  INV_X1 U3900 ( .A(n4800), .ZN(n3732) );
  AND2_X1 U3901 ( .A1(n4307), .A2(n4294), .ZN(n3422) );
  OR2_X1 U3902 ( .A1(n3597), .A2(n3596), .ZN(n4415) );
  NAND2_X1 U3903 ( .A1(n3428), .A2(n5696), .ZN(n3838) );
  NAND2_X1 U3904 ( .A1(n3675), .A2(n3674), .ZN(n3676) );
  AND4_X1 U3905 ( .A1(n3402), .A2(n3401), .A3(n3400), .A4(n3399), .ZN(n3403)
         );
  AND4_X1 U3906 ( .A1(n3219), .A2(n3218), .A3(n3217), .A4(n3216), .ZN(n3220)
         );
  MUX2_X1 U3907 ( .A(n3462), .B(n3227), .S(EBX_REG_1__SCAN_IN), .Z(n3226) );
  AND2_X1 U3908 ( .A1(n3483), .A2(n4508), .ZN(n4268) );
  AND2_X1 U3909 ( .A1(n4021), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4022)
         );
  INV_X1 U3910 ( .A(n3957), .ZN(n3855) );
  OR2_X1 U3911 ( .A1(n5145), .A2(n3836), .ZN(n5619) );
  OR2_X1 U3912 ( .A1(n5696), .A2(n6636), .ZN(n4020) );
  OR2_X1 U3913 ( .A1(n5849), .A2(n5410), .ZN(n5411) );
  INV_X1 U3914 ( .A(n3631), .ZN(n3587) );
  NAND2_X1 U3915 ( .A1(n3332), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3733) );
  NAND2_X1 U3916 ( .A1(n4367), .A2(n6644), .ZN(n3650) );
  AND4_X1 U3917 ( .A1(n3419), .A2(n3418), .A3(n3417), .A4(n3416), .ZN(n3420)
         );
  AND2_X1 U3918 ( .A1(n3565), .A2(n4797), .ZN(n3606) );
  AND2_X1 U3919 ( .A1(n4498), .A2(n4249), .ZN(n4203) );
  AND2_X1 U3920 ( .A1(n3379), .A2(n3378), .ZN(n3436) );
  INV_X1 U3921 ( .A(n6181), .ZN(n5237) );
  AND2_X1 U3922 ( .A1(n3241), .A2(n3240), .ZN(n4408) );
  NOR2_X1 U3923 ( .A1(n3498), .A2(n3421), .ZN(n4307) );
  NAND2_X1 U3924 ( .A1(n3428), .A2(n3427), .ZN(n3474) );
  NOR2_X1 U3925 ( .A1(n4171), .A2(n5452), .ZN(n4172) );
  NAND2_X1 U3926 ( .A1(n4022), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4042)
         );
  AND2_X1 U3927 ( .A1(n3912), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3958)
         );
  NOR2_X1 U3928 ( .A1(n3854), .A2(n3853), .ZN(n3972) );
  NAND2_X1 U3929 ( .A1(n3788), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3805)
         );
  NAND2_X1 U3930 ( .A1(n4582), .A2(n3427), .ZN(n3463) );
  OR2_X1 U3931 ( .A1(n5925), .A2(n5435), .ZN(n5898) );
  AND2_X1 U3932 ( .A1(n5849), .A2(n5407), .ZN(n5408) );
  INV_X1 U3933 ( .A(n5285), .ZN(n5286) );
  NAND2_X1 U3934 ( .A1(n4414), .A2(n4413), .ZN(n6351) );
  XNOR2_X1 U3935 ( .A(n3511), .B(n3510), .ZN(n4348) );
  OAI21_X1 U3936 ( .B1(n5220), .B2(n6709), .A(n5214), .ZN(n5252) );
  NAND2_X1 U3937 ( .A1(n3650), .A2(n3649), .ZN(n4482) );
  AND2_X1 U3938 ( .A1(n4680), .A2(n6530), .ZN(n4685) );
  INV_X1 U3939 ( .A(n4646), .ZN(n5022) );
  XNOR2_X1 U3940 ( .A(n3675), .B(n3651), .ZN(n4483) );
  AND2_X1 U3941 ( .A1(n4343), .A2(n4258), .ZN(n5473) );
  NOR2_X1 U3942 ( .A1(n3892), .A2(n5819), .ZN(n3856) );
  INV_X1 U3943 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n5240) );
  INV_X1 U3944 ( .A(n6194), .ZN(n6176) );
  OR2_X1 U3945 ( .A1(n5127), .A2(n3441), .ZN(n6181) );
  INV_X1 U3946 ( .A(n3275), .ZN(n5679) );
  INV_X1 U3947 ( .A(n4163), .ZN(n4165) );
  NAND2_X1 U3948 ( .A1(n4079), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4116)
         );
  AND2_X1 U3949 ( .A1(n5343), .A2(n5341), .ZN(n5342) );
  OR2_X1 U3950 ( .A1(n5622), .A2(n5608), .ZN(n5606) );
  AND2_X1 U3951 ( .A1(n5741), .A2(n5418), .ZN(n5419) );
  AOI21_X1 U3952 ( .B1(n5817), .B2(n5816), .A(n5780), .ZN(n5811) );
  OR2_X1 U3953 ( .A1(n5422), .A2(n6367), .ZN(n6057) );
  NAND2_X1 U3954 ( .A1(n5091), .A2(n5118), .ZN(n5148) );
  OR2_X1 U3955 ( .A1(n5158), .A2(n5084), .ZN(n5283) );
  AND2_X1 U3956 ( .A1(n4528), .A2(n4527), .ZN(n5373) );
  AND2_X1 U3957 ( .A1(n4413), .A2(n4289), .ZN(n4411) );
  OAI21_X1 U3958 ( .B1(n6724), .B2(n4474), .A(n4472), .ZN(n4492) );
  OR2_X1 U3959 ( .A1(n4977), .A2(n4920), .ZN(n5009) );
  XNOR2_X1 U3960 ( .A(n3619), .B(n3618), .ZN(n4481) );
  INV_X1 U3961 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4929) );
  OR2_X1 U3962 ( .A1(n3609), .A2(n3608), .ZN(n4217) );
  AND2_X1 U3963 ( .A1(n6645), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3493) );
  AND2_X1 U3964 ( .A1(n3856), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n4021)
         );
  NAND2_X1 U3965 ( .A1(n5267), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5127) );
  AND2_X1 U3966 ( .A1(n5267), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6194) );
  INV_X1 U3967 ( .A(n6198), .ZN(n6153) );
  INV_X1 U3968 ( .A(n6165), .ZN(n6178) );
  OAI22_X1 U3969 ( .A1(n4179), .A2(n5344), .B1(n5489), .B2(n4182), .ZN(n5493)
         );
  INV_X1 U3970 ( .A(n5689), .ZN(n6018) );
  NAND2_X1 U3971 ( .A1(n3157), .A2(n5665), .ZN(n4275) );
  AND2_X1 U3972 ( .A1(n5698), .A2(n4326), .ZN(n5720) );
  NOR2_X1 U3973 ( .A1(n4333), .A2(n6217), .ZN(n6234) );
  AOI21_X1 U3974 ( .B1(n5383), .B2(n5606), .A(n5382), .ZN(n6212) );
  NAND2_X1 U3975 ( .A1(n3678), .A2(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3677)
         );
  INV_X1 U3976 ( .A(n6096), .ZN(n6356) );
  AND2_X1 U3977 ( .A1(n5905), .A2(n5444), .ZN(n5893) );
  AND2_X1 U3978 ( .A1(n5930), .A2(n5443), .ZN(n5905) );
  OAI21_X1 U3979 ( .B1(n5277), .B2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n5810), 
        .ZN(n5803) );
  AND2_X1 U3980 ( .A1(n5823), .A2(n5779), .ZN(n5817) );
  CLKBUF_X1 U3981 ( .A(n4782), .Z(n4562) );
  AND2_X1 U3982 ( .A1(n4534), .A2(n4533), .ZN(n6419) );
  INV_X1 U3983 ( .A(n4850), .ZN(n4843) );
  NOR2_X1 U3984 ( .A1(n5203), .A2(n5978), .ZN(n4624) );
  AND2_X1 U3985 ( .A1(n4624), .A2(n4976), .ZN(n4759) );
  OR2_X1 U3986 ( .A1(n4424), .A2(n5981), .ZN(n5203) );
  INV_X1 U3987 ( .A(n6476), .ZN(n5257) );
  INV_X1 U3988 ( .A(n5009), .ZN(n4966) );
  INV_X1 U3989 ( .A(n6516), .ZN(n6520) );
  NAND2_X1 U3990 ( .A1(n4424), .A2(n6439), .ZN(n6532) );
  AND2_X1 U3991 ( .A1(n4598), .A2(n4920), .ZN(n5338) );
  INV_X1 U3992 ( .A(n4861), .ZN(n4756) );
  AND2_X1 U3993 ( .A1(n4491), .A2(n5981), .ZN(n4914) );
  NAND2_X1 U3994 ( .A1(n4204), .A2(n4205), .ZN(n6721) );
  INV_X1 U3995 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6999) );
  NAND2_X1 U3996 ( .A1(n5730), .A2(n6171), .ZN(n4174) );
  OR2_X1 U3997 ( .A1(n5127), .A2(n4189), .ZN(n6123) );
  NAND2_X1 U3998 ( .A1(n5267), .A2(n4173), .ZN(n6157) );
  INV_X1 U3999 ( .A(n6020), .ZN(n5688) );
  XNOR2_X1 U4000 ( .A(n5486), .B(n4192), .ZN(n5701) );
  INV_X1 U4001 ( .A(n6217), .ZN(n6236) );
  OR2_X1 U4002 ( .A1(n5653), .A2(n5652), .ZN(n6028) );
  NAND2_X1 U4003 ( .A1(n6238), .A2(n6602), .ZN(n6096) );
  OR2_X1 U4004 ( .A1(n5968), .A2(n5441), .ZN(n5948) );
  INV_X1 U4005 ( .A(n6066), .ZN(n6367) );
  INV_X1 U4006 ( .A(n6429), .ZN(n6403) );
  INV_X1 U4007 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6610) );
  INV_X1 U4008 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n5359) );
  AND2_X1 U4009 ( .A1(n4814), .A2(n4813), .ZN(n4854) );
  INV_X1 U4010 ( .A(n4765), .ZN(n4679) );
  OR2_X1 U4011 ( .A1(n5203), .A2(n4921), .ZN(n6470) );
  OR2_X1 U4012 ( .A1(n4977), .A2(n4976), .ZN(n5259) );
  OR2_X1 U4013 ( .A1(n5986), .A2(n5292), .ZN(n6516) );
  OR3_X1 U4014 ( .A1(n6532), .A2(n4976), .A3(n5978), .ZN(n5060) );
  INV_X1 U4015 ( .A(n4871), .ZN(n4910) );
  OR2_X1 U4016 ( .A1(n6532), .A2(n4921), .ZN(n6599) );
  OR2_X1 U4017 ( .A1(n4592), .A2(n4920), .ZN(n4861) );
  AND3_X1 U4018 ( .A1(n4726), .A2(n4725), .A3(n4927), .ZN(n4855) );
  INV_X1 U4019 ( .A(n4858), .ZN(n4918) );
  INV_X1 U4020 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3177) );
  INV_X1 U4021 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3178) );
  AND2_X2 U4022 ( .A1(n3178), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3186)
         );
  AND2_X2 U4023 ( .A1(n4358), .A2(n3186), .ZN(n3544) );
  INV_X1 U4024 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3179) );
  AND2_X2 U4025 ( .A1(n4357), .A2(n4369), .ZN(n3521) );
  AOI22_X1 U4026 ( .A1(n3544), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3521), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3184) );
  AND2_X4 U4027 ( .A1(n4358), .A2(n4463), .ZN(n3513) );
  AND2_X2 U4028 ( .A1(n4358), .A2(n4369), .ZN(n3519) );
  AOI22_X1 U4029 ( .A1(n3513), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3519), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3183) );
  INV_X1 U4030 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3180) );
  AND2_X2 U4031 ( .A1(n3180), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3185)
         );
  AND2_X2 U4032 ( .A1(n4358), .A2(n3185), .ZN(n3547) );
  AND2_X2 U4033 ( .A1(n3185), .A2(n4368), .ZN(n3407) );
  AOI22_X1 U4034 ( .A1(n3547), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3407), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3182) );
  AND2_X2 U4035 ( .A1(n4357), .A2(n3185), .ZN(n3415) );
  NOR2_X4 U4036 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4466) );
  AOI22_X1 U4037 ( .A1(n3415), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3408), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3181) );
  AND2_X2 U4038 ( .A1(n3186), .A2(n4466), .ZN(n3512) );
  AOI22_X1 U4040 ( .A1(n3512), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3536), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3190) );
  AND2_X2 U4041 ( .A1(n4466), .A2(n4463), .ZN(n3413) );
  AOI22_X1 U4042 ( .A1(n3413), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3553), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3189) );
  AOI22_X1 U4043 ( .A1(n3414), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3537), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3188) );
  AND2_X2 U4044 ( .A1(n4357), .A2(n4463), .ZN(n3518) );
  AOI22_X1 U4045 ( .A1(n3518), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3520), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3187) );
  NAND2_X2 U4046 ( .A1(n3172), .A2(n3191), .ZN(n4294) );
  NAND2_X1 U4047 ( .A1(n3413), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3195)
         );
  NAND2_X1 U4048 ( .A1(n3518), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3194)
         );
  NAND2_X1 U4049 ( .A1(n3512), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3193) );
  NAND2_X1 U4050 ( .A1(n3414), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3192) );
  NAND2_X1 U4051 ( .A1(n3547), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3199)
         );
  NAND2_X1 U4052 ( .A1(n3513), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3198)
         );
  NAND2_X1 U4053 ( .A1(n3407), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3197)
         );
  NAND2_X1 U4054 ( .A1(n3520), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3196) );
  NAND2_X1 U4055 ( .A1(n3415), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3203) );
  NAND2_X1 U4056 ( .A1(n3519), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3202) );
  NAND2_X1 U4057 ( .A1(n3536), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3201) );
  NAND2_X1 U4058 ( .A1(n3408), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3200) );
  NAND2_X1 U4059 ( .A1(n3544), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3207) );
  NAND2_X1 U4060 ( .A1(n3521), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3206) );
  NAND2_X1 U4061 ( .A1(n3553), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3205) );
  NAND2_X1 U4062 ( .A1(n3537), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3204)
         );
  NAND2_X1 U4063 ( .A1(n4508), .A2(n3482), .ZN(n3227) );
  AOI22_X1 U4064 ( .A1(n3547), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3519), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3215) );
  AOI22_X1 U4065 ( .A1(n3518), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3407), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3214) );
  AOI22_X1 U4066 ( .A1(n3513), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3520), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3213) );
  AOI22_X1 U4067 ( .A1(n3512), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3408), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3212) );
  AOI22_X1 U4068 ( .A1(n3544), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3414), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3219) );
  AOI22_X1 U4069 ( .A1(n3415), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3536), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3218) );
  AOI22_X1 U4070 ( .A1(n3521), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3553), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3217) );
  NAND2_X4 U4071 ( .A1(n3221), .A2(n3220), .ZN(n4249) );
  NAND2_X1 U4072 ( .A1(n4249), .A2(n3482), .ZN(n3224) );
  AND2_X1 U4073 ( .A1(n4313), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n3222)
         );
  AOI21_X1 U4074 ( .B1(n4275), .B2(EBX_REG_30__SCAN_IN), .A(n3222), .ZN(n4181)
         );
  MUX2_X1 U4075 ( .A(n3301), .B(n5665), .S(EBX_REG_3__SCAN_IN), .Z(n3223) );
  OAI21_X1 U4076 ( .B1(INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n4275), .A(n3223), 
        .ZN(n4556) );
  INV_X1 U4077 ( .A(n4556), .ZN(n3235) );
  NAND2_X1 U4078 ( .A1(n3224), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n3225)
         );
  NAND2_X1 U4079 ( .A1(n3227), .A2(EBX_REG_0__SCAN_IN), .ZN(n3229) );
  INV_X1 U4080 ( .A(EBX_REG_0__SCAN_IN), .ZN(n5125) );
  NAND2_X1 U4081 ( .A1(n3462), .A2(n5125), .ZN(n3228) );
  NAND2_X1 U4082 ( .A1(n3229), .A2(n3228), .ZN(n4274) );
  XNOR2_X1 U4083 ( .A(n3230), .B(n4274), .ZN(n5194) );
  INV_X1 U4084 ( .A(n3230), .ZN(n3231) );
  NAND2_X1 U4085 ( .A1(n3231), .A2(n4274), .ZN(n3232) );
  NAND2_X1 U4086 ( .A1(n4311), .A2(n3232), .ZN(n4402) );
  MUX2_X1 U4087 ( .A(n5665), .B(n3157), .S(EBX_REG_2__SCAN_IN), .Z(n3234) );
  NAND2_X1 U4088 ( .A1(n3224), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3233)
         );
  NOR2_X2 U4089 ( .A1(n4402), .A2(n4401), .ZN(n4553) );
  NAND2_X1 U4090 ( .A1(n3235), .A2(n4553), .ZN(n4554) );
  INV_X1 U4091 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6412) );
  NAND2_X1 U4092 ( .A1(n3157), .A2(n6412), .ZN(n3238) );
  INV_X1 U4093 ( .A(EBX_REG_4__SCAN_IN), .ZN(n3239) );
  NAND2_X1 U4094 ( .A1(n4306), .A2(n3239), .ZN(n3237) );
  NAND3_X1 U4095 ( .A1(n3238), .A2(n5665), .A3(n3237), .ZN(n3241) );
  NAND2_X1 U4096 ( .A1(n5344), .A2(n3239), .ZN(n3240) );
  MUX2_X1 U4097 ( .A(n3301), .B(n5665), .S(EBX_REG_5__SCAN_IN), .Z(n3244) );
  OAI21_X1 U4098 ( .B1(INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n4275), .A(n3244), 
        .ZN(n4536) );
  NOR2_X2 U4099 ( .A1(n4537), .A2(n4536), .ZN(n4549) );
  INV_X1 U4100 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n6396) );
  NAND2_X1 U4101 ( .A1(n3157), .A2(n6396), .ZN(n3246) );
  INV_X1 U4102 ( .A(EBX_REG_6__SCAN_IN), .ZN(n4550) );
  NAND2_X1 U4103 ( .A1(n4306), .A2(n4550), .ZN(n3245) );
  NAND3_X1 U4104 ( .A1(n3246), .A2(n5665), .A3(n3245), .ZN(n3248) );
  NAND2_X1 U4105 ( .A1(n5344), .A2(n4550), .ZN(n3247) );
  NAND2_X1 U4106 ( .A1(n3248), .A2(n3247), .ZN(n4548) );
  MUX2_X1 U4107 ( .A(n3301), .B(n5665), .S(EBX_REG_7__SCAN_IN), .Z(n3249) );
  OAI21_X1 U4108 ( .B1(INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n4275), .A(n3249), 
        .ZN(n4767) );
  INV_X1 U4109 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n6381) );
  NAND2_X1 U4110 ( .A1(n3157), .A2(n6381), .ZN(n3253) );
  INV_X1 U4111 ( .A(EBX_REG_8__SCAN_IN), .ZN(n5105) );
  NAND2_X1 U4112 ( .A1(n4306), .A2(n5105), .ZN(n3252) );
  NAND3_X1 U4113 ( .A1(n3253), .A2(n5665), .A3(n3252), .ZN(n3255) );
  NAND2_X1 U4114 ( .A1(n5344), .A2(n5105), .ZN(n3254) );
  AND2_X1 U4115 ( .A1(n3255), .A2(n3254), .ZN(n4703) );
  MUX2_X1 U4116 ( .A(n3301), .B(n5665), .S(EBX_REG_9__SCAN_IN), .Z(n3256) );
  OAI21_X1 U4117 ( .B1(INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n4275), .A(n3256), 
        .ZN(n5070) );
  MUX2_X1 U4118 ( .A(n5665), .B(n3157), .S(EBX_REG_10__SCAN_IN), .Z(n3258) );
  INV_X1 U4119 ( .A(n4306), .ZN(n4313) );
  NAND2_X1 U4120 ( .A1(n4313), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n3257) );
  NAND2_X1 U4121 ( .A1(n3258), .A2(n3257), .ZN(n5092) );
  INV_X1 U4122 ( .A(n3301), .ZN(n3290) );
  INV_X1 U4123 ( .A(EBX_REG_11__SCAN_IN), .ZN(n5183) );
  NAND2_X1 U4124 ( .A1(n3290), .A2(n5183), .ZN(n3261) );
  NAND2_X1 U4125 ( .A1(n5665), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n3259) );
  OAI211_X1 U4126 ( .C1(n4313), .C2(EBX_REG_11__SCAN_IN), .A(n3157), .B(n3259), 
        .ZN(n3260) );
  MUX2_X1 U4127 ( .A(n5665), .B(n3157), .S(EBX_REG_12__SCAN_IN), .Z(n3263) );
  NAND2_X1 U4128 ( .A1(n4313), .A2(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n3262) );
  AND2_X1 U4129 ( .A1(n3263), .A2(n3262), .ZN(n5149) );
  OR2_X2 U4130 ( .A1(n5148), .A2(n5149), .ZN(n5274) );
  NAND2_X1 U4131 ( .A1(n5665), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n3264) );
  OAI211_X1 U4132 ( .C1(n4313), .C2(EBX_REG_13__SCAN_IN), .A(n3157), .B(n3264), 
        .ZN(n3265) );
  OAI21_X1 U4133 ( .B1(n3301), .B2(EBX_REG_13__SCAN_IN), .A(n3265), .ZN(n5275)
         );
  MUX2_X1 U4134 ( .A(n5665), .B(n3157), .S(EBX_REG_14__SCAN_IN), .Z(n3267) );
  NAND2_X1 U4135 ( .A1(n4313), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n3266) );
  NAND2_X1 U4136 ( .A1(n3267), .A2(n3266), .ZN(n5625) );
  INV_X1 U4137 ( .A(EBX_REG_15__SCAN_IN), .ZN(n5687) );
  NAND2_X1 U4138 ( .A1(n3290), .A2(n5687), .ZN(n3270) );
  NAND2_X1 U4139 ( .A1(n5665), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n3268) );
  OAI211_X1 U4140 ( .C1(n4313), .C2(EBX_REG_15__SCAN_IN), .A(n3157), .B(n3268), 
        .ZN(n3269) );
  AND2_X1 U4141 ( .A1(n3270), .A2(n3269), .ZN(n5610) );
  MUX2_X1 U4142 ( .A(n5665), .B(n3157), .S(EBX_REG_16__SCAN_IN), .Z(n3272) );
  NAND2_X1 U4143 ( .A1(n4313), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n3271) );
  NAND2_X1 U4144 ( .A1(n3272), .A2(n3271), .ZN(n5370) );
  INV_X1 U4145 ( .A(n5370), .ZN(n5677) );
  NAND2_X1 U4146 ( .A1(n5665), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n3273) );
  OAI211_X1 U4147 ( .C1(n4313), .C2(EBX_REG_17__SCAN_IN), .A(n3157), .B(n3273), 
        .ZN(n3274) );
  OAI21_X1 U4148 ( .B1(n3301), .B2(EBX_REG_17__SCAN_IN), .A(n3274), .ZN(n5676)
         );
  INV_X1 U4149 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5961) );
  NAND2_X1 U4150 ( .A1(n3157), .A2(n5961), .ZN(n3277) );
  INV_X1 U4151 ( .A(EBX_REG_19__SCAN_IN), .ZN(n5581) );
  NAND2_X1 U4152 ( .A1(n4306), .A2(n5581), .ZN(n3276) );
  NAND3_X1 U4153 ( .A1(n3277), .A2(n5665), .A3(n3276), .ZN(n3279) );
  NAND2_X1 U4154 ( .A1(n5344), .A2(n5581), .ZN(n3278) );
  AND2_X1 U4155 ( .A1(n3279), .A2(n3278), .ZN(n5346) );
  NOR2_X2 U4156 ( .A1(n5679), .A2(n5346), .ZN(n5663) );
  INV_X1 U4157 ( .A(n4275), .ZN(n4263) );
  INV_X1 U4158 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5955) );
  NOR2_X1 U4159 ( .A1(n4313), .A2(EBX_REG_20__SCAN_IN), .ZN(n3280) );
  AOI21_X1 U4160 ( .B1(n4263), .B2(n5955), .A(n3280), .ZN(n5666) );
  OR2_X1 U4161 ( .A1(n4275), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n3281)
         );
  INV_X1 U4162 ( .A(EBX_REG_18__SCAN_IN), .ZN(n5592) );
  NAND2_X1 U4163 ( .A1(n4306), .A2(n5592), .ZN(n5345) );
  NAND2_X1 U4164 ( .A1(n3281), .A2(n5345), .ZN(n5664) );
  NAND2_X1 U4165 ( .A1(n5344), .A2(EBX_REG_20__SCAN_IN), .ZN(n3283) );
  NAND2_X1 U4166 ( .A1(n5664), .A2(n5665), .ZN(n3282) );
  OAI211_X1 U4167 ( .C1(n5666), .C2(n5664), .A(n3283), .B(n3282), .ZN(n3284)
         );
  INV_X1 U4168 ( .A(n3284), .ZN(n3285) );
  NAND2_X1 U4169 ( .A1(n5663), .A2(n3285), .ZN(n5655) );
  MUX2_X1 U4170 ( .A(n3301), .B(n5665), .S(EBX_REG_21__SCAN_IN), .Z(n3286) );
  OAI21_X1 U4171 ( .B1(INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n4275), .A(n3286), 
        .ZN(n5654) );
  INV_X1 U4172 ( .A(n3287), .ZN(n5657) );
  MUX2_X1 U4173 ( .A(n5665), .B(n3157), .S(EBX_REG_22__SCAN_IN), .Z(n3289) );
  NAND2_X1 U4174 ( .A1(n4313), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n3288) );
  AND2_X1 U4175 ( .A1(n3289), .A2(n3288), .ZN(n5571) );
  INV_X1 U4176 ( .A(EBX_REG_23__SCAN_IN), .ZN(n6022) );
  NAND2_X1 U4177 ( .A1(n3290), .A2(n6022), .ZN(n3293) );
  NAND2_X1 U4178 ( .A1(n5665), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n3291) );
  OAI211_X1 U4179 ( .C1(n4313), .C2(EBX_REG_23__SCAN_IN), .A(n3157), .B(n3291), 
        .ZN(n3292) );
  AND2_X1 U4180 ( .A1(n3293), .A2(n3292), .ZN(n5924) );
  AND2_X2 U4181 ( .A1(n5923), .A2(n5924), .ZN(n5921) );
  MUX2_X1 U4182 ( .A(n5665), .B(n3157), .S(EBX_REG_24__SCAN_IN), .Z(n3295) );
  NAND2_X1 U4183 ( .A1(n4313), .A2(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n3294) );
  NAND2_X1 U4184 ( .A1(n3295), .A2(n3294), .ZN(n5561) );
  MUX2_X1 U4185 ( .A(n3301), .B(n5665), .S(EBX_REG_25__SCAN_IN), .Z(n3296) );
  OAI21_X1 U4186 ( .B1(INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n4275), .A(n3296), 
        .ZN(n5550) );
  OR2_X2 U4187 ( .A1(n5549), .A2(n5550), .ZN(n5552) );
  INV_X1 U4188 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5743) );
  NAND2_X1 U4189 ( .A1(n3157), .A2(n5743), .ZN(n3298) );
  INV_X1 U4190 ( .A(EBX_REG_26__SCAN_IN), .ZN(n5536) );
  NAND2_X1 U4191 ( .A1(n4306), .A2(n5536), .ZN(n3297) );
  NAND3_X1 U4192 ( .A1(n3298), .A2(n5665), .A3(n3297), .ZN(n3300) );
  NAND2_X1 U4193 ( .A1(n5344), .A2(n5536), .ZN(n3299) );
  AND2_X1 U4194 ( .A1(n3300), .A2(n3299), .ZN(n5533) );
  OR2_X2 U4195 ( .A1(n5552), .A2(n5533), .ZN(n5535) );
  MUX2_X1 U4196 ( .A(n3301), .B(n5665), .S(EBX_REG_27__SCAN_IN), .Z(n3302) );
  OAI21_X1 U4197 ( .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n4275), .A(n3302), 
        .ZN(n5518) );
  NOR2_X4 U4198 ( .A1(n5535), .A2(n5518), .ZN(n5517) );
  INV_X1 U4199 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5879) );
  NAND2_X1 U4200 ( .A1(n3157), .A2(n5879), .ZN(n3303) );
  OAI211_X1 U4201 ( .C1(EBX_REG_28__SCAN_IN), .C2(n4313), .A(n3303), .B(n5665), 
        .ZN(n3305) );
  OR2_X1 U4202 ( .A1(n5665), .A2(EBX_REG_28__SCAN_IN), .ZN(n3304) );
  NAND2_X1 U4203 ( .A1(n3305), .A2(n3304), .ZN(n5504) );
  INV_X1 U4204 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5873) );
  NOR2_X1 U4205 ( .A1(n4313), .A2(EBX_REG_29__SCAN_IN), .ZN(n3306) );
  AOI21_X1 U4206 ( .B1(n4263), .B2(n5873), .A(n3306), .ZN(n5488) );
  INV_X1 U4207 ( .A(n4180), .ZN(n4179) );
  OR2_X1 U4208 ( .A1(n5665), .A2(EBX_REG_29__SCAN_IN), .ZN(n5489) );
  INV_X1 U4209 ( .A(n5506), .ZN(n4182) );
  NOR2_X1 U4210 ( .A1(n4180), .A2(n5344), .ZN(n4177) );
  AOI21_X1 U4211 ( .B1(n4181), .B2(n5493), .A(n4177), .ZN(n3308) );
  OAI22_X1 U4212 ( .A1(n4275), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        EBX_REG_31__SCAN_IN), .B2(n4313), .ZN(n3307) );
  XNOR2_X1 U4213 ( .A(n3308), .B(n3307), .ZN(n5865) );
  AOI22_X1 U4214 ( .A1(n3547), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3519), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3312) );
  AOI22_X1 U4215 ( .A1(n3518), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3407), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3311) );
  AOI22_X1 U4216 ( .A1(n3513), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3520), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3310) );
  AOI22_X1 U4217 ( .A1(n3512), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3408), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3309) );
  AOI22_X1 U4218 ( .A1(n3544), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3165), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3316) );
  AOI22_X1 U4219 ( .A1(n3415), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3536), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3315) );
  AOI22_X1 U4220 ( .A1(n3521), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3553), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3314) );
  AOI22_X1 U4221 ( .A1(n3413), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3537), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3313) );
  INV_X2 U4222 ( .A(n4582), .ZN(n3464) );
  NAND2_X1 U4223 ( .A1(n4681), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3321) );
  NAND2_X1 U4224 ( .A1(n4360), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3320) );
  NAND2_X1 U4225 ( .A1(n3321), .A2(n3320), .ZN(n3344) );
  NAND2_X1 U4226 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n6610), .ZN(n3345) );
  NAND2_X1 U4227 ( .A1(n3322), .A2(n3321), .ZN(n3363) );
  NAND2_X1 U4228 ( .A1(n6620), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3324) );
  NAND2_X1 U4229 ( .A1(n5467), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3323) );
  NAND2_X1 U4230 ( .A1(n3363), .A2(n3361), .ZN(n3325) );
  NAND2_X1 U4231 ( .A1(n3325), .A2(n3324), .ZN(n3329) );
  MUX2_X1 U4232 ( .A(n4929), .B(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .S(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n3328) );
  INV_X1 U4233 ( .A(n3328), .ZN(n3326) );
  XNOR2_X1 U4234 ( .A(n3329), .B(n3326), .ZN(n3331) );
  NOR2_X1 U4235 ( .A1(n4447), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3327)
         );
  AOI21_X1 U4236 ( .B1(n3329), .B2(n3328), .A(n3327), .ZN(n3377) );
  AND2_X1 U4237 ( .A1(n3377), .A2(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n3376)
         );
  INV_X1 U4238 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4388) );
  NAND2_X1 U4239 ( .A1(n3376), .A2(n4388), .ZN(n3330) );
  OR2_X1 U4240 ( .A1(n3733), .A2(n3451), .ZN(n3342) );
  AOI22_X1 U4241 ( .A1(n3407), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        INSTQUEUE_REG_13__5__SCAN_IN), .B2(n3518), .ZN(n3336) );
  AOI22_X1 U4242 ( .A1(n3547), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3519), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3335) );
  AOI22_X1 U4243 ( .A1(n3513), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3520), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3334) );
  AOI22_X1 U4244 ( .A1(n3512), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3408), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3333) );
  AOI22_X1 U4245 ( .A1(n3521), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3553), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3340) );
  AOI22_X1 U4246 ( .A1(n3413), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3537), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3339) );
  NAND2_X1 U4247 ( .A1(n3342), .A2(n3421), .ZN(n3356) );
  INV_X1 U4248 ( .A(n3345), .ZN(n3343) );
  XNOR2_X1 U4249 ( .A(n3344), .B(n3343), .ZN(n3433) );
  OAI21_X1 U4250 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6610), .A(n3345), 
        .ZN(n3346) );
  NOR2_X1 U4251 ( .A1(n3733), .A2(n3346), .ZN(n3352) );
  INV_X1 U4252 ( .A(n3346), .ZN(n3347) );
  NAND2_X1 U4253 ( .A1(n3463), .A2(n3347), .ZN(n3349) );
  NAND2_X1 U4254 ( .A1(n3349), .A2(n3348), .ZN(n3351) );
  INV_X1 U4255 ( .A(n3421), .ZN(n3470) );
  NAND2_X1 U4256 ( .A1(n3470), .A2(n3348), .ZN(n3350) );
  NAND2_X1 U4257 ( .A1(n3350), .A2(n3451), .ZN(n3366) );
  NAND2_X1 U4258 ( .A1(n3351), .A2(n3366), .ZN(n3355) );
  OAI211_X1 U4259 ( .C1(n3356), .C2(n3433), .A(n3352), .B(n3355), .ZN(n3354)
         );
  NAND2_X1 U4260 ( .A1(n3421), .A2(n4249), .ZN(n4290) );
  NAND3_X1 U4261 ( .A1(n3356), .A2(STATE2_REG_0__SCAN_IN), .A3(n3433), .ZN(
        n3353) );
  NAND3_X1 U4262 ( .A1(n3354), .A2(n3372), .A3(n3353), .ZN(n3360) );
  INV_X1 U4263 ( .A(n3355), .ZN(n3358) );
  INV_X1 U4264 ( .A(n3356), .ZN(n3357) );
  NAND3_X1 U4265 ( .A1(n3358), .A2(n3357), .A3(n3433), .ZN(n3359) );
  NAND2_X1 U4266 ( .A1(n3360), .A2(n3359), .ZN(n3365) );
  NAND2_X1 U4267 ( .A1(n3365), .A2(n3366), .ZN(n3364) );
  INV_X1 U4268 ( .A(n3733), .ZN(n3648) );
  INV_X1 U4269 ( .A(n3361), .ZN(n3362) );
  XNOR2_X1 U4270 ( .A(n3363), .B(n3362), .ZN(n3432) );
  NAND3_X1 U4271 ( .A1(n3364), .A2(n3648), .A3(n3432), .ZN(n3370) );
  INV_X1 U4272 ( .A(n3365), .ZN(n3368) );
  OAI21_X1 U4273 ( .B1(n3734), .B2(n3432), .A(n3366), .ZN(n3367) );
  NAND2_X1 U4274 ( .A1(n3368), .A2(n3367), .ZN(n3369) );
  NAND2_X1 U4275 ( .A1(n3370), .A2(n3369), .ZN(n3371) );
  OAI21_X1 U4276 ( .B1(n3709), .B2(n3434), .A(n3371), .ZN(n3375) );
  INV_X1 U4277 ( .A(n3434), .ZN(n3373) );
  INV_X1 U4278 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6644) );
  AOI22_X1 U4279 ( .A1(n3380), .A2(n3373), .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n6644), .ZN(n3374) );
  NAND2_X1 U4280 ( .A1(n3375), .A2(n3374), .ZN(n3384) );
  INV_X1 U4281 ( .A(n3376), .ZN(n3379) );
  OAI21_X1 U4282 ( .B1(n3377), .B2(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A(n4388), 
        .ZN(n3378) );
  NAND2_X1 U4283 ( .A1(n3380), .A2(n3436), .ZN(n3383) );
  INV_X1 U4284 ( .A(n3436), .ZN(n3381) );
  AND2_X1 U4285 ( .A1(n3493), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6641) );
  AOI22_X1 U4286 ( .A1(n3518), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3407), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3388) );
  AOI22_X1 U4287 ( .A1(n3547), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3519), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3387) );
  AOI22_X1 U4288 ( .A1(n3513), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3520), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3386) );
  AOI22_X1 U4289 ( .A1(n3512), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3408), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3385) );
  NAND4_X1 U4290 ( .A1(n3388), .A2(n3387), .A3(n3386), .A4(n3385), .ZN(n3394)
         );
  AOI22_X1 U4291 ( .A1(n3544), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3414), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3392) );
  AOI22_X1 U4292 ( .A1(n3415), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3536), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3391) );
  AOI22_X1 U4293 ( .A1(n3521), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3553), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3390) );
  AOI22_X1 U4294 ( .A1(n3413), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3537), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3389) );
  NAND4_X1 U4295 ( .A1(n3392), .A2(n3391), .A3(n3390), .A4(n3389), .ZN(n3393)
         );
  INV_X1 U4297 ( .A(n5696), .ZN(n5692) );
  AOI22_X1 U4298 ( .A1(n3512), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3407), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3398) );
  AOI22_X1 U4299 ( .A1(n3547), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3513), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3397) );
  AOI22_X1 U4300 ( .A1(n3521), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3553), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3396) );
  AOI22_X1 U4301 ( .A1(n3414), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3536), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3395) );
  AND4_X1 U4302 ( .A1(n3398), .A2(n3397), .A3(n3396), .A4(n3395), .ZN(n3404)
         );
  AOI22_X1 U4303 ( .A1(n3544), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3415), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3402) );
  AOI22_X1 U4304 ( .A1(n3518), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3408), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3401) );
  AOI22_X1 U4305 ( .A1(n3413), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3537), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3400) );
  AOI22_X1 U4306 ( .A1(n3519), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3520), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3399) );
  NAND2_X1 U4307 ( .A1(n3404), .A2(n3403), .ZN(n3423) );
  NAND2_X1 U4308 ( .A1(n4582), .A2(n3428), .ZN(n3405) );
  AOI22_X1 U4310 ( .A1(n3518), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3407), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3412) );
  AOI22_X1 U4311 ( .A1(n3547), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3519), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3411) );
  AOI22_X1 U4312 ( .A1(n3513), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3520), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3410) );
  AOI22_X1 U4313 ( .A1(n3512), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3408), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3409) );
  AOI22_X1 U4314 ( .A1(n3413), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3537), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3419) );
  AOI22_X1 U4315 ( .A1(n3521), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3553), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3418) );
  AOI22_X1 U4316 ( .A1(n3544), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3414), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3417) );
  AOI22_X1 U4317 ( .A1(n3415), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3536), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3416) );
  NAND3_X1 U4319 ( .A1(n5696), .A2(n3406), .A3(n3422), .ZN(n4200) );
  NAND2_X1 U4320 ( .A1(n6238), .A2(n5480), .ZN(n4204) );
  INV_X1 U4321 ( .A(n3473), .ZN(n3431) );
  NAND2_X1 U4322 ( .A1(n3424), .A2(n3423), .ZN(n3425) );
  NAND2_X1 U4323 ( .A1(n3425), .A2(n4503), .ZN(n3467) );
  INV_X1 U4324 ( .A(n3163), .ZN(n3430) );
  NAND2_X1 U4325 ( .A1(n3474), .A2(n4294), .ZN(n3504) );
  INV_X1 U4326 ( .A(n3463), .ZN(n4216) );
  AND3_X1 U4327 ( .A1(n3504), .A2(n4216), .A3(n4498), .ZN(n3429) );
  NAND3_X1 U4328 ( .A1(n3431), .A2(n3430), .A3(n3429), .ZN(n3481) );
  AND3_X1 U4329 ( .A1(n3434), .A2(n3433), .A3(n3432), .ZN(n3435) );
  OR2_X1 U4330 ( .A1(n5476), .A2(n5469), .ZN(n5481) );
  INV_X1 U4331 ( .A(n6641), .ZN(n6648) );
  INV_X1 U4332 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6709) );
  NOR2_X1 U4333 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6724) );
  INV_X1 U4334 ( .A(n6724), .ZN(n6652) );
  NOR3_X1 U4335 ( .A1(n6709), .A2(n6644), .A3(n6652), .ZN(n6639) );
  INV_X2 U4336 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6636) );
  NAND2_X1 U4337 ( .A1(n6644), .A2(n6636), .ZN(n3437) );
  INV_X1 U4338 ( .A(n3437), .ZN(n6655) );
  NAND2_X1 U4339 ( .A1(n5463), .A2(n6655), .ZN(n6407) );
  INV_X2 U4340 ( .A(n6407), .ZN(n6422) );
  NOR3_X1 U4341 ( .A1(STATEBS16_REG_SCAN_IN), .A2(n3437), .A3(n6645), .ZN(
        n6651) );
  OR2_X1 U4342 ( .A1(n6422), .A2(n6651), .ZN(n3438) );
  INV_X1 U4343 ( .A(READY_N), .ZN(n6718) );
  NAND2_X1 U4344 ( .A1(n6718), .A2(n6999), .ZN(n4186) );
  NAND3_X1 U4345 ( .A1(n4306), .A2(EBX_REG_31__SCAN_IN), .A3(n4186), .ZN(n3439) );
  INV_X1 U4346 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n3455) );
  NAND2_X1 U4347 ( .A1(STATE_REG_2__SCAN_IN), .A2(STATE_REG_1__SCAN_IN), .ZN(
        n6671) );
  OAI21_X1 U4348 ( .B1(STATE_REG_2__SCAN_IN), .B2(STATE_REG_1__SCAN_IN), .A(
        n6671), .ZN(n3468) );
  OR2_X1 U4349 ( .A1(n3468), .A2(STATE_REG_0__SCAN_IN), .ZN(n6662) );
  NAND2_X1 U4350 ( .A1(n3451), .A2(n6662), .ZN(n4239) );
  INV_X1 U4351 ( .A(n4186), .ZN(n3440) );
  NAND3_X1 U4352 ( .A1(n4239), .A2(n3348), .A3(n3440), .ZN(n3441) );
  INV_X1 U4353 ( .A(REIP_REG_14__SCAN_IN), .ZN(n6687) );
  INV_X1 U4354 ( .A(REIP_REG_11__SCAN_IN), .ZN(n6684) );
  INV_X1 U4355 ( .A(REIP_REG_8__SCAN_IN), .ZN(n6681) );
  INV_X1 U4356 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6676) );
  NAND3_X1 U4357 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_3__SCAN_IN), .A3(
        REIP_REG_2__SCAN_IN), .ZN(n5165) );
  NOR2_X1 U4358 ( .A1(n6676), .A2(n5165), .ZN(n6179) );
  NAND2_X1 U4359 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6179), .ZN(n5264) );
  NAND2_X1 U4360 ( .A1(REIP_REG_7__SCAN_IN), .A2(REIP_REG_6__SCAN_IN), .ZN(
        n5108) );
  NOR3_X1 U4361 ( .A1(n6681), .A2(n5264), .A3(n5108), .ZN(n5236) );
  NAND3_X1 U4362 ( .A1(n5236), .A2(REIP_REG_10__SCAN_IN), .A3(
        REIP_REG_9__SCAN_IN), .ZN(n6121) );
  NOR2_X1 U4363 ( .A1(n6684), .A2(n6121), .ZN(n5181) );
  NAND3_X1 U4364 ( .A1(REIP_REG_13__SCAN_IN), .A2(REIP_REG_12__SCAN_IN), .A3(
        n5181), .ZN(n5631) );
  NOR2_X1 U4365 ( .A1(n6687), .A2(n5631), .ZN(n3457) );
  OR2_X1 U4366 ( .A1(n6181), .A2(n3457), .ZN(n5632) );
  NAND2_X1 U4367 ( .A1(n5632), .A2(n5267), .ZN(n5613) );
  NAND3_X1 U4368 ( .A1(REIP_REG_17__SCAN_IN), .A2(REIP_REG_16__SCAN_IN), .A3(
        REIP_REG_15__SCAN_IN), .ZN(n3458) );
  INV_X1 U4369 ( .A(n3458), .ZN(n3442) );
  NOR2_X1 U4370 ( .A1(n6181), .A2(n3442), .ZN(n3443) );
  NOR2_X1 U4371 ( .A1(n5613), .A2(n3443), .ZN(n6111) );
  INV_X1 U4372 ( .A(REIP_REG_20__SCAN_IN), .ZN(n6691) );
  INV_X1 U4373 ( .A(REIP_REG_19__SCAN_IN), .ZN(n6861) );
  NOR2_X1 U4374 ( .A1(n6691), .A2(n6861), .ZN(n3459) );
  NAND2_X1 U4375 ( .A1(REIP_REG_18__SCAN_IN), .A2(n3459), .ZN(n3444) );
  NAND2_X1 U4376 ( .A1(n5237), .A2(n3444), .ZN(n3445) );
  NAND2_X1 U4377 ( .A1(n6111), .A2(n3445), .ZN(n6011) );
  AND3_X1 U4378 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .ZN(n3446) );
  NOR2_X1 U4379 ( .A1(n6181), .A2(n3446), .ZN(n3447) );
  NOR2_X1 U4380 ( .A1(n6011), .A2(n3447), .ZN(n6003) );
  NAND2_X1 U4381 ( .A1(n6181), .A2(n5267), .ZN(n5628) );
  INV_X1 U4382 ( .A(REIP_REG_24__SCAN_IN), .ZN(n7017) );
  INV_X1 U4383 ( .A(REIP_REG_26__SCAN_IN), .ZN(n7050) );
  INV_X1 U4384 ( .A(REIP_REG_25__SCAN_IN), .ZN(n6825) );
  NOR3_X1 U4385 ( .A1(n7017), .A2(n7050), .A3(n6825), .ZN(n5526) );
  INV_X1 U4386 ( .A(n5526), .ZN(n3448) );
  NAND2_X1 U4387 ( .A1(n5628), .A2(n3448), .ZN(n3449) );
  AND2_X1 U4388 ( .A1(n6003), .A2(n3449), .ZN(n5532) );
  INV_X1 U4389 ( .A(REIP_REG_28__SCAN_IN), .ZN(n7020) );
  INV_X1 U4390 ( .A(REIP_REG_27__SCAN_IN), .ZN(n7030) );
  OAI21_X1 U4391 ( .B1(n7020), .B2(n7030), .A(n5237), .ZN(n3450) );
  AND2_X1 U4392 ( .A1(n5532), .A2(n3450), .ZN(n5509) );
  OAI211_X1 U4393 ( .C1(REIP_REG_29__SCAN_IN), .C2(n6181), .A(n5509), .B(
        REIP_REG_30__SCAN_IN), .ZN(n4195) );
  NAND3_X1 U4394 ( .A1(n4195), .A2(REIP_REG_31__SCAN_IN), .A3(n5628), .ZN(
        n3454) );
  INV_X1 U4395 ( .A(n5127), .ZN(n3452) );
  OR3_X1 U4396 ( .A1(READY_N), .A2(STATEBS16_REG_SCAN_IN), .A3(n6662), .ZN(
        n6632) );
  AND2_X1 U4397 ( .A1(n6240), .A2(n6632), .ZN(n4188) );
  NAND3_X1 U4398 ( .A1(n3452), .A2(EBX_REG_31__SCAN_IN), .A3(n4188), .ZN(n3453) );
  OAI211_X1 U4399 ( .C1(n3455), .C2(n6176), .A(n3454), .B(n3453), .ZN(n3456)
         );
  AOI21_X1 U4400 ( .B1(n5865), .B2(n6153), .A(n3456), .ZN(n4176) );
  INV_X1 U4401 ( .A(REIP_REG_23__SCAN_IN), .ZN(n6694) );
  INV_X1 U4402 ( .A(REIP_REG_22__SCAN_IN), .ZN(n7106) );
  INV_X1 U4403 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6693) );
  NAND2_X1 U4404 ( .A1(n5237), .A2(n3457), .ZN(n6113) );
  NOR2_X1 U4405 ( .A1(n6113), .A2(n3458), .ZN(n5582) );
  NAND2_X1 U4406 ( .A1(n6012), .A2(n3459), .ZN(n5576) );
  NOR4_X1 U4407 ( .A1(n6694), .A2(n7106), .A3(n6693), .A4(n5576), .ZN(n5548)
         );
  AND2_X1 U4408 ( .A1(n5526), .A2(REIP_REG_27__SCAN_IN), .ZN(n3460) );
  NAND2_X1 U4409 ( .A1(n5548), .A2(n3460), .ZN(n5513) );
  NOR2_X1 U4410 ( .A1(n5513), .A2(n7020), .ZN(n5499) );
  INV_X1 U4411 ( .A(REIP_REG_31__SCAN_IN), .ZN(n7082) );
  NAND4_X1 U4412 ( .A1(n5499), .A2(REIP_REG_30__SCAN_IN), .A3(
        REIP_REG_29__SCAN_IN), .A4(n7082), .ZN(n4175) );
  INV_X2 U4413 ( .A(n4020), .ZN(n4131) );
  NAND2_X1 U4414 ( .A1(n6636), .A2(STATEBS16_REG_SCAN_IN), .ZN(n3820) );
  AOI22_X1 U4415 ( .A1(n4131), .A2(EAX_REG_31__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n4039), .ZN(n4170) );
  NAND2_X1 U4416 ( .A1(n3461), .A2(n5696), .ZN(n4244) );
  NAND2_X1 U4418 ( .A1(n3466), .A2(n3465), .ZN(n3502) );
  NOR2_X2 U4419 ( .A1(n3502), .A2(n3467), .ZN(n4264) );
  INV_X1 U4420 ( .A(n3468), .ZN(n3469) );
  NAND3_X1 U4421 ( .A1(n3506), .A2(n4264), .A3(n3471), .ZN(n3477) );
  AND2_X1 U4422 ( .A1(n4498), .A2(n4294), .ZN(n4220) );
  NAND2_X1 U4423 ( .A1(n3476), .A2(n3475), .ZN(n3496) );
  OAI21_X1 U4424 ( .B1(n3477), .B2(n3496), .A(STATE2_REG_0__SCAN_IN), .ZN(
        n3479) );
  NAND2_X1 U4425 ( .A1(n3479), .A2(n3478), .ZN(n3581) );
  NAND2_X1 U4426 ( .A1(n3581), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3488) );
  NAND2_X1 U4427 ( .A1(n3480), .A2(n3173), .ZN(n3485) );
  OR2_X2 U4428 ( .A1(n3481), .A2(n4249), .ZN(n4252) );
  NOR2_X1 U4429 ( .A1(n3498), .A2(n3482), .ZN(n3483) );
  NOR2_X1 U4430 ( .A1(n3421), .A2(n4249), .ZN(n3484) );
  AND2_X1 U4431 ( .A1(n5696), .A2(n4305), .ZN(n4259) );
  NAND2_X1 U4432 ( .A1(n4350), .A2(n4259), .ZN(n4272) );
  NAND3_X1 U4433 ( .A1(n3485), .A2(n4252), .A3(n4272), .ZN(n3486) );
  NAND2_X1 U4434 ( .A1(n3486), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3489) );
  NAND2_X1 U4435 ( .A1(n5463), .A2(n6644), .ZN(n4231) );
  INV_X1 U4436 ( .A(n4231), .ZN(n6720) );
  XNOR2_X1 U4437 ( .A(n6610), .B(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n5019)
         );
  INV_X1 U4438 ( .A(n3493), .ZN(n3634) );
  AND2_X1 U4439 ( .A1(n3634), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3487)
         );
  AOI21_X1 U4440 ( .B1(n6720), .B2(n5019), .A(n3487), .ZN(n3490) );
  NAND3_X1 U4441 ( .A1(n3488), .A2(n3489), .A3(n3490), .ZN(n3577) );
  INV_X1 U4442 ( .A(n3489), .ZN(n3492) );
  INV_X1 U4443 ( .A(n3490), .ZN(n3491) );
  NAND2_X1 U4444 ( .A1(n3492), .A2(n3171), .ZN(n3579) );
  NAND2_X1 U4445 ( .A1(n3577), .A2(n3579), .ZN(n3511) );
  NAND2_X1 U4446 ( .A1(n3581), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3495) );
  MUX2_X1 U4447 ( .A(n3493), .B(n4231), .S(n6610), .Z(n3494) );
  NAND2_X1 U4448 ( .A1(n3495), .A2(n3494), .ZN(n3576) );
  NAND2_X1 U4449 ( .A1(n4216), .A2(n4249), .ZN(n3497) );
  NAND2_X1 U4450 ( .A1(n3496), .A2(n3497), .ZN(n3500) );
  NAND2_X1 U4451 ( .A1(n3498), .A2(n3348), .ZN(n3499) );
  INV_X1 U4452 ( .A(n4324), .ZN(n3501) );
  NOR2_X1 U4453 ( .A1(n3406), .A2(n3501), .ZN(n3503) );
  OAI21_X1 U4454 ( .B1(n3503), .B2(n3502), .A(n4249), .ZN(n3508) );
  INV_X1 U4455 ( .A(n3838), .ZN(n4267) );
  NAND2_X1 U4456 ( .A1(n5463), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6647) );
  AOI21_X1 U4457 ( .B1(n4268), .B2(n4267), .A(n6647), .ZN(n3507) );
  NAND2_X1 U4458 ( .A1(n3504), .A2(n6240), .ZN(n3505) );
  NAND3_X1 U4459 ( .A1(n3508), .A2(n3507), .A3(n3168), .ZN(n3509) );
  INV_X1 U4460 ( .A(n3529), .ZN(n3578) );
  NAND2_X1 U4461 ( .A1(n3576), .A2(n3578), .ZN(n3510) );
  AOI22_X1 U4462 ( .A1(n4139), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4148), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3517) );
  AOI22_X1 U4463 ( .A1(n3772), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n4149), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3516) );
  INV_X1 U4464 ( .A(n3513), .ZN(n3535) );
  INV_X1 U4465 ( .A(n3407), .ZN(n3652) );
  INV_X1 U4466 ( .A(n3652), .ZN(n4103) );
  AOI22_X1 U4467 ( .A1(n3546), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3515) );
  AOI22_X1 U4468 ( .A1(n3414), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3554), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3514) );
  NAND4_X1 U4469 ( .A1(n3517), .A2(n3516), .A3(n3515), .A4(n3514), .ZN(n3527)
         );
  AOI22_X1 U4470 ( .A1(n4150), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4143), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3525) );
  INV_X1 U4471 ( .A(n3520), .ZN(n4372) );
  INV_X2 U4472 ( .A(n4372), .ZN(n4141) );
  AOI22_X1 U4473 ( .A1(n4140), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n4141), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3524) );
  AOI22_X1 U4474 ( .A1(n4151), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n4098), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3523) );
  AOI22_X1 U4475 ( .A1(n4142), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3158), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3522) );
  NAND4_X1 U4476 ( .A1(n3525), .A2(n3524), .A3(n3523), .A4(n3522), .ZN(n3526)
         );
  NAND2_X1 U4477 ( .A1(n4797), .A2(n4291), .ZN(n3528) );
  OAI21_X2 U4478 ( .B1(n4348), .B2(STATE2_REG_0__SCAN_IN), .A(n3528), .ZN(
        n3573) );
  XNOR2_X1 U4479 ( .A(n3576), .B(n3529), .ZN(n3611) );
  NAND2_X1 U4480 ( .A1(n3709), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3564) );
  AOI22_X1 U4481 ( .A1(n3544), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4148), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3534) );
  INV_X1 U4482 ( .A(n3652), .ZN(n3552) );
  AOI22_X1 U4483 ( .A1(n4143), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3552), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3533) );
  AOI22_X1 U4484 ( .A1(n3519), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n4141), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3532) );
  CLKBUF_X1 U4485 ( .A(n3553), .Z(n3530) );
  AOI22_X1 U4486 ( .A1(n3521), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3530), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3531) );
  NAND4_X1 U4487 ( .A1(n3534), .A2(n3533), .A3(n3532), .A4(n3531), .ZN(n3543)
         );
  AOI22_X1 U4488 ( .A1(n4150), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3546), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3541) );
  AOI22_X1 U4489 ( .A1(n3414), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3536), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3540) );
  AOI22_X1 U4490 ( .A1(n3772), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3408), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3539) );
  AOI22_X1 U4491 ( .A1(n4098), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3158), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3538) );
  NAND4_X1 U4492 ( .A1(n3541), .A2(n3540), .A3(n3539), .A4(n3538), .ZN(n3542)
         );
  AOI22_X1 U4493 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n3544), .B1(n3414), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3551) );
  AOI22_X1 U4494 ( .A1(n3546), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3519), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3550) );
  AOI22_X1 U4495 ( .A1(n4150), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3772), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3549) );
  AOI22_X1 U4496 ( .A1(n3521), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3158), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3548) );
  NAND4_X1 U4497 ( .A1(n3551), .A2(n3550), .A3(n3549), .A4(n3548), .ZN(n3560)
         );
  AOI22_X1 U4498 ( .A1(INSTQUEUE_REG_10__0__SCAN_IN), .A2(n4148), .B1(n3536), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3558) );
  AOI22_X1 U4499 ( .A1(INSTQUEUE_REG_12__0__SCAN_IN), .A2(n3552), .B1(n4141), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3557) );
  AOI22_X1 U4500 ( .A1(n3518), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3408), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3556) );
  AOI22_X1 U4501 ( .A1(n4098), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3554), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3555) );
  NAND4_X1 U4502 ( .A1(n3558), .A2(n3557), .A3(n3556), .A4(n3555), .ZN(n3559)
         );
  NAND2_X1 U4503 ( .A1(n4498), .A2(n4292), .ZN(n3561) );
  OAI211_X1 U4504 ( .C1(n3732), .C2(n3464), .A(STATE2_REG_0__SCAN_IN), .B(
        n3561), .ZN(n3562) );
  INV_X1 U4505 ( .A(n3562), .ZN(n3563) );
  NAND2_X1 U4506 ( .A1(n3564), .A2(n3563), .ZN(n3607) );
  XNOR2_X1 U4507 ( .A(n3732), .B(n4292), .ZN(n3565) );
  AOI21_X2 U4508 ( .B1(n3611), .B2(n6644), .A(n3566), .ZN(n3605) );
  NAND2_X1 U4509 ( .A1(n4797), .A2(n4800), .ZN(n3567) );
  AND2_X2 U4510 ( .A1(n3605), .A2(n3567), .ZN(n3571) );
  INV_X1 U4511 ( .A(n4797), .ZN(n3570) );
  NAND2_X1 U4512 ( .A1(n3709), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3569) );
  NOR2_X1 U4513 ( .A1(n3348), .A2(n6644), .ZN(n3600) );
  NAND2_X1 U4514 ( .A1(n3600), .A2(n4291), .ZN(n3568) );
  OAI211_X1 U4515 ( .C1(n4800), .C2(n3570), .A(n3569), .B(n3568), .ZN(n3617)
         );
  NAND2_X1 U4516 ( .A1(n3619), .A2(n3617), .ZN(n3575) );
  INV_X1 U4517 ( .A(n3571), .ZN(n3572) );
  NAND2_X1 U4518 ( .A1(n3573), .A2(n3572), .ZN(n3574) );
  NAND3_X1 U4519 ( .A1(n3578), .A2(n3577), .A3(n3576), .ZN(n3580) );
  NAND2_X1 U4520 ( .A1(n3162), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3586) );
  AND2_X1 U4521 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n3582) );
  NAND2_X1 U4522 ( .A1(n3582), .A2(n6620), .ZN(n6436) );
  INV_X1 U4523 ( .A(n3582), .ZN(n3583) );
  NAND2_X1 U4524 ( .A1(n3583), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3584) );
  NAND2_X1 U4525 ( .A1(n6436), .A2(n3584), .ZN(n4648) );
  AOI22_X1 U4526 ( .A1(n6720), .A2(n4648), .B1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n3634), .ZN(n3585) );
  NAND2_X1 U4527 ( .A1(n4450), .A2(n6644), .ZN(n3599) );
  AOI22_X1 U4528 ( .A1(n4143), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3591) );
  AOI22_X1 U4529 ( .A1(n4150), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4140), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3590) );
  AOI22_X1 U4530 ( .A1(n3546), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4141), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3589) );
  AOI22_X1 U4531 ( .A1(n3772), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4142), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3588) );
  NAND4_X1 U4532 ( .A1(n3591), .A2(n3590), .A3(n3589), .A4(n3588), .ZN(n3597)
         );
  AOI22_X1 U4533 ( .A1(n4139), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3545), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3595) );
  AOI22_X1 U4534 ( .A1(n4148), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4149), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3594) );
  AOI22_X1 U4535 ( .A1(n4151), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3530), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3593) );
  AOI22_X1 U4536 ( .A1(n4098), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3158), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3592) );
  NAND4_X1 U4537 ( .A1(n3595), .A2(n3594), .A3(n3593), .A4(n3592), .ZN(n3596)
         );
  INV_X1 U4538 ( .A(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4828) );
  INV_X1 U4539 ( .A(n4415), .ZN(n4425) );
  INV_X1 U4540 ( .A(n3600), .ZN(n3601) );
  OAI22_X1 U4541 ( .A1(n3734), .A2(n4828), .B1(n4425), .B2(n3601), .ZN(n3602)
         );
  NOR2_X2 U4542 ( .A1(n4305), .A2(n6636), .ZN(n3961) );
  NAND2_X1 U4543 ( .A1(n4483), .A2(n3961), .ZN(n3604) );
  NAND2_X1 U4544 ( .A1(n3604), .A2(n3820), .ZN(n3627) );
  INV_X1 U4545 ( .A(n3605), .ZN(n3609) );
  NOR2_X1 U4546 ( .A1(n3607), .A2(n3606), .ZN(n3608) );
  BUF_X2 U4547 ( .A(n4217), .Z(n4920) );
  NAND2_X1 U4548 ( .A1(n4920), .A2(n4267), .ZN(n3610) );
  NAND2_X1 U4549 ( .A1(n3610), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4225) );
  AND2_X1 U4551 ( .A1(n4259), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3620) );
  INV_X1 U4552 ( .A(n3620), .ZN(n3681) );
  NAND2_X1 U4553 ( .A1(PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n6636), .ZN(n3613)
         );
  NAND2_X1 U4554 ( .A1(n4131), .A2(EAX_REG_0__SCAN_IN), .ZN(n3612) );
  OAI211_X1 U4555 ( .C1(n3681), .C2(n5359), .A(n3613), .B(n3612), .ZN(n3614)
         );
  AOI21_X1 U4556 ( .B1(n5351), .B2(n3961), .A(n3614), .ZN(n4224) );
  INV_X1 U4557 ( .A(n4224), .ZN(n3615) );
  NAND2_X1 U4558 ( .A1(n6636), .A2(n6999), .ZN(n4163) );
  OR2_X1 U4559 ( .A1(n3615), .A2(n4163), .ZN(n3616) );
  NAND2_X1 U4560 ( .A1(n4227), .A2(n3616), .ZN(n4285) );
  NAND2_X1 U4561 ( .A1(n4481), .A2(n3961), .ZN(n3624) );
  AOI22_X1 U4562 ( .A1(n4131), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n6636), .ZN(n3622) );
  NAND2_X1 U4563 ( .A1(n3620), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3621) );
  AND2_X1 U4564 ( .A1(n3622), .A2(n3621), .ZN(n3623) );
  NAND2_X1 U4565 ( .A1(n3624), .A2(n3623), .ZN(n4284) );
  AND2_X2 U4566 ( .A1(n4285), .A2(n4284), .ZN(n4282) );
  OR2_X2 U4567 ( .A1(n3627), .A2(n4282), .ZN(n4399) );
  OAI21_X1 U4568 ( .B1(PHYADDRPOINTER_REG_2__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_1__SCAN_IN), .A(n3667), .ZN(n6359) );
  AOI22_X1 U4569 ( .A1(n4165), .A2(n6359), .B1(n4039), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3626) );
  NAND2_X1 U4570 ( .A1(n4131), .A2(EAX_REG_2__SCAN_IN), .ZN(n3625) );
  OAI211_X1 U4571 ( .C1(n3681), .C2(n5467), .A(n3626), .B(n3625), .ZN(n4398)
         );
  NAND2_X1 U4572 ( .A1(n4399), .A2(n4398), .ZN(n3629) );
  NAND2_X1 U4573 ( .A1(n3627), .A2(n4282), .ZN(n3628) );
  NAND2_X2 U4574 ( .A1(n3629), .A2(n3628), .ZN(n4480) );
  NAND2_X1 U4575 ( .A1(n3162), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3636) );
  NAND3_X1 U4576 ( .A1(n4929), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6486) );
  INV_X1 U4577 ( .A(n6486), .ZN(n3632) );
  NAND2_X1 U4578 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n3632), .ZN(n6483) );
  NAND2_X1 U4579 ( .A1(n4929), .A2(n6483), .ZN(n3633) );
  NOR3_X1 U4580 ( .A1(n4929), .A2(n6620), .A3(n4681), .ZN(n4721) );
  NAND2_X1 U4581 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4721), .ZN(n4911) );
  AOI22_X1 U4582 ( .A1(n6720), .A2(n5020), .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n3634), .ZN(n3635) );
  AOI22_X1 U4583 ( .A1(n4143), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3640) );
  AOI22_X1 U4584 ( .A1(n4150), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4140), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3639) );
  AOI22_X1 U4585 ( .A1(n3546), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4141), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3638) );
  AOI22_X1 U4586 ( .A1(n3772), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4142), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3637) );
  NAND4_X1 U4587 ( .A1(n3640), .A2(n3639), .A3(n3638), .A4(n3637), .ZN(n3647)
         );
  AOI22_X1 U4588 ( .A1(n4139), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3545), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3645) );
  AOI22_X1 U4589 ( .A1(n4148), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4149), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3644) );
  AOI22_X1 U4590 ( .A1(n4151), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3554), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3643) );
  INV_X1 U4591 ( .A(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3641) );
  AOI22_X1 U4592 ( .A1(n4098), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3158), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3642) );
  NAND4_X1 U4593 ( .A1(n3645), .A2(n3644), .A3(n3643), .A4(n3642), .ZN(n3646)
         );
  AOI22_X1 U4594 ( .A1(n3648), .A2(n4434), .B1(n3709), .B2(
        INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3649) );
  INV_X1 U4595 ( .A(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4824) );
  OR2_X1 U4596 ( .A1(n3734), .A2(n4824), .ZN(n3664) );
  AOI22_X1 U4597 ( .A1(n4143), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3656) );
  AOI22_X1 U4598 ( .A1(n4150), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4140), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3655) );
  AOI22_X1 U4599 ( .A1(n3546), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4141), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3654) );
  AOI22_X1 U4600 ( .A1(n3772), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4142), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3653) );
  NAND4_X1 U4601 ( .A1(n3656), .A2(n3655), .A3(n3654), .A4(n3653), .ZN(n3662)
         );
  AOI22_X1 U4602 ( .A1(n4139), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3545), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3660) );
  AOI22_X1 U4603 ( .A1(n4148), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4149), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3659) );
  AOI22_X1 U4604 ( .A1(n4151), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3530), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3658) );
  AOI22_X1 U4605 ( .A1(n4098), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3158), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3657) );
  NAND4_X1 U4606 ( .A1(n3660), .A2(n3659), .A3(n3658), .A4(n3657), .ZN(n3661)
         );
  INV_X1 U4607 ( .A(n4565), .ZN(n4518) );
  OR2_X1 U4608 ( .A1(n3733), .A2(n4518), .ZN(n3663) );
  NAND2_X1 U4609 ( .A1(n3664), .A2(n3663), .ZN(n3706) );
  XNOR2_X1 U4610 ( .A(n3705), .B(n3706), .ZN(n4433) );
  NAND2_X1 U4611 ( .A1(n4433), .A2(n3961), .ZN(n3673) );
  NAND2_X1 U4612 ( .A1(n6636), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3666)
         );
  NAND2_X1 U4613 ( .A1(n4131), .A2(EAX_REG_4__SCAN_IN), .ZN(n3665) );
  OAI211_X1 U4614 ( .C1(n3681), .C2(n4388), .A(n3666), .B(n3665), .ZN(n3671)
         );
  INV_X1 U4615 ( .A(n3677), .ZN(n3669) );
  INV_X1 U4616 ( .A(n3699), .ZN(n3668) );
  OAI21_X1 U4617 ( .B1(PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n3669), .A(n3668), 
        .ZN(n5164) );
  AND2_X1 U4618 ( .A1(n4165), .A2(n5164), .ZN(n3670) );
  AOI21_X1 U4619 ( .B1(n3671), .B2(n4163), .A(n3670), .ZN(n3672) );
  NAND2_X1 U4620 ( .A1(n3673), .A2(n3672), .ZN(n4406) );
  XNOR2_X2 U4621 ( .A(n3676), .B(n4482), .ZN(n4424) );
  NAND2_X1 U4622 ( .A1(n4424), .A2(n3961), .ZN(n3684) );
  OAI21_X1 U4623 ( .B1(PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n3678), .A(n3677), 
        .ZN(n6349) );
  AOI22_X1 U4624 ( .A1(n4165), .A2(n6349), .B1(n4039), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3680) );
  NAND2_X1 U4625 ( .A1(n4131), .A2(EAX_REG_3__SCAN_IN), .ZN(n3679) );
  OAI211_X1 U4626 ( .C1(n3681), .C2(n4447), .A(n3680), .B(n3679), .ZN(n3682)
         );
  INV_X1 U4627 ( .A(n3682), .ZN(n3683) );
  NAND2_X1 U4628 ( .A1(n3684), .A2(n3683), .ZN(n4479) );
  NAND2_X1 U4629 ( .A1(n4480), .A2(n3685), .ZN(n4405) );
  INV_X2 U4630 ( .A(n4405), .ZN(n3727) );
  INV_X1 U4631 ( .A(n3706), .ZN(n3686) );
  OR2_X1 U4632 ( .A1(n3705), .A2(n3686), .ZN(n3698) );
  INV_X1 U4633 ( .A(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4853) );
  AOI22_X1 U4634 ( .A1(n4143), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3690) );
  AOI22_X1 U4635 ( .A1(n4150), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4140), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3689) );
  AOI22_X1 U4636 ( .A1(n3546), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4141), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3688) );
  AOI22_X1 U4637 ( .A1(n3772), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4142), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3687) );
  NAND4_X1 U4638 ( .A1(n3690), .A2(n3689), .A3(n3688), .A4(n3687), .ZN(n3696)
         );
  AOI22_X1 U4639 ( .A1(n4139), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3545), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3694) );
  AOI22_X1 U4640 ( .A1(n4148), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4149), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3693) );
  AOI22_X1 U4641 ( .A1(n4151), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3554), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3692) );
  AOI22_X1 U4642 ( .A1(n4098), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3158), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3691) );
  NAND4_X1 U4643 ( .A1(n3694), .A2(n3693), .A3(n3692), .A4(n3691), .ZN(n3695)
         );
  INV_X1 U4644 ( .A(n4564), .ZN(n3697) );
  OAI22_X1 U4645 ( .A1(n3734), .A2(n4853), .B1(n3733), .B2(n3697), .ZN(n3707)
         );
  NAND2_X1 U4646 ( .A1(n4517), .A2(n3961), .ZN(n3704) );
  INV_X1 U4647 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3701) );
  OAI21_X1 U4648 ( .B1(PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n3699), .A(n3736), 
        .ZN(n6341) );
  NAND2_X1 U4649 ( .A1(n6341), .A2(n4165), .ZN(n3700) );
  OAI21_X1 U4650 ( .B1(n3701), .B2(n3820), .A(n3700), .ZN(n3702) );
  AOI21_X1 U4651 ( .B1(n4131), .B2(EAX_REG_5__SCAN_IN), .A(n3702), .ZN(n3703)
         );
  NAND2_X1 U4652 ( .A1(n3704), .A2(n3703), .ZN(n4545) );
  NAND2_X1 U4653 ( .A1(n3708), .A2(n3169), .ZN(n3728) );
  NAND2_X1 U4654 ( .A1(n3709), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3722) );
  AOI22_X1 U4655 ( .A1(n4143), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3713) );
  AOI22_X1 U4656 ( .A1(n4150), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4140), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3712) );
  AOI22_X1 U4657 ( .A1(n3546), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4141), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3711) );
  AOI22_X1 U4658 ( .A1(n3773), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4142), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3710) );
  NAND4_X1 U4659 ( .A1(n3713), .A2(n3712), .A3(n3711), .A4(n3710), .ZN(n3719)
         );
  AOI22_X1 U4660 ( .A1(n4139), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3545), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3717) );
  AOI22_X1 U4661 ( .A1(n4148), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4149), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3716) );
  AOI22_X1 U4662 ( .A1(n4151), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3530), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3715) );
  AOI22_X1 U4663 ( .A1(n4098), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3158), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3714) );
  NAND4_X1 U4664 ( .A1(n3717), .A2(n3716), .A3(n3715), .A4(n3714), .ZN(n3718)
         );
  INV_X1 U4665 ( .A(n4785), .ZN(n3720) );
  OR2_X1 U4666 ( .A1(n3733), .A2(n3720), .ZN(n3721) );
  NAND2_X1 U4667 ( .A1(n3728), .A2(n3729), .ZN(n4563) );
  NAND2_X1 U4668 ( .A1(n4563), .A2(n3961), .ZN(n3725) );
  XNOR2_X1 U4669 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .B(n3736), .ZN(n4573) );
  AOI22_X1 U4670 ( .A1(n4131), .A2(EAX_REG_6__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n6636), .ZN(n3723) );
  MUX2_X1 U4671 ( .A(n4573), .B(n3723), .S(n4163), .Z(n3724) );
  NAND2_X1 U4672 ( .A1(n3725), .A2(n3724), .ZN(n4544) );
  NAND2_X2 U4673 ( .A1(n3727), .A2(n3726), .ZN(n4706) );
  INV_X1 U4674 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4845) );
  OAI22_X1 U4675 ( .A1(n3734), .A2(n4845), .B1(n3733), .B2(n3732), .ZN(n3735)
         );
  INV_X1 U4676 ( .A(EAX_REG_7__SCAN_IN), .ZN(n3739) );
  NAND2_X1 U4677 ( .A1(n3737), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3741)
         );
  OAI21_X1 U4678 ( .B1(PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n3737), .A(n3741), 
        .ZN(n6334) );
  AOI22_X1 U4679 ( .A1(n4165), .A2(n6334), .B1(n4039), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3738) );
  OAI21_X1 U4680 ( .B1(n4020), .B2(n3739), .A(n3738), .ZN(n3740) );
  NOR2_X2 U4681 ( .A1(n4706), .A2(n4707), .ZN(n4699) );
  XOR2_X1 U4682 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .B(n3755), .Z(n5101) );
  AOI22_X1 U4683 ( .A1(INSTQUEUE_REG_12__0__SCAN_IN), .A2(n4150), .B1(n4103), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3745) );
  AOI22_X1 U4684 ( .A1(INSTQUEUE_REG_4__0__SCAN_IN), .A2(n4140), .B1(n4141), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3744) );
  AOI22_X1 U4685 ( .A1(n4139), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4142), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3743) );
  AOI22_X1 U4686 ( .A1(n3545), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4098), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3742) );
  NAND4_X1 U4687 ( .A1(n3745), .A2(n3744), .A3(n3743), .A4(n3742), .ZN(n3751)
         );
  AOI22_X1 U4688 ( .A1(n3773), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4149), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3749) );
  AOI22_X1 U4689 ( .A1(n3546), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n4143), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3748) );
  AOI22_X1 U4690 ( .A1(INSTQUEUE_REG_3__0__SCAN_IN), .A2(n4151), .B1(n3554), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3747) );
  AOI22_X1 U4691 ( .A1(n4148), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3158), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3746) );
  NAND4_X1 U4692 ( .A1(n3749), .A2(n3748), .A3(n3747), .A4(n3746), .ZN(n3750)
         );
  OR2_X1 U4693 ( .A1(n3751), .A2(n3750), .ZN(n3752) );
  AOI22_X1 U4694 ( .A1(n3961), .A2(n3752), .B1(n4039), .B2(
        PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3754) );
  NAND2_X1 U4695 ( .A1(n4131), .A2(EAX_REG_8__SCAN_IN), .ZN(n3753) );
  OAI211_X1 U4696 ( .C1(n5101), .C2(n4163), .A(n3754), .B(n3753), .ZN(n4698)
         );
  XNOR2_X1 U4697 ( .A(n3771), .B(n5240), .ZN(n5238) );
  AOI22_X1 U4698 ( .A1(n3545), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4151), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3759) );
  AOI22_X1 U4699 ( .A1(n4150), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3546), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3758) );
  AOI22_X1 U4700 ( .A1(n4139), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4148), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3757) );
  AOI22_X1 U4701 ( .A1(n4143), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3756) );
  NAND4_X1 U4702 ( .A1(n3759), .A2(n3758), .A3(n3757), .A4(n3756), .ZN(n3765)
         );
  AOI22_X1 U4703 ( .A1(n4140), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n4141), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3763) );
  AOI22_X1 U4704 ( .A1(n3773), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4142), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3762) );
  AOI22_X1 U4705 ( .A1(n4098), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3530), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3761) );
  AOI22_X1 U4706 ( .A1(n4149), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3158), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3760) );
  NAND4_X1 U4707 ( .A1(n3763), .A2(n3762), .A3(n3761), .A4(n3760), .ZN(n3764)
         );
  OAI21_X1 U4708 ( .B1(n3765), .B2(n3764), .A(n3961), .ZN(n3768) );
  NAND2_X1 U4709 ( .A1(n4131), .A2(EAX_REG_9__SCAN_IN), .ZN(n3767) );
  NAND2_X1 U4710 ( .A1(n4039), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3766)
         );
  NAND3_X1 U4711 ( .A1(n3768), .A2(n3767), .A3(n3766), .ZN(n3769) );
  AOI21_X1 U4712 ( .B1(n5238), .B2(n4165), .A(n3769), .ZN(n5068) );
  NAND2_X1 U4713 ( .A1(n3176), .A2(n3770), .ZN(n5080) );
  XNOR2_X1 U4714 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .B(n3788), .ZN(n6156)
         );
  AOI22_X1 U4715 ( .A1(n4139), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3773), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3777) );
  AOI22_X1 U4716 ( .A1(n4150), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3776) );
  AOI22_X1 U4717 ( .A1(n4140), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4141), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3775) );
  AOI22_X1 U4718 ( .A1(n4098), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3158), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3774) );
  NAND4_X1 U4719 ( .A1(n3777), .A2(n3776), .A3(n3775), .A4(n3774), .ZN(n3783)
         );
  AOI22_X1 U4720 ( .A1(n3545), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4148), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3781) );
  AOI22_X1 U4721 ( .A1(n3546), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4143), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3780) );
  AOI22_X1 U4722 ( .A1(n4149), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4142), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3779) );
  AOI22_X1 U4723 ( .A1(n4151), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n3554), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3778) );
  NAND4_X1 U4724 ( .A1(n3781), .A2(n3780), .A3(n3779), .A4(n3778), .ZN(n3782)
         );
  OAI21_X1 U4725 ( .B1(n3783), .B2(n3782), .A(n3961), .ZN(n3786) );
  NAND2_X1 U4726 ( .A1(n4131), .A2(EAX_REG_10__SCAN_IN), .ZN(n3785) );
  NAND2_X1 U4727 ( .A1(n4039), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3784)
         );
  NAND3_X1 U4728 ( .A1(n3786), .A2(n3785), .A3(n3784), .ZN(n3787) );
  AOI21_X1 U4729 ( .B1(n6156), .B2(n4165), .A(n3787), .ZN(n5079) );
  NOR2_X2 U4730 ( .A1(n5080), .A2(n5079), .ZN(n5081) );
  INV_X1 U4731 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3804) );
  XNOR2_X1 U4732 ( .A(n3805), .B(n3804), .ZN(n5180) );
  NAND2_X1 U4733 ( .A1(n5180), .A2(n4165), .ZN(n3803) );
  AOI22_X1 U4734 ( .A1(n4139), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4151), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3792) );
  AOI22_X1 U4735 ( .A1(n4148), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4149), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3791) );
  AOI22_X1 U4736 ( .A1(n4140), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4141), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3790) );
  AOI22_X1 U4737 ( .A1(n4150), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4142), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3789) );
  NAND4_X1 U4738 ( .A1(n3792), .A2(n3791), .A3(n3790), .A4(n3789), .ZN(n3798)
         );
  AOI22_X1 U4739 ( .A1(n4143), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3773), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3796) );
  AOI22_X1 U4740 ( .A1(n3546), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3795) );
  AOI22_X1 U4741 ( .A1(n4098), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3554), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3794) );
  AOI22_X1 U4742 ( .A1(n3545), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3158), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3793) );
  NAND4_X1 U4743 ( .A1(n3796), .A2(n3795), .A3(n3794), .A4(n3793), .ZN(n3797)
         );
  OAI21_X1 U4744 ( .B1(n3798), .B2(n3797), .A(n3961), .ZN(n3801) );
  NAND2_X1 U4745 ( .A1(n4131), .A2(EAX_REG_11__SCAN_IN), .ZN(n3800) );
  NAND2_X1 U4746 ( .A1(n4039), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3799)
         );
  AND3_X1 U4747 ( .A1(n3801), .A2(n3800), .A3(n3799), .ZN(n3802) );
  NAND2_X1 U4748 ( .A1(n3803), .A2(n3802), .ZN(n5115) );
  XOR2_X1 U4749 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .B(n3819), .Z(n6143) );
  AOI22_X1 U4750 ( .A1(n3545), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4149), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3809) );
  AOI22_X1 U4751 ( .A1(n4140), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n4143), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3808) );
  AOI22_X1 U4752 ( .A1(n3546), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n4141), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3807) );
  AOI22_X1 U4753 ( .A1(n4151), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n4098), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3806) );
  NAND4_X1 U4754 ( .A1(n3809), .A2(n3808), .A3(n3807), .A4(n3806), .ZN(n3815)
         );
  AOI22_X1 U4755 ( .A1(n4139), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4148), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3813) );
  AOI22_X1 U4756 ( .A1(n4150), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3812) );
  AOI22_X1 U4757 ( .A1(n3772), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n4142), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3811) );
  AOI22_X1 U4758 ( .A1(n3530), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3158), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3810) );
  NAND4_X1 U4759 ( .A1(n3813), .A2(n3812), .A3(n3811), .A4(n3810), .ZN(n3814)
         );
  OR2_X1 U4760 ( .A1(n3815), .A2(n3814), .ZN(n3816) );
  AOI22_X1 U4761 ( .A1(n3961), .A2(n3816), .B1(n4039), .B2(
        PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3818) );
  NAND2_X1 U4762 ( .A1(n4131), .A2(EAX_REG_12__SCAN_IN), .ZN(n3817) );
  OAI211_X1 U4763 ( .C1(n6143), .C2(n4163), .A(n3818), .B(n3817), .ZN(n5143)
         );
  INV_X1 U4764 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3853) );
  XNOR2_X1 U4765 ( .A(n3854), .B(n3853), .ZN(n6128) );
  NAND2_X1 U4766 ( .A1(n6128), .A2(n4165), .ZN(n3823) );
  NOR2_X1 U4767 ( .A1(n3820), .A2(n3853), .ZN(n3821) );
  AOI21_X1 U4768 ( .B1(n4131), .B2(EAX_REG_13__SCAN_IN), .A(n3821), .ZN(n3822)
         );
  NAND2_X1 U4769 ( .A1(n3823), .A2(n3822), .ZN(n3835) );
  XNOR2_X2 U4770 ( .A(n5145), .B(n3835), .ZN(n5273) );
  AOI22_X1 U4771 ( .A1(n4148), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4151), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3827) );
  AOI22_X1 U4772 ( .A1(n4139), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4140), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3826) );
  AOI22_X1 U4773 ( .A1(n3773), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4149), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3825) );
  AOI22_X1 U4774 ( .A1(n4143), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3158), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3824) );
  NAND4_X1 U4775 ( .A1(n3827), .A2(n3826), .A3(n3825), .A4(n3824), .ZN(n3833)
         );
  AOI22_X1 U4776 ( .A1(n3513), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3552), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3831) );
  AOI22_X1 U4777 ( .A1(n3545), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4142), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3830) );
  AOI22_X1 U4778 ( .A1(n4150), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4098), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3829) );
  AOI22_X1 U4779 ( .A1(n4141), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3554), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3828) );
  NAND4_X1 U4780 ( .A1(n3831), .A2(n3830), .A3(n3829), .A4(n3828), .ZN(n3832)
         );
  OR2_X1 U4781 ( .A1(n3833), .A2(n3832), .ZN(n3834) );
  AND2_X1 U4782 ( .A1(n3961), .A2(n3834), .ZN(n5272) );
  NAND2_X1 U4783 ( .A1(n5273), .A2(n5272), .ZN(n5271) );
  INV_X1 U4784 ( .A(n3835), .ZN(n3836) );
  NAND2_X1 U4785 ( .A1(n5271), .A2(n5619), .ZN(n5340) );
  NAND2_X1 U4786 ( .A1(n3464), .A2(n3421), .ZN(n3837) );
  OR2_X1 U4787 ( .A1(n3838), .A2(n3837), .ZN(n5348) );
  NAND2_X1 U4788 ( .A1(n4269), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4134) );
  AOI22_X1 U4789 ( .A1(n4143), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3842) );
  AOI22_X1 U4790 ( .A1(n4140), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4141), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3841) );
  AOI22_X1 U4791 ( .A1(n4149), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4142), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3840) );
  AOI22_X1 U4792 ( .A1(n4139), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4098), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3839) );
  NAND4_X1 U4793 ( .A1(n3842), .A2(n3841), .A3(n3840), .A4(n3839), .ZN(n3848)
         );
  AOI22_X1 U4794 ( .A1(n4150), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3546), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3846) );
  AOI22_X1 U4795 ( .A1(n4148), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3773), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3845) );
  AOI22_X1 U4796 ( .A1(n4151), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3554), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3844) );
  AOI22_X1 U4797 ( .A1(n3545), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3158), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3843) );
  NAND4_X1 U4798 ( .A1(n3846), .A2(n3845), .A3(n3844), .A4(n3843), .ZN(n3847)
         );
  NOR2_X1 U4799 ( .A1(n3848), .A2(n3847), .ZN(n3852) );
  NAND2_X1 U4800 ( .A1(n6636), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n3849)
         );
  NAND2_X1 U4801 ( .A1(n4163), .A2(n3849), .ZN(n3850) );
  AOI21_X1 U4802 ( .B1(n4131), .B2(EAX_REG_21__SCAN_IN), .A(n3850), .ZN(n3851)
         );
  OAI21_X1 U4803 ( .B1(n4134), .B2(n3852), .A(n3851), .ZN(n3860) );
  INV_X1 U4804 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3927) );
  INV_X1 U4805 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5819) );
  NOR2_X1 U4806 ( .A1(n3856), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n3857)
         );
  OR2_X1 U4807 ( .A1(n4021), .A2(n3857), .ZN(n6009) );
  INV_X1 U4808 ( .A(n6009), .ZN(n3858) );
  NAND2_X1 U4809 ( .A1(n3858), .A2(n4165), .ZN(n3859) );
  NAND2_X1 U4810 ( .A1(n3860), .A2(n3859), .ZN(n5651) );
  INV_X1 U4811 ( .A(n5651), .ZN(n3980) );
  AOI22_X1 U4812 ( .A1(n3546), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n4139), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3864) );
  AOI22_X1 U4813 ( .A1(n4148), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4143), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3863) );
  AOI22_X1 U4814 ( .A1(n3545), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3530), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3862) );
  AOI22_X1 U4815 ( .A1(n4149), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3158), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3861) );
  NAND4_X1 U4816 ( .A1(n3864), .A2(n3863), .A3(n3862), .A4(n3861), .ZN(n3872)
         );
  AOI22_X1 U4817 ( .A1(n4150), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3773), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3870) );
  AOI22_X1 U4818 ( .A1(n4140), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3869) );
  NAND2_X1 U4819 ( .A1(n4141), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3866)
         );
  NAND2_X1 U4820 ( .A1(n4098), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3865)
         );
  AND3_X1 U4821 ( .A1(n3866), .A2(n3865), .A3(n4163), .ZN(n3868) );
  AOI22_X1 U4822 ( .A1(n4151), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n4142), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3867) );
  NAND4_X1 U4823 ( .A1(n3870), .A2(n3869), .A3(n3868), .A4(n3867), .ZN(n3871)
         );
  NAND2_X1 U4824 ( .A1(n4134), .A2(n4163), .ZN(n3993) );
  OAI21_X1 U4825 ( .B1(n3872), .B2(n3871), .A(n3993), .ZN(n3875) );
  NOR2_X1 U4826 ( .A1(n5819), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3873) );
  AOI21_X1 U4827 ( .B1(n4131), .B2(EAX_REG_20__SCAN_IN), .A(n3873), .ZN(n3874)
         );
  NAND2_X1 U4828 ( .A1(n3875), .A2(n3874), .ZN(n3877) );
  XNOR2_X1 U4829 ( .A(n3892), .B(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n6013)
         );
  NAND2_X1 U4830 ( .A1(n6013), .A2(n4165), .ZN(n3876) );
  NAND2_X1 U4831 ( .A1(n3877), .A2(n3876), .ZN(n5662) );
  INV_X1 U4832 ( .A(n5662), .ZN(n3979) );
  AOI22_X1 U4833 ( .A1(n4139), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4149), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3881) );
  AOI22_X1 U4834 ( .A1(n4140), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4143), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3880) );
  AOI22_X1 U4835 ( .A1(n3546), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n4141), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3879) );
  AOI22_X1 U4836 ( .A1(n3545), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3554), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3878) );
  NAND4_X1 U4837 ( .A1(n3881), .A2(n3880), .A3(n3879), .A4(n3878), .ZN(n3887)
         );
  AOI22_X1 U4838 ( .A1(n4150), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3885) );
  AOI22_X1 U4839 ( .A1(n3773), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4142), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3884) );
  AOI22_X1 U4840 ( .A1(n4151), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4098), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3883) );
  AOI22_X1 U4841 ( .A1(n4148), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3158), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3882) );
  NAND4_X1 U4842 ( .A1(n3885), .A2(n3884), .A3(n3883), .A4(n3882), .ZN(n3886)
         );
  NOR2_X1 U4843 ( .A1(n3887), .A2(n3886), .ZN(n3891) );
  NAND2_X1 U4844 ( .A1(n6636), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3888)
         );
  NAND2_X1 U4845 ( .A1(n4163), .A2(n3888), .ZN(n3889) );
  AOI21_X1 U4846 ( .B1(n4131), .B2(EAX_REG_19__SCAN_IN), .A(n3889), .ZN(n3890)
         );
  OAI21_X1 U4847 ( .B1(n4134), .B2(n3891), .A(n3890), .ZN(n3895) );
  OAI21_X1 U4848 ( .B1(n3893), .B2(PHYADDRPOINTER_REG_19__SCAN_IN), .A(n3892), 
        .ZN(n5825) );
  OR2_X1 U4849 ( .A1(n5825), .A2(n4163), .ZN(n3894) );
  AND2_X1 U4850 ( .A1(n3895), .A2(n3894), .ZN(n5343) );
  AOI22_X1 U4851 ( .A1(n4148), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3899) );
  AOI22_X1 U4852 ( .A1(n4143), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4141), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3898) );
  AOI22_X1 U4853 ( .A1(n4142), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n4098), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3897) );
  AOI22_X1 U4854 ( .A1(n4150), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3530), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3896) );
  NAND4_X1 U4855 ( .A1(n3899), .A2(n3898), .A3(n3897), .A4(n3896), .ZN(n3907)
         );
  AOI22_X1 U4856 ( .A1(n3545), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4151), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3905) );
  NAND2_X1 U4857 ( .A1(n3546), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3901) );
  NAND2_X1 U4858 ( .A1(n4139), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3900) );
  AND3_X1 U4859 ( .A1(n3901), .A2(n3900), .A3(n4163), .ZN(n3904) );
  AOI22_X1 U4860 ( .A1(n4140), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4149), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3903) );
  AOI22_X1 U4861 ( .A1(n3773), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3158), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3902) );
  NAND4_X1 U4862 ( .A1(n3905), .A2(n3904), .A3(n3903), .A4(n3902), .ZN(n3906)
         );
  OAI21_X1 U4863 ( .B1(n3907), .B2(n3906), .A(n3993), .ZN(n3909) );
  AOI22_X1 U4864 ( .A1(n4131), .A2(EAX_REG_18__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n6636), .ZN(n3908) );
  NAND2_X1 U4865 ( .A1(n3909), .A2(n3908), .ZN(n3911) );
  XNOR2_X1 U4866 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .B(n3957), .ZN(n5835)
         );
  NAND2_X1 U4867 ( .A1(n4165), .A2(n5835), .ZN(n3910) );
  NAND2_X1 U4868 ( .A1(n3911), .A2(n3910), .ZN(n5589) );
  INV_X1 U4869 ( .A(n5589), .ZN(n3978) );
  XNOR2_X1 U4870 ( .A(n3912), .B(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5600)
         );
  AOI22_X1 U4871 ( .A1(n4139), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3545), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3916) );
  AOI22_X1 U4872 ( .A1(INSTQUEUE_REG_5__0__SCAN_IN), .A2(n4140), .B1(n3546), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3915) );
  AOI22_X1 U4873 ( .A1(INSTQUEUE_REG_12__0__SCAN_IN), .A2(n4148), .B1(n4103), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3914) );
  AOI22_X1 U4874 ( .A1(n4151), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3158), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3913) );
  NAND4_X1 U4875 ( .A1(n3916), .A2(n3915), .A3(n3914), .A4(n3913), .ZN(n3922)
         );
  AOI22_X1 U4876 ( .A1(n3773), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4149), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3920) );
  AOI22_X1 U4877 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n4150), .B1(n4141), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3919) );
  AOI22_X1 U4878 ( .A1(n4143), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n4142), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3918) );
  AOI22_X1 U4879 ( .A1(n4098), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3554), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3917) );
  NAND4_X1 U4880 ( .A1(n3920), .A2(n3919), .A3(n3918), .A4(n3917), .ZN(n3921)
         );
  NOR2_X1 U4881 ( .A1(n3922), .A2(n3921), .ZN(n3924) );
  AOI22_X1 U4882 ( .A1(n4131), .A2(EAX_REG_16__SCAN_IN), .B1(n4039), .B2(
        PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3923) );
  OAI21_X1 U4883 ( .B1(n4134), .B2(n3924), .A(n3923), .ZN(n3925) );
  AOI21_X1 U4884 ( .B1(n5600), .B2(n4165), .A(n3925), .ZN(n5383) );
  XOR2_X1 U4885 ( .A(n3927), .B(n3926), .Z(n5842) );
  INV_X1 U4886 ( .A(n5842), .ZN(n3942) );
  AOI22_X1 U4887 ( .A1(n3545), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4151), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3931) );
  AOI22_X1 U4888 ( .A1(n4139), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4149), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3930) );
  AOI22_X1 U4889 ( .A1(n4140), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3773), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3929) );
  AOI22_X1 U4890 ( .A1(n3546), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n4141), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3928) );
  NAND4_X1 U4891 ( .A1(n3931), .A2(n3930), .A3(n3929), .A4(n3928), .ZN(n3937)
         );
  AOI22_X1 U4892 ( .A1(n4150), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3935) );
  AOI22_X1 U4893 ( .A1(n4143), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4142), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3934) );
  AOI22_X1 U4894 ( .A1(n4098), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3530), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3933) );
  AOI22_X1 U4895 ( .A1(n4148), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3158), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3932) );
  NAND4_X1 U4896 ( .A1(n3935), .A2(n3934), .A3(n3933), .A4(n3932), .ZN(n3936)
         );
  OAI21_X1 U4897 ( .B1(n3937), .B2(n3936), .A(n3961), .ZN(n3940) );
  NAND2_X1 U4898 ( .A1(n4131), .A2(EAX_REG_15__SCAN_IN), .ZN(n3939) );
  NAND2_X1 U4899 ( .A1(n4039), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3938)
         );
  NAND3_X1 U4900 ( .A1(n3940), .A2(n3939), .A3(n3938), .ZN(n3941) );
  AOI21_X1 U4901 ( .B1(n3942), .B2(n4165), .A(n3941), .ZN(n5608) );
  OR2_X1 U4902 ( .A1(n5383), .A2(n5608), .ZN(n5381) );
  AOI22_X1 U4903 ( .A1(n4150), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4140), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3946) );
  AOI22_X1 U4904 ( .A1(n3546), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n4141), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3945) );
  AOI22_X1 U4905 ( .A1(n4151), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3530), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3944) );
  AOI22_X1 U4906 ( .A1(n4139), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3158), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3943) );
  NAND4_X1 U4907 ( .A1(n3946), .A2(n3945), .A3(n3944), .A4(n3943), .ZN(n3952)
         );
  AOI22_X1 U4908 ( .A1(n4148), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4149), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3950) );
  AOI22_X1 U4909 ( .A1(n4143), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3949) );
  AOI22_X1 U4910 ( .A1(n3773), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4142), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3948) );
  AOI22_X1 U4911 ( .A1(n3545), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4098), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3947) );
  NAND4_X1 U4912 ( .A1(n3950), .A2(n3949), .A3(n3948), .A4(n3947), .ZN(n3951)
         );
  NOR2_X1 U4913 ( .A1(n3952), .A2(n3951), .ZN(n3956) );
  NAND2_X1 U4914 ( .A1(n6636), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n3953)
         );
  NAND2_X1 U4915 ( .A1(n4163), .A2(n3953), .ZN(n3954) );
  AOI21_X1 U4916 ( .B1(n4131), .B2(EAX_REG_17__SCAN_IN), .A(n3954), .ZN(n3955)
         );
  OAI21_X1 U4917 ( .B1(n4134), .B2(n3956), .A(n3955), .ZN(n3960) );
  OAI21_X1 U4918 ( .B1(PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n3958), .A(n3957), 
        .ZN(n6115) );
  OR2_X1 U4919 ( .A1(n4163), .A2(n6115), .ZN(n3959) );
  NAND2_X1 U4920 ( .A1(n3960), .A2(n3959), .ZN(n5672) );
  NOR2_X1 U4921 ( .A1(n5381), .A2(n5672), .ZN(n3977) );
  INV_X1 U4922 ( .A(n3961), .ZN(n3976) );
  AOI22_X1 U4923 ( .A1(n4139), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3545), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3965) );
  AOI22_X1 U4924 ( .A1(n4143), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4149), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3964) );
  AOI22_X1 U4925 ( .A1(n4150), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4141), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3963) );
  AOI22_X1 U4926 ( .A1(n3554), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3158), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3962) );
  NAND4_X1 U4927 ( .A1(n3965), .A2(n3964), .A3(n3963), .A4(n3962), .ZN(n3971)
         );
  AOI22_X1 U4928 ( .A1(n3546), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n4140), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3969) );
  AOI22_X1 U4929 ( .A1(n4148), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3773), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3968) );
  AOI22_X1 U4930 ( .A1(n4103), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4142), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3967) );
  AOI22_X1 U4931 ( .A1(n4151), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n4098), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3966) );
  NAND4_X1 U4932 ( .A1(n3969), .A2(n3968), .A3(n3967), .A4(n3966), .ZN(n3970)
         );
  NOR2_X1 U4933 ( .A1(n3971), .A2(n3970), .ZN(n3975) );
  XNOR2_X1 U4934 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .B(n3972), .ZN(n5853)
         );
  AOI22_X1 U4935 ( .A1(n4165), .A2(n5853), .B1(n4039), .B2(
        PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3974) );
  NAND2_X1 U4936 ( .A1(n4131), .A2(EAX_REG_14__SCAN_IN), .ZN(n3973) );
  OAI211_X1 U4937 ( .C1(n3976), .C2(n3975), .A(n3974), .B(n3973), .ZN(n5620)
         );
  AND2_X1 U4938 ( .A1(n3977), .A2(n5620), .ZN(n5587) );
  AND2_X1 U4939 ( .A1(n3978), .A2(n5587), .ZN(n5341) );
  AOI22_X1 U4940 ( .A1(n4150), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4139), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3985) );
  AOI22_X1 U4941 ( .A1(n4103), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4141), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3984) );
  AOI22_X1 U4942 ( .A1(n3773), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4098), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3983) );
  AOI22_X1 U4943 ( .A1(n4140), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3530), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3982) );
  NAND4_X1 U4944 ( .A1(n3985), .A2(n3984), .A3(n3983), .A4(n3982), .ZN(n3995)
         );
  INV_X1 U4945 ( .A(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3988) );
  AOI22_X1 U4946 ( .A1(n4143), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n4149), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3987) );
  AOI21_X1 U4947 ( .B1(n3545), .B2(INSTQUEUE_REG_8__6__SCAN_IN), .A(n4165), 
        .ZN(n3986) );
  OAI211_X1 U4948 ( .C1(n3535), .C2(n3988), .A(n3987), .B(n3986), .ZN(n3989)
         );
  INV_X1 U4949 ( .A(n3989), .ZN(n3992) );
  AOI22_X1 U4950 ( .A1(n4148), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4151), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3991) );
  AOI22_X1 U4951 ( .A1(n4142), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3158), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3990) );
  NAND3_X1 U4952 ( .A1(n3992), .A2(n3991), .A3(n3990), .ZN(n3994) );
  OAI21_X1 U4953 ( .B1(n3995), .B2(n3994), .A(n3993), .ZN(n3997) );
  AOI22_X1 U4954 ( .A1(n4131), .A2(EAX_REG_22__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n6636), .ZN(n3996) );
  XOR2_X1 U4955 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .B(n4021), .Z(n5808) );
  AOI22_X1 U4956 ( .A1(n3997), .A2(n3996), .B1(n4165), .B2(n5808), .ZN(n5570)
         );
  AOI22_X1 U4957 ( .A1(INSTQUEUE_REG_6__0__SCAN_IN), .A2(n4140), .B1(n4103), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4001) );
  AOI22_X1 U4958 ( .A1(n3546), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n4141), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n4000) );
  AOI22_X1 U4959 ( .A1(INSTQUEUE_REG_5__0__SCAN_IN), .A2(n4151), .B1(n3554), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3999) );
  AOI22_X1 U4960 ( .A1(n3545), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3158), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3998) );
  NAND4_X1 U4961 ( .A1(n4001), .A2(n4000), .A3(n3999), .A4(n3998), .ZN(n4007)
         );
  AOI22_X1 U4962 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n4148), .B1(n4149), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n4005) );
  AOI22_X1 U4963 ( .A1(n4150), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4143), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4004) );
  AOI22_X1 U4964 ( .A1(n3773), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4142), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4003) );
  AOI22_X1 U4965 ( .A1(n4139), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4098), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4002) );
  NAND4_X1 U4966 ( .A1(n4005), .A2(n4004), .A3(n4003), .A4(n4002), .ZN(n4006)
         );
  NOR2_X1 U4967 ( .A1(n4007), .A2(n4006), .ZN(n4037) );
  AOI22_X1 U4968 ( .A1(n3773), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4149), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n4011) );
  AOI22_X1 U4969 ( .A1(n4143), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n4141), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4010) );
  AOI22_X1 U4970 ( .A1(n4151), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3530), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4009) );
  AOI22_X1 U4971 ( .A1(n4098), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3158), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4008) );
  NAND4_X1 U4972 ( .A1(n4011), .A2(n4010), .A3(n4009), .A4(n4008), .ZN(n4017)
         );
  AOI22_X1 U4973 ( .A1(n4139), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3545), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4015) );
  AOI22_X1 U4974 ( .A1(n3546), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n4140), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4014) );
  AOI22_X1 U4975 ( .A1(n4150), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4013) );
  AOI22_X1 U4976 ( .A1(n4148), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4142), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4012) );
  NAND4_X1 U4977 ( .A1(n4015), .A2(n4014), .A3(n4013), .A4(n4012), .ZN(n4016)
         );
  NOR2_X1 U4978 ( .A1(n4017), .A2(n4016), .ZN(n4036) );
  XNOR2_X1 U4979 ( .A(n4037), .B(n4036), .ZN(n4018) );
  NOR2_X1 U4980 ( .A1(n4134), .A2(n4018), .ZN(n4025) );
  INV_X1 U4981 ( .A(EAX_REG_23__SCAN_IN), .ZN(n6256) );
  NOR2_X1 U4982 ( .A1(n6999), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4019)
         );
  OAI22_X1 U4983 ( .A1(n4020), .A2(n6256), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4019), .ZN(n4024) );
  OR2_X1 U4984 ( .A1(n4022), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4023)
         );
  NAND2_X1 U4985 ( .A1(n4042), .A2(n4023), .ZN(n5996) );
  OAI22_X1 U4986 ( .A1(n4025), .A2(n4024), .B1(n4163), .B2(n5996), .ZN(n5797)
         );
  NOR2_X2 U4987 ( .A1(n5569), .A2(n5797), .ZN(n5559) );
  XNOR2_X1 U4988 ( .A(n4042), .B(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5785)
         );
  AOI22_X1 U4989 ( .A1(n4143), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4029) );
  AOI22_X1 U4990 ( .A1(n4150), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4140), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4028) );
  AOI22_X1 U4991 ( .A1(n3546), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n4141), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n4027) );
  AOI22_X1 U4992 ( .A1(n3773), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4142), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4026) );
  NAND4_X1 U4993 ( .A1(n4029), .A2(n4028), .A3(n4027), .A4(n4026), .ZN(n4035)
         );
  AOI22_X1 U4994 ( .A1(n4139), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3545), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n4033) );
  AOI22_X1 U4995 ( .A1(n4148), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4149), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4032) );
  AOI22_X1 U4996 ( .A1(n4151), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3530), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4031) );
  AOI22_X1 U4997 ( .A1(n4098), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n3158), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4030) );
  NAND4_X1 U4998 ( .A1(n4033), .A2(n4032), .A3(n4031), .A4(n4030), .ZN(n4034)
         );
  OR2_X1 U4999 ( .A1(n4035), .A2(n4034), .ZN(n4056) );
  NOR2_X1 U5000 ( .A1(n4037), .A2(n4036), .ZN(n4057) );
  XOR2_X1 U5001 ( .A(n4056), .B(n4057), .Z(n4038) );
  INV_X1 U5002 ( .A(n4134), .ZN(n4160) );
  NAND2_X1 U5003 ( .A1(n4038), .A2(n4160), .ZN(n4041) );
  AOI22_X1 U5004 ( .A1(n4131), .A2(EAX_REG_24__SCAN_IN), .B1(n4039), .B2(
        PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4040) );
  OAI211_X1 U5005 ( .C1(n5785), .C2(n4163), .A(n4041), .B(n4040), .ZN(n5560)
         );
  NAND2_X1 U5006 ( .A1(n5559), .A2(n5560), .ZN(n5543) );
  INV_X1 U5007 ( .A(n4042), .ZN(n4043) );
  NAND2_X1 U5008 ( .A1(n4043), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4044)
         );
  INV_X1 U5009 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5553) );
  NAND2_X1 U5010 ( .A1(n4044), .A2(n5553), .ZN(n4045) );
  NAND2_X1 U5011 ( .A1(n4078), .A2(n4045), .ZN(n5771) );
  AOI22_X1 U5012 ( .A1(n3545), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4149), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4049) );
  AOI22_X1 U5013 ( .A1(n4140), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3773), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4048) );
  AOI22_X1 U5014 ( .A1(n3513), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n4141), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n4047) );
  AOI22_X1 U5015 ( .A1(n4098), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3158), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4046) );
  NAND4_X1 U5016 ( .A1(n4049), .A2(n4048), .A3(n4047), .A4(n4046), .ZN(n4055)
         );
  AOI22_X1 U5017 ( .A1(n4139), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4148), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n4053) );
  AOI22_X1 U5018 ( .A1(n4150), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3552), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4052) );
  AOI22_X1 U5019 ( .A1(n4143), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4142), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4051) );
  AOI22_X1 U5020 ( .A1(n4151), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3530), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4050) );
  NAND4_X1 U5021 ( .A1(n4053), .A2(n4052), .A3(n4051), .A4(n4050), .ZN(n4054)
         );
  NOR2_X1 U5022 ( .A1(n4055), .A2(n4054), .ZN(n4073) );
  NAND2_X1 U5023 ( .A1(n4057), .A2(n4056), .ZN(n4072) );
  XNOR2_X1 U5024 ( .A(n4073), .B(n4072), .ZN(n4060) );
  AOI21_X1 U5025 ( .B1(PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n6636), .A(n4165), 
        .ZN(n4059) );
  NAND2_X1 U5026 ( .A1(n4131), .A2(EAX_REG_25__SCAN_IN), .ZN(n4058) );
  OAI211_X1 U5027 ( .C1(n4060), .C2(n4134), .A(n4059), .B(n4058), .ZN(n4061)
         );
  OAI21_X1 U5028 ( .B1(n4163), .B2(n5771), .A(n4061), .ZN(n5545) );
  AOI22_X1 U5029 ( .A1(n4143), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3552), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4065) );
  AOI22_X1 U5030 ( .A1(n4150), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4140), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4064) );
  AOI22_X1 U5031 ( .A1(n3513), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n4141), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n4063) );
  AOI22_X1 U5032 ( .A1(n3773), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4142), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4062) );
  NAND4_X1 U5033 ( .A1(n4065), .A2(n4064), .A3(n4063), .A4(n4062), .ZN(n4071)
         );
  AOI22_X1 U5034 ( .A1(n4139), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3545), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n4069) );
  AOI22_X1 U5035 ( .A1(n4148), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4149), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4068) );
  AOI22_X1 U5036 ( .A1(n4151), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3554), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4067) );
  AOI22_X1 U5037 ( .A1(n4098), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3158), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4066) );
  NAND4_X1 U5038 ( .A1(n4069), .A2(n4068), .A3(n4067), .A4(n4066), .ZN(n4070)
         );
  OR2_X1 U5039 ( .A1(n4071), .A2(n4070), .ZN(n4092) );
  NOR2_X1 U5040 ( .A1(n4073), .A2(n4072), .ZN(n4093) );
  XOR2_X1 U5041 ( .A(n4092), .B(n4093), .Z(n4074) );
  NAND2_X1 U5042 ( .A1(n4074), .A2(n4160), .ZN(n4077) );
  INV_X1 U5043 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5765) );
  NOR2_X1 U5044 ( .A1(n5765), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4075) );
  AOI211_X1 U5045 ( .C1(n4131), .C2(EAX_REG_26__SCAN_IN), .A(n4165), .B(n4075), 
        .ZN(n4076) );
  XNOR2_X1 U5046 ( .A(n4078), .B(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5769)
         );
  AOI22_X1 U5047 ( .A1(n4077), .A2(n4076), .B1(n4165), .B2(n5769), .ZN(n5531)
         );
  NAND2_X1 U5048 ( .A1(n5529), .A2(n5531), .ZN(n5514) );
  INV_X1 U5049 ( .A(n4079), .ZN(n4080) );
  INV_X1 U5050 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5521) );
  NAND2_X1 U5051 ( .A1(n4080), .A2(n5521), .ZN(n4081) );
  NAND2_X1 U5052 ( .A1(n4116), .A2(n4081), .ZN(n5757) );
  AOI22_X1 U5053 ( .A1(n3552), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4149), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4085) );
  AOI22_X1 U5054 ( .A1(n4150), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4140), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4084) );
  AOI22_X1 U5055 ( .A1(n3513), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n4141), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n4083) );
  AOI22_X1 U5056 ( .A1(n3545), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3554), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4082) );
  NAND4_X1 U5057 ( .A1(n4085), .A2(n4084), .A3(n4083), .A4(n4082), .ZN(n4091)
         );
  AOI22_X1 U5058 ( .A1(n4148), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3773), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4089) );
  AOI22_X1 U5059 ( .A1(n4143), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n4142), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4088) );
  AOI22_X1 U5060 ( .A1(n4151), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4098), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4087) );
  AOI22_X1 U5061 ( .A1(n4139), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3158), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4086) );
  NAND4_X1 U5062 ( .A1(n4089), .A2(n4088), .A3(n4087), .A4(n4086), .ZN(n4090)
         );
  NOR2_X1 U5063 ( .A1(n4091), .A2(n4090), .ZN(n4111) );
  NAND2_X1 U5064 ( .A1(n4093), .A2(n4092), .ZN(n4110) );
  XNOR2_X1 U5065 ( .A(n4111), .B(n4110), .ZN(n4096) );
  AOI21_X1 U5066 ( .B1(PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n6636), .A(n4165), 
        .ZN(n4095) );
  NAND2_X1 U5067 ( .A1(n4131), .A2(EAX_REG_27__SCAN_IN), .ZN(n4094) );
  OAI211_X1 U5068 ( .C1(n4096), .C2(n4134), .A(n4095), .B(n4094), .ZN(n4097)
         );
  OAI21_X1 U5069 ( .B1(n4163), .B2(n5757), .A(n4097), .ZN(n5516) );
  NOR2_X2 U5070 ( .A1(n5514), .A2(n5516), .ZN(n5515) );
  AOI22_X1 U5071 ( .A1(n4139), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3545), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n4102) );
  AOI22_X1 U5072 ( .A1(n4148), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4149), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4101) );
  AOI22_X1 U5073 ( .A1(n4151), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3530), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4100) );
  AOI22_X1 U5074 ( .A1(n4098), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3158), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4099) );
  NAND4_X1 U5075 ( .A1(n4102), .A2(n4101), .A3(n4100), .A4(n4099), .ZN(n4109)
         );
  AOI22_X1 U5076 ( .A1(n4143), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4107) );
  AOI22_X1 U5077 ( .A1(n4150), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4140), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4106) );
  AOI22_X1 U5078 ( .A1(n3513), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n4141), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n4105) );
  AOI22_X1 U5079 ( .A1(n3773), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4142), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4104) );
  NAND4_X1 U5080 ( .A1(n4107), .A2(n4106), .A3(n4105), .A4(n4104), .ZN(n4108)
         );
  OR2_X1 U5081 ( .A1(n4109), .A2(n4108), .ZN(n4129) );
  NOR2_X1 U5082 ( .A1(n4111), .A2(n4110), .ZN(n4130) );
  XOR2_X1 U5083 ( .A(n4129), .B(n4130), .Z(n4112) );
  NAND2_X1 U5084 ( .A1(n4112), .A2(n4160), .ZN(n4115) );
  INV_X1 U5085 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5746) );
  NOR2_X1 U5086 ( .A1(n5746), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4113) );
  AOI211_X1 U5087 ( .C1(n4131), .C2(EAX_REG_28__SCAN_IN), .A(n4165), .B(n4113), 
        .ZN(n4114) );
  XNOR2_X1 U5088 ( .A(n4116), .B(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5750)
         );
  AOI22_X1 U5089 ( .A1(n4115), .A2(n4114), .B1(n4165), .B2(n5750), .ZN(n5502)
         );
  NAND2_X1 U5090 ( .A1(n5515), .A2(n5502), .ZN(n5501) );
  INV_X1 U5091 ( .A(n4117), .ZN(n4118) );
  INV_X1 U5092 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5494) );
  OAI21_X1 U5093 ( .B1(n4118), .B2(PHYADDRPOINTER_REG_29__SCAN_IN), .A(n4171), 
        .ZN(n5737) );
  AOI22_X1 U5094 ( .A1(n4150), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4141), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n4122) );
  AOI22_X1 U5095 ( .A1(n4103), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4142), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4121) );
  AOI22_X1 U5096 ( .A1(n4151), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3554), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4120) );
  AOI22_X1 U5097 ( .A1(n4148), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3158), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4119) );
  NAND4_X1 U5098 ( .A1(n4122), .A2(n4121), .A3(n4120), .A4(n4119), .ZN(n4128)
         );
  AOI22_X1 U5099 ( .A1(n4139), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4149), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4126) );
  AOI22_X1 U5100 ( .A1(n3513), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n4140), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4125) );
  AOI22_X1 U5101 ( .A1(n4143), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3773), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4124) );
  AOI22_X1 U5102 ( .A1(n3545), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4098), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4123) );
  NAND4_X1 U5103 ( .A1(n4126), .A2(n4125), .A3(n4124), .A4(n4123), .ZN(n4127)
         );
  NOR2_X1 U5104 ( .A1(n4128), .A2(n4127), .ZN(n4138) );
  NAND2_X1 U5105 ( .A1(n4130), .A2(n4129), .ZN(n4137) );
  XNOR2_X1 U5106 ( .A(n4138), .B(n4137), .ZN(n4135) );
  AOI21_X1 U5107 ( .B1(PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n6636), .A(n4165), 
        .ZN(n4133) );
  NAND2_X1 U5108 ( .A1(n4131), .A2(EAX_REG_29__SCAN_IN), .ZN(n4132) );
  OAI211_X1 U5109 ( .C1(n4135), .C2(n4134), .A(n4133), .B(n4132), .ZN(n4136)
         );
  OAI21_X1 U5110 ( .B1(n4163), .B2(n5737), .A(n4136), .ZN(n5487) );
  NOR2_X2 U5111 ( .A1(n5501), .A2(n5487), .ZN(n5486) );
  NOR2_X1 U5112 ( .A1(n4138), .A2(n4137), .ZN(n4159) );
  AOI22_X1 U5113 ( .A1(n4139), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3773), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4147) );
  AOI22_X1 U5114 ( .A1(n4140), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3552), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4146) );
  AOI22_X1 U5115 ( .A1(n3513), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n4141), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n4145) );
  AOI22_X1 U5116 ( .A1(n4143), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n4142), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4144) );
  NAND4_X1 U5117 ( .A1(n4147), .A2(n4146), .A3(n4145), .A4(n4144), .ZN(n4157)
         );
  AOI22_X1 U5118 ( .A1(n3545), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4148), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n4155) );
  AOI22_X1 U5119 ( .A1(n4150), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4149), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4154) );
  AOI22_X1 U5120 ( .A1(n4151), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3530), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4153) );
  AOI22_X1 U5121 ( .A1(n4098), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3158), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4152) );
  NAND4_X1 U5122 ( .A1(n4155), .A2(n4154), .A3(n4153), .A4(n4152), .ZN(n4156)
         );
  NOR2_X1 U5123 ( .A1(n4157), .A2(n4156), .ZN(n4158) );
  XNOR2_X1 U5124 ( .A(n4159), .B(n4158), .ZN(n4161) );
  NAND2_X1 U5125 ( .A1(n4161), .A2(n4160), .ZN(n4168) );
  NAND2_X1 U5126 ( .A1(n6636), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4162)
         );
  NAND2_X1 U5127 ( .A1(n4163), .A2(n4162), .ZN(n4164) );
  AOI21_X1 U5128 ( .B1(n4131), .B2(EAX_REG_30__SCAN_IN), .A(n4164), .ZN(n4167)
         );
  XNOR2_X1 U5129 ( .A(n4171), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5449)
         );
  AND2_X1 U5130 ( .A1(n5449), .A2(n4165), .ZN(n4166) );
  AOI21_X1 U5131 ( .B1(n4168), .B2(n4167), .A(n4166), .ZN(n4192) );
  NAND2_X1 U5132 ( .A1(n5486), .A2(n4192), .ZN(n4169) );
  XOR2_X1 U5133 ( .A(n4170), .B(n4169), .Z(n5730) );
  INV_X1 U5134 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5452) );
  NOR2_X1 U5135 ( .A1(n5728), .A2(n6645), .ZN(n4173) );
  NAND3_X1 U5136 ( .A1(n4176), .A2(n4175), .A3(n4174), .ZN(U2796) );
  INV_X1 U5137 ( .A(n4181), .ZN(n4178) );
  AOI211_X1 U5138 ( .C1(n5506), .C2(n4179), .A(n4178), .B(n4177), .ZN(n4184)
         );
  AOI211_X1 U5139 ( .C1(n5344), .C2(n4182), .A(n4181), .B(n4180), .ZN(n4183)
         );
  NOR2_X1 U5140 ( .A1(n4184), .A2(n4183), .ZN(n5445) );
  AOI22_X1 U5141 ( .A1(PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n6194), .B1(n6193), 
        .B2(n5449), .ZN(n4191) );
  INV_X1 U5142 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5637) );
  AND3_X1 U5143 ( .A1(n3348), .A2(n5637), .A3(n4186), .ZN(n4187) );
  NOR2_X1 U5144 ( .A1(n4188), .A2(n4187), .ZN(n4189) );
  NAND2_X1 U5145 ( .A1(n6191), .A2(EBX_REG_30__SCAN_IN), .ZN(n4190) );
  OAI211_X1 U5146 ( .C1(n5445), .C2(n6198), .A(n4191), .B(n4190), .ZN(n4199)
         );
  INV_X1 U5147 ( .A(n5499), .ZN(n4194) );
  INV_X1 U5148 ( .A(REIP_REG_29__SCAN_IN), .ZN(n7100) );
  INV_X1 U5149 ( .A(REIP_REG_30__SCAN_IN), .ZN(n4193) );
  OAI21_X1 U5150 ( .B1(n4194), .B2(n7100), .A(n4193), .ZN(n4196) );
  OAI21_X1 U5151 ( .B1(n5701), .B2(n6157), .A(n4197), .ZN(n4198) );
  OR2_X1 U5152 ( .A1(n4199), .A2(n4198), .ZN(U2797) );
  NOR2_X1 U5153 ( .A1(n6645), .A2(n6636), .ZN(n4474) );
  NOR2_X1 U5154 ( .A1(n5476), .A2(n3451), .ZN(n5355) );
  INV_X1 U5155 ( .A(n5355), .ZN(n4338) );
  INV_X1 U5156 ( .A(n4352), .ZN(n4201) );
  NAND2_X1 U5157 ( .A1(n4201), .A2(n6240), .ZN(n6633) );
  AOI21_X1 U5158 ( .B1(n4338), .B2(n6633), .A(n6662), .ZN(n4202) );
  AND2_X1 U5159 ( .A1(n6229), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  OR2_X1 U5160 ( .A1(n6240), .A2(n4203), .ZN(n5485) );
  INV_X1 U5161 ( .A(n4204), .ZN(n6239) );
  OR2_X1 U5162 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6537) );
  INV_X1 U5163 ( .A(n6537), .ZN(n6530) );
  AND2_X1 U5164 ( .A1(n6530), .A2(n6645), .ZN(n5102) );
  NOR2_X1 U5165 ( .A1(n6239), .A2(n5102), .ZN(n5993) );
  INV_X1 U5166 ( .A(n5993), .ZN(n4206) );
  INV_X1 U5167 ( .A(n4205), .ZN(n5994) );
  NOR3_X1 U5168 ( .A1(n4206), .A2(n5994), .A3(READREQUEST_REG_SCAN_IN), .ZN(
        n4207) );
  AOI21_X1 U5169 ( .B1(n6721), .B2(n5485), .A(n4207), .ZN(U3474) );
  INV_X1 U5170 ( .A(EAX_REG_24__SCAN_IN), .ZN(n6258) );
  NAND2_X1 U5171 ( .A1(n6217), .A2(n3348), .ZN(n4336) );
  AOI22_X1 U5172 ( .A1(n4333), .A2(UWORD_REG_8__SCAN_IN), .B1(n6234), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4208) );
  OAI21_X1 U5173 ( .B1(n6258), .B2(n4336), .A(n4208), .ZN(U2899) );
  INV_X1 U5174 ( .A(EAX_REG_25__SCAN_IN), .ZN(n6260) );
  AOI22_X1 U5175 ( .A1(n4333), .A2(UWORD_REG_9__SCAN_IN), .B1(n6234), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4209) );
  OAI21_X1 U5176 ( .B1(n6260), .B2(n4336), .A(n4209), .ZN(U2898) );
  INV_X1 U5177 ( .A(EAX_REG_27__SCAN_IN), .ZN(n6265) );
  AOI22_X1 U5178 ( .A1(n4333), .A2(UWORD_REG_11__SCAN_IN), .B1(n6234), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n4210) );
  OAI21_X1 U5179 ( .B1(n6265), .B2(n4336), .A(n4210), .ZN(U2896) );
  INV_X1 U5180 ( .A(EAX_REG_28__SCAN_IN), .ZN(n6268) );
  AOI22_X1 U5181 ( .A1(n4333), .A2(UWORD_REG_12__SCAN_IN), .B1(n6234), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n4211) );
  OAI21_X1 U5182 ( .B1(n6268), .B2(n4336), .A(n4211), .ZN(U2895) );
  INV_X1 U5183 ( .A(EAX_REG_29__SCAN_IN), .ZN(n6270) );
  AOI22_X1 U5184 ( .A1(n4333), .A2(UWORD_REG_13__SCAN_IN), .B1(n6234), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n4212) );
  OAI21_X1 U5185 ( .B1(n6270), .B2(n4336), .A(n4212), .ZN(U2894) );
  INV_X1 U5186 ( .A(EAX_REG_26__SCAN_IN), .ZN(n6263) );
  AOI22_X1 U5187 ( .A1(n4333), .A2(UWORD_REG_10__SCAN_IN), .B1(n6234), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n4213) );
  OAI21_X1 U5188 ( .B1(n6263), .B2(n4336), .A(n4213), .ZN(U2897) );
  INV_X1 U5189 ( .A(EAX_REG_30__SCAN_IN), .ZN(n6274) );
  AOI22_X1 U5190 ( .A1(n4333), .A2(UWORD_REG_14__SCAN_IN), .B1(n6234), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n4214) );
  OAI21_X1 U5191 ( .B1(n6274), .B2(n4336), .A(n4214), .ZN(U2893) );
  NAND2_X1 U5192 ( .A1(n5348), .A2(n4498), .ZN(n4215) );
  AND2_X1 U5193 ( .A1(n4264), .A2(n4215), .ZN(n4250) );
  AND2_X1 U5194 ( .A1(n4250), .A2(n4216), .ZN(n6602) );
  INV_X1 U5195 ( .A(n4217), .ZN(n4219) );
  INV_X1 U5196 ( .A(n4290), .ZN(n4218) );
  NAND2_X1 U5197 ( .A1(n4219), .A2(n4218), .ZN(n4223) );
  INV_X1 U5198 ( .A(n6240), .ZN(n6723) );
  INV_X1 U5199 ( .A(n4220), .ZN(n4416) );
  OAI21_X1 U5200 ( .B1(n6723), .B2(n4292), .A(n4416), .ZN(n4221) );
  INV_X1 U5201 ( .A(n4221), .ZN(n4222) );
  NAND2_X1 U5202 ( .A1(n4223), .A2(n4222), .ZN(n4287) );
  XOR2_X1 U5203 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .B(n4287), .Z(n4280) );
  NAND2_X1 U5204 ( .A1(n4225), .A2(n4224), .ZN(n4226) );
  NAND2_X1 U5205 ( .A1(n4227), .A2(n4226), .ZN(n5133) );
  NAND3_X1 U5206 ( .A1(n6644), .A2(STATEBS16_REG_SCAN_IN), .A3(
        STATE2_REG_1__SCAN_IN), .ZN(n6653) );
  INV_X1 U5207 ( .A(n6653), .ZN(n4228) );
  NAND2_X1 U5208 ( .A1(n4228), .A2(n6530), .ZN(n6043) );
  NAND2_X1 U5209 ( .A1(n6422), .A2(REIP_REG_0__SCAN_IN), .ZN(n4277) );
  OAI21_X1 U5210 ( .B1(n5133), .B2(n6043), .A(n4277), .ZN(n4236) );
  NAND2_X1 U5211 ( .A1(n6644), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4230) );
  NAND2_X1 U5212 ( .A1(n6999), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4229) );
  AND2_X1 U5213 ( .A1(n4230), .A2(n4229), .ZN(n4299) );
  NAND2_X1 U5214 ( .A1(n6537), .A2(n4231), .ZN(n4232) );
  NAND2_X1 U5215 ( .A1(n4232), .A2(n6644), .ZN(n4233) );
  INV_X1 U5216 ( .A(PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n4234) );
  AOI21_X1 U5217 ( .B1(n4299), .B2(n6047), .A(n4234), .ZN(n4235) );
  AOI211_X1 U5218 ( .C1(n6356), .C2(n4280), .A(n4236), .B(n4235), .ZN(n4237)
         );
  INV_X1 U5219 ( .A(n4237), .ZN(U2986) );
  NAND2_X1 U5220 ( .A1(n4249), .A2(n6662), .ZN(n4238) );
  NOR2_X1 U5221 ( .A1(READY_N), .A2(n5469), .ZN(n4316) );
  NAND2_X1 U5222 ( .A1(n4238), .A2(n4316), .ZN(n4243) );
  NAND2_X1 U5223 ( .A1(n4239), .A2(n6718), .ZN(n4240) );
  INV_X1 U5224 ( .A(n4259), .ZN(n5693) );
  OAI211_X1 U5225 ( .C1(n4352), .C2(n4240), .A(n3348), .B(n5693), .ZN(n4241)
         );
  NAND2_X1 U5226 ( .A1(n5479), .A2(n4241), .ZN(n4242) );
  MUX2_X1 U5227 ( .A(n4243), .B(n4242), .S(n4503), .Z(n4247) );
  NAND2_X1 U5228 ( .A1(n4244), .A2(n3348), .ZN(n4245) );
  MUX2_X1 U5229 ( .A(n6723), .B(n4245), .S(n4324), .Z(n4262) );
  NAND2_X1 U5230 ( .A1(n4250), .A2(n4262), .ZN(n4246) );
  NAND2_X1 U5231 ( .A1(n4246), .A2(n5476), .ZN(n4343) );
  NAND2_X1 U5232 ( .A1(n4269), .A2(n4249), .ZN(n4257) );
  OR2_X1 U5233 ( .A1(n5479), .A2(n4257), .ZN(n4337) );
  NAND3_X1 U5234 ( .A1(n4247), .A2(n4343), .A3(n4337), .ZN(n4248) );
  INV_X1 U5235 ( .A(n6602), .ZN(n4255) );
  NOR2_X1 U5236 ( .A1(n4249), .A2(n3348), .ZN(n5478) );
  AND2_X1 U5237 ( .A1(n4250), .A2(n5478), .ZN(n5470) );
  INV_X1 U5238 ( .A(n5470), .ZN(n4254) );
  NOR2_X1 U5239 ( .A1(n4352), .A2(n4313), .ZN(n4340) );
  NOR2_X1 U5240 ( .A1(n4272), .A2(n4582), .ZN(n4251) );
  NOR2_X1 U5241 ( .A1(n4340), .A2(n4251), .ZN(n4253) );
  NAND4_X1 U5242 ( .A1(n4255), .A2(n4254), .A3(n4253), .A4(n4252), .ZN(n4256)
         );
  AND2_X1 U5243 ( .A1(n4203), .A2(n4503), .ZN(n4341) );
  NOR2_X1 U5244 ( .A1(n4257), .A2(n4341), .ZN(n4258) );
  NAND2_X1 U5245 ( .A1(n4276), .A2(n5473), .ZN(n6426) );
  NOR2_X1 U5246 ( .A1(n4259), .A2(n4503), .ZN(n4260) );
  NOR2_X1 U5247 ( .A1(n4341), .A2(n4260), .ZN(n4261) );
  OAI211_X1 U5248 ( .C1(n4264), .C2(n4263), .A(n4262), .B(n4261), .ZN(n4265)
         );
  NOR2_X1 U5249 ( .A1(n4266), .A2(n4265), .ZN(n4355) );
  NAND2_X1 U5250 ( .A1(n4350), .A2(n4267), .ZN(n4270) );
  NAND2_X1 U5251 ( .A1(n4269), .A2(n4268), .ZN(n4453) );
  NAND3_X1 U5252 ( .A1(n4355), .A2(n4270), .A3(n4453), .ZN(n4271) );
  OR2_X1 U5253 ( .A1(n6399), .A2(n6070), .ZN(n6074) );
  AND2_X1 U5254 ( .A1(n6074), .A2(n5352), .ZN(n4389) );
  OAI21_X1 U5255 ( .B1(n4272), .B2(n3464), .A(n6633), .ZN(n4273) );
  OAI21_X1 U5256 ( .B1(n4275), .B2(INSTADDRPOINTER_REG_0__SCAN_IN), .A(n4274), 
        .ZN(n5124) );
  NOR2_X1 U5257 ( .A1(n4276), .A2(n6422), .ZN(n4526) );
  OAI21_X1 U5258 ( .B1(n4526), .B2(n6073), .A(INSTADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n4278) );
  OAI211_X1 U5259 ( .C1(n6391), .C2(n5124), .A(n4278), .B(n4277), .ZN(n4279)
         );
  AOI211_X1 U5260 ( .C1(n6429), .C2(n4280), .A(n4389), .B(n4279), .ZN(n4281)
         );
  INV_X1 U5261 ( .A(n4281), .ZN(U3018) );
  INV_X1 U5262 ( .A(n4282), .ZN(n4283) );
  OAI21_X1 U5263 ( .B1(n4285), .B2(n4284), .A(n4283), .ZN(n5201) );
  AND2_X1 U5264 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4286) );
  NAND2_X1 U5265 ( .A1(n4287), .A2(n4286), .ZN(n4413) );
  NAND2_X1 U5266 ( .A1(n4287), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4288)
         );
  INV_X1 U5267 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4525) );
  NAND2_X1 U5268 ( .A1(n4288), .A2(n4525), .ZN(n4289) );
  NAND2_X1 U5269 ( .A1(n4481), .A2(n4218), .ZN(n4298) );
  NAND2_X1 U5270 ( .A1(n4291), .A2(n4292), .ZN(n4426) );
  OAI21_X1 U5271 ( .B1(n4292), .B2(n4291), .A(n4426), .ZN(n4293) );
  INV_X1 U5272 ( .A(n4293), .ZN(n4296) );
  NAND3_X1 U5273 ( .A1(n4503), .A2(n3421), .A3(n4294), .ZN(n4295) );
  AOI21_X1 U5274 ( .B1(n4296), .B2(n6240), .A(n4295), .ZN(n4297) );
  NAND2_X1 U5275 ( .A1(n4298), .A2(n4297), .ZN(n4412) );
  XOR2_X1 U5276 ( .A(n4411), .B(n4412), .Z(n4396) );
  NAND2_X1 U5277 ( .A1(n4396), .A2(n6356), .ZN(n4303) );
  INV_X1 U5278 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6710) );
  NOR2_X1 U5279 ( .A1(n6407), .A2(n6710), .ZN(n4390) );
  INV_X1 U5280 ( .A(n4299), .ZN(n4300) );
  NOR2_X1 U5281 ( .A1(n6360), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n4301)
         );
  AOI211_X1 U5282 ( .C1(n6350), .C2(PHYADDRPOINTER_REG_1__SCAN_IN), .A(n4390), 
        .B(n4301), .ZN(n4302) );
  OAI211_X1 U5283 ( .C1(n6043), .C2(n5201), .A(n4303), .B(n4302), .ZN(U2985)
         );
  INV_X1 U5284 ( .A(n5473), .ZN(n4304) );
  OR2_X1 U5285 ( .A1(n5479), .A2(n4304), .ZN(n4309) );
  AND3_X1 U5286 ( .A1(n4305), .A2(n4582), .A3(n5692), .ZN(n4320) );
  NAND4_X1 U5287 ( .A1(n4307), .A2(n4508), .A3(n4320), .A4(n4306), .ZN(n4308)
         );
  NAND2_X1 U5288 ( .A1(n4309), .A2(n4308), .ZN(n4310) );
  AND2_X2 U5289 ( .A1(n4310), .A2(n6641), .ZN(n6023) );
  NAND2_X1 U5290 ( .A1(n6023), .A2(n5696), .ZN(n5691) );
  INV_X1 U5291 ( .A(EBX_REG_1__SCAN_IN), .ZN(n4315) );
  INV_X1 U5292 ( .A(n5194), .ZN(n4314) );
  INV_X1 U5293 ( .A(n4311), .ZN(n4312) );
  AOI21_X1 U5294 ( .B1(n4314), .B2(n4313), .A(n4312), .ZN(n4393) );
  OAI222_X1 U5295 ( .A1(n5201), .A2(n5691), .B1(n6023), .B2(n4315), .C1(n5689), 
        .C2(n4393), .ZN(U2858) );
  NAND2_X1 U5296 ( .A1(n5479), .A2(n5470), .ZN(n4319) );
  INV_X1 U5297 ( .A(n4252), .ZN(n4317) );
  NAND2_X1 U5298 ( .A1(n4317), .A2(n4316), .ZN(n4318) );
  NAND2_X1 U5299 ( .A1(n4319), .A2(n4318), .ZN(n4345) );
  AND2_X1 U5300 ( .A1(n4350), .A2(n4320), .ZN(n4321) );
  OAI21_X1 U5301 ( .B1(n4345), .B2(n4321), .A(n6641), .ZN(n4323) );
  AND2_X1 U5302 ( .A1(n4340), .A2(n6718), .ZN(n4322) );
  NAND2_X1 U5303 ( .A1(n6238), .A2(n4322), .ZN(n6272) );
  NAND2_X1 U5304 ( .A1(n4324), .A2(n5696), .ZN(n4325) );
  INV_X1 U5305 ( .A(n4325), .ZN(n4326) );
  INV_X1 U5306 ( .A(DATAI_1_), .ZN(n7005) );
  INV_X1 U5307 ( .A(EAX_REG_1__SCAN_IN), .ZN(n6280) );
  OAI222_X1 U5308 ( .A1(n5201), .A2(n6024), .B1(n5291), .B2(n7005), .C1(n5698), 
        .C2(n6280), .ZN(U2890) );
  OAI222_X1 U5309 ( .A1(n5133), .A2(n5691), .B1(n5125), .B2(n6023), .C1(n5689), 
        .C2(n5124), .ZN(U2859) );
  INV_X1 U5310 ( .A(EAX_REG_19__SCAN_IN), .ZN(n6248) );
  AOI22_X1 U5311 ( .A1(n4333), .A2(UWORD_REG_3__SCAN_IN), .B1(n6229), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n4327) );
  OAI21_X1 U5312 ( .B1(n6248), .B2(n4336), .A(n4327), .ZN(U2904) );
  INV_X1 U5313 ( .A(EAX_REG_21__SCAN_IN), .ZN(n6252) );
  AOI22_X1 U5314 ( .A1(n4333), .A2(UWORD_REG_5__SCAN_IN), .B1(n6229), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n4328) );
  OAI21_X1 U5315 ( .B1(n6252), .B2(n4336), .A(n4328), .ZN(U2902) );
  INV_X1 U5316 ( .A(EAX_REG_18__SCAN_IN), .ZN(n6246) );
  AOI22_X1 U5317 ( .A1(n4333), .A2(UWORD_REG_2__SCAN_IN), .B1(n6229), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n4329) );
  OAI21_X1 U5318 ( .B1(n6246), .B2(n4336), .A(n4329), .ZN(U2905) );
  AOI22_X1 U5319 ( .A1(n4333), .A2(UWORD_REG_7__SCAN_IN), .B1(n6229), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n4330) );
  OAI21_X1 U5320 ( .B1(n6256), .B2(n4336), .A(n4330), .ZN(U2900) );
  INV_X1 U5321 ( .A(EAX_REG_20__SCAN_IN), .ZN(n6250) );
  AOI22_X1 U5322 ( .A1(n4333), .A2(UWORD_REG_4__SCAN_IN), .B1(n6229), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n4331) );
  OAI21_X1 U5323 ( .B1(n6250), .B2(n4336), .A(n4331), .ZN(U2903) );
  INV_X1 U5324 ( .A(EAX_REG_17__SCAN_IN), .ZN(n6244) );
  AOI22_X1 U5325 ( .A1(n4333), .A2(UWORD_REG_1__SCAN_IN), .B1(n6229), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n4332) );
  OAI21_X1 U5326 ( .B1(n6244), .B2(n4336), .A(n4332), .ZN(U2906) );
  INV_X1 U5327 ( .A(EAX_REG_22__SCAN_IN), .ZN(n6254) );
  AOI22_X1 U5328 ( .A1(n4333), .A2(UWORD_REG_6__SCAN_IN), .B1(n6229), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n4334) );
  OAI21_X1 U5329 ( .B1(n6254), .B2(n4336), .A(n4334), .ZN(U2901) );
  INV_X1 U5330 ( .A(EAX_REG_16__SCAN_IN), .ZN(n6242) );
  AOI22_X1 U5331 ( .A1(n4333), .A2(UWORD_REG_0__SCAN_IN), .B1(n6229), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n4335) );
  OAI21_X1 U5332 ( .B1(n6242), .B2(n4336), .A(n4335), .ZN(U2907) );
  INV_X1 U5333 ( .A(DATAI_0_), .ZN(n7036) );
  INV_X1 U5334 ( .A(EAX_REG_0__SCAN_IN), .ZN(n6277) );
  OAI222_X1 U5335 ( .A1(n5133), .A2(n6024), .B1(n5291), .B2(n7036), .C1(n5698), 
        .C2(n6277), .ZN(U2891) );
  INV_X1 U5336 ( .A(n4337), .ZN(n4347) );
  AOI21_X1 U5337 ( .B1(n4338), .B2(n4352), .A(n6662), .ZN(n4339) );
  OAI211_X1 U5338 ( .C1(n4340), .C2(n4339), .A(n5479), .B(n6718), .ZN(n4344)
         );
  INV_X1 U5339 ( .A(n4341), .ZN(n4342) );
  NAND3_X1 U5340 ( .A1(n4344), .A2(n4343), .A3(n4342), .ZN(n4346) );
  INV_X1 U5341 ( .A(FLUSH_REG_SCAN_IN), .ZN(n7067) );
  NAND2_X1 U5342 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4474), .ZN(n6707) );
  OAI22_X1 U5343 ( .A1(n4467), .A2(n6648), .B1(n7067), .B2(n6707), .ZN(n4383)
         );
  AOI21_X1 U5344 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n6644), .A(n4383), .ZN(
        n5466) );
  INV_X1 U5345 ( .A(n4350), .ZN(n4351) );
  AND2_X1 U5346 ( .A1(n4352), .A2(n4351), .ZN(n4353) );
  AND2_X1 U5347 ( .A1(n4252), .A2(n4353), .ZN(n4354) );
  NAND2_X1 U5348 ( .A1(n4355), .A2(n4354), .ZN(n5350) );
  INV_X1 U5349 ( .A(n5350), .ZN(n4356) );
  OR2_X1 U5350 ( .A1(n4349), .A2(n4356), .ZN(n4362) );
  NOR2_X1 U5351 ( .A1(n4358), .A2(n4357), .ZN(n4363) );
  NOR2_X1 U5352 ( .A1(n5348), .A2(n4363), .ZN(n4359) );
  AOI21_X1 U5353 ( .B1(n5355), .B2(n4360), .A(n4359), .ZN(n4361) );
  NAND2_X1 U5354 ( .A1(n4362), .A2(n4361), .ZN(n6615) );
  INV_X1 U5355 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5857) );
  AOI22_X1 U5356 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n5857), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n4525), .ZN(n5460) );
  INV_X1 U5357 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5352) );
  NOR2_X1 U5358 ( .A1(n6645), .A2(n5352), .ZN(n5458) );
  INV_X1 U5359 ( .A(n4363), .ZN(n4364) );
  AOI222_X1 U5360 ( .A1(n6615), .A2(n5463), .B1(n5460), .B2(n5458), .C1(n4364), 
        .C2(n6637), .ZN(n4366) );
  NAND2_X1 U5361 ( .A1(n5466), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4365) );
  OAI21_X1 U5362 ( .B1(n5466), .B2(n4366), .A(n4365), .ZN(U3460) );
  NAND2_X1 U5363 ( .A1(n6189), .A2(n5350), .ZN(n4379) );
  OR2_X1 U5364 ( .A1(n5473), .A2(n5470), .ZN(n4456) );
  INV_X1 U5365 ( .A(n4368), .ZN(n5457) );
  AOI21_X1 U5366 ( .B1(n5457), .B2(n4369), .A(n4463), .ZN(n4370) );
  NAND3_X1 U5367 ( .A1(n4456), .A2(n4370), .A3(n3652), .ZN(n4377) );
  AND2_X1 U5368 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4373) );
  INV_X1 U5369 ( .A(n4373), .ZN(n4371) );
  XNOR2_X1 U5370 ( .A(n4371), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4375)
         );
  INV_X1 U5371 ( .A(n4453), .ZN(n4374) );
  OAI211_X1 U5372 ( .C1(n4373), .C2(n4447), .A(n3535), .B(n4372), .ZN(n4380)
         );
  AOI22_X1 U5373 ( .A1(n5355), .A2(n4375), .B1(n4374), .B2(n4380), .ZN(n4376)
         );
  AND2_X1 U5374 ( .A1(n4377), .A2(n4376), .ZN(n4378) );
  NAND2_X1 U5375 ( .A1(n4379), .A2(n4378), .ZN(n4446) );
  AOI22_X1 U5376 ( .A1(n4446), .A2(n5463), .B1(n6637), .B2(n4380), .ZN(n4382)
         );
  NAND2_X1 U5377 ( .A1(n5466), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4381) );
  OAI21_X1 U5378 ( .B1(n5466), .B2(n4382), .A(n4381), .ZN(U3456) );
  INV_X1 U5379 ( .A(n5466), .ZN(n5358) );
  NAND2_X1 U5380 ( .A1(n6709), .A2(n4383), .ZN(n4387) );
  INV_X1 U5381 ( .A(n4922), .ZN(n4970) );
  OR2_X1 U5382 ( .A1(n4384), .A2(n4970), .ZN(n4385) );
  XNOR2_X1 U5383 ( .A(n4385), .B(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n5174)
         );
  NOR2_X1 U5384 ( .A1(n4252), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4386) );
  NAND2_X1 U5385 ( .A1(n5174), .A2(n4386), .ZN(n4470) );
  OAI22_X1 U5386 ( .A1(n5358), .A2(n4388), .B1(n4387), .B2(n4470), .ZN(U3455)
         );
  OAI21_X1 U5387 ( .B1(n4526), .B2(n4389), .A(INSTADDRPOINTER_REG_1__SCAN_IN), 
        .ZN(n4392) );
  INV_X1 U5388 ( .A(n4390), .ZN(n4391) );
  OAI211_X1 U5389 ( .C1(n6391), .C2(n4393), .A(n4392), .B(n4391), .ZN(n4395)
         );
  NOR2_X1 U5390 ( .A1(n6073), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4532)
         );
  NOR3_X1 U5391 ( .A1(n5438), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n4532), 
        .ZN(n4394) );
  AOI211_X1 U5392 ( .C1(n4396), .C2(n6429), .A(n4395), .B(n4394), .ZN(n4397)
         );
  INV_X1 U5393 ( .A(n4397), .ZN(U3017) );
  NOR2_X1 U5394 ( .A1(n4399), .A2(n4398), .ZN(n4400) );
  NOR2_X1 U5395 ( .A1(n4480), .A2(n4400), .ZN(n6355) );
  INV_X1 U5396 ( .A(n6355), .ZN(n5142) );
  AND2_X1 U5397 ( .A1(n4402), .A2(n4401), .ZN(n4403) );
  NOR2_X1 U5398 ( .A1(n4553), .A2(n4403), .ZN(n6423) );
  INV_X1 U5399 ( .A(n6023), .ZN(n5668) );
  AOI22_X1 U5400 ( .A1(n6018), .A2(n6423), .B1(EBX_REG_2__SCAN_IN), .B2(n5668), 
        .ZN(n4404) );
  OAI21_X1 U5401 ( .B1(n5142), .B2(n5691), .A(n4404), .ZN(U2857) );
  INV_X1 U5402 ( .A(DATAI_2_), .ZN(n7091) );
  INV_X1 U5403 ( .A(EAX_REG_2__SCAN_IN), .ZN(n6283) );
  OAI222_X1 U5404 ( .A1(n5142), .A2(n6024), .B1(n5291), .B2(n7091), .C1(n5698), 
        .C2(n6283), .ZN(U2889) );
  AOI21_X1 U5405 ( .B1(n4480), .B2(n4479), .A(n4406), .ZN(n4407) );
  NOR2_X1 U5406 ( .A1(n3727), .A2(n4407), .ZN(n4444) );
  INV_X1 U5407 ( .A(n4444), .ZN(n5176) );
  NAND2_X1 U5408 ( .A1(n4554), .A2(n4408), .ZN(n4409) );
  AND2_X1 U5409 ( .A1(n4537), .A2(n4409), .ZN(n6405) );
  AOI22_X1 U5410 ( .A1(n6018), .A2(n6405), .B1(EBX_REG_4__SCAN_IN), .B2(n5668), 
        .ZN(n4410) );
  OAI21_X1 U5411 ( .B1(n5176), .B2(n5691), .A(n4410), .ZN(U2855) );
  NAND2_X1 U5412 ( .A1(n4412), .A2(n4411), .ZN(n4414) );
  NAND2_X1 U5413 ( .A1(n6351), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4419)
         );
  XNOR2_X1 U5414 ( .A(n4426), .B(n4415), .ZN(n4417) );
  OAI21_X1 U5415 ( .B1(n4417), .B2(n6723), .A(n4416), .ZN(n4418) );
  AOI21_X1 U5416 ( .B1(n4483), .B2(n4218), .A(n4418), .ZN(n6352) );
  NAND2_X1 U5417 ( .A1(n4419), .A2(n6352), .ZN(n4423) );
  INV_X1 U5418 ( .A(n6351), .ZN(n4421) );
  INV_X1 U5419 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4420) );
  NAND2_X1 U5420 ( .A1(n4421), .A2(n4420), .ZN(n4422) );
  AND2_X1 U5421 ( .A1(n4423), .A2(n4422), .ZN(n6343) );
  NAND2_X1 U5422 ( .A1(n4424), .A2(n4218), .ZN(n4430) );
  NAND2_X1 U5423 ( .A1(n4426), .A2(n4425), .ZN(n4435) );
  INV_X1 U5424 ( .A(n4434), .ZN(n4427) );
  XNOR2_X1 U5425 ( .A(n4435), .B(n4427), .ZN(n4428) );
  NAND2_X1 U5426 ( .A1(n4428), .A2(n6240), .ZN(n4429) );
  NAND2_X1 U5427 ( .A1(n4430), .A2(n4429), .ZN(n4431) );
  INV_X1 U5428 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6417) );
  XNOR2_X1 U5429 ( .A(n4431), .B(n6417), .ZN(n6344) );
  NAND2_X1 U5430 ( .A1(n6343), .A2(n6344), .ZN(n6342) );
  NAND2_X1 U5431 ( .A1(n4431), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4432)
         );
  NAND2_X1 U5432 ( .A1(n6342), .A2(n4432), .ZN(n4440) );
  NAND2_X1 U5433 ( .A1(n4433), .A2(n4218), .ZN(n4438) );
  NAND2_X1 U5434 ( .A1(n4435), .A2(n4434), .ZN(n4567) );
  XNOR2_X1 U5435 ( .A(n4567), .B(n4565), .ZN(n4436) );
  NAND2_X1 U5436 ( .A1(n4436), .A2(n6240), .ZN(n4437) );
  NAND2_X1 U5437 ( .A1(n4438), .A2(n4437), .ZN(n4514) );
  XNOR2_X1 U5438 ( .A(n4514), .B(n6412), .ZN(n4439) );
  NAND2_X1 U5439 ( .A1(n4440), .A2(n4439), .ZN(n4516) );
  OR2_X1 U5440 ( .A1(n4440), .A2(n4439), .ZN(n4441) );
  NAND2_X1 U5441 ( .A1(n4516), .A2(n4441), .ZN(n6404) );
  INV_X1 U5442 ( .A(n6043), .ZN(n6337) );
  AOI22_X1 U5443 ( .A1(n6350), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .B1(n6422), 
        .B2(REIP_REG_4__SCAN_IN), .ZN(n4442) );
  OAI21_X1 U5444 ( .B1(n5164), .B2(n6360), .A(n4442), .ZN(n4443) );
  AOI21_X1 U5445 ( .B1(n4444), .B2(n6337), .A(n4443), .ZN(n4445) );
  OAI21_X1 U5446 ( .B1(n6096), .B2(n6404), .A(n4445), .ZN(U2982) );
  INV_X1 U5447 ( .A(DATAI_4_), .ZN(n7098) );
  INV_X1 U5448 ( .A(EAX_REG_4__SCAN_IN), .ZN(n6289) );
  OAI222_X1 U5449 ( .A1(n5176), .A2(n6024), .B1(n5291), .B2(n7098), .C1(n5698), 
        .C2(n6289), .ZN(U2887) );
  OR2_X1 U5450 ( .A1(n4446), .A2(n4467), .ZN(n4449) );
  NAND2_X1 U5451 ( .A1(n4467), .A2(n4447), .ZN(n4448) );
  NAND2_X1 U5452 ( .A1(n4449), .A2(n4448), .ZN(n6627) );
  NAND2_X1 U5453 ( .A1(n5134), .A2(n5350), .ZN(n4458) );
  XNOR2_X1 U5454 ( .A(n4368), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4455)
         );
  XNOR2_X1 U5455 ( .A(n5467), .B(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4451)
         );
  NAND2_X1 U5456 ( .A1(n5355), .A2(n4451), .ZN(n4452) );
  OAI21_X1 U5457 ( .B1(n4455), .B2(n4453), .A(n4452), .ZN(n4454) );
  AOI21_X1 U5458 ( .B1(n4456), .B2(n4455), .A(n4454), .ZN(n4457) );
  NAND2_X1 U5459 ( .A1(n4458), .A2(n4457), .ZN(n5464) );
  NAND2_X1 U5460 ( .A1(n5464), .A2(n6614), .ZN(n4460) );
  NAND2_X1 U5461 ( .A1(n4467), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4459) );
  NAND2_X1 U5462 ( .A1(n4460), .A2(n4459), .ZN(n6621) );
  NAND2_X1 U5463 ( .A1(n6621), .A2(n6645), .ZN(n4461) );
  OR2_X1 U5464 ( .A1(n6627), .A2(n4461), .ZN(n4465) );
  NOR2_X1 U5465 ( .A1(FLUSH_REG_SCAN_IN), .A2(n6645), .ZN(n4462) );
  NAND2_X1 U5466 ( .A1(n4463), .A2(n4462), .ZN(n4464) );
  NAND2_X1 U5467 ( .A1(n4465), .A2(n4464), .ZN(n6609) );
  INV_X1 U5468 ( .A(n4466), .ZN(n4471) );
  MUX2_X1 U5469 ( .A(n4467), .B(n7067), .S(STATE2_REG_1__SCAN_IN), .Z(n4468)
         );
  NAND2_X1 U5470 ( .A1(n4468), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4469) );
  NAND2_X1 U5471 ( .A1(n4470), .A2(n4469), .ZN(n6601) );
  AOI21_X1 U5472 ( .B1(n6609), .B2(n4471), .A(n6601), .ZN(n4475) );
  AND2_X1 U5473 ( .A1(n4475), .A2(n7067), .ZN(n4473) );
  OAI21_X1 U5474 ( .B1(n4473), .B2(n6707), .A(n4646), .ZN(n6434) );
  NAND2_X1 U5475 ( .A1(n4475), .A2(n4474), .ZN(n6643) );
  INV_X1 U5476 ( .A(n6643), .ZN(n4477) );
  INV_X1 U5477 ( .A(n5351), .ZN(n6533) );
  AND2_X1 U5478 ( .A1(n6709), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5988) );
  OAI22_X1 U5479 ( .A1(n4920), .A2(n6537), .B1(n6533), .B2(n5988), .ZN(n4476)
         );
  OAI21_X1 U5480 ( .B1(n4477), .B2(n4476), .A(n6434), .ZN(n4478) );
  OAI21_X1 U5481 ( .B1(n6434), .B2(n6610), .A(n4478), .ZN(U3465) );
  XOR2_X1 U5482 ( .A(n4480), .B(n4479), .Z(n6346) );
  INV_X1 U5483 ( .A(n6346), .ZN(n4557) );
  INV_X1 U5484 ( .A(DATAI_3_), .ZN(n6902) );
  INV_X1 U5485 ( .A(EAX_REG_3__SCAN_IN), .ZN(n6286) );
  OAI222_X1 U5486 ( .A1(n4557), .A2(n6024), .B1(n5291), .B2(n6902), .C1(n5698), 
        .C2(n6286), .ZN(U2888) );
  NAND2_X1 U5487 ( .A1(n5978), .A2(n4920), .ZN(n4921) );
  INV_X1 U5488 ( .A(n4482), .ZN(n4919) );
  NOR2_X1 U5489 ( .A1(n4921), .A2(n4919), .ZN(n4484) );
  AND2_X1 U5490 ( .A1(n4484), .A2(n5981), .ZN(n4858) );
  INV_X1 U5491 ( .A(n6043), .ZN(n6354) );
  NAND2_X1 U5492 ( .A1(n6354), .A2(DATAI_31_), .ZN(n6600) );
  INV_X1 U5493 ( .A(n5981), .ZN(n6439) );
  INV_X1 U5494 ( .A(n5978), .ZN(n4485) );
  NOR3_X1 U5495 ( .A1(n6439), .A2(n4919), .A3(n4485), .ZN(n4486) );
  AND2_X1 U5496 ( .A1(n6530), .A2(n6999), .ZN(n5016) );
  INV_X1 U5497 ( .A(n5016), .ZN(n5991) );
  OAI21_X1 U5498 ( .B1(n4486), .B2(n6043), .A(n5991), .ZN(n4489) );
  INV_X1 U5499 ( .A(n4349), .ZN(n5195) );
  AND2_X1 U5500 ( .A1(n5134), .A2(n5195), .ZN(n4727) );
  INV_X1 U5501 ( .A(n4727), .ZN(n4923) );
  NAND2_X1 U5502 ( .A1(n6189), .A2(n5351), .ZN(n4593) );
  OR2_X1 U5503 ( .A1(n4923), .A2(n4593), .ZN(n4487) );
  NAND2_X1 U5504 ( .A1(n4487), .A2(n4911), .ZN(n4493) );
  INV_X1 U5505 ( .A(n4493), .ZN(n4488) );
  NAND2_X1 U5506 ( .A1(n4489), .A2(n4488), .ZN(n4490) );
  AOI21_X1 U5507 ( .B1(n6610), .B2(STATE2_REG_3__SCAN_IN), .A(n4646), .ZN(
        n6481) );
  OAI211_X1 U5508 ( .C1(n4721), .C2(n6530), .A(n4490), .B(n6481), .ZN(n4915)
         );
  NAND2_X1 U5509 ( .A1(n4915), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4497)
         );
  NAND2_X1 U5510 ( .A1(n6354), .A2(DATAI_23_), .ZN(n6591) );
  INV_X1 U5511 ( .A(n6591), .ZN(n6519) );
  NAND2_X1 U5512 ( .A1(n5978), .A2(n4976), .ZN(n5292) );
  NOR2_X1 U5513 ( .A1(n5292), .A2(n4919), .ZN(n4491) );
  NAND3_X1 U5514 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n6644), .A3(n4492), .ZN(
        n4615) );
  NOR2_X1 U5515 ( .A1(n4615), .A2(n5692), .ZN(n6517) );
  INV_X1 U5516 ( .A(n6517), .ZN(n6590) );
  AOI22_X1 U5517 ( .A1(n4493), .A2(n6530), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4721), .ZN(n4912) );
  INV_X1 U5518 ( .A(DATAI_7_), .ZN(n7104) );
  NOR2_X2 U5519 ( .A1(n7104), .A2(n4646), .ZN(n6595) );
  INV_X1 U5520 ( .A(n6595), .ZN(n4494) );
  OAI22_X1 U5521 ( .A1(n6590), .A2(n4911), .B1(n4912), .B2(n4494), .ZN(n4495)
         );
  AOI21_X1 U5522 ( .B1(n6519), .B2(n4914), .A(n4495), .ZN(n4496) );
  OAI211_X1 U5523 ( .C1(n4918), .C2(n6600), .A(n4497), .B(n4496), .ZN(U3147)
         );
  NAND2_X1 U5524 ( .A1(n6354), .A2(DATAI_24_), .ZN(n6528) );
  NAND2_X1 U5525 ( .A1(n4915), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4502)
         );
  NAND2_X1 U5526 ( .A1(n6354), .A2(DATAI_16_), .ZN(n6546) );
  INV_X1 U5527 ( .A(n6546), .ZN(n5328) );
  NOR2_X1 U5528 ( .A1(n4615), .A2(n4498), .ZN(n6477) );
  INV_X1 U5529 ( .A(n6477), .ZN(n6527) );
  NOR2_X2 U5530 ( .A1(n7036), .A2(n4646), .ZN(n6543) );
  INV_X1 U5531 ( .A(n6543), .ZN(n4499) );
  OAI22_X1 U5532 ( .A1(n6527), .A2(n4911), .B1(n4912), .B2(n4499), .ZN(n4500)
         );
  AOI21_X1 U5533 ( .B1(n5328), .B2(n4914), .A(n4500), .ZN(n4501) );
  OAI211_X1 U5534 ( .C1(n4918), .C2(n6528), .A(n4502), .B(n4501), .ZN(U3140)
         );
  NAND2_X1 U5535 ( .A1(n6337), .A2(DATAI_26_), .ZN(n6560) );
  NAND2_X1 U5536 ( .A1(n4915), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4507)
         );
  NAND2_X1 U5537 ( .A1(n6354), .A2(DATAI_18_), .ZN(n6555) );
  INV_X1 U5538 ( .A(n6555), .ZN(n6496) );
  NOR2_X1 U5539 ( .A1(n4615), .A2(n4503), .ZN(n6495) );
  INV_X1 U5540 ( .A(n6495), .ZN(n6554) );
  NOR2_X2 U5541 ( .A1(n7091), .A2(n4646), .ZN(n6557) );
  INV_X1 U5542 ( .A(n6557), .ZN(n4504) );
  OAI22_X1 U5543 ( .A1(n6554), .A2(n4911), .B1(n4912), .B2(n4504), .ZN(n4505)
         );
  AOI21_X1 U5544 ( .B1(n6496), .B2(n4914), .A(n4505), .ZN(n4506) );
  OAI211_X1 U5545 ( .C1(n4918), .C2(n6560), .A(n4507), .B(n4506), .ZN(U3142)
         );
  NAND2_X1 U5546 ( .A1(n6337), .A2(DATAI_27_), .ZN(n6567) );
  NAND2_X1 U5547 ( .A1(n4915), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4512)
         );
  NAND2_X1 U5548 ( .A1(n6337), .A2(DATAI_19_), .ZN(n6562) );
  INV_X1 U5549 ( .A(n6562), .ZN(n6500) );
  NOR2_X1 U5550 ( .A1(n4615), .A2(n4508), .ZN(n6499) );
  INV_X1 U5551 ( .A(n6499), .ZN(n6561) );
  NOR2_X2 U5552 ( .A1(n6902), .A2(n4646), .ZN(n6564) );
  INV_X1 U5553 ( .A(n6564), .ZN(n4509) );
  OAI22_X1 U5554 ( .A1(n6561), .A2(n4911), .B1(n4912), .B2(n4509), .ZN(n4510)
         );
  AOI21_X1 U5555 ( .B1(n6500), .B2(n4914), .A(n4510), .ZN(n4511) );
  OAI211_X1 U5556 ( .C1(n4918), .C2(n6567), .A(n4512), .B(n4511), .ZN(U3143)
         );
  XNOR2_X1 U5557 ( .A(n4405), .B(n4545), .ZN(n6336) );
  INV_X1 U5558 ( .A(n6336), .ZN(n4560) );
  AOI22_X1 U5559 ( .A1(n5720), .A2(DATAI_5_), .B1(n6213), .B2(
        EAX_REG_5__SCAN_IN), .ZN(n4513) );
  OAI21_X1 U5560 ( .B1(n4560), .B2(n6024), .A(n4513), .ZN(U2886) );
  NAND2_X1 U5561 ( .A1(n4514), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4515)
         );
  NAND2_X1 U5562 ( .A1(n4516), .A2(n4515), .ZN(n4523) );
  NAND2_X1 U5563 ( .A1(n4517), .A2(n4218), .ZN(n4522) );
  OR2_X1 U5564 ( .A1(n4567), .A2(n4518), .ZN(n4519) );
  XNOR2_X1 U5565 ( .A(n4519), .B(n4564), .ZN(n4520) );
  NAND2_X1 U5566 ( .A1(n4520), .A2(n6240), .ZN(n4521) );
  NAND2_X1 U5567 ( .A1(n4522), .A2(n4521), .ZN(n4561) );
  INV_X1 U5568 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4531) );
  XNOR2_X1 U5569 ( .A(n4561), .B(n4531), .ZN(n4524) );
  NAND2_X1 U5570 ( .A1(n4523), .A2(n4524), .ZN(n4782) );
  OAI21_X1 U5571 ( .B1(n4523), .B2(n4524), .A(n4562), .ZN(n6335) );
  NAND2_X1 U5572 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4535) );
  INV_X1 U5573 ( .A(n4535), .ZN(n6402) );
  AOI21_X1 U5574 ( .B1(INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .A(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n6420) );
  INV_X1 U5575 ( .A(n6420), .ZN(n6401) );
  NAND2_X1 U5576 ( .A1(n6402), .A2(n6401), .ZN(n4530) );
  NOR2_X1 U5577 ( .A1(n4531), .A2(n4530), .ZN(n5096) );
  INV_X1 U5578 ( .A(n4534), .ZN(n5423) );
  NOR2_X1 U5579 ( .A1(n4420), .A2(n4525), .ZN(n6421) );
  INV_X1 U5580 ( .A(n4526), .ZN(n4528) );
  NAND2_X1 U5581 ( .A1(n6070), .A2(n5352), .ZN(n4527) );
  OAI21_X1 U5582 ( .B1(n5423), .B2(n6421), .A(n5373), .ZN(n6398) );
  INV_X1 U5583 ( .A(n6398), .ZN(n6432) );
  OAI21_X1 U5584 ( .B1(n5438), .B2(n5096), .A(n6432), .ZN(n4529) );
  INV_X1 U5585 ( .A(n4529), .ZN(n6395) );
  AOI221_X1 U5586 ( .B1(n6426), .B2(n4531), .C1(n4530), .C2(n4531), .A(n6395), 
        .ZN(n4542) );
  INV_X1 U5587 ( .A(n4532), .ZN(n4533) );
  NAND3_X1 U5588 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n6419), .ZN(n5095) );
  NOR3_X1 U5589 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n4535), .A3(n5095), 
        .ZN(n4541) );
  AOI21_X1 U5590 ( .B1(n4537), .B2(n4536), .A(n4549), .ZN(n4538) );
  INV_X1 U5591 ( .A(n4538), .ZN(n6175) );
  INV_X1 U5592 ( .A(REIP_REG_5__SCAN_IN), .ZN(n4539) );
  OAI22_X1 U5593 ( .A1(n6391), .A2(n6175), .B1(n6407), .B2(n4539), .ZN(n4540)
         );
  NOR3_X1 U5594 ( .A1(n4542), .A2(n4541), .A3(n4540), .ZN(n4543) );
  OAI21_X1 U5595 ( .B1(n6403), .B2(n6335), .A(n4543), .ZN(U3013) );
  AOI21_X1 U5596 ( .B1(n3727), .B2(n4545), .A(n4544), .ZN(n4547) );
  INV_X1 U5597 ( .A(n4706), .ZN(n4546) );
  NOR2_X1 U5598 ( .A1(n4547), .A2(n4546), .ZN(n4576) );
  INV_X1 U5599 ( .A(n5691), .ZN(n6020) );
  OAI21_X1 U5600 ( .B1(n4549), .B2(n4548), .A(n4768), .ZN(n6392) );
  OAI22_X1 U5601 ( .A1(n5689), .A2(n6392), .B1(n4550), .B2(n6023), .ZN(n4551)
         );
  AOI21_X1 U5602 ( .B1(n4576), .B2(n6020), .A(n4551), .ZN(n4552) );
  INV_X1 U5603 ( .A(n4552), .ZN(U2853) );
  INV_X1 U5604 ( .A(n4553), .ZN(n4555) );
  AOI21_X1 U5605 ( .B1(n4556), .B2(n4555), .A(n3243), .ZN(n6413) );
  INV_X1 U5606 ( .A(n6413), .ZN(n6197) );
  INV_X1 U5607 ( .A(EBX_REG_3__SCAN_IN), .ZN(n4558) );
  OAI222_X1 U5608 ( .A1(n6197), .A2(n5689), .B1(n4558), .B2(n6023), .C1(n4557), 
        .C2(n5688), .ZN(U2856) );
  INV_X1 U5609 ( .A(n4576), .ZN(n5270) );
  INV_X1 U5610 ( .A(DATAI_6_), .ZN(n6989) );
  INV_X1 U5611 ( .A(EAX_REG_6__SCAN_IN), .ZN(n6295) );
  OAI222_X1 U5612 ( .A1(n5270), .A2(n6024), .B1(n5291), .B2(n6989), .C1(n5698), 
        .C2(n6295), .ZN(U2885) );
  INV_X1 U5613 ( .A(EBX_REG_5__SCAN_IN), .ZN(n4559) );
  OAI222_X1 U5614 ( .A1(n6175), .A2(n5689), .B1(n5688), .B2(n4560), .C1(n4559), 
        .C2(n6023), .ZN(U2854) );
  NAND2_X1 U5615 ( .A1(n4561), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4780)
         );
  NAND2_X1 U5616 ( .A1(n4562), .A2(n4780), .ZN(n4572) );
  NAND3_X1 U5617 ( .A1(n4796), .A2(n4218), .A3(n4563), .ZN(n4570) );
  NAND2_X1 U5618 ( .A1(n4565), .A2(n4564), .ZN(n4566) );
  OR2_X1 U5619 ( .A1(n4567), .A2(n4566), .ZN(n4784) );
  XNOR2_X1 U5620 ( .A(n4784), .B(n4785), .ZN(n4568) );
  NAND2_X1 U5621 ( .A1(n4568), .A2(n6240), .ZN(n4569) );
  NAND2_X1 U5622 ( .A1(n4570), .A2(n4569), .ZN(n4779) );
  XNOR2_X1 U5623 ( .A(n4779), .B(n6396), .ZN(n4790) );
  NAND2_X1 U5624 ( .A1(n4572), .A2(n4790), .ZN(n4571) );
  OAI21_X1 U5625 ( .B1(n4572), .B2(n4790), .A(n4571), .ZN(n6390) );
  INV_X1 U5626 ( .A(n4573), .ZN(n5261) );
  AOI22_X1 U5627 ( .A1(n6350), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .B1(n6422), 
        .B2(REIP_REG_6__SCAN_IN), .ZN(n4574) );
  OAI21_X1 U5628 ( .B1(n5261), .B2(n6360), .A(n4574), .ZN(n4575) );
  AOI21_X1 U5629 ( .B1(n4576), .B2(n6337), .A(n4575), .ZN(n4577) );
  OAI21_X1 U5630 ( .B1(n6390), .B2(n6096), .A(n4577), .ZN(U2980) );
  NAND2_X1 U5631 ( .A1(n6337), .A2(DATAI_30_), .ZN(n6588) );
  NAND2_X1 U5632 ( .A1(n4915), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4581)
         );
  NAND2_X1 U5633 ( .A1(n6337), .A2(DATAI_22_), .ZN(n6583) );
  INV_X1 U5634 ( .A(n6583), .ZN(n5318) );
  NOR2_X1 U5635 ( .A1(n4615), .A2(n3428), .ZN(n6511) );
  INV_X1 U5636 ( .A(n6511), .ZN(n6582) );
  NOR2_X2 U5637 ( .A1(n6989), .A2(n4646), .ZN(n6585) );
  INV_X1 U5638 ( .A(n6585), .ZN(n4578) );
  OAI22_X1 U5639 ( .A1(n6582), .A2(n4911), .B1(n4912), .B2(n4578), .ZN(n4579)
         );
  AOI21_X1 U5640 ( .B1(n5318), .B2(n4914), .A(n4579), .ZN(n4580) );
  OAI211_X1 U5641 ( .C1(n4918), .C2(n6588), .A(n4581), .B(n4580), .ZN(U3146)
         );
  AND2_X1 U5642 ( .A1(n6354), .A2(DATAI_28_), .ZN(n6504) );
  INV_X1 U5643 ( .A(n6504), .ZN(n6569) );
  NAND2_X1 U5644 ( .A1(n4915), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4586)
         );
  NAND2_X1 U5645 ( .A1(n6337), .A2(DATAI_20_), .ZN(n6574) );
  INV_X1 U5646 ( .A(n6574), .ZN(n5314) );
  NOR2_X1 U5647 ( .A1(n4615), .A2(n4582), .ZN(n6503) );
  INV_X1 U5648 ( .A(n6503), .ZN(n6568) );
  NOR2_X2 U5649 ( .A1(n7098), .A2(n4646), .ZN(n6571) );
  INV_X1 U5650 ( .A(n6571), .ZN(n4583) );
  OAI22_X1 U5651 ( .A1(n6568), .A2(n4911), .B1(n4912), .B2(n4583), .ZN(n4584)
         );
  AOI21_X1 U5652 ( .B1(n5314), .B2(n4914), .A(n4584), .ZN(n4585) );
  OAI211_X1 U5653 ( .C1(n4918), .C2(n6569), .A(n4586), .B(n4585), .ZN(U3144)
         );
  NAND2_X1 U5654 ( .A1(n6337), .A2(DATAI_25_), .ZN(n6548) );
  NAND2_X1 U5655 ( .A1(n4915), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4590)
         );
  NAND2_X1 U5656 ( .A1(n6337), .A2(DATAI_17_), .ZN(n6553) );
  INV_X1 U5657 ( .A(n6553), .ZN(n6492) );
  NOR2_X1 U5658 ( .A1(n4615), .A2(n3451), .ZN(n6491) );
  INV_X1 U5659 ( .A(n6491), .ZN(n6547) );
  NOR2_X2 U5660 ( .A1(n7005), .A2(n4646), .ZN(n6550) );
  INV_X1 U5661 ( .A(n6550), .ZN(n4587) );
  OAI22_X1 U5662 ( .A1(n6547), .A2(n4911), .B1(n4912), .B2(n4587), .ZN(n4588)
         );
  AOI21_X1 U5663 ( .B1(n6492), .B2(n4914), .A(n4588), .ZN(n4589) );
  OAI211_X1 U5664 ( .C1(n4918), .C2(n6548), .A(n4590), .B(n4589), .ZN(U3141)
         );
  NOR2_X1 U5665 ( .A1(n5978), .A2(n4919), .ZN(n4591) );
  INV_X1 U5666 ( .A(n4598), .ZN(n4592) );
  NAND2_X1 U5667 ( .A1(n4681), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4969) );
  NOR2_X1 U5668 ( .A1(n4929), .A2(n4969), .ZN(n5297) );
  INV_X1 U5669 ( .A(n4593), .ZN(n4683) );
  AND2_X1 U5670 ( .A1(n5134), .A2(n4349), .ZN(n5293) );
  AND2_X1 U5671 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5297), .ZN(n4616)
         );
  AOI21_X1 U5672 ( .B1(n4683), .B2(n5293), .A(n4616), .ZN(n4597) );
  NAND2_X1 U5673 ( .A1(n4598), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5985) );
  NAND3_X1 U5674 ( .A1(n6530), .A2(n4597), .A3(n5985), .ZN(n4594) );
  OAI211_X1 U5675 ( .C1(n6530), .C2(n5297), .A(n6481), .B(n4594), .ZN(n4614)
         );
  NAND2_X1 U5676 ( .A1(n6530), .A2(n5985), .ZN(n4596) );
  NAND2_X1 U5677 ( .A1(STATE2_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4595) );
  OAI22_X1 U5678 ( .A1(n4597), .A2(n4596), .B1(n4969), .B2(n4595), .ZN(n4613)
         );
  AOI22_X1 U5679 ( .A1(INSTQUEUE_REG_13__3__SCAN_IN), .A2(n4614), .B1(n6564), 
        .B2(n4613), .ZN(n4600) );
  INV_X1 U5680 ( .A(n6567), .ZN(n5223) );
  AOI22_X1 U5681 ( .A1(n5338), .A2(n5223), .B1(n6499), .B2(n4616), .ZN(n4599)
         );
  OAI211_X1 U5682 ( .C1(n6562), .C2(n4861), .A(n4600), .B(n4599), .ZN(U3127)
         );
  AOI22_X1 U5683 ( .A1(INSTQUEUE_REG_13__6__SCAN_IN), .A2(n4614), .B1(n6585), 
        .B2(n4613), .ZN(n4602) );
  INV_X1 U5684 ( .A(n6588), .ZN(n6512) );
  AOI22_X1 U5685 ( .A1(n5338), .A2(n6512), .B1(n6511), .B2(n4616), .ZN(n4601)
         );
  OAI211_X1 U5686 ( .C1(n6583), .C2(n4861), .A(n4602), .B(n4601), .ZN(U3130)
         );
  AOI22_X1 U5687 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n4614), .B1(n6571), 
        .B2(n4613), .ZN(n4604) );
  AOI22_X1 U5688 ( .A1(n5338), .A2(n6504), .B1(n6503), .B2(n4616), .ZN(n4603)
         );
  OAI211_X1 U5689 ( .C1(n6574), .C2(n4861), .A(n4604), .B(n4603), .ZN(U3128)
         );
  AOI22_X1 U5690 ( .A1(INSTQUEUE_REG_13__2__SCAN_IN), .A2(n4614), .B1(n6557), 
        .B2(n4613), .ZN(n4606) );
  INV_X1 U5691 ( .A(n6560), .ZN(n5234) );
  AOI22_X1 U5692 ( .A1(n5338), .A2(n5234), .B1(n6495), .B2(n4616), .ZN(n4605)
         );
  OAI211_X1 U5693 ( .C1(n6555), .C2(n4861), .A(n4606), .B(n4605), .ZN(U3126)
         );
  AOI22_X1 U5694 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n4614), .B1(n6543), 
        .B2(n4613), .ZN(n4608) );
  INV_X1 U5695 ( .A(n6528), .ZN(n6478) );
  AOI22_X1 U5696 ( .A1(n5338), .A2(n6478), .B1(n6477), .B2(n4616), .ZN(n4607)
         );
  OAI211_X1 U5697 ( .C1(n6546), .C2(n4861), .A(n4608), .B(n4607), .ZN(U3124)
         );
  AOI22_X1 U5698 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n4614), .B1(n6595), 
        .B2(n4613), .ZN(n4610) );
  INV_X1 U5699 ( .A(n6600), .ZN(n5230) );
  AOI22_X1 U5700 ( .A1(n5338), .A2(n5230), .B1(n6517), .B2(n4616), .ZN(n4609)
         );
  OAI211_X1 U5701 ( .C1(n6591), .C2(n4861), .A(n4610), .B(n4609), .ZN(U3131)
         );
  AOI22_X1 U5702 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n4614), .B1(n6550), 
        .B2(n4613), .ZN(n4612) );
  INV_X1 U5703 ( .A(n6548), .ZN(n5250) );
  AOI22_X1 U5704 ( .A1(n5338), .A2(n5250), .B1(n6491), .B2(n4616), .ZN(n4611)
         );
  OAI211_X1 U5705 ( .C1(n6553), .C2(n4861), .A(n4612), .B(n4611), .ZN(U3125)
         );
  NAND2_X1 U5706 ( .A1(n6337), .A2(DATAI_21_), .ZN(n6581) );
  INV_X1 U5707 ( .A(DATAI_5_), .ZN(n7086) );
  NOR2_X2 U5708 ( .A1(n7086), .A2(n4646), .ZN(n6578) );
  AOI22_X1 U5709 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(n4614), .B1(n6578), 
        .B2(n4613), .ZN(n4618) );
  NAND2_X1 U5710 ( .A1(n6337), .A2(DATAI_29_), .ZN(n6576) );
  INV_X1 U5711 ( .A(n6576), .ZN(n5218) );
  NOR2_X2 U5712 ( .A1(n4615), .A2(n3470), .ZN(n6507) );
  AOI22_X1 U5713 ( .A1(n5338), .A2(n5218), .B1(n6507), .B2(n4616), .ZN(n4617)
         );
  OAI211_X1 U5714 ( .C1(n6581), .C2(n4861), .A(n4618), .B(n4617), .ZN(U3129)
         );
  NAND2_X1 U5715 ( .A1(n4624), .A2(n4920), .ZN(n4850) );
  INV_X1 U5716 ( .A(n5134), .ZN(n5982) );
  NAND2_X1 U5717 ( .A1(n5982), .A2(n4349), .ZN(n5015) );
  OR2_X1 U5718 ( .A1(n5015), .A2(n6189), .ZN(n4816) );
  INV_X1 U5719 ( .A(n4816), .ZN(n4619) );
  NAND3_X1 U5720 ( .A1(n4929), .A2(n6620), .A3(n4681), .ZN(n4811) );
  NOR2_X1 U5721 ( .A1(n6610), .A2(n4811), .ZN(n4641) );
  AOI21_X1 U5722 ( .B1(n4619), .B2(n5351), .A(n4641), .ZN(n4622) );
  AOI21_X1 U5723 ( .B1(n4624), .B2(STATEBS16_REG_SCAN_IN), .A(n6537), .ZN(
        n4621) );
  AOI22_X1 U5724 ( .A1(n4622), .A2(n4621), .B1(n6537), .B2(n4811), .ZN(n4620)
         );
  NAND2_X1 U5725 ( .A1(n6481), .A2(n4620), .ZN(n4640) );
  INV_X1 U5726 ( .A(n4621), .ZN(n4623) );
  OAI22_X1 U5727 ( .A1(n4623), .A2(n4622), .B1(n6636), .B2(n4811), .ZN(n4639)
         );
  AOI22_X1 U5728 ( .A1(INSTQUEUE_REG_1__6__SCAN_IN), .A2(n4640), .B1(n6585), 
        .B2(n4639), .ZN(n4626) );
  AOI22_X1 U5729 ( .A1(n4759), .A2(n5318), .B1(n6511), .B2(n4641), .ZN(n4625)
         );
  OAI211_X1 U5730 ( .C1(n6588), .C2(n4850), .A(n4626), .B(n4625), .ZN(U3034)
         );
  AOI22_X1 U5731 ( .A1(INSTQUEUE_REG_1__1__SCAN_IN), .A2(n4640), .B1(n6550), 
        .B2(n4639), .ZN(n4628) );
  AOI22_X1 U5732 ( .A1(n4759), .A2(n6492), .B1(n6491), .B2(n4641), .ZN(n4627)
         );
  OAI211_X1 U5733 ( .C1(n6548), .C2(n4850), .A(n4628), .B(n4627), .ZN(U3029)
         );
  AOI22_X1 U5734 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(n4640), .B1(n6578), 
        .B2(n4639), .ZN(n4630) );
  INV_X1 U5735 ( .A(n6581), .ZN(n6508) );
  AOI22_X1 U5736 ( .A1(n4759), .A2(n6508), .B1(n6507), .B2(n4641), .ZN(n4629)
         );
  OAI211_X1 U5737 ( .C1(n6576), .C2(n4850), .A(n4630), .B(n4629), .ZN(U3033)
         );
  AOI22_X1 U5738 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n4640), .B1(n6571), 
        .B2(n4639), .ZN(n4632) );
  AOI22_X1 U5739 ( .A1(n4759), .A2(n5314), .B1(n6503), .B2(n4641), .ZN(n4631)
         );
  OAI211_X1 U5740 ( .C1(n6569), .C2(n4850), .A(n4632), .B(n4631), .ZN(U3032)
         );
  AOI22_X1 U5741 ( .A1(INSTQUEUE_REG_1__2__SCAN_IN), .A2(n4640), .B1(n6557), 
        .B2(n4639), .ZN(n4634) );
  AOI22_X1 U5742 ( .A1(n4759), .A2(n6496), .B1(n6495), .B2(n4641), .ZN(n4633)
         );
  OAI211_X1 U5743 ( .C1(n6560), .C2(n4850), .A(n4634), .B(n4633), .ZN(U3030)
         );
  AOI22_X1 U5744 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(n4640), .B1(n6595), 
        .B2(n4639), .ZN(n4636) );
  AOI22_X1 U5745 ( .A1(n4759), .A2(n6519), .B1(n6517), .B2(n4641), .ZN(n4635)
         );
  OAI211_X1 U5746 ( .C1(n6600), .C2(n4850), .A(n4636), .B(n4635), .ZN(U3035)
         );
  AOI22_X1 U5747 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n4640), .B1(n6543), 
        .B2(n4639), .ZN(n4638) );
  AOI22_X1 U5748 ( .A1(n4759), .A2(n5328), .B1(n6477), .B2(n4641), .ZN(n4637)
         );
  OAI211_X1 U5749 ( .C1(n6528), .C2(n4850), .A(n4638), .B(n4637), .ZN(U3028)
         );
  AOI22_X1 U5750 ( .A1(INSTQUEUE_REG_1__3__SCAN_IN), .A2(n4640), .B1(n6564), 
        .B2(n4639), .ZN(n4643) );
  AOI22_X1 U5751 ( .A1(n4759), .A2(n6500), .B1(n6499), .B2(n4641), .ZN(n4642)
         );
  OAI211_X1 U5752 ( .C1(n6567), .C2(n4850), .A(n4643), .B(n4642), .ZN(U3031)
         );
  NAND3_X1 U5753 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n4929), .A3(n6620), .ZN(n6446) );
  NOR2_X1 U5754 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6446), .ZN(n4760)
         );
  INV_X1 U5755 ( .A(n6470), .ZN(n4644) );
  NOR2_X1 U5756 ( .A1(n4759), .A2(n4644), .ZN(n4645) );
  INV_X1 U5757 ( .A(n6189), .ZN(n5987) );
  NOR2_X1 U5758 ( .A1(n5134), .A2(n4349), .ZN(n4867) );
  NAND2_X1 U5759 ( .A1(n5987), .A2(n4867), .ZN(n6442) );
  OAI21_X1 U5760 ( .B1(n4645), .B2(n5016), .A(n6442), .ZN(n4647) );
  AND2_X1 U5761 ( .A1(n4648), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5296) );
  OAI21_X1 U5762 ( .B1(n5019), .B2(n6636), .A(n5022), .ZN(n4724) );
  NOR2_X1 U5763 ( .A1(n5296), .A2(n4724), .ZN(n4870) );
  OAI221_X1 U5764 ( .B1(n4760), .B2(n6709), .C1(n4760), .C2(n4647), .A(n4870), 
        .ZN(n4765) );
  INV_X1 U5765 ( .A(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4654) );
  OR2_X1 U5766 ( .A1(n6442), .A2(n6537), .ZN(n4650) );
  NOR2_X1 U5767 ( .A1(n4648), .A2(n6636), .ZN(n5303) );
  NAND2_X1 U5768 ( .A1(n5303), .A2(n5019), .ZN(n4872) );
  OR2_X1 U5769 ( .A1(n4872), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4649)
         );
  NAND2_X1 U5770 ( .A1(n4650), .A2(n4649), .ZN(n4761) );
  AOI22_X1 U5771 ( .A1(n6499), .A2(n4760), .B1(n6564), .B2(n4761), .ZN(n4651)
         );
  OAI21_X1 U5772 ( .B1(n6470), .B2(n6562), .A(n4651), .ZN(n4652) );
  AOI21_X1 U5773 ( .B1(n4759), .B2(n5223), .A(n4652), .ZN(n4653) );
  OAI21_X1 U5774 ( .B1(n4679), .B2(n4654), .A(n4653), .ZN(U3039) );
  INV_X1 U5775 ( .A(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4658) );
  AOI22_X1 U5776 ( .A1(n6511), .A2(n4760), .B1(n6585), .B2(n4761), .ZN(n4655)
         );
  OAI21_X1 U5777 ( .B1(n6470), .B2(n6583), .A(n4655), .ZN(n4656) );
  AOI21_X1 U5778 ( .B1(n4759), .B2(n6512), .A(n4656), .ZN(n4657) );
  OAI21_X1 U5779 ( .B1(n4679), .B2(n4658), .A(n4657), .ZN(U3042) );
  INV_X1 U5780 ( .A(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4662) );
  AOI22_X1 U5781 ( .A1(n6477), .A2(n4760), .B1(n6543), .B2(n4761), .ZN(n4659)
         );
  OAI21_X1 U5782 ( .B1(n6470), .B2(n6546), .A(n4659), .ZN(n4660) );
  AOI21_X1 U5783 ( .B1(n4759), .B2(n6478), .A(n4660), .ZN(n4661) );
  OAI21_X1 U5784 ( .B1(n4679), .B2(n4662), .A(n4661), .ZN(U3036) );
  INV_X1 U5785 ( .A(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4666) );
  AOI22_X1 U5786 ( .A1(n6503), .A2(n4760), .B1(n6571), .B2(n4761), .ZN(n4663)
         );
  OAI21_X1 U5787 ( .B1(n6470), .B2(n6574), .A(n4663), .ZN(n4664) );
  AOI21_X1 U5788 ( .B1(n4759), .B2(n6504), .A(n4664), .ZN(n4665) );
  OAI21_X1 U5789 ( .B1(n4679), .B2(n4666), .A(n4665), .ZN(U3040) );
  INV_X1 U5790 ( .A(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4670) );
  AOI22_X1 U5791 ( .A1(n6495), .A2(n4760), .B1(n6557), .B2(n4761), .ZN(n4667)
         );
  OAI21_X1 U5792 ( .B1(n6470), .B2(n6555), .A(n4667), .ZN(n4668) );
  AOI21_X1 U5793 ( .B1(n4759), .B2(n5234), .A(n4668), .ZN(n4669) );
  OAI21_X1 U5794 ( .B1(n4679), .B2(n4670), .A(n4669), .ZN(U3038) );
  INV_X1 U5795 ( .A(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4674) );
  AOI22_X1 U5796 ( .A1(n6517), .A2(n4760), .B1(n6595), .B2(n4761), .ZN(n4671)
         );
  OAI21_X1 U5797 ( .B1(n6470), .B2(n6591), .A(n4671), .ZN(n4672) );
  AOI21_X1 U5798 ( .B1(n4759), .B2(n5230), .A(n4672), .ZN(n4673) );
  OAI21_X1 U5799 ( .B1(n4679), .B2(n4674), .A(n4673), .ZN(U3043) );
  INV_X1 U5800 ( .A(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4678) );
  AOI22_X1 U5801 ( .A1(n6491), .A2(n4760), .B1(n6550), .B2(n4761), .ZN(n4675)
         );
  OAI21_X1 U5802 ( .B1(n6470), .B2(n6553), .A(n4675), .ZN(n4676) );
  AOI21_X1 U5803 ( .B1(n4759), .B2(n5250), .A(n4676), .ZN(n4677) );
  OAI21_X1 U5804 ( .B1(n4679), .B2(n4678), .A(n4677), .ZN(U3037) );
  OR3_X1 U5805 ( .A1(n6532), .A2(n5978), .A3(n6999), .ZN(n4680) );
  INV_X1 U5806 ( .A(n5015), .ZN(n4682) );
  NAND3_X1 U5807 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6620), .A3(n4681), .ZN(n5018) );
  NOR2_X1 U5808 ( .A1(n6610), .A2(n5018), .ZN(n4688) );
  AOI21_X1 U5809 ( .B1(n4683), .B2(n4682), .A(n4688), .ZN(n4687) );
  AOI22_X1 U5810 ( .A1(n4685), .A2(n4687), .B1(n6537), .B2(n5018), .ZN(n4684)
         );
  NAND2_X1 U5811 ( .A1(n6481), .A2(n4684), .ZN(n4774) );
  INV_X1 U5812 ( .A(n4685), .ZN(n4686) );
  OAI22_X1 U5813 ( .A1(n4687), .A2(n4686), .B1(n6636), .B2(n5018), .ZN(n4773)
         );
  AOI22_X1 U5814 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n4774), .B1(n6595), 
        .B2(n4773), .ZN(n4691) );
  INV_X1 U5815 ( .A(n4688), .ZN(n4775) );
  OAI22_X1 U5816 ( .A1(n4874), .A2(n6591), .B1(n6590), .B2(n4775), .ZN(n4689)
         );
  AOI21_X1 U5817 ( .B1(n5230), .B2(n5032), .A(n4689), .ZN(n4690) );
  NAND2_X1 U5818 ( .A1(n4691), .A2(n4690), .ZN(U3099) );
  AOI22_X1 U5819 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n4774), .B1(n6585), 
        .B2(n4773), .ZN(n4694) );
  OAI22_X1 U5820 ( .A1(n4874), .A2(n6583), .B1(n6582), .B2(n4775), .ZN(n4692)
         );
  AOI21_X1 U5821 ( .B1(n6512), .B2(n5032), .A(n4692), .ZN(n4693) );
  NAND2_X1 U5822 ( .A1(n4694), .A2(n4693), .ZN(U3098) );
  AOI22_X1 U5823 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4774), .B1(n6571), 
        .B2(n4773), .ZN(n4697) );
  OAI22_X1 U5824 ( .A1(n4874), .A2(n6574), .B1(n6568), .B2(n4775), .ZN(n4695)
         );
  AOI21_X1 U5825 ( .B1(n6504), .B2(n5032), .A(n4695), .ZN(n4696) );
  NAND2_X1 U5826 ( .A1(n4697), .A2(n4696), .ZN(U3096) );
  INV_X1 U5827 ( .A(n4698), .ZN(n4701) );
  INV_X1 U5828 ( .A(n4705), .ZN(n4700) );
  AOI21_X1 U5829 ( .B1(n4701), .B2(n4700), .A(n3176), .ZN(n4808) );
  INV_X1 U5830 ( .A(n4808), .ZN(n5112) );
  INV_X1 U5831 ( .A(n5069), .ZN(n4702) );
  AOI21_X1 U5832 ( .B1(n4703), .B2(n4770), .A(n4702), .ZN(n6377) );
  AOI22_X1 U5833 ( .A1(n6377), .A2(n6018), .B1(EBX_REG_8__SCAN_IN), .B2(n5668), 
        .ZN(n4704) );
  OAI21_X1 U5834 ( .B1(n5112), .B2(n5691), .A(n4704), .ZN(U2851) );
  AOI21_X1 U5835 ( .B1(n4707), .B2(n4706), .A(n4705), .ZN(n6331) );
  INV_X1 U5836 ( .A(n6331), .ZN(n4771) );
  OAI222_X1 U5837 ( .A1(n4771), .A2(n6024), .B1(n5291), .B2(n7104), .C1(n5698), 
        .C2(n3739), .ZN(U2884) );
  AOI22_X1 U5838 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n4774), .B1(n6557), 
        .B2(n4773), .ZN(n4710) );
  OAI22_X1 U5839 ( .A1(n4874), .A2(n6555), .B1(n6554), .B2(n4775), .ZN(n4708)
         );
  INV_X1 U5840 ( .A(n4708), .ZN(n4709) );
  OAI211_X1 U5841 ( .C1(n6560), .C2(n5060), .A(n4710), .B(n4709), .ZN(U3094)
         );
  AOI22_X1 U5842 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n4774), .B1(n6550), 
        .B2(n4773), .ZN(n4713) );
  OAI22_X1 U5843 ( .A1(n4874), .A2(n6553), .B1(n6547), .B2(n4775), .ZN(n4711)
         );
  INV_X1 U5844 ( .A(n4711), .ZN(n4712) );
  OAI211_X1 U5845 ( .C1(n6548), .C2(n5060), .A(n4713), .B(n4712), .ZN(U3093)
         );
  AOI22_X1 U5846 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n4774), .B1(n6564), 
        .B2(n4773), .ZN(n4716) );
  OAI22_X1 U5847 ( .A1(n4874), .A2(n6562), .B1(n6561), .B2(n4775), .ZN(n4714)
         );
  INV_X1 U5848 ( .A(n4714), .ZN(n4715) );
  OAI211_X1 U5849 ( .C1(n6567), .C2(n5060), .A(n4716), .B(n4715), .ZN(U3095)
         );
  AOI22_X1 U5850 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n4774), .B1(n6543), 
        .B2(n4773), .ZN(n4719) );
  OAI22_X1 U5851 ( .A1(n4874), .A2(n6546), .B1(n6527), .B2(n4775), .ZN(n4717)
         );
  INV_X1 U5852 ( .A(n4717), .ZN(n4718) );
  OAI211_X1 U5853 ( .C1(n6528), .C2(n5060), .A(n4719), .B(n4718), .ZN(U3092)
         );
  INV_X1 U5854 ( .A(DATAI_8_), .ZN(n7008) );
  INV_X1 U5855 ( .A(EAX_REG_8__SCAN_IN), .ZN(n6300) );
  OAI222_X1 U5856 ( .A1(n5112), .A2(n6024), .B1(n5291), .B2(n7008), .C1(n5698), 
        .C2(n6300), .ZN(U2883) );
  OAI21_X1 U5857 ( .B1(n4756), .B2(n4858), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n4720) );
  NAND3_X1 U5858 ( .A1(n4923), .A2(n6530), .A3(n4720), .ZN(n4726) );
  INV_X1 U5859 ( .A(n4721), .ZN(n4722) );
  NOR2_X1 U5860 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4722), .ZN(n4857)
         );
  OAI21_X1 U5861 ( .B1(n6709), .B2(n4857), .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), 
        .ZN(n4723) );
  INV_X1 U5862 ( .A(n4723), .ZN(n4725) );
  NOR2_X1 U5863 ( .A1(n5303), .A2(n4724), .ZN(n4927) );
  INV_X1 U5864 ( .A(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4733) );
  AND2_X1 U5865 ( .A1(n4727), .A2(n6530), .ZN(n4930) );
  NAND2_X1 U5866 ( .A1(n4930), .A2(n6189), .ZN(n4729) );
  AND2_X1 U5867 ( .A1(n5296), .A2(n5019), .ZN(n4931) );
  NAND2_X1 U5868 ( .A1(n4931), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4728) );
  NAND2_X1 U5869 ( .A1(n4729), .A2(n4728), .ZN(n4856) );
  AOI22_X1 U5870 ( .A1(n6495), .A2(n4857), .B1(n6557), .B2(n4856), .ZN(n4730)
         );
  OAI21_X1 U5871 ( .B1(n4918), .B2(n6555), .A(n4730), .ZN(n4731) );
  AOI21_X1 U5872 ( .B1(n5234), .B2(n4756), .A(n4731), .ZN(n4732) );
  OAI21_X1 U5873 ( .B1(n4855), .B2(n4733), .A(n4732), .ZN(U3134) );
  INV_X1 U5874 ( .A(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4737) );
  AOI22_X1 U5875 ( .A1(n6491), .A2(n4857), .B1(n6550), .B2(n4856), .ZN(n4734)
         );
  OAI21_X1 U5876 ( .B1(n6553), .B2(n4918), .A(n4734), .ZN(n4735) );
  AOI21_X1 U5877 ( .B1(n5250), .B2(n4756), .A(n4735), .ZN(n4736) );
  OAI21_X1 U5878 ( .B1(n4855), .B2(n4737), .A(n4736), .ZN(U3133) );
  INV_X1 U5879 ( .A(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4741) );
  AOI22_X1 U5880 ( .A1(n6499), .A2(n4857), .B1(n6564), .B2(n4856), .ZN(n4738)
         );
  OAI21_X1 U5881 ( .B1(n4918), .B2(n6562), .A(n4738), .ZN(n4739) );
  AOI21_X1 U5882 ( .B1(n5223), .B2(n4756), .A(n4739), .ZN(n4740) );
  OAI21_X1 U5883 ( .B1(n4855), .B2(n4741), .A(n4740), .ZN(U3135) );
  INV_X1 U5884 ( .A(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4745) );
  AOI22_X1 U5885 ( .A1(n6503), .A2(n4857), .B1(n6571), .B2(n4856), .ZN(n4742)
         );
  OAI21_X1 U5886 ( .B1(n4918), .B2(n6574), .A(n4742), .ZN(n4743) );
  AOI21_X1 U5887 ( .B1(n6504), .B2(n4756), .A(n4743), .ZN(n4744) );
  OAI21_X1 U5888 ( .B1(n4855), .B2(n4745), .A(n4744), .ZN(U3136) );
  INV_X1 U5889 ( .A(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4749) );
  AOI22_X1 U5890 ( .A1(n6511), .A2(n4857), .B1(n6585), .B2(n4856), .ZN(n4746)
         );
  OAI21_X1 U5891 ( .B1(n4918), .B2(n6583), .A(n4746), .ZN(n4747) );
  AOI21_X1 U5892 ( .B1(n6512), .B2(n4756), .A(n4747), .ZN(n4748) );
  OAI21_X1 U5893 ( .B1(n4855), .B2(n4749), .A(n4748), .ZN(U3138) );
  INV_X1 U5894 ( .A(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4753) );
  AOI22_X1 U5895 ( .A1(n6517), .A2(n4857), .B1(n6595), .B2(n4856), .ZN(n4750)
         );
  OAI21_X1 U5896 ( .B1(n4918), .B2(n6591), .A(n4750), .ZN(n4751) );
  AOI21_X1 U5897 ( .B1(n5230), .B2(n4756), .A(n4751), .ZN(n4752) );
  OAI21_X1 U5898 ( .B1(n4855), .B2(n4753), .A(n4752), .ZN(U3139) );
  INV_X1 U5899 ( .A(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4758) );
  AOI22_X1 U5900 ( .A1(n6578), .A2(n4856), .B1(n6507), .B2(n4857), .ZN(n4754)
         );
  OAI21_X1 U5901 ( .B1(n6581), .B2(n4918), .A(n4754), .ZN(n4755) );
  AOI21_X1 U5902 ( .B1(n5218), .B2(n4756), .A(n4755), .ZN(n4757) );
  OAI21_X1 U5903 ( .B1(n4855), .B2(n4758), .A(n4757), .ZN(U3137) );
  NAND2_X1 U5904 ( .A1(n4759), .A2(n5218), .ZN(n4763) );
  AOI22_X1 U5905 ( .A1(n6578), .A2(n4761), .B1(n6507), .B2(n4760), .ZN(n4762)
         );
  OAI211_X1 U5906 ( .C1(n6470), .C2(n6581), .A(n4763), .B(n4762), .ZN(n4764)
         );
  AOI21_X1 U5907 ( .B1(n4765), .B2(INSTQUEUE_REG_2__5__SCAN_IN), .A(n4764), 
        .ZN(n4766) );
  INV_X1 U5908 ( .A(n4766), .ZN(U3041) );
  NAND2_X1 U5909 ( .A1(n4768), .A2(n4767), .ZN(n4769) );
  NAND2_X1 U5910 ( .A1(n4770), .A2(n4769), .ZN(n6382) );
  INV_X1 U5911 ( .A(EBX_REG_7__SCAN_IN), .ZN(n4772) );
  OAI222_X1 U5912 ( .A1(n6382), .A2(n5689), .B1(n4772), .B2(n6023), .C1(n4771), 
        .C2(n5688), .ZN(U2852) );
  AOI22_X1 U5913 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n4774), .B1(n6578), 
        .B2(n4773), .ZN(n4778) );
  INV_X1 U5914 ( .A(n6507), .ZN(n6575) );
  OAI22_X1 U5915 ( .A1(n4874), .A2(n6581), .B1(n6575), .B2(n4775), .ZN(n4776)
         );
  AOI21_X1 U5916 ( .B1(n5218), .B2(n5032), .A(n4776), .ZN(n4777) );
  NAND2_X1 U5917 ( .A1(n4778), .A2(n4777), .ZN(U3097) );
  NAND2_X1 U5918 ( .A1(n4779), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4791)
         );
  AND2_X1 U5919 ( .A1(n4780), .A2(n4791), .ZN(n4781) );
  NAND2_X1 U5920 ( .A1(n4782), .A2(n4781), .ZN(n6326) );
  NAND2_X1 U5921 ( .A1(n4783), .A2(n4218), .ZN(n4789) );
  INV_X1 U5922 ( .A(n4784), .ZN(n4786) );
  NAND2_X1 U5923 ( .A1(n4786), .A2(n4785), .ZN(n4799) );
  XNOR2_X1 U5924 ( .A(n4799), .B(n4800), .ZN(n4787) );
  NAND2_X1 U5925 ( .A1(n4787), .A2(n6240), .ZN(n4788) );
  NAND2_X1 U5926 ( .A1(n4789), .A2(n4788), .ZN(n4794) );
  INV_X1 U5927 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6388) );
  XNOR2_X1 U5928 ( .A(n4794), .B(n6388), .ZN(n6328) );
  INV_X1 U5929 ( .A(n4790), .ZN(n4792) );
  NAND2_X1 U5930 ( .A1(n4792), .A2(n4791), .ZN(n6325) );
  AND2_X1 U5931 ( .A1(n6328), .A2(n6325), .ZN(n4793) );
  NAND2_X1 U5932 ( .A1(n6326), .A2(n4793), .ZN(n6327) );
  NAND2_X1 U5933 ( .A1(n4794), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4795)
         );
  NAND2_X1 U5934 ( .A1(n6327), .A2(n4795), .ZN(n4803) );
  AND3_X1 U5935 ( .A1(n4797), .A2(n4218), .A3(n4800), .ZN(n4798) );
  INV_X1 U5936 ( .A(n4799), .ZN(n4801) );
  NAND3_X1 U5937 ( .A1(n4801), .A2(n6240), .A3(n4800), .ZN(n4802) );
  NAND2_X1 U5938 ( .A1(n5158), .A2(n4802), .ZN(n5073) );
  XNOR2_X1 U5939 ( .A(n5073), .B(n6381), .ZN(n4804) );
  NAND2_X1 U5940 ( .A1(n4803), .A2(n4804), .ZN(n5156) );
  OAI21_X1 U5941 ( .B1(n4803), .B2(n4804), .A(n5074), .ZN(n6375) );
  INV_X1 U5942 ( .A(n5101), .ZN(n4806) );
  AOI22_X1 U5943 ( .A1(n6350), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .B1(n6422), 
        .B2(REIP_REG_8__SCAN_IN), .ZN(n4805) );
  OAI21_X1 U5944 ( .B1(n6360), .B2(n4806), .A(n4805), .ZN(n4807) );
  AOI21_X1 U5945 ( .B1(n4808), .B2(n6354), .A(n4807), .ZN(n4809) );
  OAI21_X1 U5946 ( .B1(n6375), .B2(n6096), .A(n4809), .ZN(U2978) );
  NOR3_X1 U5947 ( .A1(n4843), .A2(n4914), .A3(n6537), .ZN(n4810) );
  OAI21_X1 U5948 ( .B1(n4810), .B2(n5016), .A(n4816), .ZN(n4814) );
  NOR2_X1 U5949 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4811), .ZN(n4846)
         );
  INV_X1 U5950 ( .A(n4846), .ZN(n4812) );
  NOR2_X1 U5951 ( .A1(n5019), .A2(n5020), .ZN(n5204) );
  OAI21_X1 U5952 ( .B1(n5204), .B2(n6636), .A(n5022), .ZN(n5212) );
  AOI211_X1 U5953 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4812), .A(n5296), .B(
        n5212), .ZN(n4813) );
  INV_X1 U5954 ( .A(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4820) );
  INV_X1 U5955 ( .A(n4914), .ZN(n4841) );
  NAND2_X1 U5956 ( .A1(n5204), .A2(n5303), .ZN(n4815) );
  OAI21_X1 U5957 ( .B1(n4816), .B2(n6537), .A(n4815), .ZN(n4847) );
  AOI22_X1 U5958 ( .A1(n6511), .A2(n4846), .B1(n6585), .B2(n4847), .ZN(n4817)
         );
  OAI21_X1 U5959 ( .B1(n4841), .B2(n6588), .A(n4817), .ZN(n4818) );
  AOI21_X1 U5960 ( .B1(n4843), .B2(n5318), .A(n4818), .ZN(n4819) );
  OAI21_X1 U5961 ( .B1(n4854), .B2(n4820), .A(n4819), .ZN(U3026) );
  AOI22_X1 U5962 ( .A1(n6503), .A2(n4846), .B1(n6571), .B2(n4847), .ZN(n4821)
         );
  OAI21_X1 U5963 ( .B1(n4841), .B2(n6569), .A(n4821), .ZN(n4822) );
  AOI21_X1 U5964 ( .B1(n4843), .B2(n5314), .A(n4822), .ZN(n4823) );
  OAI21_X1 U5965 ( .B1(n4854), .B2(n4824), .A(n4823), .ZN(U3024) );
  AOI22_X1 U5966 ( .A1(n6495), .A2(n4846), .B1(n6557), .B2(n4847), .ZN(n4825)
         );
  OAI21_X1 U5967 ( .B1(n4841), .B2(n6560), .A(n4825), .ZN(n4826) );
  AOI21_X1 U5968 ( .B1(n4843), .B2(n6496), .A(n4826), .ZN(n4827) );
  OAI21_X1 U5969 ( .B1(n4854), .B2(n4828), .A(n4827), .ZN(U3022) );
  INV_X1 U5970 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4832) );
  AOI22_X1 U5971 ( .A1(n6491), .A2(n4846), .B1(n6550), .B2(n4847), .ZN(n4829)
         );
  OAI21_X1 U5972 ( .B1(n4841), .B2(n6548), .A(n4829), .ZN(n4830) );
  AOI21_X1 U5973 ( .B1(n4843), .B2(n6492), .A(n4830), .ZN(n4831) );
  OAI21_X1 U5974 ( .B1(n4854), .B2(n4832), .A(n4831), .ZN(U3021) );
  INV_X1 U5975 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4836) );
  AOI22_X1 U5976 ( .A1(n6477), .A2(n4846), .B1(n6543), .B2(n4847), .ZN(n4833)
         );
  OAI21_X1 U5977 ( .B1(n6528), .B2(n4841), .A(n4833), .ZN(n4834) );
  AOI21_X1 U5978 ( .B1(n4843), .B2(n5328), .A(n4834), .ZN(n4835) );
  OAI21_X1 U5979 ( .B1(n4854), .B2(n4836), .A(n4835), .ZN(U3020) );
  AOI22_X1 U5980 ( .A1(n6499), .A2(n4846), .B1(n6564), .B2(n4847), .ZN(n4837)
         );
  OAI21_X1 U5981 ( .B1(n4841), .B2(n6567), .A(n4837), .ZN(n4838) );
  AOI21_X1 U5982 ( .B1(n4843), .B2(n6500), .A(n4838), .ZN(n4839) );
  OAI21_X1 U5983 ( .B1(n4854), .B2(n3641), .A(n4839), .ZN(U3023) );
  AOI22_X1 U5984 ( .A1(n6517), .A2(n4846), .B1(n6595), .B2(n4847), .ZN(n4840)
         );
  OAI21_X1 U5985 ( .B1(n4841), .B2(n6600), .A(n4840), .ZN(n4842) );
  AOI21_X1 U5986 ( .B1(n4843), .B2(n6519), .A(n4842), .ZN(n4844) );
  OAI21_X1 U5987 ( .B1(n4854), .B2(n4845), .A(n4844), .ZN(U3027) );
  AOI22_X1 U5988 ( .A1(n6578), .A2(n4847), .B1(n6507), .B2(n4846), .ZN(n4849)
         );
  NAND2_X1 U5989 ( .A1(n4914), .A2(n5218), .ZN(n4848) );
  OAI211_X1 U5990 ( .C1(n4850), .C2(n6581), .A(n4849), .B(n4848), .ZN(n4851)
         );
  INV_X1 U5991 ( .A(n4851), .ZN(n4852) );
  OAI21_X1 U5992 ( .B1(n4854), .B2(n4853), .A(n4852), .ZN(U3025) );
  INV_X1 U5993 ( .A(n4855), .ZN(n4863) );
  AOI22_X1 U5994 ( .A1(n6477), .A2(n4857), .B1(n6543), .B2(n4856), .ZN(n4860)
         );
  NAND2_X1 U5995 ( .A1(n4858), .A2(n5328), .ZN(n4859) );
  OAI211_X1 U5996 ( .C1(n4861), .C2(n6528), .A(n4860), .B(n4859), .ZN(n4862)
         );
  AOI21_X1 U5997 ( .B1(n4863), .B2(INSTQUEUE_REG_14__0__SCAN_IN), .A(n4862), 
        .ZN(n4864) );
  INV_X1 U5998 ( .A(n4864), .ZN(U3132) );
  NAND3_X1 U5999 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n6620), .ZN(n6540) );
  NOR2_X1 U6000 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6540), .ZN(n4903)
         );
  NAND2_X1 U6001 ( .A1(n6599), .A2(n4874), .ZN(n4865) );
  NAND2_X1 U6002 ( .A1(n4865), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4866) );
  NAND2_X1 U6003 ( .A1(n4866), .A2(n6530), .ZN(n4873) );
  INV_X1 U6004 ( .A(n4873), .ZN(n4868) );
  NAND2_X1 U6005 ( .A1(n4867), .A2(n6189), .ZN(n6534) );
  AOI22_X1 U6006 ( .A1(n4868), .A2(n6534), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4929), .ZN(n4869) );
  OAI211_X1 U6007 ( .C1(n4903), .C2(n6709), .A(n4870), .B(n4869), .ZN(n4871)
         );
  INV_X1 U6008 ( .A(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n4878) );
  OAI22_X1 U6009 ( .A1(n4873), .A2(n6534), .B1(n4929), .B2(n4872), .ZN(n4907)
         );
  INV_X1 U6010 ( .A(n4874), .ZN(n4904) );
  AOI22_X1 U6011 ( .A1(n4904), .A2(n5234), .B1(n6495), .B2(n4903), .ZN(n4875)
         );
  OAI21_X1 U6012 ( .B1(n6555), .B2(n6599), .A(n4875), .ZN(n4876) );
  AOI21_X1 U6013 ( .B1(n4907), .B2(n6557), .A(n4876), .ZN(n4877) );
  OAI21_X1 U6014 ( .B1(n4910), .B2(n4878), .A(n4877), .ZN(U3102) );
  INV_X1 U6015 ( .A(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4882) );
  AOI22_X1 U6016 ( .A1(n4904), .A2(n6478), .B1(n6477), .B2(n4903), .ZN(n4879)
         );
  OAI21_X1 U6017 ( .B1(n6546), .B2(n6599), .A(n4879), .ZN(n4880) );
  AOI21_X1 U6018 ( .B1(n4907), .B2(n6543), .A(n4880), .ZN(n4881) );
  OAI21_X1 U6019 ( .B1(n4910), .B2(n4882), .A(n4881), .ZN(U3100) );
  INV_X1 U6020 ( .A(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n4886) );
  AOI22_X1 U6021 ( .A1(n4904), .A2(n5250), .B1(n6491), .B2(n4903), .ZN(n4883)
         );
  OAI21_X1 U6022 ( .B1(n6553), .B2(n6599), .A(n4883), .ZN(n4884) );
  AOI21_X1 U6023 ( .B1(n4907), .B2(n6550), .A(n4884), .ZN(n4885) );
  OAI21_X1 U6024 ( .B1(n4910), .B2(n4886), .A(n4885), .ZN(U3101) );
  INV_X1 U6025 ( .A(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4890) );
  AOI22_X1 U6026 ( .A1(n4904), .A2(n6512), .B1(n6511), .B2(n4903), .ZN(n4887)
         );
  OAI21_X1 U6027 ( .B1(n6583), .B2(n6599), .A(n4887), .ZN(n4888) );
  AOI21_X1 U6028 ( .B1(n4907), .B2(n6585), .A(n4888), .ZN(n4889) );
  OAI21_X1 U6029 ( .B1(n4910), .B2(n4890), .A(n4889), .ZN(U3106) );
  INV_X1 U6030 ( .A(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4894) );
  AOI22_X1 U6031 ( .A1(n4904), .A2(n5218), .B1(n6507), .B2(n4903), .ZN(n4891)
         );
  OAI21_X1 U6032 ( .B1(n6581), .B2(n6599), .A(n4891), .ZN(n4892) );
  AOI21_X1 U6033 ( .B1(n4907), .B2(n6578), .A(n4892), .ZN(n4893) );
  OAI21_X1 U6034 ( .B1(n4910), .B2(n4894), .A(n4893), .ZN(U3105) );
  INV_X1 U6035 ( .A(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4898) );
  AOI22_X1 U6036 ( .A1(n4904), .A2(n6504), .B1(n6503), .B2(n4903), .ZN(n4895)
         );
  OAI21_X1 U6037 ( .B1(n6574), .B2(n6599), .A(n4895), .ZN(n4896) );
  AOI21_X1 U6038 ( .B1(n4907), .B2(n6571), .A(n4896), .ZN(n4897) );
  OAI21_X1 U6039 ( .B1(n4910), .B2(n4898), .A(n4897), .ZN(U3104) );
  INV_X1 U6040 ( .A(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4902) );
  AOI22_X1 U6041 ( .A1(n4904), .A2(n5230), .B1(n6517), .B2(n4903), .ZN(n4899)
         );
  OAI21_X1 U6042 ( .B1(n6591), .B2(n6599), .A(n4899), .ZN(n4900) );
  AOI21_X1 U6043 ( .B1(n4907), .B2(n6595), .A(n4900), .ZN(n4901) );
  OAI21_X1 U6044 ( .B1(n4910), .B2(n4902), .A(n4901), .ZN(U3107) );
  INV_X1 U6045 ( .A(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4909) );
  AOI22_X1 U6046 ( .A1(n4904), .A2(n5223), .B1(n6499), .B2(n4903), .ZN(n4905)
         );
  OAI21_X1 U6047 ( .B1(n6562), .B2(n6599), .A(n4905), .ZN(n4906) );
  AOI21_X1 U6048 ( .B1(n4907), .B2(n6564), .A(n4906), .ZN(n4908) );
  OAI21_X1 U6049 ( .B1(n4910), .B2(n4909), .A(n4908), .ZN(U3103) );
  INV_X1 U6050 ( .A(n6578), .ZN(n5308) );
  OAI22_X1 U6051 ( .A1(n5308), .A2(n4912), .B1(n4911), .B2(n6575), .ZN(n4913)
         );
  AOI21_X1 U6052 ( .B1(n6508), .B2(n4914), .A(n4913), .ZN(n4917) );
  NAND2_X1 U6053 ( .A1(n4915), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4916)
         );
  OAI211_X1 U6054 ( .C1(n4918), .C2(n6576), .A(n4917), .B(n4916), .ZN(U3145)
         );
  NOR2_X1 U6055 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6486), .ZN(n4962)
         );
  INV_X1 U6056 ( .A(n4962), .ZN(n4926) );
  NAND2_X1 U6057 ( .A1(n5981), .A2(n4919), .ZN(n5986) );
  AOI21_X1 U6058 ( .B1(n5009), .B2(n6525), .A(n6999), .ZN(n4924) );
  NOR2_X1 U6059 ( .A1(n4923), .A2(n4922), .ZN(n6482) );
  NOR2_X1 U6060 ( .A1(n4924), .A2(n6482), .ZN(n4925) );
  AOI22_X1 U6061 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n4926), .B1(n6530), .B2(
        n4925), .ZN(n4928) );
  INV_X1 U6062 ( .A(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4937) );
  NAND2_X1 U6063 ( .A1(n4930), .A2(n5987), .ZN(n4933) );
  NAND2_X1 U6064 ( .A1(n4931), .A2(n4929), .ZN(n4932) );
  NAND2_X1 U6065 ( .A1(n4933), .A2(n4932), .ZN(n4963) );
  AOI22_X1 U6066 ( .A1(n6511), .A2(n4962), .B1(n6585), .B2(n4963), .ZN(n4934)
         );
  OAI21_X1 U6067 ( .B1(n6525), .B2(n6583), .A(n4934), .ZN(n4935) );
  AOI21_X1 U6068 ( .B1(n4966), .B2(n6512), .A(n4935), .ZN(n4936) );
  OAI21_X1 U6069 ( .B1(n3170), .B2(n4937), .A(n4936), .ZN(U3074) );
  INV_X1 U6070 ( .A(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4941) );
  AOI22_X1 U6071 ( .A1(n6491), .A2(n4962), .B1(n6550), .B2(n4963), .ZN(n4938)
         );
  OAI21_X1 U6072 ( .B1(n6525), .B2(n6553), .A(n4938), .ZN(n4939) );
  AOI21_X1 U6073 ( .B1(n4966), .B2(n5250), .A(n4939), .ZN(n4940) );
  OAI21_X1 U6074 ( .B1(n3170), .B2(n4941), .A(n4940), .ZN(U3069) );
  INV_X1 U6075 ( .A(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4945) );
  AOI22_X1 U6076 ( .A1(n6499), .A2(n4962), .B1(n6564), .B2(n4963), .ZN(n4942)
         );
  OAI21_X1 U6077 ( .B1(n6525), .B2(n6562), .A(n4942), .ZN(n4943) );
  AOI21_X1 U6078 ( .B1(n4966), .B2(n5223), .A(n4943), .ZN(n4944) );
  OAI21_X1 U6079 ( .B1(n3170), .B2(n4945), .A(n4944), .ZN(U3071) );
  INV_X1 U6080 ( .A(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4949) );
  AOI22_X1 U6081 ( .A1(n6477), .A2(n4962), .B1(n6543), .B2(n4963), .ZN(n4946)
         );
  OAI21_X1 U6082 ( .B1(n6546), .B2(n6525), .A(n4946), .ZN(n4947) );
  AOI21_X1 U6083 ( .B1(n6478), .B2(n4966), .A(n4947), .ZN(n4948) );
  OAI21_X1 U6084 ( .B1(n3170), .B2(n4949), .A(n4948), .ZN(U3068) );
  INV_X1 U6085 ( .A(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4953) );
  AOI22_X1 U6086 ( .A1(n6495), .A2(n4962), .B1(n6557), .B2(n4963), .ZN(n4950)
         );
  OAI21_X1 U6087 ( .B1(n6525), .B2(n6555), .A(n4950), .ZN(n4951) );
  AOI21_X1 U6088 ( .B1(n4966), .B2(n5234), .A(n4951), .ZN(n4952) );
  OAI21_X1 U6089 ( .B1(n3170), .B2(n4953), .A(n4952), .ZN(U3070) );
  INV_X1 U6090 ( .A(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4957) );
  AOI22_X1 U6091 ( .A1(n6517), .A2(n4962), .B1(n6595), .B2(n4963), .ZN(n4954)
         );
  OAI21_X1 U6092 ( .B1(n6525), .B2(n6591), .A(n4954), .ZN(n4955) );
  AOI21_X1 U6093 ( .B1(n4966), .B2(n5230), .A(n4955), .ZN(n4956) );
  OAI21_X1 U6094 ( .B1(n3170), .B2(n4957), .A(n4956), .ZN(U3075) );
  INV_X1 U6095 ( .A(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4961) );
  AOI22_X1 U6096 ( .A1(n6503), .A2(n4962), .B1(n6571), .B2(n4963), .ZN(n4958)
         );
  OAI21_X1 U6097 ( .B1(n6525), .B2(n6574), .A(n4958), .ZN(n4959) );
  AOI21_X1 U6098 ( .B1(n4966), .B2(n6504), .A(n4959), .ZN(n4960) );
  OAI21_X1 U6099 ( .B1(n3170), .B2(n4961), .A(n4960), .ZN(U3072) );
  INV_X1 U6100 ( .A(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4968) );
  AOI22_X1 U6101 ( .A1(n6578), .A2(n4963), .B1(n4962), .B2(n6507), .ZN(n4964)
         );
  OAI21_X1 U6102 ( .B1(n6525), .B2(n6581), .A(n4964), .ZN(n4965) );
  AOI21_X1 U6103 ( .B1(n4966), .B2(n5218), .A(n4965), .ZN(n4967) );
  OAI21_X1 U6104 ( .B1(n3170), .B2(n4968), .A(n4967), .ZN(U3073) );
  OR2_X1 U6105 ( .A1(n4969), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5208)
         );
  INV_X1 U6106 ( .A(n6481), .ZN(n6536) );
  OAI21_X1 U6107 ( .B1(n4977), .B2(n6999), .A(n6530), .ZN(n4975) );
  NAND2_X1 U6108 ( .A1(n5293), .A2(n4970), .ZN(n5209) );
  NOR2_X1 U6109 ( .A1(n6610), .A2(n5208), .ZN(n5006) );
  INV_X1 U6110 ( .A(n5006), .ZN(n4971) );
  OAI21_X1 U6111 ( .B1(n5209), .B2(n6533), .A(n4971), .ZN(n4973) );
  NOR2_X1 U6112 ( .A1(n4975), .A2(n4973), .ZN(n4972) );
  AOI211_X2 U6113 ( .C1(n5208), .C2(n6537), .A(n6536), .B(n4972), .ZN(n5014)
         );
  INV_X1 U6114 ( .A(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4981) );
  INV_X1 U6115 ( .A(n4973), .ZN(n4974) );
  OAI22_X1 U6116 ( .A1(n4975), .A2(n4974), .B1(n5208), .B2(n6636), .ZN(n5011)
         );
  INV_X1 U6117 ( .A(n5259), .ZN(n5007) );
  AOI22_X1 U6118 ( .A1(n5007), .A2(n5230), .B1(n6517), .B2(n5006), .ZN(n4978)
         );
  OAI21_X1 U6119 ( .B1(n5009), .B2(n6591), .A(n4978), .ZN(n4979) );
  AOI21_X1 U6120 ( .B1(n6595), .B2(n5011), .A(n4979), .ZN(n4980) );
  OAI21_X1 U6121 ( .B1(n5014), .B2(n4981), .A(n4980), .ZN(U3067) );
  INV_X1 U6122 ( .A(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4985) );
  AOI22_X1 U6123 ( .A1(n5007), .A2(n5250), .B1(n6491), .B2(n5006), .ZN(n4982)
         );
  OAI21_X1 U6124 ( .B1(n5009), .B2(n6553), .A(n4982), .ZN(n4983) );
  AOI21_X1 U6125 ( .B1(n6550), .B2(n5011), .A(n4983), .ZN(n4984) );
  OAI21_X1 U6126 ( .B1(n5014), .B2(n4985), .A(n4984), .ZN(U3061) );
  INV_X1 U6127 ( .A(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4989) );
  AOI22_X1 U6128 ( .A1(n5007), .A2(n6512), .B1(n6511), .B2(n5006), .ZN(n4986)
         );
  OAI21_X1 U6129 ( .B1(n5009), .B2(n6583), .A(n4986), .ZN(n4987) );
  AOI21_X1 U6130 ( .B1(n6585), .B2(n5011), .A(n4987), .ZN(n4988) );
  OAI21_X1 U6131 ( .B1(n5014), .B2(n4989), .A(n4988), .ZN(U3066) );
  INV_X1 U6132 ( .A(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4993) );
  AOI22_X1 U6133 ( .A1(n5007), .A2(n5218), .B1(n6507), .B2(n5006), .ZN(n4990)
         );
  OAI21_X1 U6134 ( .B1(n5009), .B2(n6581), .A(n4990), .ZN(n4991) );
  AOI21_X1 U6135 ( .B1(n6578), .B2(n5011), .A(n4991), .ZN(n4992) );
  OAI21_X1 U6136 ( .B1(n5014), .B2(n4993), .A(n4992), .ZN(U3065) );
  INV_X1 U6137 ( .A(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4997) );
  AOI22_X1 U6138 ( .A1(n5007), .A2(n5234), .B1(n6495), .B2(n5006), .ZN(n4994)
         );
  OAI21_X1 U6139 ( .B1(n5009), .B2(n6555), .A(n4994), .ZN(n4995) );
  AOI21_X1 U6140 ( .B1(n6557), .B2(n5011), .A(n4995), .ZN(n4996) );
  OAI21_X1 U6141 ( .B1(n5014), .B2(n4997), .A(n4996), .ZN(U3062) );
  INV_X1 U6142 ( .A(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n5001) );
  AOI22_X1 U6143 ( .A1(n5007), .A2(n5223), .B1(n6499), .B2(n5006), .ZN(n4998)
         );
  OAI21_X1 U6144 ( .B1(n5009), .B2(n6562), .A(n4998), .ZN(n4999) );
  AOI21_X1 U6145 ( .B1(n6564), .B2(n5011), .A(n4999), .ZN(n5000) );
  OAI21_X1 U6146 ( .B1(n5014), .B2(n5001), .A(n5000), .ZN(U3063) );
  INV_X1 U6147 ( .A(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n5005) );
  AOI22_X1 U6148 ( .A1(n5007), .A2(n6478), .B1(n6477), .B2(n5006), .ZN(n5002)
         );
  OAI21_X1 U6149 ( .B1(n5009), .B2(n6546), .A(n5002), .ZN(n5003) );
  AOI21_X1 U6150 ( .B1(n6543), .B2(n5011), .A(n5003), .ZN(n5004) );
  OAI21_X1 U6151 ( .B1(n5014), .B2(n5005), .A(n5004), .ZN(U3060) );
  INV_X1 U6152 ( .A(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n5013) );
  AOI22_X1 U6153 ( .A1(n5007), .A2(n6504), .B1(n6503), .B2(n5006), .ZN(n5008)
         );
  OAI21_X1 U6154 ( .B1(n5009), .B2(n6574), .A(n5008), .ZN(n5010) );
  AOI21_X1 U6155 ( .B1(n6571), .B2(n5011), .A(n5010), .ZN(n5012) );
  OAI21_X1 U6156 ( .B1(n5014), .B2(n5013), .A(n5012), .ZN(U3064) );
  NOR3_X1 U6157 ( .A1(n5032), .A2(n6520), .A3(n6537), .ZN(n5017) );
  OR2_X1 U6158 ( .A1(n5987), .A2(n5015), .ZN(n5026) );
  OAI21_X1 U6159 ( .B1(n5017), .B2(n5016), .A(n5026), .ZN(n5025) );
  NOR2_X1 U6160 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5018), .ZN(n5062)
         );
  INV_X1 U6161 ( .A(n5062), .ZN(n5023) );
  INV_X1 U6162 ( .A(n5019), .ZN(n5021) );
  AND2_X1 U6163 ( .A1(n5021), .A2(n5020), .ZN(n5295) );
  OAI21_X1 U6164 ( .B1(n5295), .B2(n6636), .A(n5022), .ZN(n5302) );
  AOI211_X1 U6165 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5023), .A(n5296), .B(
        n5302), .ZN(n5024) );
  NAND2_X1 U6166 ( .A1(n5025), .A2(n5024), .ZN(n5066) );
  INV_X1 U6167 ( .A(n5066), .ZN(n5035) );
  INV_X1 U6168 ( .A(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n5034) );
  INV_X1 U6169 ( .A(n5026), .ZN(n5027) );
  NAND2_X1 U6170 ( .A1(n5027), .A2(n6530), .ZN(n5029) );
  NAND2_X1 U6171 ( .A1(n5295), .A2(n5303), .ZN(n5028) );
  NAND2_X1 U6172 ( .A1(n5029), .A2(n5028), .ZN(n5061) );
  AOI22_X1 U6173 ( .A1(n6578), .A2(n5061), .B1(n6507), .B2(n5062), .ZN(n5030)
         );
  OAI21_X1 U6174 ( .B1(n6576), .B2(n6516), .A(n5030), .ZN(n5031) );
  AOI21_X1 U6175 ( .B1(n6508), .B2(n5032), .A(n5031), .ZN(n5033) );
  OAI21_X1 U6176 ( .B1(n5035), .B2(n5034), .A(n5033), .ZN(U3089) );
  NOR2_X1 U6177 ( .A1(n5060), .A2(n6591), .ZN(n5038) );
  AOI22_X1 U6178 ( .A1(n6517), .A2(n5062), .B1(n6595), .B2(n5061), .ZN(n5036)
         );
  OAI21_X1 U6179 ( .B1(n6600), .B2(n6516), .A(n5036), .ZN(n5037) );
  AOI211_X1 U6180 ( .C1(n5066), .C2(INSTQUEUE_REG_8__7__SCAN_IN), .A(n5038), 
        .B(n5037), .ZN(n5039) );
  INV_X1 U6181 ( .A(n5039), .ZN(U3091) );
  NOR2_X1 U6182 ( .A1(n5060), .A2(n6553), .ZN(n5042) );
  AOI22_X1 U6183 ( .A1(n6491), .A2(n5062), .B1(n6550), .B2(n5061), .ZN(n5040)
         );
  OAI21_X1 U6184 ( .B1(n6548), .B2(n6516), .A(n5040), .ZN(n5041) );
  AOI211_X1 U6185 ( .C1(n5066), .C2(INSTQUEUE_REG_8__1__SCAN_IN), .A(n5042), 
        .B(n5041), .ZN(n5043) );
  INV_X1 U6186 ( .A(n5043), .ZN(U3085) );
  NOR2_X1 U6187 ( .A1(n5060), .A2(n6555), .ZN(n5046) );
  AOI22_X1 U6188 ( .A1(n6495), .A2(n5062), .B1(n6557), .B2(n5061), .ZN(n5044)
         );
  OAI21_X1 U6189 ( .B1(n6560), .B2(n6516), .A(n5044), .ZN(n5045) );
  AOI211_X1 U6190 ( .C1(n5066), .C2(INSTQUEUE_REG_8__2__SCAN_IN), .A(n5046), 
        .B(n5045), .ZN(n5047) );
  INV_X1 U6191 ( .A(n5047), .ZN(U3086) );
  NOR2_X1 U6192 ( .A1(n5060), .A2(n6574), .ZN(n5050) );
  AOI22_X1 U6193 ( .A1(n6503), .A2(n5062), .B1(n6571), .B2(n5061), .ZN(n5048)
         );
  OAI21_X1 U6194 ( .B1(n6569), .B2(n6516), .A(n5048), .ZN(n5049) );
  AOI211_X1 U6195 ( .C1(n5066), .C2(INSTQUEUE_REG_8__4__SCAN_IN), .A(n5050), 
        .B(n5049), .ZN(n5051) );
  INV_X1 U6196 ( .A(n5051), .ZN(U3088) );
  NOR2_X1 U6197 ( .A1(n5060), .A2(n6562), .ZN(n5054) );
  AOI22_X1 U6198 ( .A1(n6499), .A2(n5062), .B1(n6564), .B2(n5061), .ZN(n5052)
         );
  OAI21_X1 U6199 ( .B1(n6567), .B2(n6516), .A(n5052), .ZN(n5053) );
  AOI211_X1 U6200 ( .C1(n5066), .C2(INSTQUEUE_REG_8__3__SCAN_IN), .A(n5054), 
        .B(n5053), .ZN(n5055) );
  INV_X1 U6201 ( .A(n5055), .ZN(U3087) );
  NOR2_X1 U6202 ( .A1(n5060), .A2(n6583), .ZN(n5058) );
  AOI22_X1 U6203 ( .A1(n6511), .A2(n5062), .B1(n6585), .B2(n5061), .ZN(n5056)
         );
  OAI21_X1 U6204 ( .B1(n6588), .B2(n6516), .A(n5056), .ZN(n5057) );
  AOI211_X1 U6205 ( .C1(n5066), .C2(INSTQUEUE_REG_8__6__SCAN_IN), .A(n5058), 
        .B(n5057), .ZN(n5059) );
  INV_X1 U6206 ( .A(n5059), .ZN(U3090) );
  NOR2_X1 U6207 ( .A1(n5060), .A2(n6546), .ZN(n5065) );
  AOI22_X1 U6208 ( .A1(n6477), .A2(n5062), .B1(n6543), .B2(n5061), .ZN(n5063)
         );
  OAI21_X1 U6209 ( .B1(n6528), .B2(n6516), .A(n5063), .ZN(n5064) );
  AOI211_X1 U6210 ( .C1(n5066), .C2(INSTQUEUE_REG_8__0__SCAN_IN), .A(n5065), 
        .B(n5064), .ZN(n5067) );
  INV_X1 U6211 ( .A(n5067), .ZN(U3084) );
  OAI21_X1 U6212 ( .B1(n3176), .B2(n3770), .A(n5080), .ZN(n5244) );
  INV_X1 U6213 ( .A(DATAI_9_), .ZN(n6811) );
  INV_X1 U6214 ( .A(EAX_REG_9__SCAN_IN), .ZN(n6303) );
  OAI222_X1 U6215 ( .A1(n5244), .A2(n6024), .B1(n5291), .B2(n6811), .C1(n5698), 
        .C2(n6303), .ZN(U2882) );
  AOI21_X1 U6216 ( .B1(n5070), .B2(n5069), .A(n5093), .ZN(n6369) );
  INV_X1 U6217 ( .A(n6369), .ZN(n5072) );
  INV_X1 U6218 ( .A(EBX_REG_9__SCAN_IN), .ZN(n5071) );
  OAI222_X1 U6219 ( .A1(n5072), .A2(n5689), .B1(n6023), .B2(n5071), .C1(n5244), 
        .C2(n5688), .ZN(U2850) );
  NAND2_X1 U6220 ( .A1(n5073), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n5154)
         );
  NAND2_X1 U6221 ( .A1(n5074), .A2(n5154), .ZN(n5085) );
  INV_X1 U6222 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n5372) );
  OR2_X1 U6223 ( .A1(n5158), .A2(n5372), .ZN(n5153) );
  NAND2_X1 U6224 ( .A1(n5158), .A2(n5372), .ZN(n5152) );
  NAND2_X1 U6225 ( .A1(n5153), .A2(n5152), .ZN(n5075) );
  XNOR2_X1 U6226 ( .A(n5085), .B(n5075), .ZN(n6371) );
  NAND2_X1 U6227 ( .A1(n6371), .A2(n6356), .ZN(n5078) );
  AND2_X1 U6228 ( .A1(n6422), .A2(REIP_REG_9__SCAN_IN), .ZN(n6368) );
  NOR2_X1 U6229 ( .A1(n6360), .A2(n5238), .ZN(n5076) );
  AOI211_X1 U6230 ( .C1(n6350), .C2(PHYADDRPOINTER_REG_9__SCAN_IN), .A(n6368), 
        .B(n5076), .ZN(n5077) );
  OAI211_X1 U6231 ( .C1(n6043), .C2(n5244), .A(n5078), .B(n5077), .ZN(U2977)
         );
  AND2_X1 U6232 ( .A1(n5080), .A2(n5079), .ZN(n5082) );
  OR2_X1 U6233 ( .A1(n5082), .A2(n5116), .ZN(n6158) );
  AOI22_X1 U6234 ( .A1(n5720), .A2(DATAI_10_), .B1(n6213), .B2(
        EAX_REG_10__SCAN_IN), .ZN(n5083) );
  OAI21_X1 U6235 ( .B1(n6158), .B2(n6024), .A(n5083), .ZN(U2881) );
  INV_X1 U6236 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5084) );
  NAND2_X1 U6237 ( .A1(n5158), .A2(n5084), .ZN(n5151) );
  NAND2_X1 U6238 ( .A1(n5283), .A2(n5151), .ZN(n5088) );
  NAND2_X1 U6239 ( .A1(n5085), .A2(n5152), .ZN(n5086) );
  NAND2_X1 U6240 ( .A1(n5086), .A2(n5153), .ZN(n5087) );
  XOR2_X1 U6241 ( .A(n5088), .B(n5087), .Z(n5192) );
  NAND2_X1 U6242 ( .A1(INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n6378) );
  INV_X1 U6243 ( .A(n6378), .ZN(n5097) );
  NAND2_X1 U6244 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n5096), .ZN(n5376)
         );
  NAND4_X1 U6245 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_6__SCAN_IN), .A3(n6421), .A4(n6402), .ZN(n5375) );
  INV_X1 U6246 ( .A(n5375), .ZN(n5089) );
  NOR2_X1 U6247 ( .A1(n5423), .A2(n5089), .ZN(n5090) );
  INV_X1 U6248 ( .A(n5373), .ZN(n5427) );
  AOI211_X1 U6249 ( .C1(n6399), .C2(n5376), .A(n5090), .B(n5427), .ZN(n6389)
         );
  OAI21_X1 U6250 ( .B1(n5438), .B2(n5097), .A(n6389), .ZN(n6370) );
  NOR2_X1 U6251 ( .A1(n5093), .A2(n5092), .ZN(n5094) );
  OR2_X1 U6252 ( .A1(n5091), .A2(n5094), .ZN(n6149) );
  INV_X1 U6253 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6683) );
  OAI22_X1 U6254 ( .A1(n6149), .A2(n6391), .B1(n6683), .B2(n6407), .ZN(n5099)
         );
  NAND2_X1 U6255 ( .A1(n6426), .A2(n5095), .ZN(n6400) );
  NAND2_X1 U6256 ( .A1(n5096), .A2(n6400), .ZN(n6397) );
  NOR2_X1 U6257 ( .A1(n6396), .A2(n6397), .ZN(n6384) );
  NAND2_X1 U6258 ( .A1(n5097), .A2(n6384), .ZN(n6374) );
  AOI221_X1 U6259 ( .B1(INSTADDRPOINTER_REG_9__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .C1(n5372), .C2(n5084), .A(n6374), 
        .ZN(n5098) );
  AOI211_X1 U6260 ( .C1(INSTADDRPOINTER_REG_10__SCAN_IN), .C2(n6370), .A(n5099), .B(n5098), .ZN(n5100) );
  OAI21_X1 U6261 ( .B1(n5192), .B2(n6403), .A(n5100), .ZN(U3008) );
  NAND2_X1 U6262 ( .A1(n6193), .A2(n5101), .ZN(n5104) );
  NAND2_X1 U6263 ( .A1(n6194), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n5103)
         );
  NAND2_X1 U6264 ( .A1(n5267), .A2(n5102), .ZN(n6165) );
  NAND3_X1 U6265 ( .A1(n5104), .A2(n5103), .A3(n6165), .ZN(n5107) );
  NOR2_X1 U6266 ( .A1(n6123), .A2(n5105), .ZN(n5106) );
  AOI211_X1 U6267 ( .C1(n6377), .C2(n6153), .A(n5107), .B(n5106), .ZN(n5111)
         );
  NAND3_X1 U6268 ( .A1(n5237), .A2(REIP_REG_5__SCAN_IN), .A3(n6179), .ZN(n6166) );
  OAI21_X1 U6269 ( .B1(n5108), .B2(n6166), .A(n6681), .ZN(n5109) );
  OAI21_X1 U6270 ( .B1(n6181), .B2(n5236), .A(n5267), .ZN(n6155) );
  NAND2_X1 U6271 ( .A1(n5109), .A2(n6155), .ZN(n5110) );
  OAI211_X1 U6272 ( .C1(n5112), .C2(n6157), .A(n5111), .B(n5110), .ZN(U2819)
         );
  INV_X1 U6273 ( .A(EBX_REG_10__SCAN_IN), .ZN(n5113) );
  OAI222_X1 U6274 ( .A1(n6158), .A2(n5691), .B1(n5113), .B2(n6023), .C1(n5689), 
        .C2(n6149), .ZN(U2849) );
  NOR2_X1 U6275 ( .A1(n5116), .A2(n5115), .ZN(n5117) );
  OR2_X1 U6276 ( .A1(n5114), .A2(n5117), .ZN(n5187) );
  OR2_X1 U6277 ( .A1(n5091), .A2(n5118), .ZN(n5119) );
  AND2_X1 U6278 ( .A1(n5148), .A2(n5119), .ZN(n6362) );
  NOR2_X1 U6279 ( .A1(n6023), .A2(n5183), .ZN(n5120) );
  AOI21_X1 U6280 ( .B1(n6362), .B2(n6018), .A(n5120), .ZN(n5121) );
  OAI21_X1 U6281 ( .B1(n5187), .B2(n5691), .A(n5121), .ZN(U2848) );
  INV_X1 U6282 ( .A(n5478), .ZN(n5122) );
  OR2_X1 U6283 ( .A1(n5127), .A2(n5122), .ZN(n5123) );
  NAND2_X1 U6284 ( .A1(n5123), .A2(n6157), .ZN(n6200) );
  INV_X1 U6285 ( .A(n6200), .ZN(n5202) );
  OAI22_X1 U6286 ( .A1(n5125), .A2(n6123), .B1(n6198), .B2(n5124), .ZN(n5131)
         );
  INV_X1 U6287 ( .A(n4203), .ZN(n5126) );
  NOR2_X1 U6288 ( .A1(n5127), .A2(n5126), .ZN(n6190) );
  INV_X1 U6289 ( .A(n6190), .ZN(n5129) );
  OAI21_X1 U6290 ( .B1(n6194), .B2(n6193), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n5128) );
  OAI21_X1 U6291 ( .B1(n5129), .B2(n6533), .A(n5128), .ZN(n5130) );
  AOI211_X1 U6292 ( .C1(REIP_REG_0__SCAN_IN), .C2(n5628), .A(n5131), .B(n5130), 
        .ZN(n5132) );
  OAI21_X1 U6293 ( .B1(n5202), .B2(n5133), .A(n5132), .ZN(U2827) );
  NAND2_X1 U6294 ( .A1(n5237), .A2(n6710), .ZN(n5193) );
  NAND2_X1 U6295 ( .A1(n5193), .A2(n5267), .ZN(n6188) );
  AOI22_X1 U6296 ( .A1(n6190), .A2(n5134), .B1(n6153), .B2(n6423), .ZN(n5139)
         );
  INV_X1 U6297 ( .A(n6359), .ZN(n5135) );
  AOI22_X1 U6298 ( .A1(PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n6194), .B1(n6193), 
        .B2(n5135), .ZN(n5138) );
  INV_X1 U6299 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6187) );
  NAND3_X1 U6300 ( .A1(n5237), .A2(REIP_REG_1__SCAN_IN), .A3(n6187), .ZN(n5137) );
  NAND2_X1 U6301 ( .A1(n6191), .A2(EBX_REG_2__SCAN_IN), .ZN(n5136) );
  NAND4_X1 U6302 ( .A1(n5139), .A2(n5138), .A3(n5137), .A4(n5136), .ZN(n5140)
         );
  AOI21_X1 U6303 ( .B1(REIP_REG_2__SCAN_IN), .B2(n6188), .A(n5140), .ZN(n5141)
         );
  OAI21_X1 U6304 ( .B1(n5142), .B2(n5202), .A(n5141), .ZN(U2825) );
  OR2_X1 U6305 ( .A1(n5114), .A2(n5143), .ZN(n5144) );
  NAND2_X1 U6306 ( .A1(n5145), .A2(n5144), .ZN(n6145) );
  AOI22_X1 U6307 ( .A1(n5720), .A2(DATAI_12_), .B1(n6213), .B2(
        EAX_REG_12__SCAN_IN), .ZN(n5146) );
  OAI21_X1 U6308 ( .B1(n6145), .B2(n6024), .A(n5146), .ZN(U2879) );
  INV_X1 U6309 ( .A(n5274), .ZN(n5147) );
  AOI21_X1 U6310 ( .B1(n5149), .B2(n5148), .A(n5147), .ZN(n6135) );
  AOI22_X1 U6311 ( .A1(n6135), .A2(n6018), .B1(EBX_REG_12__SCAN_IN), .B2(n5668), .ZN(n5150) );
  OAI21_X1 U6312 ( .B1(n6145), .B2(n5691), .A(n5150), .ZN(U2847) );
  AND2_X1 U6313 ( .A1(n5152), .A2(n5151), .ZN(n5278) );
  AND2_X1 U6314 ( .A1(n5154), .A2(n5153), .ZN(n5155) );
  NAND2_X1 U6315 ( .A1(n5156), .A2(n5155), .ZN(n5282) );
  NAND2_X1 U6316 ( .A1(n5278), .A2(n5282), .ZN(n5157) );
  NAND2_X1 U6317 ( .A1(n5157), .A2(n5283), .ZN(n5160) );
  INV_X1 U6318 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5284) );
  XNOR2_X1 U6319 ( .A(n5849), .B(n5284), .ZN(n5159) );
  XNOR2_X1 U6320 ( .A(n5160), .B(n5159), .ZN(n6363) );
  NAND2_X1 U6321 ( .A1(n6363), .A2(n6356), .ZN(n5163) );
  AND2_X1 U6322 ( .A1(n6422), .A2(REIP_REG_11__SCAN_IN), .ZN(n6361) );
  NOR2_X1 U6323 ( .A1(n6360), .A2(n5180), .ZN(n5161) );
  AOI211_X1 U6324 ( .C1(n6350), .C2(PHYADDRPOINTER_REG_11__SCAN_IN), .A(n6361), 
        .B(n5161), .ZN(n5162) );
  OAI211_X1 U6325 ( .C1(n6043), .C2(n5187), .A(n5163), .B(n5162), .ZN(U2975)
         );
  NOR3_X1 U6326 ( .A1(n6181), .A2(REIP_REG_4__SCAN_IN), .A3(n5165), .ZN(n5173)
         );
  INV_X1 U6327 ( .A(n6405), .ZN(n5171) );
  INV_X1 U6328 ( .A(n5164), .ZN(n5168) );
  INV_X1 U6329 ( .A(n5267), .ZN(n5629) );
  OAI21_X1 U6330 ( .B1(n5629), .B2(n5165), .A(n5628), .ZN(n6203) );
  OAI22_X1 U6331 ( .A1(n6203), .A2(n6676), .B1(n5166), .B2(n6176), .ZN(n5167)
         );
  AOI211_X1 U6332 ( .C1(n6193), .C2(n5168), .A(n5167), .B(n6178), .ZN(n5170)
         );
  NAND2_X1 U6333 ( .A1(n6191), .A2(EBX_REG_4__SCAN_IN), .ZN(n5169) );
  OAI211_X1 U6334 ( .C1(n5171), .C2(n6198), .A(n5170), .B(n5169), .ZN(n5172)
         );
  AOI211_X1 U6335 ( .C1(n6190), .C2(n5174), .A(n5173), .B(n5172), .ZN(n5175)
         );
  OAI21_X1 U6336 ( .B1(n5176), .B2(n5202), .A(n5175), .ZN(U2823) );
  INV_X1 U6337 ( .A(DATAI_11_), .ZN(n5177) );
  INV_X1 U6338 ( .A(EAX_REG_11__SCAN_IN), .ZN(n6309) );
  OAI222_X1 U6339 ( .A1(n5187), .A2(n6024), .B1(n5291), .B2(n5177), .C1(n5698), 
        .C2(n6309), .ZN(U2880) );
  INV_X1 U6340 ( .A(n6121), .ZN(n5178) );
  NAND3_X1 U6341 ( .A1(n5237), .A2(n6684), .A3(n5178), .ZN(n5179) );
  OAI21_X1 U6342 ( .B1(n5180), .B2(n6186), .A(n5179), .ZN(n5185) );
  OAI21_X1 U6343 ( .B1(n6181), .B2(n5181), .A(n5267), .ZN(n6142) );
  AOI22_X1 U6344 ( .A1(PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n6194), .B1(
        REIP_REG_11__SCAN_IN), .B2(n6142), .ZN(n5182) );
  OAI211_X1 U6345 ( .C1(n6123), .C2(n5183), .A(n5182), .B(n6165), .ZN(n5184)
         );
  AOI211_X1 U6346 ( .C1(n6362), .C2(n6153), .A(n5185), .B(n5184), .ZN(n5186)
         );
  OAI21_X1 U6347 ( .B1(n5187), .B2(n6157), .A(n5186), .ZN(U2816) );
  INV_X1 U6348 ( .A(n6158), .ZN(n5190) );
  AOI22_X1 U6349 ( .A1(n6350), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .B1(n6422), 
        .B2(REIP_REG_10__SCAN_IN), .ZN(n5188) );
  OAI21_X1 U6350 ( .B1(n6360), .B2(n6156), .A(n5188), .ZN(n5189) );
  AOI21_X1 U6351 ( .B1(n5190), .B2(n6354), .A(n5189), .ZN(n5191) );
  OAI21_X1 U6352 ( .B1(n5192), .B2(n6096), .A(n5191), .ZN(U2976) );
  INV_X1 U6353 ( .A(n5193), .ZN(n5199) );
  AOI22_X1 U6354 ( .A1(n5195), .A2(n6190), .B1(n6153), .B2(n5194), .ZN(n5197)
         );
  AOI22_X1 U6355 ( .A1(n6194), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .B1(n5629), 
        .B2(REIP_REG_1__SCAN_IN), .ZN(n5196) );
  OAI211_X1 U6356 ( .C1(PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n6186), .A(n5197), 
        .B(n5196), .ZN(n5198) );
  AOI211_X1 U6357 ( .C1(n6191), .C2(EBX_REG_1__SCAN_IN), .A(n5199), .B(n5198), 
        .ZN(n5200) );
  OAI21_X1 U6358 ( .B1(n5202), .B2(n5201), .A(n5200), .ZN(U2826) );
  INV_X1 U6359 ( .A(n5204), .ZN(n5207) );
  INV_X1 U6360 ( .A(n5296), .ZN(n5206) );
  NAND3_X1 U6361 ( .A1(n5987), .A2(n6530), .A3(n5293), .ZN(n5205) );
  OAI21_X1 U6362 ( .B1(n5207), .B2(n5206), .A(n5205), .ZN(n5253) );
  INV_X1 U6363 ( .A(n5253), .ZN(n5216) );
  NOR2_X1 U6364 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5208), .ZN(n5220)
         );
  INV_X1 U6365 ( .A(n5209), .ZN(n5211) );
  AOI21_X1 U6366 ( .B1(n5259), .B2(n6476), .A(n6999), .ZN(n5210) );
  NOR3_X1 U6367 ( .A1(n5211), .A2(n5210), .A3(n6537), .ZN(n5213) );
  NOR3_X1 U6368 ( .A1(n5303), .A2(n5213), .A3(n5212), .ZN(n5214) );
  AOI22_X1 U6369 ( .A1(n6507), .A2(n5220), .B1(INSTQUEUE_REG_4__5__SCAN_IN), 
        .B2(n5252), .ZN(n5215) );
  OAI21_X1 U6370 ( .B1(n5308), .B2(n5216), .A(n5215), .ZN(n5217) );
  AOI21_X1 U6371 ( .B1(n5218), .B2(n5257), .A(n5217), .ZN(n5219) );
  OAI21_X1 U6372 ( .B1(n6581), .B2(n5259), .A(n5219), .ZN(U3057) );
  INV_X1 U6373 ( .A(n5220), .ZN(n5255) );
  AOI22_X1 U6374 ( .A1(n5253), .A2(n6564), .B1(INSTQUEUE_REG_4__3__SCAN_IN), 
        .B2(n5252), .ZN(n5221) );
  OAI21_X1 U6375 ( .B1(n6561), .B2(n5255), .A(n5221), .ZN(n5222) );
  AOI21_X1 U6376 ( .B1(n5223), .B2(n5257), .A(n5222), .ZN(n5224) );
  OAI21_X1 U6377 ( .B1(n6562), .B2(n5259), .A(n5224), .ZN(U3055) );
  AOI22_X1 U6378 ( .A1(n5253), .A2(n6543), .B1(INSTQUEUE_REG_4__0__SCAN_IN), 
        .B2(n5252), .ZN(n5225) );
  OAI21_X1 U6379 ( .B1(n6527), .B2(n5255), .A(n5225), .ZN(n5226) );
  AOI21_X1 U6380 ( .B1(n6478), .B2(n5257), .A(n5226), .ZN(n5227) );
  OAI21_X1 U6381 ( .B1(n6546), .B2(n5259), .A(n5227), .ZN(U3052) );
  AOI22_X1 U6382 ( .A1(n5253), .A2(n6595), .B1(INSTQUEUE_REG_4__7__SCAN_IN), 
        .B2(n5252), .ZN(n5228) );
  OAI21_X1 U6383 ( .B1(n6590), .B2(n5255), .A(n5228), .ZN(n5229) );
  AOI21_X1 U6384 ( .B1(n5230), .B2(n5257), .A(n5229), .ZN(n5231) );
  OAI21_X1 U6385 ( .B1(n6591), .B2(n5259), .A(n5231), .ZN(U3059) );
  AOI22_X1 U6386 ( .A1(n5253), .A2(n6557), .B1(INSTQUEUE_REG_4__2__SCAN_IN), 
        .B2(n5252), .ZN(n5232) );
  OAI21_X1 U6387 ( .B1(n6554), .B2(n5255), .A(n5232), .ZN(n5233) );
  AOI21_X1 U6388 ( .B1(n5234), .B2(n5257), .A(n5233), .ZN(n5235) );
  OAI21_X1 U6389 ( .B1(n6555), .B2(n5259), .A(n5235), .ZN(U3054) );
  NAND2_X1 U6390 ( .A1(n5237), .A2(n5236), .ZN(n6150) );
  OAI22_X1 U6391 ( .A1(n6150), .A2(REIP_REG_9__SCAN_IN), .B1(n5238), .B2(n6186), .ZN(n5242) );
  AOI22_X1 U6392 ( .A1(EBX_REG_9__SCAN_IN), .A2(n6191), .B1(
        REIP_REG_9__SCAN_IN), .B2(n6155), .ZN(n5239) );
  OAI211_X1 U6393 ( .C1(n6176), .C2(n5240), .A(n5239), .B(n6165), .ZN(n5241)
         );
  AOI211_X1 U6394 ( .C1(n6369), .C2(n6153), .A(n5242), .B(n5241), .ZN(n5243)
         );
  OAI21_X1 U6395 ( .B1(n6157), .B2(n5244), .A(n5243), .ZN(U2818) );
  AOI22_X1 U6396 ( .A1(n5253), .A2(n6571), .B1(INSTQUEUE_REG_4__4__SCAN_IN), 
        .B2(n5252), .ZN(n5245) );
  OAI21_X1 U6397 ( .B1(n6568), .B2(n5255), .A(n5245), .ZN(n5246) );
  AOI21_X1 U6398 ( .B1(n6504), .B2(n5257), .A(n5246), .ZN(n5247) );
  OAI21_X1 U6399 ( .B1(n6574), .B2(n5259), .A(n5247), .ZN(U3056) );
  AOI22_X1 U6400 ( .A1(n5253), .A2(n6550), .B1(INSTQUEUE_REG_4__1__SCAN_IN), 
        .B2(n5252), .ZN(n5248) );
  OAI21_X1 U6401 ( .B1(n6547), .B2(n5255), .A(n5248), .ZN(n5249) );
  AOI21_X1 U6402 ( .B1(n5250), .B2(n5257), .A(n5249), .ZN(n5251) );
  OAI21_X1 U6403 ( .B1(n6553), .B2(n5259), .A(n5251), .ZN(U3053) );
  AOI22_X1 U6404 ( .A1(n5253), .A2(n6585), .B1(INSTQUEUE_REG_4__6__SCAN_IN), 
        .B2(n5252), .ZN(n5254) );
  OAI21_X1 U6405 ( .B1(n6582), .B2(n5255), .A(n5254), .ZN(n5256) );
  AOI21_X1 U6406 ( .B1(n6512), .B2(n5257), .A(n5256), .ZN(n5258) );
  OAI21_X1 U6407 ( .B1(n6583), .B2(n5259), .A(n5258), .ZN(U3058) );
  OAI22_X1 U6408 ( .A1(n5261), .A2(n6186), .B1(n6176), .B2(n5260), .ZN(n5263)
         );
  OAI22_X1 U6409 ( .A1(n6123), .A2(n4550), .B1(n6198), .B2(n6392), .ZN(n5262)
         );
  NOR2_X1 U6410 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6166), .ZN(n6172) );
  NOR4_X1 U6411 ( .A1(n5263), .A2(n5262), .A3(n6178), .A4(n6172), .ZN(n5269)
         );
  INV_X1 U6412 ( .A(n5264), .ZN(n5266) );
  INV_X1 U6413 ( .A(n5628), .ZN(n5265) );
  AOI21_X1 U6414 ( .B1(n5267), .B2(n5266), .A(n5265), .ZN(n6183) );
  NAND2_X1 U6415 ( .A1(n6183), .A2(REIP_REG_6__SCAN_IN), .ZN(n5268) );
  OAI211_X1 U6416 ( .C1(n5270), .C2(n6157), .A(n5269), .B(n5268), .ZN(U2821)
         );
  OAI21_X1 U6417 ( .B1(n5273), .B2(n5272), .A(n5271), .ZN(n6127) );
  AOI21_X1 U6418 ( .B1(n5275), .B2(n5274), .A(n5626), .ZN(n6126) );
  AOI22_X1 U6419 ( .A1(n6126), .A2(n6018), .B1(EBX_REG_13__SCAN_IN), .B2(n5668), .ZN(n5276) );
  OAI21_X1 U6420 ( .B1(n6127), .B2(n5691), .A(n5276), .ZN(U2846) );
  AND2_X1 U6421 ( .A1(n5158), .A2(n5284), .ZN(n5280) );
  INV_X1 U6422 ( .A(n5278), .ZN(n5279) );
  NOR2_X1 U6423 ( .A1(n5280), .A2(n5279), .ZN(n5281) );
  NAND2_X1 U6424 ( .A1(n5282), .A2(n5281), .ZN(n5287) );
  INV_X1 U6425 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5396) );
  NOR2_X1 U6426 ( .A1(n5849), .A2(n5396), .ZN(n5392) );
  NAND2_X1 U6427 ( .A1(n5849), .A2(n5396), .ZN(n5390) );
  XNOR2_X1 U6428 ( .A(n5158), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5360)
         );
  XNOR2_X1 U6429 ( .A(n5361), .B(n5360), .ZN(n6085) );
  NAND2_X1 U6430 ( .A1(n6085), .A2(n6356), .ZN(n5290) );
  AND2_X1 U6431 ( .A1(n6422), .A2(REIP_REG_13__SCAN_IN), .ZN(n6083) );
  NOR2_X1 U6432 ( .A1(n6360), .A2(n6128), .ZN(n5288) );
  AOI211_X1 U6433 ( .C1(n6350), .C2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n6083), 
        .B(n5288), .ZN(n5289) );
  OAI211_X1 U6434 ( .C1(n6043), .C2(n6127), .A(n5290), .B(n5289), .ZN(U2973)
         );
  INV_X1 U6435 ( .A(DATAI_13_), .ZN(n7097) );
  INV_X1 U6436 ( .A(EAX_REG_13__SCAN_IN), .ZN(n6315) );
  OAI222_X1 U6437 ( .A1(n6127), .A2(n6024), .B1(n5291), .B2(n7097), .C1(n6315), 
        .C2(n5698), .ZN(U2878) );
  INV_X1 U6438 ( .A(n5293), .ZN(n5294) );
  NOR2_X1 U6439 ( .A1(n5987), .A2(n5294), .ZN(n5299) );
  AOI22_X1 U6440 ( .A1(n5299), .A2(n6530), .B1(n5296), .B2(n5295), .ZN(n5311)
         );
  NAND2_X1 U6441 ( .A1(n6610), .A2(n5297), .ZN(n5336) );
  INV_X1 U6442 ( .A(n5336), .ZN(n5306) );
  INV_X1 U6443 ( .A(n5338), .ZN(n5298) );
  AOI21_X1 U6444 ( .B1(n5298), .B2(n6592), .A(n6999), .ZN(n5300) );
  NOR3_X1 U6445 ( .A1(n5300), .A2(n5299), .A3(n6537), .ZN(n5301) );
  AOI211_X1 U6446 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5336), .A(n5302), .B(
        n5301), .ZN(n5305) );
  INV_X1 U6447 ( .A(n5303), .ZN(n5304) );
  NAND2_X1 U6448 ( .A1(n5305), .A2(n5304), .ZN(n5333) );
  AOI22_X1 U6449 ( .A1(n6507), .A2(n5306), .B1(INSTQUEUE_REG_12__5__SCAN_IN), 
        .B2(n5333), .ZN(n5307) );
  OAI21_X1 U6450 ( .B1(n5308), .B2(n5311), .A(n5307), .ZN(n5309) );
  AOI21_X1 U6451 ( .B1(n6508), .B2(n5338), .A(n5309), .ZN(n5310) );
  OAI21_X1 U6452 ( .B1(n6576), .B2(n6592), .A(n5310), .ZN(U3121) );
  INV_X1 U6453 ( .A(n5311), .ZN(n5334) );
  AOI22_X1 U6454 ( .A1(n5334), .A2(n6571), .B1(INSTQUEUE_REG_12__4__SCAN_IN), 
        .B2(n5333), .ZN(n5312) );
  OAI21_X1 U6455 ( .B1(n6568), .B2(n5336), .A(n5312), .ZN(n5313) );
  AOI21_X1 U6456 ( .B1(n5314), .B2(n5338), .A(n5313), .ZN(n5315) );
  OAI21_X1 U6457 ( .B1(n6569), .B2(n6592), .A(n5315), .ZN(U3120) );
  AOI22_X1 U6458 ( .A1(n5334), .A2(n6585), .B1(INSTQUEUE_REG_12__6__SCAN_IN), 
        .B2(n5333), .ZN(n5316) );
  OAI21_X1 U6459 ( .B1(n6582), .B2(n5336), .A(n5316), .ZN(n5317) );
  AOI21_X1 U6460 ( .B1(n5318), .B2(n5338), .A(n5317), .ZN(n5319) );
  OAI21_X1 U6461 ( .B1(n6588), .B2(n6592), .A(n5319), .ZN(U3122) );
  AOI22_X1 U6462 ( .A1(n5334), .A2(n6550), .B1(INSTQUEUE_REG_12__1__SCAN_IN), 
        .B2(n5333), .ZN(n5320) );
  OAI21_X1 U6463 ( .B1(n6547), .B2(n5336), .A(n5320), .ZN(n5321) );
  AOI21_X1 U6464 ( .B1(n6492), .B2(n5338), .A(n5321), .ZN(n5322) );
  OAI21_X1 U6465 ( .B1(n6548), .B2(n6592), .A(n5322), .ZN(U3117) );
  AOI22_X1 U6466 ( .A1(n5334), .A2(n6557), .B1(INSTQUEUE_REG_12__2__SCAN_IN), 
        .B2(n5333), .ZN(n5323) );
  OAI21_X1 U6467 ( .B1(n6554), .B2(n5336), .A(n5323), .ZN(n5324) );
  AOI21_X1 U6468 ( .B1(n6496), .B2(n5338), .A(n5324), .ZN(n5325) );
  OAI21_X1 U6469 ( .B1(n6560), .B2(n6592), .A(n5325), .ZN(U3118) );
  AOI22_X1 U6470 ( .A1(n5334), .A2(n6543), .B1(INSTQUEUE_REG_12__0__SCAN_IN), 
        .B2(n5333), .ZN(n5326) );
  OAI21_X1 U6471 ( .B1(n6527), .B2(n5336), .A(n5326), .ZN(n5327) );
  AOI21_X1 U6472 ( .B1(n5328), .B2(n5338), .A(n5327), .ZN(n5329) );
  OAI21_X1 U6473 ( .B1(n6528), .B2(n6592), .A(n5329), .ZN(U3116) );
  AOI22_X1 U6474 ( .A1(n5334), .A2(n6595), .B1(INSTQUEUE_REG_12__7__SCAN_IN), 
        .B2(n5333), .ZN(n5330) );
  OAI21_X1 U6475 ( .B1(n6590), .B2(n5336), .A(n5330), .ZN(n5331) );
  AOI21_X1 U6476 ( .B1(n6519), .B2(n5338), .A(n5331), .ZN(n5332) );
  OAI21_X1 U6477 ( .B1(n6600), .B2(n6592), .A(n5332), .ZN(U3123) );
  AOI22_X1 U6478 ( .A1(n5334), .A2(n6564), .B1(INSTQUEUE_REG_12__3__SCAN_IN), 
        .B2(n5333), .ZN(n5335) );
  OAI21_X1 U6479 ( .B1(n6561), .B2(n5336), .A(n5335), .ZN(n5337) );
  AOI21_X1 U6480 ( .B1(n6500), .B2(n5338), .A(n5337), .ZN(n5339) );
  OAI21_X1 U6481 ( .B1(n6567), .B2(n6592), .A(n5339), .ZN(U3119) );
  AND2_X1 U6482 ( .A1(n5650), .A2(n5341), .ZN(n5588) );
  NAND2_X1 U6483 ( .A1(n5650), .A2(n5342), .ZN(n5661) );
  MUX2_X1 U6484 ( .A(n5664), .B(n5345), .S(n5344), .Z(n5591) );
  NOR2_X1 U6485 ( .A1(n5679), .A2(n5591), .ZN(n5590) );
  XNOR2_X1 U6486 ( .A(n5590), .B(n5346), .ZN(n5965) );
  AOI22_X1 U6487 ( .A1(n5965), .A2(n6018), .B1(EBX_REG_19__SCAN_IN), .B2(n5668), .ZN(n5347) );
  OAI21_X1 U6488 ( .B1(n6035), .B2(n5691), .A(n5347), .ZN(U2840) );
  NOR2_X1 U6489 ( .A1(n5348), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n5349)
         );
  AOI21_X1 U6490 ( .B1(n5351), .B2(n5350), .A(n5349), .ZN(n6613) );
  INV_X1 U6491 ( .A(n5463), .ZN(n5354) );
  AOI22_X1 U6492 ( .A1(n6637), .A2(n5359), .B1(STATE2_REG_1__SCAN_IN), .B2(
        n5352), .ZN(n5353) );
  OAI21_X1 U6493 ( .B1(n6613), .B2(n5354), .A(n5353), .ZN(n5356) );
  AND2_X1 U6494 ( .A1(n5355), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n6611)
         );
  AOI22_X1 U6495 ( .A1(n5358), .A2(n5356), .B1(n5463), .B2(n6611), .ZN(n5357)
         );
  OAI21_X1 U6496 ( .B1(n5359), .B2(n5358), .A(n5357), .ZN(U3461) );
  NAND2_X1 U6497 ( .A1(n5361), .A2(n5360), .ZN(n5364) );
  INV_X1 U6498 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5362) );
  NAND2_X1 U6499 ( .A1(n5849), .A2(n5362), .ZN(n5363) );
  NAND2_X1 U6500 ( .A1(n5364), .A2(n5363), .ZN(n5847) );
  INV_X1 U6501 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5848) );
  OAI21_X2 U6502 ( .B1(n5847), .B2(n5366), .A(n5365), .ZN(n5839) );
  INV_X1 U6503 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n6064) );
  NOR2_X1 U6504 ( .A1(n5849), .A2(n6064), .ZN(n5368) );
  NAND2_X1 U6505 ( .A1(n5849), .A2(n6064), .ZN(n5367) );
  OAI21_X2 U6506 ( .B1(n5839), .B2(n5368), .A(n5367), .ZN(n6039) );
  INV_X1 U6507 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5409) );
  NOR2_X1 U6508 ( .A1(n5277), .A2(n5409), .ZN(n6041) );
  NOR2_X1 U6509 ( .A1(n5849), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n6040)
         );
  NOR2_X1 U6510 ( .A1(n6041), .A2(n6040), .ZN(n5369) );
  XNOR2_X1 U6511 ( .A(n6039), .B(n5369), .ZN(n5388) );
  XNOR2_X1 U6512 ( .A(n5678), .B(n5370), .ZN(n5683) );
  INV_X1 U6513 ( .A(REIP_REG_16__SCAN_IN), .ZN(n5371) );
  NOR2_X1 U6514 ( .A1(n6407), .A2(n5371), .ZN(n5384) );
  INV_X1 U6515 ( .A(n5438), .ZN(n5951) );
  NAND2_X1 U6516 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n6082) );
  NOR2_X1 U6517 ( .A1(n5362), .A2(n6082), .ZN(n6076) );
  NAND2_X1 U6518 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n6076), .ZN(n5422) );
  NOR3_X1 U6519 ( .A1(n5372), .A2(n5084), .A3(n6378), .ZN(n5374) );
  AOI22_X1 U6520 ( .A1(n5438), .A2(n5373), .B1(n5374), .B2(n6389), .ZN(n6364)
         );
  AOI21_X1 U6521 ( .B1(n5951), .B2(n5422), .A(n6364), .ZN(n6065) );
  INV_X1 U6522 ( .A(n5374), .ZN(n5377) );
  NOR2_X1 U6523 ( .A1(n5375), .A2(n5377), .ZN(n5424) );
  NAND2_X1 U6524 ( .A1(n5424), .A2(n6419), .ZN(n5394) );
  NOR2_X1 U6525 ( .A1(n5377), .A2(n5376), .ZN(n5425) );
  NAND2_X1 U6526 ( .A1(n6399), .A2(n5425), .ZN(n6071) );
  NAND2_X1 U6527 ( .A1(n5394), .A2(n6071), .ZN(n6066) );
  NAND2_X1 U6528 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5439) );
  OAI21_X1 U6529 ( .B1(INSTADDRPOINTER_REG_15__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .A(n5439), .ZN(n5378) );
  OAI22_X1 U6530 ( .A1(n6065), .A2(n5409), .B1(n6057), .B2(n5378), .ZN(n5379)
         );
  AOI211_X1 U6531 ( .C1(n6424), .C2(n5683), .A(n5384), .B(n5379), .ZN(n5380)
         );
  OAI21_X1 U6532 ( .B1(n5388), .B2(n6403), .A(n5380), .ZN(U3002) );
  INV_X1 U6533 ( .A(n5673), .ZN(n5382) );
  AOI21_X1 U6534 ( .B1(n6350), .B2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n5384), 
        .ZN(n5385) );
  OAI21_X1 U6535 ( .B1(n5600), .B2(n6360), .A(n5385), .ZN(n5386) );
  AOI21_X1 U6536 ( .B1(n6212), .B2(n6337), .A(n5386), .ZN(n5387) );
  OAI21_X1 U6537 ( .B1(n5388), .B2(n6096), .A(n5387), .ZN(U2970) );
  INV_X1 U6538 ( .A(n5390), .ZN(n5391) );
  NOR2_X1 U6539 ( .A1(n5392), .A2(n5391), .ZN(n5393) );
  XNOR2_X1 U6540 ( .A(n5389), .B(n5393), .ZN(n5405) );
  AOI21_X1 U6541 ( .B1(n6426), .B2(n5394), .A(INSTADDRPOINTER_REG_11__SCAN_IN), 
        .ZN(n5395) );
  OAI21_X1 U6542 ( .B1(n6364), .B2(n5395), .A(INSTADDRPOINTER_REG_12__SCAN_IN), 
        .ZN(n5399) );
  NAND3_X1 U6543 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n5396), .A3(n6066), .ZN(n5398) );
  AOI22_X1 U6544 ( .A1(n6135), .A2(n6424), .B1(n6422), .B2(
        REIP_REG_12__SCAN_IN), .ZN(n5397) );
  AND3_X1 U6545 ( .A1(n5399), .A2(n5398), .A3(n5397), .ZN(n5400) );
  OAI21_X1 U6546 ( .B1(n5405), .B2(n6403), .A(n5400), .ZN(U3006) );
  INV_X1 U6547 ( .A(n6360), .ZN(n5843) );
  INV_X1 U6548 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n6136) );
  INV_X1 U6549 ( .A(REIP_REG_12__SCAN_IN), .ZN(n5401) );
  OAI22_X1 U6550 ( .A1(n6047), .A2(n6136), .B1(n6407), .B2(n5401), .ZN(n5403)
         );
  NOR2_X1 U6551 ( .A1(n6145), .A2(n6043), .ZN(n5402) );
  AOI211_X1 U6552 ( .C1(n5843), .C2(n6143), .A(n5403), .B(n5402), .ZN(n5404)
         );
  OAI21_X1 U6553 ( .B1(n5405), .B2(n6096), .A(n5404), .ZN(U2974) );
  INV_X1 U6554 ( .A(EBX_REG_30__SCAN_IN), .ZN(n5406) );
  OAI222_X1 U6555 ( .A1(n5688), .A2(n5701), .B1(n5406), .B2(n6023), .C1(n5689), 
        .C2(n5445), .ZN(U2829) );
  AND2_X1 U6556 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5440) );
  NAND2_X1 U6557 ( .A1(n5440), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5407) );
  INV_X1 U6558 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5952) );
  INV_X1 U6559 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6055) );
  AND3_X1 U6560 ( .A1(n5952), .A2(n5409), .A3(n6055), .ZN(n5410) );
  NOR2_X1 U6561 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5413) );
  INV_X1 U6562 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5933) );
  INV_X1 U6563 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5412) );
  NAND4_X1 U6564 ( .A1(n5413), .A2(n5933), .A3(n5412), .A4(n5955), .ZN(n5416)
         );
  AND2_X1 U6565 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5791) );
  AND2_X1 U6566 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5954) );
  AND2_X1 U6567 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5443) );
  NAND2_X1 U6568 ( .A1(n3159), .A2(n3167), .ZN(n5414) );
  NAND2_X1 U6569 ( .A1(n5414), .A2(n5849), .ZN(n5415) );
  OAI21_X2 U6570 ( .B1(n5823), .B2(n5416), .A(n5415), .ZN(n5775) );
  XNOR2_X1 U6571 ( .A(n5849), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5774)
         );
  NAND2_X2 U6572 ( .A1(n5775), .A2(n5774), .ZN(n5773) );
  INV_X1 U6573 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5907) );
  NAND2_X1 U6574 ( .A1(n5849), .A2(n5907), .ZN(n5417) );
  NAND2_X2 U6575 ( .A1(n5773), .A2(n5417), .ZN(n5741) );
  NAND2_X1 U6576 ( .A1(n5849), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5761) );
  AND2_X1 U6577 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5874) );
  NAND2_X1 U6578 ( .A1(n5754), .A2(n5874), .ZN(n5734) );
  NOR2_X2 U6579 ( .A1(n5734), .A2(n5873), .ZN(n5725) );
  OR2_X1 U6580 ( .A1(n5849), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5762)
         );
  INV_X1 U6581 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5892) );
  NAND2_X1 U6582 ( .A1(n5879), .A2(n5892), .ZN(n5883) );
  NOR2_X1 U6583 ( .A1(n5762), .A2(n5883), .ZN(n5732) );
  NAND2_X1 U6584 ( .A1(n5732), .A2(n5873), .ZN(n5723) );
  INV_X1 U6585 ( .A(n5723), .ZN(n5418) );
  NOR2_X1 U6586 ( .A1(n5422), .A2(n5439), .ZN(n5426) );
  AOI21_X1 U6587 ( .B1(n5424), .B2(n5426), .A(n5423), .ZN(n5430) );
  AOI21_X1 U6588 ( .B1(n5426), .B2(n5425), .A(n6426), .ZN(n5428) );
  OR2_X1 U6589 ( .A1(n5428), .A2(n5427), .ZN(n5429) );
  NOR2_X1 U6590 ( .A1(n5430), .A2(n5429), .ZN(n6056) );
  AND2_X1 U6591 ( .A1(n5954), .A2(n5440), .ZN(n5431) );
  OR2_X1 U6592 ( .A1(n5438), .A2(n5431), .ZN(n5432) );
  NAND2_X1 U6593 ( .A1(n6056), .A2(n5432), .ZN(n5945) );
  NOR2_X1 U6594 ( .A1(n5438), .A2(n5791), .ZN(n5433) );
  OR2_X1 U6595 ( .A1(n5945), .A2(n5433), .ZN(n5925) );
  OR2_X1 U6596 ( .A1(n6419), .A2(n6399), .ZN(n5949) );
  INV_X1 U6597 ( .A(n5443), .ZN(n5434) );
  AND2_X1 U6598 ( .A1(n5949), .A2(n5434), .ZN(n5435) );
  NAND2_X1 U6599 ( .A1(n5914), .A2(n5438), .ZN(n5858) );
  AND2_X1 U6600 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5444) );
  NAND2_X1 U6601 ( .A1(n5914), .A2(n5444), .ZN(n5436) );
  NAND2_X1 U6602 ( .A1(n5858), .A2(n5436), .ZN(n5888) );
  INV_X1 U6603 ( .A(n5874), .ZN(n5882) );
  NAND2_X1 U6604 ( .A1(n5858), .A2(n5882), .ZN(n5437) );
  AND2_X1 U6605 ( .A1(n5888), .A2(n5437), .ZN(n5870) );
  OAI211_X1 U6606 ( .C1(INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n5438), .A(n5870), .B(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5859) );
  NAND2_X1 U6607 ( .A1(n6052), .A2(n5440), .ZN(n5968) );
  INV_X1 U6608 ( .A(n5954), .ZN(n5441) );
  INV_X1 U6609 ( .A(n5791), .ZN(n5442) );
  NOR2_X1 U6610 ( .A1(n5948), .A2(n5442), .ZN(n5930) );
  NAND3_X1 U6611 ( .A1(n5893), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(n5874), .ZN(n5863) );
  NAND2_X1 U6612 ( .A1(n5863), .A2(n5420), .ZN(n5447) );
  NAND2_X1 U6613 ( .A1(n6422), .A2(REIP_REG_30__SCAN_IN), .ZN(n5450) );
  AOI21_X1 U6614 ( .B1(n5859), .B2(n5447), .A(n5446), .ZN(n5448) );
  OAI21_X1 U6615 ( .B1(n5456), .B2(n6403), .A(n5448), .ZN(U2988) );
  NAND2_X1 U6616 ( .A1(n5843), .A2(n5449), .ZN(n5451) );
  OAI211_X1 U6617 ( .C1(n6047), .C2(n5452), .A(n5451), .B(n5450), .ZN(n5453)
         );
  AOI21_X1 U6618 ( .B1(n5454), .B2(n6354), .A(n5453), .ZN(n5455) );
  OAI21_X1 U6619 ( .B1(n5456), .B2(n6096), .A(n5455), .ZN(U2956) );
  AOI21_X1 U6620 ( .B1(n6637), .B2(n5457), .A(n5466), .ZN(n5468) );
  INV_X1 U6621 ( .A(n5458), .ZN(n5461) );
  NAND3_X1 U6622 ( .A1(n6637), .A2(n4368), .A3(n5467), .ZN(n5459) );
  OAI21_X1 U6623 ( .B1(n5461), .B2(n5460), .A(n5459), .ZN(n5462) );
  AOI21_X1 U6624 ( .B1(n5464), .B2(n5463), .A(n5462), .ZN(n5465) );
  OAI22_X1 U6625 ( .A1(n5468), .A2(n5467), .B1(n5466), .B2(n5465), .ZN(U3459)
         );
  INV_X1 U6626 ( .A(n5469), .ZN(n5477) );
  OR2_X1 U6627 ( .A1(n6602), .A2(n5480), .ZN(n5471) );
  NOR2_X1 U6628 ( .A1(n5471), .A2(n5470), .ZN(n5472) );
  OR2_X1 U6629 ( .A1(n5479), .A2(n5472), .ZN(n5475) );
  NAND2_X1 U6630 ( .A1(n5479), .A2(n5473), .ZN(n5474) );
  OAI211_X1 U6631 ( .C1(n5477), .C2(n5476), .A(n5475), .B(n5474), .ZN(n6603)
         );
  OR2_X1 U6632 ( .A1(n5479), .A2(n5478), .ZN(n5484) );
  INV_X1 U6633 ( .A(n5480), .ZN(n5482) );
  NAND2_X1 U6634 ( .A1(n5482), .A2(n5481), .ZN(n5483) );
  NAND2_X1 U6635 ( .A1(n5484), .A2(n5483), .ZN(n6090) );
  AOI21_X1 U6636 ( .B1(n5485), .B2(n6662), .A(READY_N), .ZN(n6722) );
  NOR2_X1 U6637 ( .A1(n6090), .A2(n6722), .ZN(n6604) );
  OR2_X1 U6638 ( .A1(n6604), .A2(n6648), .ZN(n6095) );
  MUX2_X1 U6639 ( .A(n6603), .B(MORE_REG_SCAN_IN), .S(n6095), .Z(U3471) );
  AOI21_X1 U6640 ( .B1(n5487), .B2(n5501), .A(n5486), .ZN(n5739) );
  INV_X1 U6641 ( .A(n5739), .ZN(n5704) );
  NAND2_X1 U6642 ( .A1(n5488), .A2(n5665), .ZN(n5490) );
  NAND2_X1 U6643 ( .A1(n5490), .A2(n5489), .ZN(n5491) );
  NOR2_X1 U6644 ( .A1(n5506), .A2(n5491), .ZN(n5492) );
  OR2_X1 U6645 ( .A1(n5493), .A2(n5492), .ZN(n5868) );
  OAI22_X1 U6646 ( .A1(n5494), .A2(n6176), .B1(n6186), .B2(n5737), .ZN(n5496)
         );
  NOR2_X1 U6647 ( .A1(n5509), .A2(n7100), .ZN(n5495) );
  AOI211_X1 U6648 ( .C1(EBX_REG_29__SCAN_IN), .C2(n6191), .A(n5496), .B(n5495), 
        .ZN(n5497) );
  OAI21_X1 U6649 ( .B1(n5868), .B2(n6198), .A(n5497), .ZN(n5498) );
  OAI21_X1 U6650 ( .B1(n5704), .B2(n6157), .A(n5500), .ZN(U2798) );
  OAI21_X1 U6651 ( .B1(n5515), .B2(n5502), .A(n5501), .ZN(n5747) );
  INV_X1 U6652 ( .A(n5747), .ZN(n5503) );
  NAND2_X1 U6653 ( .A1(n5503), .A2(n6171), .ZN(n5512) );
  NOR2_X1 U6654 ( .A1(n5517), .A2(n5504), .ZN(n5505) );
  OR2_X1 U6655 ( .A1(n5506), .A2(n5505), .ZN(n5640) );
  INV_X1 U6656 ( .A(n5640), .ZN(n5881) );
  AOI22_X1 U6657 ( .A1(PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n6194), .B1(n6193), 
        .B2(n5750), .ZN(n5508) );
  NAND2_X1 U6658 ( .A1(n6191), .A2(EBX_REG_28__SCAN_IN), .ZN(n5507) );
  OAI211_X1 U6659 ( .C1(n5509), .C2(n7020), .A(n5508), .B(n5507), .ZN(n5510)
         );
  AOI21_X1 U6660 ( .B1(n5881), .B2(n6153), .A(n5510), .ZN(n5511) );
  OAI211_X1 U6661 ( .C1(REIP_REG_28__SCAN_IN), .C2(n5513), .A(n5512), .B(n5511), .ZN(U2799) );
  AOI21_X1 U6662 ( .B1(n5516), .B2(n5530), .A(n5515), .ZN(n5759) );
  INV_X1 U6663 ( .A(n5759), .ZN(n5709) );
  INV_X1 U6664 ( .A(n5517), .ZN(n5520) );
  NAND2_X1 U6665 ( .A1(n5535), .A2(n5518), .ZN(n5519) );
  NAND2_X1 U6666 ( .A1(n5520), .A2(n5519), .ZN(n5889) );
  INV_X1 U6667 ( .A(n5889), .ZN(n5525) );
  OAI22_X1 U6668 ( .A1(n5521), .A2(n6176), .B1(n6186), .B2(n5757), .ZN(n5522)
         );
  AOI21_X1 U6669 ( .B1(n6191), .B2(EBX_REG_27__SCAN_IN), .A(n5522), .ZN(n5523)
         );
  OAI21_X1 U6670 ( .B1(n5532), .B2(n7030), .A(n5523), .ZN(n5524) );
  AOI21_X1 U6671 ( .B1(n5525), .B2(n6153), .A(n5524), .ZN(n5528) );
  NAND3_X1 U6672 ( .A1(n5548), .A2(n5526), .A3(n7030), .ZN(n5527) );
  OAI211_X1 U6673 ( .C1(n5709), .C2(n6157), .A(n5528), .B(n5527), .ZN(U2800)
         );
  OAI21_X1 U6674 ( .B1(n5544), .B2(n5531), .A(n5530), .ZN(n5766) );
  INV_X1 U6675 ( .A(n5548), .ZN(n5562) );
  NAND2_X1 U6676 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_25__SCAN_IN), .ZN(
        n5547) );
  OAI21_X1 U6677 ( .B1(n5562), .B2(n5547), .A(n7050), .ZN(n5541) );
  INV_X1 U6678 ( .A(n5532), .ZN(n5540) );
  NAND2_X1 U6679 ( .A1(n5552), .A2(n5533), .ZN(n5534) );
  NAND2_X1 U6680 ( .A1(n5535), .A2(n5534), .ZN(n5900) );
  OAI22_X1 U6681 ( .A1(n5536), .A2(n6123), .B1(n5765), .B2(n6176), .ZN(n5537)
         );
  AOI21_X1 U6682 ( .B1(n6193), .B2(n5769), .A(n5537), .ZN(n5538) );
  OAI21_X1 U6683 ( .B1(n5900), .B2(n6198), .A(n5538), .ZN(n5539) );
  AOI21_X1 U6684 ( .B1(n5541), .B2(n5540), .A(n5539), .ZN(n5542) );
  OAI21_X1 U6685 ( .B1(n5766), .B2(n6157), .A(n5542), .ZN(U2801) );
  AOI21_X1 U6686 ( .B1(n5545), .B2(n5543), .A(n5544), .ZN(n5546) );
  INV_X1 U6687 ( .A(n5546), .ZN(n5778) );
  OAI211_X1 U6688 ( .C1(REIP_REG_24__SCAN_IN), .C2(REIP_REG_25__SCAN_IN), .A(
        n5548), .B(n5547), .ZN(n5558) );
  NAND2_X1 U6689 ( .A1(n5549), .A2(n5550), .ZN(n5551) );
  NAND2_X1 U6690 ( .A1(n5552), .A2(n5551), .ZN(n5645) );
  INV_X1 U6691 ( .A(n5645), .ZN(n5910) );
  OAI22_X1 U6692 ( .A1(n5553), .A2(n6176), .B1(n6186), .B2(n5771), .ZN(n5554)
         );
  AOI21_X1 U6693 ( .B1(n6191), .B2(EBX_REG_25__SCAN_IN), .A(n5554), .ZN(n5555)
         );
  OAI21_X1 U6694 ( .B1(n6003), .B2(n6825), .A(n5555), .ZN(n5556) );
  AOI21_X1 U6695 ( .B1(n5910), .B2(n6153), .A(n5556), .ZN(n5557) );
  OAI211_X1 U6696 ( .C1(n5778), .C2(n6157), .A(n5558), .B(n5557), .ZN(U2802)
         );
  OAI21_X1 U6697 ( .B1(n5796), .B2(n5560), .A(n5543), .ZN(n5784) );
  OAI21_X1 U6698 ( .B1(n5921), .B2(n5561), .A(n5549), .ZN(n5647) );
  INV_X1 U6699 ( .A(n5647), .ZN(n5918) );
  INV_X1 U6700 ( .A(EBX_REG_24__SCAN_IN), .ZN(n5563) );
  OAI22_X1 U6701 ( .A1(n6123), .A2(n5563), .B1(REIP_REG_24__SCAN_IN), .B2(
        n5562), .ZN(n5566) );
  AOI22_X1 U6702 ( .A1(PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n6194), .B1(n5785), 
        .B2(n6193), .ZN(n5564) );
  OAI21_X1 U6703 ( .B1(n6003), .B2(n7017), .A(n5564), .ZN(n5565) );
  AOI211_X1 U6704 ( .C1(n5918), .C2(n6153), .A(n5566), .B(n5565), .ZN(n5567)
         );
  OAI21_X1 U6705 ( .B1(n5784), .B2(n6157), .A(n5567), .ZN(U2803) );
  OAI21_X1 U6706 ( .B1(n5652), .B2(n5570), .A(n5569), .ZN(n5805) );
  NOR2_X1 U6707 ( .A1(n6693), .A2(n5576), .ZN(n5995) );
  AND2_X1 U6708 ( .A1(n5657), .A2(n5571), .ZN(n5572) );
  OR2_X1 U6709 ( .A1(n5572), .A2(n5923), .ZN(n5936) );
  AOI22_X1 U6710 ( .A1(PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n6194), .B1(n6193), 
        .B2(n5808), .ZN(n5574) );
  NAND2_X1 U6711 ( .A1(n6191), .A2(EBX_REG_22__SCAN_IN), .ZN(n5573) );
  OAI211_X1 U6712 ( .C1(n5936), .C2(n6198), .A(n5574), .B(n5573), .ZN(n5575)
         );
  AOI21_X1 U6713 ( .B1(n5995), .B2(n7106), .A(n5575), .ZN(n5578) );
  NOR2_X1 U6714 ( .A1(REIP_REG_21__SCAN_IN), .A2(n5576), .ZN(n6006) );
  OAI21_X1 U6715 ( .B1(n6006), .B2(n6011), .A(REIP_REG_22__SCAN_IN), .ZN(n5577) );
  OAI211_X1 U6716 ( .C1(n5805), .C2(n6157), .A(n5578), .B(n5577), .ZN(U2805)
         );
  AOI22_X1 U6717 ( .A1(n6861), .A2(n6012), .B1(PHYADDRPOINTER_REG_19__SCAN_IN), 
        .B2(n6194), .ZN(n5586) );
  INV_X1 U6718 ( .A(n5825), .ZN(n5579) );
  AOI21_X1 U6719 ( .B1(n6193), .B2(n5579), .A(n6178), .ZN(n5580) );
  OAI21_X1 U6720 ( .B1(n5581), .B2(n6123), .A(n5580), .ZN(n5584) );
  INV_X1 U6721 ( .A(REIP_REG_18__SCAN_IN), .ZN(n7073) );
  NAND2_X1 U6722 ( .A1(n5582), .A2(n7073), .ZN(n5594) );
  AOI21_X1 U6723 ( .B1(n5594), .B2(n6111), .A(n6861), .ZN(n5583) );
  AOI211_X1 U6724 ( .C1(n6153), .C2(n5965), .A(n5584), .B(n5583), .ZN(n5585)
         );
  OAI211_X1 U6725 ( .C1(n6035), .C2(n6157), .A(n5586), .B(n5585), .ZN(U2808)
         );
  NAND2_X1 U6726 ( .A1(n5650), .A2(n5587), .ZN(n5675) );
  AOI21_X1 U6727 ( .B1(n5589), .B2(n5675), .A(n5588), .ZN(n6204) );
  INV_X1 U6728 ( .A(n6204), .ZN(n5837) );
  AOI21_X1 U6729 ( .B1(n5679), .B2(n5591), .A(n5590), .ZN(n5671) );
  INV_X1 U6730 ( .A(n5835), .ZN(n5593) );
  OAI22_X1 U6731 ( .A1(n6186), .A2(n5593), .B1(n6123), .B2(n5592), .ZN(n5597)
         );
  AOI21_X1 U6732 ( .B1(n6194), .B2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n6178), 
        .ZN(n5595) );
  OAI211_X1 U6733 ( .C1(n6111), .C2(n7073), .A(n5595), .B(n5594), .ZN(n5596)
         );
  AOI211_X1 U6734 ( .C1(n5671), .C2(n6153), .A(n5597), .B(n5596), .ZN(n5598)
         );
  OAI21_X1 U6735 ( .B1(n5837), .B2(n6157), .A(n5598), .ZN(U2809) );
  INV_X1 U6736 ( .A(n6212), .ZN(n5686) );
  NAND2_X1 U6737 ( .A1(n6194), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5599)
         );
  OAI211_X1 U6738 ( .C1(n6186), .C2(n5600), .A(n6165), .B(n5599), .ZN(n5604)
         );
  NAND2_X1 U6739 ( .A1(REIP_REG_16__SCAN_IN), .A2(REIP_REG_15__SCAN_IN), .ZN(
        n6112) );
  OAI21_X1 U6740 ( .B1(REIP_REG_16__SCAN_IN), .B2(REIP_REG_15__SCAN_IN), .A(
        n6112), .ZN(n5602) );
  AOI22_X1 U6741 ( .A1(EBX_REG_16__SCAN_IN), .A2(n6191), .B1(
        REIP_REG_16__SCAN_IN), .B2(n5613), .ZN(n5601) );
  OAI21_X1 U6742 ( .B1(n6113), .B2(n5602), .A(n5601), .ZN(n5603) );
  AOI211_X1 U6743 ( .C1(n6153), .C2(n5683), .A(n5604), .B(n5603), .ZN(n5605)
         );
  OAI21_X1 U6744 ( .B1(n5686), .B2(n6157), .A(n5605), .ZN(U2811) );
  INV_X1 U6745 ( .A(n5606), .ZN(n5607) );
  AOI21_X1 U6746 ( .B1(n5608), .B2(n5622), .A(n5607), .ZN(n5844) );
  INV_X1 U6747 ( .A(n5844), .ZN(n5719) );
  OR2_X1 U6748 ( .A1(n5609), .A2(n5610), .ZN(n5611) );
  NAND2_X1 U6749 ( .A1(n5678), .A2(n5611), .ZN(n6058) );
  INV_X1 U6750 ( .A(n6058), .ZN(n5617) );
  AOI21_X1 U6751 ( .B1(n5842), .B2(n6193), .A(n6178), .ZN(n5612) );
  OAI21_X1 U6752 ( .B1(n3927), .B2(n6176), .A(n5612), .ZN(n5616) );
  AOI22_X1 U6753 ( .A1(EBX_REG_15__SCAN_IN), .A2(n6191), .B1(
        REIP_REG_15__SCAN_IN), .B2(n5613), .ZN(n5614) );
  OAI21_X1 U6754 ( .B1(REIP_REG_15__SCAN_IN), .B2(n6113), .A(n5614), .ZN(n5615) );
  AOI211_X1 U6755 ( .C1(n5617), .C2(n6153), .A(n5616), .B(n5615), .ZN(n5618)
         );
  OAI21_X1 U6756 ( .B1(n5719), .B2(n6157), .A(n5618), .ZN(U2812) );
  INV_X1 U6757 ( .A(n5619), .ZN(n5621) );
  NOR2_X1 U6758 ( .A1(n5621), .A2(n5620), .ZN(n5624) );
  INV_X1 U6759 ( .A(n5622), .ZN(n5623) );
  AOI21_X1 U6760 ( .B1(n5624), .B2(n5271), .A(n5623), .ZN(n5855) );
  INV_X1 U6761 ( .A(n5855), .ZN(n5722) );
  NOR2_X1 U6762 ( .A1(n5626), .A2(n5625), .ZN(n5627) );
  OR2_X1 U6763 ( .A1(n5609), .A2(n5627), .ZN(n6068) );
  INV_X1 U6764 ( .A(n6068), .ZN(n5635) );
  OAI21_X1 U6765 ( .B1(n5629), .B2(n5631), .A(n5628), .ZN(n6134) );
  OAI22_X1 U6766 ( .A1(n6134), .A2(n6687), .B1(n5853), .B2(n6186), .ZN(n5634)
         );
  AOI22_X1 U6767 ( .A1(EBX_REG_14__SCAN_IN), .A2(n6191), .B1(
        PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n6194), .ZN(n5630) );
  OAI211_X1 U6768 ( .C1(n5632), .C2(n5631), .A(n5630), .B(n6165), .ZN(n5633)
         );
  AOI211_X1 U6769 ( .C1(n5635), .C2(n6153), .A(n5634), .B(n5633), .ZN(n5636)
         );
  OAI21_X1 U6770 ( .B1(n5722), .B2(n6157), .A(n5636), .ZN(U2813) );
  INV_X1 U6771 ( .A(n5865), .ZN(n5638) );
  OAI22_X1 U6772 ( .A1(n5638), .A2(n5689), .B1(n6023), .B2(n5637), .ZN(U2828)
         );
  INV_X1 U6773 ( .A(EBX_REG_29__SCAN_IN), .ZN(n5639) );
  OAI222_X1 U6774 ( .A1(n5688), .A2(n5704), .B1(n5639), .B2(n6023), .C1(n5868), 
        .C2(n5689), .ZN(U2830) );
  INV_X1 U6775 ( .A(EBX_REG_28__SCAN_IN), .ZN(n5641) );
  OAI222_X1 U6776 ( .A1(n5688), .A2(n5747), .B1(n5641), .B2(n6023), .C1(n5640), 
        .C2(n5689), .ZN(U2831) );
  INV_X1 U6777 ( .A(EBX_REG_27__SCAN_IN), .ZN(n5642) );
  OAI222_X1 U6778 ( .A1(n5688), .A2(n5709), .B1(n5642), .B2(n6023), .C1(n5889), 
        .C2(n5689), .ZN(U2832) );
  INV_X1 U6779 ( .A(n5900), .ZN(n5643) );
  AOI22_X1 U6780 ( .A1(n5643), .A2(n6018), .B1(EBX_REG_26__SCAN_IN), .B2(n5668), .ZN(n5644) );
  OAI21_X1 U6781 ( .B1(n5766), .B2(n5691), .A(n5644), .ZN(U2833) );
  INV_X1 U6782 ( .A(EBX_REG_25__SCAN_IN), .ZN(n5646) );
  OAI222_X1 U6783 ( .A1(n5778), .A2(n5691), .B1(n5646), .B2(n6023), .C1(n5645), 
        .C2(n5689), .ZN(U2834) );
  OAI222_X1 U6784 ( .A1(n5688), .A2(n5784), .B1(n6023), .B2(n5563), .C1(n5647), 
        .C2(n5689), .ZN(U2835) );
  INV_X1 U6785 ( .A(EBX_REG_22__SCAN_IN), .ZN(n5648) );
  OAI222_X1 U6786 ( .A1(n5688), .A2(n5805), .B1(n6023), .B2(n5648), .C1(n5936), 
        .C2(n5689), .ZN(U2837) );
  NAND2_X1 U6787 ( .A1(n5650), .A2(n5649), .ZN(n5659) );
  AND2_X1 U6788 ( .A1(n5659), .A2(n5651), .ZN(n5653) );
  INV_X1 U6789 ( .A(EBX_REG_21__SCAN_IN), .ZN(n5658) );
  NAND2_X1 U6790 ( .A1(n5655), .A2(n5654), .ZN(n5656) );
  NAND2_X1 U6791 ( .A1(n5657), .A2(n5656), .ZN(n6004) );
  OAI222_X1 U6792 ( .A1(n6028), .A2(n5691), .B1(n5658), .B2(n6023), .C1(n5689), 
        .C2(n6004), .ZN(U2838) );
  INV_X1 U6793 ( .A(n5659), .ZN(n5660) );
  INV_X1 U6794 ( .A(n6032), .ZN(n5670) );
  MUX2_X1 U6795 ( .A(n5665), .B(n5664), .S(n5663), .Z(n5667) );
  XNOR2_X1 U6796 ( .A(n5667), .B(n5666), .ZN(n6010) );
  AOI22_X1 U6797 ( .A1(n6010), .A2(n6018), .B1(EBX_REG_20__SCAN_IN), .B2(n5668), .ZN(n5669) );
  OAI21_X1 U6798 ( .B1(n5670), .B2(n5691), .A(n5669), .ZN(U2839) );
  INV_X1 U6799 ( .A(n5671), .ZN(n5972) );
  OAI222_X1 U6800 ( .A1(n5972), .A2(n5689), .B1(n6023), .B2(n5592), .C1(n5837), 
        .C2(n5688), .ZN(U2841) );
  NAND2_X1 U6801 ( .A1(n5673), .A2(n5672), .ZN(n5674) );
  NAND2_X1 U6802 ( .A1(n5675), .A2(n5674), .ZN(n6044) );
  OAI21_X1 U6803 ( .B1(n5678), .B2(n5677), .A(n5676), .ZN(n5680) );
  NAND2_X1 U6804 ( .A1(n5680), .A2(n5679), .ZN(n6116) );
  INV_X1 U6805 ( .A(EBX_REG_17__SCAN_IN), .ZN(n6120) );
  OAI22_X1 U6806 ( .A1(n6116), .A2(n5689), .B1(n6120), .B2(n6023), .ZN(n5681)
         );
  AOI21_X1 U6807 ( .B1(n6207), .B2(n6020), .A(n5681), .ZN(n5682) );
  INV_X1 U6808 ( .A(n5682), .ZN(U2842) );
  INV_X1 U6809 ( .A(EBX_REG_16__SCAN_IN), .ZN(n5685) );
  INV_X1 U6810 ( .A(n5683), .ZN(n5684) );
  OAI222_X1 U6811 ( .A1(n5686), .A2(n5691), .B1(n6023), .B2(n5685), .C1(n5689), 
        .C2(n5684), .ZN(U2843) );
  OAI222_X1 U6812 ( .A1(n5719), .A2(n5688), .B1(n5687), .B2(n6023), .C1(n5689), 
        .C2(n6058), .ZN(U2844) );
  INV_X1 U6813 ( .A(EBX_REG_14__SCAN_IN), .ZN(n5690) );
  OAI222_X1 U6814 ( .A1(n5722), .A2(n5691), .B1(n6023), .B2(n5690), .C1(n6068), 
        .C2(n5689), .ZN(U2845) );
  NAND3_X1 U6815 ( .A1(n5730), .A2(n5692), .A3(n5698), .ZN(n5695) );
  NOR2_X2 U6816 ( .A1(n6213), .A2(n5693), .ZN(n6210) );
  AOI22_X1 U6817 ( .A1(n6210), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n6213), .ZN(n5694) );
  NAND2_X1 U6818 ( .A1(n5695), .A2(n5694), .ZN(U2860) );
  AOI22_X1 U6819 ( .A1(n6210), .A2(DATAI_30_), .B1(EAX_REG_30__SCAN_IN), .B2(
        n6213), .ZN(n5700) );
  AND2_X1 U6820 ( .A1(n3470), .A2(n5696), .ZN(n5697) );
  NAND2_X1 U6821 ( .A1(n6214), .A2(DATAI_14_), .ZN(n5699) );
  OAI211_X1 U6822 ( .C1(n5701), .C2(n6024), .A(n5700), .B(n5699), .ZN(U2861)
         );
  AOI22_X1 U6823 ( .A1(n6210), .A2(DATAI_29_), .B1(EAX_REG_29__SCAN_IN), .B2(
        n6213), .ZN(n5703) );
  NAND2_X1 U6824 ( .A1(n6214), .A2(DATAI_13_), .ZN(n5702) );
  OAI211_X1 U6825 ( .C1(n5704), .C2(n6024), .A(n5703), .B(n5702), .ZN(U2862)
         );
  AOI22_X1 U6826 ( .A1(n6210), .A2(DATAI_28_), .B1(EAX_REG_28__SCAN_IN), .B2(
        n6213), .ZN(n5706) );
  NAND2_X1 U6827 ( .A1(n6214), .A2(DATAI_12_), .ZN(n5705) );
  OAI211_X1 U6828 ( .C1(n5747), .C2(n6024), .A(n5706), .B(n5705), .ZN(U2863)
         );
  AOI22_X1 U6829 ( .A1(n6210), .A2(DATAI_27_), .B1(EAX_REG_27__SCAN_IN), .B2(
        n6213), .ZN(n5708) );
  NAND2_X1 U6830 ( .A1(n6214), .A2(DATAI_11_), .ZN(n5707) );
  OAI211_X1 U6831 ( .C1(n5709), .C2(n6024), .A(n5708), .B(n5707), .ZN(U2864)
         );
  AOI22_X1 U6832 ( .A1(n6210), .A2(DATAI_26_), .B1(EAX_REG_26__SCAN_IN), .B2(
        n6213), .ZN(n5711) );
  NAND2_X1 U6833 ( .A1(n6214), .A2(DATAI_10_), .ZN(n5710) );
  OAI211_X1 U6834 ( .C1(n5766), .C2(n6024), .A(n5711), .B(n5710), .ZN(U2865)
         );
  AOI22_X1 U6835 ( .A1(n6210), .A2(DATAI_25_), .B1(EAX_REG_25__SCAN_IN), .B2(
        n6213), .ZN(n5713) );
  NAND2_X1 U6836 ( .A1(n6214), .A2(DATAI_9_), .ZN(n5712) );
  OAI211_X1 U6837 ( .C1(n5778), .C2(n6024), .A(n5713), .B(n5712), .ZN(U2866)
         );
  AOI22_X1 U6838 ( .A1(n6210), .A2(DATAI_24_), .B1(EAX_REG_24__SCAN_IN), .B2(
        n6213), .ZN(n5715) );
  NAND2_X1 U6839 ( .A1(n6214), .A2(DATAI_8_), .ZN(n5714) );
  OAI211_X1 U6840 ( .C1(n5784), .C2(n6024), .A(n5715), .B(n5714), .ZN(U2867)
         );
  AOI22_X1 U6841 ( .A1(n6210), .A2(DATAI_22_), .B1(EAX_REG_22__SCAN_IN), .B2(
        n6213), .ZN(n5717) );
  NAND2_X1 U6842 ( .A1(n6214), .A2(DATAI_6_), .ZN(n5716) );
  OAI211_X1 U6843 ( .C1(n5805), .C2(n6024), .A(n5717), .B(n5716), .ZN(U2869)
         );
  AOI22_X1 U6844 ( .A1(n5720), .A2(DATAI_15_), .B1(n6213), .B2(
        EAX_REG_15__SCAN_IN), .ZN(n5718) );
  OAI21_X1 U6845 ( .B1(n5719), .B2(n6024), .A(n5718), .ZN(U2876) );
  AOI22_X1 U6846 ( .A1(n5720), .A2(DATAI_14_), .B1(n6213), .B2(
        EAX_REG_14__SCAN_IN), .ZN(n5721) );
  OAI21_X1 U6847 ( .B1(n5722), .B2(n6024), .A(n5721), .ZN(U2877) );
  NOR3_X1 U6848 ( .A1(n5773), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(n5723), 
        .ZN(n5724) );
  AOI21_X1 U6849 ( .B1(n5725), .B2(INSTADDRPOINTER_REG_30__SCAN_IN), .A(n5724), 
        .ZN(n5726) );
  XNOR2_X1 U6850 ( .A(n5726), .B(n5857), .ZN(n5867) );
  NAND2_X1 U6851 ( .A1(n6422), .A2(REIP_REG_31__SCAN_IN), .ZN(n5861) );
  NAND2_X1 U6852 ( .A1(n6350), .A2(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5727)
         );
  OAI211_X1 U6853 ( .C1(n6360), .C2(n5728), .A(n5861), .B(n5727), .ZN(n5729)
         );
  OAI21_X1 U6854 ( .B1(n5867), .B2(n6096), .A(n5731), .ZN(U2955) );
  NAND2_X1 U6855 ( .A1(n5741), .A2(n5732), .ZN(n5733) );
  NAND2_X1 U6856 ( .A1(n5734), .A2(n5733), .ZN(n5735) );
  XNOR2_X1 U6857 ( .A(n5735), .B(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5877)
         );
  NAND2_X1 U6858 ( .A1(n6422), .A2(REIP_REG_29__SCAN_IN), .ZN(n5869) );
  NAND2_X1 U6859 ( .A1(n6350), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5736)
         );
  OAI211_X1 U6860 ( .C1(n6360), .C2(n5737), .A(n5869), .B(n5736), .ZN(n5738)
         );
  AOI21_X1 U6861 ( .B1(n5739), .B2(n6354), .A(n5738), .ZN(n5740) );
  OAI21_X1 U6862 ( .B1(n5877), .B2(n6096), .A(n5740), .ZN(U2957) );
  INV_X1 U6863 ( .A(n5741), .ZN(n5764) );
  NAND3_X1 U6864 ( .A1(n5764), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .A3(n5849), .ZN(n5744) );
  INV_X1 U6865 ( .A(n5762), .ZN(n5742) );
  NAND3_X1 U6866 ( .A1(n5775), .A2(n5742), .A3(n5907), .ZN(n5752) );
  AOI22_X1 U6867 ( .A1(n5744), .A2(n5752), .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n5743), .ZN(n5745) );
  XNOR2_X1 U6868 ( .A(n5745), .B(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5886)
         );
  NAND2_X1 U6869 ( .A1(n6422), .A2(REIP_REG_28__SCAN_IN), .ZN(n5878) );
  OAI21_X1 U6870 ( .B1(n6047), .B2(n5746), .A(n5878), .ZN(n5749) );
  NOR2_X1 U6871 ( .A1(n5747), .A2(n6043), .ZN(n5748) );
  AOI211_X1 U6872 ( .C1(n5843), .C2(n5750), .A(n5749), .B(n5748), .ZN(n5751)
         );
  OAI21_X1 U6873 ( .B1(n6096), .B2(n5886), .A(n5751), .ZN(U2958) );
  INV_X1 U6874 ( .A(n5752), .ZN(n5753) );
  NOR2_X1 U6875 ( .A1(n5754), .A2(n5753), .ZN(n5755) );
  XNOR2_X1 U6876 ( .A(n5755), .B(n5892), .ZN(n5895) );
  NAND2_X1 U6877 ( .A1(n6422), .A2(REIP_REG_27__SCAN_IN), .ZN(n5887) );
  NAND2_X1 U6878 ( .A1(n6350), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5756)
         );
  OAI211_X1 U6879 ( .C1(n6360), .C2(n5757), .A(n5887), .B(n5756), .ZN(n5758)
         );
  AOI21_X1 U6880 ( .B1(n5759), .B2(n6354), .A(n5758), .ZN(n5760) );
  OAI21_X1 U6881 ( .B1(n5895), .B2(n6096), .A(n5760), .ZN(U2959) );
  NAND2_X1 U6882 ( .A1(n5762), .A2(n5761), .ZN(n5763) );
  XNOR2_X1 U6883 ( .A(n5764), .B(n5763), .ZN(n5904) );
  NAND2_X1 U6884 ( .A1(n6422), .A2(REIP_REG_26__SCAN_IN), .ZN(n5896) );
  OAI21_X1 U6885 ( .B1(n6047), .B2(n5765), .A(n5896), .ZN(n5768) );
  NOR2_X1 U6886 ( .A1(n5766), .A2(n6043), .ZN(n5767) );
  AOI211_X1 U6887 ( .C1(n5843), .C2(n5769), .A(n5768), .B(n5767), .ZN(n5770)
         );
  OAI21_X1 U6888 ( .B1(n5904), .B2(n6096), .A(n5770), .ZN(U2960) );
  AND2_X1 U6889 ( .A1(n6422), .A2(REIP_REG_25__SCAN_IN), .ZN(n5909) );
  NOR2_X1 U6890 ( .A1(n6360), .A2(n5771), .ZN(n5772) );
  AOI211_X1 U6891 ( .C1(n6350), .C2(PHYADDRPOINTER_REG_25__SCAN_IN), .A(n5909), 
        .B(n5772), .ZN(n5777) );
  OAI21_X1 U6892 ( .B1(n5775), .B2(n5774), .A(n5773), .ZN(n5906) );
  NAND2_X1 U6893 ( .A1(n5906), .A2(n6356), .ZN(n5776) );
  OAI211_X1 U6894 ( .C1(n5778), .C2(n6043), .A(n5777), .B(n5776), .ZN(U2961)
         );
  OAI21_X1 U6895 ( .B1(n5794), .B2(n5961), .A(n5849), .ZN(n5779) );
  XNOR2_X1 U6896 ( .A(n5849), .B(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5816)
         );
  NOR2_X1 U6897 ( .A1(n5849), .A2(n5955), .ZN(n5780) );
  XNOR2_X1 U6898 ( .A(n5849), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5812)
         );
  NOR2_X1 U6899 ( .A1(n5849), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5801)
         );
  NAND2_X1 U6900 ( .A1(n5781), .A2(n5801), .ZN(n5792) );
  NAND3_X1 U6901 ( .A1(n5849), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5782) );
  OAI22_X1 U6902 ( .A1(n5792), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .B1(n5803), .B2(n5782), .ZN(n5783) );
  XNOR2_X1 U6903 ( .A(n5783), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5920)
         );
  INV_X1 U6904 ( .A(n5784), .ZN(n5789) );
  INV_X1 U6905 ( .A(n5785), .ZN(n5787) );
  AND2_X1 U6906 ( .A1(n6422), .A2(REIP_REG_24__SCAN_IN), .ZN(n5917) );
  AOI21_X1 U6907 ( .B1(n6350), .B2(PHYADDRPOINTER_REG_24__SCAN_IN), .A(n5917), 
        .ZN(n5786) );
  OAI21_X1 U6908 ( .B1(n5787), .B2(n6360), .A(n5786), .ZN(n5788) );
  AOI21_X1 U6909 ( .B1(n5789), .B2(n6354), .A(n5788), .ZN(n5790) );
  OAI21_X1 U6910 ( .B1(n5920), .B2(n6096), .A(n5790), .ZN(U2962) );
  NAND3_X1 U6911 ( .A1(n5849), .A2(n5791), .A3(n5954), .ZN(n5793) );
  OAI21_X1 U6912 ( .B1(n5794), .B2(n5793), .A(n5792), .ZN(n5795) );
  XNOR2_X1 U6913 ( .A(n5795), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5932)
         );
  AOI21_X1 U6914 ( .B1(n5797), .B2(n5569), .A(n5796), .ZN(n6025) );
  NAND2_X1 U6915 ( .A1(n6422), .A2(REIP_REG_23__SCAN_IN), .ZN(n5927) );
  NAND2_X1 U6916 ( .A1(n6350), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5798)
         );
  OAI211_X1 U6917 ( .C1(n6360), .C2(n5996), .A(n5927), .B(n5798), .ZN(n5799)
         );
  AOI21_X1 U6918 ( .B1(n6025), .B2(n6354), .A(n5799), .ZN(n5800) );
  OAI21_X1 U6919 ( .B1(n5932), .B2(n6096), .A(n5800), .ZN(U2963) );
  AOI21_X1 U6920 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n5849), .A(n5801), 
        .ZN(n5802) );
  XNOR2_X1 U6921 ( .A(n5803), .B(n5802), .ZN(n5941) );
  INV_X1 U6922 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5804) );
  NAND2_X1 U6923 ( .A1(n6422), .A2(REIP_REG_22__SCAN_IN), .ZN(n5935) );
  OAI21_X1 U6924 ( .B1(n6047), .B2(n5804), .A(n5935), .ZN(n5807) );
  NOR2_X1 U6925 ( .A1(n5805), .A2(n6043), .ZN(n5806) );
  AOI211_X1 U6926 ( .C1(n5843), .C2(n5808), .A(n5807), .B(n5806), .ZN(n5809)
         );
  OAI21_X1 U6927 ( .B1(n5941), .B2(n6096), .A(n5809), .ZN(U2964) );
  OAI21_X1 U6928 ( .B1(n5812), .B2(n5811), .A(n5810), .ZN(n5942) );
  NAND2_X1 U6929 ( .A1(n5942), .A2(n6356), .ZN(n5815) );
  NOR2_X1 U6930 ( .A1(n6407), .A2(n6693), .ZN(n5944) );
  NOR2_X1 U6931 ( .A1(n6360), .A2(n6009), .ZN(n5813) );
  AOI211_X1 U6932 ( .C1(n6350), .C2(PHYADDRPOINTER_REG_21__SCAN_IN), .A(n5944), 
        .B(n5813), .ZN(n5814) );
  OAI211_X1 U6933 ( .C1(n6043), .C2(n6028), .A(n5815), .B(n5814), .ZN(U2965)
         );
  XNOR2_X1 U6934 ( .A(n5817), .B(n5816), .ZN(n5959) );
  NAND2_X1 U6935 ( .A1(n5843), .A2(n6013), .ZN(n5818) );
  NAND2_X1 U6936 ( .A1(n6422), .A2(REIP_REG_20__SCAN_IN), .ZN(n5953) );
  OAI211_X1 U6937 ( .C1(n6047), .C2(n5819), .A(n5818), .B(n5953), .ZN(n5820)
         );
  AOI21_X1 U6938 ( .B1(n6032), .B2(n6354), .A(n5820), .ZN(n5821) );
  OAI21_X1 U6939 ( .B1(n5959), .B2(n6096), .A(n5821), .ZN(U2966) );
  OAI21_X1 U6940 ( .B1(n3156), .B2(n5961), .A(n5823), .ZN(n5824) );
  XNOR2_X1 U6941 ( .A(n5824), .B(n5277), .ZN(n5960) );
  NAND2_X1 U6942 ( .A1(n5960), .A2(n6356), .ZN(n5828) );
  AND2_X1 U6943 ( .A1(n6422), .A2(REIP_REG_19__SCAN_IN), .ZN(n5964) );
  NOR2_X1 U6944 ( .A1(n6360), .A2(n5825), .ZN(n5826) );
  AOI211_X1 U6945 ( .C1(n6350), .C2(PHYADDRPOINTER_REG_19__SCAN_IN), .A(n5964), 
        .B(n5826), .ZN(n5827) );
  OAI211_X1 U6946 ( .C1(n6043), .C2(n6035), .A(n5828), .B(n5827), .ZN(U2967)
         );
  INV_X1 U6947 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5833) );
  NAND2_X1 U6948 ( .A1(n6422), .A2(REIP_REG_18__SCAN_IN), .ZN(n5971) );
  NAND2_X1 U6949 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n6041), .ZN(n5830) );
  NAND3_X1 U6950 ( .A1(n6040), .A2(n6055), .A3(n6039), .ZN(n5829) );
  OAI21_X1 U6951 ( .B1(n5830), .B2(n6039), .A(n5829), .ZN(n5831) );
  XOR2_X1 U6952 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .B(n5831), .Z(n5969) );
  NAND2_X1 U6953 ( .A1(n6356), .A2(n5969), .ZN(n5832) );
  OAI211_X1 U6954 ( .C1(n6047), .C2(n5833), .A(n5971), .B(n5832), .ZN(n5834)
         );
  AOI21_X1 U6955 ( .B1(n5843), .B2(n5835), .A(n5834), .ZN(n5836) );
  OAI21_X1 U6956 ( .B1(n5837), .B2(n6043), .A(n5836), .ZN(U2968) );
  XNOR2_X1 U6957 ( .A(n5849), .B(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5838)
         );
  XNOR2_X1 U6958 ( .A(n5839), .B(n5838), .ZN(n6059) );
  INV_X1 U6959 ( .A(REIP_REG_15__SCAN_IN), .ZN(n5840) );
  OAI22_X1 U6960 ( .A1(n6047), .A2(n3927), .B1(n6407), .B2(n5840), .ZN(n5841)
         );
  AOI21_X1 U6961 ( .B1(n5843), .B2(n5842), .A(n5841), .ZN(n5846) );
  NAND2_X1 U6962 ( .A1(n5844), .A2(n6354), .ZN(n5845) );
  OAI211_X1 U6963 ( .C1(n6059), .C2(n6096), .A(n5846), .B(n5845), .ZN(U2971)
         );
  XNOR2_X1 U6964 ( .A(n5849), .B(n5848), .ZN(n5850) );
  XNOR2_X1 U6965 ( .A(n5851), .B(n5850), .ZN(n6067) );
  AOI22_X1 U6966 ( .A1(n6350), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .B1(n6422), 
        .B2(REIP_REG_14__SCAN_IN), .ZN(n5852) );
  OAI21_X1 U6967 ( .B1(n5853), .B2(n6360), .A(n5852), .ZN(n5854) );
  AOI21_X1 U6968 ( .B1(n5855), .B2(n6354), .A(n5854), .ZN(n5856) );
  OAI21_X1 U6969 ( .B1(n6067), .B2(n6096), .A(n5856), .ZN(U2972) );
  NAND2_X1 U6970 ( .A1(n5857), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5862) );
  NAND3_X1 U6971 ( .A1(n5859), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .A3(n5858), .ZN(n5860) );
  OAI211_X1 U6972 ( .C1(n5863), .C2(n5862), .A(n5861), .B(n5860), .ZN(n5864)
         );
  AOI21_X1 U6973 ( .B1(n5865), .B2(n6424), .A(n5864), .ZN(n5866) );
  OAI21_X1 U6974 ( .B1(n5867), .B2(n6403), .A(n5866), .ZN(U2987) );
  INV_X1 U6975 ( .A(n5868), .ZN(n5872) );
  OAI21_X1 U6976 ( .B1(n5870), .B2(n5873), .A(n5869), .ZN(n5871) );
  AOI21_X1 U6977 ( .B1(n5872), .B2(n6424), .A(n5871), .ZN(n5876) );
  NAND3_X1 U6978 ( .A1(n5893), .A2(n5874), .A3(n5873), .ZN(n5875) );
  OAI211_X1 U6979 ( .C1(n5877), .C2(n6403), .A(n5876), .B(n5875), .ZN(U2989)
         );
  OAI21_X1 U6980 ( .B1(n5888), .B2(n5879), .A(n5878), .ZN(n5880) );
  AOI21_X1 U6981 ( .B1(n5881), .B2(n6424), .A(n5880), .ZN(n5885) );
  NAND3_X1 U6982 ( .A1(n5893), .A2(n5883), .A3(n5882), .ZN(n5884) );
  OAI211_X1 U6983 ( .C1(n5886), .C2(n6403), .A(n5885), .B(n5884), .ZN(U2990)
         );
  OAI21_X1 U6984 ( .B1(n5888), .B2(n5892), .A(n5887), .ZN(n5891) );
  NOR2_X1 U6985 ( .A1(n5889), .A2(n6391), .ZN(n5890) );
  AOI211_X1 U6986 ( .C1(n5893), .C2(n5892), .A(n5891), .B(n5890), .ZN(n5894)
         );
  OAI21_X1 U6987 ( .B1(n5895), .B2(n6403), .A(n5894), .ZN(U2991) );
  XNOR2_X1 U6988 ( .A(n5907), .B(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5902)
         );
  INV_X1 U6989 ( .A(n5896), .ZN(n5897) );
  AOI21_X1 U6990 ( .B1(n5898), .B2(INSTADDRPOINTER_REG_26__SCAN_IN), .A(n5897), 
        .ZN(n5899) );
  OAI21_X1 U6991 ( .B1(n5900), .B2(n6391), .A(n5899), .ZN(n5901) );
  AOI21_X1 U6992 ( .B1(n5905), .B2(n5902), .A(n5901), .ZN(n5903) );
  OAI21_X1 U6993 ( .B1(n5904), .B2(n6403), .A(n5903), .ZN(U2992) );
  INV_X1 U6994 ( .A(n5905), .ZN(n5913) );
  NAND2_X1 U6995 ( .A1(n5906), .A2(n6429), .ZN(n5912) );
  NOR2_X1 U6996 ( .A1(n5914), .A2(n5907), .ZN(n5908) );
  AOI211_X1 U6997 ( .C1(n5910), .C2(n6424), .A(n5909), .B(n5908), .ZN(n5911)
         );
  OAI211_X1 U6998 ( .C1(INSTADDRPOINTER_REG_25__SCAN_IN), .C2(n5913), .A(n5912), .B(n5911), .ZN(U2993) );
  AOI21_X1 U6999 ( .B1(n5930), .B2(INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5915) );
  NOR2_X1 U7000 ( .A1(n5915), .A2(n5914), .ZN(n5916) );
  AOI211_X1 U7001 ( .C1(n6424), .C2(n5918), .A(n5917), .B(n5916), .ZN(n5919)
         );
  OAI21_X1 U7002 ( .B1(n5920), .B2(n6403), .A(n5919), .ZN(U2994) );
  INV_X1 U7003 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5929) );
  INV_X1 U7004 ( .A(n5921), .ZN(n5922) );
  OAI21_X1 U7005 ( .B1(n5924), .B2(n5923), .A(n5922), .ZN(n5999) );
  NAND2_X1 U7006 ( .A1(n5925), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5926) );
  OAI211_X1 U7007 ( .C1(n5999), .C2(n6391), .A(n5927), .B(n5926), .ZN(n5928)
         );
  AOI21_X1 U7008 ( .B1(n5930), .B2(n5929), .A(n5928), .ZN(n5931) );
  OAI21_X1 U7009 ( .B1(n5932), .B2(n6403), .A(n5931), .ZN(U2995) );
  INV_X1 U7010 ( .A(n5948), .ZN(n5939) );
  XNOR2_X1 U7011 ( .A(n5933), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5938)
         );
  NAND2_X1 U7012 ( .A1(n5945), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5934) );
  OAI211_X1 U7013 ( .C1(n5936), .C2(n6391), .A(n5935), .B(n5934), .ZN(n5937)
         );
  AOI21_X1 U7014 ( .B1(n5939), .B2(n5938), .A(n5937), .ZN(n5940) );
  OAI21_X1 U7015 ( .B1(n5941), .B2(n6403), .A(n5940), .ZN(U2996) );
  NAND2_X1 U7016 ( .A1(n5942), .A2(n6429), .ZN(n5947) );
  NOR2_X1 U7017 ( .A1(n6004), .A2(n6391), .ZN(n5943) );
  AOI211_X1 U7018 ( .C1(INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n5945), .A(n5944), .B(n5943), .ZN(n5946) );
  OAI211_X1 U7019 ( .C1(INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n5948), .A(n5947), .B(n5946), .ZN(U2997) );
  INV_X1 U7020 ( .A(n5949), .ZN(n5950) );
  OAI21_X1 U7021 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n5950), .A(n6056), 
        .ZN(n5974) );
  AOI21_X1 U7022 ( .B1(n5952), .B2(n5951), .A(n5974), .ZN(n5962) );
  OAI21_X1 U7023 ( .B1(n5962), .B2(n5955), .A(n5953), .ZN(n5957) );
  AOI211_X1 U7024 ( .C1(n5961), .C2(n5955), .A(n5954), .B(n5968), .ZN(n5956)
         );
  AOI211_X1 U7025 ( .C1(n6424), .C2(n6010), .A(n5957), .B(n5956), .ZN(n5958)
         );
  OAI21_X1 U7026 ( .B1(n5959), .B2(n6403), .A(n5958), .ZN(U2998) );
  NAND2_X1 U7027 ( .A1(n5960), .A2(n6429), .ZN(n5967) );
  NOR2_X1 U7028 ( .A1(n5962), .A2(n5961), .ZN(n5963) );
  AOI211_X1 U7029 ( .C1(n6424), .C2(n5965), .A(n5964), .B(n5963), .ZN(n5966)
         );
  OAI211_X1 U7030 ( .C1(INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n5968), .A(n5967), .B(n5966), .ZN(U2999) );
  NAND2_X1 U7031 ( .A1(n6429), .A2(n5969), .ZN(n5970) );
  OAI211_X1 U7032 ( .C1(n5972), .C2(n6391), .A(n5971), .B(n5970), .ZN(n5973)
         );
  AOI21_X1 U7033 ( .B1(INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n5974), .A(n5973), 
        .ZN(n5977) );
  NOR2_X1 U7034 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n6055), .ZN(n5975)
         );
  NAND2_X1 U7035 ( .A1(n6052), .A2(n5975), .ZN(n5976) );
  NAND2_X1 U7036 ( .A1(n5977), .A2(n5976), .ZN(U3000) );
  INV_X1 U7037 ( .A(n6438), .ZN(n6531) );
  OAI211_X1 U7038 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n5978), .A(n6531), .B(
        n6530), .ZN(n5979) );
  OAI21_X1 U7039 ( .B1(n5988), .B2(n4349), .A(n5979), .ZN(n5980) );
  MUX2_X1 U7040 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n5980), .S(n6434), 
        .Z(U3464) );
  XNOR2_X1 U7041 ( .A(n5981), .B(n6438), .ZN(n5983) );
  OAI22_X1 U7042 ( .A1(n5983), .A2(n6537), .B1(n5982), .B2(n5988), .ZN(n5984)
         );
  MUX2_X1 U7043 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n5984), .S(n6434), 
        .Z(U3463) );
  INV_X1 U7044 ( .A(n4424), .ZN(n5990) );
  NAND2_X1 U7045 ( .A1(n5985), .A2(n6532), .ZN(n6441) );
  NOR2_X1 U7046 ( .A1(n5986), .A2(n6531), .ZN(n6488) );
  NOR2_X1 U7047 ( .A1(n6441), .A2(n6488), .ZN(n5989) );
  OAI222_X1 U7048 ( .A1(n5991), .A2(n5990), .B1(n6537), .B2(n5989), .C1(n5988), 
        .C2(n5987), .ZN(n5992) );
  MUX2_X1 U7049 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n5992), .S(n6434), 
        .Z(U3462) );
  INV_X1 U7050 ( .A(MEMORYFETCH_REG_SCAN_IN), .ZN(n7054) );
  OAI21_X1 U7051 ( .B1(n5994), .B2(n7054), .A(n5993), .ZN(U2788) );
  AOI21_X1 U7052 ( .B1(REIP_REG_22__SCAN_IN), .B2(n5995), .A(
        REIP_REG_23__SCAN_IN), .ZN(n6002) );
  INV_X1 U7053 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5997) );
  OAI22_X1 U7054 ( .A1(n5997), .A2(n6176), .B1(n5996), .B2(n6186), .ZN(n5998)
         );
  AOI21_X1 U7055 ( .B1(EBX_REG_23__SCAN_IN), .B2(n6191), .A(n5998), .ZN(n6001)
         );
  INV_X1 U7056 ( .A(n5999), .ZN(n6019) );
  AOI22_X1 U7057 ( .A1(n6025), .A2(n6171), .B1(n6019), .B2(n6153), .ZN(n6000)
         );
  OAI211_X1 U7058 ( .C1(n6003), .C2(n6002), .A(n6001), .B(n6000), .ZN(U2804)
         );
  AOI22_X1 U7059 ( .A1(EBX_REG_21__SCAN_IN), .A2(n6191), .B1(
        PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n6194), .ZN(n6008) );
  OAI22_X1 U7060 ( .A1(n6028), .A2(n6157), .B1(n6198), .B2(n6004), .ZN(n6005)
         );
  AOI211_X1 U7061 ( .C1(REIP_REG_21__SCAN_IN), .C2(n6011), .A(n6006), .B(n6005), .ZN(n6007) );
  OAI211_X1 U7062 ( .C1(n6009), .C2(n6186), .A(n6008), .B(n6007), .ZN(U2806)
         );
  AOI22_X1 U7063 ( .A1(EBX_REG_20__SCAN_IN), .A2(n6191), .B1(
        PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n6194), .ZN(n6017) );
  AOI22_X1 U7064 ( .A1(n6032), .A2(n6171), .B1(n6153), .B2(n6010), .ZN(n6016)
         );
  OAI221_X1 U7065 ( .B1(REIP_REG_20__SCAN_IN), .B2(n6012), .C1(
        REIP_REG_20__SCAN_IN), .C2(REIP_REG_19__SCAN_IN), .A(n6011), .ZN(n6015) );
  NAND2_X1 U7066 ( .A1(n6013), .A2(n6193), .ZN(n6014) );
  NAND4_X1 U7067 ( .A1(n6017), .A2(n6016), .A3(n6015), .A4(n6014), .ZN(U2807)
         );
  AOI22_X1 U7068 ( .A1(n6025), .A2(n6020), .B1(n6019), .B2(n6018), .ZN(n6021)
         );
  OAI21_X1 U7069 ( .B1(n6023), .B2(n6022), .A(n6021), .ZN(U2836) );
  INV_X1 U7070 ( .A(n6024), .ZN(n6211) );
  AOI22_X1 U7071 ( .A1(n6025), .A2(n6211), .B1(n6210), .B2(DATAI_23_), .ZN(
        n6027) );
  AOI22_X1 U7072 ( .A1(n6214), .A2(DATAI_7_), .B1(n6213), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n6026) );
  NAND2_X1 U7073 ( .A1(n6027), .A2(n6026), .ZN(U2868) );
  INV_X1 U7074 ( .A(n6028), .ZN(n6029) );
  AOI22_X1 U7075 ( .A1(n6029), .A2(n6211), .B1(n6210), .B2(DATAI_21_), .ZN(
        n6031) );
  AOI22_X1 U7076 ( .A1(n6214), .A2(DATAI_5_), .B1(n6213), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n6030) );
  NAND2_X1 U7077 ( .A1(n6031), .A2(n6030), .ZN(U2870) );
  AOI22_X1 U7078 ( .A1(n6032), .A2(n6211), .B1(n6210), .B2(DATAI_20_), .ZN(
        n6034) );
  AOI22_X1 U7079 ( .A1(n6214), .A2(DATAI_4_), .B1(n6213), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n6033) );
  NAND2_X1 U7080 ( .A1(n6034), .A2(n6033), .ZN(U2871) );
  INV_X1 U7081 ( .A(n6035), .ZN(n6036) );
  AOI22_X1 U7082 ( .A1(n6036), .A2(n6211), .B1(n6210), .B2(DATAI_19_), .ZN(
        n6038) );
  AOI22_X1 U7083 ( .A1(n6214), .A2(DATAI_3_), .B1(n6213), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n6037) );
  NAND2_X1 U7084 ( .A1(n6038), .A2(n6037), .ZN(U2872) );
  INV_X1 U7085 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n6048) );
  MUX2_X1 U7086 ( .A(n6041), .B(n6040), .S(n6039), .Z(n6042) );
  XNOR2_X1 U7087 ( .A(n6042), .B(n6055), .ZN(n6049) );
  OAI22_X1 U7088 ( .A1(n6044), .A2(n6043), .B1(n6115), .B2(n6360), .ZN(n6045)
         );
  AOI21_X1 U7089 ( .B1(n6049), .B2(n6356), .A(n6045), .ZN(n6046) );
  NAND2_X1 U7090 ( .A1(n6422), .A2(REIP_REG_17__SCAN_IN), .ZN(n6053) );
  OAI211_X1 U7091 ( .C1(n6048), .C2(n6047), .A(n6046), .B(n6053), .ZN(U2969)
         );
  INV_X1 U7092 ( .A(n6049), .ZN(n6050) );
  OAI22_X1 U7093 ( .A1(n6050), .A2(n6403), .B1(n6391), .B2(n6116), .ZN(n6051)
         );
  AOI21_X1 U7094 ( .B1(n6052), .B2(n6055), .A(n6051), .ZN(n6054) );
  OAI211_X1 U7095 ( .C1(n6056), .C2(n6055), .A(n6054), .B(n6053), .ZN(U3001)
         );
  INV_X1 U7096 ( .A(n6057), .ZN(n6062) );
  OAI22_X1 U7097 ( .A1(n6058), .A2(n6391), .B1(n5840), .B2(n6407), .ZN(n6061)
         );
  NOR2_X1 U7098 ( .A1(n6059), .A2(n6403), .ZN(n6060) );
  AOI211_X1 U7099 ( .C1(n6064), .C2(n6062), .A(n6061), .B(n6060), .ZN(n6063)
         );
  OAI21_X1 U7100 ( .B1(n6065), .B2(n6064), .A(n6063), .ZN(U3003) );
  NAND2_X1 U7101 ( .A1(n6076), .A2(n6066), .ZN(n6081) );
  OAI222_X1 U7102 ( .A1(n6068), .A2(n6391), .B1(n6407), .B2(n6687), .C1(n6403), 
        .C2(n6067), .ZN(n6069) );
  INV_X1 U7103 ( .A(n6069), .ZN(n6080) );
  INV_X1 U7104 ( .A(n6070), .ZN(n6072) );
  AOI21_X1 U7105 ( .B1(n6072), .B2(n6071), .A(INSTADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n6078) );
  INV_X1 U7106 ( .A(n6073), .ZN(n6077) );
  AOI21_X1 U7107 ( .B1(n6074), .B2(n6082), .A(n6364), .ZN(n6075) );
  OAI21_X1 U7108 ( .B1(n6077), .B2(n6076), .A(n6075), .ZN(n6084) );
  OAI21_X1 U7109 ( .B1(n6078), .B2(n6084), .A(INSTADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n6079) );
  OAI211_X1 U7110 ( .C1(INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n6081), .A(n6080), .B(n6079), .ZN(U3004) );
  OR2_X1 U7111 ( .A1(n6082), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n6088)
         );
  AOI21_X1 U7112 ( .B1(n6126), .B2(n6424), .A(n6083), .ZN(n6087) );
  AOI22_X1 U7113 ( .A1(n6085), .A2(n6429), .B1(INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n6084), .ZN(n6086) );
  OAI211_X1 U7114 ( .C1(n6367), .C2(n6088), .A(n6087), .B(n6086), .ZN(U3005)
         );
  INV_X1 U7115 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6673) );
  INV_X1 U7116 ( .A(STATE_REG_0__SCAN_IN), .ZN(n6993) );
  AOI21_X1 U7117 ( .B1(STATE_REG_1__SCAN_IN), .B2(n6673), .A(n6993), .ZN(n6093) );
  INV_X1 U7118 ( .A(ADS_N_REG_SCAN_IN), .ZN(n6089) );
  NAND2_X1 U7119 ( .A1(n6993), .A2(STATE_REG_1__SCAN_IN), .ZN(n7122) );
  INV_X2 U7120 ( .A(n7122), .ZN(n7123) );
  AOI21_X1 U7121 ( .B1(n6093), .B2(n6089), .A(n7123), .ZN(U2789) );
  OAI21_X1 U7122 ( .B1(n6090), .B2(n6648), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n6091) );
  OAI21_X1 U7123 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6647), .A(n6091), .ZN(
        U2790) );
  NOR2_X1 U7124 ( .A1(STATE_REG_0__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n6094) );
  OAI21_X1 U7125 ( .B1(n6094), .B2(D_C_N_REG_SCAN_IN), .A(n7122), .ZN(n6092)
         );
  OAI21_X1 U7126 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n7122), .A(n6092), .ZN(
        U2791) );
  OAI21_X1 U7127 ( .B1(BS16_N), .B2(n6094), .A(n3155), .ZN(n6704) );
  OAI21_X1 U7128 ( .B1(n3155), .B2(n6999), .A(n6704), .ZN(U2792) );
  INV_X1 U7129 ( .A(n6095), .ZN(n6097) );
  OAI21_X1 U7130 ( .B1(n6097), .B2(n7067), .A(n6096), .ZN(U2793) );
  INV_X1 U7131 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n7034) );
  NOR4_X1 U7132 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(DATAWIDTH_REG_8__SCAN_IN), .A3(DATAWIDTH_REG_11__SCAN_IN), .A4(DATAWIDTH_REG_23__SCAN_IN), .ZN(n6107)
         );
  AOI211_X1 U7133 ( .C1(DATAWIDTH_REG_1__SCAN_IN), .C2(
        DATAWIDTH_REG_0__SCAN_IN), .A(DATAWIDTH_REG_17__SCAN_IN), .B(
        DATAWIDTH_REG_7__SCAN_IN), .ZN(n6106) );
  NOR4_X1 U7134 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(DATAWIDTH_REG_13__SCAN_IN), .A3(DATAWIDTH_REG_20__SCAN_IN), .A4(DATAWIDTH_REG_22__SCAN_IN), .ZN(n6098)
         );
  INV_X1 U7135 ( .A(DATAWIDTH_REG_12__SCAN_IN), .ZN(n7060) );
  INV_X1 U7136 ( .A(DATAWIDTH_REG_4__SCAN_IN), .ZN(n7051) );
  NAND3_X1 U7137 ( .A1(n6098), .A2(n7060), .A3(n7051), .ZN(n6104) );
  NOR4_X1 U7138 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(DATAWIDTH_REG_6__SCAN_IN), 
        .A3(DATAWIDTH_REG_10__SCAN_IN), .A4(DATAWIDTH_REG_21__SCAN_IN), .ZN(
        n6102) );
  NOR4_X1 U7139 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(DATAWIDTH_REG_14__SCAN_IN), .A3(DATAWIDTH_REG_15__SCAN_IN), .A4(DATAWIDTH_REG_3__SCAN_IN), .ZN(n6101) );
  NOR4_X1 U7140 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(
        DATAWIDTH_REG_29__SCAN_IN), .A3(DATAWIDTH_REG_30__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n6100) );
  NOR4_X1 U7141 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(
        DATAWIDTH_REG_25__SCAN_IN), .A3(DATAWIDTH_REG_26__SCAN_IN), .A4(
        DATAWIDTH_REG_27__SCAN_IN), .ZN(n6099) );
  NAND4_X1 U7142 ( .A1(n6102), .A2(n6101), .A3(n6100), .A4(n6099), .ZN(n6103)
         );
  NOR4_X1 U7143 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(
        DATAWIDTH_REG_16__SCAN_IN), .A3(n6104), .A4(n6103), .ZN(n6105) );
  NAND3_X1 U7144 ( .A1(n6107), .A2(n6106), .A3(n6105), .ZN(n6716) );
  NOR3_X1 U7145 ( .A1(REIP_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .A3(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6109) );
  INV_X1 U7146 ( .A(n6109), .ZN(n6108) );
  NOR2_X1 U7147 ( .A1(n6716), .A2(REIP_REG_1__SCAN_IN), .ZN(n6714) );
  AOI22_X1 U7148 ( .A1(n7034), .A2(n6716), .B1(n6108), .B2(n6714), .ZN(U2794)
         );
  INV_X1 U7149 ( .A(n6716), .ZN(n6713) );
  INV_X1 U7150 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n7107) );
  AOI21_X1 U7151 ( .B1(n6710), .B2(n7107), .A(n6109), .ZN(n6110) );
  INV_X1 U7152 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n7015) );
  AOI22_X1 U7153 ( .A1(n6713), .A2(n6110), .B1(n7015), .B2(n6716), .ZN(U2795)
         );
  INV_X1 U7154 ( .A(REIP_REG_17__SCAN_IN), .ZN(n7088) );
  AOI221_X1 U7155 ( .B1(n6113), .B2(n7088), .C1(n6112), .C2(n7088), .A(n6111), 
        .ZN(n6114) );
  AOI211_X1 U7156 ( .C1(n6194), .C2(PHYADDRPOINTER_REG_17__SCAN_IN), .A(n6178), 
        .B(n6114), .ZN(n6119) );
  OAI22_X1 U7157 ( .A1(n6116), .A2(n6198), .B1(n6115), .B2(n6186), .ZN(n6117)
         );
  AOI21_X1 U7158 ( .B1(n6207), .B2(n6171), .A(n6117), .ZN(n6118) );
  OAI211_X1 U7159 ( .C1(n6120), .C2(n6123), .A(n6119), .B(n6118), .ZN(U2810)
         );
  NOR3_X1 U7160 ( .A1(n6181), .A2(n6121), .A3(n6684), .ZN(n6141) );
  AOI21_X1 U7161 ( .B1(REIP_REG_12__SCAN_IN), .B2(n6141), .A(
        REIP_REG_13__SCAN_IN), .ZN(n6133) );
  INV_X1 U7162 ( .A(EBX_REG_13__SCAN_IN), .ZN(n6124) );
  AOI21_X1 U7163 ( .B1(n6194), .B2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n6178), 
        .ZN(n6122) );
  OAI21_X1 U7164 ( .B1(n6124), .B2(n6123), .A(n6122), .ZN(n6125) );
  AOI21_X1 U7165 ( .B1(n6126), .B2(n6153), .A(n6125), .ZN(n6132) );
  INV_X1 U7166 ( .A(n6127), .ZN(n6130) );
  INV_X1 U7167 ( .A(n6128), .ZN(n6129) );
  AOI22_X1 U7168 ( .A1(n6130), .A2(n6171), .B1(n6193), .B2(n6129), .ZN(n6131)
         );
  OAI211_X1 U7169 ( .C1(n6134), .C2(n6133), .A(n6132), .B(n6131), .ZN(U2814)
         );
  INV_X1 U7170 ( .A(n6135), .ZN(n6139) );
  OAI21_X1 U7171 ( .B1(n6176), .B2(n6136), .A(n6165), .ZN(n6137) );
  AOI21_X1 U7172 ( .B1(n6191), .B2(EBX_REG_12__SCAN_IN), .A(n6137), .ZN(n6138)
         );
  OAI21_X1 U7173 ( .B1(n6139), .B2(n6198), .A(n6138), .ZN(n6140) );
  AOI221_X1 U7174 ( .B1(n6142), .B2(REIP_REG_12__SCAN_IN), .C1(n6141), .C2(
        n5401), .A(n6140), .ZN(n6148) );
  INV_X1 U7175 ( .A(n6143), .ZN(n6144) );
  OAI22_X1 U7176 ( .A1(n6145), .A2(n6157), .B1(n6186), .B2(n6144), .ZN(n6146)
         );
  INV_X1 U7177 ( .A(n6146), .ZN(n6147) );
  NAND2_X1 U7178 ( .A1(n6148), .A2(n6147), .ZN(U2815) );
  INV_X1 U7179 ( .A(n6149), .ZN(n6154) );
  INV_X1 U7180 ( .A(n6150), .ZN(n6152) );
  INV_X1 U7181 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6682) );
  AOI22_X1 U7182 ( .A1(REIP_REG_10__SCAN_IN), .A2(REIP_REG_9__SCAN_IN), .B1(
        n6683), .B2(n6682), .ZN(n6151) );
  AOI22_X1 U7183 ( .A1(n6154), .A2(n6153), .B1(n6152), .B2(n6151), .ZN(n6163)
         );
  AOI22_X1 U7184 ( .A1(PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n6194), .B1(
        REIP_REG_10__SCAN_IN), .B2(n6155), .ZN(n6162) );
  AOI21_X1 U7185 ( .B1(n6191), .B2(EBX_REG_10__SCAN_IN), .A(n6178), .ZN(n6161)
         );
  OAI22_X1 U7186 ( .A1(n6158), .A2(n6157), .B1(n6186), .B2(n6156), .ZN(n6159)
         );
  INV_X1 U7187 ( .A(n6159), .ZN(n6160) );
  NAND4_X1 U7188 ( .A1(n6163), .A2(n6162), .A3(n6161), .A4(n6160), .ZN(U2817)
         );
  NAND2_X1 U7189 ( .A1(n6194), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n6164)
         );
  OAI211_X1 U7190 ( .C1(n6198), .C2(n6382), .A(n6165), .B(n6164), .ZN(n6168)
         );
  INV_X1 U7191 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6679) );
  NOR3_X1 U7192 ( .A1(n6166), .A2(n6679), .A3(REIP_REG_7__SCAN_IN), .ZN(n6167)
         );
  AOI211_X1 U7193 ( .C1(n6191), .C2(EBX_REG_7__SCAN_IN), .A(n6168), .B(n6167), 
        .ZN(n6169) );
  INV_X1 U7194 ( .A(n6169), .ZN(n6170) );
  AOI21_X1 U7195 ( .B1(n6331), .B2(n6171), .A(n6170), .ZN(n6174) );
  OAI21_X1 U7196 ( .B1(n6183), .B2(n6172), .A(REIP_REG_7__SCAN_IN), .ZN(n6173)
         );
  OAI211_X1 U7197 ( .C1(n6186), .C2(n6334), .A(n6174), .B(n6173), .ZN(U2820)
         );
  OAI22_X1 U7198 ( .A1(n6176), .A2(n3701), .B1(n6198), .B2(n6175), .ZN(n6177)
         );
  AOI211_X1 U7199 ( .C1(n6191), .C2(EBX_REG_5__SCAN_IN), .A(n6178), .B(n6177), 
        .ZN(n6185) );
  INV_X1 U7200 ( .A(n6179), .ZN(n6180) );
  OAI21_X1 U7201 ( .B1(n6181), .B2(n6180), .A(n4539), .ZN(n6182) );
  AOI22_X1 U7202 ( .A1(n6336), .A2(n6200), .B1(n6183), .B2(n6182), .ZN(n6184)
         );
  OAI211_X1 U7203 ( .C1(n6341), .C2(n6186), .A(n6185), .B(n6184), .ZN(U2822)
         );
  INV_X1 U7204 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6675) );
  OR2_X1 U7205 ( .A1(n6188), .A2(n6187), .ZN(n6202) );
  AOI22_X1 U7206 ( .A1(EBX_REG_3__SCAN_IN), .A2(n6191), .B1(n6190), .B2(n6189), 
        .ZN(n6196) );
  INV_X1 U7207 ( .A(n6349), .ZN(n6192) );
  AOI22_X1 U7208 ( .A1(PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n6194), .B1(n6193), 
        .B2(n6192), .ZN(n6195) );
  OAI211_X1 U7209 ( .C1(n6198), .C2(n6197), .A(n6196), .B(n6195), .ZN(n6199)
         );
  AOI21_X1 U7210 ( .B1(n6346), .B2(n6200), .A(n6199), .ZN(n6201) );
  OAI221_X1 U7211 ( .B1(n6203), .B2(n6675), .C1(n6203), .C2(n6202), .A(n6201), 
        .ZN(U2824) );
  AOI22_X1 U7212 ( .A1(n6204), .A2(n6211), .B1(n6210), .B2(DATAI_18_), .ZN(
        n6206) );
  AOI22_X1 U7213 ( .A1(n6214), .A2(DATAI_2_), .B1(n6213), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n6205) );
  NAND2_X1 U7214 ( .A1(n6206), .A2(n6205), .ZN(U2873) );
  AOI22_X1 U7215 ( .A1(n6207), .A2(n6211), .B1(n6210), .B2(DATAI_17_), .ZN(
        n6209) );
  AOI22_X1 U7216 ( .A1(n6214), .A2(DATAI_1_), .B1(n6213), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n6208) );
  NAND2_X1 U7217 ( .A1(n6209), .A2(n6208), .ZN(U2874) );
  AOI22_X1 U7218 ( .A1(n6212), .A2(n6211), .B1(n6210), .B2(DATAI_16_), .ZN(
        n6216) );
  AOI22_X1 U7219 ( .A1(n6214), .A2(DATAI_0_), .B1(n6213), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n6215) );
  NAND2_X1 U7220 ( .A1(n6216), .A2(n6215), .ZN(U2875) );
  INV_X1 U7221 ( .A(EAX_REG_15__SCAN_IN), .ZN(n6324) );
  AOI22_X1 U7222 ( .A1(n4333), .A2(LWORD_REG_15__SCAN_IN), .B1(n6229), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6218) );
  OAI21_X1 U7223 ( .B1(n6324), .B2(n6236), .A(n6218), .ZN(U2908) );
  INV_X1 U7224 ( .A(EAX_REG_14__SCAN_IN), .ZN(n6319) );
  AOI22_X1 U7225 ( .A1(n4333), .A2(LWORD_REG_14__SCAN_IN), .B1(n6229), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n6219) );
  OAI21_X1 U7226 ( .B1(n6319), .B2(n6236), .A(n6219), .ZN(U2909) );
  AOI22_X1 U7227 ( .A1(n4333), .A2(LWORD_REG_13__SCAN_IN), .B1(n6229), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n6220) );
  OAI21_X1 U7228 ( .B1(n6315), .B2(n6236), .A(n6220), .ZN(U2910) );
  INV_X1 U7229 ( .A(EAX_REG_12__SCAN_IN), .ZN(n6312) );
  AOI22_X1 U7230 ( .A1(n4333), .A2(LWORD_REG_12__SCAN_IN), .B1(n6229), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6221) );
  OAI21_X1 U7231 ( .B1(n6312), .B2(n6236), .A(n6221), .ZN(U2911) );
  AOI22_X1 U7232 ( .A1(n4333), .A2(LWORD_REG_11__SCAN_IN), .B1(n6229), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n6222) );
  OAI21_X1 U7233 ( .B1(n6309), .B2(n6236), .A(n6222), .ZN(U2912) );
  INV_X1 U7234 ( .A(EAX_REG_10__SCAN_IN), .ZN(n6306) );
  AOI22_X1 U7235 ( .A1(n4333), .A2(LWORD_REG_10__SCAN_IN), .B1(n6229), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n6223) );
  OAI21_X1 U7236 ( .B1(n6306), .B2(n6236), .A(n6223), .ZN(U2913) );
  AOI22_X1 U7237 ( .A1(n4333), .A2(LWORD_REG_9__SCAN_IN), .B1(n6229), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n6224) );
  OAI21_X1 U7238 ( .B1(n6303), .B2(n6236), .A(n6224), .ZN(U2914) );
  AOI22_X1 U7239 ( .A1(n4333), .A2(LWORD_REG_8__SCAN_IN), .B1(n6229), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n6225) );
  OAI21_X1 U7240 ( .B1(n6300), .B2(n6236), .A(n6225), .ZN(U2915) );
  AOI22_X1 U7241 ( .A1(n4333), .A2(LWORD_REG_7__SCAN_IN), .B1(n6229), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n6226) );
  OAI21_X1 U7242 ( .B1(n3739), .B2(n6236), .A(n6226), .ZN(U2916) );
  AOI22_X1 U7243 ( .A1(n4333), .A2(LWORD_REG_6__SCAN_IN), .B1(n6229), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n6227) );
  OAI21_X1 U7244 ( .B1(n6295), .B2(n6236), .A(n6227), .ZN(U2917) );
  INV_X1 U7245 ( .A(EAX_REG_5__SCAN_IN), .ZN(n6292) );
  AOI22_X1 U7246 ( .A1(n4333), .A2(LWORD_REG_5__SCAN_IN), .B1(n6229), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n6228) );
  OAI21_X1 U7247 ( .B1(n6292), .B2(n6236), .A(n6228), .ZN(U2918) );
  AOI22_X1 U7248 ( .A1(n4333), .A2(LWORD_REG_4__SCAN_IN), .B1(n6229), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n6230) );
  OAI21_X1 U7249 ( .B1(n6289), .B2(n6236), .A(n6230), .ZN(U2919) );
  AOI22_X1 U7250 ( .A1(n4333), .A2(LWORD_REG_3__SCAN_IN), .B1(n6234), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n6231) );
  OAI21_X1 U7251 ( .B1(n6286), .B2(n6236), .A(n6231), .ZN(U2920) );
  AOI22_X1 U7252 ( .A1(n4333), .A2(LWORD_REG_2__SCAN_IN), .B1(n6234), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n6232) );
  OAI21_X1 U7253 ( .B1(n6283), .B2(n6236), .A(n6232), .ZN(U2921) );
  AOI22_X1 U7254 ( .A1(n4333), .A2(LWORD_REG_1__SCAN_IN), .B1(n6234), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n6233) );
  OAI21_X1 U7255 ( .B1(n6280), .B2(n6236), .A(n6233), .ZN(U2922) );
  AOI22_X1 U7256 ( .A1(n4333), .A2(LWORD_REG_0__SCAN_IN), .B1(n6234), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n6235) );
  OAI21_X1 U7257 ( .B1(n6277), .B2(n6236), .A(n6235), .ZN(U2923) );
  INV_X1 U7258 ( .A(n6633), .ZN(n6237) );
  NAND2_X2 U7259 ( .A1(n6238), .A2(n6237), .ZN(n6323) );
  OAI21_X1 U7260 ( .B1(n6240), .B2(n6718), .A(n6239), .ZN(n6317) );
  INV_X1 U7261 ( .A(n6272), .ZN(n6320) );
  AND2_X1 U7262 ( .A1(n6320), .A2(DATAI_0_), .ZN(n6275) );
  AOI21_X1 U7263 ( .B1(UWORD_REG_0__SCAN_IN), .B2(n6321), .A(n6275), .ZN(n6241) );
  OAI21_X1 U7264 ( .B1(n6242), .B2(n6323), .A(n6241), .ZN(U2924) );
  AND2_X1 U7265 ( .A1(n6320), .A2(DATAI_1_), .ZN(n6278) );
  AOI21_X1 U7266 ( .B1(UWORD_REG_1__SCAN_IN), .B2(n6321), .A(n6278), .ZN(n6243) );
  OAI21_X1 U7267 ( .B1(n6244), .B2(n6323), .A(n6243), .ZN(U2925) );
  AND2_X1 U7268 ( .A1(n6320), .A2(DATAI_2_), .ZN(n6281) );
  AOI21_X1 U7269 ( .B1(UWORD_REG_2__SCAN_IN), .B2(n6321), .A(n6281), .ZN(n6245) );
  OAI21_X1 U7270 ( .B1(n6246), .B2(n6323), .A(n6245), .ZN(U2926) );
  AND2_X1 U7271 ( .A1(n6320), .A2(DATAI_3_), .ZN(n6284) );
  AOI21_X1 U7272 ( .B1(UWORD_REG_3__SCAN_IN), .B2(n6321), .A(n6284), .ZN(n6247) );
  OAI21_X1 U7273 ( .B1(n6248), .B2(n6323), .A(n6247), .ZN(U2927) );
  AND2_X1 U7274 ( .A1(n6320), .A2(DATAI_4_), .ZN(n6287) );
  AOI21_X1 U7275 ( .B1(UWORD_REG_4__SCAN_IN), .B2(n6321), .A(n6287), .ZN(n6249) );
  OAI21_X1 U7276 ( .B1(n6250), .B2(n6323), .A(n6249), .ZN(U2928) );
  NOR2_X1 U7277 ( .A1(n6272), .A2(n7086), .ZN(n6290) );
  AOI21_X1 U7278 ( .B1(UWORD_REG_5__SCAN_IN), .B2(n6321), .A(n6290), .ZN(n6251) );
  OAI21_X1 U7279 ( .B1(n6252), .B2(n6323), .A(n6251), .ZN(U2929) );
  AND2_X1 U7280 ( .A1(n6320), .A2(DATAI_6_), .ZN(n6293) );
  AOI21_X1 U7281 ( .B1(UWORD_REG_6__SCAN_IN), .B2(n6321), .A(n6293), .ZN(n6253) );
  OAI21_X1 U7282 ( .B1(n6254), .B2(n6323), .A(n6253), .ZN(U2930) );
  AND2_X1 U7283 ( .A1(n6320), .A2(DATAI_7_), .ZN(n6296) );
  AOI21_X1 U7284 ( .B1(UWORD_REG_7__SCAN_IN), .B2(n6321), .A(n6296), .ZN(n6255) );
  OAI21_X1 U7285 ( .B1(n6256), .B2(n6323), .A(n6255), .ZN(U2931) );
  AND2_X1 U7286 ( .A1(n6320), .A2(DATAI_8_), .ZN(n6298) );
  AOI21_X1 U7287 ( .B1(UWORD_REG_8__SCAN_IN), .B2(n6321), .A(n6298), .ZN(n6257) );
  OAI21_X1 U7288 ( .B1(n6258), .B2(n6323), .A(n6257), .ZN(U2932) );
  AND2_X1 U7289 ( .A1(n6320), .A2(DATAI_9_), .ZN(n6301) );
  AOI21_X1 U7290 ( .B1(UWORD_REG_9__SCAN_IN), .B2(n6321), .A(n6301), .ZN(n6259) );
  OAI21_X1 U7291 ( .B1(n6260), .B2(n6323), .A(n6259), .ZN(U2933) );
  INV_X1 U7292 ( .A(DATAI_10_), .ZN(n6261) );
  NOR2_X1 U7293 ( .A1(n6272), .A2(n6261), .ZN(n6304) );
  AOI21_X1 U7294 ( .B1(UWORD_REG_10__SCAN_IN), .B2(n6321), .A(n6304), .ZN(
        n6262) );
  OAI21_X1 U7295 ( .B1(n6263), .B2(n6323), .A(n6262), .ZN(U2934) );
  AND2_X1 U7296 ( .A1(n6320), .A2(DATAI_11_), .ZN(n6307) );
  AOI21_X1 U7297 ( .B1(UWORD_REG_11__SCAN_IN), .B2(n6321), .A(n6307), .ZN(
        n6264) );
  OAI21_X1 U7298 ( .B1(n6265), .B2(n6323), .A(n6264), .ZN(U2935) );
  INV_X1 U7299 ( .A(DATAI_12_), .ZN(n6266) );
  NOR2_X1 U7300 ( .A1(n6272), .A2(n6266), .ZN(n6310) );
  AOI21_X1 U7301 ( .B1(UWORD_REG_12__SCAN_IN), .B2(n6321), .A(n6310), .ZN(
        n6267) );
  OAI21_X1 U7302 ( .B1(n6268), .B2(n6323), .A(n6267), .ZN(U2936) );
  AND2_X1 U7303 ( .A1(n6320), .A2(DATAI_13_), .ZN(n6313) );
  AOI21_X1 U7304 ( .B1(UWORD_REG_13__SCAN_IN), .B2(n6321), .A(n6313), .ZN(
        n6269) );
  OAI21_X1 U7305 ( .B1(n6270), .B2(n6323), .A(n6269), .ZN(U2937) );
  INV_X1 U7306 ( .A(DATAI_14_), .ZN(n6271) );
  NOR2_X1 U7307 ( .A1(n6272), .A2(n6271), .ZN(n6316) );
  AOI21_X1 U7308 ( .B1(UWORD_REG_14__SCAN_IN), .B2(n6321), .A(n6316), .ZN(
        n6273) );
  OAI21_X1 U7309 ( .B1(n6274), .B2(n6323), .A(n6273), .ZN(U2938) );
  AOI21_X1 U7310 ( .B1(LWORD_REG_0__SCAN_IN), .B2(n6321), .A(n6275), .ZN(n6276) );
  OAI21_X1 U7311 ( .B1(n6277), .B2(n6323), .A(n6276), .ZN(U2939) );
  AOI21_X1 U7312 ( .B1(LWORD_REG_1__SCAN_IN), .B2(n6321), .A(n6278), .ZN(n6279) );
  OAI21_X1 U7313 ( .B1(n6280), .B2(n6323), .A(n6279), .ZN(U2940) );
  AOI21_X1 U7314 ( .B1(LWORD_REG_2__SCAN_IN), .B2(n6321), .A(n6281), .ZN(n6282) );
  OAI21_X1 U7315 ( .B1(n6283), .B2(n6323), .A(n6282), .ZN(U2941) );
  AOI21_X1 U7316 ( .B1(LWORD_REG_3__SCAN_IN), .B2(n6321), .A(n6284), .ZN(n6285) );
  OAI21_X1 U7317 ( .B1(n6286), .B2(n6323), .A(n6285), .ZN(U2942) );
  AOI21_X1 U7318 ( .B1(LWORD_REG_4__SCAN_IN), .B2(n6321), .A(n6287), .ZN(n6288) );
  OAI21_X1 U7319 ( .B1(n6289), .B2(n6323), .A(n6288), .ZN(U2943) );
  AOI21_X1 U7320 ( .B1(LWORD_REG_5__SCAN_IN), .B2(n6321), .A(n6290), .ZN(n6291) );
  OAI21_X1 U7321 ( .B1(n6292), .B2(n6323), .A(n6291), .ZN(U2944) );
  AOI21_X1 U7322 ( .B1(LWORD_REG_6__SCAN_IN), .B2(n6321), .A(n6293), .ZN(n6294) );
  OAI21_X1 U7323 ( .B1(n6295), .B2(n6323), .A(n6294), .ZN(U2945) );
  AOI21_X1 U7324 ( .B1(LWORD_REG_7__SCAN_IN), .B2(n6321), .A(n6296), .ZN(n6297) );
  OAI21_X1 U7325 ( .B1(n3739), .B2(n6323), .A(n6297), .ZN(U2946) );
  AOI21_X1 U7326 ( .B1(LWORD_REG_8__SCAN_IN), .B2(n6321), .A(n6298), .ZN(n6299) );
  OAI21_X1 U7327 ( .B1(n6300), .B2(n6323), .A(n6299), .ZN(U2947) );
  AOI21_X1 U7328 ( .B1(LWORD_REG_9__SCAN_IN), .B2(n6321), .A(n6301), .ZN(n6302) );
  OAI21_X1 U7329 ( .B1(n6303), .B2(n6323), .A(n6302), .ZN(U2948) );
  AOI21_X1 U7330 ( .B1(LWORD_REG_10__SCAN_IN), .B2(n6317), .A(n6304), .ZN(
        n6305) );
  OAI21_X1 U7331 ( .B1(n6306), .B2(n6323), .A(n6305), .ZN(U2949) );
  AOI21_X1 U7332 ( .B1(LWORD_REG_11__SCAN_IN), .B2(n6317), .A(n6307), .ZN(
        n6308) );
  OAI21_X1 U7333 ( .B1(n6309), .B2(n6323), .A(n6308), .ZN(U2950) );
  AOI21_X1 U7334 ( .B1(LWORD_REG_12__SCAN_IN), .B2(n6317), .A(n6310), .ZN(
        n6311) );
  OAI21_X1 U7335 ( .B1(n6312), .B2(n6323), .A(n6311), .ZN(U2951) );
  AOI21_X1 U7336 ( .B1(LWORD_REG_13__SCAN_IN), .B2(n6317), .A(n6313), .ZN(
        n6314) );
  OAI21_X1 U7337 ( .B1(n6315), .B2(n6323), .A(n6314), .ZN(U2952) );
  AOI21_X1 U7338 ( .B1(LWORD_REG_14__SCAN_IN), .B2(n6317), .A(n6316), .ZN(
        n6318) );
  OAI21_X1 U7339 ( .B1(n6319), .B2(n6323), .A(n6318), .ZN(U2953) );
  AOI22_X1 U7340 ( .A1(n6321), .A2(LWORD_REG_15__SCAN_IN), .B1(n6320), .B2(
        DATAI_15_), .ZN(n6322) );
  OAI21_X1 U7341 ( .B1(n6324), .B2(n6323), .A(n6322), .ZN(U2954) );
  AOI22_X1 U7342 ( .A1(n6422), .A2(REIP_REG_7__SCAN_IN), .B1(n6350), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n6333) );
  AND2_X1 U7343 ( .A1(n6326), .A2(n6325), .ZN(n6329) );
  OAI21_X1 U7344 ( .B1(n6329), .B2(n6328), .A(n3160), .ZN(n6330) );
  INV_X1 U7345 ( .A(n6330), .ZN(n6385) );
  AOI22_X1 U7346 ( .A1(n6385), .A2(n6356), .B1(n6354), .B2(n6331), .ZN(n6332)
         );
  OAI211_X1 U7347 ( .C1(n6360), .C2(n6334), .A(n6333), .B(n6332), .ZN(U2979)
         );
  AOI22_X1 U7348 ( .A1(n6422), .A2(REIP_REG_5__SCAN_IN), .B1(n6350), .B2(
        PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n6340) );
  INV_X1 U7349 ( .A(n6335), .ZN(n6338) );
  AOI22_X1 U7350 ( .A1(n6338), .A2(n6356), .B1(n6337), .B2(n6336), .ZN(n6339)
         );
  OAI211_X1 U7351 ( .C1(n6360), .C2(n6341), .A(n6340), .B(n6339), .ZN(U2981)
         );
  AOI22_X1 U7352 ( .A1(n6422), .A2(REIP_REG_3__SCAN_IN), .B1(n6350), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n6348) );
  OAI21_X1 U7353 ( .B1(n3164), .B2(n6343), .A(n3161), .ZN(n6345) );
  INV_X1 U7354 ( .A(n6345), .ZN(n6414) );
  AOI22_X1 U7355 ( .A1(n6346), .A2(n6354), .B1(n6356), .B2(n6414), .ZN(n6347)
         );
  OAI211_X1 U7356 ( .C1(n6360), .C2(n6349), .A(n6348), .B(n6347), .ZN(U2983)
         );
  AOI22_X1 U7357 ( .A1(n6422), .A2(REIP_REG_2__SCAN_IN), .B1(n6350), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6358) );
  XOR2_X1 U7358 ( .A(n6351), .B(INSTADDRPOINTER_REG_2__SCAN_IN), .Z(n6353) );
  XNOR2_X1 U7359 ( .A(n6353), .B(n6352), .ZN(n6430) );
  AOI22_X1 U7360 ( .A1(n6356), .A2(n6430), .B1(n6355), .B2(n6354), .ZN(n6357)
         );
  OAI211_X1 U7361 ( .C1(n6360), .C2(n6359), .A(n6358), .B(n6357), .ZN(U2984)
         );
  AOI21_X1 U7362 ( .B1(n6362), .B2(n6424), .A(n6361), .ZN(n6366) );
  AOI22_X1 U7363 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n6364), .B1(n6429), .B2(n6363), .ZN(n6365) );
  OAI211_X1 U7364 ( .C1(INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n6367), .A(n6366), .B(n6365), .ZN(U3007) );
  AOI21_X1 U7365 ( .B1(n6369), .B2(n6424), .A(n6368), .ZN(n6373) );
  AOI22_X1 U7366 ( .A1(n6371), .A2(n6429), .B1(INSTADDRPOINTER_REG_9__SCAN_IN), 
        .B2(n6370), .ZN(n6372) );
  OAI211_X1 U7367 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n6374), .A(n6373), 
        .B(n6372), .ZN(U3009) );
  INV_X1 U7368 ( .A(n6375), .ZN(n6376) );
  AOI222_X1 U7369 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6422), .B1(n6424), .B2(
        n6377), .C1(n6429), .C2(n6376), .ZN(n6380) );
  OAI211_X1 U7370 ( .C1(INSTADDRPOINTER_REG_7__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .A(n6384), .B(n6378), .ZN(n6379) );
  OAI211_X1 U7371 ( .C1(n6389), .C2(n6381), .A(n6380), .B(n6379), .ZN(U3010)
         );
  INV_X1 U7372 ( .A(n6382), .ZN(n6383) );
  AOI22_X1 U7373 ( .A1(n6424), .A2(n6383), .B1(n6422), .B2(REIP_REG_7__SCAN_IN), .ZN(n6387) );
  AOI22_X1 U7374 ( .A1(n6385), .A2(n6429), .B1(n6384), .B2(n6388), .ZN(n6386)
         );
  OAI211_X1 U7375 ( .C1(n6389), .C2(n6388), .A(n6387), .B(n6386), .ZN(U3011)
         );
  OAI222_X1 U7376 ( .A1(n6392), .A2(n6391), .B1(n6407), .B2(n6679), .C1(n6403), 
        .C2(n6390), .ZN(n6393) );
  INV_X1 U7377 ( .A(n6393), .ZN(n6394) );
  OAI221_X1 U7378 ( .B1(INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n6397), .C1(n6396), .C2(n6395), .A(n6394), .ZN(U3012) );
  AOI21_X1 U7379 ( .B1(n6399), .B2(n6420), .A(n6398), .ZN(n6416) );
  NAND2_X1 U7380 ( .A1(n6401), .A2(n6400), .ZN(n6418) );
  AOI211_X1 U7381 ( .C1(n6417), .C2(n6412), .A(n6402), .B(n6418), .ZN(n6410)
         );
  NOR2_X1 U7382 ( .A1(n6404), .A2(n6403), .ZN(n6409) );
  NAND2_X1 U7383 ( .A1(n6424), .A2(n6405), .ZN(n6406) );
  OAI21_X1 U7384 ( .B1(n6676), .B2(n6407), .A(n6406), .ZN(n6408) );
  NOR3_X1 U7385 ( .A1(n6410), .A2(n6409), .A3(n6408), .ZN(n6411) );
  OAI21_X1 U7386 ( .B1(n6416), .B2(n6412), .A(n6411), .ZN(U3014) );
  AOI222_X1 U7387 ( .A1(n6414), .A2(n6429), .B1(n6424), .B2(n6413), .C1(n6422), 
        .C2(REIP_REG_3__SCAN_IN), .ZN(n6415) );
  OAI221_X1 U7388 ( .B1(INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n6418), .C1(n6417), .C2(n6416), .A(n6415), .ZN(U3015) );
  NAND2_X1 U7389 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n6419), .ZN(n6433)
         );
  AOI21_X1 U7390 ( .B1(n6421), .B2(INSTADDRPOINTER_REG_0__SCAN_IN), .A(n6420), 
        .ZN(n6427) );
  AOI22_X1 U7391 ( .A1(n6424), .A2(n6423), .B1(n6422), .B2(REIP_REG_2__SCAN_IN), .ZN(n6425) );
  OAI21_X1 U7392 ( .B1(n6427), .B2(n6426), .A(n6425), .ZN(n6428) );
  AOI21_X1 U7393 ( .B1(n6430), .B2(n6429), .A(n6428), .ZN(n6431) );
  OAI221_X1 U7394 ( .B1(INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n6433), .C1(n4420), .C2(n6432), .A(n6431), .ZN(U3016) );
  INV_X1 U7395 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6435) );
  NOR2_X1 U7396 ( .A1(n6435), .A2(n6434), .ZN(U3019) );
  INV_X1 U7397 ( .A(n6436), .ZN(n6526) );
  NAND2_X1 U7398 ( .A1(n6526), .A2(n4929), .ZN(n6469) );
  OAI22_X1 U7399 ( .A1(n6476), .A2(n6546), .B1(n6527), .B2(n6469), .ZN(n6437)
         );
  INV_X1 U7400 ( .A(n6437), .ZN(n6450) );
  NAND2_X1 U7401 ( .A1(n6439), .A2(n6438), .ZN(n6440) );
  OAI21_X1 U7402 ( .B1(n6441), .B2(n6440), .A(n6530), .ZN(n6448) );
  OR2_X1 U7403 ( .A1(n6442), .A2(n6533), .ZN(n6443) );
  AND2_X1 U7404 ( .A1(n6443), .A2(n6469), .ZN(n6447) );
  INV_X1 U7405 ( .A(n6447), .ZN(n6445) );
  AOI21_X1 U7406 ( .B1(n6537), .B2(n6446), .A(n6536), .ZN(n6444) );
  OAI21_X1 U7407 ( .B1(n6448), .B2(n6445), .A(n6444), .ZN(n6473) );
  OAI22_X1 U7408 ( .A1(n6448), .A2(n6447), .B1(n6446), .B2(n6636), .ZN(n6472)
         );
  AOI22_X1 U7409 ( .A1(INSTQUEUE_REG_3__0__SCAN_IN), .A2(n6473), .B1(n6543), 
        .B2(n6472), .ZN(n6449) );
  OAI211_X1 U7410 ( .C1(n6528), .C2(n6470), .A(n6450), .B(n6449), .ZN(U3044)
         );
  OAI22_X1 U7411 ( .A1(n6470), .A2(n6548), .B1(n6547), .B2(n6469), .ZN(n6451)
         );
  INV_X1 U7412 ( .A(n6451), .ZN(n6453) );
  AOI22_X1 U7413 ( .A1(INSTQUEUE_REG_3__1__SCAN_IN), .A2(n6473), .B1(n6550), 
        .B2(n6472), .ZN(n6452) );
  OAI211_X1 U7414 ( .C1(n6553), .C2(n6476), .A(n6453), .B(n6452), .ZN(U3045)
         );
  OAI22_X1 U7415 ( .A1(n6470), .A2(n6560), .B1(n6554), .B2(n6469), .ZN(n6454)
         );
  INV_X1 U7416 ( .A(n6454), .ZN(n6456) );
  AOI22_X1 U7417 ( .A1(INSTQUEUE_REG_3__2__SCAN_IN), .A2(n6473), .B1(n6557), 
        .B2(n6472), .ZN(n6455) );
  OAI211_X1 U7418 ( .C1(n6555), .C2(n6476), .A(n6456), .B(n6455), .ZN(U3046)
         );
  OAI22_X1 U7419 ( .A1(n6476), .A2(n6562), .B1(n6561), .B2(n6469), .ZN(n6457)
         );
  INV_X1 U7420 ( .A(n6457), .ZN(n6459) );
  AOI22_X1 U7421 ( .A1(INSTQUEUE_REG_3__3__SCAN_IN), .A2(n6473), .B1(n6564), 
        .B2(n6472), .ZN(n6458) );
  OAI211_X1 U7422 ( .C1(n6470), .C2(n6567), .A(n6459), .B(n6458), .ZN(U3047)
         );
  OAI22_X1 U7423 ( .A1(n6470), .A2(n6569), .B1(n6568), .B2(n6469), .ZN(n6460)
         );
  INV_X1 U7424 ( .A(n6460), .ZN(n6462) );
  AOI22_X1 U7425 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n6473), .B1(n6571), 
        .B2(n6472), .ZN(n6461) );
  OAI211_X1 U7426 ( .C1(n6574), .C2(n6476), .A(n6462), .B(n6461), .ZN(U3048)
         );
  OAI22_X1 U7427 ( .A1(n6470), .A2(n6576), .B1(n6575), .B2(n6469), .ZN(n6463)
         );
  INV_X1 U7428 ( .A(n6463), .ZN(n6465) );
  AOI22_X1 U7429 ( .A1(INSTQUEUE_REG_3__5__SCAN_IN), .A2(n6473), .B1(n6578), 
        .B2(n6472), .ZN(n6464) );
  OAI211_X1 U7430 ( .C1(n6581), .C2(n6476), .A(n6465), .B(n6464), .ZN(U3049)
         );
  OAI22_X1 U7431 ( .A1(n6470), .A2(n6588), .B1(n6582), .B2(n6469), .ZN(n6466)
         );
  INV_X1 U7432 ( .A(n6466), .ZN(n6468) );
  AOI22_X1 U7433 ( .A1(INSTQUEUE_REG_3__6__SCAN_IN), .A2(n6473), .B1(n6585), 
        .B2(n6472), .ZN(n6467) );
  OAI211_X1 U7434 ( .C1(n6583), .C2(n6476), .A(n6468), .B(n6467), .ZN(U3050)
         );
  OAI22_X1 U7435 ( .A1(n6470), .A2(n6600), .B1(n6590), .B2(n6469), .ZN(n6471)
         );
  INV_X1 U7436 ( .A(n6471), .ZN(n6475) );
  AOI22_X1 U7437 ( .A1(INSTQUEUE_REG_3__7__SCAN_IN), .A2(n6473), .B1(n6595), 
        .B2(n6472), .ZN(n6474) );
  OAI211_X1 U7438 ( .C1(n6591), .C2(n6476), .A(n6475), .B(n6474), .ZN(U3051)
         );
  INV_X1 U7439 ( .A(n6525), .ZN(n6513) );
  INV_X1 U7440 ( .A(n6483), .ZN(n6518) );
  AOI22_X1 U7441 ( .A1(n6513), .A2(n6478), .B1(n6518), .B2(n6477), .ZN(n6490)
         );
  NAND2_X1 U7442 ( .A1(n6530), .A2(n6488), .ZN(n6479) );
  NAND2_X1 U7443 ( .A1(n6479), .A2(n6486), .ZN(n6480) );
  NAND2_X1 U7444 ( .A1(n6481), .A2(n6480), .ZN(n6522) );
  INV_X1 U7445 ( .A(n6482), .ZN(n6484) );
  OAI21_X1 U7446 ( .B1(n6484), .B2(n6533), .A(n6483), .ZN(n6485) );
  NAND2_X1 U7447 ( .A1(n6485), .A2(n6530), .ZN(n6487) );
  OAI22_X1 U7448 ( .A1(n6488), .A2(n6487), .B1(n6486), .B2(n6636), .ZN(n6521)
         );
  AOI22_X1 U7449 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n6522), .B1(n6543), 
        .B2(n6521), .ZN(n6489) );
  OAI211_X1 U7450 ( .C1(n6546), .C2(n6516), .A(n6490), .B(n6489), .ZN(U3076)
         );
  AOI22_X1 U7451 ( .A1(n6520), .A2(n6492), .B1(n6518), .B2(n6491), .ZN(n6494)
         );
  AOI22_X1 U7452 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n6522), .B1(n6550), 
        .B2(n6521), .ZN(n6493) );
  OAI211_X1 U7453 ( .C1(n6548), .C2(n6525), .A(n6494), .B(n6493), .ZN(U3077)
         );
  AOI22_X1 U7454 ( .A1(n6520), .A2(n6496), .B1(n6518), .B2(n6495), .ZN(n6498)
         );
  AOI22_X1 U7455 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n6522), .B1(n6557), 
        .B2(n6521), .ZN(n6497) );
  OAI211_X1 U7456 ( .C1(n6560), .C2(n6525), .A(n6498), .B(n6497), .ZN(U3078)
         );
  AOI22_X1 U7457 ( .A1(n6520), .A2(n6500), .B1(n6518), .B2(n6499), .ZN(n6502)
         );
  AOI22_X1 U7458 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n6522), .B1(n6564), 
        .B2(n6521), .ZN(n6501) );
  OAI211_X1 U7459 ( .C1(n6567), .C2(n6525), .A(n6502), .B(n6501), .ZN(U3079)
         );
  AOI22_X1 U7460 ( .A1(n6513), .A2(n6504), .B1(n6518), .B2(n6503), .ZN(n6506)
         );
  AOI22_X1 U7461 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n6522), .B1(n6571), 
        .B2(n6521), .ZN(n6505) );
  OAI211_X1 U7462 ( .C1(n6574), .C2(n6516), .A(n6506), .B(n6505), .ZN(U3080)
         );
  AOI22_X1 U7463 ( .A1(n6520), .A2(n6508), .B1(n6518), .B2(n6507), .ZN(n6510)
         );
  AOI22_X1 U7464 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n6522), .B1(n6578), 
        .B2(n6521), .ZN(n6509) );
  OAI211_X1 U7465 ( .C1(n6576), .C2(n6525), .A(n6510), .B(n6509), .ZN(U3081)
         );
  AOI22_X1 U7466 ( .A1(n6513), .A2(n6512), .B1(n6518), .B2(n6511), .ZN(n6515)
         );
  AOI22_X1 U7467 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n6522), .B1(n6585), 
        .B2(n6521), .ZN(n6514) );
  OAI211_X1 U7468 ( .C1(n6583), .C2(n6516), .A(n6515), .B(n6514), .ZN(U3082)
         );
  AOI22_X1 U7469 ( .A1(n6520), .A2(n6519), .B1(n6518), .B2(n6517), .ZN(n6524)
         );
  AOI22_X1 U7470 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n6522), .B1(n6595), 
        .B2(n6521), .ZN(n6523) );
  OAI211_X1 U7471 ( .C1(n6600), .C2(n6525), .A(n6524), .B(n6523), .ZN(U3083)
         );
  NAND2_X1 U7472 ( .A1(n6526), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6589) );
  OAI22_X1 U7473 ( .A1(n6599), .A2(n6528), .B1(n6527), .B2(n6589), .ZN(n6529)
         );
  INV_X1 U7474 ( .A(n6529), .ZN(n6545) );
  OAI21_X1 U7475 ( .B1(n6532), .B2(n6531), .A(n6530), .ZN(n6542) );
  OR2_X1 U7476 ( .A1(n6534), .A2(n6533), .ZN(n6535) );
  AND2_X1 U7477 ( .A1(n6535), .A2(n6589), .ZN(n6541) );
  INV_X1 U7478 ( .A(n6541), .ZN(n6539) );
  AOI21_X1 U7479 ( .B1(n6537), .B2(n6540), .A(n6536), .ZN(n6538) );
  OAI21_X1 U7480 ( .B1(n6542), .B2(n6539), .A(n6538), .ZN(n6596) );
  OAI22_X1 U7481 ( .A1(n6542), .A2(n6541), .B1(n6540), .B2(n6636), .ZN(n6594)
         );
  AOI22_X1 U7482 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6596), .B1(n6543), 
        .B2(n6594), .ZN(n6544) );
  OAI211_X1 U7483 ( .C1(n6546), .C2(n6592), .A(n6545), .B(n6544), .ZN(U3108)
         );
  OAI22_X1 U7484 ( .A1(n6599), .A2(n6548), .B1(n6547), .B2(n6589), .ZN(n6549)
         );
  INV_X1 U7485 ( .A(n6549), .ZN(n6552) );
  AOI22_X1 U7486 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6596), .B1(n6550), 
        .B2(n6594), .ZN(n6551) );
  OAI211_X1 U7487 ( .C1(n6553), .C2(n6592), .A(n6552), .B(n6551), .ZN(U3109)
         );
  OAI22_X1 U7488 ( .A1(n6592), .A2(n6555), .B1(n6554), .B2(n6589), .ZN(n6556)
         );
  INV_X1 U7489 ( .A(n6556), .ZN(n6559) );
  AOI22_X1 U7490 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6596), .B1(n6557), 
        .B2(n6594), .ZN(n6558) );
  OAI211_X1 U7491 ( .C1(n6560), .C2(n6599), .A(n6559), .B(n6558), .ZN(U3110)
         );
  OAI22_X1 U7492 ( .A1(n6592), .A2(n6562), .B1(n6561), .B2(n6589), .ZN(n6563)
         );
  INV_X1 U7493 ( .A(n6563), .ZN(n6566) );
  AOI22_X1 U7494 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6596), .B1(n6564), 
        .B2(n6594), .ZN(n6565) );
  OAI211_X1 U7495 ( .C1(n6567), .C2(n6599), .A(n6566), .B(n6565), .ZN(U3111)
         );
  OAI22_X1 U7496 ( .A1(n6599), .A2(n6569), .B1(n6568), .B2(n6589), .ZN(n6570)
         );
  INV_X1 U7497 ( .A(n6570), .ZN(n6573) );
  AOI22_X1 U7498 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6596), .B1(n6571), 
        .B2(n6594), .ZN(n6572) );
  OAI211_X1 U7499 ( .C1(n6574), .C2(n6592), .A(n6573), .B(n6572), .ZN(U3112)
         );
  OAI22_X1 U7500 ( .A1(n6599), .A2(n6576), .B1(n6575), .B2(n6589), .ZN(n6577)
         );
  INV_X1 U7501 ( .A(n6577), .ZN(n6580) );
  AOI22_X1 U7502 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6596), .B1(n6578), 
        .B2(n6594), .ZN(n6579) );
  OAI211_X1 U7503 ( .C1(n6581), .C2(n6592), .A(n6580), .B(n6579), .ZN(U3113)
         );
  OAI22_X1 U7504 ( .A1(n6592), .A2(n6583), .B1(n6582), .B2(n6589), .ZN(n6584)
         );
  INV_X1 U7505 ( .A(n6584), .ZN(n6587) );
  AOI22_X1 U7506 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6596), .B1(n6585), 
        .B2(n6594), .ZN(n6586) );
  OAI211_X1 U7507 ( .C1(n6588), .C2(n6599), .A(n6587), .B(n6586), .ZN(U3114)
         );
  OAI22_X1 U7508 ( .A1(n6592), .A2(n6591), .B1(n6590), .B2(n6589), .ZN(n6593)
         );
  INV_X1 U7509 ( .A(n6593), .ZN(n6598) );
  AOI22_X1 U7510 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6596), .B1(n6595), 
        .B2(n6594), .ZN(n6597) );
  OAI211_X1 U7511 ( .C1(n6600), .C2(n6599), .A(n6598), .B(n6597), .ZN(U3115)
         );
  INV_X1 U7512 ( .A(n6601), .ZN(n6607) );
  NOR2_X1 U7513 ( .A1(n6603), .A2(n6602), .ZN(n6606) );
  OAI21_X1 U7514 ( .B1(FLUSH_REG_SCAN_IN), .B2(MORE_REG_SCAN_IN), .A(n6604), 
        .ZN(n6605) );
  NAND3_X1 U7515 ( .A1(n6607), .A2(n6606), .A3(n6605), .ZN(n6608) );
  NOR2_X1 U7516 ( .A1(n6609), .A2(n6608), .ZN(n6630) );
  NOR2_X1 U7517 ( .A1(n6611), .A2(n6610), .ZN(n6612) );
  AND2_X1 U7518 ( .A1(n6613), .A2(n6612), .ZN(n6617) );
  NAND2_X1 U7519 ( .A1(n6617), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6619) );
  NAND2_X1 U7520 ( .A1(n6615), .A2(n6614), .ZN(n6616) );
  OAI21_X1 U7521 ( .B1(n6617), .B2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(n6616), 
        .ZN(n6618) );
  OAI211_X1 U7522 ( .C1(n6621), .C2(n6620), .A(n6619), .B(n6618), .ZN(n6623)
         );
  NAND2_X1 U7523 ( .A1(n6621), .A2(n6620), .ZN(n6622) );
  NAND2_X1 U7524 ( .A1(n6623), .A2(n6622), .ZN(n6625) );
  NAND2_X1 U7525 ( .A1(n6627), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6624) );
  NAND2_X1 U7526 ( .A1(n6625), .A2(n6624), .ZN(n6626) );
  OAI21_X1 U7527 ( .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n6627), .A(n6626), 
        .ZN(n6628) );
  NAND2_X1 U7528 ( .A1(n6628), .A2(n6435), .ZN(n6629) );
  NAND2_X1 U7529 ( .A1(n6630), .A2(n6629), .ZN(n6640) );
  NAND2_X1 U7530 ( .A1(READY_N), .A2(n4333), .ZN(n6631) );
  OAI21_X1 U7531 ( .B1(n6640), .B2(n6648), .A(n6631), .ZN(n6635) );
  OR2_X1 U7532 ( .A1(n6633), .A2(n6632), .ZN(n6634) );
  AOI21_X1 U7533 ( .B1(READY_N), .B2(n6636), .A(n6706), .ZN(n6646) );
  AOI211_X1 U7534 ( .C1(n6724), .C2(n6637), .A(STATE2_REG_0__SCAN_IN), .B(
        n6706), .ZN(n6638) );
  AOI211_X1 U7535 ( .C1(n6641), .C2(n6640), .A(n6639), .B(n6638), .ZN(n6642)
         );
  OAI221_X1 U7536 ( .B1(n6644), .B2(n6646), .C1(n6644), .C2(n6643), .A(n6642), 
        .ZN(U3148) );
  NOR3_X1 U7537 ( .A1(n6655), .A2(n6646), .A3(n6645), .ZN(n6650) );
  AOI221_X1 U7538 ( .B1(READY_N), .B2(n6648), .C1(n6647), .C2(n6648), .A(n6706), .ZN(n6649) );
  OR3_X1 U7539 ( .A1(n6651), .A2(n6650), .A3(n6649), .ZN(U3149) );
  OAI211_X1 U7540 ( .C1(STATE2_REG_2__SCAN_IN), .C2(n6718), .A(n6707), .B(
        n6652), .ZN(n6654) );
  OAI21_X1 U7541 ( .B1(n6655), .B2(n6654), .A(n6653), .ZN(U3150) );
  INV_X1 U7542 ( .A(n3155), .ZN(n6656) );
  AND2_X1 U7543 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6656), .ZN(U3151) );
  AND2_X1 U7544 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6656), .ZN(U3152) );
  AND2_X1 U7545 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6656), .ZN(U3153) );
  AND2_X1 U7546 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6656), .ZN(U3154) );
  AND2_X1 U7547 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6656), .ZN(U3155) );
  AND2_X1 U7548 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6656), .ZN(U3156) );
  AND2_X1 U7549 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6656), .ZN(U3157) );
  AND2_X1 U7550 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6656), .ZN(U3158) );
  AND2_X1 U7551 ( .A1(n6656), .A2(DATAWIDTH_REG_23__SCAN_IN), .ZN(U3159) );
  INV_X1 U7552 ( .A(DATAWIDTH_REG_22__SCAN_IN), .ZN(n6832) );
  NOR2_X1 U7553 ( .A1(n3155), .A2(n6832), .ZN(U3160) );
  AND2_X1 U7554 ( .A1(n6656), .A2(DATAWIDTH_REG_21__SCAN_IN), .ZN(U3161) );
  INV_X1 U7555 ( .A(DATAWIDTH_REG_20__SCAN_IN), .ZN(n7024) );
  NOR2_X1 U7556 ( .A1(n3155), .A2(n7024), .ZN(U3162) );
  INV_X1 U7557 ( .A(DATAWIDTH_REG_19__SCAN_IN), .ZN(n7057) );
  NOR2_X1 U7558 ( .A1(n3155), .A2(n7057), .ZN(U3163) );
  INV_X1 U7559 ( .A(DATAWIDTH_REG_18__SCAN_IN), .ZN(n7002) );
  NOR2_X1 U7560 ( .A1(n3155), .A2(n7002), .ZN(U3164) );
  INV_X1 U7561 ( .A(DATAWIDTH_REG_17__SCAN_IN), .ZN(n7037) );
  NOR2_X1 U7562 ( .A1(n3155), .A2(n7037), .ZN(U3165) );
  INV_X1 U7563 ( .A(DATAWIDTH_REG_16__SCAN_IN), .ZN(n7056) );
  NOR2_X1 U7564 ( .A1(n3155), .A2(n7056), .ZN(U3166) );
  AND2_X1 U7565 ( .A1(n6656), .A2(DATAWIDTH_REG_15__SCAN_IN), .ZN(U3167) );
  INV_X1 U7566 ( .A(DATAWIDTH_REG_14__SCAN_IN), .ZN(n7009) );
  NOR2_X1 U7567 ( .A1(n3155), .A2(n7009), .ZN(U3168) );
  AND2_X1 U7568 ( .A1(n6656), .A2(DATAWIDTH_REG_13__SCAN_IN), .ZN(U3169) );
  NOR2_X1 U7569 ( .A1(n3155), .A2(n7060), .ZN(U3170) );
  INV_X1 U7570 ( .A(DATAWIDTH_REG_11__SCAN_IN), .ZN(n6992) );
  NOR2_X1 U7571 ( .A1(n3155), .A2(n6992), .ZN(U3171) );
  INV_X1 U7572 ( .A(DATAWIDTH_REG_10__SCAN_IN), .ZN(n6986) );
  NOR2_X1 U7573 ( .A1(n3155), .A2(n6986), .ZN(U3172) );
  INV_X1 U7574 ( .A(DATAWIDTH_REG_9__SCAN_IN), .ZN(n7040) );
  NOR2_X1 U7575 ( .A1(n3155), .A2(n7040), .ZN(U3173) );
  INV_X1 U7576 ( .A(DATAWIDTH_REG_8__SCAN_IN), .ZN(n7070) );
  NOR2_X1 U7577 ( .A1(n3155), .A2(n7070), .ZN(U3174) );
  INV_X1 U7578 ( .A(DATAWIDTH_REG_7__SCAN_IN), .ZN(n6990) );
  NOR2_X1 U7579 ( .A1(n3155), .A2(n6990), .ZN(U3175) );
  INV_X1 U7580 ( .A(DATAWIDTH_REG_6__SCAN_IN), .ZN(n7083) );
  NOR2_X1 U7581 ( .A1(n3155), .A2(n7083), .ZN(U3176) );
  INV_X1 U7582 ( .A(DATAWIDTH_REG_5__SCAN_IN), .ZN(n7075) );
  NOR2_X1 U7583 ( .A1(n3155), .A2(n7075), .ZN(U3177) );
  NOR2_X1 U7584 ( .A1(n3155), .A2(n7051), .ZN(U3178) );
  AND2_X1 U7585 ( .A1(n6656), .A2(DATAWIDTH_REG_3__SCAN_IN), .ZN(U3179) );
  INV_X1 U7586 ( .A(DATAWIDTH_REG_2__SCAN_IN), .ZN(n7090) );
  NOR2_X1 U7587 ( .A1(n3155), .A2(n7090), .ZN(U3180) );
  INV_X1 U7588 ( .A(n6671), .ZN(n6658) );
  AOI22_X1 U7589 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .B1(
        STATE_REG_2__SCAN_IN), .B2(HOLD), .ZN(n6672) );
  INV_X1 U7590 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6663) );
  OAI221_X1 U7591 ( .B1(n6673), .B2(NA_N), .C1(n6673), .C2(n6663), .A(n6993), 
        .ZN(n6666) );
  INV_X1 U7592 ( .A(HOLD), .ZN(n7031) );
  NOR2_X1 U7593 ( .A1(n6663), .A2(n7031), .ZN(n6660) );
  INV_X1 U7594 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n7003) );
  OAI21_X1 U7595 ( .B1(n6660), .B2(n7003), .A(n7122), .ZN(n6657) );
  OAI211_X1 U7596 ( .C1(n6658), .C2(n6672), .A(n6666), .B(n6657), .ZN(U3181)
         );
  NOR2_X1 U7597 ( .A1(n6993), .A2(n7003), .ZN(n6668) );
  NAND2_X1 U7598 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n6659) );
  OAI21_X1 U7599 ( .B1(n6668), .B2(n6660), .A(n6659), .ZN(n6661) );
  OAI211_X1 U7600 ( .C1(n6663), .C2(n6718), .A(n6662), .B(n6661), .ZN(U3182)
         );
  NOR2_X1 U7601 ( .A1(NA_N), .A2(n6718), .ZN(n6664) );
  OAI21_X1 U7602 ( .B1(n6664), .B2(n6663), .A(n7003), .ZN(n6665) );
  AOI21_X1 U7603 ( .B1(n6673), .B2(n6665), .A(n7031), .ZN(n6667) );
  OAI21_X1 U7604 ( .B1(n6993), .B2(n6667), .A(n6666), .ZN(n6670) );
  INV_X1 U7605 ( .A(NA_N), .ZN(n6967) );
  NAND4_X1 U7606 ( .A1(STATE_REG_1__SCAN_IN), .A2(READY_N), .A3(n6668), .A4(
        n6967), .ZN(n6669) );
  OAI211_X1 U7607 ( .C1(n6672), .C2(n6671), .A(n6670), .B(n6669), .ZN(U3183)
         );
  NAND2_X1 U7608 ( .A1(n7123), .A2(n6673), .ZN(n6700) );
  INV_X1 U7609 ( .A(ADDRESS_REG_0__SCAN_IN), .ZN(n7006) );
  OAI222_X1 U7610 ( .A1(n6700), .A2(n6187), .B1(n7006), .B2(n7123), .C1(n6710), 
        .C2(n6696), .ZN(U3184) );
  INV_X1 U7611 ( .A(ADDRESS_REG_1__SCAN_IN), .ZN(n6834) );
  OAI222_X1 U7612 ( .A1(n6696), .A2(n6187), .B1(n6834), .B2(n7123), .C1(n6675), 
        .C2(n6697), .ZN(U3185) );
  INV_X1 U7613 ( .A(ADDRESS_REG_2__SCAN_IN), .ZN(n6674) );
  OAI222_X1 U7614 ( .A1(n6696), .A2(n6675), .B1(n6674), .B2(n7123), .C1(n6676), 
        .C2(n6697), .ZN(U3186) );
  INV_X1 U7615 ( .A(ADDRESS_REG_3__SCAN_IN), .ZN(n6984) );
  OAI222_X1 U7616 ( .A1(n6696), .A2(n6676), .B1(n6984), .B2(n7123), .C1(n4539), 
        .C2(n6700), .ZN(U3187) );
  INV_X1 U7617 ( .A(ADDRESS_REG_4__SCAN_IN), .ZN(n6677) );
  OAI222_X1 U7618 ( .A1(n6700), .A2(n6679), .B1(n6677), .B2(n7123), .C1(n4539), 
        .C2(n6696), .ZN(U3188) );
  INV_X1 U7619 ( .A(ADDRESS_REG_5__SCAN_IN), .ZN(n6678) );
  INV_X1 U7620 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6680) );
  OAI222_X1 U7621 ( .A1(n6696), .A2(n6679), .B1(n6678), .B2(n7123), .C1(n6680), 
        .C2(n6697), .ZN(U3189) );
  INV_X1 U7622 ( .A(ADDRESS_REG_6__SCAN_IN), .ZN(n7076) );
  OAI222_X1 U7623 ( .A1(n6696), .A2(n6680), .B1(n7076), .B2(n7123), .C1(n6681), 
        .C2(n6700), .ZN(U3190) );
  INV_X1 U7624 ( .A(ADDRESS_REG_7__SCAN_IN), .ZN(n6836) );
  OAI222_X1 U7625 ( .A1(n6697), .A2(n6682), .B1(n6836), .B2(n7123), .C1(n6681), 
        .C2(n6696), .ZN(U3191) );
  INV_X1 U7626 ( .A(ADDRESS_REG_8__SCAN_IN), .ZN(n7023) );
  OAI222_X1 U7627 ( .A1(n6696), .A2(n6682), .B1(n7023), .B2(n7123), .C1(n6683), 
        .C2(n6700), .ZN(U3192) );
  INV_X1 U7628 ( .A(ADDRESS_REG_9__SCAN_IN), .ZN(n7033) );
  OAI222_X1 U7629 ( .A1(n6696), .A2(n6683), .B1(n7033), .B2(n7123), .C1(n6684), 
        .C2(n6697), .ZN(U3193) );
  INV_X1 U7630 ( .A(ADDRESS_REG_10__SCAN_IN), .ZN(n6831) );
  OAI222_X1 U7631 ( .A1(n6696), .A2(n6684), .B1(n6831), .B2(n7123), .C1(n5401), 
        .C2(n6697), .ZN(U3194) );
  INV_X1 U7632 ( .A(ADDRESS_REG_11__SCAN_IN), .ZN(n7021) );
  INV_X1 U7633 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6686) );
  OAI222_X1 U7634 ( .A1(n6696), .A2(n5401), .B1(n7021), .B2(n7123), .C1(n6686), 
        .C2(n6700), .ZN(U3195) );
  INV_X1 U7635 ( .A(ADDRESS_REG_12__SCAN_IN), .ZN(n6685) );
  OAI222_X1 U7636 ( .A1(n6696), .A2(n6686), .B1(n6685), .B2(n7123), .C1(n6687), 
        .C2(n6700), .ZN(U3196) );
  INV_X1 U7637 ( .A(ADDRESS_REG_13__SCAN_IN), .ZN(n6688) );
  OAI222_X1 U7638 ( .A1(n6700), .A2(n5840), .B1(n6688), .B2(n7123), .C1(n6687), 
        .C2(n6696), .ZN(U3197) );
  INV_X1 U7639 ( .A(ADDRESS_REG_14__SCAN_IN), .ZN(n6837) );
  OAI222_X1 U7640 ( .A1(n6696), .A2(n5840), .B1(n6837), .B2(n7123), .C1(n5371), 
        .C2(n6700), .ZN(U3198) );
  INV_X1 U7641 ( .A(ADDRESS_REG_15__SCAN_IN), .ZN(n6689) );
  OAI222_X1 U7642 ( .A1(n6696), .A2(n5371), .B1(n6689), .B2(n7123), .C1(n7088), 
        .C2(n6697), .ZN(U3199) );
  INV_X1 U7643 ( .A(ADDRESS_REG_16__SCAN_IN), .ZN(n6823) );
  OAI222_X1 U7644 ( .A1(n6696), .A2(n7088), .B1(n6823), .B2(n7123), .C1(n7073), 
        .C2(n6697), .ZN(U3200) );
  INV_X1 U7645 ( .A(ADDRESS_REG_17__SCAN_IN), .ZN(n7069) );
  OAI222_X1 U7646 ( .A1(n6697), .A2(n6861), .B1(n7069), .B2(n7123), .C1(n7073), 
        .C2(n6696), .ZN(U3201) );
  INV_X1 U7647 ( .A(ADDRESS_REG_18__SCAN_IN), .ZN(n6690) );
  OAI222_X1 U7648 ( .A1(n6696), .A2(n6861), .B1(n6690), .B2(n7123), .C1(n6691), 
        .C2(n6697), .ZN(U3202) );
  INV_X1 U7649 ( .A(ADDRESS_REG_19__SCAN_IN), .ZN(n6872) );
  OAI222_X1 U7650 ( .A1(n6696), .A2(n6691), .B1(n6872), .B2(n7123), .C1(n6693), 
        .C2(n6697), .ZN(U3203) );
  INV_X1 U7651 ( .A(ADDRESS_REG_20__SCAN_IN), .ZN(n6692) );
  OAI222_X1 U7652 ( .A1(n6696), .A2(n6693), .B1(n6692), .B2(n7123), .C1(n7106), 
        .C2(n6697), .ZN(U3204) );
  INV_X1 U7653 ( .A(ADDRESS_REG_21__SCAN_IN), .ZN(n6820) );
  OAI222_X1 U7654 ( .A1(n6696), .A2(n7106), .B1(n6820), .B2(n7123), .C1(n6694), 
        .C2(n6697), .ZN(U3205) );
  INV_X1 U7655 ( .A(ADDRESS_REG_22__SCAN_IN), .ZN(n6968) );
  OAI222_X1 U7656 ( .A1(n6696), .A2(n6694), .B1(n6968), .B2(n7123), .C1(n7017), 
        .C2(n6697), .ZN(U3206) );
  INV_X1 U7657 ( .A(ADDRESS_REG_23__SCAN_IN), .ZN(n6964) );
  OAI222_X1 U7658 ( .A1(n6697), .A2(n6825), .B1(n6964), .B2(n7123), .C1(n7017), 
        .C2(n6696), .ZN(U3207) );
  INV_X1 U7659 ( .A(ADDRESS_REG_24__SCAN_IN), .ZN(n7066) );
  OAI222_X1 U7660 ( .A1(n6696), .A2(n6825), .B1(n7066), .B2(n7123), .C1(n7050), 
        .C2(n6697), .ZN(U3208) );
  INV_X1 U7661 ( .A(ADDRESS_REG_25__SCAN_IN), .ZN(n6695) );
  OAI222_X1 U7662 ( .A1(n6696), .A2(n7050), .B1(n6695), .B2(n7123), .C1(n7030), 
        .C2(n6697), .ZN(U3209) );
  INV_X1 U7663 ( .A(ADDRESS_REG_26__SCAN_IN), .ZN(n6864) );
  OAI222_X1 U7664 ( .A1(n6696), .A2(n7030), .B1(n6864), .B2(n7123), .C1(n7020), 
        .C2(n6697), .ZN(U3210) );
  INV_X1 U7665 ( .A(ADDRESS_REG_27__SCAN_IN), .ZN(n6970) );
  OAI222_X1 U7666 ( .A1(n6696), .A2(n7020), .B1(n6970), .B2(n7123), .C1(n7100), 
        .C2(n6697), .ZN(U3211) );
  INV_X1 U7667 ( .A(ADDRESS_REG_28__SCAN_IN), .ZN(n6698) );
  OAI222_X1 U7668 ( .A1(n6696), .A2(n7100), .B1(n6698), .B2(n7123), .C1(n4193), 
        .C2(n6697), .ZN(U3212) );
  INV_X1 U7669 ( .A(ADDRESS_REG_29__SCAN_IN), .ZN(n6699) );
  OAI222_X1 U7670 ( .A1(n6700), .A2(n7082), .B1(n6699), .B2(n7123), .C1(n4193), 
        .C2(n6696), .ZN(U3213) );
  OAI22_X1 U7671 ( .A1(n7122), .A2(BYTEENABLE_REG_2__SCAN_IN), .B1(
        BE_N_REG_2__SCAN_IN), .B2(n7123), .ZN(n6701) );
  INV_X1 U7672 ( .A(n6701), .ZN(U3446) );
  INV_X1 U7673 ( .A(BE_N_REG_1__SCAN_IN), .ZN(n6870) );
  AOI22_X1 U7674 ( .A1(n7123), .A2(n7034), .B1(n6870), .B2(n7122), .ZN(U3447)
         );
  OAI22_X1 U7675 ( .A1(n7122), .A2(BYTEENABLE_REG_0__SCAN_IN), .B1(
        BE_N_REG_0__SCAN_IN), .B2(n7123), .ZN(n6702) );
  INV_X1 U7676 ( .A(n6702), .ZN(U3448) );
  OAI21_X1 U7677 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(n3155), .A(n6704), .ZN(
        n6703) );
  INV_X1 U7678 ( .A(n6703), .ZN(U3451) );
  OAI21_X1 U7679 ( .B1(n3155), .B2(n7107), .A(n6704), .ZN(U3452) );
  INV_X1 U7680 ( .A(n6706), .ZN(n6708) );
  OAI221_X1 U7681 ( .B1(n6709), .B2(STATE2_REG_0__SCAN_IN), .C1(n6709), .C2(
        n6708), .A(n6707), .ZN(U3453) );
  AOI21_X1 U7682 ( .B1(REIP_REG_0__SCAN_IN), .B2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6711) );
  AOI22_X1 U7683 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .B1(
        n6711), .B2(n6710), .ZN(n6712) );
  INV_X1 U7684 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n7018) );
  AOI22_X1 U7685 ( .A1(n6713), .A2(n6712), .B1(n7018), .B2(n6716), .ZN(U3468)
         );
  INV_X1 U7686 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n7103) );
  INV_X1 U7687 ( .A(REIP_REG_0__SCAN_IN), .ZN(n6715) );
  AOI22_X1 U7688 ( .A1(n7103), .A2(n6716), .B1(n6715), .B2(n6714), .ZN(U3469)
         );
  INV_X1 U7689 ( .A(READREQUEST_REG_SCAN_IN), .ZN(n7059) );
  OAI22_X1 U7690 ( .A1(n7122), .A2(n7059), .B1(W_R_N_REG_SCAN_IN), .B2(n7123), 
        .ZN(n6717) );
  INV_X1 U7691 ( .A(n6717), .ZN(U3470) );
  AND2_X1 U7692 ( .A1(n6718), .A2(n4333), .ZN(n6719) );
  NOR4_X1 U7693 ( .A1(n6721), .A2(n6720), .A3(n6530), .A4(n6719), .ZN(n6728)
         );
  OAI211_X1 U7694 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n6723), .A(n6722), .B(
        STATE2_REG_2__SCAN_IN), .ZN(n6725) );
  AOI21_X1 U7695 ( .B1(n6725), .B2(STATE2_REG_0__SCAN_IN), .A(n6724), .ZN(
        n6727) );
  NAND2_X1 U7696 ( .A1(n6728), .A2(REQUESTPENDING_REG_SCAN_IN), .ZN(n6726) );
  OAI21_X1 U7697 ( .B1(n6728), .B2(n6727), .A(n6726), .ZN(U3472) );
  INV_X1 U7698 ( .A(M_IO_N_REG_SCAN_IN), .ZN(n6903) );
  AOI22_X1 U7699 ( .A1(n7123), .A2(n7054), .B1(n6903), .B2(n7122), .ZN(U3473)
         );
  AOI22_X1 U7700 ( .A1(keyinput_f41), .A2(D_C_N_REG_SCAN_IN), .B1(READY_N), 
        .B2(keyinput_f35), .ZN(n6729) );
  OAI221_X1 U7701 ( .B1(keyinput_f41), .B2(D_C_N_REG_SCAN_IN), .C1(READY_N), 
        .C2(keyinput_f35), .A(n6729), .ZN(n6736) );
  AOI22_X1 U7702 ( .A1(DATAI_26_), .A2(keyinput_f5), .B1(REIP_REG_31__SCAN_IN), 
        .B2(keyinput_f51), .ZN(n6730) );
  OAI221_X1 U7703 ( .B1(DATAI_26_), .B2(keyinput_f5), .C1(REIP_REG_31__SCAN_IN), .C2(keyinput_f51), .A(n6730), .ZN(n6735) );
  AOI22_X1 U7704 ( .A1(keyinput_f111), .A2(DATAWIDTH_REG_7__SCAN_IN), .B1(
        DATAI_8_), .B2(keyinput_f23), .ZN(n6731) );
  OAI221_X1 U7705 ( .B1(keyinput_f111), .B2(DATAWIDTH_REG_7__SCAN_IN), .C1(
        DATAI_8_), .C2(keyinput_f23), .A(n6731), .ZN(n6734) );
  AOI22_X1 U7706 ( .A1(keyinput_f82), .A2(ADDRESS_REG_18__SCAN_IN), .B1(
        keyinput_f80), .B2(ADDRESS_REG_20__SCAN_IN), .ZN(n6732) );
  OAI221_X1 U7707 ( .B1(keyinput_f82), .B2(ADDRESS_REG_18__SCAN_IN), .C1(
        keyinput_f80), .C2(ADDRESS_REG_20__SCAN_IN), .A(n6732), .ZN(n6733) );
  NOR4_X1 U7708 ( .A1(n6736), .A2(n6735), .A3(n6734), .A4(n6733), .ZN(n6897)
         );
  AOI22_X1 U7709 ( .A1(keyinput_f75), .A2(ADDRESS_REG_25__SCAN_IN), .B1(
        keyinput_f98), .B2(ADDRESS_REG_2__SCAN_IN), .ZN(n6737) );
  OAI221_X1 U7710 ( .B1(keyinput_f75), .B2(ADDRESS_REG_25__SCAN_IN), .C1(
        keyinput_f98), .C2(ADDRESS_REG_2__SCAN_IN), .A(n6737), .ZN(n6762) );
  OAI22_X1 U7711 ( .A1(DATAI_19_), .A2(keyinput_f12), .B1(DATAI_1_), .B2(
        keyinput_f30), .ZN(n6738) );
  AOI221_X1 U7712 ( .B1(DATAI_19_), .B2(keyinput_f12), .C1(keyinput_f30), .C2(
        DATAI_1_), .A(n6738), .ZN(n6742) );
  AOI22_X1 U7713 ( .A1(keyinput_f121), .A2(DATAWIDTH_REG_17__SCAN_IN), .B1(
        DATAI_5_), .B2(keyinput_f26), .ZN(n6739) );
  OAI221_X1 U7714 ( .B1(keyinput_f121), .B2(DATAWIDTH_REG_17__SCAN_IN), .C1(
        DATAI_5_), .C2(keyinput_f26), .A(n6739), .ZN(n6740) );
  AOI21_X1 U7715 ( .B1(keyinput_f25), .B2(n6989), .A(n6740), .ZN(n6741) );
  OAI211_X1 U7716 ( .C1(keyinput_f25), .C2(n6989), .A(n6742), .B(n6741), .ZN(
        n6761) );
  OAI22_X1 U7717 ( .A1(DATAI_18_), .A2(keyinput_f13), .B1(
        DATAWIDTH_REG_18__SCAN_IN), .B2(keyinput_f122), .ZN(n6743) );
  AOI221_X1 U7718 ( .B1(DATAI_18_), .B2(keyinput_f13), .C1(keyinput_f122), 
        .C2(DATAWIDTH_REG_18__SCAN_IN), .A(n6743), .ZN(n6750) );
  OAI22_X1 U7719 ( .A1(DATAI_12_), .A2(keyinput_f19), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(keyinput_f77), .ZN(n6744) );
  AOI221_X1 U7720 ( .B1(DATAI_12_), .B2(keyinput_f19), .C1(keyinput_f77), .C2(
        ADDRESS_REG_23__SCAN_IN), .A(n6744), .ZN(n6749) );
  OAI22_X1 U7721 ( .A1(STATE_REG_2__SCAN_IN), .A2(keyinput_f101), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(keyinput_f91), .ZN(n6745) );
  AOI221_X1 U7722 ( .B1(STATE_REG_2__SCAN_IN), .B2(keyinput_f101), .C1(
        keyinput_f91), .C2(ADDRESS_REG_9__SCAN_IN), .A(n6745), .ZN(n6748) );
  OAI22_X1 U7723 ( .A1(DATAI_25_), .A2(keyinput_f6), .B1(keyinput_f44), .B2(
        MORE_REG_SCAN_IN), .ZN(n6746) );
  AOI221_X1 U7724 ( .B1(DATAI_25_), .B2(keyinput_f6), .C1(MORE_REG_SCAN_IN), 
        .C2(keyinput_f44), .A(n6746), .ZN(n6747) );
  NAND4_X1 U7725 ( .A1(n6750), .A2(n6749), .A3(n6748), .A4(n6747), .ZN(n6760)
         );
  OAI22_X1 U7726 ( .A1(MEMORYFETCH_REG_SCAN_IN), .A2(keyinput_f32), .B1(
        BE_N_REG_2__SCAN_IN), .B2(keyinput_f68), .ZN(n6751) );
  AOI221_X1 U7727 ( .B1(MEMORYFETCH_REG_SCAN_IN), .B2(keyinput_f32), .C1(
        keyinput_f68), .C2(BE_N_REG_2__SCAN_IN), .A(n6751), .ZN(n6758) );
  OAI22_X1 U7728 ( .A1(keyinput_f97), .A2(ADDRESS_REG_3__SCAN_IN), .B1(
        keyinput_f47), .B2(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6752) );
  AOI221_X1 U7729 ( .B1(keyinput_f97), .B2(ADDRESS_REG_3__SCAN_IN), .C1(
        BYTEENABLE_REG_0__SCAN_IN), .C2(keyinput_f47), .A(n6752), .ZN(n6757)
         );
  OAI22_X1 U7730 ( .A1(DATAI_11_), .A2(keyinput_f20), .B1(DATAI_22_), .B2(
        keyinput_f9), .ZN(n6753) );
  AOI221_X1 U7731 ( .B1(DATAI_11_), .B2(keyinput_f20), .C1(keyinput_f9), .C2(
        DATAI_22_), .A(n6753), .ZN(n6756) );
  OAI22_X1 U7732 ( .A1(keyinput_f112), .A2(DATAWIDTH_REG_8__SCAN_IN), .B1(
        keyinput_f115), .B2(DATAWIDTH_REG_11__SCAN_IN), .ZN(n6754) );
  AOI221_X1 U7733 ( .B1(keyinput_f112), .B2(DATAWIDTH_REG_8__SCAN_IN), .C1(
        DATAWIDTH_REG_11__SCAN_IN), .C2(keyinput_f115), .A(n6754), .ZN(n6755)
         );
  NAND4_X1 U7734 ( .A1(n6758), .A2(n6757), .A3(n6756), .A4(n6755), .ZN(n6759)
         );
  NOR4_X1 U7735 ( .A1(n6762), .A2(n6761), .A3(n6760), .A4(n6759), .ZN(n6896)
         );
  OAI22_X1 U7736 ( .A1(keyinput_f73), .A2(ADDRESS_REG_27__SCAN_IN), .B1(
        keyinput_f72), .B2(ADDRESS_REG_28__SCAN_IN), .ZN(n6763) );
  AOI221_X1 U7737 ( .B1(keyinput_f73), .B2(ADDRESS_REG_27__SCAN_IN), .C1(
        ADDRESS_REG_28__SCAN_IN), .C2(keyinput_f72), .A(n6763), .ZN(n6770) );
  OAI22_X1 U7738 ( .A1(REIP_REG_23__SCAN_IN), .A2(keyinput_f59), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(keyinput_f85), .ZN(n6764) );
  AOI221_X1 U7739 ( .B1(REIP_REG_23__SCAN_IN), .B2(keyinput_f59), .C1(
        keyinput_f85), .C2(ADDRESS_REG_15__SCAN_IN), .A(n6764), .ZN(n6769) );
  OAI22_X1 U7740 ( .A1(keyinput_f48), .A2(BYTEENABLE_REG_1__SCAN_IN), .B1(
        keyinput_f127), .B2(DATAWIDTH_REG_23__SCAN_IN), .ZN(n6765) );
  AOI221_X1 U7741 ( .B1(keyinput_f48), .B2(BYTEENABLE_REG_1__SCAN_IN), .C1(
        DATAWIDTH_REG_23__SCAN_IN), .C2(keyinput_f127), .A(n6765), .ZN(n6768)
         );
  OAI22_X1 U7742 ( .A1(DATAI_24_), .A2(keyinput_f7), .B1(keyinput_f34), .B2(
        BS16_N), .ZN(n6766) );
  AOI221_X1 U7743 ( .B1(DATAI_24_), .B2(keyinput_f7), .C1(BS16_N), .C2(
        keyinput_f34), .A(n6766), .ZN(n6767) );
  NAND4_X1 U7744 ( .A1(n6770), .A2(n6769), .A3(n6768), .A4(n6767), .ZN(n6798)
         );
  OAI22_X1 U7745 ( .A1(DATAI_0_), .A2(keyinput_f31), .B1(DATAI_16_), .B2(
        keyinput_f15), .ZN(n6771) );
  AOI221_X1 U7746 ( .B1(DATAI_0_), .B2(keyinput_f31), .C1(keyinput_f15), .C2(
        DATAI_16_), .A(n6771), .ZN(n6778) );
  OAI22_X1 U7747 ( .A1(STATE_REG_0__SCAN_IN), .A2(keyinput_f103), .B1(
        keyinput_f46), .B2(W_R_N_REG_SCAN_IN), .ZN(n6772) );
  AOI221_X1 U7748 ( .B1(STATE_REG_0__SCAN_IN), .B2(keyinput_f103), .C1(
        W_R_N_REG_SCAN_IN), .C2(keyinput_f46), .A(n6772), .ZN(n6777) );
  OAI22_X1 U7749 ( .A1(keyinput_f96), .A2(ADDRESS_REG_4__SCAN_IN), .B1(
        keyinput_f38), .B2(ADS_N_REG_SCAN_IN), .ZN(n6773) );
  AOI221_X1 U7750 ( .B1(keyinput_f96), .B2(ADDRESS_REG_4__SCAN_IN), .C1(
        ADS_N_REG_SCAN_IN), .C2(keyinput_f38), .A(n6773), .ZN(n6776) );
  OAI22_X1 U7751 ( .A1(keyinput_f88), .A2(ADDRESS_REG_12__SCAN_IN), .B1(
        keyinput_f87), .B2(ADDRESS_REG_13__SCAN_IN), .ZN(n6774) );
  AOI221_X1 U7752 ( .B1(keyinput_f88), .B2(ADDRESS_REG_12__SCAN_IN), .C1(
        ADDRESS_REG_13__SCAN_IN), .C2(keyinput_f87), .A(n6774), .ZN(n6775) );
  NAND4_X1 U7753 ( .A1(n6778), .A2(n6777), .A3(n6776), .A4(n6775), .ZN(n6797)
         );
  OAI22_X1 U7754 ( .A1(DATAI_30_), .A2(keyinput_f1), .B1(keyinput_f105), .B2(
        DATAWIDTH_REG_1__SCAN_IN), .ZN(n6779) );
  AOI221_X1 U7755 ( .B1(DATAI_30_), .B2(keyinput_f1), .C1(
        DATAWIDTH_REG_1__SCAN_IN), .C2(keyinput_f105), .A(n6779), .ZN(n6786)
         );
  OAI22_X1 U7756 ( .A1(REIP_REG_22__SCAN_IN), .A2(keyinput_f60), .B1(
        BYTEENABLE_REG_2__SCAN_IN), .B2(keyinput_f49), .ZN(n6780) );
  AOI221_X1 U7757 ( .B1(REIP_REG_22__SCAN_IN), .B2(keyinput_f60), .C1(
        keyinput_f49), .C2(BYTEENABLE_REG_2__SCAN_IN), .A(n6780), .ZN(n6785)
         );
  OAI22_X1 U7758 ( .A1(STATEBS16_REG_SCAN_IN), .A2(keyinput_f43), .B1(
        DATAI_28_), .B2(keyinput_f3), .ZN(n6781) );
  AOI221_X1 U7759 ( .B1(STATEBS16_REG_SCAN_IN), .B2(keyinput_f43), .C1(
        keyinput_f3), .C2(DATAI_28_), .A(n6781), .ZN(n6784) );
  OAI22_X1 U7760 ( .A1(REIP_REG_24__SCAN_IN), .A2(keyinput_f58), .B1(
        keyinput_f62), .B2(REIP_REG_20__SCAN_IN), .ZN(n6782) );
  AOI221_X1 U7761 ( .B1(REIP_REG_24__SCAN_IN), .B2(keyinput_f58), .C1(
        REIP_REG_20__SCAN_IN), .C2(keyinput_f62), .A(n6782), .ZN(n6783) );
  NAND4_X1 U7762 ( .A1(n6786), .A2(n6785), .A3(n6784), .A4(n6783), .ZN(n6796)
         );
  OAI22_X1 U7763 ( .A1(keyinput_f95), .A2(ADDRESS_REG_5__SCAN_IN), .B1(
        keyinput_f78), .B2(ADDRESS_REG_22__SCAN_IN), .ZN(n6787) );
  AOI221_X1 U7764 ( .B1(keyinput_f95), .B2(ADDRESS_REG_5__SCAN_IN), .C1(
        ADDRESS_REG_22__SCAN_IN), .C2(keyinput_f78), .A(n6787), .ZN(n6794) );
  OAI22_X1 U7765 ( .A1(keyinput_f123), .A2(DATAWIDTH_REG_19__SCAN_IN), .B1(
        keyinput_f120), .B2(DATAWIDTH_REG_16__SCAN_IN), .ZN(n6788) );
  AOI221_X1 U7766 ( .B1(keyinput_f123), .B2(DATAWIDTH_REG_19__SCAN_IN), .C1(
        DATAWIDTH_REG_16__SCAN_IN), .C2(keyinput_f120), .A(n6788), .ZN(n6793)
         );
  OAI22_X1 U7767 ( .A1(REQUESTPENDING_REG_SCAN_IN), .A2(keyinput_f42), .B1(
        keyinput_f116), .B2(DATAWIDTH_REG_12__SCAN_IN), .ZN(n6789) );
  AOI221_X1 U7768 ( .B1(REQUESTPENDING_REG_SCAN_IN), .B2(keyinput_f42), .C1(
        DATAWIDTH_REG_12__SCAN_IN), .C2(keyinput_f116), .A(n6789), .ZN(n6792)
         );
  OAI22_X1 U7769 ( .A1(STATE_REG_1__SCAN_IN), .A2(keyinput_f102), .B1(DATAI_2_), .B2(keyinput_f29), .ZN(n6790) );
  AOI221_X1 U7770 ( .B1(STATE_REG_1__SCAN_IN), .B2(keyinput_f102), .C1(
        keyinput_f29), .C2(DATAI_2_), .A(n6790), .ZN(n6791) );
  NAND4_X1 U7771 ( .A1(n6794), .A2(n6793), .A3(n6792), .A4(n6791), .ZN(n6795)
         );
  NOR4_X1 U7772 ( .A1(n6798), .A2(n6797), .A3(n6796), .A4(n6795), .ZN(n6895)
         );
  OAI22_X1 U7773 ( .A1(keyinput_f71), .A2(ADDRESS_REG_29__SCAN_IN), .B1(
        keyinput_f33), .B2(NA_N), .ZN(n6799) );
  AOI221_X1 U7774 ( .B1(keyinput_f71), .B2(ADDRESS_REG_29__SCAN_IN), .C1(NA_N), 
        .C2(keyinput_f33), .A(n6799), .ZN(n6806) );
  OAI22_X1 U7775 ( .A1(DATAI_15_), .A2(keyinput_f16), .B1(keyinput_f70), .B2(
        BE_N_REG_0__SCAN_IN), .ZN(n6800) );
  AOI221_X1 U7776 ( .B1(DATAI_15_), .B2(keyinput_f16), .C1(BE_N_REG_0__SCAN_IN), .C2(keyinput_f70), .A(n6800), .ZN(n6805) );
  OAI22_X1 U7777 ( .A1(REIP_REG_18__SCAN_IN), .A2(keyinput_f64), .B1(
        FLUSH_REG_SCAN_IN), .B2(keyinput_f45), .ZN(n6801) );
  AOI221_X1 U7778 ( .B1(REIP_REG_18__SCAN_IN), .B2(keyinput_f64), .C1(
        keyinput_f45), .C2(FLUSH_REG_SCAN_IN), .A(n6801), .ZN(n6804) );
  OAI22_X1 U7779 ( .A1(REIP_REG_21__SCAN_IN), .A2(keyinput_f61), .B1(
        keyinput_f108), .B2(DATAWIDTH_REG_4__SCAN_IN), .ZN(n6802) );
  AOI221_X1 U7780 ( .B1(REIP_REG_21__SCAN_IN), .B2(keyinput_f61), .C1(
        DATAWIDTH_REG_4__SCAN_IN), .C2(keyinput_f108), .A(n6802), .ZN(n6803)
         );
  NAND4_X1 U7781 ( .A1(n6806), .A2(n6805), .A3(n6804), .A4(n6803), .ZN(n6893)
         );
  OAI22_X1 U7782 ( .A1(keyinput_f109), .A2(DATAWIDTH_REG_5__SCAN_IN), .B1(
        keyinput_f67), .B2(BE_N_REG_3__SCAN_IN), .ZN(n6807) );
  AOI221_X1 U7783 ( .B1(keyinput_f109), .B2(DATAWIDTH_REG_5__SCAN_IN), .C1(
        BE_N_REG_3__SCAN_IN), .C2(keyinput_f67), .A(n6807), .ZN(n6817) );
  INV_X1 U7784 ( .A(keyinput_f117), .ZN(n6809) );
  OAI22_X1 U7785 ( .A1(n5371), .A2(keyinput_f66), .B1(n6809), .B2(
        DATAWIDTH_REG_13__SCAN_IN), .ZN(n6808) );
  AOI221_X1 U7786 ( .B1(n5371), .B2(keyinput_f66), .C1(
        DATAWIDTH_REG_13__SCAN_IN), .C2(n6809), .A(n6808), .ZN(n6816) );
  OAI22_X1 U7787 ( .A1(n6811), .A2(keyinput_f22), .B1(n7059), .B2(keyinput_f37), .ZN(n6810) );
  AOI221_X1 U7788 ( .B1(n6811), .B2(keyinput_f22), .C1(keyinput_f37), .C2(
        n7059), .A(n6810), .ZN(n6815) );
  INV_X1 U7789 ( .A(DATAI_20_), .ZN(n6813) );
  OAI22_X1 U7790 ( .A1(n6813), .A2(keyinput_f11), .B1(n7024), .B2(
        keyinput_f124), .ZN(n6812) );
  AOI221_X1 U7791 ( .B1(n6813), .B2(keyinput_f11), .C1(keyinput_f124), .C2(
        n7024), .A(n6812), .ZN(n6814) );
  NAND4_X1 U7792 ( .A1(n6817), .A2(n6816), .A3(n6815), .A4(n6814), .ZN(n6892)
         );
  AOI22_X1 U7793 ( .A1(n6271), .A2(keyinput_f17), .B1(keyinput_f40), .B2(n6903), .ZN(n6818) );
  OAI221_X1 U7794 ( .B1(n6271), .B2(keyinput_f17), .C1(n6903), .C2(
        keyinput_f40), .A(n6818), .ZN(n6829) );
  INV_X1 U7795 ( .A(DATAI_21_), .ZN(n7101) );
  AOI22_X1 U7796 ( .A1(n7101), .A2(keyinput_f10), .B1(keyinput_f79), .B2(n6820), .ZN(n6819) );
  OAI221_X1 U7797 ( .B1(n7101), .B2(keyinput_f10), .C1(n6820), .C2(
        keyinput_f79), .A(n6819), .ZN(n6828) );
  INV_X1 U7798 ( .A(CODEFETCH_REG_SCAN_IN), .ZN(n6822) );
  AOI22_X1 U7799 ( .A1(n6823), .A2(keyinput_f84), .B1(n6822), .B2(keyinput_f39), .ZN(n6821) );
  OAI221_X1 U7800 ( .B1(n6823), .B2(keyinput_f84), .C1(n6822), .C2(
        keyinput_f39), .A(n6821), .ZN(n6827) );
  AOI22_X1 U7801 ( .A1(n6825), .A2(keyinput_f57), .B1(keyinput_f21), .B2(n6261), .ZN(n6824) );
  OAI221_X1 U7802 ( .B1(n6825), .B2(keyinput_f57), .C1(n6261), .C2(
        keyinput_f21), .A(n6824), .ZN(n6826) );
  NOR4_X1 U7803 ( .A1(n6829), .A2(n6828), .A3(n6827), .A4(n6826), .ZN(n6844)
         );
  OAI22_X1 U7804 ( .A1(keyinput_f126), .A2(n6832), .B1(n6831), .B2(
        keyinput_f90), .ZN(n6830) );
  AOI221_X1 U7805 ( .B1(n6832), .B2(keyinput_f126), .C1(n6831), .C2(
        keyinput_f90), .A(n6830), .ZN(n6843) );
  OAI22_X1 U7806 ( .A1(keyinput_f50), .A2(n7015), .B1(n6834), .B2(keyinput_f99), .ZN(n6833) );
  AOI221_X1 U7807 ( .B1(n7015), .B2(keyinput_f50), .C1(n6834), .C2(
        keyinput_f99), .A(n6833), .ZN(n6842) );
  OAI22_X1 U7808 ( .A1(n6836), .A2(keyinput_f93), .B1(n7066), .B2(keyinput_f76), .ZN(n6835) );
  AOI221_X1 U7809 ( .B1(n6836), .B2(keyinput_f93), .C1(keyinput_f76), .C2(
        n7066), .A(n6835), .ZN(n6839) );
  XOR2_X1 U7810 ( .A(n6837), .B(keyinput_f86), .Z(n6838) );
  OAI211_X1 U7811 ( .C1(n7031), .C2(keyinput_f36), .A(n6839), .B(n6838), .ZN(
        n6840) );
  AOI21_X1 U7812 ( .B1(n7031), .B2(keyinput_f36), .A(n6840), .ZN(n6841) );
  NAND4_X1 U7813 ( .A1(n6844), .A2(n6843), .A3(n6842), .A4(n6841), .ZN(n6891)
         );
  INV_X1 U7814 ( .A(keyinput_f119), .ZN(n6846) );
  OAI22_X1 U7815 ( .A1(n7098), .A2(keyinput_f27), .B1(n6846), .B2(
        DATAWIDTH_REG_15__SCAN_IN), .ZN(n6845) );
  AOI221_X1 U7816 ( .B1(n7098), .B2(keyinput_f27), .C1(
        DATAWIDTH_REG_15__SCAN_IN), .C2(n6846), .A(n6845), .ZN(n6889) );
  OAI22_X1 U7817 ( .A1(n7020), .A2(keyinput_f54), .B1(n7006), .B2(
        keyinput_f100), .ZN(n6847) );
  AOI221_X1 U7818 ( .B1(n7020), .B2(keyinput_f54), .C1(keyinput_f100), .C2(
        n7006), .A(n6847), .ZN(n6888) );
  INV_X1 U7819 ( .A(DATAI_29_), .ZN(n6852) );
  OAI22_X1 U7820 ( .A1(n7069), .A2(keyinput_f83), .B1(n7021), .B2(keyinput_f89), .ZN(n6848) );
  AOI221_X1 U7821 ( .B1(n7069), .B2(keyinput_f83), .C1(keyinput_f89), .C2(
        n7021), .A(n6848), .ZN(n6850) );
  XNOR2_X1 U7822 ( .A(keyinput_f107), .B(DATAWIDTH_REG_3__SCAN_IN), .ZN(n6849)
         );
  OAI211_X1 U7823 ( .C1(n6852), .C2(keyinput_f2), .A(n6850), .B(n6849), .ZN(
        n6851) );
  AOI21_X1 U7824 ( .B1(n6852), .B2(keyinput_f2), .A(n6851), .ZN(n6887) );
  INV_X1 U7825 ( .A(DATAI_27_), .ZN(n6965) );
  INV_X1 U7826 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6854) );
  AOI22_X1 U7827 ( .A1(n6965), .A2(keyinput_f4), .B1(keyinput_f104), .B2(n6854), .ZN(n6853) );
  OAI221_X1 U7828 ( .B1(n6965), .B2(keyinput_f4), .C1(n6854), .C2(
        keyinput_f104), .A(n6853), .ZN(n6885) );
  INV_X1 U7829 ( .A(DATAI_31_), .ZN(n6972) );
  AOI22_X1 U7830 ( .A1(n7088), .A2(keyinput_f65), .B1(n6972), .B2(keyinput_f0), 
        .ZN(n6855) );
  OAI221_X1 U7831 ( .B1(n7088), .B2(keyinput_f65), .C1(n6972), .C2(keyinput_f0), .A(n6855), .ZN(n6884) );
  OAI22_X1 U7832 ( .A1(keyinput_f114), .A2(n6986), .B1(n7076), .B2(
        keyinput_f94), .ZN(n6856) );
  AOI221_X1 U7833 ( .B1(n6986), .B2(keyinput_f114), .C1(n7076), .C2(
        keyinput_f94), .A(n6856), .ZN(n6859) );
  XOR2_X1 U7834 ( .A(keyinput_f125), .B(DATAWIDTH_REG_21__SCAN_IN), .Z(n6857)
         );
  AOI21_X1 U7835 ( .B1(keyinput_f56), .B2(n7050), .A(n6857), .ZN(n6858) );
  OAI211_X1 U7836 ( .C1(keyinput_f56), .C2(n7050), .A(n6859), .B(n6858), .ZN(
        n6883) );
  INV_X1 U7837 ( .A(DATAI_17_), .ZN(n6973) );
  OAI22_X1 U7838 ( .A1(n6861), .A2(keyinput_f63), .B1(n6973), .B2(keyinput_f14), .ZN(n6860) );
  AOI221_X1 U7839 ( .B1(n6861), .B2(keyinput_f63), .C1(keyinput_f14), .C2(
        n6973), .A(n6860), .ZN(n6881) );
  XNOR2_X1 U7840 ( .A(keyinput_f118), .B(n7009), .ZN(n6868) );
  XNOR2_X1 U7841 ( .A(keyinput_f113), .B(n7040), .ZN(n6867) );
  AOI22_X1 U7842 ( .A1(n7104), .A2(keyinput_f24), .B1(n7097), .B2(keyinput_f18), .ZN(n6862) );
  OAI221_X1 U7843 ( .B1(n7104), .B2(keyinput_f24), .C1(n7097), .C2(
        keyinput_f18), .A(n6862), .ZN(n6866) );
  INV_X1 U7844 ( .A(DATAI_23_), .ZN(n7072) );
  AOI22_X1 U7845 ( .A1(n6864), .A2(keyinput_f74), .B1(n7072), .B2(keyinput_f8), 
        .ZN(n6863) );
  OAI221_X1 U7846 ( .B1(n6864), .B2(keyinput_f74), .C1(n7072), .C2(keyinput_f8), .A(n6863), .ZN(n6865) );
  NOR4_X1 U7847 ( .A1(n6868), .A2(n6867), .A3(n6866), .A4(n6865), .ZN(n6880)
         );
  OAI22_X1 U7848 ( .A1(keyinput_f106), .A2(n7090), .B1(n6870), .B2(
        keyinput_f69), .ZN(n6869) );
  AOI221_X1 U7849 ( .B1(n7090), .B2(keyinput_f106), .C1(n6870), .C2(
        keyinput_f69), .A(n6869), .ZN(n6879) );
  AOI22_X1 U7850 ( .A1(n6872), .A2(keyinput_f81), .B1(n7030), .B2(keyinput_f55), .ZN(n6871) );
  OAI221_X1 U7851 ( .B1(n6872), .B2(keyinput_f81), .C1(n7030), .C2(
        keyinput_f55), .A(n6871), .ZN(n6877) );
  AOI22_X1 U7852 ( .A1(n4193), .A2(keyinput_f52), .B1(keyinput_f110), .B2(
        n7083), .ZN(n6873) );
  OAI221_X1 U7853 ( .B1(n4193), .B2(keyinput_f52), .C1(n7083), .C2(
        keyinput_f110), .A(n6873), .ZN(n6876) );
  AOI22_X1 U7854 ( .A1(n7023), .A2(keyinput_f92), .B1(n7100), .B2(keyinput_f53), .ZN(n6874) );
  OAI221_X1 U7855 ( .B1(n7023), .B2(keyinput_f92), .C1(n7100), .C2(
        keyinput_f53), .A(n6874), .ZN(n6875) );
  NOR3_X1 U7856 ( .A1(n6877), .A2(n6876), .A3(n6875), .ZN(n6878) );
  NAND4_X1 U7857 ( .A1(n6881), .A2(n6880), .A3(n6879), .A4(n6878), .ZN(n6882)
         );
  NOR4_X1 U7858 ( .A1(n6885), .A2(n6884), .A3(n6883), .A4(n6882), .ZN(n6886)
         );
  NAND4_X1 U7859 ( .A1(n6889), .A2(n6888), .A3(n6887), .A4(n6886), .ZN(n6890)
         );
  NOR4_X1 U7860 ( .A1(n6893), .A2(n6892), .A3(n6891), .A4(n6890), .ZN(n6894)
         );
  NAND4_X1 U7861 ( .A1(n6897), .A2(n6896), .A3(n6895), .A4(n6894), .ZN(n6899)
         );
  AOI21_X1 U7862 ( .B1(keyinput_f28), .B2(n6899), .A(keyinput_g28), .ZN(n6901)
         );
  INV_X1 U7863 ( .A(keyinput_f28), .ZN(n6898) );
  AOI21_X1 U7864 ( .B1(n6899), .B2(n6898), .A(n6902), .ZN(n6900) );
  AOI22_X1 U7865 ( .A1(n6902), .A2(n6901), .B1(keyinput_g28), .B2(n6900), .ZN(
        n7121) );
  XNOR2_X1 U7866 ( .A(n6903), .B(keyinput_g40), .ZN(n6910) );
  AOI22_X1 U7867 ( .A1(ADDRESS_REG_21__SCAN_IN), .A2(keyinput_g79), .B1(
        DATAI_20_), .B2(keyinput_g11), .ZN(n6904) );
  OAI221_X1 U7868 ( .B1(ADDRESS_REG_21__SCAN_IN), .B2(keyinput_g79), .C1(
        DATAI_20_), .C2(keyinput_g11), .A(n6904), .ZN(n6909) );
  AOI22_X1 U7869 ( .A1(ADDRESS_REG_28__SCAN_IN), .A2(keyinput_g72), .B1(
        REIP_REG_23__SCAN_IN), .B2(keyinput_g59), .ZN(n6905) );
  OAI221_X1 U7870 ( .B1(ADDRESS_REG_28__SCAN_IN), .B2(keyinput_g72), .C1(
        REIP_REG_23__SCAN_IN), .C2(keyinput_g59), .A(n6905), .ZN(n6908) );
  AOI22_X1 U7871 ( .A1(ADDRESS_REG_1__SCAN_IN), .A2(keyinput_g99), .B1(
        DATAI_16_), .B2(keyinput_g15), .ZN(n6906) );
  OAI221_X1 U7872 ( .B1(ADDRESS_REG_1__SCAN_IN), .B2(keyinput_g99), .C1(
        DATAI_16_), .C2(keyinput_g15), .A(n6906), .ZN(n6907) );
  NOR4_X1 U7873 ( .A1(n6910), .A2(n6909), .A3(n6908), .A4(n6907), .ZN(n6938)
         );
  AOI22_X1 U7874 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(keyinput_g126), .B1(
        REIP_REG_25__SCAN_IN), .B2(keyinput_g57), .ZN(n6911) );
  OAI221_X1 U7875 ( .B1(DATAWIDTH_REG_22__SCAN_IN), .B2(keyinput_g126), .C1(
        REIP_REG_25__SCAN_IN), .C2(keyinput_g57), .A(n6911), .ZN(n6918) );
  AOI22_X1 U7876 ( .A1(ADDRESS_REG_4__SCAN_IN), .A2(keyinput_g96), .B1(
        DATAI_10_), .B2(keyinput_g21), .ZN(n6912) );
  OAI221_X1 U7877 ( .B1(ADDRESS_REG_4__SCAN_IN), .B2(keyinput_g96), .C1(
        DATAI_10_), .C2(keyinput_g21), .A(n6912), .ZN(n6917) );
  AOI22_X1 U7878 ( .A1(ADS_N_REG_SCAN_IN), .A2(keyinput_g38), .B1(DATAI_29_), 
        .B2(keyinput_g2), .ZN(n6913) );
  OAI221_X1 U7879 ( .B1(ADS_N_REG_SCAN_IN), .B2(keyinput_g38), .C1(DATAI_29_), 
        .C2(keyinput_g2), .A(n6913), .ZN(n6916) );
  AOI22_X1 U7880 ( .A1(BE_N_REG_0__SCAN_IN), .A2(keyinput_g70), .B1(DATAI_9_), 
        .B2(keyinput_g22), .ZN(n6914) );
  OAI221_X1 U7881 ( .B1(BE_N_REG_0__SCAN_IN), .B2(keyinput_g70), .C1(DATAI_9_), 
        .C2(keyinput_g22), .A(n6914), .ZN(n6915) );
  NOR4_X1 U7882 ( .A1(n6918), .A2(n6917), .A3(n6916), .A4(n6915), .ZN(n6937)
         );
  AOI22_X1 U7883 ( .A1(ADDRESS_REG_19__SCAN_IN), .A2(keyinput_g81), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(keyinput_g75), .ZN(n6919) );
  OAI221_X1 U7884 ( .B1(ADDRESS_REG_19__SCAN_IN), .B2(keyinput_g81), .C1(
        ADDRESS_REG_25__SCAN_IN), .C2(keyinput_g75), .A(n6919), .ZN(n6926) );
  AOI22_X1 U7885 ( .A1(BE_N_REG_1__SCAN_IN), .A2(keyinput_g69), .B1(DATAI_22_), 
        .B2(keyinput_g9), .ZN(n6920) );
  OAI221_X1 U7886 ( .B1(BE_N_REG_1__SCAN_IN), .B2(keyinput_g69), .C1(DATAI_22_), .C2(keyinput_g9), .A(n6920), .ZN(n6925) );
  AOI22_X1 U7887 ( .A1(D_C_N_REG_SCAN_IN), .A2(keyinput_g41), .B1(
        CODEFETCH_REG_SCAN_IN), .B2(keyinput_g39), .ZN(n6921) );
  OAI221_X1 U7888 ( .B1(D_C_N_REG_SCAN_IN), .B2(keyinput_g41), .C1(
        CODEFETCH_REG_SCAN_IN), .C2(keyinput_g39), .A(n6921), .ZN(n6924) );
  AOI22_X1 U7889 ( .A1(ADDRESS_REG_20__SCAN_IN), .A2(keyinput_g80), .B1(
        REIP_REG_16__SCAN_IN), .B2(keyinput_g66), .ZN(n6922) );
  OAI221_X1 U7890 ( .B1(ADDRESS_REG_20__SCAN_IN), .B2(keyinput_g80), .C1(
        REIP_REG_16__SCAN_IN), .C2(keyinput_g66), .A(n6922), .ZN(n6923) );
  NOR4_X1 U7891 ( .A1(n6926), .A2(n6925), .A3(n6924), .A4(n6923), .ZN(n6936)
         );
  AOI22_X1 U7892 ( .A1(ADDRESS_REG_16__SCAN_IN), .A2(keyinput_g84), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(keyinput_g88), .ZN(n6927) );
  OAI221_X1 U7893 ( .B1(ADDRESS_REG_16__SCAN_IN), .B2(keyinput_g84), .C1(
        ADDRESS_REG_12__SCAN_IN), .C2(keyinput_g88), .A(n6927), .ZN(n6934) );
  AOI22_X1 U7894 ( .A1(ADDRESS_REG_14__SCAN_IN), .A2(keyinput_g86), .B1(
        DATAWIDTH_REG_23__SCAN_IN), .B2(keyinput_g127), .ZN(n6928) );
  OAI221_X1 U7895 ( .B1(ADDRESS_REG_14__SCAN_IN), .B2(keyinput_g86), .C1(
        DATAWIDTH_REG_23__SCAN_IN), .C2(keyinput_g127), .A(n6928), .ZN(n6933)
         );
  AOI22_X1 U7896 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(keyinput_g125), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(keyinput_g71), .ZN(n6929) );
  OAI221_X1 U7897 ( .B1(DATAWIDTH_REG_21__SCAN_IN), .B2(keyinput_g125), .C1(
        ADDRESS_REG_29__SCAN_IN), .C2(keyinput_g71), .A(n6929), .ZN(n6932) );
  AOI22_X1 U7898 ( .A1(ADDRESS_REG_2__SCAN_IN), .A2(keyinput_g98), .B1(
        DATAI_24_), .B2(keyinput_g7), .ZN(n6930) );
  OAI221_X1 U7899 ( .B1(ADDRESS_REG_2__SCAN_IN), .B2(keyinput_g98), .C1(
        DATAI_24_), .C2(keyinput_g7), .A(n6930), .ZN(n6931) );
  NOR4_X1 U7900 ( .A1(n6934), .A2(n6933), .A3(n6932), .A4(n6931), .ZN(n6935)
         );
  NAND4_X1 U7901 ( .A1(n6938), .A2(n6937), .A3(n6936), .A4(n6935), .ZN(n7119)
         );
  AOI22_X1 U7902 ( .A1(DATAWIDTH_REG_0__SCAN_IN), .A2(keyinput_g104), .B1(
        DATAI_28_), .B2(keyinput_g3), .ZN(n6939) );
  OAI221_X1 U7903 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(keyinput_g104), .C1(
        DATAI_28_), .C2(keyinput_g3), .A(n6939), .ZN(n6946) );
  AOI22_X1 U7904 ( .A1(ADDRESS_REG_13__SCAN_IN), .A2(keyinput_g87), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(keyinput_g85), .ZN(n6940) );
  OAI221_X1 U7905 ( .B1(ADDRESS_REG_13__SCAN_IN), .B2(keyinput_g87), .C1(
        ADDRESS_REG_15__SCAN_IN), .C2(keyinput_g85), .A(n6940), .ZN(n6945) );
  AOI22_X1 U7906 ( .A1(ADDRESS_REG_10__SCAN_IN), .A2(keyinput_g90), .B1(
        BE_N_REG_2__SCAN_IN), .B2(keyinput_g68), .ZN(n6941) );
  OAI221_X1 U7907 ( .B1(ADDRESS_REG_10__SCAN_IN), .B2(keyinput_g90), .C1(
        BE_N_REG_2__SCAN_IN), .C2(keyinput_g68), .A(n6941), .ZN(n6944) );
  AOI22_X1 U7908 ( .A1(ADDRESS_REG_5__SCAN_IN), .A2(keyinput_g95), .B1(
        DATAI_11_), .B2(keyinput_g20), .ZN(n6942) );
  OAI221_X1 U7909 ( .B1(ADDRESS_REG_5__SCAN_IN), .B2(keyinput_g95), .C1(
        DATAI_11_), .C2(keyinput_g20), .A(n6942), .ZN(n6943) );
  NOR4_X1 U7910 ( .A1(n6946), .A2(n6945), .A3(n6944), .A4(n6943), .ZN(n6981)
         );
  AOI22_X1 U7911 ( .A1(ADDRESS_REG_7__SCAN_IN), .A2(keyinput_g93), .B1(
        REIP_REG_21__SCAN_IN), .B2(keyinput_g61), .ZN(n6947) );
  OAI221_X1 U7912 ( .B1(ADDRESS_REG_7__SCAN_IN), .B2(keyinput_g93), .C1(
        REIP_REG_21__SCAN_IN), .C2(keyinput_g61), .A(n6947), .ZN(n6954) );
  AOI22_X1 U7913 ( .A1(ADDRESS_REG_26__SCAN_IN), .A2(keyinput_g74), .B1(
        STATE_REG_2__SCAN_IN), .B2(keyinput_g101), .ZN(n6948) );
  OAI221_X1 U7914 ( .B1(ADDRESS_REG_26__SCAN_IN), .B2(keyinput_g74), .C1(
        STATE_REG_2__SCAN_IN), .C2(keyinput_g101), .A(n6948), .ZN(n6953) );
  AOI22_X1 U7915 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(keyinput_g117), .B1(
        W_R_N_REG_SCAN_IN), .B2(keyinput_g46), .ZN(n6949) );
  OAI221_X1 U7916 ( .B1(DATAWIDTH_REG_13__SCAN_IN), .B2(keyinput_g117), .C1(
        W_R_N_REG_SCAN_IN), .C2(keyinput_g46), .A(n6949), .ZN(n6952) );
  AOI22_X1 U7917 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(keyinput_g119), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(keyinput_g82), .ZN(n6950) );
  OAI221_X1 U7918 ( .B1(DATAWIDTH_REG_15__SCAN_IN), .B2(keyinput_g119), .C1(
        ADDRESS_REG_18__SCAN_IN), .C2(keyinput_g82), .A(n6950), .ZN(n6951) );
  NOR4_X1 U7919 ( .A1(n6954), .A2(n6953), .A3(n6952), .A4(n6951), .ZN(n6980)
         );
  AOI22_X1 U7920 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(keyinput_g107), .B1(
        BE_N_REG_3__SCAN_IN), .B2(keyinput_g67), .ZN(n6955) );
  OAI221_X1 U7921 ( .B1(DATAWIDTH_REG_3__SCAN_IN), .B2(keyinput_g107), .C1(
        BE_N_REG_3__SCAN_IN), .C2(keyinput_g67), .A(n6955), .ZN(n6962) );
  AOI22_X1 U7922 ( .A1(STATE_REG_1__SCAN_IN), .A2(keyinput_g102), .B1(READY_N), 
        .B2(keyinput_g35), .ZN(n6956) );
  OAI221_X1 U7923 ( .B1(STATE_REG_1__SCAN_IN), .B2(keyinput_g102), .C1(READY_N), .C2(keyinput_g35), .A(n6956), .ZN(n6961) );
  AOI22_X1 U7924 ( .A1(DATAI_15_), .A2(keyinput_g16), .B1(REIP_REG_20__SCAN_IN), .B2(keyinput_g62), .ZN(n6957) );
  OAI221_X1 U7925 ( .B1(DATAI_15_), .B2(keyinput_g16), .C1(
        REIP_REG_20__SCAN_IN), .C2(keyinput_g62), .A(n6957), .ZN(n6960) );
  AOI22_X1 U7926 ( .A1(BS16_N), .A2(keyinput_g34), .B1(REIP_REG_19__SCAN_IN), 
        .B2(keyinput_g63), .ZN(n6958) );
  OAI221_X1 U7927 ( .B1(BS16_N), .B2(keyinput_g34), .C1(REIP_REG_19__SCAN_IN), 
        .C2(keyinput_g63), .A(n6958), .ZN(n6959) );
  NOR4_X1 U7928 ( .A1(n6962), .A2(n6961), .A3(n6960), .A4(n6959), .ZN(n6979)
         );
  AOI22_X1 U7929 ( .A1(n6965), .A2(keyinput_g4), .B1(keyinput_g77), .B2(n6964), 
        .ZN(n6963) );
  OAI221_X1 U7930 ( .B1(n6965), .B2(keyinput_g4), .C1(n6964), .C2(keyinput_g77), .A(n6963), .ZN(n6977) );
  AOI22_X1 U7931 ( .A1(n6968), .A2(keyinput_g78), .B1(keyinput_g33), .B2(n6967), .ZN(n6966) );
  OAI221_X1 U7932 ( .B1(n6968), .B2(keyinput_g78), .C1(n6967), .C2(
        keyinput_g33), .A(n6966), .ZN(n6976) );
  AOI22_X1 U7933 ( .A1(n4193), .A2(keyinput_g52), .B1(keyinput_g73), .B2(n6970), .ZN(n6969) );
  OAI221_X1 U7934 ( .B1(n4193), .B2(keyinput_g52), .C1(n6970), .C2(
        keyinput_g73), .A(n6969), .ZN(n6975) );
  AOI22_X1 U7935 ( .A1(n6973), .A2(keyinput_g14), .B1(n6972), .B2(keyinput_g0), 
        .ZN(n6971) );
  OAI221_X1 U7936 ( .B1(n6973), .B2(keyinput_g14), .C1(n6972), .C2(keyinput_g0), .A(n6971), .ZN(n6974) );
  NOR4_X1 U7937 ( .A1(n6977), .A2(n6976), .A3(n6975), .A4(n6974), .ZN(n6978)
         );
  NAND4_X1 U7938 ( .A1(n6981), .A2(n6980), .A3(n6979), .A4(n6978), .ZN(n7118)
         );
  INV_X1 U7939 ( .A(DATAI_18_), .ZN(n6983) );
  AOI22_X1 U7940 ( .A1(n6984), .A2(keyinput_g97), .B1(n6983), .B2(keyinput_g13), .ZN(n6982) );
  OAI221_X1 U7941 ( .B1(n6984), .B2(keyinput_g97), .C1(n6983), .C2(
        keyinput_g13), .A(n6982), .ZN(n6997) );
  INV_X1 U7942 ( .A(DATAI_19_), .ZN(n6987) );
  AOI22_X1 U7943 ( .A1(n6987), .A2(keyinput_g12), .B1(keyinput_g114), .B2(
        n6986), .ZN(n6985) );
  OAI221_X1 U7944 ( .B1(n6987), .B2(keyinput_g12), .C1(n6986), .C2(
        keyinput_g114), .A(n6985), .ZN(n6996) );
  AOI22_X1 U7945 ( .A1(n6990), .A2(keyinput_g111), .B1(n6989), .B2(
        keyinput_g25), .ZN(n6988) );
  OAI221_X1 U7946 ( .B1(n6990), .B2(keyinput_g111), .C1(n6989), .C2(
        keyinput_g25), .A(n6988), .ZN(n6995) );
  AOI22_X1 U7947 ( .A1(n6993), .A2(keyinput_g103), .B1(keyinput_g115), .B2(
        n6992), .ZN(n6991) );
  OAI221_X1 U7948 ( .B1(n6993), .B2(keyinput_g103), .C1(n6992), .C2(
        keyinput_g115), .A(n6991), .ZN(n6994) );
  NOR4_X1 U7949 ( .A1(n6997), .A2(n6996), .A3(n6995), .A4(n6994), .ZN(n7048)
         );
  INV_X1 U7950 ( .A(DATAI_30_), .ZN(n7000) );
  AOI22_X1 U7951 ( .A1(n7000), .A2(keyinput_g1), .B1(n6999), .B2(keyinput_g43), 
        .ZN(n6998) );
  OAI221_X1 U7952 ( .B1(n7000), .B2(keyinput_g1), .C1(n6999), .C2(keyinput_g43), .A(n6998), .ZN(n7013) );
  AOI22_X1 U7953 ( .A1(n7003), .A2(keyinput_g42), .B1(keyinput_g122), .B2(
        n7002), .ZN(n7001) );
  OAI221_X1 U7954 ( .B1(n7003), .B2(keyinput_g42), .C1(n7002), .C2(
        keyinput_g122), .A(n7001), .ZN(n7012) );
  AOI22_X1 U7955 ( .A1(n7006), .A2(keyinput_g100), .B1(n7005), .B2(
        keyinput_g30), .ZN(n7004) );
  OAI221_X1 U7956 ( .B1(n7006), .B2(keyinput_g100), .C1(n7005), .C2(
        keyinput_g30), .A(n7004), .ZN(n7011) );
  AOI22_X1 U7957 ( .A1(n7009), .A2(keyinput_g118), .B1(n7008), .B2(
        keyinput_g23), .ZN(n7007) );
  OAI221_X1 U7958 ( .B1(n7009), .B2(keyinput_g118), .C1(n7008), .C2(
        keyinput_g23), .A(n7007), .ZN(n7010) );
  NOR4_X1 U7959 ( .A1(n7013), .A2(n7012), .A3(n7011), .A4(n7010), .ZN(n7047)
         );
  AOI22_X1 U7960 ( .A1(n7015), .A2(keyinput_g50), .B1(n6271), .B2(keyinput_g17), .ZN(n7014) );
  OAI221_X1 U7961 ( .B1(n7015), .B2(keyinput_g50), .C1(n6271), .C2(
        keyinput_g17), .A(n7014), .ZN(n7028) );
  AOI22_X1 U7962 ( .A1(n7018), .A2(keyinput_g49), .B1(n7017), .B2(keyinput_g58), .ZN(n7016) );
  OAI221_X1 U7963 ( .B1(n7018), .B2(keyinput_g49), .C1(n7017), .C2(
        keyinput_g58), .A(n7016), .ZN(n7027) );
  AOI22_X1 U7964 ( .A1(n7021), .A2(keyinput_g89), .B1(n7020), .B2(keyinput_g54), .ZN(n7019) );
  OAI221_X1 U7965 ( .B1(n7021), .B2(keyinput_g89), .C1(n7020), .C2(
        keyinput_g54), .A(n7019), .ZN(n7026) );
  AOI22_X1 U7966 ( .A1(n7024), .A2(keyinput_g124), .B1(keyinput_g92), .B2(
        n7023), .ZN(n7022) );
  OAI221_X1 U7967 ( .B1(n7024), .B2(keyinput_g124), .C1(n7023), .C2(
        keyinput_g92), .A(n7022), .ZN(n7025) );
  NOR4_X1 U7968 ( .A1(n7028), .A2(n7027), .A3(n7026), .A4(n7025), .ZN(n7046)
         );
  AOI22_X1 U7969 ( .A1(n7031), .A2(keyinput_g36), .B1(n7030), .B2(keyinput_g55), .ZN(n7029) );
  OAI221_X1 U7970 ( .B1(n7031), .B2(keyinput_g36), .C1(n7030), .C2(
        keyinput_g55), .A(n7029), .ZN(n7044) );
  AOI22_X1 U7971 ( .A1(n7034), .A2(keyinput_g48), .B1(n7033), .B2(keyinput_g91), .ZN(n7032) );
  OAI221_X1 U7972 ( .B1(n7034), .B2(keyinput_g48), .C1(n7033), .C2(
        keyinput_g91), .A(n7032), .ZN(n7043) );
  AOI22_X1 U7973 ( .A1(n7037), .A2(keyinput_g121), .B1(n7036), .B2(
        keyinput_g31), .ZN(n7035) );
  OAI221_X1 U7974 ( .B1(n7037), .B2(keyinput_g121), .C1(n7036), .C2(
        keyinput_g31), .A(n7035), .ZN(n7042) );
  INV_X1 U7975 ( .A(MORE_REG_SCAN_IN), .ZN(n7039) );
  AOI22_X1 U7976 ( .A1(n7040), .A2(keyinput_g113), .B1(n7039), .B2(
        keyinput_g44), .ZN(n7038) );
  OAI221_X1 U7977 ( .B1(n7040), .B2(keyinput_g113), .C1(n7039), .C2(
        keyinput_g44), .A(n7038), .ZN(n7041) );
  NOR4_X1 U7978 ( .A1(n7044), .A2(n7043), .A3(n7042), .A4(n7041), .ZN(n7045)
         );
  NAND4_X1 U7979 ( .A1(n7048), .A2(n7047), .A3(n7046), .A4(n7045), .ZN(n7117)
         );
  AOI22_X1 U7980 ( .A1(n7051), .A2(keyinput_g108), .B1(n7050), .B2(
        keyinput_g56), .ZN(n7049) );
  OAI221_X1 U7981 ( .B1(n7051), .B2(keyinput_g108), .C1(n7050), .C2(
        keyinput_g56), .A(n7049), .ZN(n7064) );
  INV_X1 U7982 ( .A(DATAI_25_), .ZN(n7053) );
  AOI22_X1 U7983 ( .A1(n7054), .A2(keyinput_g32), .B1(n7053), .B2(keyinput_g6), 
        .ZN(n7052) );
  OAI221_X1 U7984 ( .B1(n7054), .B2(keyinput_g32), .C1(n7053), .C2(keyinput_g6), .A(n7052), .ZN(n7063) );
  AOI22_X1 U7985 ( .A1(n7057), .A2(keyinput_g123), .B1(keyinput_g120), .B2(
        n7056), .ZN(n7055) );
  OAI221_X1 U7986 ( .B1(n7057), .B2(keyinput_g123), .C1(n7056), .C2(
        keyinput_g120), .A(n7055), .ZN(n7062) );
  AOI22_X1 U7987 ( .A1(n7060), .A2(keyinput_g116), .B1(n7059), .B2(
        keyinput_g37), .ZN(n7058) );
  OAI221_X1 U7988 ( .B1(n7060), .B2(keyinput_g116), .C1(n7059), .C2(
        keyinput_g37), .A(n7058), .ZN(n7061) );
  NOR4_X1 U7989 ( .A1(n7064), .A2(n7063), .A3(n7062), .A4(n7061), .ZN(n7115)
         );
  AOI22_X1 U7990 ( .A1(n7067), .A2(keyinput_g45), .B1(keyinput_g76), .B2(n7066), .ZN(n7065) );
  OAI221_X1 U7991 ( .B1(n7067), .B2(keyinput_g45), .C1(n7066), .C2(
        keyinput_g76), .A(n7065), .ZN(n7080) );
  AOI22_X1 U7992 ( .A1(n7070), .A2(keyinput_g112), .B1(keyinput_g83), .B2(
        n7069), .ZN(n7068) );
  OAI221_X1 U7993 ( .B1(n7070), .B2(keyinput_g112), .C1(n7069), .C2(
        keyinput_g83), .A(n7068), .ZN(n7079) );
  AOI22_X1 U7994 ( .A1(n7073), .A2(keyinput_g64), .B1(keyinput_g8), .B2(n7072), 
        .ZN(n7071) );
  OAI221_X1 U7995 ( .B1(n7073), .B2(keyinput_g64), .C1(n7072), .C2(keyinput_g8), .A(n7071), .ZN(n7078) );
  AOI22_X1 U7996 ( .A1(n7076), .A2(keyinput_g94), .B1(n7075), .B2(
        keyinput_g109), .ZN(n7074) );
  OAI221_X1 U7997 ( .B1(n7076), .B2(keyinput_g94), .C1(n7075), .C2(
        keyinput_g109), .A(n7074), .ZN(n7077) );
  NOR4_X1 U7998 ( .A1(n7080), .A2(n7079), .A3(n7078), .A4(n7077), .ZN(n7114)
         );
  AOI22_X1 U7999 ( .A1(n7083), .A2(keyinput_g110), .B1(n7082), .B2(
        keyinput_g51), .ZN(n7081) );
  OAI221_X1 U8000 ( .B1(n7083), .B2(keyinput_g110), .C1(n7082), .C2(
        keyinput_g51), .A(n7081), .ZN(n7095) );
  INV_X1 U8001 ( .A(DATAI_26_), .ZN(n7085) );
  AOI22_X1 U8002 ( .A1(n7086), .A2(keyinput_g26), .B1(n7085), .B2(keyinput_g5), 
        .ZN(n7084) );
  OAI221_X1 U8003 ( .B1(n7086), .B2(keyinput_g26), .C1(n7085), .C2(keyinput_g5), .A(n7084), .ZN(n7094) );
  AOI22_X1 U8004 ( .A1(n6266), .A2(keyinput_g19), .B1(n7088), .B2(keyinput_g65), .ZN(n7087) );
  OAI221_X1 U8005 ( .B1(n6266), .B2(keyinput_g19), .C1(n7088), .C2(
        keyinput_g65), .A(n7087), .ZN(n7093) );
  AOI22_X1 U8006 ( .A1(n7091), .A2(keyinput_g29), .B1(keyinput_g106), .B2(
        n7090), .ZN(n7089) );
  OAI221_X1 U8007 ( .B1(n7091), .B2(keyinput_g29), .C1(n7090), .C2(
        keyinput_g106), .A(n7089), .ZN(n7092) );
  NOR4_X1 U8008 ( .A1(n7095), .A2(n7094), .A3(n7093), .A4(n7092), .ZN(n7113)
         );
  AOI22_X1 U8009 ( .A1(n7098), .A2(keyinput_g27), .B1(n7097), .B2(keyinput_g18), .ZN(n7096) );
  OAI221_X1 U8010 ( .B1(n7098), .B2(keyinput_g27), .C1(n7097), .C2(
        keyinput_g18), .A(n7096), .ZN(n7111) );
  AOI22_X1 U8011 ( .A1(n7101), .A2(keyinput_g10), .B1(n7100), .B2(keyinput_g53), .ZN(n7099) );
  OAI221_X1 U8012 ( .B1(n7101), .B2(keyinput_g10), .C1(n7100), .C2(
        keyinput_g53), .A(n7099), .ZN(n7110) );
  AOI22_X1 U8013 ( .A1(n7104), .A2(keyinput_g24), .B1(keyinput_g47), .B2(n7103), .ZN(n7102) );
  OAI221_X1 U8014 ( .B1(n7104), .B2(keyinput_g24), .C1(n7103), .C2(
        keyinput_g47), .A(n7102), .ZN(n7109) );
  AOI22_X1 U8015 ( .A1(n7107), .A2(keyinput_g105), .B1(n7106), .B2(
        keyinput_g60), .ZN(n7105) );
  OAI221_X1 U8016 ( .B1(n7107), .B2(keyinput_g105), .C1(n7106), .C2(
        keyinput_g60), .A(n7105), .ZN(n7108) );
  NOR4_X1 U8017 ( .A1(n7111), .A2(n7110), .A3(n7109), .A4(n7108), .ZN(n7112)
         );
  NAND4_X1 U8018 ( .A1(n7115), .A2(n7114), .A3(n7113), .A4(n7112), .ZN(n7116)
         );
  NOR4_X1 U8019 ( .A1(n7119), .A2(n7118), .A3(n7117), .A4(n7116), .ZN(n7120)
         );
  NOR2_X1 U8020 ( .A1(n7121), .A2(n7120), .ZN(n7125) );
  AOI22_X1 U8021 ( .A1(n7123), .A2(BYTEENABLE_REG_3__SCAN_IN), .B1(
        BE_N_REG_3__SCAN_IN), .B2(n7122), .ZN(n7124) );
  XNOR2_X1 U8022 ( .A(n7125), .B(n7124), .ZN(U3445) );
  AND2_X2 U4039 ( .A1(n3185), .A2(n4466), .ZN(n3536) );
  AND2_X2 U3690 ( .A1(n4466), .A2(n4369), .ZN(n3408) );
  NAND2_X1 U4318 ( .A1(n3175), .A2(n3420), .ZN(n3498) );
  AOI21_X1 U3682 ( .B1(n4244), .B2(n6240), .A(n3166), .ZN(n3506) );
  CLKBUF_X1 U3721 ( .A(n3581), .Z(n3162) );
  CLKBUF_X1 U3723 ( .A(n3461), .Z(n3406) );
  CLKBUF_X1 U3775 ( .A(n3553), .Z(n3554) );
  CLKBUF_X1 U3789 ( .A(n3423), .Z(n4305) );
  CLKBUF_X1 U3871 ( .A(n3611), .Z(n5351) );
  CLKBUF_X1 U4296 ( .A(n5340), .Z(n5650) );
  OR2_X1 U4309 ( .A1(n3394), .A2(n3393), .ZN(n5696) );
  CLKBUF_X1 U4417 ( .A(n5559), .Z(n5796) );
  CLKBUF_X1 U4550 ( .A(n5081), .Z(n5116) );
endmodule

