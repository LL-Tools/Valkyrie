

module b14_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, keyinput_128, keyinput_129, 
        keyinput_130, keyinput_131, keyinput_132, keyinput_133, keyinput_134, 
        keyinput_135, keyinput_136, keyinput_137, keyinput_138, keyinput_139, 
        keyinput_140, keyinput_141, keyinput_142, keyinput_143, keyinput_144, 
        keyinput_145, keyinput_146, keyinput_147, keyinput_148, keyinput_149, 
        keyinput_150, keyinput_151, keyinput_152, keyinput_153, keyinput_154, 
        keyinput_155, keyinput_156, keyinput_157, keyinput_158, keyinput_159, 
        keyinput_160, keyinput_161, keyinput_162, keyinput_163, keyinput_164, 
        keyinput_165, keyinput_166, keyinput_167, keyinput_168, keyinput_169, 
        keyinput_170, keyinput_171, keyinput_172, keyinput_173, keyinput_174, 
        keyinput_175, keyinput_176, keyinput_177, keyinput_178, keyinput_179, 
        keyinput_180, keyinput_181, keyinput_182, keyinput_183, keyinput_184, 
        keyinput_185, keyinput_186, keyinput_187, keyinput_188, keyinput_189, 
        keyinput_190, keyinput_191, keyinput_192, keyinput_193, keyinput_194, 
        keyinput_195, keyinput_196, keyinput_197, keyinput_198, keyinput_199, 
        keyinput_200, keyinput_201, keyinput_202, keyinput_203, keyinput_204, 
        keyinput_205, keyinput_206, keyinput_207, keyinput_208, keyinput_209, 
        keyinput_210, keyinput_211, keyinput_212, keyinput_213, keyinput_214, 
        keyinput_215, keyinput_216, keyinput_217, keyinput_218, keyinput_219, 
        keyinput_220, keyinput_221, keyinput_222, keyinput_223, keyinput_224, 
        keyinput_225, keyinput_226, keyinput_227, keyinput_228, keyinput_229, 
        keyinput_230, keyinput_231, keyinput_232, keyinput_233, keyinput_234, 
        keyinput_235, keyinput_236, keyinput_237, keyinput_238, keyinput_239, 
        keyinput_240, keyinput_241, keyinput_242, keyinput_243, keyinput_244, 
        keyinput_245, keyinput_246, keyinput_247, keyinput_248, keyinput_249, 
        keyinput_250, keyinput_251, keyinput_252, keyinput_253, keyinput_254, 
        keyinput_255, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, 
        DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, 
        DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, 
        DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, 
        DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, 
        DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, U3352, U3351, U3350, U3349, 
        U3348, U3347, U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, 
        U3338, U3337, U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, 
        U3328, U3327, U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, 
        U3320, U3319, U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, 
        U3310, U3309, U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, 
        U3300, U3299, U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, 
        U3467, U3469, U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, 
        U3487, U3489, U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, 
        U3506, U3507, U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, 
        U3516, U3517, U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, 
        U3526, U3527, U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, 
        U3536, U3537, U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, 
        U3546, U3547, U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, 
        U3284, U3283, U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, 
        U3274, U3273, U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, 
        U3264, U3263, U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, 
        U3255, U3254, U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, 
        U3245, U3244, U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, 
        U3554, U3555, U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, 
        U3564, U3565, U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, 
        U3574, U3575, U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, 
        U3237, U3236, U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, 
        U3227, U3226, U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, 
        U3217, U3216, U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, 
        U4043 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, keyinput_128, keyinput_129, keyinput_130,
         keyinput_131, keyinput_132, keyinput_133, keyinput_134, keyinput_135,
         keyinput_136, keyinput_137, keyinput_138, keyinput_139, keyinput_140,
         keyinput_141, keyinput_142, keyinput_143, keyinput_144, keyinput_145,
         keyinput_146, keyinput_147, keyinput_148, keyinput_149, keyinput_150,
         keyinput_151, keyinput_152, keyinput_153, keyinput_154, keyinput_155,
         keyinput_156, keyinput_157, keyinput_158, keyinput_159, keyinput_160,
         keyinput_161, keyinput_162, keyinput_163, keyinput_164, keyinput_165,
         keyinput_166, keyinput_167, keyinput_168, keyinput_169, keyinput_170,
         keyinput_171, keyinput_172, keyinput_173, keyinput_174, keyinput_175,
         keyinput_176, keyinput_177, keyinput_178, keyinput_179, keyinput_180,
         keyinput_181, keyinput_182, keyinput_183, keyinput_184, keyinput_185,
         keyinput_186, keyinput_187, keyinput_188, keyinput_189, keyinput_190,
         keyinput_191, keyinput_192, keyinput_193, keyinput_194, keyinput_195,
         keyinput_196, keyinput_197, keyinput_198, keyinput_199, keyinput_200,
         keyinput_201, keyinput_202, keyinput_203, keyinput_204, keyinput_205,
         keyinput_206, keyinput_207, keyinput_208, keyinput_209, keyinput_210,
         keyinput_211, keyinput_212, keyinput_213, keyinput_214, keyinput_215,
         keyinput_216, keyinput_217, keyinput_218, keyinput_219, keyinput_220,
         keyinput_221, keyinput_222, keyinput_223, keyinput_224, keyinput_225,
         keyinput_226, keyinput_227, keyinput_228, keyinput_229, keyinput_230,
         keyinput_231, keyinput_232, keyinput_233, keyinput_234, keyinput_235,
         keyinput_236, keyinput_237, keyinput_238, keyinput_239, keyinput_240,
         keyinput_241, keyinput_242, keyinput_243, keyinput_244, keyinput_245,
         keyinput_246, keyinput_247, keyinput_248, keyinput_249, keyinput_250,
         keyinput_251, keyinput_252, keyinput_253, keyinput_254, keyinput_255,
         DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475,
         n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485,
         n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495,
         n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505,
         n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515,
         n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525,
         n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535,
         n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545,
         n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555,
         n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565,
         n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575,
         n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585,
         n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595,
         n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605,
         n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615,
         n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625,
         n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635,
         n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645,
         n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655,
         n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665,
         n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675,
         n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685,
         n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695,
         n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705,
         n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715,
         n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725,
         n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735,
         n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745,
         n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755,
         n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765,
         n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775,
         n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785,
         n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795,
         n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805,
         n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815,
         n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825,
         n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835,
         n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845,
         n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855,
         n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865,
         n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875,
         n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885,
         n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895,
         n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905,
         n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915,
         n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925,
         n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935,
         n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945,
         n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955,
         n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965,
         n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975,
         n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985,
         n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995,
         n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005,
         n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015,
         n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025,
         n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035,
         n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045,
         n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055,
         n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065,
         n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075,
         n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085,
         n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095,
         n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105,
         n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115,
         n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125,
         n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135,
         n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145,
         n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155,
         n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165,
         n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175,
         n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185,
         n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195,
         n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205,
         n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215,
         n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225,
         n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235,
         n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245,
         n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255,
         n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265,
         n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275,
         n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285,
         n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295,
         n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305,
         n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315,
         n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325,
         n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335,
         n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345,
         n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355,
         n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365,
         n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375,
         n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385,
         n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395,
         n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405,
         n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415,
         n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425,
         n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435,
         n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445,
         n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455,
         n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465,
         n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475,
         n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485,
         n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495,
         n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505,
         n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515,
         n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525,
         n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535,
         n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545,
         n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555,
         n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565,
         n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575,
         n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585,
         n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595,
         n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605,
         n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615,
         n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625,
         n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635,
         n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645,
         n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655,
         n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665,
         n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675,
         n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685,
         n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695,
         n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705,
         n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715,
         n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725,
         n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735,
         n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745,
         n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755,
         n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765,
         n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775,
         n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785,
         n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795,
         n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805,
         n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815,
         n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825,
         n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835,
         n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845,
         n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855,
         n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865,
         n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875,
         n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885,
         n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895,
         n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905,
         n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915,
         n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925,
         n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935,
         n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945,
         n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955,
         n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965,
         n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975,
         n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985,
         n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995,
         n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005,
         n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015,
         n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4026,
         n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036,
         n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046,
         n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056,
         n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066,
         n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076,
         n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086,
         n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096,
         n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106,
         n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116,
         n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126,
         n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136,
         n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146,
         n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156,
         n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166,
         n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176,
         n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186,
         n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196,
         n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206,
         n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216,
         n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226,
         n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236,
         n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246,
         n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256,
         n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266,
         n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276,
         n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286,
         n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296,
         n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306,
         n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316,
         n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326,
         n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336,
         n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346,
         n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356,
         n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366,
         n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376,
         n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386,
         n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396,
         n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406,
         n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416,
         n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426,
         n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436,
         n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446,
         n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456,
         n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466,
         n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476,
         n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486,
         n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496,
         n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506,
         n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516,
         n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526,
         n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536,
         n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546,
         n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556,
         n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
         n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576,
         n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586,
         n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596,
         n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606,
         n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616,
         n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626,
         n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636,
         n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646,
         n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656,
         n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666,
         n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676,
         n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686,
         n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696,
         n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706,
         n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716,
         n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726,
         n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736,
         n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746,
         n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756,
         n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766,
         n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776,
         n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786,
         n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796,
         n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806,
         n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816,
         n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826,
         n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836,
         n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846,
         n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856,
         n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866,
         n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876,
         n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886,
         n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896,
         n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906,
         n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916,
         n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926,
         n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936,
         n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946,
         n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956,
         n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966,
         n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976,
         n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986,
         n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996,
         n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006,
         n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016,
         n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026,
         n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036,
         n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046,
         n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056,
         n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066,
         n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076,
         n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086,
         n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096,
         n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106,
         n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116,
         n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126,
         n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136,
         n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146,
         n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156,
         n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166,
         n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176,
         n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186,
         n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196,
         n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206,
         n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216,
         n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226,
         n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236,
         n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246,
         n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256,
         n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266,
         n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276,
         n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286,
         n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296,
         n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306,
         n5307, n5308, n5309, n5310, n5311;

  BUF_X1 U2503 ( .A(n4969), .Z(n2467) );
  INV_X1 U2504 ( .A(n3327), .ZN(n3859) );
  INV_X1 U2505 ( .A(n2965), .ZN(n3876) );
  INV_X1 U2506 ( .A(n3891), .ZN(n3882) );
  INV_X1 U2507 ( .A(n2935), .ZN(n2466) );
  XNOR2_X2 U2508 ( .A(n2804), .B(n4506), .ZN(n2855) );
  XNOR2_X2 U2509 ( .A(n2754), .B(IR_REG_2__SCAN_IN), .ZN(n5022) );
  AND2_X2 U2510 ( .A1(n2943), .A2(n2959), .ZN(n3327) );
  NAND3_X2 U2511 ( .A1(n4956), .A2(n2879), .A3(n4955), .ZN(n2943) );
  NOR2_X1 U2512 ( .A1(n3864), .A2(n3863), .ZN(n3955) );
  AOI21_X1 U2513 ( .B1(n3965), .B2(n3962), .A(n3961), .ZN(n3932) );
  OR2_X1 U2514 ( .A1(n4063), .A2(n4103), .ZN(n3086) );
  AND2_X2 U2515 ( .A1(n3066), .A2(n5260), .ZN(n5301) );
  CLKBUF_X1 U2516 ( .A(n5003), .Z(n5036) );
  NAND2_X2 U2517 ( .A1(n2972), .A2(n2971), .ZN(n3087) );
  AND4_X1 U2518 ( .A1(n2931), .A2(n2930), .A3(n2929), .A4(n2928), .ZN(n5049)
         );
  AND2_X2 U2520 ( .A1(n2925), .A2(n2926), .ZN(n2966) );
  NAND2_X1 U2521 ( .A1(n4958), .A2(n3077), .ZN(n5283) );
  OR2_X1 U2522 ( .A1(n2873), .A2(n2810), .ZN(n2806) );
  NOR2_X1 U2523 ( .A1(n2711), .A2(n2662), .ZN(n2522) );
  INV_X1 U2524 ( .A(IR_REG_23__SCAN_IN), .ZN(n2797) );
  INV_X1 U2525 ( .A(IR_REG_24__SCAN_IN), .ZN(n4496) );
  INV_X1 U2526 ( .A(IR_REG_11__SCAN_IN), .ZN(n4470) );
  INV_X1 U2527 ( .A(IR_REG_19__SCAN_IN), .ZN(n4485) );
  INV_X1 U2528 ( .A(IR_REG_20__SCAN_IN), .ZN(n4486) );
  XNOR2_X1 U2529 ( .A(n2750), .B(IR_REG_1__SCAN_IN), .ZN(n4969) );
  INV_X1 U2530 ( .A(n2742), .ZN(n2710) );
  INV_X1 U2531 ( .A(IR_REG_6__SCAN_IN), .ZN(n4250) );
  INV_X1 U2532 ( .A(IR_REG_8__SCAN_IN), .ZN(n4255) );
  NAND2_X1 U2533 ( .A1(n4613), .A2(n2849), .ZN(n2850) );
  NAND2_X1 U2534 ( .A1(n2941), .A2(n4957), .ZN(n2959) );
  NAND3_X1 U2535 ( .A1(n4255), .A2(n4250), .A3(n4254), .ZN(n2711) );
  NOR2_X1 U2536 ( .A1(n2586), .A2(n2585), .ZN(n2584) );
  INV_X1 U2537 ( .A(n2592), .ZN(n2585) );
  NAND2_X1 U2538 ( .A1(n4962), .A2(REG1_REG_15__SCAN_IN), .ZN(n2614) );
  NAND2_X1 U2539 ( .A1(n2914), .A2(n4485), .ZN(n2919) );
  INV_X1 U2540 ( .A(n2917), .ZN(n2914) );
  OR2_X1 U2541 ( .A1(n2682), .A2(n2486), .ZN(n2679) );
  AOI21_X1 U2542 ( .B1(n2684), .B2(n2686), .A(n2683), .ZN(n2682) );
  INV_X1 U2543 ( .A(n2687), .ZN(n2684) );
  OR2_X1 U2544 ( .A1(n2685), .A2(n2486), .ZN(n2680) );
  INV_X1 U2545 ( .A(n2686), .ZN(n2685) );
  NOR2_X1 U2546 ( .A1(n2688), .A2(n4068), .ZN(n2687) );
  NOR2_X1 U2547 ( .A1(n2468), .A2(n3669), .ZN(n2688) );
  NAND2_X1 U2548 ( .A1(n2959), .A2(n3070), .ZN(n2575) );
  NAND2_X1 U2549 ( .A1(n4957), .A2(n2576), .ZN(n2974) );
  NAND2_X1 U2550 ( .A1(n5049), .A2(n2973), .ZN(n4108) );
  NAND2_X1 U2551 ( .A1(n2921), .A2(n2924), .ZN(n2926) );
  MUX2_X1 U2552 ( .A(IR_REG_31__SCAN_IN), .B(n2923), .S(IR_REG_29__SCAN_IN), 
        .Z(n2924) );
  AND2_X1 U2553 ( .A1(n2611), .A2(n4265), .ZN(n2610) );
  AOI21_X1 U2554 ( .B1(n4407), .B2(n4408), .A(n2551), .ZN(n2550) );
  XNOR2_X1 U2555 ( .A(n5228), .B(keyinput_13), .ZN(n2551) );
  NAND2_X1 U2556 ( .A1(n4409), .A2(n2548), .ZN(n2547) );
  XNOR2_X1 U2557 ( .A(n4410), .B(n2549), .ZN(n2548) );
  NOR2_X1 U2558 ( .A1(n2545), .A2(n2544), .ZN(n2543) );
  XNOR2_X1 U2559 ( .A(n4428), .B(keyinput_29), .ZN(n2544) );
  NOR2_X1 U2560 ( .A1(n2546), .A2(n4427), .ZN(n2545) );
  AND2_X1 U2561 ( .A1(U3149), .A2(keyinput_32), .ZN(n2542) );
  AOI21_X1 U2562 ( .B1(n2538), .B2(n4475), .A(n2536), .ZN(n2535) );
  INV_X1 U2563 ( .A(n4477), .ZN(n2536) );
  INV_X1 U2564 ( .A(n2538), .ZN(n2537) );
  NAND2_X1 U2565 ( .A1(n2532), .A2(n2497), .ZN(n2531) );
  OAI21_X1 U2566 ( .B1(n4509), .B2(n2534), .A(n2533), .ZN(n2532) );
  INV_X1 U2567 ( .A(IR_REG_16__SCAN_IN), .ZN(n2716) );
  INV_X1 U2568 ( .A(n5193), .ZN(n2593) );
  INV_X1 U2569 ( .A(n2824), .ZN(n2649) );
  INV_X1 U2570 ( .A(n2667), .ZN(n2666) );
  OAI21_X1 U2571 ( .B1(n4739), .B2(n2668), .A(n4667), .ZN(n2667) );
  INV_X1 U2572 ( .A(n4666), .ZN(n2668) );
  AND2_X1 U2573 ( .A1(n4766), .A2(n4682), .ZN(n4748) );
  OR2_X1 U2574 ( .A1(n4779), .A2(n4680), .ZN(n4766) );
  AND2_X1 U2575 ( .A1(n2679), .A2(n2677), .ZN(n2676) );
  INV_X1 U2576 ( .A(n4649), .ZN(n2677) );
  INV_X1 U2577 ( .A(n2659), .ZN(n2658) );
  OAI21_X1 U2578 ( .B1(n3635), .B2(n2660), .A(n2661), .ZN(n2659) );
  NAND2_X1 U2579 ( .A1(n4564), .A2(n3686), .ZN(n2661) );
  INV_X1 U2580 ( .A(n3639), .ZN(n2660) );
  NOR2_X1 U2581 ( .A1(n3548), .A2(n4080), .ZN(n3561) );
  NOR2_X1 U2582 ( .A1(n3274), .A2(n2694), .ZN(n2693) );
  INV_X1 U2583 ( .A(n3247), .ZN(n2694) );
  NAND2_X1 U2584 ( .A1(n2691), .A2(n2693), .ZN(n2690) );
  NAND2_X1 U2585 ( .A1(n3289), .A2(n3244), .ZN(n2691) );
  NAND2_X1 U2586 ( .A1(n2654), .A2(n3112), .ZN(n2652) );
  OAI21_X1 U2587 ( .B1(n2792), .B2(IR_REG_22__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2798) );
  INV_X1 U2588 ( .A(IR_REG_3__SCAN_IN), .ZN(n4456) );
  NAND2_X1 U2589 ( .A1(n3523), .A2(n3522), .ZN(n3524) );
  OR2_X1 U2590 ( .A1(n3313), .A2(n4234), .ZN(n3338) );
  OAI21_X1 U2591 ( .B1(n5236), .B2(n5232), .A(n5233), .ZN(n3752) );
  INV_X1 U2592 ( .A(n3879), .ZN(n3892) );
  OR2_X1 U2593 ( .A1(n2606), .A2(n2603), .ZN(n2602) );
  INV_X1 U2594 ( .A(n2607), .ZN(n2603) );
  AND2_X1 U2595 ( .A1(n3914), .A2(n2608), .ZN(n2606) );
  NAND2_X1 U2596 ( .A1(n2605), .A2(n2607), .ZN(n2604) );
  INV_X1 U2597 ( .A(n3973), .ZN(n2605) );
  NAND2_X1 U2598 ( .A1(n4574), .A2(n3844), .ZN(n2944) );
  AOI21_X1 U2599 ( .B1(n3079), .B2(n3800), .A(n2946), .ZN(n2947) );
  AND2_X1 U2600 ( .A1(n3597), .A2(n2590), .ZN(n2589) );
  NAND2_X1 U2601 ( .A1(n2705), .A2(n2593), .ZN(n2590) );
  NAND2_X1 U2602 ( .A1(n2587), .A2(n2477), .ZN(n2586) );
  NAND2_X1 U2603 ( .A1(n2588), .A2(n5215), .ZN(n2587) );
  NAND2_X2 U2604 ( .A1(n3327), .A2(n3129), .ZN(n3891) );
  NAND2_X1 U2605 ( .A1(n3524), .A2(n3525), .ZN(n3594) );
  NOR2_X1 U2606 ( .A1(n5019), .A2(n2475), .ZN(n2819) );
  NAND2_X1 U2607 ( .A1(n5023), .A2(n2756), .ZN(n2757) );
  NAND2_X1 U2608 ( .A1(n2826), .A2(n2474), .ZN(n2981) );
  NAND2_X1 U2609 ( .A1(n2996), .A2(n2824), .ZN(n2825) );
  NOR2_X1 U2610 ( .A1(n2884), .A2(n2829), .ZN(n2830) );
  AND2_X1 U2611 ( .A1(n3193), .A2(REG2_REG_7__SCAN_IN), .ZN(n2829) );
  OR2_X1 U2612 ( .A1(n3018), .A2(n3440), .ZN(n2644) );
  INV_X1 U2613 ( .A(REG3_REG_10__SCAN_IN), .ZN(n3402) );
  NOR2_X1 U2614 ( .A1(n3055), .A2(n2833), .ZN(n2834) );
  AND2_X1 U2615 ( .A1(n3326), .A2(REG2_REG_9__SCAN_IN), .ZN(n2833) );
  OR2_X1 U2616 ( .A1(n2837), .A2(n4965), .ZN(n2632) );
  NAND2_X1 U2617 ( .A1(n2632), .A2(REG2_REG_12__SCAN_IN), .ZN(n2630) );
  NAND2_X1 U2618 ( .A1(n3477), .A2(n2624), .ZN(n2623) );
  NAND2_X1 U2619 ( .A1(n4966), .A2(REG1_REG_11__SCAN_IN), .ZN(n2624) );
  NOR2_X1 U2620 ( .A1(n4587), .A2(n2620), .ZN(n4585) );
  INV_X1 U2621 ( .A(n2621), .ZN(n2620) );
  AOI21_X1 U2622 ( .B1(n4964), .B2(REG1_REG_13__SCAN_IN), .A(n2775), .ZN(n2621) );
  NAND2_X1 U2623 ( .A1(n2846), .A2(n2845), .ZN(n2629) );
  NAND2_X1 U2624 ( .A1(n2629), .A2(REG2_REG_14__SCAN_IN), .ZN(n2628) );
  INV_X1 U2626 ( .A(n4642), .ZN(n2639) );
  XNOR2_X1 U2627 ( .A(n2850), .B(n4623), .ZN(n4628) );
  AND2_X1 U2628 ( .A1(n2473), .A2(n5297), .ZN(n2558) );
  AND2_X1 U2629 ( .A1(n4729), .A2(n4730), .ZN(n4732) );
  OR2_X1 U2630 ( .A1(n4034), .A2(n4685), .ZN(n4724) );
  AND2_X1 U2631 ( .A1(n3854), .A2(REG3_REG_25__SCAN_IN), .ZN(n3795) );
  OAI21_X1 U2632 ( .B1(n4862), .B2(n2513), .A(n2512), .ZN(n4779) );
  AOI21_X1 U2633 ( .B1(n4678), .B2(n4677), .A(n4679), .ZN(n2512) );
  INV_X1 U2634 ( .A(n4678), .ZN(n2513) );
  OAI21_X1 U2635 ( .B1(n4792), .B2(n4660), .A(n4659), .ZN(n4777) );
  NAND2_X1 U2636 ( .A1(n4838), .A2(n4696), .ZN(n4654) );
  OR2_X1 U2637 ( .A1(n4838), .A2(n4696), .ZN(n4652) );
  AND2_X1 U2638 ( .A1(n4674), .A2(n2516), .ZN(n2515) );
  NAND2_X1 U2639 ( .A1(n4068), .A2(n2517), .ZN(n2516) );
  AND2_X1 U2640 ( .A1(n4013), .A2(n5251), .ZN(n4649) );
  AOI21_X1 U2641 ( .B1(n2687), .B2(n2468), .A(n2487), .ZN(n2686) );
  INV_X1 U2642 ( .A(n5194), .ZN(n3711) );
  NOR2_X1 U2643 ( .A1(n3338), .A2(n3402), .ZN(n3385) );
  NAND2_X1 U2644 ( .A1(n3245), .A2(n2695), .ZN(n3285) );
  INV_X1 U2645 ( .A(n2691), .ZN(n2695) );
  OR2_X1 U2646 ( .A1(n2945), .A2(n5047), .ZN(n3129) );
  AND2_X1 U2647 ( .A1(n4574), .A2(n3079), .ZN(n3107) );
  AND2_X1 U2648 ( .A1(n2974), .A2(n5006), .ZN(n2574) );
  NAND2_X1 U2649 ( .A1(n2967), .A2(REG3_REG_1__SCAN_IN), .ZN(n2930) );
  AND2_X1 U2650 ( .A1(n2943), .A2(n2882), .ZN(n2951) );
  NAND2_X1 U2651 ( .A1(n2880), .A2(n2879), .ZN(n2910) );
  INV_X1 U2652 ( .A(IR_REG_15__SCAN_IN), .ZN(n2722) );
  NAND2_X1 U2653 ( .A1(n4264), .A2(n4470), .ZN(n2714) );
  NAND2_X1 U2654 ( .A1(n2709), .A2(n4259), .ZN(n2662) );
  NOR2_X1 U2655 ( .A1(IR_REG_1__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2752)
         );
  INV_X1 U2656 ( .A(n2580), .ZN(n2579) );
  OAI21_X1 U2657 ( .B1(n3175), .B2(n2581), .A(n3218), .ZN(n2580) );
  AND4_X1 U2658 ( .A1(n3532), .A2(n3531), .A3(n3530), .A4(n3529), .ZN(n3668)
         );
  NAND2_X1 U2659 ( .A1(n3176), .A2(n3175), .ZN(n3231) );
  MUX2_X1 U2660 ( .A(n5022), .B(DATAI_2_), .S(n3025), .Z(n4113) );
  AND4_X1 U2661 ( .A1(n3099), .A2(n3098), .A3(n3097), .A4(n3096), .ZN(n3246)
         );
  INV_X1 U2662 ( .A(n3668), .ZN(n4562) );
  NAND2_X1 U2663 ( .A1(n2966), .A2(REG2_REG_2__SCAN_IN), .ZN(n2972) );
  XNOR2_X1 U2664 ( .A(n2830), .B(n5134), .ZN(n3018) );
  XNOR2_X1 U2665 ( .A(n2623), .B(n2622), .ZN(n4575) );
  NAND2_X1 U2666 ( .A1(n2496), .A2(n2614), .ZN(n2613) );
  NOR2_X1 U2667 ( .A1(n2815), .A2(n2495), .ZN(n5000) );
  NAND2_X1 U2668 ( .A1(n4634), .A2(n2618), .ZN(n2815) );
  NAND2_X1 U2669 ( .A1(n2619), .A2(n2782), .ZN(n2618) );
  NAND2_X1 U2670 ( .A1(n2657), .A2(n3639), .ZN(n3678) );
  NAND2_X1 U2671 ( .A1(n3636), .A2(n3635), .ZN(n2657) );
  INV_X1 U2672 ( .A(keyinput_14), .ZN(n2549) );
  NOR2_X1 U2673 ( .A1(n2550), .A2(n2547), .ZN(n4414) );
  AOI211_X1 U2674 ( .C1(n4425), .C2(n4426), .A(n4424), .B(n4423), .ZN(n2546)
         );
  NOR3_X1 U2675 ( .A1(n2543), .A2(n4430), .A3(n2542), .ZN(n4431) );
  INV_X1 U2676 ( .A(keyinput_184), .ZN(n2626) );
  NAND2_X1 U2677 ( .A1(n2529), .A2(n2527), .ZN(n2526) );
  XNOR2_X1 U2678 ( .A(n4447), .B(n2528), .ZN(n2527) );
  NAND2_X1 U2679 ( .A1(n4445), .A2(n4446), .ZN(n2529) );
  INV_X1 U2680 ( .A(keyinput_50), .ZN(n2528) );
  XNOR2_X1 U2681 ( .A(n2626), .B(IR_REG_1__SCAN_IN), .ZN(n4242) );
  NAND2_X1 U2682 ( .A1(n2525), .A2(n2523), .ZN(n4449) );
  XNOR2_X1 U2683 ( .A(n2524), .B(REG3_REG_20__SCAN_IN), .ZN(n2523) );
  NAND2_X1 U2684 ( .A1(n2526), .A2(n4448), .ZN(n2525) );
  INV_X1 U2685 ( .A(keyinput_53), .ZN(n2524) );
  XNOR2_X1 U2686 ( .A(n2625), .B(IR_REG_1__SCAN_IN), .ZN(n4461) );
  INV_X1 U2687 ( .A(keyinput_56), .ZN(n2625) );
  AND2_X1 U2688 ( .A1(n4474), .A2(n2539), .ZN(n2538) );
  NAND2_X1 U2689 ( .A1(n2541), .A2(n4467), .ZN(n2539) );
  OAI21_X1 U2690 ( .B1(n4468), .B2(n2537), .A(n2535), .ZN(n2540) );
  OR2_X1 U2691 ( .A1(n4508), .A2(n4507), .ZN(n2534) );
  NOR2_X1 U2692 ( .A1(n4512), .A2(n4511), .ZN(n2533) );
  NAND2_X1 U2693 ( .A1(n2703), .A2(n2790), .ZN(n2791) );
  NAND2_X1 U2694 ( .A1(n2701), .A2(n2700), .ZN(n2699) );
  INV_X1 U2695 ( .A(IR_REG_25__SCAN_IN), .ZN(n2700) );
  INV_X1 U2696 ( .A(n2791), .ZN(n2701) );
  AND2_X1 U2697 ( .A1(n2787), .A2(n2611), .ZN(n2566) );
  NOR2_X1 U2698 ( .A1(n2786), .A2(n2785), .ZN(n2787) );
  INV_X1 U2699 ( .A(IR_REG_2__SCAN_IN), .ZN(n4245) );
  XNOR2_X1 U2700 ( .A(n3330), .B(n3892), .ZN(n3371) );
  NAND2_X1 U2701 ( .A1(n3329), .A2(n3328), .ZN(n3330) );
  OR2_X1 U2702 ( .A1(n2702), .A2(n2481), .ZN(n2592) );
  INV_X1 U2703 ( .A(n2594), .ZN(n2588) );
  AOI21_X1 U2704 ( .B1(n2531), .B2(n4534), .A(n2530), .ZN(n4535) );
  OR2_X1 U2705 ( .A1(n4533), .A2(n2498), .ZN(n2530) );
  NAND2_X1 U2706 ( .A1(n2887), .A2(n2769), .ZN(n2770) );
  NOR2_X1 U2707 ( .A1(n4723), .A2(n4685), .ZN(n4710) );
  INV_X1 U2708 ( .A(n4146), .ZN(n4683) );
  AND2_X1 U2709 ( .A1(n4012), .A2(n4011), .ZN(n4678) );
  INV_X1 U2710 ( .A(n4005), .ZN(n2517) );
  AND2_X1 U2711 ( .A1(n3778), .A2(n5266), .ZN(n2565) );
  NOR2_X1 U2712 ( .A1(n4877), .A2(n5217), .ZN(n3779) );
  NAND2_X1 U2713 ( .A1(n3569), .A2(n2569), .ZN(n3652) );
  AND2_X1 U2714 ( .A1(n2570), .A2(n3687), .ZN(n2569) );
  AND2_X1 U2715 ( .A1(n3568), .A2(n3637), .ZN(n2570) );
  INV_X1 U2716 ( .A(REG3_REG_9__SCAN_IN), .ZN(n4234) );
  NOR2_X1 U2717 ( .A1(n3187), .A2(n3186), .ZN(n3204) );
  OAI21_X1 U2718 ( .B1(n3086), .B2(n2506), .A(n2503), .ZN(n5078) );
  AND2_X1 U2719 ( .A1(n2504), .A2(n4107), .ZN(n2503) );
  NAND2_X1 U2720 ( .A1(n4075), .A2(n2505), .ZN(n2504) );
  INV_X1 U2721 ( .A(n4108), .ZN(n2505) );
  NAND2_X1 U2722 ( .A1(n5078), .A2(n5079), .ZN(n5077) );
  NOR2_X1 U2723 ( .A1(n3287), .A2(n3286), .ZN(n3248) );
  AND3_X1 U2724 ( .A1(n2697), .A2(n2713), .A3(n2566), .ZN(n2873) );
  NOR2_X1 U2725 ( .A1(n2699), .A2(n2698), .ZN(n2697) );
  NAND2_X1 U2726 ( .A1(n4285), .A2(n2788), .ZN(n2698) );
  INV_X1 U2727 ( .A(IR_REG_21__SCAN_IN), .ZN(n2788) );
  INV_X1 U2728 ( .A(IR_REG_14__SCAN_IN), .ZN(n4269) );
  INV_X1 U2729 ( .A(IR_REG_12__SCAN_IN), .ZN(n4264) );
  INV_X1 U2730 ( .A(IR_REG_9__SCAN_IN), .ZN(n4259) );
  NOR2_X1 U2731 ( .A1(n2711), .A2(IR_REG_5__SCAN_IN), .ZN(n2663) );
  INV_X2 U2732 ( .A(IR_REG_7__SCAN_IN), .ZN(n4254) );
  AND2_X1 U2733 ( .A1(n3154), .A2(n3177), .ZN(n2578) );
  NAND2_X1 U2734 ( .A1(n3731), .A2(n2595), .ZN(n2594) );
  INV_X1 U2735 ( .A(n3733), .ZN(n2595) );
  NAND2_X1 U2736 ( .A1(n2591), .A2(n2589), .ZN(n3732) );
  NAND2_X1 U2737 ( .A1(n3594), .A2(n2592), .ZN(n2591) );
  NAND2_X1 U2738 ( .A1(n2601), .A2(n2599), .ZN(n3949) );
  AOI21_X1 U2739 ( .B1(n2602), .B2(n2604), .A(n2600), .ZN(n2599) );
  INV_X1 U2740 ( .A(n3863), .ZN(n2600) );
  AND2_X1 U2741 ( .A1(n3949), .A2(n3954), .ZN(n3951) );
  OR2_X1 U2742 ( .A1(n3838), .A2(n4381), .ZN(n3852) );
  NAND2_X1 U2743 ( .A1(n3155), .A2(n3154), .ZN(n3176) );
  NOR2_X1 U2744 ( .A1(n3757), .A2(n3756), .ZN(n3819) );
  OR2_X1 U2745 ( .A1(n3972), .A2(n3973), .ZN(n2609) );
  NAND2_X1 U2746 ( .A1(n3368), .A2(n3376), .ZN(n3419) );
  OR2_X1 U2747 ( .A1(n3358), .A2(n3357), .ZN(n3359) );
  XNOR2_X1 U2748 ( .A(n3028), .B(n3879), .ZN(n3030) );
  NAND2_X1 U2749 ( .A1(n3030), .A2(n3029), .ZN(n3142) );
  INV_X1 U2750 ( .A(n3718), .ZN(n3741) );
  INV_X1 U2751 ( .A(n4865), .ZN(n4651) );
  NAND2_X1 U2752 ( .A1(n3941), .A2(n3942), .ZN(n3940) );
  NOR2_X1 U2753 ( .A1(n3466), .A2(n3527), .ZN(n3528) );
  NAND2_X1 U2754 ( .A1(n3594), .A2(n2702), .ZN(n5188) );
  XNOR2_X1 U2755 ( .A(REG0_REG_3__SCAN_IN), .B(keyinput_122), .ZN(n2553) );
  AND4_X1 U2756 ( .A1(n3607), .A2(n3606), .A3(n3605), .A4(n3604), .ZN(n3777)
         );
  AND4_X1 U2757 ( .A1(n3589), .A2(n3588), .A3(n3587), .A4(n3586), .ZN(n4888)
         );
  AND4_X1 U2758 ( .A1(n3391), .A2(n3390), .A3(n3389), .A4(n3388), .ZN(n3638)
         );
  AND4_X1 U2759 ( .A1(n3343), .A2(n3342), .A3(n3341), .A4(n3340), .ZN(n3536)
         );
  AND4_X1 U2760 ( .A1(n3093), .A2(n3092), .A3(n3091), .A4(n3090), .ZN(n3923)
         );
  NAND2_X1 U2761 ( .A1(n5024), .A2(n5025), .ZN(n5023) );
  OR2_X1 U2762 ( .A1(n2999), .A2(n2998), .ZN(n2996) );
  OAI21_X1 U2763 ( .B1(n5117), .B2(n3006), .A(n3001), .ZN(n2762) );
  OAI21_X1 U2764 ( .B1(n2648), .B2(n2469), .A(n2646), .ZN(n2827) );
  AOI21_X1 U2765 ( .B1(n2822), .B2(n2647), .A(n2483), .ZN(n2646) );
  OR2_X1 U2766 ( .A1(n3483), .A2(n3482), .ZN(n3480) );
  NAND2_X1 U2767 ( .A1(n2631), .A2(n2630), .ZN(n4590) );
  AND2_X1 U2768 ( .A1(n2628), .A2(n2627), .ZN(n4616) );
  OR2_X1 U2769 ( .A1(n4616), .A2(n4615), .ZN(n4613) );
  AND2_X1 U2770 ( .A1(n2612), .A2(n2614), .ZN(n2780) );
  NAND2_X1 U2771 ( .A1(n2780), .A2(n4623), .ZN(n2781) );
  INV_X1 U2772 ( .A(n2640), .ZN(n2637) );
  NAND2_X1 U2773 ( .A1(n4960), .A2(REG2_REG_17__SCAN_IN), .ZN(n2640) );
  NOR2_X1 U2774 ( .A1(n2480), .A2(n2597), .ZN(n2596) );
  INV_X1 U2775 ( .A(n2717), .ZN(n2597) );
  NOR2_X1 U2776 ( .A1(n5229), .A2(n5248), .ZN(n2617) );
  NOR2_X1 U2777 ( .A1(n4710), .A2(n4709), .ZN(n4708) );
  AND2_X1 U2778 ( .A1(n4710), .A2(n4709), .ZN(n2511) );
  INV_X1 U2779 ( .A(n4711), .ZN(n2509) );
  AND2_X1 U2780 ( .A1(n4732), .A2(n4713), .ZN(n4715) );
  OR2_X1 U2781 ( .A1(n4033), .A2(n4686), .ZN(n4709) );
  NAND2_X1 U2782 ( .A1(n2665), .A2(n2664), .ZN(n4706) );
  AOI21_X1 U2783 ( .B1(n2666), .B2(n2668), .A(n2484), .ZN(n2664) );
  OAI21_X1 U2784 ( .B1(n4748), .B2(n4684), .A(n4683), .ZN(n4725) );
  INV_X1 U2785 ( .A(n4753), .ZN(n4741) );
  OR2_X1 U2786 ( .A1(n4748), .A2(n4747), .ZN(n4750) );
  NOR2_X1 U2787 ( .A1(n4048), .A2(n4784), .ZN(n2568) );
  AOI22_X1 U2788 ( .A1(n4777), .A2(n4663), .B1(n4662), .B2(n4661), .ZN(n4759)
         );
  INV_X1 U2789 ( .A(n4661), .ZN(n4784) );
  NAND2_X1 U2790 ( .A1(n4812), .A2(n2568), .ZN(n4785) );
  NAND2_X1 U2791 ( .A1(n4812), .A2(n4802), .ZN(n4793) );
  AND2_X1 U2792 ( .A1(n4845), .A2(n4828), .ZN(n4812) );
  AOI21_X1 U2793 ( .B1(n2470), .B2(n2671), .A(n2485), .ZN(n2670) );
  INV_X1 U2794 ( .A(n4656), .ZN(n2671) );
  AND2_X1 U2795 ( .A1(n3779), .A2(n2564), .ZN(n4845) );
  AND2_X1 U2796 ( .A1(n2471), .A2(n4847), .ZN(n2564) );
  NAND2_X1 U2797 ( .A1(n4676), .A2(n4856), .ZN(n4862) );
  NAND2_X1 U2798 ( .A1(n3779), .A2(n2471), .ZN(n4867) );
  NAND2_X1 U2799 ( .A1(n3779), .A2(n2565), .ZN(n5265) );
  AND2_X1 U2800 ( .A1(n4044), .A2(n4043), .ZN(n4856) );
  NAND2_X1 U2801 ( .A1(n2675), .A2(n2674), .ZN(n5264) );
  AOI21_X1 U2802 ( .B1(n2676), .B2(n2680), .A(n2488), .ZN(n2674) );
  INV_X1 U2803 ( .A(n5238), .ZN(n3778) );
  NAND2_X1 U2804 ( .A1(n2514), .A2(n4068), .ZN(n4882) );
  NAND2_X1 U2805 ( .A1(n3705), .A2(n4005), .ZN(n2514) );
  OR2_X1 U2806 ( .A1(n3710), .A2(n3774), .ZN(n4877) );
  NAND2_X1 U2807 ( .A1(n4007), .A2(n4078), .ZN(n3660) );
  AOI21_X1 U2808 ( .B1(n2658), .B2(n2660), .A(n2489), .ZN(n2656) );
  NOR2_X1 U2809 ( .A1(n3652), .A2(n3665), .ZN(n3712) );
  OAI21_X1 U2810 ( .B1(n3552), .B2(n2502), .A(n2500), .ZN(n4007) );
  AND2_X1 U2811 ( .A1(n2501), .A2(n4099), .ZN(n2500) );
  NAND2_X1 U2812 ( .A1(n4096), .A2(n3544), .ZN(n2501) );
  AND2_X1 U2813 ( .A1(n3385), .A2(n3384), .ZN(n3425) );
  NAND2_X1 U2814 ( .A1(n3569), .A2(n2570), .ZN(n3685) );
  NAND2_X1 U2815 ( .A1(n3569), .A2(n3568), .ZN(n3623) );
  AND2_X1 U2816 ( .A1(n3563), .A2(n3562), .ZN(n3628) );
  AND2_X1 U2817 ( .A1(n3616), .A2(n3644), .ZN(n4077) );
  AND2_X1 U2818 ( .A1(n3501), .A2(n3500), .ZN(n3569) );
  NAND2_X1 U2819 ( .A1(n3552), .A2(n4080), .ZN(n3646) );
  OR2_X1 U2820 ( .A1(n3542), .A2(n3541), .ZN(n3548) );
  AOI21_X1 U2821 ( .B1(n3491), .B2(n4126), .A(n4124), .ZN(n3493) );
  NOR2_X1 U2822 ( .A1(n3437), .A2(n3438), .ZN(n3501) );
  NAND2_X1 U2823 ( .A1(n3290), .A2(n4118), .ZN(n3266) );
  AND2_X1 U2824 ( .A1(n2690), .A2(n2696), .ZN(n2689) );
  INV_X1 U2825 ( .A(n2693), .ZN(n2692) );
  OR2_X1 U2826 ( .A1(n3273), .A2(n3272), .ZN(n2696) );
  NAND2_X1 U2827 ( .A1(n3248), .A2(n3272), .ZN(n3277) );
  NAND2_X1 U2828 ( .A1(n2555), .A2(n3267), .ZN(n3437) );
  INV_X1 U2829 ( .A(n3277), .ZN(n2555) );
  INV_X1 U2830 ( .A(n3271), .ZN(n3272) );
  NAND2_X1 U2831 ( .A1(n3095), .A2(REG3_REG_5__SCAN_IN), .ZN(n3187) );
  NAND2_X1 U2832 ( .A1(n3237), .A2(n4079), .ZN(n2521) );
  NAND2_X1 U2833 ( .A1(n2521), .A2(n2519), .ZN(n3290) );
  NOR2_X1 U2834 ( .A1(n3289), .A2(n2520), .ZN(n2519) );
  INV_X1 U2835 ( .A(n4115), .ZN(n2520) );
  OR2_X1 U2836 ( .A1(n5087), .A2(n3243), .ZN(n3287) );
  AND2_X1 U2837 ( .A1(n2652), .A2(n3113), .ZN(n2651) );
  INV_X1 U2838 ( .A(n5048), .ZN(n4839) );
  AND2_X1 U2839 ( .A1(n4115), .A2(n4117), .ZN(n4079) );
  NAND2_X1 U2840 ( .A1(n2561), .A2(n2563), .ZN(n5087) );
  NOR2_X1 U2841 ( .A1(n2562), .A2(n5090), .ZN(n2561) );
  NAND2_X1 U2842 ( .A1(n4063), .A2(n3107), .ZN(n3109) );
  NAND2_X1 U2843 ( .A1(n2563), .A2(n2560), .ZN(n5089) );
  INV_X1 U2844 ( .A(n2562), .ZN(n2560) );
  INV_X1 U2845 ( .A(n2973), .ZN(n3080) );
  AND3_X1 U2846 ( .A1(n4905), .A2(n4904), .A3(n4903), .ZN(n4941) );
  NAND2_X1 U2847 ( .A1(n2805), .A2(n2807), .ZN(n4989) );
  OR2_X1 U2848 ( .A1(n2806), .A2(n4505), .ZN(n2807) );
  INV_X1 U2849 ( .A(IR_REG_22__SCAN_IN), .ZN(n2790) );
  NAND2_X1 U2850 ( .A1(n2919), .A2(IR_REG_31__SCAN_IN), .ZN(n2915) );
  NAND2_X1 U2851 ( .A1(n2720), .A2(n2717), .ZN(n2912) );
  NAND2_X1 U2852 ( .A1(n2713), .A2(n2712), .ZN(n2727) );
  NOR2_X1 U2853 ( .A1(IR_REG_2__SCAN_IN), .A2(IR_REG_1__SCAN_IN), .ZN(n2573)
         );
  NOR2_X1 U2854 ( .A1(IR_REG_4__SCAN_IN), .A2(IR_REG_3__SCAN_IN), .ZN(n2572)
         );
  AND2_X1 U2855 ( .A1(n2749), .A2(n2748), .ZN(n3088) );
  AND2_X1 U2856 ( .A1(n3885), .A2(n3871), .ZN(n4733) );
  AND2_X1 U2857 ( .A1(n2609), .A2(n2608), .ZN(n3915) );
  AND4_X1 U2858 ( .A1(n3353), .A2(n3352), .A3(n3351), .A4(n3350), .ZN(n3630)
         );
  NAND2_X1 U2859 ( .A1(n3732), .A2(n2594), .ZN(n5216) );
  NAND2_X1 U2860 ( .A1(n4000), .A2(DATAI_24_), .ZN(n4661) );
  NAND2_X1 U2861 ( .A1(n2598), .A2(n2602), .ZN(n3864) );
  INV_X1 U2862 ( .A(n3498), .ZN(n3500) );
  NAND2_X1 U2863 ( .A1(n4000), .A2(DATAI_22_), .ZN(n4828) );
  INV_X1 U2864 ( .A(n5244), .ZN(n3980) );
  INV_X1 U2865 ( .A(n3576), .ZN(n3629) );
  NAND2_X1 U2866 ( .A1(n2583), .A2(n2582), .ZN(n5236) );
  OR2_X1 U2867 ( .A1(n2479), .A2(n2586), .ZN(n2582) );
  NAND2_X1 U2868 ( .A1(n3594), .A2(n2584), .ZN(n2583) );
  AND4_X1 U2869 ( .A1(n3192), .A2(n3191), .A3(n3190), .A4(n3189), .ZN(n3319)
         );
  NAND2_X1 U2870 ( .A1(n3231), .A2(n3177), .ZN(n3217) );
  INV_X1 U2871 ( .A(n5192), .ZN(n5239) );
  AND2_X1 U2872 ( .A1(n3596), .A2(n3595), .ZN(n5193) );
  INV_X1 U2873 ( .A(n3403), .ZN(n5231) );
  OAI21_X1 U2874 ( .B1(n2554), .B2(n2499), .A(n2552), .ZN(n4555) );
  AND2_X1 U2875 ( .A1(n4553), .A2(n4552), .ZN(n2552) );
  AOI211_X1 U2876 ( .C1(n4547), .C2(n4548), .A(n4546), .B(n4545), .ZN(n2554)
         );
  INV_X1 U2877 ( .A(n4886), .ZN(n4648) );
  NAND2_X1 U2878 ( .A1(n3209), .A2(n2706), .ZN(n4568) );
  NAND4_X1 U2879 ( .A1(n3048), .A2(n3047), .A3(n3046), .A4(n3045), .ZN(n4573)
         );
  NAND2_X1 U2880 ( .A1(n2940), .A2(n2939), .ZN(n4574) );
  AND3_X1 U2881 ( .A1(n2938), .A2(n2937), .A3(n2936), .ZN(n2940) );
  INV_X1 U2882 ( .A(U4043), .ZN(n5017) );
  AND2_X1 U2883 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n2708)
         );
  XNOR2_X1 U2884 ( .A(n2757), .B(n5075), .ZN(n3011) );
  NAND2_X1 U2885 ( .A1(n3011), .A2(REG1_REG_3__SCAN_IN), .ZN(n3010) );
  INV_X1 U2886 ( .A(n2644), .ZN(n3017) );
  OAI21_X1 U2887 ( .B1(n3018), .B2(n2642), .A(n2641), .ZN(n3055) );
  NAND2_X1 U2888 ( .A1(n2645), .A2(REG2_REG_8__SCAN_IN), .ZN(n2642) );
  INV_X1 U2889 ( .A(n3056), .ZN(n2645) );
  INV_X1 U2890 ( .A(n2831), .ZN(n2643) );
  NOR2_X1 U2891 ( .A1(n2630), .A2(n2838), .ZN(n4579) );
  AOI21_X1 U2892 ( .B1(n4575), .B2(REG1_REG_12__SCAN_IN), .A(n2476), .ZN(n4587) );
  NAND2_X1 U2893 ( .A1(n2627), .A2(n2629), .ZN(n4604) );
  NOR2_X1 U2894 ( .A1(n2628), .A2(n2847), .ZN(n4603) );
  AOI22_X1 U2895 ( .A1(n4600), .A2(REG1_REG_14__SCAN_IN), .B1(n2777), .B2(
        n4963), .ZN(n4611) );
  OAI21_X1 U2896 ( .B1(n2780), .B2(n4623), .A(n2781), .ZN(n4622) );
  NAND2_X1 U2897 ( .A1(n4626), .A2(n2851), .ZN(n4641) );
  INV_X1 U2898 ( .A(n4626), .ZN(n2633) );
  NAND2_X1 U2899 ( .A1(n4628), .A2(n2636), .ZN(n2635) );
  NOR2_X1 U2900 ( .A1(n2637), .A2(REG2_REG_16__SCAN_IN), .ZN(n2636) );
  INV_X1 U2901 ( .A(n4632), .ZN(n5038) );
  XNOR2_X1 U2902 ( .A(n2616), .B(n2615), .ZN(n5008) );
  INV_X1 U2903 ( .A(n5002), .ZN(n2615) );
  NOR2_X1 U2904 ( .A1(n5000), .A2(n2617), .ZN(n2616) );
  OR2_X1 U2905 ( .A1(n2473), .A2(n5297), .ZN(n2556) );
  NAND2_X1 U2906 ( .A1(n4732), .A2(n2558), .ZN(n2557) );
  OR2_X1 U2907 ( .A1(n4732), .A2(n5297), .ZN(n2559) );
  AOI21_X1 U2908 ( .B1(n2510), .B2(n5256), .A(n2507), .ZN(n4910) );
  NAND2_X1 U2909 ( .A1(n2509), .A2(n2508), .ZN(n2507) );
  OR2_X1 U2910 ( .A1(n2511), .A2(n4708), .ZN(n2510) );
  NAND2_X1 U2911 ( .A1(n4712), .A2(n4839), .ZN(n2508) );
  NAND2_X1 U2912 ( .A1(n4738), .A2(n4666), .ZN(n4721) );
  NAND2_X1 U2913 ( .A1(n4812), .A2(n2567), .ZN(n4921) );
  AND2_X1 U2914 ( .A1(n2568), .A2(n4772), .ZN(n2567) );
  NAND2_X1 U2915 ( .A1(n2672), .A2(n2470), .ZN(n4810) );
  NAND2_X1 U2916 ( .A1(n2673), .A2(n4656), .ZN(n2672) );
  NAND2_X1 U2917 ( .A1(n2678), .A2(n2679), .ZN(n4650) );
  OR2_X1 U2918 ( .A1(n3701), .A2(n2680), .ZN(n2678) );
  NAND2_X1 U2919 ( .A1(n2681), .A2(n2686), .ZN(n4880) );
  NAND2_X1 U2920 ( .A1(n3701), .A2(n2687), .ZN(n2681) );
  AOI21_X1 U2921 ( .B1(n3701), .B2(n3669), .A(n2468), .ZN(n3775) );
  NAND2_X1 U2922 ( .A1(n2575), .A2(n2974), .ZN(n3690) );
  NAND2_X1 U2923 ( .A1(n3285), .A2(n3247), .ZN(n3275) );
  AND2_X1 U2924 ( .A1(n5258), .A2(n3118), .ZN(n5268) );
  INV_X1 U2925 ( .A(n4897), .ZN(n5298) );
  NAND2_X1 U2926 ( .A1(n3086), .A2(n4108), .ZN(n3121) );
  NAND2_X1 U2927 ( .A1(n2951), .A2(n2933), .ZN(n5260) );
  NOR2_X1 U2928 ( .A1(n4900), .A2(n4899), .ZN(n4901) );
  NAND2_X1 U2929 ( .A1(n2921), .A2(IR_REG_31__SCAN_IN), .ZN(n2875) );
  XNOR2_X1 U2930 ( .A(n2789), .B(IR_REG_24__SCAN_IN), .ZN(n4956) );
  AND2_X1 U2931 ( .A1(n2778), .A2(n2724), .ZN(n4962) );
  AND2_X1 U2932 ( .A1(n2713), .A2(n2611), .ZN(n2725) );
  NAND2_X1 U2933 ( .A1(n2753), .A2(IR_REG_31__SCAN_IN), .ZN(n2754) );
  INV_X1 U2934 ( .A(n2752), .ZN(n2753) );
  NOR2_X4 U2935 ( .A1(n2927), .A2(n2926), .ZN(n2967) );
  AND2_X1 U2936 ( .A1(n3668), .A2(n3711), .ZN(n2468) );
  XNOR2_X1 U2937 ( .A(n3087), .B(n4113), .ZN(n4075) );
  INV_X1 U2938 ( .A(n4075), .ZN(n2506) );
  OR2_X1 U2939 ( .A1(n2813), .A2(n2812), .ZN(n4089) );
  OR2_X1 U2940 ( .A1(n2998), .A2(n2650), .ZN(n2469) );
  AOI21_X1 U2942 ( .B1(n3594), .B2(n3593), .A(n2705), .ZN(n3598) );
  AND2_X1 U2943 ( .A1(n2482), .A2(n4811), .ZN(n2470) );
  AND2_X1 U2944 ( .A1(n2565), .A2(n4868), .ZN(n2471) );
  MUX2_X1 U2945 ( .A(n4963), .B(DATAI_14_), .S(n3025), .Z(n3665) );
  AND2_X1 U2946 ( .A1(n4698), .A2(n4713), .ZN(n2472) );
  AND2_X1 U2947 ( .A1(n2472), .A2(n5295), .ZN(n2473) );
  NAND2_X2 U2948 ( .A1(n2943), .A2(n2942), .ZN(n2965) );
  NAND2_X1 U2949 ( .A1(n2710), .A2(n2709), .ZN(n2740) );
  NAND4_X1 U2950 ( .A1(n3318), .A2(n3317), .A3(n3316), .A4(n3315), .ZN(n3325)
         );
  OR2_X1 U2951 ( .A1(n2825), .A2(n4967), .ZN(n2474) );
  AND2_X1 U2952 ( .A1(n5022), .A2(REG2_REG_2__SCAN_IN), .ZN(n2475) );
  NOR2_X1 U2953 ( .A1(n2792), .A2(n2699), .ZN(n2803) );
  AND2_X1 U2954 ( .A1(n2623), .A2(n4965), .ZN(n2476) );
  AND2_X1 U2955 ( .A1(n2713), .A2(n2566), .ZN(n2809) );
  AND2_X1 U2956 ( .A1(n2710), .A2(n2663), .ZN(n2735) );
  NAND2_X1 U2957 ( .A1(n3740), .A2(n3739), .ZN(n2477) );
  OR2_X1 U2958 ( .A1(n2792), .A2(n2791), .ZN(n2478) );
  INV_X1 U2959 ( .A(IR_REG_10__SCAN_IN), .ZN(n2712) );
  NAND2_X1 U2960 ( .A1(n4628), .A2(n4627), .ZN(n4626) );
  AND2_X1 U2961 ( .A1(n2589), .A2(n5215), .ZN(n2479) );
  NOR2_X1 U2962 ( .A1(n2913), .A2(n2810), .ZN(n2480) );
  INV_X1 U2963 ( .A(n5006), .ZN(n4959) );
  NAND2_X1 U2964 ( .A1(n2919), .A2(n2918), .ZN(n5006) );
  AND2_X1 U2965 ( .A1(n3593), .A2(n2593), .ZN(n2481) );
  INV_X1 U2966 ( .A(n3177), .ZN(n2581) );
  AND2_X1 U2967 ( .A1(n2844), .A2(n4963), .ZN(n2847) );
  INV_X1 U2968 ( .A(n2847), .ZN(n2627) );
  INV_X1 U2969 ( .A(n4967), .ZN(n2650) );
  NAND2_X1 U2970 ( .A1(n2715), .A2(IR_REG_31__SCAN_IN), .ZN(n2720) );
  NOR2_X1 U2971 ( .A1(n4921), .A2(n4741), .ZN(n4729) );
  AND2_X1 U2972 ( .A1(n3779), .A2(n3778), .ZN(n4695) );
  NAND2_X1 U2973 ( .A1(n4855), .A2(n4847), .ZN(n2482) );
  INV_X1 U2974 ( .A(n5049), .ZN(n3064) );
  INV_X1 U2975 ( .A(n2713), .ZN(n2733) );
  INV_X1 U2976 ( .A(IR_REG_31__SCAN_IN), .ZN(n2810) );
  MUX2_X1 U2977 ( .A(IR_REG_0__SCAN_IN), .B(DATAI_0_), .S(n3025), .Z(n3079) );
  INV_X1 U2978 ( .A(n3079), .ZN(n2563) );
  AND2_X1 U2979 ( .A1(n2649), .A2(n4967), .ZN(n2483) );
  AND2_X1 U2980 ( .A1(n4669), .A2(n4668), .ZN(n2484) );
  NAND2_X1 U2981 ( .A1(n2631), .A2(n2632), .ZN(n4578) );
  AND2_X1 U2982 ( .A1(n4840), .A2(n4658), .ZN(n2485) );
  AND2_X1 U2983 ( .A1(n3777), .A2(n4885), .ZN(n2486) );
  NAND2_X1 U2984 ( .A1(n4590), .A2(n2842), .ZN(n4591) );
  AND2_X1 U2985 ( .A1(n3648), .A2(n3645), .ZN(n4096) );
  INV_X1 U2986 ( .A(n4096), .ZN(n2502) );
  NOR2_X1 U2987 ( .A1(n4561), .A2(n3774), .ZN(n2487) );
  INV_X1 U2988 ( .A(n3677), .ZN(n4564) );
  AND4_X1 U2989 ( .A1(n3429), .A2(n3428), .A3(n3427), .A4(n3426), .ZN(n3677)
         );
  INV_X1 U2990 ( .A(IR_REG_5__SCAN_IN), .ZN(n2709) );
  NOR2_X1 U2991 ( .A1(n4648), .A2(n5238), .ZN(n2488) );
  OR2_X1 U2992 ( .A1(n4611), .A2(n2613), .ZN(n2612) );
  AND2_X1 U2993 ( .A1(n2837), .A2(n4965), .ZN(n2838) );
  AND2_X1 U2994 ( .A1(n3677), .A2(n3687), .ZN(n2489) );
  AND2_X1 U2995 ( .A1(n4098), .A2(n3643), .ZN(n4080) );
  AND4_X1 U2996 ( .A1(n3470), .A2(n3469), .A3(n3468), .A4(n3467), .ZN(n3702)
         );
  AND2_X1 U2997 ( .A1(n2672), .A2(n2482), .ZN(n2490) );
  NAND2_X1 U2998 ( .A1(n2577), .A2(n2579), .ZN(n3201) );
  INV_X1 U2999 ( .A(IR_REG_0__SCAN_IN), .ZN(n2571) );
  XNOR2_X1 U3000 ( .A(n2915), .B(n4486), .ZN(n2941) );
  INV_X1 U3001 ( .A(n4883), .ZN(n2683) );
  AND2_X1 U3002 ( .A1(n3245), .A2(n3244), .ZN(n3284) );
  NAND2_X1 U3003 ( .A1(n3025), .A2(DATAI_23_), .ZN(n4802) );
  NOR2_X1 U3004 ( .A1(n2886), .A2(n2885), .ZN(n2884) );
  NAND2_X1 U3005 ( .A1(n3025), .A2(DATAI_20_), .ZN(n4868) );
  AND2_X1 U3006 ( .A1(n4881), .A2(n4136), .ZN(n4068) );
  INV_X1 U3007 ( .A(n4068), .ZN(n2518) );
  AND2_X1 U3008 ( .A1(n2644), .A2(n2643), .ZN(n2491) );
  AND2_X1 U3009 ( .A1(n2521), .A2(n4115), .ZN(n2492) );
  NAND2_X1 U3010 ( .A1(n3627), .A2(n3549), .ZN(n2493) );
  NAND2_X1 U3011 ( .A1(n3025), .A2(DATAI_21_), .ZN(n4847) );
  NAND2_X1 U3012 ( .A1(n3122), .A2(n3111), .ZN(n5076) );
  NAND2_X1 U3013 ( .A1(n2575), .A2(n2574), .ZN(n3068) );
  AND2_X1 U3014 ( .A1(n3072), .A2(n3071), .ZN(n4860) );
  AND2_X1 U3015 ( .A1(n2563), .A2(n3080), .ZN(n2494) );
  NAND2_X1 U3016 ( .A1(n3110), .A2(n2506), .ZN(n3122) );
  OR2_X1 U3017 ( .A1(n2814), .A2(n2617), .ZN(n2495) );
  OR2_X1 U3018 ( .A1(n4962), .A2(REG1_REG_15__SCAN_IN), .ZN(n2496) );
  AND2_X1 U3019 ( .A1(n3025), .A2(DATAI_25_), .ZN(n4760) );
  INV_X1 U3020 ( .A(n4960), .ZN(n2619) );
  INV_X1 U3021 ( .A(n4965), .ZN(n2622) );
  AND4_X1 U3022 ( .A1(n4524), .A2(n4523), .A3(n4522), .A4(n4521), .ZN(n2497)
         );
  AND2_X1 U3023 ( .A1(D_REG_16__SCAN_IN), .A2(keyinput_103), .ZN(n2498) );
  OR2_X1 U3024 ( .A1(n4550), .A2(n2553), .ZN(n2499) );
  OAI21_X2 U3025 ( .B1(n3705), .B2(n2518), .A(n2515), .ZN(n4859) );
  NAND2_X1 U3026 ( .A1(n4859), .A2(n4858), .ZN(n4676) );
  AND2_X2 U3027 ( .A1(n2710), .A2(n2522), .ZN(n2713) );
  NAND2_X2 U3028 ( .A1(n4105), .A2(n4108), .ZN(n4063) );
  AOI21_X1 U3029 ( .B1(n2540), .B2(n4483), .A(n4482), .ZN(n4490) );
  INV_X1 U3030 ( .A(n4475), .ZN(n2541) );
  NAND2_X1 U3031 ( .A1(n4732), .A2(n2472), .ZN(n5296) );
  NAND3_X1 U3032 ( .A1(n2559), .A2(n2557), .A3(n2556), .ZN(n5304) );
  NAND2_X1 U3033 ( .A1(n3131), .A2(n3080), .ZN(n2562) );
  NAND3_X1 U3034 ( .A1(n2573), .A2(n2572), .A3(n2571), .ZN(n2742) );
  NAND2_X1 U3035 ( .A1(n2806), .A2(n4505), .ZN(n2805) );
  INV_X1 U3036 ( .A(n2974), .ZN(n2949) );
  INV_X1 U3037 ( .A(n3070), .ZN(n2576) );
  NAND2_X1 U3038 ( .A1(n3155), .A2(n2578), .ZN(n2577) );
  NAND2_X1 U3039 ( .A1(n2720), .A2(n2596), .ZN(n2917) );
  OR2_X1 U3040 ( .A1(n3972), .A2(n2604), .ZN(n2598) );
  NAND2_X1 U3041 ( .A1(n3972), .A2(n2602), .ZN(n2601) );
  INV_X1 U3042 ( .A(n2609), .ZN(n3971) );
  NAND2_X1 U3043 ( .A1(n3850), .A2(n3851), .ZN(n2607) );
  NAND2_X1 U3044 ( .A1(n3836), .A2(n3837), .ZN(n2608) );
  NAND2_X1 U3045 ( .A1(n2713), .A2(n2610), .ZN(n2715) );
  NOR2_X2 U3046 ( .A1(n2714), .A2(IR_REG_10__SCAN_IN), .ZN(n2611) );
  INV_X1 U3047 ( .A(n2838), .ZN(n2631) );
  NAND2_X1 U3048 ( .A1(n2851), .A2(n2639), .ZN(n2638) );
  NAND2_X1 U3049 ( .A1(n2638), .A2(n2640), .ZN(n2634) );
  NOR2_X1 U3050 ( .A1(n2633), .A2(n2638), .ZN(n4640) );
  NAND2_X1 U3051 ( .A1(n2635), .A2(n2634), .ZN(n2857) );
  NAND2_X1 U3052 ( .A1(n2831), .A2(n2645), .ZN(n2641) );
  NOR2_X1 U3053 ( .A1(n5032), .A2(n2822), .ZN(n2999) );
  INV_X1 U3054 ( .A(n2469), .ZN(n2647) );
  INV_X1 U3055 ( .A(n5032), .ZN(n2648) );
  NAND2_X1 U3056 ( .A1(n2653), .A2(n2651), .ZN(n3116) );
  NAND3_X1 U3057 ( .A1(n3110), .A2(n2506), .A3(n3112), .ZN(n2653) );
  INV_X1 U3058 ( .A(n3111), .ZN(n2654) );
  NAND2_X1 U3059 ( .A1(n3636), .A2(n2658), .ZN(n2655) );
  NAND2_X1 U3060 ( .A1(n2655), .A2(n2656), .ZN(n3640) );
  NAND2_X1 U3061 ( .A1(n4740), .A2(n2666), .ZN(n2665) );
  NAND2_X1 U3062 ( .A1(n4740), .A2(n4739), .ZN(n4738) );
  NAND2_X1 U3063 ( .A1(n4833), .A2(n2470), .ZN(n2669) );
  NAND2_X1 U3064 ( .A1(n2669), .A2(n2670), .ZN(n4792) );
  INV_X1 U3065 ( .A(n4833), .ZN(n2673) );
  NAND2_X1 U3066 ( .A1(n3701), .A2(n2676), .ZN(n2675) );
  OAI21_X1 U3067 ( .B1(n3245), .B2(n2692), .A(n2689), .ZN(n3547) );
  NAND2_X1 U3068 ( .A1(n2809), .A2(n2788), .ZN(n2792) );
  OAI211_X1 U3069 ( .C1(n2467), .C2(REG1_REG_1__SCAN_IN), .A(n2751), .B(n2708), 
        .ZN(n2991) );
  NAND2_X1 U3070 ( .A1(n2467), .A2(REG1_REG_1__SCAN_IN), .ZN(n2751) );
  NAND2_X1 U3071 ( .A1(n2805), .A2(IR_REG_31__SCAN_IN), .ZN(n2804) );
  NOR2_X1 U3072 ( .A1(n4725), .A2(n4724), .ZN(n4723) );
  NAND2_X1 U3073 ( .A1(n2966), .A2(REG2_REG_1__SCAN_IN), .ZN(n2931) );
  MUX2_X1 U3074 ( .A(n2467), .B(DATAI_1_), .S(n3025), .Z(n2973) );
  AND3_X1 U3075 ( .A1(n2970), .A2(n2969), .A3(n2968), .ZN(n2971) );
  NAND2_X1 U3076 ( .A1(n3712), .A2(n3711), .ZN(n3710) );
  NOR2_X1 U3077 ( .A1(n3561), .A2(n2707), .ZN(n3562) );
  INV_X1 U3078 ( .A(n3561), .ZN(n3549) );
  AND2_X1 U3079 ( .A1(n2705), .A2(n3593), .ZN(n2702) );
  AND2_X1 U3080 ( .A1(n2797), .A2(n4496), .ZN(n2703) );
  NAND2_X1 U3081 ( .A1(n4825), .A2(n4697), .ZN(n4656) );
  XNOR2_X1 U3082 ( .A(n4568), .B(n3506), .ZN(n3510) );
  INV_X1 U3083 ( .A(n4838), .ZN(n4653) );
  NOR2_X1 U3084 ( .A1(n3380), .A2(n3379), .ZN(n3368) );
  OR2_X1 U3085 ( .A1(n4797), .A2(n4823), .ZN(n2704) );
  XOR2_X1 U3086 ( .A(n3584), .B(n3879), .Z(n2705) );
  AND3_X1 U3087 ( .A1(n3208), .A2(n3207), .A3(n3206), .ZN(n2706) );
  INV_X1 U3088 ( .A(n4868), .ZN(n4696) );
  AND2_X1 U3089 ( .A1(n4567), .A2(n3560), .ZN(n2707) );
  OR2_X1 U3090 ( .A1(n4834), .A2(n4021), .ZN(n4677) );
  NAND2_X1 U3091 ( .A1(n2973), .A2(n3327), .ZN(n2963) );
  OAI21_X1 U3092 ( .B1(n5049), .B2(n2965), .A(n2963), .ZN(n2964) );
  INV_X1 U3093 ( .A(n4593), .ZN(n2842) );
  INV_X1 U3094 ( .A(IR_REG_26__SCAN_IN), .ZN(n4285) );
  NAND2_X1 U3095 ( .A1(n2927), .A2(n2926), .ZN(n2935) );
  AND2_X1 U3096 ( .A1(n3490), .A2(n3489), .ZN(n4126) );
  INV_X1 U3097 ( .A(n4847), .ZN(n4697) );
  INV_X1 U3098 ( .A(IR_REG_13__SCAN_IN), .ZN(n4265) );
  XNOR2_X1 U3099 ( .A(n3146), .B(n3892), .ZN(n3151) );
  NAND2_X1 U3100 ( .A1(n3375), .A2(n3374), .ZN(n3376) );
  AND2_X1 U3101 ( .A1(n3795), .A2(REG3_REG_26__SCAN_IN), .ZN(n3870) );
  INV_X1 U3102 ( .A(n4828), .ZN(n4658) );
  INV_X1 U3103 ( .A(n4079), .ZN(n3114) );
  INV_X1 U3104 ( .A(n4113), .ZN(n3131) );
  INV_X1 U3105 ( .A(n4570), .ZN(n3273) );
  INV_X1 U3106 ( .A(n3376), .ZN(n3377) );
  INV_X1 U3107 ( .A(n4840), .ZN(n4657) );
  NOR2_X1 U3108 ( .A1(n3951), .A2(n3955), .ZN(n3941) );
  NOR2_X1 U3109 ( .A1(n3852), .A2(n3956), .ZN(n3854) );
  AND2_X1 U3110 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n3095) );
  INV_X1 U3111 ( .A(n4825), .ZN(n4855) );
  OR2_X1 U3112 ( .A1(n3821), .A2(n3974), .ZN(n3838) );
  AND2_X1 U3113 ( .A1(n2934), .A2(n5260), .ZN(n3975) );
  AND4_X1 U3114 ( .A1(n3799), .A2(n3798), .A3(n3797), .A4(n3796), .ZN(n4781)
         );
  NOR2_X1 U3115 ( .A1(n2820), .A2(n3007), .ZN(n2821) );
  NOR2_X1 U3116 ( .A1(n3255), .A2(n2835), .ZN(n3483) );
  INV_X1 U3117 ( .A(n4135), .ZN(n4044) );
  NAND2_X1 U3118 ( .A1(n3702), .A2(n3654), .ZN(n3666) );
  INV_X1 U3119 ( .A(n4887), .ZN(n4866) );
  INV_X1 U3120 ( .A(n3560), .ZN(n3567) );
  XNOR2_X1 U3121 ( .A(n2793), .B(IR_REG_26__SCAN_IN), .ZN(n2879) );
  AOI21_X1 U3122 ( .B1(n3869), .B2(n3868), .A(n3867), .ZN(n3909) );
  AND2_X1 U3123 ( .A1(n3898), .A2(n3886), .ZN(n4716) );
  NOR2_X1 U3124 ( .A1(n3585), .A2(n4367), .ZN(n3602) );
  NAND2_X1 U3125 ( .A1(n3425), .A2(REG3_REG_13__SCAN_IN), .ZN(n3466) );
  NAND2_X1 U3126 ( .A1(REG3_REG_18__SCAN_IN), .A2(n3741), .ZN(n3757) );
  INV_X1 U3127 ( .A(n3975), .ZN(n5237) );
  INV_X1 U3128 ( .A(n4781), .ZN(n4664) );
  AND4_X1 U3129 ( .A1(n3746), .A2(n3745), .A3(n3744), .A4(n3743), .ZN(n4886)
         );
  NOR2_X1 U3130 ( .A1(n2986), .A2(n2818), .ZN(n5021) );
  OR2_X1 U3131 ( .A1(n4054), .A2(n4797), .ZN(n4811) );
  INV_X1 U3132 ( .A(n5283), .ZN(n5292) );
  INV_X1 U3133 ( .A(n4860), .ZN(n5256) );
  INV_X1 U3134 ( .A(n5275), .ZN(n5202) );
  INV_X1 U3135 ( .A(n5273), .ZN(n5303) );
  NAND2_X1 U3136 ( .A1(n3068), .A2(n5046), .ZN(n5275) );
  AND2_X1 U3137 ( .A1(n4907), .A2(n4153), .ZN(n4940) );
  AND2_X1 U3138 ( .A1(n2767), .A2(n2766), .ZN(n3193) );
  OR2_X1 U3139 ( .A1(n2953), .A2(n2952), .ZN(n5192) );
  AND2_X1 U3140 ( .A1(n3141), .A2(n3140), .ZN(n5244) );
  NAND4_X1 U3141 ( .A1(n3825), .A2(n3824), .A3(n3823), .A4(n3822), .ZN(n4825)
         );
  NAND4_X1 U3142 ( .A1(n3762), .A2(n3761), .A3(n3760), .A4(n3759), .ZN(n4838)
         );
  OR2_X1 U3143 ( .A1(n2858), .A2(n2920), .ZN(n5042) );
  INV_X1 U3144 ( .A(n5268), .ZN(n4876) );
  INV_X1 U3145 ( .A(n5307), .ZN(n5305) );
  INV_X1 U3146 ( .A(n5311), .ZN(n5308) );
  INV_X1 U3147 ( .A(n4988), .ZN(n4987) );
  INV_X1 U31480 ( .A(n2926), .ZN(n4954) );
  INV_X1 U31490 ( .A(n4089), .ZN(n4957) );
  AND2_X1 U3150 ( .A1(n2732), .A2(n2731), .ZN(n4966) );
  INV_X1 U3151 ( .A(n3088), .ZN(n5075) );
  INV_X1 U3152 ( .A(REG1_REG_18__SCAN_IN), .ZN(n5248) );
  NAND3_X1 U3153 ( .A1(n4269), .A2(n2716), .A3(n2722), .ZN(n2785) );
  NAND2_X1 U3154 ( .A1(n2785), .A2(IR_REG_31__SCAN_IN), .ZN(n2717) );
  OAI21_X1 U3155 ( .B1(n2912), .B2(IR_REG_17__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2718) );
  XNOR2_X1 U3156 ( .A(n2718), .B(IR_REG_18__SCAN_IN), .ZN(n5001) );
  MUX2_X1 U3157 ( .A(n5248), .B(REG1_REG_18__SCAN_IN), .S(n5001), .Z(n2816) );
  INV_X1 U3158 ( .A(IR_REG_17__SCAN_IN), .ZN(n2719) );
  XNOR2_X1 U3159 ( .A(n2912), .B(n2719), .ZN(n4960) );
  NAND2_X1 U3160 ( .A1(n2720), .A2(n4269), .ZN(n2721) );
  NAND2_X1 U3161 ( .A1(n2721), .A2(IR_REG_31__SCAN_IN), .ZN(n2723) );
  NAND2_X1 U3162 ( .A1(n2723), .A2(n2722), .ZN(n2778) );
  OR2_X1 U3163 ( .A1(n2723), .A2(n2722), .ZN(n2724) );
  OR2_X1 U3164 ( .A1(n2725), .A2(n2810), .ZN(n2726) );
  XNOR2_X1 U3165 ( .A(n2726), .B(IR_REG_13__SCAN_IN), .ZN(n4964) );
  NOR2_X1 U3166 ( .A1(n4964), .A2(REG1_REG_13__SCAN_IN), .ZN(n2775) );
  AND2_X1 U3167 ( .A1(n2727), .A2(IR_REG_31__SCAN_IN), .ZN(n2730) );
  INV_X1 U3168 ( .A(n2730), .ZN(n2728) );
  NAND2_X1 U3169 ( .A1(n2728), .A2(n4470), .ZN(n2731) );
  NAND2_X1 U3170 ( .A1(n2731), .A2(IR_REG_31__SCAN_IN), .ZN(n2729) );
  XNOR2_X1 U3171 ( .A(n2729), .B(IR_REG_12__SCAN_IN), .ZN(n4965) );
  INV_X1 U3172 ( .A(REG1_REG_11__SCAN_IN), .ZN(n5163) );
  NAND2_X1 U3173 ( .A1(n2730), .A2(IR_REG_11__SCAN_IN), .ZN(n2732) );
  INV_X1 U3174 ( .A(n4966), .ZN(n3488) );
  NAND2_X1 U3175 ( .A1(n2733), .A2(IR_REG_31__SCAN_IN), .ZN(n2734) );
  XNOR2_X1 U3176 ( .A(n2734), .B(IR_REG_10__SCAN_IN), .ZN(n3360) );
  NOR2_X1 U3177 ( .A1(n2735), .A2(n2810), .ZN(n2736) );
  MUX2_X1 U3178 ( .A(n2810), .B(n2736), .S(IR_REG_9__SCAN_IN), .Z(n2737) );
  INV_X1 U3179 ( .A(n2737), .ZN(n2738) );
  AND2_X1 U3180 ( .A1(n2733), .A2(n2738), .ZN(n3326) );
  NAND2_X1 U3181 ( .A1(n3326), .A2(REG1_REG_9__SCAN_IN), .ZN(n2772) );
  INV_X1 U3182 ( .A(REG1_REG_9__SCAN_IN), .ZN(n2739) );
  MUX2_X1 U3183 ( .A(REG1_REG_9__SCAN_IN), .B(n2739), .S(n3326), .Z(n3058) );
  OAI21_X1 U3184 ( .B1(n2740), .B2(IR_REG_6__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2765) );
  NAND2_X1 U3185 ( .A1(n2765), .A2(n4254), .ZN(n2767) );
  NAND2_X1 U3186 ( .A1(n2767), .A2(IR_REG_31__SCAN_IN), .ZN(n2741) );
  XNOR2_X1 U3187 ( .A(n2741), .B(IR_REG_8__SCAN_IN), .ZN(n3302) );
  INV_X1 U3188 ( .A(REG1_REG_5__SCAN_IN), .ZN(n5117) );
  NAND2_X1 U3189 ( .A1(n2742), .A2(IR_REG_31__SCAN_IN), .ZN(n2743) );
  MUX2_X1 U3190 ( .A(IR_REG_31__SCAN_IN), .B(n2743), .S(IR_REG_5__SCAN_IN), 
        .Z(n2744) );
  AND2_X1 U3191 ( .A1(n2744), .A2(n2740), .ZN(n4968) );
  INV_X1 U3192 ( .A(n4968), .ZN(n3006) );
  NAND2_X1 U3193 ( .A1(n2752), .A2(n4245), .ZN(n2745) );
  NAND2_X1 U3194 ( .A1(n2745), .A2(IR_REG_31__SCAN_IN), .ZN(n2747) );
  NAND2_X1 U3195 ( .A1(n2747), .A2(n4456), .ZN(n2749) );
  NAND2_X1 U3196 ( .A1(n2749), .A2(IR_REG_31__SCAN_IN), .ZN(n2746) );
  XNOR2_X1 U3197 ( .A(n2746), .B(IR_REG_4__SCAN_IN), .ZN(n3094) );
  OR2_X1 U3198 ( .A1(n2747), .A2(n4456), .ZN(n2748) );
  INV_X1 U3199 ( .A(REG1_REG_1__SCAN_IN), .ZN(n2990) );
  NAND2_X1 U3200 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2750)
         );
  INV_X1 U3201 ( .A(n2467), .ZN(n2995) );
  OAI21_X1 U3202 ( .B1(n2990), .B2(n2995), .A(n2991), .ZN(n5025) );
  INV_X1 U3203 ( .A(REG1_REG_2__SCAN_IN), .ZN(n2755) );
  MUX2_X1 U3204 ( .A(REG1_REG_2__SCAN_IN), .B(n2755), .S(n5022), .Z(n5024) );
  NAND2_X1 U3205 ( .A1(n5022), .A2(REG1_REG_2__SCAN_IN), .ZN(n2756) );
  NAND2_X1 U3206 ( .A1(n3088), .A2(n2757), .ZN(n2758) );
  NAND2_X1 U3207 ( .A1(n2758), .A2(n3010), .ZN(n2759) );
  NAND2_X1 U3208 ( .A1(n3094), .A2(n2759), .ZN(n2760) );
  INV_X1 U3209 ( .A(n3094), .ZN(n5105) );
  XNOR2_X1 U32100 ( .A(n2759), .B(n5105), .ZN(n5039) );
  NAND2_X1 U32110 ( .A1(REG1_REG_4__SCAN_IN), .A2(n5039), .ZN(n5037) );
  NAND2_X1 U32120 ( .A1(n2760), .A2(n5037), .ZN(n3003) );
  MUX2_X1 U32130 ( .A(REG1_REG_5__SCAN_IN), .B(n5117), .S(n4968), .Z(n3002) );
  NAND2_X1 U32140 ( .A1(n3003), .A2(n3002), .ZN(n3001) );
  NAND2_X1 U32150 ( .A1(n2740), .A2(IR_REG_31__SCAN_IN), .ZN(n2761) );
  XNOR2_X1 U32160 ( .A(n2761), .B(IR_REG_6__SCAN_IN), .ZN(n4967) );
  XNOR2_X1 U32170 ( .A(n2762), .B(n4967), .ZN(n2978) );
  INV_X1 U32180 ( .A(REG1_REG_6__SCAN_IN), .ZN(n2764) );
  INV_X1 U32190 ( .A(n2762), .ZN(n2763) );
  OAI22_X1 U32200 ( .A1(n2978), .A2(n2764), .B1(n2763), .B2(n2650), .ZN(n2889)
         );
  INV_X1 U32210 ( .A(REG1_REG_7__SCAN_IN), .ZN(n2768) );
  OR2_X1 U32220 ( .A1(n2765), .A2(n4254), .ZN(n2766) );
  MUX2_X1 U32230 ( .A(REG1_REG_7__SCAN_IN), .B(n2768), .S(n3193), .Z(n2888) );
  NAND2_X1 U32240 ( .A1(n2889), .A2(n2888), .ZN(n2887) );
  NAND2_X1 U32250 ( .A1(n3193), .A2(REG1_REG_7__SCAN_IN), .ZN(n2769) );
  NAND2_X1 U32260 ( .A1(n3302), .A2(n2770), .ZN(n2771) );
  INV_X1 U32270 ( .A(n3302), .ZN(n5134) );
  XNOR2_X1 U32280 ( .A(n2770), .B(n5134), .ZN(n3020) );
  NAND2_X1 U32290 ( .A1(REG1_REG_8__SCAN_IN), .A2(n3020), .ZN(n3019) );
  NAND2_X1 U32300 ( .A1(n2771), .A2(n3019), .ZN(n3059) );
  NAND2_X1 U32310 ( .A1(n3058), .A2(n3059), .ZN(n3057) );
  NAND2_X1 U32320 ( .A1(n2772), .A2(n3057), .ZN(n2773) );
  NAND2_X1 U32330 ( .A1(n3360), .A2(n2773), .ZN(n2774) );
  INV_X1 U32340 ( .A(n3360), .ZN(n5151) );
  XNOR2_X1 U32350 ( .A(n2773), .B(n5151), .ZN(n3259) );
  NAND2_X1 U32360 ( .A1(REG1_REG_10__SCAN_IN), .A2(n3259), .ZN(n3258) );
  NAND2_X1 U32370 ( .A1(n2774), .A2(n3258), .ZN(n3479) );
  MUX2_X1 U32380 ( .A(REG1_REG_11__SCAN_IN), .B(n5163), .S(n4966), .Z(n3478)
         );
  NAND2_X1 U32390 ( .A1(n3479), .A2(n3478), .ZN(n3477) );
  AOI21_X1 U32400 ( .B1(n4964), .B2(REG1_REG_13__SCAN_IN), .A(n4585), .ZN(
        n2776) );
  XNOR2_X1 U32410 ( .A(n2720), .B(IR_REG_14__SCAN_IN), .ZN(n4963) );
  XNOR2_X1 U32420 ( .A(n2776), .B(n4963), .ZN(n4600) );
  INV_X1 U32430 ( .A(n2776), .ZN(n2777) );
  NAND2_X1 U32440 ( .A1(n2778), .A2(IR_REG_31__SCAN_IN), .ZN(n2779) );
  XNOR2_X1 U32450 ( .A(n2779), .B(IR_REG_16__SCAN_IN), .ZN(n4961) );
  INV_X1 U32460 ( .A(n4961), .ZN(n4623) );
  NOR2_X1 U32470 ( .A1(n4622), .A2(REG1_REG_16__SCAN_IN), .ZN(n4637) );
  INV_X1 U32480 ( .A(n2781), .ZN(n4636) );
  INV_X1 U32490 ( .A(REG1_REG_17__SCAN_IN), .ZN(n2782) );
  OR2_X1 U32500 ( .A1(n4960), .A2(n2782), .ZN(n2784) );
  NAND2_X1 U32510 ( .A1(n4960), .A2(n2782), .ZN(n2783) );
  NAND2_X1 U32520 ( .A1(n2784), .A2(n2783), .ZN(n4635) );
  OAI21_X1 U32530 ( .B1(n4637), .B2(n4636), .A(n4635), .ZN(n4634) );
  NOR2_X2 U32540 ( .A1(IR_REG_18__SCAN_IN), .A2(IR_REG_17__SCAN_IN), .ZN(n2913) );
  NAND4_X1 U32550 ( .A1(n2913), .A2(n4486), .A3(n4485), .A4(n4265), .ZN(n2786)
         );
  NAND2_X1 U32560 ( .A1(n2798), .A2(n2797), .ZN(n2800) );
  NAND2_X1 U32570 ( .A1(n2800), .A2(IR_REG_31__SCAN_IN), .ZN(n2789) );
  OR2_X1 U32580 ( .A1(n2803), .A2(n2810), .ZN(n2793) );
  NAND2_X1 U32590 ( .A1(n2478), .A2(IR_REG_31__SCAN_IN), .ZN(n2794) );
  MUX2_X1 U32600 ( .A(IR_REG_31__SCAN_IN), .B(n2794), .S(IR_REG_25__SCAN_IN), 
        .Z(n2796) );
  INV_X1 U32610 ( .A(n2803), .ZN(n2795) );
  NAND2_X1 U32620 ( .A1(n2796), .A2(n2795), .ZN(n2895) );
  INV_X1 U32630 ( .A(n2895), .ZN(n4955) );
  OR2_X1 U32640 ( .A1(n2798), .A2(n2797), .ZN(n2799) );
  NAND2_X1 U32650 ( .A1(n2800), .A2(n2799), .ZN(n3136) );
  NAND2_X1 U32660 ( .A1(n3136), .A2(STATE_REG_SCAN_IN), .ZN(n4970) );
  INV_X1 U32670 ( .A(n4970), .ZN(n2882) );
  INV_X1 U32680 ( .A(n2951), .ZN(n2802) );
  INV_X1 U32690 ( .A(n3136), .ZN(n2801) );
  NAND2_X1 U32700 ( .A1(n2801), .A2(STATE_REG_SCAN_IN), .ZN(n4156) );
  NAND2_X1 U32710 ( .A1(n2802), .A2(n4156), .ZN(n2859) );
  INV_X1 U32720 ( .A(IR_REG_27__SCAN_IN), .ZN(n4505) );
  INV_X1 U32730 ( .A(IR_REG_28__SCAN_IN), .ZN(n4506) );
  NAND2_X1 U32740 ( .A1(n2792), .A2(IR_REG_31__SCAN_IN), .ZN(n2808) );
  XNOR2_X1 U32750 ( .A(n2808), .B(n2790), .ZN(n3070) );
  NOR2_X1 U32760 ( .A1(n2809), .A2(n2810), .ZN(n2811) );
  MUX2_X1 U32770 ( .A(n2810), .B(n2811), .S(IR_REG_21__SCAN_IN), .Z(n2813) );
  INV_X1 U32780 ( .A(n2792), .ZN(n2812) );
  NAND2_X1 U32790 ( .A1(n2949), .A2(n3136), .ZN(n2861) );
  NAND3_X1 U32800 ( .A1(n2859), .A2(n3025), .A3(n2861), .ZN(n2858) );
  INV_X1 U32810 ( .A(n4989), .ZN(n5013) );
  OR2_X1 U32820 ( .A1(n2858), .A2(n5013), .ZN(n4632) );
  NOR2_X1 U32830 ( .A1(n5001), .A2(REG1_REG_18__SCAN_IN), .ZN(n2814) );
  AOI211_X1 U32840 ( .C1(n2816), .C2(n2815), .A(n4632), .B(n5000), .ZN(n2867)
         );
  INV_X1 U32850 ( .A(REG2_REG_10__SCAN_IN), .ZN(n3257) );
  INV_X1 U32860 ( .A(REG2_REG_8__SCAN_IN), .ZN(n3440) );
  NAND2_X1 U32870 ( .A1(n4969), .A2(REG2_REG_1__SCAN_IN), .ZN(n2817) );
  OAI21_X1 U32880 ( .B1(n2467), .B2(REG2_REG_1__SCAN_IN), .A(n2817), .ZN(n2987) );
  NAND2_X1 U32890 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(
        n5012) );
  NOR2_X1 U32900 ( .A1(n2987), .A2(n5012), .ZN(n2986) );
  INV_X1 U32910 ( .A(n2817), .ZN(n2818) );
  XNOR2_X1 U32920 ( .A(n5022), .B(REG2_REG_2__SCAN_IN), .ZN(n5020) );
  NOR2_X1 U32930 ( .A1(n5021), .A2(n5020), .ZN(n5019) );
  NOR2_X1 U32940 ( .A1(n2819), .A2(n5075), .ZN(n2820) );
  INV_X1 U32950 ( .A(REG2_REG_3__SCAN_IN), .ZN(n3009) );
  XNOR2_X1 U32960 ( .A(n2819), .B(n5075), .ZN(n3008) );
  NOR2_X1 U32970 ( .A1(n3009), .A2(n3008), .ZN(n3007) );
  NOR2_X1 U32980 ( .A1(n2821), .A2(n5105), .ZN(n2822) );
  INV_X1 U32990 ( .A(REG2_REG_4__SCAN_IN), .ZN(n5034) );
  XOR2_X1 U33000 ( .A(n2821), .B(n3094), .Z(n5033) );
  NOR2_X1 U33010 ( .A1(n5034), .A2(n5033), .ZN(n5032) );
  INV_X1 U33020 ( .A(REG2_REG_5__SCAN_IN), .ZN(n2823) );
  MUX2_X1 U33030 ( .A(n2823), .B(REG2_REG_5__SCAN_IN), .S(n4968), .Z(n2998) );
  NAND2_X1 U33040 ( .A1(n4968), .A2(REG2_REG_5__SCAN_IN), .ZN(n2824) );
  INV_X1 U33050 ( .A(n2827), .ZN(n2826) );
  INV_X1 U33060 ( .A(REG2_REG_6__SCAN_IN), .ZN(n3250) );
  NOR2_X1 U33070 ( .A1(n2981), .A2(n3250), .ZN(n2980) );
  NOR2_X1 U33080 ( .A1(n2827), .A2(n2980), .ZN(n2886) );
  NAND2_X1 U33090 ( .A1(n3193), .A2(REG2_REG_7__SCAN_IN), .ZN(n2828) );
  OAI21_X1 U33100 ( .B1(n3193), .B2(REG2_REG_7__SCAN_IN), .A(n2828), .ZN(n2885) );
  NOR2_X1 U33110 ( .A1(n2830), .A2(n5134), .ZN(n2831) );
  NAND2_X1 U33120 ( .A1(n3326), .A2(REG2_REG_9__SCAN_IN), .ZN(n2832) );
  OAI21_X1 U33130 ( .B1(n3326), .B2(REG2_REG_9__SCAN_IN), .A(n2832), .ZN(n3056) );
  XNOR2_X1 U33140 ( .A(n2834), .B(n5151), .ZN(n3256) );
  NOR2_X1 U33150 ( .A1(n3257), .A2(n3256), .ZN(n3255) );
  NOR2_X1 U33160 ( .A1(n2834), .A2(n5151), .ZN(n2835) );
  INV_X1 U33170 ( .A(REG2_REG_11__SCAN_IN), .ZN(n3572) );
  MUX2_X1 U33180 ( .A(n3572), .B(REG2_REG_11__SCAN_IN), .S(n4966), .Z(n3482)
         );
  NAND2_X1 U33190 ( .A1(n4966), .A2(REG2_REG_11__SCAN_IN), .ZN(n2836) );
  NAND2_X1 U33200 ( .A1(n3480), .A2(n2836), .ZN(n2837) );
  INV_X1 U33210 ( .A(REG2_REG_12__SCAN_IN), .ZN(n4580) );
  INV_X1 U33220 ( .A(REG2_REG_13__SCAN_IN), .ZN(n2839) );
  OR2_X1 U33230 ( .A1(n4964), .A2(n2839), .ZN(n2841) );
  NAND2_X1 U33240 ( .A1(n4964), .A2(n2839), .ZN(n2840) );
  AND2_X1 U33250 ( .A1(n2841), .A2(n2840), .ZN(n4593) );
  NAND2_X1 U33260 ( .A1(n4964), .A2(REG2_REG_13__SCAN_IN), .ZN(n2843) );
  NAND2_X1 U33270 ( .A1(n4591), .A2(n2843), .ZN(n2844) );
  INV_X1 U33280 ( .A(n2844), .ZN(n2846) );
  INV_X1 U33290 ( .A(n4963), .ZN(n2845) );
  INV_X1 U33300 ( .A(REG2_REG_14__SCAN_IN), .ZN(n4605) );
  NAND2_X1 U33310 ( .A1(n4962), .A2(REG2_REG_15__SCAN_IN), .ZN(n2849) );
  OR2_X1 U33320 ( .A1(n4962), .A2(REG2_REG_15__SCAN_IN), .ZN(n2848) );
  NAND2_X1 U33330 ( .A1(n2849), .A2(n2848), .ZN(n4615) );
  INV_X1 U33340 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4627) );
  OR2_X1 U33350 ( .A1(n2850), .A2(n4961), .ZN(n2851) );
  INV_X1 U33360 ( .A(REG2_REG_17__SCAN_IN), .ZN(n2853) );
  NOR2_X1 U33370 ( .A1(n4960), .A2(n2853), .ZN(n2852) );
  AOI21_X1 U33380 ( .B1(n2853), .B2(n4960), .A(n2852), .ZN(n4642) );
  INV_X1 U33390 ( .A(REG2_REG_18__SCAN_IN), .ZN(n2854) );
  INV_X1 U33400 ( .A(n5001), .ZN(n5229) );
  AOI22_X1 U33410 ( .A1(n5001), .A2(n2854), .B1(REG2_REG_18__SCAN_IN), .B2(
        n5229), .ZN(n2856) );
  NOR2_X1 U33420 ( .A1(n2857), .A2(n2856), .ZN(n4997) );
  INV_X1 U33430 ( .A(n2858), .ZN(n4993) );
  INV_X1 U33440 ( .A(n2855), .ZN(n2920) );
  NAND3_X1 U33450 ( .A1(n4993), .A2(n5013), .A3(n2920), .ZN(n5031) );
  AOI211_X1 U33460 ( .C1(n2857), .C2(n2856), .A(n4997), .B(n5031), .ZN(n2866)
         );
  INV_X1 U33470 ( .A(n2859), .ZN(n2860) );
  AOI21_X1 U33480 ( .B1(n4000), .B2(n2861), .A(n2860), .ZN(n5003) );
  INV_X1 U33490 ( .A(REG3_REG_18__SCAN_IN), .ZN(n2862) );
  NOR2_X1 U33500 ( .A1(STATE_REG_SCAN_IN), .A2(n2862), .ZN(n2863) );
  AOI21_X1 U33510 ( .B1(n5036), .B2(ADDR_REG_18__SCAN_IN), .A(n2863), .ZN(
        n2864) );
  OAI21_X1 U33520 ( .B1(n5229), .B2(n5042), .A(n2864), .ZN(n2865) );
  OR3_X1 U3353 ( .A1(n2867), .A2(n2866), .A3(n2865), .ZN(U3258) );
  NOR2_X2 U33540 ( .A1(n2943), .A2(n4970), .ZN(U4043) );
  INV_X2 U3355 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  INV_X1 U3356 ( .A(DATAI_22_), .ZN(n2868) );
  MUX2_X1 U3357 ( .A(n2868), .B(n3070), .S(STATE_REG_SCAN_IN), .Z(n2869) );
  INV_X1 U3358 ( .A(n2869), .ZN(U3330) );
  INV_X1 U3359 ( .A(n2879), .ZN(n2896) );
  INV_X1 U3360 ( .A(DATAI_26_), .ZN(n2870) );
  MUX2_X1 U3361 ( .A(n2896), .B(n2870), .S(U3149), .Z(n2871) );
  INV_X1 U3362 ( .A(n2871), .ZN(U3326) );
  INV_X1 U3363 ( .A(DATAI_30_), .ZN(n2876) );
  NOR2_X1 U3364 ( .A1(IR_REG_27__SCAN_IN), .A2(IR_REG_28__SCAN_IN), .ZN(n2872)
         );
  NAND2_X1 U3365 ( .A1(n2873), .A2(n2872), .ZN(n2922) );
  INV_X1 U3366 ( .A(n2922), .ZN(n2874) );
  INV_X1 U3367 ( .A(IR_REG_29__SCAN_IN), .ZN(n4292) );
  NAND2_X1 U3368 ( .A1(n2874), .A2(n4292), .ZN(n2921) );
  INV_X1 U3369 ( .A(IR_REG_30__SCAN_IN), .ZN(n4510) );
  XNOR2_X2 U3370 ( .A(n2875), .B(n4510), .ZN(n2927) );
  MUX2_X1 U3371 ( .A(n2876), .B(n2927), .S(STATE_REG_SCAN_IN), .Z(n2877) );
  INV_X1 U3372 ( .A(n2877), .ZN(U3322) );
  NAND2_X1 U3373 ( .A1(n2895), .A2(B_REG_SCAN_IN), .ZN(n2878) );
  MUX2_X1 U3374 ( .A(n2878), .B(B_REG_SCAN_IN), .S(n4956), .Z(n2880) );
  NAND2_X1 U3375 ( .A1(n2910), .A2(n2951), .ZN(n4988) );
  INV_X1 U3376 ( .A(D_REG_0__SCAN_IN), .ZN(n4514) );
  INV_X1 U3377 ( .A(n4956), .ZN(n2881) );
  NAND2_X1 U3378 ( .A1(n2896), .A2(n2881), .ZN(n2909) );
  INV_X1 U3379 ( .A(n2909), .ZN(n2883) );
  AOI22_X1 U3380 ( .A1(n4988), .A2(n4514), .B1(n2883), .B2(n2882), .ZN(U3458)
         );
  AOI211_X1 U3381 ( .C1(n2886), .C2(n2885), .A(n2884), .B(n5031), .ZN(n2894)
         );
  INV_X1 U3382 ( .A(n3193), .ZN(n5127) );
  OAI211_X1 U3383 ( .C1(n2889), .C2(n2888), .A(n5038), .B(n2887), .ZN(n2892)
         );
  INV_X1 U3384 ( .A(REG3_REG_7__SCAN_IN), .ZN(n4434) );
  NOR2_X1 U3385 ( .A1(STATE_REG_SCAN_IN), .A2(n4434), .ZN(n2890) );
  AOI21_X1 U3386 ( .B1(n5003), .B2(ADDR_REG_7__SCAN_IN), .A(n2890), .ZN(n2891)
         );
  OAI211_X1 U3387 ( .C1(n5042), .C2(n5127), .A(n2892), .B(n2891), .ZN(n2893)
         );
  OR2_X1 U3388 ( .A1(n2894), .A2(n2893), .ZN(U3247) );
  NOR2_X1 U3389 ( .A1(n5036), .A2(U4043), .ZN(U3148) );
  NAND2_X1 U3390 ( .A1(n2896), .A2(n2895), .ZN(n4952) );
  OAI21_X1 U3391 ( .B1(n2910), .B2(D_REG_1__SCAN_IN), .A(n4952), .ZN(n4905) );
  INV_X1 U3392 ( .A(n4905), .ZN(n2908) );
  NOR2_X1 U3393 ( .A1(D_REG_2__SCAN_IN), .A2(D_REG_3__SCAN_IN), .ZN(n2900) );
  NOR4_X1 U3394 ( .A1(D_REG_12__SCAN_IN), .A2(D_REG_5__SCAN_IN), .A3(
        D_REG_7__SCAN_IN), .A4(D_REG_10__SCAN_IN), .ZN(n2899) );
  NOR4_X1 U3395 ( .A1(D_REG_8__SCAN_IN), .A2(D_REG_14__SCAN_IN), .A3(
        D_REG_6__SCAN_IN), .A4(D_REG_17__SCAN_IN), .ZN(n2898) );
  NOR4_X1 U3396 ( .A1(D_REG_9__SCAN_IN), .A2(D_REG_22__SCAN_IN), .A3(
        D_REG_20__SCAN_IN), .A4(D_REG_11__SCAN_IN), .ZN(n2897) );
  NAND4_X1 U3397 ( .A1(n2900), .A2(n2899), .A3(n2898), .A4(n2897), .ZN(n2907)
         );
  NOR4_X1 U3398 ( .A1(D_REG_30__SCAN_IN), .A2(D_REG_31__SCAN_IN), .A3(
        D_REG_28__SCAN_IN), .A4(D_REG_25__SCAN_IN), .ZN(n2904) );
  NOR4_X1 U3399 ( .A1(D_REG_29__SCAN_IN), .A2(D_REG_26__SCAN_IN), .A3(
        D_REG_24__SCAN_IN), .A4(D_REG_27__SCAN_IN), .ZN(n2903) );
  NOR4_X1 U3400 ( .A1(D_REG_16__SCAN_IN), .A2(D_REG_15__SCAN_IN), .A3(
        D_REG_13__SCAN_IN), .A4(D_REG_4__SCAN_IN), .ZN(n2902) );
  NOR4_X1 U3401 ( .A1(D_REG_23__SCAN_IN), .A2(D_REG_21__SCAN_IN), .A3(
        D_REG_19__SCAN_IN), .A4(D_REG_18__SCAN_IN), .ZN(n2901) );
  NAND4_X1 U3402 ( .A1(n2904), .A2(n2903), .A3(n2902), .A4(n2901), .ZN(n2906)
         );
  INV_X1 U3403 ( .A(n2910), .ZN(n2905) );
  OAI21_X1 U3404 ( .B1(n2907), .B2(n2906), .A(n2905), .ZN(n4904) );
  AND2_X1 U3405 ( .A1(n2908), .A2(n4904), .ZN(n3065) );
  OAI21_X1 U3406 ( .B1(n2910), .B2(D_REG_0__SCAN_IN), .A(n2909), .ZN(n4907) );
  INV_X1 U3407 ( .A(n4907), .ZN(n2911) );
  NAND2_X1 U3408 ( .A1(n3065), .A2(n2911), .ZN(n2953) );
  INV_X1 U3409 ( .A(n2941), .ZN(n4958) );
  NAND2_X1 U3410 ( .A1(n3070), .A2(n4089), .ZN(n5047) );
  INV_X1 U3411 ( .A(n5047), .ZN(n3077) );
  NOR2_X1 U3412 ( .A1(n5283), .A2(U3149), .ZN(n2916) );
  NAND2_X1 U3413 ( .A1(n2953), .A2(n2916), .ZN(n3140) );
  NAND2_X1 U3414 ( .A1(n2917), .A2(IR_REG_19__SCAN_IN), .ZN(n2918) );
  NAND2_X1 U3415 ( .A1(n2941), .A2(n5006), .ZN(n2945) );
  NAND2_X1 U3416 ( .A1(n2945), .A2(n3077), .ZN(n2950) );
  NAND2_X1 U3417 ( .A1(n2953), .A2(n2950), .ZN(n3138) );
  NAND2_X1 U3418 ( .A1(n2945), .A2(n2949), .ZN(n3137) );
  NAND2_X1 U3419 ( .A1(n2951), .A2(n3137), .ZN(n4906) );
  INV_X1 U3420 ( .A(n4906), .ZN(n4153) );
  NAND3_X1 U3421 ( .A1(n3140), .A2(n3138), .A3(n4153), .ZN(n3050) );
  INV_X1 U3422 ( .A(n3050), .ZN(n2956) );
  INV_X1 U3423 ( .A(REG3_REG_0__SCAN_IN), .ZN(n4996) );
  OR2_X1 U3424 ( .A1(n2953), .A2(n4906), .ZN(n3403) );
  NAND2_X1 U3425 ( .A1(n2855), .A2(n2949), .ZN(n5048) );
  NAND2_X1 U3426 ( .A1(n5231), .A2(n4839), .ZN(n3976) );
  INV_X1 U3427 ( .A(n3976), .ZN(n3049) );
  INV_X1 U3428 ( .A(n2927), .ZN(n2925) );
  NAND2_X1 U3429 ( .A1(n2922), .A2(IR_REG_31__SCAN_IN), .ZN(n2923) );
  AND2_X2 U3430 ( .A1(n4954), .A2(n2927), .ZN(n3043) );
  NAND2_X1 U3431 ( .A1(n3043), .A2(REG1_REG_1__SCAN_IN), .ZN(n2929) );
  NAND2_X1 U3432 ( .A1(n2466), .A2(REG0_REG_1__SCAN_IN), .ZN(n2928) );
  NAND2_X1 U3433 ( .A1(n2951), .A2(n5292), .ZN(n2932) );
  OR2_X1 U3434 ( .A1(n2953), .A2(n2932), .ZN(n2934) );
  NAND2_X1 U3435 ( .A1(n2941), .A2(n4959), .ZN(n5056) );
  OR2_X1 U3436 ( .A1(n5056), .A2(n5047), .ZN(n4903) );
  INV_X1 U3437 ( .A(n4903), .ZN(n2933) );
  AOI22_X1 U3438 ( .A1(n3049), .A2(n3064), .B1(n3079), .B2(n5237), .ZN(n2955)
         );
  INV_X1 U3439 ( .A(REG1_REG_0__SCAN_IN), .ZN(n5052) );
  NAND2_X1 U3440 ( .A1(n3044), .A2(REG0_REG_0__SCAN_IN), .ZN(n2938) );
  NAND2_X1 U3441 ( .A1(n2966), .A2(REG2_REG_0__SCAN_IN), .ZN(n2937) );
  NAND2_X1 U3442 ( .A1(n3043), .A2(REG1_REG_0__SCAN_IN), .ZN(n2936) );
  NAND2_X1 U3443 ( .A1(n2967), .A2(REG3_REG_0__SCAN_IN), .ZN(n2939) );
  INV_X1 U3444 ( .A(n2959), .ZN(n2942) );
  NAND2_X1 U3446 ( .A1(n3079), .A2(n3327), .ZN(n2960) );
  OAI211_X1 U3447 ( .C1(n2943), .C2(n5052), .A(n2944), .B(n2960), .ZN(n2958)
         );
  NAND2_X1 U3448 ( .A1(n4574), .A2(n3882), .ZN(n2948) );
  NOR2_X1 U3449 ( .A1(n2943), .A2(n2571), .ZN(n2946) );
  NAND2_X1 U3450 ( .A1(n2948), .A2(n2947), .ZN(n2957) );
  XOR2_X1 U3451 ( .A(n2958), .B(n2957), .Z(n5011) );
  NAND3_X1 U3452 ( .A1(n2951), .A2(n2974), .A3(n2950), .ZN(n2952) );
  NAND2_X1 U3453 ( .A1(n5011), .A2(n5239), .ZN(n2954) );
  OAI211_X1 U3454 ( .C1(n2956), .C2(n4996), .A(n2955), .B(n2954), .ZN(U3229)
         );
  NAND2_X1 U3455 ( .A1(n2958), .A2(n2957), .ZN(n2962) );
  AND2_X4 U3456 ( .A1(n3068), .A2(n2959), .ZN(n3879) );
  NAND2_X1 U3457 ( .A1(n2960), .A2(n3879), .ZN(n2961) );
  NAND2_X1 U34580 ( .A1(n2962), .A2(n2961), .ZN(n3031) );
  XNOR2_X1 U34590 ( .A(n2964), .B(n3879), .ZN(n3033) );
  OAI22_X1 U3460 ( .A1(n5049), .A2(n3891), .B1(n3080), .B2(n2965), .ZN(n3034)
         );
  XNOR2_X1 U3461 ( .A(n3033), .B(n3034), .ZN(n3032) );
  XNOR2_X1 U3462 ( .A(n3031), .B(n3032), .ZN(n2977) );
  NAND2_X1 U3463 ( .A1(n3044), .A2(REG0_REG_2__SCAN_IN), .ZN(n2970) );
  NAND2_X1 U3464 ( .A1(n3043), .A2(REG1_REG_2__SCAN_IN), .ZN(n2969) );
  NAND2_X1 U3465 ( .A1(n2967), .A2(REG3_REG_2__SCAN_IN), .ZN(n2968) );
  AOI22_X1 U3466 ( .A1(n3049), .A2(n3087), .B1(n2973), .B2(n5237), .ZN(n2976)
         );
  OR2_X1 U34670 ( .A1(n2855), .A2(n2974), .ZN(n4887) );
  NAND2_X1 U3468 ( .A1(n5231), .A2(n4866), .ZN(n3977) );
  INV_X1 U34690 ( .A(n3977), .ZN(n3051) );
  AOI22_X1 U3470 ( .A1(n3051), .A2(n4574), .B1(REG3_REG_1__SCAN_IN), .B2(n3050), .ZN(n2975) );
  OAI211_X1 U34710 ( .C1(n2977), .C2(n5192), .A(n2976), .B(n2975), .ZN(U3219)
         );
  XNOR2_X1 U3472 ( .A(n2978), .B(REG1_REG_6__SCAN_IN), .ZN(n2984) );
  AND2_X1 U34730 ( .A1(REG3_REG_6__SCAN_IN), .A2(U3149), .ZN(n3221) );
  AOI21_X1 U3474 ( .B1(n5003), .B2(ADDR_REG_6__SCAN_IN), .A(n3221), .ZN(n2979)
         );
  OAI21_X1 U34750 ( .B1(n2650), .B2(n5042), .A(n2979), .ZN(n2983) );
  AOI211_X1 U3476 ( .C1(n3250), .C2(n2981), .A(n2980), .B(n5031), .ZN(n2982)
         );
  AOI211_X1 U34770 ( .C1(n5038), .C2(n2984), .A(n2983), .B(n2982), .ZN(n2985)
         );
  INV_X1 U3478 ( .A(n2985), .ZN(U3246) );
  AOI211_X1 U34790 ( .C1(n5012), .C2(n2987), .A(n2986), .B(n5031), .ZN(n2989)
         );
  INV_X1 U3480 ( .A(REG3_REG_1__SCAN_IN), .ZN(n4220) );
  NOR2_X1 U34810 ( .A1(STATE_REG_SCAN_IN), .A2(n4220), .ZN(n2988) );
  AOI211_X1 U3482 ( .C1(n5003), .C2(ADDR_REG_1__SCAN_IN), .A(n2989), .B(n2988), 
        .ZN(n2994) );
  MUX2_X1 U34830 ( .A(REG1_REG_1__SCAN_IN), .B(n2990), .S(n2467), .Z(n2992) );
  OAI211_X1 U3484 ( .C1(n2708), .C2(n2992), .A(n5038), .B(n2991), .ZN(n2993)
         );
  OAI211_X1 U34850 ( .C1(n5042), .C2(n2995), .A(n2994), .B(n2993), .ZN(U3241)
         );
  INV_X1 U3486 ( .A(REG3_REG_5__SCAN_IN), .ZN(n4370) );
  NOR2_X1 U34870 ( .A1(STATE_REG_SCAN_IN), .A2(n4370), .ZN(n3226) );
  INV_X1 U3488 ( .A(n2996), .ZN(n2997) );
  AOI211_X1 U34890 ( .C1(n2999), .C2(n2998), .A(n2997), .B(n5031), .ZN(n3000)
         );
  AOI211_X1 U3490 ( .C1(n5003), .C2(ADDR_REG_5__SCAN_IN), .A(n3226), .B(n3000), 
        .ZN(n3005) );
  OAI211_X1 U34910 ( .C1(n3003), .C2(n3002), .A(n5038), .B(n3001), .ZN(n3004)
         );
  OAI211_X1 U3492 ( .C1(n5042), .C2(n3006), .A(n3005), .B(n3004), .ZN(U3245)
         );
  AOI211_X1 U34930 ( .C1(n3009), .C2(n3008), .A(n3007), .B(n5031), .ZN(n3016)
         );
  OAI211_X1 U3494 ( .C1(REG1_REG_3__SCAN_IN), .C2(n3011), .A(n5038), .B(n3010), 
        .ZN(n3014) );
  INV_X1 U34950 ( .A(REG3_REG_3__SCAN_IN), .ZN(n5096) );
  NOR2_X1 U3496 ( .A1(STATE_REG_SCAN_IN), .A2(n5096), .ZN(n3012) );
  AOI21_X1 U34970 ( .B1(n5036), .B2(ADDR_REG_3__SCAN_IN), .A(n3012), .ZN(n3013) );
  OAI211_X1 U3498 ( .C1(n5042), .C2(n5075), .A(n3014), .B(n3013), .ZN(n3015)
         );
  OR2_X1 U34990 ( .A1(n3016), .A2(n3015), .ZN(U3243) );
  AOI211_X1 U3500 ( .C1(n3440), .C2(n3018), .A(n3017), .B(n5031), .ZN(n3024)
         );
  OAI211_X1 U35010 ( .C1(n3020), .C2(REG1_REG_8__SCAN_IN), .A(n5038), .B(n3019), .ZN(n3022) );
  INV_X1 U3502 ( .A(REG3_REG_8__SCAN_IN), .ZN(n4443) );
  NOR2_X1 U35030 ( .A1(STATE_REG_SCAN_IN), .A2(n4443), .ZN(n3321) );
  AOI21_X1 U3504 ( .B1(n5036), .B2(ADDR_REG_8__SCAN_IN), .A(n3321), .ZN(n3021)
         );
  OAI211_X1 U35050 ( .C1(n5042), .C2(n5134), .A(n3022), .B(n3021), .ZN(n3023)
         );
  OR2_X1 U35060 ( .A1(n3024), .A2(n3023), .ZN(U3248) );
  NAND2_X1 U35070 ( .A1(n3087), .A2(n3800), .ZN(n3027) );
  NAND2_X1 U35080 ( .A1(n4113), .A2(n3327), .ZN(n3026) );
  NAND2_X1 U35090 ( .A1(n3027), .A2(n3026), .ZN(n3028) );
  AOI22_X1 U35100 ( .A1(n3087), .A2(n3882), .B1(n4113), .B2(n3844), .ZN(n3029)
         );
  OAI21_X1 U35110 ( .B1(n3030), .B2(n3029), .A(n3142), .ZN(n3042) );
  NAND2_X1 U35120 ( .A1(n3032), .A2(n3031), .ZN(n3037) );
  INV_X1 U35130 ( .A(n3033), .ZN(n3035) );
  NAND2_X1 U35140 ( .A1(n3035), .A2(n3034), .ZN(n3036) );
  NAND2_X1 U35150 ( .A1(n3037), .A2(n3036), .ZN(n3038) );
  INV_X1 U35160 ( .A(n3038), .ZN(n3040) );
  INV_X1 U35170 ( .A(n3042), .ZN(n3039) );
  NAND2_X1 U35180 ( .A1(n3040), .A2(n3039), .ZN(n3143) );
  INV_X1 U35190 ( .A(n3143), .ZN(n3041) );
  AOI21_X1 U35200 ( .B1(n3042), .B2(n3038), .A(n3041), .ZN(n3054) );
  NAND2_X1 U35210 ( .A1(n2967), .A2(n5096), .ZN(n3048) );
  NAND2_X1 U35220 ( .A1(n3043), .A2(REG1_REG_3__SCAN_IN), .ZN(n3047) );
  NAND2_X1 U35230 ( .A1(n3044), .A2(REG0_REG_3__SCAN_IN), .ZN(n3046) );
  NAND2_X1 U35240 ( .A1(n2966), .A2(REG2_REG_3__SCAN_IN), .ZN(n3045) );
  AOI22_X1 U35250 ( .A1(n3049), .A2(n4573), .B1(n4113), .B2(n5237), .ZN(n3053)
         );
  AOI22_X1 U35260 ( .A1(n3051), .A2(n3064), .B1(REG3_REG_2__SCAN_IN), .B2(
        n3050), .ZN(n3052) );
  OAI211_X1 U35270 ( .C1(n3054), .C2(n5192), .A(n3053), .B(n3052), .ZN(U3234)
         );
  AOI211_X1 U35280 ( .C1(n2491), .C2(n3056), .A(n3055), .B(n5031), .ZN(n3063)
         );
  INV_X1 U35290 ( .A(n3326), .ZN(n5143) );
  OAI211_X1 U35300 ( .C1(n3059), .C2(n3058), .A(n5038), .B(n3057), .ZN(n3061)
         );
  AND2_X1 U35310 ( .A1(U3149), .A2(REG3_REG_9__SCAN_IN), .ZN(n3345) );
  AOI21_X1 U35320 ( .B1(n5036), .B2(ADDR_REG_9__SCAN_IN), .A(n3345), .ZN(n3060) );
  OAI211_X1 U35330 ( .C1(n5042), .C2(n5143), .A(n3061), .B(n3060), .ZN(n3062)
         );
  OR2_X1 U35340 ( .A1(n3063), .A2(n3062), .ZN(U3249) );
  NAND2_X1 U35350 ( .A1(n3080), .A2(n3064), .ZN(n4105) );
  XNOR2_X1 U35360 ( .A(n4063), .B(n3107), .ZN(n5062) );
  NAND2_X1 U35370 ( .A1(n3065), .A2(n4940), .ZN(n3066) );
  OR2_X1 U35380 ( .A1(n5056), .A2(n4089), .ZN(n3117) );
  INV_X1 U35390 ( .A(n3117), .ZN(n3067) );
  AND2_X1 U35400 ( .A1(n5258), .A2(n3067), .ZN(n5099) );
  INV_X1 U35410 ( .A(n5099), .ZN(n3700) );
  INV_X1 U35420 ( .A(n4574), .ZN(n3069) );
  NAND2_X1 U35430 ( .A1(n3069), .A2(n3079), .ZN(n4103) );
  XNOR2_X1 U35440 ( .A(n4063), .B(n4103), .ZN(n3075) );
  NAND2_X1 U35450 ( .A1(n4958), .A2(n4957), .ZN(n3072) );
  NAND2_X1 U35460 ( .A1(n4959), .A2(n2576), .ZN(n3071) );
  AOI22_X1 U35470 ( .A1(n4866), .A2(n4574), .B1(n3087), .B2(n4839), .ZN(n3073)
         );
  OAI21_X1 U35480 ( .B1(n3080), .B2(n5283), .A(n3073), .ZN(n3074) );
  AOI21_X1 U35490 ( .B1(n3075), .B2(n5256), .A(n3074), .ZN(n3076) );
  OAI21_X1 U35500 ( .B1(n5062), .B2(n3068), .A(n3076), .ZN(n5063) );
  NAND2_X1 U35510 ( .A1(n5063), .A2(n5258), .ZN(n3085) );
  AND2_X1 U35520 ( .A1(n5258), .A2(n5006), .ZN(n4818) );
  NAND2_X1 U35530 ( .A1(n2973), .A2(n3079), .ZN(n3078) );
  NAND2_X1 U35540 ( .A1(n2941), .A2(n3077), .ZN(n5273) );
  NAND2_X1 U35550 ( .A1(n3078), .A2(n5303), .ZN(n3081) );
  NOR2_X1 U35560 ( .A1(n3081), .A2(n2494), .ZN(n5064) );
  INV_X1 U35570 ( .A(REG2_REG_1__SCAN_IN), .ZN(n3082) );
  OAI22_X1 U35580 ( .A1(n5258), .A2(n3082), .B1(n4220), .B2(n5260), .ZN(n3083)
         );
  AOI21_X1 U35590 ( .B1(n4818), .B2(n5064), .A(n3083), .ZN(n3084) );
  OAI211_X1 U35600 ( .C1(n5062), .C2(n3700), .A(n3085), .B(n3084), .ZN(U3289)
         );
  INV_X1 U35610 ( .A(n3087), .ZN(n4112) );
  NAND2_X1 U35620 ( .A1(n4112), .A2(n4113), .ZN(n4107) );
  INV_X1 U35630 ( .A(n4573), .ZN(n3159) );
  MUX2_X1 U35640 ( .A(n3088), .B(DATAI_3_), .S(n3025), .Z(n5090) );
  NAND2_X1 U35650 ( .A1(n3159), .A2(n5090), .ZN(n4114) );
  INV_X1 U35660 ( .A(n5090), .ZN(n5084) );
  NAND2_X1 U35670 ( .A1(n4573), .A2(n5084), .ZN(n4110) );
  AND2_X1 U35680 ( .A1(n4114), .A2(n4110), .ZN(n5079) );
  NAND2_X1 U35690 ( .A1(n5077), .A2(n4114), .ZN(n3237) );
  NAND2_X1 U35700 ( .A1(n2966), .A2(REG2_REG_4__SCAN_IN), .ZN(n3093) );
  NAND2_X1 U35710 ( .A1(n3043), .A2(REG1_REG_4__SCAN_IN), .ZN(n3092) );
  NOR2_X1 U35720 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n3089) );
  NOR2_X1 U35730 ( .A1(n3095), .A2(n3089), .ZN(n3104) );
  NAND2_X1 U35740 ( .A1(n2967), .A2(n3104), .ZN(n3091) );
  NAND2_X1 U35750 ( .A1(n3044), .A2(REG0_REG_4__SCAN_IN), .ZN(n3090) );
  MUX2_X1 U35760 ( .A(n3094), .B(DATAI_4_), .S(n3025), .Z(n3243) );
  NAND2_X1 U35770 ( .A1(n3923), .A2(n3243), .ZN(n4115) );
  INV_X1 U35780 ( .A(n3923), .ZN(n4572) );
  INV_X1 U35790 ( .A(n3243), .ZN(n3147) );
  NAND2_X1 U35800 ( .A1(n4572), .A2(n3147), .ZN(n4117) );
  XNOR2_X1 U35810 ( .A(n3237), .B(n4079), .ZN(n3102) );
  NAND2_X1 U3582 ( .A1(n2966), .A2(REG2_REG_5__SCAN_IN), .ZN(n3099) );
  NAND2_X1 U3583 ( .A1(n3043), .A2(REG1_REG_5__SCAN_IN), .ZN(n3098) );
  OAI21_X1 U3584 ( .B1(n3095), .B2(REG3_REG_5__SCAN_IN), .A(n3187), .ZN(n3288)
         );
  INV_X1 U3585 ( .A(n3288), .ZN(n3235) );
  NAND2_X1 U3586 ( .A1(n2967), .A2(n3235), .ZN(n3097) );
  NAND2_X1 U3587 ( .A1(n3044), .A2(REG0_REG_5__SCAN_IN), .ZN(n3096) );
  INV_X1 U3588 ( .A(n3246), .ZN(n4571) );
  AOI22_X1 U3589 ( .A1(n4571), .A2(n4839), .B1(n4866), .B2(n4573), .ZN(n3100)
         );
  OAI21_X1 U3590 ( .B1(n3147), .B2(n5283), .A(n3100), .ZN(n3101) );
  AOI21_X1 U3591 ( .B1(n3102), .B2(n5256), .A(n3101), .ZN(n5109) );
  AOI21_X1 U3592 ( .B1(n5087), .B2(n3243), .A(n5273), .ZN(n3103) );
  NAND2_X1 U3593 ( .A1(n3103), .A2(n3287), .ZN(n5108) );
  INV_X1 U3594 ( .A(n5108), .ZN(n3106) );
  INV_X1 U3595 ( .A(n3104), .ZN(n3163) );
  OAI22_X1 U3596 ( .A1(n5258), .A2(n5034), .B1(n3163), .B2(n5260), .ZN(n3105)
         );
  AOI21_X1 U3597 ( .B1(n3106), .B2(n4818), .A(n3105), .ZN(n3120) );
  NAND2_X1 U3598 ( .A1(n3064), .A2(n2973), .ZN(n3108) );
  NAND2_X1 U3599 ( .A1(n3109), .A2(n3108), .ZN(n3123) );
  INV_X1 U3600 ( .A(n3123), .ZN(n3110) );
  NAND2_X1 U3601 ( .A1(n4112), .A2(n3131), .ZN(n3111) );
  NAND2_X1 U3602 ( .A1(n4573), .A2(n5090), .ZN(n3112) );
  NAND2_X1 U3603 ( .A1(n3159), .A2(n5084), .ZN(n3113) );
  INV_X1 U3604 ( .A(n3116), .ZN(n3115) );
  NAND2_X1 U3605 ( .A1(n3115), .A2(n3114), .ZN(n3245) );
  NAND2_X1 U3606 ( .A1(n3116), .A2(n4079), .ZN(n5106) );
  NAND2_X1 U3607 ( .A1(n3068), .A2(n3117), .ZN(n3118) );
  NAND3_X1 U3608 ( .A1(n3245), .A2(n5106), .A3(n5268), .ZN(n3119) );
  OAI211_X1 U3609 ( .C1(n5109), .C2(n5301), .A(n3120), .B(n3119), .ZN(U3286)
         );
  XOR2_X1 U3610 ( .A(n4075), .B(n3121), .Z(n3128) );
  NAND2_X1 U3611 ( .A1(n3123), .A2(n4075), .ZN(n3124) );
  NAND2_X1 U3612 ( .A1(n3122), .A2(n3124), .ZN(n5071) );
  INV_X1 U3613 ( .A(n3068), .ZN(n5086) );
  AOI22_X1 U3614 ( .A1(n3064), .A2(n4866), .B1(n4839), .B2(n4573), .ZN(n3125)
         );
  OAI21_X1 U3615 ( .B1(n3131), .B2(n5283), .A(n3125), .ZN(n3126) );
  AOI21_X1 U3616 ( .B1(n5071), .B2(n5086), .A(n3126), .ZN(n3127) );
  OAI21_X1 U3617 ( .B1(n3128), .B2(n4860), .A(n3127), .ZN(n5069) );
  INV_X1 U3618 ( .A(n5069), .ZN(n3135) );
  INV_X1 U3619 ( .A(n3129), .ZN(n3130) );
  NAND2_X1 U3620 ( .A1(n5258), .A2(n3130), .ZN(n4897) );
  OAI21_X1 U3621 ( .B1(n2494), .B2(n3131), .A(n5089), .ZN(n5068) );
  INV_X1 U3622 ( .A(n5260), .ZN(n5097) );
  AOI22_X1 U3623 ( .A1(n5301), .A2(REG2_REG_2__SCAN_IN), .B1(
        REG3_REG_2__SCAN_IN), .B2(n5097), .ZN(n3132) );
  OAI21_X1 U3624 ( .B1(n4897), .B2(n5068), .A(n3132), .ZN(n3133) );
  AOI21_X1 U3625 ( .B1(n5071), .B2(n5099), .A(n3133), .ZN(n3134) );
  OAI21_X1 U3626 ( .B1(n3135), .B2(n5301), .A(n3134), .ZN(U3288) );
  NAND4_X1 U3627 ( .A1(n3138), .A2(n3137), .A3(n2943), .A4(n3136), .ZN(n3139)
         );
  NAND2_X1 U3628 ( .A1(n3139), .A2(STATE_REG_SCAN_IN), .ZN(n3141) );
  NAND2_X1 U3629 ( .A1(n3143), .A2(n3142), .ZN(n3920) );
  NAND2_X1 U3630 ( .A1(n4573), .A2(n3800), .ZN(n3145) );
  NAND2_X1 U3631 ( .A1(n5090), .A2(n3327), .ZN(n3144) );
  NAND2_X1 U3632 ( .A1(n3145), .A2(n3144), .ZN(n3146) );
  AOI22_X1 U3633 ( .A1(n4573), .A2(n3882), .B1(n5090), .B2(n3844), .ZN(n3152)
         );
  XNOR2_X1 U3634 ( .A(n3151), .B(n3152), .ZN(n3921) );
  NAND2_X1 U3635 ( .A1(n3920), .A2(n3921), .ZN(n3155) );
  OAI22_X1 U3636 ( .A1(n3923), .A2(n2965), .B1(n3147), .B2(n3859), .ZN(n3148)
         );
  XNOR2_X1 U3637 ( .A(n3148), .B(n3879), .ZN(n3172) );
  OR2_X1 U3638 ( .A1(n3923), .A2(n3891), .ZN(n3150) );
  NAND2_X1 U3639 ( .A1(n3243), .A2(n3800), .ZN(n3149) );
  NAND2_X1 U3640 ( .A1(n3150), .A2(n3149), .ZN(n3173) );
  XNOR2_X1 U3641 ( .A(n3172), .B(n3173), .ZN(n3156) );
  INV_X1 U3642 ( .A(n3151), .ZN(n3153) );
  NAND2_X1 U3643 ( .A1(n3153), .A2(n3152), .ZN(n3157) );
  AND2_X1 U3644 ( .A1(n3156), .A2(n3157), .ZN(n3154) );
  INV_X1 U3645 ( .A(n3176), .ZN(n3230) );
  AOI21_X1 U3646 ( .B1(n3155), .B2(n3157), .A(n3156), .ZN(n3158) );
  OR3_X1 U3647 ( .A1(n3230), .A2(n3158), .A3(n5192), .ZN(n3162) );
  INV_X1 U3648 ( .A(REG3_REG_4__SCAN_IN), .ZN(n4447) );
  NOR2_X1 U3649 ( .A1(n4447), .A2(STATE_REG_SCAN_IN), .ZN(n5035) );
  OAI22_X1 U3650 ( .A1(n3159), .A2(n3977), .B1(n3976), .B2(n3246), .ZN(n3160)
         );
  AOI211_X1 U3651 ( .C1(n3243), .C2(n5237), .A(n5035), .B(n3160), .ZN(n3161)
         );
  OAI211_X1 U3652 ( .C1(n5244), .C2(n3163), .A(n3162), .B(n3161), .ZN(U3227)
         );
  MUX2_X1 U3653 ( .A(n4968), .B(DATAI_5_), .S(n3025), .Z(n3286) );
  INV_X1 U3654 ( .A(n3286), .ZN(n3294) );
  OAI22_X1 U3655 ( .A1(n3246), .A2(n2965), .B1(n3294), .B2(n3859), .ZN(n3164)
         );
  XNOR2_X1 U3656 ( .A(n3164), .B(n3879), .ZN(n3167) );
  OR2_X1 U3657 ( .A1(n3246), .A2(n3891), .ZN(n3166) );
  NAND2_X1 U3658 ( .A1(n3286), .A2(n3876), .ZN(n3165) );
  AND2_X1 U3659 ( .A1(n3166), .A2(n3165), .ZN(n3168) );
  NAND2_X1 U3660 ( .A1(n3167), .A2(n3168), .ZN(n3177) );
  INV_X1 U3661 ( .A(n3167), .ZN(n3170) );
  INV_X1 U3662 ( .A(n3168), .ZN(n3169) );
  NAND2_X1 U3663 ( .A1(n3170), .A2(n3169), .ZN(n3171) );
  NAND2_X1 U3664 ( .A1(n3177), .A2(n3171), .ZN(n3228) );
  INV_X1 U3665 ( .A(n3172), .ZN(n3174) );
  AND2_X1 U3666 ( .A1(n3174), .A2(n3173), .ZN(n3229) );
  NOR2_X1 U3667 ( .A1(n3228), .A2(n3229), .ZN(n3175) );
  NAND2_X1 U3668 ( .A1(n3043), .A2(REG1_REG_6__SCAN_IN), .ZN(n3181) );
  NAND2_X1 U3669 ( .A1(n2466), .A2(REG0_REG_6__SCAN_IN), .ZN(n3180) );
  XNOR2_X1 U3670 ( .A(n3187), .B(REG3_REG_6__SCAN_IN), .ZN(n3216) );
  NAND2_X1 U3671 ( .A1(n2967), .A2(n3216), .ZN(n3179) );
  NAND2_X1 U3672 ( .A1(n2966), .A2(REG2_REG_6__SCAN_IN), .ZN(n3178) );
  NAND4_X1 U3673 ( .A1(n3181), .A2(n3180), .A3(n3179), .A4(n3178), .ZN(n4570)
         );
  NAND2_X1 U3674 ( .A1(n4570), .A2(n3876), .ZN(n3183) );
  MUX2_X1 U3675 ( .A(n4967), .B(DATAI_6_), .S(n3025), .Z(n3271) );
  NAND2_X1 U3676 ( .A1(n3271), .A2(n3327), .ZN(n3182) );
  NAND2_X1 U3677 ( .A1(n3183), .A2(n3182), .ZN(n3184) );
  XNOR2_X1 U3678 ( .A(n3184), .B(n3892), .ZN(n3197) );
  AOI22_X1 U3679 ( .A1(n4570), .A2(n3882), .B1(n3271), .B2(n3844), .ZN(n3198)
         );
  XNOR2_X1 U3680 ( .A(n3197), .B(n3198), .ZN(n3218) );
  NAND2_X1 U3681 ( .A1(n3043), .A2(REG1_REG_7__SCAN_IN), .ZN(n3192) );
  NAND2_X1 U3682 ( .A1(n2966), .A2(REG2_REG_7__SCAN_IN), .ZN(n3191) );
  INV_X1 U3683 ( .A(n3187), .ZN(n3185) );
  AOI21_X1 U3684 ( .B1(n3185), .B2(REG3_REG_6__SCAN_IN), .A(
        REG3_REG_7__SCAN_IN), .ZN(n3188) );
  NAND2_X1 U3685 ( .A1(REG3_REG_7__SCAN_IN), .A2(REG3_REG_6__SCAN_IN), .ZN(
        n3186) );
  OR2_X1 U3686 ( .A1(n3188), .A2(n3204), .ZN(n3278) );
  INV_X1 U3687 ( .A(n3278), .ZN(n3212) );
  NAND2_X1 U3688 ( .A1(n2967), .A2(n3212), .ZN(n3190) );
  NAND2_X1 U3689 ( .A1(n3044), .A2(REG0_REG_7__SCAN_IN), .ZN(n3189) );
  MUX2_X1 U3690 ( .A(n3193), .B(DATAI_7_), .S(n3025), .Z(n3433) );
  INV_X1 U3691 ( .A(n3433), .ZN(n3267) );
  OAI22_X1 U3692 ( .A1(n3319), .A2(n2965), .B1(n3267), .B2(n3859), .ZN(n3194)
         );
  XNOR2_X1 U3693 ( .A(n3194), .B(n3879), .ZN(n3299) );
  OR2_X1 U3694 ( .A1(n3319), .A2(n3891), .ZN(n3196) );
  NAND2_X1 U3695 ( .A1(n3433), .A2(n3876), .ZN(n3195) );
  NAND2_X1 U3696 ( .A1(n3196), .A2(n3195), .ZN(n3300) );
  XNOR2_X1 U3697 ( .A(n3299), .B(n3300), .ZN(n3202) );
  INV_X1 U3698 ( .A(n3197), .ZN(n3199) );
  NAND2_X1 U3699 ( .A1(n3199), .A2(n3198), .ZN(n3203) );
  AND2_X1 U3700 ( .A1(n3202), .A2(n3203), .ZN(n3200) );
  NAND2_X1 U3701 ( .A1(n3201), .A2(n3200), .ZN(n3367) );
  NAND2_X1 U3702 ( .A1(n3367), .A2(n5239), .ZN(n3215) );
  AOI21_X1 U3703 ( .B1(n3201), .B2(n3203), .A(n3202), .ZN(n3214) );
  OAI22_X1 U3704 ( .A1(n3975), .A2(n3267), .B1(STATE_REG_SCAN_IN), .B2(n4434), 
        .ZN(n3211) );
  NAND2_X1 U3705 ( .A1(n3204), .A2(REG3_REG_8__SCAN_IN), .ZN(n3313) );
  OR2_X1 U3706 ( .A1(n3204), .A2(REG3_REG_8__SCAN_IN), .ZN(n3205) );
  AND2_X1 U3707 ( .A1(n3313), .A2(n3205), .ZN(n3298) );
  NAND2_X1 U3708 ( .A1(n2967), .A2(n3298), .ZN(n3209) );
  NAND2_X1 U3709 ( .A1(n3043), .A2(REG1_REG_8__SCAN_IN), .ZN(n3208) );
  NAND2_X1 U3710 ( .A1(n2966), .A2(REG2_REG_8__SCAN_IN), .ZN(n3207) );
  NAND2_X1 U3711 ( .A1(n3044), .A2(REG0_REG_8__SCAN_IN), .ZN(n3206) );
  INV_X1 U3712 ( .A(n4568), .ZN(n3507) );
  OAI22_X1 U3713 ( .A1(n3273), .A2(n3977), .B1(n3976), .B2(n3507), .ZN(n3210)
         );
  AOI211_X1 U3714 ( .C1(n3212), .C2(n3980), .A(n3211), .B(n3210), .ZN(n3213)
         );
  OAI21_X1 U3715 ( .B1(n3215), .B2(n3214), .A(n3213), .ZN(U3210) );
  INV_X1 U3716 ( .A(n3216), .ZN(n3249) );
  OAI21_X1 U3717 ( .B1(n3218), .B2(n3217), .A(n3201), .ZN(n3219) );
  NAND2_X1 U3718 ( .A1(n3219), .A2(n5239), .ZN(n3223) );
  OAI22_X1 U3719 ( .A1(n3246), .A2(n3977), .B1(n3976), .B2(n3319), .ZN(n3220)
         );
  AOI211_X1 U3720 ( .C1(n3271), .C2(n5237), .A(n3221), .B(n3220), .ZN(n3222)
         );
  OAI211_X1 U3721 ( .C1(n5244), .C2(n3249), .A(n3223), .B(n3222), .ZN(U3236)
         );
  OR2_X1 U3722 ( .A1(n3923), .A2(n4887), .ZN(n3225) );
  NAND2_X1 U3723 ( .A1(n4570), .A2(n4839), .ZN(n3224) );
  NAND2_X1 U3724 ( .A1(n3225), .A2(n3224), .ZN(n3291) );
  AOI21_X1 U3725 ( .B1(n5231), .B2(n3291), .A(n3226), .ZN(n3227) );
  OAI21_X1 U3726 ( .B1(n3975), .B2(n3294), .A(n3227), .ZN(n3234) );
  OAI21_X1 U3727 ( .B1(n3230), .B2(n3229), .A(n3228), .ZN(n3232) );
  AOI21_X1 U3728 ( .B1(n3232), .B2(n3231), .A(n5192), .ZN(n3233) );
  AOI211_X1 U3729 ( .C1(n3235), .C2(n3980), .A(n3234), .B(n3233), .ZN(n3236)
         );
  INV_X1 U3730 ( .A(n3236), .ZN(U3224) );
  NAND2_X1 U3731 ( .A1(n3246), .A2(n3286), .ZN(n4093) );
  NAND2_X1 U3732 ( .A1(n4571), .A2(n3294), .ZN(n3265) );
  NAND2_X1 U3733 ( .A1(n4093), .A2(n3265), .ZN(n3289) );
  NAND2_X1 U3734 ( .A1(n3290), .A2(n3265), .ZN(n3238) );
  NAND2_X1 U3735 ( .A1(n3273), .A2(n3271), .ZN(n4120) );
  NAND2_X1 U3736 ( .A1(n4570), .A2(n3272), .ZN(n4094) );
  NAND2_X1 U3737 ( .A1(n4120), .A2(n4094), .ZN(n4058) );
  XNOR2_X1 U3738 ( .A(n3238), .B(n4058), .ZN(n3239) );
  NAND2_X1 U3739 ( .A1(n3239), .A2(n5256), .ZN(n3242) );
  OAI22_X1 U3740 ( .A1(n3246), .A2(n4887), .B1(n3319), .B2(n5048), .ZN(n3240)
         );
  INV_X1 U3741 ( .A(n3240), .ZN(n3241) );
  OAI211_X1 U3742 ( .C1(n5283), .C2(n3272), .A(n3242), .B(n3241), .ZN(n5121)
         );
  INV_X1 U3743 ( .A(n5121), .ZN(n3254) );
  NAND2_X1 U3744 ( .A1(n4572), .A2(n3243), .ZN(n3244) );
  NAND2_X1 U3745 ( .A1(n3246), .A2(n3294), .ZN(n3247) );
  XNOR2_X1 U3746 ( .A(n3275), .B(n4058), .ZN(n5123) );
  OAI21_X1 U3747 ( .B1(n3248), .B2(n3272), .A(n3277), .ZN(n5120) );
  NOR2_X1 U3748 ( .A1(n5120), .A2(n4897), .ZN(n3252) );
  OAI22_X1 U3749 ( .A1(n5258), .A2(n3250), .B1(n3249), .B2(n5260), .ZN(n3251)
         );
  AOI211_X1 U3750 ( .C1(n5123), .C2(n5268), .A(n3252), .B(n3251), .ZN(n3253)
         );
  OAI21_X1 U3751 ( .B1(n5301), .B2(n3254), .A(n3253), .ZN(U3284) );
  AOI211_X1 U3752 ( .C1(n3257), .C2(n3256), .A(n3255), .B(n5031), .ZN(n3264)
         );
  OAI211_X1 U3753 ( .C1(n3259), .C2(REG1_REG_10__SCAN_IN), .A(n5038), .B(n3258), .ZN(n3262) );
  NOR2_X1 U3754 ( .A1(STATE_REG_SCAN_IN), .A2(n3402), .ZN(n3260) );
  AOI21_X1 U3755 ( .B1(n5003), .B2(ADDR_REG_10__SCAN_IN), .A(n3260), .ZN(n3261) );
  OAI211_X1 U3756 ( .C1(n5042), .C2(n5151), .A(n3262), .B(n3261), .ZN(n3263)
         );
  OR2_X1 U3757 ( .A1(n3264), .A2(n3263), .ZN(U3250) );
  AND2_X1 U3758 ( .A1(n3265), .A2(n4094), .ZN(n4118) );
  NAND2_X1 U3759 ( .A1(n3266), .A2(n4120), .ZN(n3443) );
  NAND2_X1 U3760 ( .A1(n3319), .A2(n3433), .ZN(n4121) );
  INV_X1 U3761 ( .A(n3319), .ZN(n4569) );
  NAND2_X1 U3762 ( .A1(n4569), .A2(n3267), .ZN(n3490) );
  NAND2_X1 U3763 ( .A1(n4121), .A2(n3490), .ZN(n3508) );
  XNOR2_X1 U3764 ( .A(n3443), .B(n3508), .ZN(n3270) );
  OAI22_X1 U3765 ( .A1(n3273), .A2(n4887), .B1(n3507), .B2(n5048), .ZN(n3268)
         );
  AOI21_X1 U3766 ( .B1(n3433), .B2(n5292), .A(n3268), .ZN(n3269) );
  OAI21_X1 U3767 ( .B1(n3270), .B2(n4860), .A(n3269), .ZN(n5128) );
  INV_X1 U3768 ( .A(n5128), .ZN(n3283) );
  NOR2_X1 U3769 ( .A1(n4570), .A2(n3271), .ZN(n3274) );
  INV_X1 U3770 ( .A(n3508), .ZN(n4082) );
  XNOR2_X1 U3771 ( .A(n3547), .B(n4082), .ZN(n5130) );
  NAND2_X1 U3772 ( .A1(n5130), .A2(n5268), .ZN(n3282) );
  INV_X1 U3773 ( .A(n3437), .ZN(n3276) );
  AOI211_X1 U3774 ( .C1(n3433), .C2(n3277), .A(n5273), .B(n3276), .ZN(n5129)
         );
  INV_X1 U3775 ( .A(REG2_REG_7__SCAN_IN), .ZN(n3279) );
  OAI22_X1 U3776 ( .A1(n5258), .A2(n3279), .B1(n3278), .B2(n5260), .ZN(n3280)
         );
  AOI21_X1 U3777 ( .B1(n5129), .B2(n4818), .A(n3280), .ZN(n3281) );
  OAI211_X1 U3778 ( .C1(n3283), .C2(n5301), .A(n3282), .B(n3281), .ZN(U3283)
         );
  OAI21_X1 U3779 ( .B1(n3284), .B2(n3289), .A(n3285), .ZN(n5116) );
  XNOR2_X1 U3780 ( .A(n3287), .B(n3286), .ZN(n5113) );
  OAI22_X1 U3781 ( .A1(n5113), .A2(n4897), .B1(n3288), .B2(n5260), .ZN(n3296)
         );
  INV_X1 U3782 ( .A(n3289), .ZN(n4081) );
  OAI211_X1 U3783 ( .C1(n2492), .C2(n4081), .A(n3290), .B(n5256), .ZN(n3293)
         );
  INV_X1 U3784 ( .A(n3291), .ZN(n3292) );
  OAI211_X1 U3785 ( .C1(n5283), .C2(n3294), .A(n3293), .B(n3292), .ZN(n5114)
         );
  MUX2_X1 U3786 ( .A(n5114), .B(REG2_REG_5__SCAN_IN), .S(n5301), .Z(n3295) );
  AOI211_X1 U3787 ( .C1(n5268), .C2(n5116), .A(n3296), .B(n3295), .ZN(n3297)
         );
  INV_X1 U3788 ( .A(n3297), .ZN(U3285) );
  INV_X1 U3789 ( .A(n3298), .ZN(n3439) );
  INV_X1 U3790 ( .A(n3367), .ZN(n3308) );
  INV_X1 U3791 ( .A(n3299), .ZN(n3301) );
  AND2_X1 U3792 ( .A1(n3301), .A2(n3300), .ZN(n3310) );
  NAND2_X1 U3793 ( .A1(n4568), .A2(n3876), .ZN(n3304) );
  MUX2_X1 U3794 ( .A(n3302), .B(DATAI_8_), .S(n3025), .Z(n3438) );
  NAND2_X1 U3795 ( .A1(n3438), .A2(n3327), .ZN(n3303) );
  NAND2_X1 U3796 ( .A1(n3304), .A2(n3303), .ZN(n3305) );
  XNOR2_X1 U3797 ( .A(n3305), .B(n3879), .ZN(n3307) );
  AOI22_X1 U3798 ( .A1(n4568), .A2(n3882), .B1(n3438), .B2(n3844), .ZN(n3306)
         );
  NAND2_X1 U3799 ( .A1(n3307), .A2(n3306), .ZN(n3333) );
  OAI21_X1 U3800 ( .B1(n3307), .B2(n3306), .A(n3333), .ZN(n3309) );
  OAI21_X1 U3801 ( .B1(n3308), .B2(n3310), .A(n3309), .ZN(n3311) );
  NOR2_X1 U3802 ( .A1(n3310), .A2(n3309), .ZN(n3332) );
  NAND2_X1 U3803 ( .A1(n3367), .A2(n3332), .ZN(n3331) );
  AOI21_X1 U3804 ( .B1(n3311), .B2(n3331), .A(n5192), .ZN(n3312) );
  INV_X1 U3805 ( .A(n3312), .ZN(n3323) );
  NAND2_X1 U3806 ( .A1(n2966), .A2(REG2_REG_9__SCAN_IN), .ZN(n3318) );
  NAND2_X1 U3807 ( .A1(n3043), .A2(REG1_REG_9__SCAN_IN), .ZN(n3317) );
  NAND2_X1 U3808 ( .A1(n3313), .A2(n4234), .ZN(n3314) );
  AND2_X1 U3809 ( .A1(n3338), .A2(n3314), .ZN(n3324) );
  NAND2_X1 U3810 ( .A1(n2967), .A2(n3324), .ZN(n3316) );
  NAND2_X1 U3811 ( .A1(n2466), .A2(REG0_REG_9__SCAN_IN), .ZN(n3315) );
  INV_X1 U3812 ( .A(n3325), .ZN(n3492) );
  OAI22_X1 U3813 ( .A1(n3319), .A2(n3977), .B1(n3976), .B2(n3492), .ZN(n3320)
         );
  AOI211_X1 U3814 ( .C1(n3438), .C2(n5237), .A(n3321), .B(n3320), .ZN(n3322)
         );
  OAI211_X1 U3815 ( .C1(n5244), .C2(n3439), .A(n3323), .B(n3322), .ZN(U3218)
         );
  INV_X1 U3816 ( .A(n3324), .ZN(n3502) );
  NAND2_X1 U3817 ( .A1(n3325), .A2(n3876), .ZN(n3329) );
  MUX2_X1 U3818 ( .A(n3326), .B(DATAI_9_), .S(n4000), .Z(n3498) );
  NAND2_X1 U3819 ( .A1(n3498), .A2(n3327), .ZN(n3328) );
  AOI22_X1 U3820 ( .A1(n3325), .A2(n3882), .B1(n3498), .B2(n3844), .ZN(n3372)
         );
  XNOR2_X1 U3821 ( .A(n3371), .B(n3372), .ZN(n3336) );
  NAND2_X1 U3822 ( .A1(n3331), .A2(n3333), .ZN(n3335) );
  AND2_X1 U3823 ( .A1(n3336), .A2(n3332), .ZN(n3365) );
  NAND2_X1 U3824 ( .A1(n3367), .A2(n3365), .ZN(n3378) );
  INV_X1 U3825 ( .A(n3336), .ZN(n3334) );
  OR2_X1 U3826 ( .A1(n3334), .A2(n3333), .ZN(n3375) );
  AND2_X1 U3827 ( .A1(n3378), .A2(n3375), .ZN(n3398) );
  OAI21_X1 U3828 ( .B1(n3336), .B2(n3335), .A(n3398), .ZN(n3337) );
  NAND2_X1 U3829 ( .A1(n3337), .A2(n5239), .ZN(n3347) );
  NAND2_X1 U3830 ( .A1(n2966), .A2(REG2_REG_10__SCAN_IN), .ZN(n3343) );
  NAND2_X1 U3831 ( .A1(n3043), .A2(REG1_REG_10__SCAN_IN), .ZN(n3342) );
  AND2_X1 U3832 ( .A1(n3338), .A2(n3402), .ZN(n3339) );
  NOR2_X1 U3833 ( .A1(n3385), .A2(n3339), .ZN(n3555) );
  NAND2_X1 U3834 ( .A1(n2967), .A2(n3555), .ZN(n3341) );
  NAND2_X1 U3835 ( .A1(n2466), .A2(REG0_REG_10__SCAN_IN), .ZN(n3340) );
  OAI22_X1 U3836 ( .A1(n3507), .A2(n4887), .B1(n3536), .B2(n5048), .ZN(n3497)
         );
  NOR2_X1 U3837 ( .A1(n3975), .A2(n3500), .ZN(n3344) );
  AOI211_X1 U3838 ( .C1(n5231), .C2(n3497), .A(n3345), .B(n3344), .ZN(n3346)
         );
  OAI211_X1 U3839 ( .C1(n5244), .C2(n3502), .A(n3347), .B(n3346), .ZN(U3228)
         );
  INV_X1 U3840 ( .A(REG3_REG_11__SCAN_IN), .ZN(n3348) );
  XNOR2_X1 U3841 ( .A(n3385), .B(n3348), .ZN(n3349) );
  INV_X1 U3842 ( .A(n3349), .ZN(n3571) );
  NAND2_X1 U3843 ( .A1(n2966), .A2(REG2_REG_11__SCAN_IN), .ZN(n3353) );
  NAND2_X1 U3844 ( .A1(n3043), .A2(REG1_REG_11__SCAN_IN), .ZN(n3352) );
  NAND2_X1 U3845 ( .A1(n2967), .A2(n3349), .ZN(n3351) );
  NAND2_X1 U3846 ( .A1(n3044), .A2(REG0_REG_11__SCAN_IN), .ZN(n3350) );
  MUX2_X1 U3847 ( .A(n4966), .B(DATAI_11_), .S(n3025), .Z(n3576) );
  OAI22_X1 U3848 ( .A1(n3630), .A2(n2965), .B1(n3629), .B2(n3859), .ZN(n3354)
         );
  XNOR2_X1 U3849 ( .A(n3354), .B(n3879), .ZN(n3358) );
  OR2_X1 U3850 ( .A1(n3630), .A2(n3891), .ZN(n3356) );
  NAND2_X1 U3851 ( .A1(n3576), .A2(n3876), .ZN(n3355) );
  AND2_X1 U3852 ( .A1(n3356), .A2(n3355), .ZN(n3357) );
  NAND2_X1 U3853 ( .A1(n3358), .A2(n3357), .ZN(n3418) );
  NAND2_X1 U3854 ( .A1(n3418), .A2(n3359), .ZN(n3380) );
  MUX2_X1 U3855 ( .A(n3360), .B(DATAI_10_), .S(n4000), .Z(n3560) );
  OAI22_X1 U3856 ( .A1(n3536), .A2(n2965), .B1(n3567), .B2(n3859), .ZN(n3361)
         );
  XNOR2_X1 U3857 ( .A(n3361), .B(n3879), .ZN(n3370) );
  INV_X1 U3858 ( .A(n3370), .ZN(n3364) );
  OR2_X1 U3859 ( .A1(n3536), .A2(n3891), .ZN(n3363) );
  NAND2_X1 U3860 ( .A1(n3560), .A2(n3876), .ZN(n3362) );
  NAND2_X1 U3861 ( .A1(n3363), .A2(n3362), .ZN(n3369) );
  AND2_X1 U3862 ( .A1(n3364), .A2(n3369), .ZN(n3379) );
  AND2_X1 U3863 ( .A1(n3365), .A2(n3368), .ZN(n3366) );
  NAND2_X1 U3864 ( .A1(n3367), .A2(n3366), .ZN(n3421) );
  XNOR2_X1 U3865 ( .A(n3370), .B(n3369), .ZN(n3400) );
  INV_X1 U3866 ( .A(n3371), .ZN(n3373) );
  NAND2_X1 U3867 ( .A1(n3373), .A2(n3372), .ZN(n3397) );
  AND2_X1 U3868 ( .A1(n3400), .A2(n3397), .ZN(n3374) );
  NAND2_X1 U3869 ( .A1(n3421), .A2(n3419), .ZN(n3417) );
  NAND2_X1 U3870 ( .A1(n3378), .A2(n3377), .ZN(n3399) );
  INV_X1 U3871 ( .A(n3379), .ZN(n3382) );
  INV_X1 U3872 ( .A(n3380), .ZN(n3381) );
  AOI21_X1 U3873 ( .B1(n3399), .B2(n3382), .A(n3381), .ZN(n3383) );
  OAI21_X1 U3874 ( .B1(n3417), .B2(n3383), .A(n5239), .ZN(n3396) );
  NAND2_X1 U3875 ( .A1(n2966), .A2(REG2_REG_12__SCAN_IN), .ZN(n3391) );
  NAND2_X1 U3876 ( .A1(n3043), .A2(REG1_REG_12__SCAN_IN), .ZN(n3390) );
  AND2_X1 U3877 ( .A1(REG3_REG_12__SCAN_IN), .A2(REG3_REG_11__SCAN_IN), .ZN(
        n3384) );
  AOI21_X1 U3878 ( .B1(n3385), .B2(REG3_REG_11__SCAN_IN), .A(
        REG3_REG_12__SCAN_IN), .ZN(n3386) );
  OR2_X1 U3879 ( .A1(n3425), .A2(n3386), .ZN(n3625) );
  INV_X1 U3880 ( .A(n3625), .ZN(n3387) );
  NAND2_X1 U3881 ( .A1(n2967), .A2(n3387), .ZN(n3389) );
  NAND2_X1 U3882 ( .A1(n2466), .A2(REG0_REG_12__SCAN_IN), .ZN(n3388) );
  OR2_X1 U3883 ( .A1(n3638), .A2(n5048), .ZN(n3393) );
  OR2_X1 U3884 ( .A1(n3536), .A2(n4887), .ZN(n3392) );
  NAND2_X1 U3885 ( .A1(n3393), .A2(n3392), .ZN(n3575) );
  AND2_X1 U3886 ( .A1(U3149), .A2(REG3_REG_11__SCAN_IN), .ZN(n3485) );
  NOR2_X1 U3887 ( .A1(n3975), .A2(n3629), .ZN(n3394) );
  AOI211_X1 U3888 ( .C1(n5231), .C2(n3575), .A(n3485), .B(n3394), .ZN(n3395)
         );
  OAI211_X1 U3889 ( .C1(n5244), .C2(n3571), .A(n3396), .B(n3395), .ZN(U3233)
         );
  INV_X1 U3890 ( .A(n3555), .ZN(n3407) );
  AND2_X1 U3891 ( .A1(n3398), .A2(n3397), .ZN(n3401) );
  OAI211_X1 U3892 ( .C1(n3401), .C2(n3400), .A(n5239), .B(n3399), .ZN(n3406)
         );
  INV_X1 U3893 ( .A(n3630), .ZN(n4566) );
  AOI22_X1 U3894 ( .A1(n4566), .A2(n4839), .B1(n4866), .B2(n3325), .ZN(n3553)
         );
  OAI22_X1 U3895 ( .A1(n3553), .A2(n3403), .B1(STATE_REG_SCAN_IN), .B2(n3402), 
        .ZN(n3404) );
  AOI21_X1 U3896 ( .B1(n3560), .B2(n5237), .A(n3404), .ZN(n3405) );
  OAI211_X1 U3897 ( .C1(n5244), .C2(n3407), .A(n3406), .B(n3405), .ZN(U3214)
         );
  INV_X1 U3898 ( .A(n3418), .ZN(n3416) );
  MUX2_X1 U3899 ( .A(n4965), .B(DATAI_12_), .S(n3025), .Z(n3624) );
  INV_X1 U3900 ( .A(n3624), .ZN(n3637) );
  OAI22_X1 U3901 ( .A1(n3638), .A2(n2965), .B1(n3637), .B2(n3859), .ZN(n3408)
         );
  XNOR2_X1 U3902 ( .A(n3408), .B(n3879), .ZN(n3411) );
  OR2_X1 U3903 ( .A1(n3638), .A2(n3891), .ZN(n3410) );
  NAND2_X1 U3904 ( .A1(n3624), .A2(n3876), .ZN(n3409) );
  AND2_X1 U3905 ( .A1(n3410), .A2(n3409), .ZN(n3412) );
  NAND2_X1 U3906 ( .A1(n3411), .A2(n3412), .ZN(n3460) );
  INV_X1 U3907 ( .A(n3411), .ZN(n3414) );
  INV_X1 U3908 ( .A(n3412), .ZN(n3413) );
  NAND2_X1 U3909 ( .A1(n3414), .A2(n3413), .ZN(n3415) );
  AND2_X1 U3910 ( .A1(n3460), .A2(n3415), .ZN(n3422) );
  NOR3_X1 U3911 ( .A1(n3417), .A2(n3416), .A3(n3422), .ZN(n3424) );
  AND2_X1 U3912 ( .A1(n3419), .A2(n3418), .ZN(n3420) );
  NAND2_X1 U3913 ( .A1(n3421), .A2(n3420), .ZN(n3423) );
  NAND2_X1 U3914 ( .A1(n3423), .A2(n3422), .ZN(n3461) );
  INV_X1 U3915 ( .A(n3461), .ZN(n3459) );
  OAI21_X1 U3916 ( .B1(n3424), .B2(n3459), .A(n5239), .ZN(n3432) );
  AND2_X1 U3917 ( .A1(REG3_REG_12__SCAN_IN), .A2(U3149), .ZN(n4576) );
  OAI21_X1 U3918 ( .B1(n3425), .B2(REG3_REG_13__SCAN_IN), .A(n3466), .ZN(n3476) );
  INV_X1 U3919 ( .A(n3476), .ZN(n3697) );
  NAND2_X1 U3920 ( .A1(n2967), .A2(n3697), .ZN(n3429) );
  NAND2_X1 U3921 ( .A1(n3043), .A2(REG1_REG_13__SCAN_IN), .ZN(n3428) );
  NAND2_X1 U3922 ( .A1(n3044), .A2(REG0_REG_13__SCAN_IN), .ZN(n3427) );
  NAND2_X1 U3923 ( .A1(n2966), .A2(REG2_REG_13__SCAN_IN), .ZN(n3426) );
  OAI22_X1 U3924 ( .A1(n3630), .A2(n3977), .B1(n3976), .B2(n3677), .ZN(n3430)
         );
  AOI211_X1 U3925 ( .C1(n3624), .C2(n5237), .A(n4576), .B(n3430), .ZN(n3431)
         );
  OAI211_X1 U3926 ( .C1(n5244), .C2(n3625), .A(n3432), .B(n3431), .ZN(U3221)
         );
  INV_X1 U3927 ( .A(n3438), .ZN(n3506) );
  INV_X1 U3928 ( .A(n3510), .ZN(n4076) );
  NAND2_X1 U3929 ( .A1(n3547), .A2(n3508), .ZN(n3434) );
  NAND2_X1 U3930 ( .A1(n4569), .A2(n3433), .ZN(n3511) );
  NAND2_X1 U3931 ( .A1(n3434), .A2(n3511), .ZN(n3436) );
  NOR2_X1 U3932 ( .A1(n3436), .A2(n4076), .ZN(n3435) );
  AOI21_X1 U3933 ( .B1(n4076), .B2(n3436), .A(n3435), .ZN(n5135) );
  AOI21_X1 U3934 ( .B1(n3438), .B2(n3437), .A(n3501), .ZN(n5138) );
  INV_X2 U3935 ( .A(n5301), .ZN(n5258) );
  OAI22_X1 U3936 ( .A1(n5258), .A2(n3440), .B1(n3439), .B2(n5260), .ZN(n3441)
         );
  AOI21_X1 U3937 ( .B1(n5138), .B2(n5298), .A(n3441), .ZN(n3449) );
  INV_X1 U3938 ( .A(n4121), .ZN(n3442) );
  OR2_X2 U3939 ( .A1(n3443), .A2(n3442), .ZN(n3491) );
  NAND2_X1 U3940 ( .A1(n3491), .A2(n3490), .ZN(n3444) );
  XNOR2_X1 U3941 ( .A(n3444), .B(n3510), .ZN(n3445) );
  NAND2_X1 U3942 ( .A1(n3445), .A2(n5256), .ZN(n3447) );
  AOI22_X1 U3943 ( .A1(n4569), .A2(n4866), .B1(n4839), .B2(n3325), .ZN(n3446)
         );
  OAI211_X1 U3944 ( .C1(n5283), .C2(n3506), .A(n3447), .B(n3446), .ZN(n5137)
         );
  NAND2_X1 U3945 ( .A1(n5137), .A2(n5258), .ZN(n3448) );
  OAI211_X1 U3946 ( .C1(n5135), .C2(n4876), .A(n3449), .B(n3448), .ZN(U3282)
         );
  INV_X1 U3947 ( .A(n3460), .ZN(n3458) );
  MUX2_X1 U3948 ( .A(n4964), .B(DATAI_13_), .S(n3025), .Z(n3686) );
  INV_X1 U3949 ( .A(n3686), .ZN(n3687) );
  OAI22_X1 U3950 ( .A1(n3677), .A2(n2965), .B1(n3687), .B2(n3859), .ZN(n3450)
         );
  XNOR2_X1 U3951 ( .A(n3450), .B(n3879), .ZN(n3453) );
  OR2_X1 U3952 ( .A1(n3677), .A2(n3891), .ZN(n3452) );
  NAND2_X1 U3953 ( .A1(n3686), .A2(n3876), .ZN(n3451) );
  AND2_X1 U3954 ( .A1(n3452), .A2(n3451), .ZN(n3454) );
  NAND2_X1 U3955 ( .A1(n3453), .A2(n3454), .ZN(n3522) );
  INV_X1 U3956 ( .A(n3453), .ZN(n3456) );
  INV_X1 U3957 ( .A(n3454), .ZN(n3455) );
  NAND2_X1 U3958 ( .A1(n3456), .A2(n3455), .ZN(n3457) );
  AND2_X1 U3959 ( .A1(n3522), .A2(n3457), .ZN(n3462) );
  NOR3_X1 U3960 ( .A1(n3459), .A2(n3458), .A3(n3462), .ZN(n3465) );
  NAND2_X1 U3961 ( .A1(n3461), .A2(n3460), .ZN(n3463) );
  NAND2_X1 U3962 ( .A1(n3463), .A2(n3462), .ZN(n3523) );
  INV_X1 U3963 ( .A(n3523), .ZN(n3464) );
  OAI21_X1 U3964 ( .B1(n3465), .B2(n3464), .A(n5239), .ZN(n3475) );
  INV_X1 U3965 ( .A(REG3_REG_14__SCAN_IN), .ZN(n3527) );
  AOI21_X1 U3966 ( .B1(n3466), .B2(n3527), .A(n3528), .ZN(n3518) );
  NAND2_X1 U3967 ( .A1(n2967), .A2(n3518), .ZN(n3470) );
  NAND2_X1 U3968 ( .A1(n3043), .A2(REG1_REG_14__SCAN_IN), .ZN(n3469) );
  NAND2_X1 U3969 ( .A1(n3044), .A2(REG0_REG_14__SCAN_IN), .ZN(n3468) );
  NAND2_X1 U3970 ( .A1(n2966), .A2(REG2_REG_14__SCAN_IN), .ZN(n3467) );
  OR2_X1 U3971 ( .A1(n3702), .A2(n5048), .ZN(n3472) );
  OR2_X1 U3972 ( .A1(n3638), .A2(n4887), .ZN(n3471) );
  NAND2_X1 U3973 ( .A1(n3472), .A2(n3471), .ZN(n3688) );
  INV_X1 U3974 ( .A(REG3_REG_13__SCAN_IN), .ZN(n4451) );
  NOR2_X1 U3975 ( .A1(STATE_REG_SCAN_IN), .A2(n4451), .ZN(n4596) );
  NOR2_X1 U3976 ( .A1(n3975), .A2(n3687), .ZN(n3473) );
  AOI211_X1 U3977 ( .C1(n5231), .C2(n3688), .A(n4596), .B(n3473), .ZN(n3474)
         );
  OAI211_X1 U3978 ( .C1(n3476), .C2(n5244), .A(n3475), .B(n3474), .ZN(U3231)
         );
  OAI211_X1 U3979 ( .C1(n3479), .C2(n3478), .A(n3477), .B(n5038), .ZN(n3487)
         );
  INV_X1 U3980 ( .A(n3480), .ZN(n3481) );
  AOI211_X1 U3981 ( .C1(n3483), .C2(n3482), .A(n3481), .B(n5031), .ZN(n3484)
         );
  AOI211_X1 U3982 ( .C1(n5036), .C2(ADDR_REG_11__SCAN_IN), .A(n3485), .B(n3484), .ZN(n3486) );
  OAI211_X1 U3983 ( .C1(n5042), .C2(n3488), .A(n3487), .B(n3486), .ZN(U3251)
         );
  NAND2_X1 U3984 ( .A1(n4568), .A2(n3506), .ZN(n3489) );
  NOR2_X1 U3985 ( .A1(n4568), .A2(n3506), .ZN(n4124) );
  NAND2_X1 U3986 ( .A1(n3492), .A2(n3498), .ZN(n4123) );
  NAND2_X1 U3987 ( .A1(n3493), .A2(n4123), .ZN(n3551) );
  INV_X1 U3988 ( .A(n3551), .ZN(n3495) );
  NAND2_X1 U3989 ( .A1(n3325), .A2(n3500), .ZN(n4128) );
  NAND2_X1 U3990 ( .A1(n3492), .A2(n3500), .ZN(n3538) );
  NAND2_X1 U3991 ( .A1(n3325), .A2(n3498), .ZN(n3539) );
  NAND2_X1 U3992 ( .A1(n3538), .A2(n3539), .ZN(n4059) );
  OAI21_X1 U3993 ( .B1(n3493), .B2(n4059), .A(n5256), .ZN(n3494) );
  AOI21_X1 U3994 ( .B1(n3495), .B2(n4128), .A(n3494), .ZN(n3496) );
  AOI211_X1 U3995 ( .C1(n5292), .C2(n3498), .A(n3497), .B(n3496), .ZN(n5144)
         );
  INV_X1 U3996 ( .A(n3569), .ZN(n3499) );
  OAI21_X1 U3997 ( .B1(n3501), .B2(n3500), .A(n3499), .ZN(n5145) );
  INV_X1 U3998 ( .A(n5145), .ZN(n3505) );
  INV_X1 U3999 ( .A(REG2_REG_9__SCAN_IN), .ZN(n3503) );
  OAI22_X1 U4000 ( .A1(n5258), .A2(n3503), .B1(n3502), .B2(n5260), .ZN(n3504)
         );
  AOI21_X1 U4001 ( .B1(n3505), .B2(n5298), .A(n3504), .ZN(n3517) );
  NAND2_X1 U4002 ( .A1(n3507), .A2(n3506), .ZN(n3509) );
  AND2_X1 U4003 ( .A1(n3508), .A2(n3509), .ZN(n3537) );
  NAND2_X1 U4004 ( .A1(n3547), .A2(n3537), .ZN(n3514) );
  INV_X1 U4005 ( .A(n3509), .ZN(n3513) );
  AND2_X1 U4006 ( .A1(n3511), .A2(n3510), .ZN(n3512) );
  OR2_X1 U4007 ( .A1(n3513), .A2(n3512), .ZN(n3540) );
  AND2_X1 U4008 ( .A1(n3514), .A2(n3540), .ZN(n3515) );
  XOR2_X1 U4009 ( .A(n4059), .B(n3515), .Z(n5147) );
  NAND2_X1 U4010 ( .A1(n5147), .A2(n5268), .ZN(n3516) );
  OAI211_X1 U4011 ( .C1(n5144), .C2(n5301), .A(n3517), .B(n3516), .ZN(U3281)
         );
  INV_X1 U4012 ( .A(n3518), .ZN(n3655) );
  INV_X1 U4013 ( .A(n3665), .ZN(n3654) );
  OAI22_X1 U4014 ( .A1(n3702), .A2(n2965), .B1(n3654), .B2(n3859), .ZN(n3519)
         );
  XNOR2_X1 U4015 ( .A(n3519), .B(n3879), .ZN(n3583) );
  OR2_X1 U4016 ( .A1(n3702), .A2(n3891), .ZN(n3521) );
  NAND2_X1 U4017 ( .A1(n3665), .A2(n3876), .ZN(n3520) );
  NAND2_X1 U4018 ( .A1(n3521), .A2(n3520), .ZN(n3581) );
  XNOR2_X1 U4019 ( .A(n3583), .B(n3581), .ZN(n3525) );
  OAI21_X1 U4020 ( .B1(n3525), .B2(n3524), .A(n3594), .ZN(n3526) );
  NAND2_X1 U4021 ( .A1(n3526), .A2(n5239), .ZN(n3535) );
  NOR2_X1 U4022 ( .A1(STATE_REG_SCAN_IN), .A2(n3527), .ZN(n4601) );
  NAND2_X1 U4023 ( .A1(n3528), .A2(REG3_REG_15__SCAN_IN), .ZN(n3585) );
  OAI21_X1 U4024 ( .B1(n3528), .B2(REG3_REG_15__SCAN_IN), .A(n3585), .ZN(n5199) );
  INV_X1 U4025 ( .A(n5199), .ZN(n3713) );
  NAND2_X1 U4026 ( .A1(n2967), .A2(n3713), .ZN(n3532) );
  NAND2_X1 U4027 ( .A1(n3043), .A2(REG1_REG_15__SCAN_IN), .ZN(n3531) );
  NAND2_X1 U4028 ( .A1(n2466), .A2(REG0_REG_15__SCAN_IN), .ZN(n3530) );
  NAND2_X1 U4029 ( .A1(n2966), .A2(REG2_REG_15__SCAN_IN), .ZN(n3529) );
  OAI22_X1 U4030 ( .A1(n3668), .A2(n3976), .B1(n3977), .B2(n3677), .ZN(n3533)
         );
  AOI211_X1 U4031 ( .C1(n3665), .C2(n5237), .A(n4601), .B(n3533), .ZN(n3534)
         );
  OAI211_X1 U4032 ( .C1(n5244), .C2(n3655), .A(n3535), .B(n3534), .ZN(U3212)
         );
  NAND2_X1 U4033 ( .A1(n3536), .A2(n3560), .ZN(n4098) );
  INV_X1 U4034 ( .A(n3536), .ZN(n4567) );
  NAND2_X1 U4035 ( .A1(n4567), .A2(n3567), .ZN(n3643) );
  AND2_X1 U4036 ( .A1(n3537), .A2(n3538), .ZN(n3545) );
  NAND2_X1 U4037 ( .A1(n3547), .A2(n3545), .ZN(n3543) );
  INV_X1 U4038 ( .A(n3538), .ZN(n3542) );
  AND2_X1 U4039 ( .A1(n3540), .A2(n3539), .ZN(n3541) );
  AND2_X1 U4040 ( .A1(n3543), .A2(n3548), .ZN(n3550) );
  INV_X1 U4041 ( .A(n4080), .ZN(n3544) );
  AND2_X1 U4042 ( .A1(n3545), .A2(n3544), .ZN(n3546) );
  NAND2_X1 U40430 ( .A1(n3547), .A2(n3546), .ZN(n3627) );
  AOI21_X1 U4044 ( .B1(n4080), .B2(n3550), .A(n2493), .ZN(n5155) );
  INV_X1 U4045 ( .A(n5155), .ZN(n3559) );
  NAND2_X1 U4046 ( .A1(n3551), .A2(n4128), .ZN(n3552) );
  OAI211_X1 U4047 ( .C1(n4080), .C2(n3552), .A(n3646), .B(n5256), .ZN(n3554)
         );
  OAI211_X1 U4048 ( .C1(n5283), .C2(n3567), .A(n3554), .B(n3553), .ZN(n5153)
         );
  XNOR2_X1 U4049 ( .A(n3569), .B(n3567), .ZN(n5152) );
  AOI22_X1 U4050 ( .A1(n5301), .A2(REG2_REG_10__SCAN_IN), .B1(n3555), .B2(
        n5097), .ZN(n3556) );
  OAI21_X1 U4051 ( .B1(n5152), .B2(n4897), .A(n3556), .ZN(n3557) );
  AOI21_X1 U4052 ( .B1(n5153), .B2(n5258), .A(n3557), .ZN(n3558) );
  OAI21_X1 U4053 ( .B1(n3559), .B2(n4876), .A(n3558), .ZN(U3280) );
  NAND2_X1 U4054 ( .A1(n3630), .A2(n3576), .ZN(n3616) );
  NAND2_X1 U4055 ( .A1(n4566), .A2(n3629), .ZN(n3644) );
  NAND2_X1 U4056 ( .A1(n3627), .A2(n3562), .ZN(n3565) );
  INV_X1 U4057 ( .A(n4077), .ZN(n3563) );
  AND2_X1 U4058 ( .A1(n3627), .A2(n3628), .ZN(n3564) );
  AOI21_X1 U4059 ( .B1(n4077), .B2(n3565), .A(n3564), .ZN(n5160) );
  NAND2_X1 U4060 ( .A1(n3569), .A2(n3567), .ZN(n3566) );
  NAND2_X1 U4061 ( .A1(n3566), .A2(n3576), .ZN(n3570) );
  AND2_X1 U4062 ( .A1(n3629), .A2(n3567), .ZN(n3568) );
  NAND2_X1 U4063 ( .A1(n3570), .A2(n3623), .ZN(n5159) );
  INV_X1 U4064 ( .A(n5159), .ZN(n3574) );
  OAI22_X1 U4065 ( .A1(n5258), .A2(n3572), .B1(n3571), .B2(n5260), .ZN(n3573)
         );
  AOI21_X1 U4066 ( .B1(n3574), .B2(n5298), .A(n3573), .ZN(n3580) );
  NAND2_X1 U4067 ( .A1(n3646), .A2(n3643), .ZN(n3613) );
  XNOR2_X1 U4068 ( .A(n3613), .B(n4077), .ZN(n3578) );
  AOI21_X1 U4069 ( .B1(n3576), .B2(n5292), .A(n3575), .ZN(n3577) );
  OAI21_X1 U4070 ( .B1(n3578), .B2(n4860), .A(n3577), .ZN(n5161) );
  NAND2_X1 U4071 ( .A1(n5161), .A2(n5258), .ZN(n3579) );
  OAI211_X1 U4072 ( .C1(n5160), .C2(n4876), .A(n3580), .B(n3579), .ZN(U3279)
         );
  INV_X1 U4073 ( .A(n3581), .ZN(n3582) );
  NAND2_X1 U4074 ( .A1(n3583), .A2(n3582), .ZN(n3593) );
  MUX2_X1 U4075 ( .A(n4962), .B(DATAI_15_), .S(n3025), .Z(n5194) );
  OAI22_X1 U4076 ( .A1(n3668), .A2(n2965), .B1(n3711), .B2(n3859), .ZN(n3584)
         );
  NAND2_X1 U4077 ( .A1(n2966), .A2(REG2_REG_16__SCAN_IN), .ZN(n3589) );
  NAND2_X1 U4078 ( .A1(n3043), .A2(REG1_REG_16__SCAN_IN), .ZN(n3588) );
  INV_X1 U4079 ( .A(REG3_REG_16__SCAN_IN), .ZN(n4367) );
  AOI21_X1 U4080 ( .B1(n3585), .B2(n4367), .A(n3602), .ZN(n3671) );
  NAND2_X1 U4081 ( .A1(n2967), .A2(n3671), .ZN(n3587) );
  NAND2_X1 U4082 ( .A1(n3044), .A2(REG0_REG_16__SCAN_IN), .ZN(n3586) );
  MUX2_X1 U4083 ( .A(n4961), .B(DATAI_16_), .S(n3025), .Z(n3774) );
  INV_X1 U4084 ( .A(n3774), .ZN(n3664) );
  OAI22_X1 U4085 ( .A1(n4888), .A2(n2965), .B1(n3664), .B2(n3859), .ZN(n3590)
         );
  XNOR2_X1 U4086 ( .A(n3590), .B(n3879), .ZN(n3731) );
  OR2_X1 U4087 ( .A1(n4888), .A2(n3891), .ZN(n3592) );
  NAND2_X1 U4088 ( .A1(n3774), .A2(n3876), .ZN(n3591) );
  NAND2_X1 U4089 ( .A1(n3592), .A2(n3591), .ZN(n3733) );
  XNOR2_X1 U4090 ( .A(n3731), .B(n3733), .ZN(n3597) );
  NOR2_X1 U4091 ( .A1(n3598), .A2(n3597), .ZN(n3600) );
  OR2_X1 U4092 ( .A1(n3668), .A2(n3891), .ZN(n3596) );
  NAND2_X1 U4093 ( .A1(n5194), .A2(n3876), .ZN(n3595) );
  NAND2_X1 U4094 ( .A1(n5188), .A2(n5193), .ZN(n5190) );
  INV_X1 U4095 ( .A(n3732), .ZN(n3599) );
  AOI21_X1 U4096 ( .B1(n3600), .B2(n5190), .A(n3599), .ZN(n3611) );
  NOR2_X1 U4097 ( .A1(n4367), .A2(STATE_REG_SCAN_IN), .ZN(n4625) );
  INV_X1 U4098 ( .A(n4625), .ZN(n3601) );
  OAI21_X1 U4099 ( .B1(n3975), .B2(n3664), .A(n3601), .ZN(n3609) );
  NAND2_X1 U4100 ( .A1(n3602), .A2(REG3_REG_17__SCAN_IN), .ZN(n3718) );
  OAI21_X1 U4101 ( .B1(REG3_REG_17__SCAN_IN), .B2(n3602), .A(n3718), .ZN(n5221) );
  INV_X1 U4102 ( .A(n5221), .ZN(n3603) );
  NAND2_X1 U4103 ( .A1(n2967), .A2(n3603), .ZN(n3607) );
  NAND2_X1 U4104 ( .A1(n3043), .A2(REG1_REG_17__SCAN_IN), .ZN(n3606) );
  NAND2_X1 U4105 ( .A1(n2466), .A2(REG0_REG_17__SCAN_IN), .ZN(n3605) );
  NAND2_X1 U4106 ( .A1(n2966), .A2(REG2_REG_17__SCAN_IN), .ZN(n3604) );
  OAI22_X1 U4107 ( .A1(n3668), .A2(n3977), .B1(n3976), .B2(n3777), .ZN(n3608)
         );
  AOI211_X1 U4108 ( .C1(n3671), .C2(n3980), .A(n3609), .B(n3608), .ZN(n3610)
         );
  OAI21_X1 U4109 ( .B1(n3611), .B2(n5192), .A(n3610), .ZN(U3223) );
  OAI22_X1 U4110 ( .A1(n3630), .A2(n4887), .B1(n3677), .B2(n5048), .ZN(n3621)
         );
  INV_X1 U4111 ( .A(n3644), .ZN(n3612) );
  NOR2_X1 U4112 ( .A1(n3613), .A2(n3612), .ZN(n3681) );
  INV_X1 U4113 ( .A(n3681), .ZN(n3614) );
  NAND2_X1 U4114 ( .A1(n3638), .A2(n3624), .ZN(n3615) );
  INV_X1 U4115 ( .A(n3638), .ZN(n4565) );
  NAND2_X1 U4116 ( .A1(n4565), .A2(n3637), .ZN(n3679) );
  NAND2_X1 U4117 ( .A1(n3615), .A2(n3679), .ZN(n3635) );
  INV_X1 U4118 ( .A(n3635), .ZN(n4064) );
  AOI21_X1 U4119 ( .B1(n3614), .B2(n3616), .A(n4064), .ZN(n3619) );
  INV_X1 U4120 ( .A(n3679), .ZN(n3617) );
  NAND2_X1 U4121 ( .A1(n3616), .A2(n3615), .ZN(n3680) );
  NOR3_X1 U4122 ( .A1(n3681), .A2(n3617), .A3(n3680), .ZN(n3618) );
  NOR3_X1 U4123 ( .A1(n3619), .A2(n3618), .A3(n4860), .ZN(n3620) );
  AOI211_X1 U4124 ( .C1(n5292), .C2(n3624), .A(n3621), .B(n3620), .ZN(n5166)
         );
  INV_X1 U4125 ( .A(n3685), .ZN(n3622) );
  AOI211_X1 U4126 ( .C1(n3624), .C2(n3623), .A(n5273), .B(n3622), .ZN(n5168)
         );
  OAI22_X1 U4127 ( .A1(n5258), .A2(n4580), .B1(n3625), .B2(n5260), .ZN(n3626)
         );
  AOI21_X1 U4128 ( .B1(n5168), .B2(n4818), .A(n3626), .ZN(n3634) );
  NAND2_X1 U4129 ( .A1(n3628), .A2(n3627), .ZN(n3632) );
  NAND2_X1 U4130 ( .A1(n3630), .A2(n3629), .ZN(n3631) );
  NAND2_X1 U4131 ( .A1(n3632), .A2(n3631), .ZN(n3636) );
  XNOR2_X1 U4132 ( .A(n3636), .B(n3635), .ZN(n5169) );
  NAND2_X1 U4133 ( .A1(n5169), .A2(n5268), .ZN(n3633) );
  OAI211_X1 U4134 ( .C1(n5166), .C2(n5301), .A(n3634), .B(n3633), .ZN(U3278)
         );
  NAND2_X1 U4135 ( .A1(n3638), .A2(n3637), .ZN(n3639) );
  NAND2_X1 U4136 ( .A1(n3702), .A2(n3665), .ZN(n4003) );
  INV_X1 U4137 ( .A(n3702), .ZN(n4563) );
  NAND2_X1 U4138 ( .A1(n4563), .A2(n3654), .ZN(n4004) );
  NAND2_X1 U4139 ( .A1(n4003), .A2(n4004), .ZN(n3659) );
  NAND2_X1 U4140 ( .A1(n3640), .A2(n3659), .ZN(n3667) );
  OAI21_X1 U4141 ( .B1(n3640), .B2(n3659), .A(n3667), .ZN(n3641) );
  INV_X1 U4142 ( .A(n3641), .ZN(n5181) );
  NAND2_X1 U4143 ( .A1(n4564), .A2(n3687), .ZN(n3642) );
  AND2_X1 U4144 ( .A1(n3679), .A2(n3642), .ZN(n3648) );
  AND2_X1 U4145 ( .A1(n3644), .A2(n3643), .ZN(n3645) );
  NOR2_X1 U4146 ( .A1(n4564), .A2(n3687), .ZN(n3647) );
  AOI21_X1 U4147 ( .B1(n3680), .B2(n3648), .A(n3647), .ZN(n4099) );
  XNOR2_X1 U4148 ( .A(n4007), .B(n3659), .ZN(n3651) );
  OAI22_X1 U4149 ( .A1(n3668), .A2(n5048), .B1(n3677), .B2(n4887), .ZN(n3649)
         );
  AOI21_X1 U4150 ( .B1(n3665), .B2(n5292), .A(n3649), .ZN(n3650) );
  OAI21_X1 U4151 ( .B1(n3651), .B2(n4860), .A(n3650), .ZN(n5183) );
  INV_X1 U4152 ( .A(n3652), .ZN(n3684) );
  INV_X1 U4153 ( .A(n3712), .ZN(n3653) );
  OAI21_X1 U4154 ( .B1(n3684), .B2(n3654), .A(n3653), .ZN(n5180) );
  NOR2_X1 U4155 ( .A1(n5180), .A2(n4897), .ZN(n3657) );
  OAI22_X1 U4156 ( .A1(n5258), .A2(n4605), .B1(n3655), .B2(n5260), .ZN(n3656)
         );
  AOI211_X1 U4157 ( .C1(n5183), .C2(n5258), .A(n3657), .B(n3656), .ZN(n3658)
         );
  OAI21_X1 U4158 ( .B1(n5181), .B2(n4876), .A(n3658), .ZN(U3276) );
  INV_X1 U4159 ( .A(n3659), .ZN(n4078) );
  NAND2_X1 U4160 ( .A1(n3660), .A2(n4003), .ZN(n3708) );
  NAND2_X1 U4161 ( .A1(n3668), .A2(n5194), .ZN(n4006) );
  NAND2_X1 U4162 ( .A1(n4562), .A2(n3711), .ZN(n4005) );
  NAND2_X1 U4163 ( .A1(n4006), .A2(n4005), .ZN(n3707) );
  OR2_X2 U4164 ( .A1(n3708), .A2(n3707), .ZN(n3705) );
  OR2_X1 U4165 ( .A1(n4888), .A2(n3774), .ZN(n4881) );
  NAND2_X1 U4166 ( .A1(n4888), .A2(n3774), .ZN(n4136) );
  NAND3_X1 U4167 ( .A1(n3705), .A2(n2518), .A3(n4005), .ZN(n3661) );
  NAND3_X1 U4168 ( .A1(n4882), .A2(n5256), .A3(n3661), .ZN(n3663) );
  INV_X1 U4169 ( .A(n3777), .ZN(n4560) );
  AOI22_X1 U4170 ( .A1(n4866), .A2(n4562), .B1(n4560), .B2(n4839), .ZN(n3662)
         );
  OAI211_X1 U4171 ( .C1(n5283), .C2(n3664), .A(n3663), .B(n3662), .ZN(n5208)
         );
  INV_X1 U4172 ( .A(n5208), .ZN(n3676) );
  NAND2_X1 U4173 ( .A1(n3667), .A2(n3666), .ZN(n3701) );
  NAND2_X1 U4174 ( .A1(n4562), .A2(n5194), .ZN(n3669) );
  XNOR2_X1 U4175 ( .A(n3775), .B(n4068), .ZN(n5210) );
  NAND2_X1 U4176 ( .A1(n5210), .A2(n5268), .ZN(n3675) );
  INV_X1 U4177 ( .A(n4877), .ZN(n3670) );
  AOI211_X1 U4178 ( .C1(n3774), .C2(n3710), .A(n5273), .B(n3670), .ZN(n5209)
         );
  INV_X1 U4179 ( .A(n3671), .ZN(n3672) );
  OAI22_X1 U4180 ( .A1(n5258), .A2(n4627), .B1(n3672), .B2(n5260), .ZN(n3673)
         );
  AOI21_X1 U4181 ( .B1(n5209), .B2(n4818), .A(n3673), .ZN(n3674) );
  OAI211_X1 U4182 ( .C1(n5301), .C2(n3676), .A(n3675), .B(n3674), .ZN(U3274)
         );
  XNOR2_X1 U4183 ( .A(n3677), .B(n3687), .ZN(n4069) );
  XNOR2_X1 U4184 ( .A(n3678), .B(n4069), .ZN(n5173) );
  OAI21_X1 U4185 ( .B1(n3681), .B2(n3680), .A(n3679), .ZN(n3682) );
  XNOR2_X1 U4186 ( .A(n3682), .B(n4069), .ZN(n3683) );
  NOR2_X1 U4187 ( .A1(n3683), .A2(n4860), .ZN(n3691) );
  AOI211_X1 U4188 ( .C1(n3686), .C2(n3685), .A(n5273), .B(n3684), .ZN(n3689)
         );
  NOR2_X1 U4189 ( .A1(n3687), .A2(n5283), .ZN(n3692) );
  NOR4_X1 U4190 ( .A1(n3691), .A2(n3689), .A3(n3692), .A4(n3688), .ZN(n5174)
         );
  OAI21_X1 U4191 ( .B1(n5173), .B2(n3690), .A(n5174), .ZN(n3696) );
  INV_X1 U4192 ( .A(n3691), .ZN(n3694) );
  INV_X1 U4193 ( .A(n3692), .ZN(n3693) );
  NAND3_X1 U4194 ( .A1(n3694), .A2(n4959), .A3(n3693), .ZN(n3695) );
  NAND3_X1 U4195 ( .A1(n3696), .A2(n5258), .A3(n3695), .ZN(n3699) );
  AOI22_X1 U4196 ( .A1(n5301), .A2(REG2_REG_13__SCAN_IN), .B1(n5097), .B2(
        n3697), .ZN(n3698) );
  OAI211_X1 U4197 ( .C1(n5173), .C2(n3700), .A(n3699), .B(n3698), .ZN(U3277)
         );
  INV_X1 U4198 ( .A(n3707), .ZN(n4065) );
  XNOR2_X1 U4199 ( .A(n3701), .B(n4065), .ZN(n5203) );
  OR2_X1 U4200 ( .A1(n4888), .A2(n5048), .ZN(n3704) );
  OR2_X1 U4201 ( .A1(n3702), .A2(n4887), .ZN(n3703) );
  NAND2_X1 U4202 ( .A1(n3704), .A2(n3703), .ZN(n5187) );
  INV_X1 U4203 ( .A(n3705), .ZN(n3706) );
  AOI211_X1 U4204 ( .C1(n3708), .C2(n3707), .A(n4860), .B(n3706), .ZN(n3709)
         );
  AOI211_X1 U4205 ( .C1(n5292), .C2(n5194), .A(n5187), .B(n3709), .ZN(n5201)
         );
  INV_X1 U4206 ( .A(n5201), .ZN(n3716) );
  OAI211_X1 U4207 ( .C1(n3712), .C2(n3711), .A(n5303), .B(n3710), .ZN(n5200)
         );
  INV_X1 U4208 ( .A(n4818), .ZN(n4872) );
  AOI22_X1 U4209 ( .A1(n5301), .A2(REG2_REG_15__SCAN_IN), .B1(n5097), .B2(
        n3713), .ZN(n3714) );
  OAI21_X1 U4210 ( .B1(n5200), .B2(n4872), .A(n3714), .ZN(n3715) );
  AOI21_X1 U4211 ( .B1(n3716), .B2(n5258), .A(n3715), .ZN(n3717) );
  OAI21_X1 U4212 ( .B1(n5203), .B2(n4876), .A(n3717), .ZN(U3275) );
  INV_X1 U4213 ( .A(REG3_REG_19__SCAN_IN), .ZN(n4206) );
  XNOR2_X1 U4214 ( .A(n4206), .B(n3757), .ZN(n5261) );
  INV_X1 U4215 ( .A(n5261), .ZN(n3767) );
  NAND2_X1 U4216 ( .A1(n2967), .A2(n3767), .ZN(n3722) );
  NAND2_X1 U4217 ( .A1(n3043), .A2(REG1_REG_19__SCAN_IN), .ZN(n3721) );
  NAND2_X1 U4218 ( .A1(n2466), .A2(REG0_REG_19__SCAN_IN), .ZN(n3720) );
  NAND2_X1 U4219 ( .A1(n2966), .A2(REG2_REG_19__SCAN_IN), .ZN(n3719) );
  NAND4_X1 U4220 ( .A1(n3722), .A2(n3721), .A3(n3720), .A4(n3719), .ZN(n4865)
         );
  NAND2_X1 U4221 ( .A1(n4865), .A2(n3844), .ZN(n3725) );
  INV_X1 U4222 ( .A(DATAI_19_), .ZN(n3723) );
  MUX2_X1 U4223 ( .A(n5006), .B(n3723), .S(n3025), .Z(n5266) );
  OR2_X1 U4224 ( .A1(n5266), .A2(n3859), .ZN(n3724) );
  NAND2_X1 U4225 ( .A1(n3725), .A2(n3724), .ZN(n3726) );
  XNOR2_X1 U4226 ( .A(n3726), .B(n3892), .ZN(n3730) );
  NAND2_X1 U4227 ( .A1(n4865), .A2(n3882), .ZN(n3728) );
  OR2_X1 U4228 ( .A1(n5266), .A2(n2965), .ZN(n3727) );
  NAND2_X1 U4229 ( .A1(n3728), .A2(n3727), .ZN(n3729) );
  NOR2_X1 U4230 ( .A1(n3730), .A2(n3729), .ZN(n3810) );
  AOI21_X1 U4231 ( .B1(n3730), .B2(n3729), .A(n3810), .ZN(n3753) );
  OR2_X1 U4232 ( .A1(n3777), .A2(n3891), .ZN(n3735) );
  MUX2_X1 U4233 ( .A(n4960), .B(DATAI_17_), .S(n3025), .Z(n5217) );
  NAND2_X1 U4234 ( .A1(n5217), .A2(n3876), .ZN(n3734) );
  NAND2_X1 U4235 ( .A1(n3735), .A2(n3734), .ZN(n3738) );
  INV_X1 U4236 ( .A(n5217), .ZN(n4885) );
  OAI22_X1 U4237 ( .A1(n3777), .A2(n2965), .B1(n4885), .B2(n3859), .ZN(n3736)
         );
  XNOR2_X1 U4238 ( .A(n3736), .B(n3892), .ZN(n3737) );
  XOR2_X1 U4239 ( .A(n3738), .B(n3737), .Z(n5215) );
  INV_X1 U4240 ( .A(n3737), .ZN(n3740) );
  INV_X1 U4241 ( .A(n3738), .ZN(n3739) );
  NAND2_X1 U4242 ( .A1(n2966), .A2(REG2_REG_18__SCAN_IN), .ZN(n3746) );
  NAND2_X1 U4243 ( .A1(n3043), .A2(REG1_REG_18__SCAN_IN), .ZN(n3745) );
  OAI21_X1 U4244 ( .B1(REG3_REG_18__SCAN_IN), .B2(n3741), .A(n3757), .ZN(n5243) );
  INV_X1 U4245 ( .A(n5243), .ZN(n3742) );
  NAND2_X1 U4246 ( .A1(n2967), .A2(n3742), .ZN(n3744) );
  NAND2_X1 U4247 ( .A1(n3044), .A2(REG0_REG_18__SCAN_IN), .ZN(n3743) );
  MUX2_X1 U4248 ( .A(n5001), .B(DATAI_18_), .S(n3025), .Z(n5238) );
  OAI22_X1 U4249 ( .A1(n4886), .A2(n2965), .B1(n3778), .B2(n3859), .ZN(n3747)
         );
  XNOR2_X1 U4250 ( .A(n3747), .B(n3879), .ZN(n3750) );
  OR2_X1 U4251 ( .A1(n4886), .A2(n3891), .ZN(n3749) );
  NAND2_X1 U4252 ( .A1(n5238), .A2(n3876), .ZN(n3748) );
  AND2_X1 U4253 ( .A1(n3749), .A2(n3748), .ZN(n3751) );
  NOR2_X1 U4254 ( .A1(n3750), .A2(n3751), .ZN(n5232) );
  NAND2_X1 U4255 ( .A1(n3751), .A2(n3750), .ZN(n5233) );
  NAND2_X1 U4256 ( .A1(n3752), .A2(n3753), .ZN(n3812) );
  OAI21_X1 U4257 ( .B1(n3753), .B2(n3752), .A(n3812), .ZN(n3754) );
  INV_X1 U4258 ( .A(n3754), .ZN(n3769) );
  NAND2_X1 U4259 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n5004) );
  OR2_X1 U4260 ( .A1(n4886), .A2(n4887), .ZN(n3764) );
  NAND2_X1 U4261 ( .A1(n3043), .A2(REG1_REG_20__SCAN_IN), .ZN(n3762) );
  NAND2_X1 U4262 ( .A1(n2966), .A2(REG2_REG_20__SCAN_IN), .ZN(n3761) );
  INV_X1 U4263 ( .A(n3757), .ZN(n3755) );
  AOI21_X1 U4264 ( .B1(n3755), .B2(REG3_REG_19__SCAN_IN), .A(
        REG3_REG_20__SCAN_IN), .ZN(n3758) );
  NAND2_X1 U4265 ( .A1(REG3_REG_19__SCAN_IN), .A2(REG3_REG_20__SCAN_IN), .ZN(
        n3756) );
  NOR2_X1 U4266 ( .A1(n3758), .A2(n3819), .ZN(n4870) );
  NAND2_X1 U4267 ( .A1(n2967), .A2(n4870), .ZN(n3760) );
  NAND2_X1 U4268 ( .A1(n3044), .A2(REG0_REG_20__SCAN_IN), .ZN(n3759) );
  NAND2_X1 U4269 ( .A1(n4838), .A2(n4839), .ZN(n3763) );
  NAND2_X1 U4270 ( .A1(n3764), .A2(n3763), .ZN(n5254) );
  NAND2_X1 U4271 ( .A1(n5231), .A2(n5254), .ZN(n3765) );
  OAI211_X1 U4272 ( .C1(n3975), .C2(n5266), .A(n5004), .B(n3765), .ZN(n3766)
         );
  AOI21_X1 U4273 ( .B1(n3980), .B2(n3767), .A(n3766), .ZN(n3768) );
  OAI21_X1 U4274 ( .B1(n3769), .B2(n5192), .A(n3768), .ZN(U3216) );
  NAND2_X1 U4275 ( .A1(n4560), .A2(n4885), .ZN(n3776) );
  AND2_X1 U4276 ( .A1(n4881), .A2(n3776), .ZN(n4008) );
  NAND2_X1 U4277 ( .A1(n3777), .A2(n5217), .ZN(n4014) );
  INV_X1 U4278 ( .A(n4014), .ZN(n3770) );
  AOI21_X1 U4279 ( .B1(n4882), .B2(n4008), .A(n3770), .ZN(n3771) );
  NAND2_X1 U4280 ( .A1(n4886), .A2(n5238), .ZN(n4013) );
  NAND2_X1 U4281 ( .A1(n4648), .A2(n3778), .ZN(n5251) );
  NAND2_X1 U4282 ( .A1(n3771), .A2(n4649), .ZN(n5252) );
  OAI211_X1 U4283 ( .C1(n3771), .C2(n4649), .A(n5252), .B(n5256), .ZN(n3773)
         );
  OAI22_X1 U4284 ( .A1(n4651), .A2(n5048), .B1(n3777), .B2(n4887), .ZN(n5230)
         );
  INV_X1 U4285 ( .A(n5230), .ZN(n3772) );
  OAI211_X1 U4286 ( .C1(n5283), .C2(n3778), .A(n3773), .B(n3772), .ZN(n5245)
         );
  INV_X1 U4287 ( .A(n5245), .ZN(n3783) );
  INV_X1 U4288 ( .A(n4888), .ZN(n4561) );
  NAND2_X1 U4289 ( .A1(n4014), .A2(n3776), .ZN(n4883) );
  XNOR2_X1 U4290 ( .A(n4650), .B(n4649), .ZN(n5247) );
  NAND2_X1 U4291 ( .A1(n5247), .A2(n5268), .ZN(n3782) );
  INV_X1 U4292 ( .A(n3779), .ZN(n4879) );
  AOI211_X1 U4293 ( .C1(n5238), .C2(n4879), .A(n5273), .B(n4695), .ZN(n5246)
         );
  OAI22_X1 U4294 ( .A1(n5258), .A2(n2854), .B1(n5243), .B2(n5260), .ZN(n3780)
         );
  AOI21_X1 U4295 ( .B1(n5246), .B2(n4818), .A(n3780), .ZN(n3781) );
  OAI211_X1 U4296 ( .C1(n5301), .C2(n3783), .A(n3782), .B(n3781), .ZN(U3272)
         );
  NAND2_X1 U4297 ( .A1(n2966), .A2(REG2_REG_26__SCAN_IN), .ZN(n3789) );
  NAND2_X1 U4298 ( .A1(n3043), .A2(REG1_REG_26__SCAN_IN), .ZN(n3788) );
  NAND2_X1 U4299 ( .A1(n3819), .A2(REG3_REG_21__SCAN_IN), .ZN(n3821) );
  INV_X1 U4300 ( .A(REG3_REG_22__SCAN_IN), .ZN(n3974) );
  INV_X1 U4301 ( .A(REG3_REG_23__SCAN_IN), .ZN(n4381) );
  INV_X1 U4302 ( .A(REG3_REG_24__SCAN_IN), .ZN(n3956) );
  NOR2_X1 U4303 ( .A1(n3795), .A2(REG3_REG_26__SCAN_IN), .ZN(n3784) );
  OR2_X1 U4304 ( .A1(n3870), .A2(n3784), .ZN(n4743) );
  INV_X1 U4305 ( .A(n4743), .ZN(n3785) );
  NAND2_X1 U4306 ( .A1(n2967), .A2(n3785), .ZN(n3787) );
  NAND2_X1 U4307 ( .A1(n3044), .A2(REG0_REG_26__SCAN_IN), .ZN(n3786) );
  NAND4_X1 U4308 ( .A1(n3789), .A2(n3788), .A3(n3787), .A4(n3786), .ZN(n4769)
         );
  NAND2_X1 U4309 ( .A1(n4769), .A2(n3800), .ZN(n3791) );
  NAND2_X1 U4310 ( .A1(n3025), .A2(DATAI_26_), .ZN(n4753) );
  OR2_X1 U4311 ( .A1(n4753), .A2(n3859), .ZN(n3790) );
  NAND2_X1 U4312 ( .A1(n3791), .A2(n3790), .ZN(n3792) );
  XNOR2_X1 U4313 ( .A(n3792), .B(n3879), .ZN(n3984) );
  INV_X1 U4314 ( .A(n3984), .ZN(n3869) );
  NOR2_X1 U4315 ( .A1(n4753), .A2(n2965), .ZN(n3793) );
  AOI21_X1 U4316 ( .B1(n4769), .B2(n3882), .A(n3793), .ZN(n3983) );
  INV_X1 U4317 ( .A(n3983), .ZN(n3868) );
  NAND2_X1 U4318 ( .A1(n2966), .A2(REG2_REG_25__SCAN_IN), .ZN(n3799) );
  NAND2_X1 U4319 ( .A1(n3043), .A2(REG1_REG_25__SCAN_IN), .ZN(n3798) );
  NOR2_X1 U4320 ( .A1(n3854), .A2(REG3_REG_25__SCAN_IN), .ZN(n3794) );
  OR2_X1 U4321 ( .A1(n3795), .A2(n3794), .ZN(n4761) );
  INV_X1 U4322 ( .A(n4761), .ZN(n3946) );
  NAND2_X1 U4323 ( .A1(n2967), .A2(n3946), .ZN(n3797) );
  NAND2_X1 U4324 ( .A1(n3044), .A2(REG0_REG_25__SCAN_IN), .ZN(n3796) );
  OR2_X1 U4325 ( .A1(n4781), .A2(n3891), .ZN(n3802) );
  NAND2_X1 U4326 ( .A1(n4760), .A2(n3800), .ZN(n3801) );
  NAND2_X1 U4327 ( .A1(n3802), .A2(n3801), .ZN(n3866) );
  INV_X1 U4328 ( .A(n4760), .ZN(n4772) );
  OAI22_X1 U4329 ( .A1(n4781), .A2(n2965), .B1(n4772), .B2(n3859), .ZN(n3803)
         );
  XNOR2_X1 U4330 ( .A(n3803), .B(n3892), .ZN(n3865) );
  NAND2_X1 U4331 ( .A1(n2966), .A2(REG2_REG_22__SCAN_IN), .ZN(n3808) );
  NAND2_X1 U4332 ( .A1(n3043), .A2(REG1_REG_22__SCAN_IN), .ZN(n3807) );
  NAND2_X1 U4333 ( .A1(n3821), .A2(n3974), .ZN(n3804) );
  AND2_X1 U4334 ( .A1(n3838), .A2(n3804), .ZN(n4814) );
  NAND2_X1 U4335 ( .A1(n2967), .A2(n4814), .ZN(n3806) );
  NAND2_X1 U4336 ( .A1(n2466), .A2(REG0_REG_22__SCAN_IN), .ZN(n3805) );
  NAND4_X1 U4337 ( .A1(n3808), .A2(n3807), .A3(n3806), .A4(n3805), .ZN(n4840)
         );
  OAI22_X1 U4338 ( .A1(n4657), .A2(n3891), .B1(n4828), .B2(n2965), .ZN(n3834)
         );
  INV_X1 U4339 ( .A(n3834), .ZN(n3837) );
  OAI22_X1 U4340 ( .A1(n4657), .A2(n2965), .B1(n4828), .B2(n3859), .ZN(n3809)
         );
  XNOR2_X1 U4341 ( .A(n3809), .B(n3892), .ZN(n3835) );
  INV_X1 U4342 ( .A(n3835), .ZN(n3836) );
  INV_X1 U4343 ( .A(n3810), .ZN(n3811) );
  NAND2_X1 U4344 ( .A1(n3812), .A2(n3811), .ZN(n3965) );
  NAND2_X1 U4345 ( .A1(n4838), .A2(n3844), .ZN(n3814) );
  OR2_X1 U4346 ( .A1(n4868), .A2(n3859), .ZN(n3813) );
  NAND2_X1 U4347 ( .A1(n3814), .A2(n3813), .ZN(n3815) );
  XNOR2_X1 U4348 ( .A(n3815), .B(n3879), .ZN(n3818) );
  NOR2_X1 U4349 ( .A1(n4868), .A2(n2965), .ZN(n3816) );
  AOI21_X1 U4350 ( .B1(n4838), .B2(n3882), .A(n3816), .ZN(n3817) );
  OR2_X1 U4351 ( .A1(n3818), .A2(n3817), .ZN(n3962) );
  AND2_X1 U4352 ( .A1(n3818), .A2(n3817), .ZN(n3961) );
  NAND2_X1 U4353 ( .A1(n2966), .A2(REG2_REG_21__SCAN_IN), .ZN(n3825) );
  NAND2_X1 U4354 ( .A1(n3043), .A2(REG1_REG_21__SCAN_IN), .ZN(n3824) );
  OR2_X1 U4355 ( .A1(n3819), .A2(REG3_REG_21__SCAN_IN), .ZN(n3820) );
  AND2_X1 U4356 ( .A1(n3821), .A2(n3820), .ZN(n4849) );
  NAND2_X1 U4357 ( .A1(n2967), .A2(n4849), .ZN(n3823) );
  NAND2_X1 U4358 ( .A1(n2466), .A2(REG0_REG_21__SCAN_IN), .ZN(n3822) );
  NAND2_X1 U4359 ( .A1(n4825), .A2(n3876), .ZN(n3827) );
  OR2_X1 U4360 ( .A1(n4847), .A2(n3859), .ZN(n3826) );
  NAND2_X1 U4361 ( .A1(n3827), .A2(n3826), .ZN(n3828) );
  XNOR2_X1 U4362 ( .A(n3828), .B(n3879), .ZN(n3830) );
  NOR2_X1 U4363 ( .A1(n4847), .A2(n2965), .ZN(n3829) );
  AOI21_X1 U4364 ( .B1(n4825), .B2(n3882), .A(n3829), .ZN(n3831) );
  NAND2_X1 U4365 ( .A1(n3830), .A2(n3831), .ZN(n3929) );
  NAND2_X1 U4366 ( .A1(n3932), .A2(n3929), .ZN(n3934) );
  INV_X1 U4367 ( .A(n3830), .ZN(n3833) );
  INV_X1 U4368 ( .A(n3831), .ZN(n3832) );
  NAND2_X1 U4369 ( .A1(n3833), .A2(n3832), .ZN(n3931) );
  NAND2_X1 U4370 ( .A1(n3934), .A2(n3931), .ZN(n3972) );
  XNOR2_X1 U4371 ( .A(n3835), .B(n3834), .ZN(n3973) );
  NAND2_X1 U4372 ( .A1(n2966), .A2(REG2_REG_23__SCAN_IN), .ZN(n3843) );
  NAND2_X1 U4373 ( .A1(n3043), .A2(REG1_REG_23__SCAN_IN), .ZN(n3842) );
  NAND2_X1 U4374 ( .A1(n3838), .A2(n4381), .ZN(n3839) );
  AND2_X1 U4375 ( .A1(n3852), .A2(n3839), .ZN(n4805) );
  NAND2_X1 U4376 ( .A1(n2967), .A2(n4805), .ZN(n3841) );
  NAND2_X1 U4377 ( .A1(n3044), .A2(REG0_REG_23__SCAN_IN), .ZN(n3840) );
  NAND4_X1 U4378 ( .A1(n3843), .A2(n3842), .A3(n3841), .A4(n3840), .ZN(n4824)
         );
  NAND2_X1 U4379 ( .A1(n4824), .A2(n3844), .ZN(n3846) );
  OR2_X1 U4380 ( .A1(n4802), .A2(n3859), .ZN(n3845) );
  NAND2_X1 U4381 ( .A1(n3846), .A2(n3845), .ZN(n3847) );
  XNOR2_X1 U4382 ( .A(n3847), .B(n3892), .ZN(n3850) );
  NOR2_X1 U4383 ( .A1(n4802), .A2(n2965), .ZN(n3848) );
  AOI21_X1 U4384 ( .B1(n4824), .B2(n3882), .A(n3848), .ZN(n3849) );
  XNOR2_X1 U4385 ( .A(n3850), .B(n3849), .ZN(n3914) );
  INV_X1 U4386 ( .A(n3849), .ZN(n3851) );
  NAND2_X1 U4387 ( .A1(n2966), .A2(REG2_REG_24__SCAN_IN), .ZN(n3858) );
  NAND2_X1 U4388 ( .A1(n3043), .A2(REG1_REG_24__SCAN_IN), .ZN(n3857) );
  AND2_X1 U4389 ( .A1(n3852), .A2(n3956), .ZN(n3853) );
  NOR2_X1 U4390 ( .A1(n3854), .A2(n3853), .ZN(n4787) );
  NAND2_X1 U4391 ( .A1(n2967), .A2(n4787), .ZN(n3856) );
  NAND2_X1 U4392 ( .A1(n2466), .A2(REG0_REG_24__SCAN_IN), .ZN(n3855) );
  NAND4_X1 U4393 ( .A1(n3858), .A2(n3857), .A3(n3856), .A4(n3855), .ZN(n4799)
         );
  INV_X1 U4394 ( .A(n4799), .ZN(n4662) );
  OAI22_X1 U4395 ( .A1(n4662), .A2(n2965), .B1(n4661), .B2(n3859), .ZN(n3860)
         );
  XOR2_X1 U4396 ( .A(n3892), .B(n3860), .Z(n3863) );
  NAND2_X1 U4397 ( .A1(n4799), .A2(n3882), .ZN(n3862) );
  OR2_X1 U4398 ( .A1(n4661), .A2(n2965), .ZN(n3861) );
  NAND2_X1 U4399 ( .A1(n3862), .A2(n3861), .ZN(n3954) );
  XOR2_X1 U4400 ( .A(n3866), .B(n3865), .Z(n3942) );
  OAI21_X1 U4401 ( .B1(n3866), .B2(n3865), .A(n3940), .ZN(n3986) );
  AOI21_X1 U4402 ( .B1(n3984), .B2(n3983), .A(n3986), .ZN(n3867) );
  NAND2_X1 U4403 ( .A1(n2966), .A2(REG2_REG_27__SCAN_IN), .ZN(n3875) );
  NAND2_X1 U4404 ( .A1(n3043), .A2(REG1_REG_27__SCAN_IN), .ZN(n3874) );
  NAND2_X1 U4405 ( .A1(n3870), .A2(REG3_REG_27__SCAN_IN), .ZN(n3885) );
  OR2_X1 U4406 ( .A1(n3870), .A2(REG3_REG_27__SCAN_IN), .ZN(n3871) );
  NAND2_X1 U4407 ( .A1(n2967), .A2(n4733), .ZN(n3873) );
  NAND2_X1 U4408 ( .A1(n2466), .A2(REG0_REG_27__SCAN_IN), .ZN(n3872) );
  NAND4_X1 U4409 ( .A1(n3875), .A2(n3874), .A3(n3873), .A4(n3872), .ZN(n4669)
         );
  NAND2_X1 U4410 ( .A1(n4669), .A2(n3876), .ZN(n3878) );
  NAND2_X1 U4411 ( .A1(n4000), .A2(DATAI_27_), .ZN(n4730) );
  OR2_X1 U4412 ( .A1(n4730), .A2(n3859), .ZN(n3877) );
  NAND2_X1 U4413 ( .A1(n3878), .A2(n3877), .ZN(n3880) );
  XNOR2_X1 U4414 ( .A(n3880), .B(n3879), .ZN(n3883) );
  NOR2_X1 U4415 ( .A1(n4730), .A2(n2965), .ZN(n3881) );
  AOI21_X1 U4416 ( .B1(n4669), .B2(n3882), .A(n3881), .ZN(n3884) );
  XNOR2_X1 U4417 ( .A(n3883), .B(n3884), .ZN(n3908) );
  OAI22_X1 U4418 ( .A1(n3909), .A2(n3908), .B1(n3884), .B2(n3883), .ZN(n3897)
         );
  NAND2_X1 U4419 ( .A1(n3043), .A2(REG1_REG_28__SCAN_IN), .ZN(n3890) );
  NAND2_X1 U4420 ( .A1(n2466), .A2(REG0_REG_28__SCAN_IN), .ZN(n3889) );
  INV_X1 U4421 ( .A(REG3_REG_28__SCAN_IN), .ZN(n4440) );
  OR2_X1 U4422 ( .A1(n3885), .A2(n4440), .ZN(n3898) );
  NAND2_X1 U4423 ( .A1(n3885), .A2(n4440), .ZN(n3886) );
  NAND2_X1 U4424 ( .A1(n2967), .A2(n4716), .ZN(n3888) );
  NAND2_X1 U4425 ( .A1(n2966), .A2(REG2_REG_28__SCAN_IN), .ZN(n3887) );
  NAND4_X1 U4426 ( .A1(n3890), .A2(n3889), .A3(n3888), .A4(n3887), .ZN(n4159)
         );
  INV_X1 U4427 ( .A(n4159), .ZN(n4722) );
  NAND2_X1 U4428 ( .A1(n3025), .A2(DATAI_28_), .ZN(n4713) );
  OAI22_X1 U4429 ( .A1(n4722), .A2(n3891), .B1(n4713), .B2(n2965), .ZN(n3895)
         );
  OAI22_X1 U4430 ( .A1(n4722), .A2(n2965), .B1(n4713), .B2(n3859), .ZN(n3893)
         );
  XNOR2_X1 U4431 ( .A(n3893), .B(n3892), .ZN(n3894) );
  XOR2_X1 U4432 ( .A(n3895), .B(n3894), .Z(n3896) );
  XNOR2_X1 U4433 ( .A(n3897), .B(n3896), .ZN(n3906) );
  OAI22_X1 U4434 ( .A1(n3975), .A2(n4713), .B1(STATE_REG_SCAN_IN), .B2(n4440), 
        .ZN(n3904) );
  INV_X1 U4435 ( .A(n4669), .ZN(n4707) );
  NAND2_X1 U4436 ( .A1(n3043), .A2(REG1_REG_29__SCAN_IN), .ZN(n3902) );
  NAND2_X1 U4437 ( .A1(n3044), .A2(REG0_REG_29__SCAN_IN), .ZN(n3901) );
  INV_X1 U4438 ( .A(n3898), .ZN(n4672) );
  NAND2_X1 U4439 ( .A1(n2967), .A2(n4672), .ZN(n3900) );
  NAND2_X1 U4440 ( .A1(n2966), .A2(REG2_REG_29__SCAN_IN), .ZN(n3899) );
  NAND4_X1 U4441 ( .A1(n3902), .A2(n3901), .A3(n3900), .A4(n3899), .ZN(n4712)
         );
  INV_X1 U4442 ( .A(n4712), .ZN(n4030) );
  OAI22_X1 U4443 ( .A1(n4707), .A2(n3977), .B1(n3976), .B2(n4030), .ZN(n3903)
         );
  AOI211_X1 U4444 ( .C1(n4716), .C2(n3980), .A(n3904), .B(n3903), .ZN(n3905)
         );
  OAI21_X1 U4445 ( .B1(n3906), .B2(n5192), .A(n3905), .ZN(U3217) );
  INV_X1 U4446 ( .A(DATAI_28_), .ZN(n4402) );
  MUX2_X1 U4447 ( .A(n4402), .B(n2855), .S(STATE_REG_SCAN_IN), .Z(n3907) );
  INV_X1 U4448 ( .A(n3907), .ZN(U3324) );
  XNOR2_X1 U4449 ( .A(n3909), .B(n3908), .ZN(n3913) );
  INV_X1 U4450 ( .A(REG3_REG_27__SCAN_IN), .ZN(n4380) );
  OAI22_X1 U4451 ( .A1(n3975), .A2(n4730), .B1(STATE_REG_SCAN_IN), .B2(n4380), 
        .ZN(n3911) );
  INV_X1 U4452 ( .A(n4769), .ZN(n4028) );
  OAI22_X1 U4453 ( .A1(n4028), .A2(n3977), .B1(n3976), .B2(n4722), .ZN(n3910)
         );
  AOI211_X1 U4454 ( .C1(n4733), .C2(n3980), .A(n3911), .B(n3910), .ZN(n3912)
         );
  OAI21_X1 U4455 ( .B1(n3913), .B2(n5192), .A(n3912), .ZN(U3211) );
  XNOR2_X1 U4456 ( .A(n3915), .B(n3914), .ZN(n3919) );
  OAI22_X1 U4457 ( .A1(n3975), .A2(n4802), .B1(STATE_REG_SCAN_IN), .B2(n4381), 
        .ZN(n3917) );
  OAI22_X1 U4458 ( .A1(n4662), .A2(n3976), .B1(n3977), .B2(n4657), .ZN(n3916)
         );
  AOI211_X1 U4459 ( .C1(n4805), .C2(n3980), .A(n3917), .B(n3916), .ZN(n3918)
         );
  OAI21_X1 U4460 ( .B1(n3919), .B2(n5192), .A(n3918), .ZN(U3213) );
  OAI21_X1 U4461 ( .B1(n3921), .B2(n3920), .A(n3155), .ZN(n3922) );
  NAND2_X1 U4462 ( .A1(n3922), .A2(n5239), .ZN(n3928) );
  OR2_X1 U4463 ( .A1(n3923), .A2(n5048), .ZN(n3925) );
  NAND2_X1 U4464 ( .A1(n3087), .A2(n4866), .ZN(n3924) );
  NAND2_X1 U4465 ( .A1(n3925), .A2(n3924), .ZN(n5081) );
  AOI22_X1 U4466 ( .A1(n5237), .A2(n5090), .B1(n5231), .B2(n5081), .ZN(n3927)
         );
  MUX2_X1 U4467 ( .A(n5244), .B(STATE_REG_SCAN_IN), .S(REG3_REG_3__SCAN_IN), 
        .Z(n3926) );
  NAND3_X1 U4468 ( .A1(n3928), .A2(n3927), .A3(n3926), .ZN(U3215) );
  AOI21_X1 U4469 ( .B1(n3931), .B2(n3929), .A(n3932), .ZN(n3930) );
  INV_X1 U4470 ( .A(n3930), .ZN(n3935) );
  INV_X1 U4471 ( .A(n3931), .ZN(n3933) );
  AOI22_X1 U4472 ( .A1(n3935), .A2(n3934), .B1(n3933), .B2(n3932), .ZN(n3939)
         );
  INV_X1 U4473 ( .A(REG3_REG_21__SCAN_IN), .ZN(n4221) );
  OAI22_X1 U4474 ( .A1(n3975), .A2(n4847), .B1(STATE_REG_SCAN_IN), .B2(n4221), 
        .ZN(n3937) );
  OAI22_X1 U4475 ( .A1(n4653), .A2(n3977), .B1(n3976), .B2(n4657), .ZN(n3936)
         );
  AOI211_X1 U4476 ( .C1(n4849), .C2(n3980), .A(n3937), .B(n3936), .ZN(n3938)
         );
  OAI21_X1 U4477 ( .B1(n3939), .B2(n5192), .A(n3938), .ZN(U3220) );
  OAI21_X1 U4478 ( .B1(n3942), .B2(n3941), .A(n3940), .ZN(n3943) );
  INV_X1 U4479 ( .A(n3943), .ZN(n3948) );
  INV_X1 U4480 ( .A(REG3_REG_25__SCAN_IN), .ZN(n4368) );
  OAI22_X1 U4481 ( .A1(n3975), .A2(n4772), .B1(STATE_REG_SCAN_IN), .B2(n4368), 
        .ZN(n3945) );
  OAI22_X1 U4482 ( .A1(n4662), .A2(n3977), .B1(n3976), .B2(n4028), .ZN(n3944)
         );
  AOI211_X1 U4483 ( .C1(n3946), .C2(n3980), .A(n3945), .B(n3944), .ZN(n3947)
         );
  OAI21_X1 U4484 ( .B1(n3948), .B2(n5192), .A(n3947), .ZN(U3222) );
  INV_X1 U4485 ( .A(n3955), .ZN(n3950) );
  AOI21_X1 U4486 ( .B1(n3950), .B2(n3949), .A(n3954), .ZN(n3952) );
  NOR2_X1 U4487 ( .A1(n3952), .A2(n3951), .ZN(n3953) );
  AOI21_X1 U4488 ( .B1(n3955), .B2(n3954), .A(n3953), .ZN(n3960) );
  OAI22_X1 U4489 ( .A1(n3975), .A2(n4661), .B1(STATE_REG_SCAN_IN), .B2(n3956), 
        .ZN(n3958) );
  INV_X1 U4490 ( .A(n4824), .ZN(n4049) );
  OAI22_X1 U4491 ( .A1(n4049), .A2(n3977), .B1(n3976), .B2(n4781), .ZN(n3957)
         );
  AOI211_X1 U4492 ( .C1(n4787), .C2(n3980), .A(n3958), .B(n3957), .ZN(n3959)
         );
  OAI21_X1 U4493 ( .B1(n3960), .B2(n5192), .A(n3959), .ZN(U3226) );
  INV_X1 U4494 ( .A(n3961), .ZN(n3963) );
  NAND2_X1 U4495 ( .A1(n3963), .A2(n3962), .ZN(n3964) );
  XNOR2_X1 U4496 ( .A(n3965), .B(n3964), .ZN(n3970) );
  INV_X1 U4497 ( .A(REG3_REG_20__SCAN_IN), .ZN(n3966) );
  OAI22_X1 U4498 ( .A1(n3975), .A2(n4868), .B1(STATE_REG_SCAN_IN), .B2(n3966), 
        .ZN(n3968) );
  OAI22_X1 U4499 ( .A1(n4651), .A2(n3977), .B1(n3976), .B2(n4855), .ZN(n3967)
         );
  AOI211_X1 U4500 ( .C1(n4870), .C2(n3980), .A(n3968), .B(n3967), .ZN(n3969)
         );
  OAI21_X1 U4501 ( .B1(n3970), .B2(n5192), .A(n3969), .ZN(U3230) );
  AOI21_X1 U4502 ( .B1(n3973), .B2(n3972), .A(n3971), .ZN(n3982) );
  OAI22_X1 U4503 ( .A1(n3975), .A2(n4828), .B1(STATE_REG_SCAN_IN), .B2(n3974), 
        .ZN(n3979) );
  OAI22_X1 U4504 ( .A1(n4855), .A2(n3977), .B1(n3976), .B2(n4049), .ZN(n3978)
         );
  AOI211_X1 U4505 ( .C1(n4814), .C2(n3980), .A(n3979), .B(n3978), .ZN(n3981)
         );
  OAI21_X1 U4506 ( .B1(n3982), .B2(n5192), .A(n3981), .ZN(U3232) );
  XNOR2_X1 U4507 ( .A(n3984), .B(n3983), .ZN(n3985) );
  XNOR2_X1 U4508 ( .A(n3986), .B(n3985), .ZN(n3993) );
  OR2_X1 U4509 ( .A1(n4781), .A2(n4887), .ZN(n3988) );
  NAND2_X1 U4510 ( .A1(n4669), .A2(n4839), .ZN(n3987) );
  NAND2_X1 U4511 ( .A1(n3988), .A2(n3987), .ZN(n4751) );
  AOI22_X1 U4512 ( .A1(n5231), .A2(n4751), .B1(REG3_REG_26__SCAN_IN), .B2(
        U3149), .ZN(n3990) );
  NAND2_X1 U4513 ( .A1(n5237), .A2(n4741), .ZN(n3989) );
  OAI211_X1 U4514 ( .C1(n5244), .C2(n4743), .A(n3990), .B(n3989), .ZN(n3991)
         );
  INV_X1 U4515 ( .A(n3991), .ZN(n3992) );
  OAI21_X1 U4516 ( .B1(n3993), .B2(n5192), .A(n3992), .ZN(U3237) );
  NAND2_X1 U4517 ( .A1(n3043), .A2(REG1_REG_31__SCAN_IN), .ZN(n3996) );
  NAND2_X1 U4518 ( .A1(n2966), .A2(REG2_REG_31__SCAN_IN), .ZN(n3995) );
  NAND2_X1 U4519 ( .A1(n2466), .A2(REG0_REG_31__SCAN_IN), .ZN(n3994) );
  AND3_X1 U4520 ( .A1(n3996), .A2(n3995), .A3(n3994), .ZN(n5282) );
  AND2_X1 U4521 ( .A1(n4000), .A2(DATAI_31_), .ZN(n5297) );
  NAND2_X1 U4522 ( .A1(n5282), .A2(n5297), .ZN(n4002) );
  NAND2_X1 U4523 ( .A1(n3043), .A2(REG1_REG_30__SCAN_IN), .ZN(n3999) );
  NAND2_X1 U4524 ( .A1(n2966), .A2(REG2_REG_30__SCAN_IN), .ZN(n3998) );
  NAND2_X1 U4525 ( .A1(n3044), .A2(REG0_REG_30__SCAN_IN), .ZN(n3997) );
  NAND3_X1 U4526 ( .A1(n3999), .A2(n3998), .A3(n3997), .ZN(n4692) );
  NAND2_X1 U4527 ( .A1(n4000), .A2(DATAI_30_), .ZN(n5295) );
  NAND2_X1 U4528 ( .A1(n4692), .A2(n5295), .ZN(n4001) );
  NAND2_X1 U4529 ( .A1(n4002), .A2(n4001), .ZN(n4144) );
  INV_X1 U4530 ( .A(n4144), .ZN(n4042) );
  INV_X1 U4531 ( .A(n5297), .ZN(n4041) );
  INV_X1 U4532 ( .A(n5282), .ZN(n4158) );
  NAND2_X1 U4533 ( .A1(n4003), .A2(n4006), .ZN(n4101) );
  NAND2_X1 U4534 ( .A1(n4005), .A2(n4004), .ZN(n4129) );
  NAND2_X1 U4535 ( .A1(n4129), .A2(n4006), .ZN(n4134) );
  OAI21_X1 U4536 ( .B1(n4007), .B2(n4101), .A(n4134), .ZN(n4009) );
  AND2_X1 U4537 ( .A1(n4838), .A2(n4868), .ZN(n4135) );
  NAND2_X1 U4538 ( .A1(n4865), .A2(n5266), .ZN(n4056) );
  AND2_X1 U4539 ( .A1(n5251), .A2(n4056), .ZN(n4015) );
  NAND2_X1 U4540 ( .A1(n4008), .A2(n4015), .ZN(n4673) );
  AOI211_X1 U4541 ( .C1(n4009), .C2(n4136), .A(n4135), .B(n4673), .ZN(n4023)
         );
  NAND2_X1 U4542 ( .A1(n4825), .A2(n4847), .ZN(n4794) );
  NOR2_X1 U4543 ( .A1(n4840), .A2(n4828), .ZN(n4797) );
  OR2_X1 U4544 ( .A1(n4794), .A2(n4797), .ZN(n4012) );
  NAND2_X1 U4545 ( .A1(n4840), .A2(n4828), .ZN(n4053) );
  NAND2_X1 U4546 ( .A1(n4824), .A2(n4802), .ZN(n4010) );
  AND2_X1 U4547 ( .A1(n4053), .A2(n4010), .ZN(n4011) );
  NAND2_X1 U4548 ( .A1(n4014), .A2(n4013), .ZN(n4016) );
  NAND2_X1 U4549 ( .A1(n4016), .A2(n4015), .ZN(n4018) );
  INV_X1 U4550 ( .A(n5266), .ZN(n4017) );
  NAND2_X1 U4551 ( .A1(n4651), .A2(n4017), .ZN(n4057) );
  NAND2_X1 U4552 ( .A1(n4018), .A2(n4057), .ZN(n4675) );
  NAND2_X1 U4553 ( .A1(n4675), .A2(n4044), .ZN(n4019) );
  NAND2_X1 U4554 ( .A1(n4653), .A2(n4696), .ZN(n4043) );
  NAND2_X1 U4555 ( .A1(n4019), .A2(n4043), .ZN(n4834) );
  NOR2_X1 U4556 ( .A1(n4825), .A2(n4847), .ZN(n4020) );
  OR2_X1 U4557 ( .A1(n4797), .A2(n4020), .ZN(n4021) );
  NOR2_X1 U4558 ( .A1(n4799), .A2(n4661), .ZN(n4680) );
  NOR2_X1 U4559 ( .A1(n4824), .A2(n4802), .ZN(n4679) );
  NOR2_X1 U4560 ( .A1(n4680), .A2(n4679), .ZN(n4140) );
  INV_X1 U4561 ( .A(n4140), .ZN(n4022) );
  AOI221_X1 U4562 ( .B1(n4023), .B2(n4678), .C1(n4677), .C2(n4678), .A(n4022), 
        .ZN(n4027) );
  OR2_X1 U4563 ( .A1(n4781), .A2(n4760), .ZN(n4024) );
  NAND2_X1 U4564 ( .A1(n4799), .A2(n4661), .ZN(n4765) );
  NAND2_X1 U4565 ( .A1(n4024), .A2(n4765), .ZN(n4681) );
  NOR2_X1 U4566 ( .A1(n4159), .A2(n4713), .ZN(n4686) );
  NOR2_X1 U4567 ( .A1(n4669), .A2(n4730), .ZN(n4685) );
  NOR2_X1 U4568 ( .A1(n4686), .A2(n4685), .ZN(n4032) );
  NAND2_X1 U4569 ( .A1(n3025), .A2(DATAI_29_), .ZN(n4698) );
  INV_X1 U4570 ( .A(n4698), .ZN(n4699) );
  OR2_X1 U4571 ( .A1(n5282), .A2(n5297), .ZN(n4092) );
  OR2_X1 U4572 ( .A1(n4692), .A2(n5295), .ZN(n4026) );
  NAND2_X1 U4573 ( .A1(n4092), .A2(n4026), .ZN(n4045) );
  AOI21_X1 U4574 ( .B1(n4030), .B2(n4699), .A(n4045), .ZN(n4031) );
  OAI211_X1 U4575 ( .C1(n4027), .C2(n4681), .A(n4032), .B(n4031), .ZN(n4038)
         );
  NAND2_X1 U4576 ( .A1(n4028), .A2(n4741), .ZN(n4055) );
  NAND2_X1 U4577 ( .A1(n4781), .A2(n4760), .ZN(n4746) );
  NAND2_X1 U4578 ( .A1(n4055), .A2(n4746), .ZN(n4684) );
  AND2_X1 U4579 ( .A1(n4159), .A2(n4713), .ZN(n4033) );
  INV_X1 U4580 ( .A(n4033), .ZN(n4029) );
  OAI21_X1 U4581 ( .B1(n4030), .B2(n4699), .A(n4029), .ZN(n4145) );
  OAI21_X1 U4582 ( .B1(n4032), .B2(n4145), .A(n4031), .ZN(n4149) );
  INV_X1 U4583 ( .A(n4709), .ZN(n4036) );
  NAND2_X1 U4584 ( .A1(n4669), .A2(n4730), .ZN(n4141) );
  INV_X1 U4585 ( .A(n4141), .ZN(n4034) );
  INV_X1 U4586 ( .A(n4724), .ZN(n4035) );
  XNOR2_X1 U4587 ( .A(n4712), .B(n4698), .ZN(n4688) );
  INV_X1 U4588 ( .A(n4688), .ZN(n4067) );
  AND2_X1 U4589 ( .A1(n4769), .A2(n4753), .ZN(n4146) );
  AND4_X1 U4590 ( .A1(n4036), .A2(n4035), .A3(n4067), .A4(n4683), .ZN(n4037)
         );
  OAI22_X1 U4591 ( .A1(n4038), .A2(n4684), .B1(n4149), .B2(n4037), .ZN(n4039)
         );
  OAI21_X1 U4592 ( .B1(n4158), .B2(n5295), .A(n4039), .ZN(n4040) );
  OAI21_X1 U4593 ( .B1(n4042), .B2(n4041), .A(n4040), .ZN(n4091) );
  NOR2_X1 U4594 ( .A1(n4045), .A2(n4144), .ZN(n4046) );
  AND2_X1 U4595 ( .A1(n4856), .A2(n4046), .ZN(n4052) );
  INV_X1 U4596 ( .A(n4765), .ZN(n4047) );
  NOR2_X1 U4597 ( .A1(n4680), .A2(n4047), .ZN(n4778) );
  NOR2_X1 U4598 ( .A1(n4709), .A2(n4724), .ZN(n4051) );
  INV_X1 U4599 ( .A(n4802), .ZN(n4048) );
  AND2_X1 U4600 ( .A1(n4824), .A2(n4048), .ZN(n4660) );
  INV_X1 U4601 ( .A(n4660), .ZN(n4050) );
  NAND2_X1 U4602 ( .A1(n4049), .A2(n4802), .ZN(n4659) );
  NAND2_X1 U4603 ( .A1(n4050), .A2(n4659), .ZN(n4798) );
  NAND4_X1 U4604 ( .A1(n4052), .A2(n4778), .A3(n4051), .A4(n4798), .ZN(n4062)
         );
  INV_X1 U4605 ( .A(n4053), .ZN(n4054) );
  INV_X1 U4606 ( .A(n4811), .ZN(n4820) );
  NAND2_X1 U4607 ( .A1(n4683), .A2(n4055), .ZN(n4739) );
  INV_X1 U4608 ( .A(n4739), .ZN(n4749) );
  NAND2_X1 U4609 ( .A1(n4057), .A2(n4056), .ZN(n5263) );
  NOR2_X1 U4610 ( .A1(n5263), .A2(n4058), .ZN(n4060) );
  NAND4_X1 U4611 ( .A1(n4820), .A2(n4749), .A3(n4060), .A4(n4059), .ZN(n4061)
         );
  NOR2_X1 U4612 ( .A1(n4062), .A2(n4061), .ZN(n4088) );
  INV_X1 U4613 ( .A(n4063), .ZN(n4066) );
  NAND4_X1 U4614 ( .A1(n4066), .A2(n4065), .A3(n4064), .A4(n5079), .ZN(n4074)
         );
  NAND2_X1 U4615 ( .A1(n2563), .A2(n4574), .ZN(n4104) );
  AND2_X1 U4616 ( .A1(n4103), .A2(n4104), .ZN(n5051) );
  NAND3_X1 U4617 ( .A1(n4068), .A2(n4067), .A3(n5051), .ZN(n4073) );
  XNOR2_X1 U4618 ( .A(n4664), .B(n4772), .ZN(n4767) );
  INV_X1 U4619 ( .A(n4767), .ZN(n4071) );
  XNOR2_X1 U4620 ( .A(n4825), .B(n4847), .ZN(n4836) );
  INV_X1 U4621 ( .A(n4836), .ZN(n4070) );
  NAND3_X1 U4622 ( .A1(n4071), .A2(n4070), .A3(n4069), .ZN(n4072) );
  NOR3_X1 U4623 ( .A1(n4074), .A2(n4073), .A3(n4072), .ZN(n4087) );
  AND2_X1 U4624 ( .A1(n4076), .A2(n4075), .ZN(n4086) );
  NAND4_X1 U4625 ( .A1(n2683), .A2(n4078), .A3(n4649), .A4(n4077), .ZN(n4084)
         );
  NAND4_X1 U4626 ( .A1(n4082), .A2(n4081), .A3(n4080), .A4(n4079), .ZN(n4083)
         );
  NOR2_X1 U4627 ( .A1(n4084), .A2(n4083), .ZN(n4085) );
  NAND4_X1 U4628 ( .A1(n4088), .A2(n4087), .A3(n4086), .A4(n4085), .ZN(n4090)
         );
  MUX2_X1 U4629 ( .A(n4091), .B(n4090), .S(n4089), .Z(n4151) );
  NAND2_X1 U4630 ( .A1(n4092), .A2(n4144), .ZN(n4148) );
  INV_X1 U4631 ( .A(n4093), .ZN(n4095) );
  NAND4_X1 U4632 ( .A1(n4095), .A2(n4126), .A3(n4094), .A4(n4128), .ZN(n4097)
         );
  AOI21_X1 U4633 ( .B1(n4098), .B2(n4097), .A(n2502), .ZN(n4102) );
  INV_X1 U4634 ( .A(n4099), .ZN(n4100) );
  OR3_X1 U4635 ( .A1(n4102), .A2(n4101), .A3(n4100), .ZN(n4133) );
  INV_X1 U4636 ( .A(n4103), .ZN(n4106) );
  OAI211_X1 U4637 ( .C1(n4106), .C2(n4957), .A(n4105), .B(n4104), .ZN(n4109)
         );
  NAND3_X1 U4638 ( .A1(n4109), .A2(n4108), .A3(n4107), .ZN(n4111) );
  OAI211_X1 U4639 ( .C1(n4113), .C2(n4112), .A(n4111), .B(n4110), .ZN(n4116)
         );
  NAND3_X1 U4640 ( .A1(n4116), .A2(n4115), .A3(n4114), .ZN(n4119) );
  NAND3_X1 U4641 ( .A1(n4119), .A2(n4118), .A3(n4117), .ZN(n4122) );
  NAND3_X1 U4642 ( .A1(n4122), .A2(n4121), .A3(n4120), .ZN(n4127) );
  INV_X1 U4643 ( .A(n4123), .ZN(n4125) );
  AOI211_X1 U4644 ( .C1(n4127), .C2(n4126), .A(n4125), .B(n4124), .ZN(n4131)
         );
  INV_X1 U4645 ( .A(n4128), .ZN(n4130) );
  NOR4_X1 U4646 ( .A1(n4131), .A2(n4130), .A3(n2502), .A4(n4129), .ZN(n4132)
         );
  AOI21_X1 U4647 ( .B1(n4134), .B2(n4133), .A(n4132), .ZN(n4137) );
  AOI211_X1 U4648 ( .C1(n4137), .C2(n4136), .A(n4135), .B(n4673), .ZN(n4138)
         );
  OAI21_X1 U4649 ( .B1(n4138), .B2(n4677), .A(n4678), .ZN(n4139) );
  AOI21_X1 U4650 ( .B1(n4140), .B2(n4139), .A(n4681), .ZN(n4142) );
  OAI21_X1 U4651 ( .B1(n4142), .B2(n4684), .A(n4141), .ZN(n4143) );
  NOR4_X1 U4652 ( .A1(n4146), .A2(n4145), .A3(n4144), .A4(n4143), .ZN(n4147)
         );
  AOI21_X1 U4653 ( .B1(n4149), .B2(n4148), .A(n4147), .ZN(n4150) );
  MUX2_X1 U4654 ( .A(n4151), .B(n4150), .S(n2941), .Z(n4152) );
  XNOR2_X1 U4655 ( .A(n4152), .B(n5006), .ZN(n4157) );
  NAND3_X1 U4656 ( .A1(n4153), .A2(n4866), .A3(n5013), .ZN(n4154) );
  OAI211_X1 U4657 ( .C1(n2576), .C2(n4156), .A(n4154), .B(B_REG_SCAN_IN), .ZN(
        n4155) );
  OAI21_X1 U4658 ( .B1(n4157), .B2(n4156), .A(n4155), .ZN(U3239) );
  MUX2_X1 U4659 ( .A(DATAO_REG_31__SCAN_IN), .B(n4158), .S(U4043), .Z(U3581)
         );
  MUX2_X1 U4660 ( .A(n4692), .B(DATAO_REG_30__SCAN_IN), .S(n5017), .Z(U3580)
         );
  MUX2_X1 U4661 ( .A(n4712), .B(DATAO_REG_29__SCAN_IN), .S(n5017), .Z(U3579)
         );
  MUX2_X1 U4662 ( .A(n4159), .B(DATAO_REG_28__SCAN_IN), .S(n5017), .Z(U3578)
         );
  MUX2_X1 U4663 ( .A(n4669), .B(DATAO_REG_27__SCAN_IN), .S(n5017), .Z(U3577)
         );
  MUX2_X1 U4664 ( .A(n4769), .B(DATAO_REG_26__SCAN_IN), .S(n5017), .Z(U3576)
         );
  XNOR2_X1 U4665 ( .A(DATAI_21_), .B(keyinput_138), .ZN(n4165) );
  XNOR2_X1 U4666 ( .A(DATAI_20_), .B(keyinput_139), .ZN(n4161) );
  XNOR2_X1 U4667 ( .A(DATAI_22_), .B(keyinput_137), .ZN(n4160) );
  NAND2_X1 U4668 ( .A1(n4161), .A2(n4160), .ZN(n4164) );
  XNOR2_X1 U4669 ( .A(DATAI_19_), .B(keyinput_140), .ZN(n4163) );
  XNOR2_X1 U4670 ( .A(DATAI_23_), .B(keyinput_136), .ZN(n4162) );
  NOR4_X1 U4671 ( .A1(n4165), .A2(n4164), .A3(n4163), .A4(n4162), .ZN(n4178)
         );
  XOR2_X1 U4672 ( .A(DATAI_26_), .B(keyinput_133), .Z(n4168) );
  XOR2_X1 U4673 ( .A(DATAI_27_), .B(keyinput_132), .Z(n4167) );
  XNOR2_X1 U4674 ( .A(DATAI_24_), .B(keyinput_135), .ZN(n4166) );
  NOR3_X1 U4675 ( .A1(n4168), .A2(n4167), .A3(n4166), .ZN(n4175) );
  XOR2_X1 U4676 ( .A(DATAI_28_), .B(keyinput_131), .Z(n4174) );
  XOR2_X1 U4677 ( .A(DATAI_25_), .B(keyinput_134), .Z(n4173) );
  XNOR2_X1 U4678 ( .A(keyinput_129), .B(DATAI_30_), .ZN(n4171) );
  XNOR2_X1 U4679 ( .A(keyinput_128), .B(DATAI_31_), .ZN(n4170) );
  XOR2_X1 U4680 ( .A(DATAI_29_), .B(keyinput_130), .Z(n4169) );
  OAI21_X1 U4681 ( .B1(n4171), .B2(n4170), .A(n4169), .ZN(n4172) );
  NAND4_X1 U4682 ( .A1(n4175), .A2(n4174), .A3(n4173), .A4(n4172), .ZN(n4177)
         );
  XNOR2_X1 U4683 ( .A(DATAI_18_), .B(keyinput_141), .ZN(n4176) );
  AOI21_X1 U4684 ( .B1(n4178), .B2(n4177), .A(n4176), .ZN(n4182) );
  XOR2_X1 U4685 ( .A(DATAI_15_), .B(keyinput_144), .Z(n4181) );
  XOR2_X1 U4686 ( .A(DATAI_17_), .B(keyinput_142), .Z(n4180) );
  XNOR2_X1 U4687 ( .A(DATAI_16_), .B(keyinput_143), .ZN(n4179) );
  NOR4_X1 U4688 ( .A1(n4182), .A2(n4181), .A3(n4180), .A4(n4179), .ZN(n4186)
         );
  XOR2_X1 U4689 ( .A(DATAI_14_), .B(keyinput_145), .Z(n4185) );
  XNOR2_X1 U4690 ( .A(DATAI_12_), .B(keyinput_147), .ZN(n4184) );
  XNOR2_X1 U4691 ( .A(DATAI_13_), .B(keyinput_146), .ZN(n4183) );
  NOR4_X1 U4692 ( .A1(n4186), .A2(n4185), .A3(n4184), .A4(n4183), .ZN(n4189)
         );
  INV_X1 U4693 ( .A(DATAI_11_), .ZN(n4418) );
  XNOR2_X1 U4694 ( .A(n4418), .B(keyinput_148), .ZN(n4188) );
  XOR2_X1 U4695 ( .A(DATAI_10_), .B(keyinput_149), .Z(n4187) );
  OAI21_X1 U4696 ( .B1(n4189), .B2(n4188), .A(n4187), .ZN(n4192) );
  XNOR2_X1 U4697 ( .A(DATAI_9_), .B(keyinput_150), .ZN(n4191) );
  XNOR2_X1 U4698 ( .A(DATAI_8_), .B(keyinput_151), .ZN(n4190) );
  NAND3_X1 U4699 ( .A1(n4192), .A2(n4191), .A3(n4190), .ZN(n4196) );
  INV_X1 U4700 ( .A(DATAI_7_), .ZN(n5126) );
  XNOR2_X1 U4701 ( .A(n5126), .B(keyinput_152), .ZN(n4195) );
  XNOR2_X1 U4702 ( .A(DATAI_5_), .B(keyinput_154), .ZN(n4194) );
  XNOR2_X1 U4703 ( .A(DATAI_6_), .B(keyinput_153), .ZN(n4193) );
  NAND4_X1 U4704 ( .A1(n4196), .A2(n4195), .A3(n4194), .A4(n4193), .ZN(n4199)
         );
  XNOR2_X1 U4705 ( .A(DATAI_3_), .B(keyinput_156), .ZN(n4198) );
  XNOR2_X1 U4706 ( .A(DATAI_4_), .B(keyinput_155), .ZN(n4197) );
  NAND3_X1 U4707 ( .A1(n4199), .A2(n4198), .A3(n4197), .ZN(n4205) );
  XNOR2_X1 U4708 ( .A(DATAI_2_), .B(keyinput_157), .ZN(n4204) );
  XOR2_X1 U4709 ( .A(DATAI_1_), .B(keyinput_158), .Z(n4202) );
  XNOR2_X1 U4710 ( .A(STATE_REG_SCAN_IN), .B(keyinput_160), .ZN(n4201) );
  XNOR2_X1 U4711 ( .A(DATAI_0_), .B(keyinput_159), .ZN(n4200) );
  NAND3_X1 U4712 ( .A1(n4202), .A2(n4201), .A3(n4200), .ZN(n4203) );
  AOI21_X1 U4713 ( .B1(n4205), .B2(n4204), .A(n4203), .ZN(n4216) );
  XNOR2_X1 U4714 ( .A(REG3_REG_7__SCAN_IN), .B(keyinput_161), .ZN(n4215) );
  XNOR2_X1 U4715 ( .A(n4206), .B(keyinput_167), .ZN(n4210) );
  XNOR2_X1 U4716 ( .A(keyinput_163), .B(REG3_REG_14__SCAN_IN), .ZN(n4209) );
  XNOR2_X1 U4717 ( .A(REG3_REG_3__SCAN_IN), .B(keyinput_166), .ZN(n4208) );
  XNOR2_X1 U4718 ( .A(REG3_REG_23__SCAN_IN), .B(keyinput_164), .ZN(n4207) );
  NAND4_X1 U4719 ( .A1(n4210), .A2(n4209), .A3(n4208), .A4(n4207), .ZN(n4213)
         );
  XNOR2_X1 U4720 ( .A(REG3_REG_27__SCAN_IN), .B(keyinput_162), .ZN(n4212) );
  XNOR2_X1 U4721 ( .A(REG3_REG_10__SCAN_IN), .B(keyinput_165), .ZN(n4211) );
  NOR3_X1 U4722 ( .A1(n4213), .A2(n4212), .A3(n4211), .ZN(n4214) );
  OAI21_X1 U4723 ( .B1(n4216), .B2(n4215), .A(n4214), .ZN(n4219) );
  XNOR2_X1 U4724 ( .A(REG3_REG_28__SCAN_IN), .B(keyinput_168), .ZN(n4218) );
  XNOR2_X1 U4725 ( .A(REG3_REG_8__SCAN_IN), .B(keyinput_169), .ZN(n4217) );
  AOI21_X1 U4726 ( .B1(n4219), .B2(n4218), .A(n4217), .ZN(n4233) );
  OAI22_X1 U4727 ( .A1(REG3_REG_25__SCAN_IN), .A2(keyinput_173), .B1(
        REG3_REG_12__SCAN_IN), .B2(keyinput_172), .ZN(n4232) );
  OAI22_X1 U4728 ( .A1(n4220), .A2(keyinput_170), .B1(REG3_REG_16__SCAN_IN), 
        .B2(keyinput_174), .ZN(n4231) );
  INV_X1 U4729 ( .A(REG3_REG_17__SCAN_IN), .ZN(n4643) );
  OAI22_X1 U4730 ( .A1(keyinput_171), .A2(n4221), .B1(n4643), .B2(keyinput_176), .ZN(n4229) );
  NOR2_X1 U4731 ( .A1(n4370), .A2(keyinput_175), .ZN(n4228) );
  NOR2_X1 U4732 ( .A1(REG3_REG_24__SCAN_IN), .A2(keyinput_177), .ZN(n4227) );
  AOI22_X1 U4733 ( .A1(n4221), .A2(keyinput_171), .B1(keyinput_170), .B2(n4220), .ZN(n4225) );
  AOI22_X1 U4734 ( .A1(n4643), .A2(keyinput_176), .B1(n4370), .B2(keyinput_175), .ZN(n4224) );
  AOI22_X1 U4735 ( .A1(REG3_REG_25__SCAN_IN), .A2(keyinput_173), .B1(
        REG3_REG_24__SCAN_IN), .B2(keyinput_177), .ZN(n4223) );
  AOI22_X1 U4736 ( .A1(REG3_REG_16__SCAN_IN), .A2(keyinput_174), .B1(
        REG3_REG_12__SCAN_IN), .B2(keyinput_172), .ZN(n4222) );
  NAND4_X1 U4737 ( .A1(n4225), .A2(n4224), .A3(n4223), .A4(n4222), .ZN(n4226)
         );
  OR4_X1 U4738 ( .A1(n4229), .A2(n4228), .A3(n4227), .A4(n4226), .ZN(n4230) );
  NOR4_X1 U4739 ( .A1(n4233), .A2(n4232), .A3(n4231), .A4(n4230), .ZN(n4238)
         );
  XOR2_X1 U4740 ( .A(REG3_REG_4__SCAN_IN), .B(keyinput_178), .Z(n4237) );
  XNOR2_X1 U4741 ( .A(n4234), .B(keyinput_179), .ZN(n4236) );
  XNOR2_X1 U4742 ( .A(REG3_REG_0__SCAN_IN), .B(keyinput_180), .ZN(n4235) );
  OAI211_X1 U4743 ( .C1(n4238), .C2(n4237), .A(n4236), .B(n4235), .ZN(n4241)
         );
  XOR2_X1 U4744 ( .A(REG3_REG_20__SCAN_IN), .B(keyinput_181), .Z(n4240) );
  XOR2_X1 U4745 ( .A(keyinput_182), .B(REG3_REG_13__SCAN_IN), .Z(n4239) );
  AOI21_X1 U4746 ( .B1(n4241), .B2(n4240), .A(n4239), .ZN(n4244) );
  XNOR2_X1 U4747 ( .A(IR_REG_0__SCAN_IN), .B(keyinput_183), .ZN(n4243) );
  OAI21_X1 U4748 ( .B1(n4244), .B2(n4243), .A(n4242), .ZN(n4253) );
  XNOR2_X1 U4749 ( .A(n4456), .B(keyinput_186), .ZN(n4249) );
  XNOR2_X1 U4750 ( .A(n4245), .B(keyinput_185), .ZN(n4248) );
  XNOR2_X1 U4751 ( .A(IR_REG_4__SCAN_IN), .B(keyinput_187), .ZN(n4247) );
  XNOR2_X1 U4752 ( .A(IR_REG_5__SCAN_IN), .B(keyinput_188), .ZN(n4246) );
  NOR4_X1 U4753 ( .A1(n4249), .A2(n4248), .A3(n4247), .A4(n4246), .ZN(n4252)
         );
  XNOR2_X1 U4754 ( .A(n4250), .B(keyinput_189), .ZN(n4251) );
  AOI21_X1 U4755 ( .B1(n4253), .B2(n4252), .A(n4251), .ZN(n4258) );
  XNOR2_X1 U4756 ( .A(n4254), .B(keyinput_190), .ZN(n4257) );
  XNOR2_X1 U4757 ( .A(n4255), .B(keyinput_191), .ZN(n4256) );
  OAI21_X1 U4758 ( .B1(n4258), .B2(n4257), .A(n4256), .ZN(n4263) );
  XNOR2_X1 U4759 ( .A(n4259), .B(keyinput_192), .ZN(n4262) );
  XOR2_X1 U4760 ( .A(IR_REG_10__SCAN_IN), .B(keyinput_193), .Z(n4261) );
  XNOR2_X1 U4761 ( .A(n4470), .B(keyinput_194), .ZN(n4260) );
  NAND4_X1 U4762 ( .A1(n4263), .A2(n4262), .A3(n4261), .A4(n4260), .ZN(n4268)
         );
  XNOR2_X1 U4763 ( .A(n4264), .B(keyinput_195), .ZN(n4267) );
  XNOR2_X1 U4764 ( .A(n4265), .B(keyinput_196), .ZN(n4266) );
  AOI21_X1 U4765 ( .B1(n4268), .B2(n4267), .A(n4266), .ZN(n4273) );
  XNOR2_X1 U4766 ( .A(n4269), .B(keyinput_197), .ZN(n4272) );
  XNOR2_X1 U4767 ( .A(IR_REG_16__SCAN_IN), .B(keyinput_199), .ZN(n4271) );
  XNOR2_X1 U4768 ( .A(IR_REG_15__SCAN_IN), .B(keyinput_198), .ZN(n4270) );
  NOR4_X1 U4769 ( .A1(n4273), .A2(n4272), .A3(n4271), .A4(n4270), .ZN(n4280)
         );
  XNOR2_X1 U4770 ( .A(IR_REG_18__SCAN_IN), .B(keyinput_201), .ZN(n4277) );
  XNOR2_X1 U4771 ( .A(IR_REG_17__SCAN_IN), .B(keyinput_200), .ZN(n4276) );
  XNOR2_X1 U4772 ( .A(IR_REG_19__SCAN_IN), .B(keyinput_202), .ZN(n4275) );
  XNOR2_X1 U4773 ( .A(IR_REG_20__SCAN_IN), .B(keyinput_203), .ZN(n4274) );
  NAND4_X1 U4774 ( .A1(n4277), .A2(n4276), .A3(n4275), .A4(n4274), .ZN(n4279)
         );
  XNOR2_X1 U4775 ( .A(IR_REG_21__SCAN_IN), .B(keyinput_204), .ZN(n4278) );
  OAI21_X1 U4776 ( .B1(n4280), .B2(n4279), .A(n4278), .ZN(n4284) );
  XNOR2_X1 U4777 ( .A(n2790), .B(keyinput_205), .ZN(n4283) );
  XNOR2_X1 U4778 ( .A(IR_REG_24__SCAN_IN), .B(keyinput_207), .ZN(n4282) );
  XNOR2_X1 U4779 ( .A(IR_REG_23__SCAN_IN), .B(keyinput_206), .ZN(n4281) );
  AOI211_X1 U4780 ( .C1(n4284), .C2(n4283), .A(n4282), .B(n4281), .ZN(n4288)
         );
  XNOR2_X1 U4781 ( .A(IR_REG_25__SCAN_IN), .B(keyinput_208), .ZN(n4287) );
  XNOR2_X1 U4782 ( .A(n4285), .B(keyinput_209), .ZN(n4286) );
  OAI21_X1 U4783 ( .B1(n4288), .B2(n4287), .A(n4286), .ZN(n4291) );
  XNOR2_X1 U4784 ( .A(IR_REG_27__SCAN_IN), .B(keyinput_210), .ZN(n4290) );
  XNOR2_X1 U4785 ( .A(IR_REG_28__SCAN_IN), .B(keyinput_211), .ZN(n4289) );
  NAND3_X1 U4786 ( .A1(n4291), .A2(n4290), .A3(n4289), .ZN(n4295) );
  XNOR2_X1 U4787 ( .A(n4292), .B(keyinput_212), .ZN(n4294) );
  XNOR2_X1 U4788 ( .A(IR_REG_30__SCAN_IN), .B(keyinput_213), .ZN(n4293) );
  NAND3_X1 U4789 ( .A1(n4295), .A2(n4294), .A3(n4293), .ZN(n4309) );
  INV_X1 U4790 ( .A(D_REG_3__SCAN_IN), .ZN(n4973) );
  OAI22_X1 U4791 ( .A1(n4973), .A2(keyinput_218), .B1(D_REG_0__SCAN_IN), .B2(
        keyinput_215), .ZN(n4296) );
  AOI221_X1 U4792 ( .B1(n4973), .B2(keyinput_218), .C1(keyinput_215), .C2(
        D_REG_0__SCAN_IN), .A(n4296), .ZN(n4308) );
  OAI22_X1 U4793 ( .A1(D_REG_1__SCAN_IN), .A2(keyinput_216), .B1(
        D_REG_4__SCAN_IN), .B2(keyinput_219), .ZN(n4297) );
  AOI221_X1 U4794 ( .B1(D_REG_1__SCAN_IN), .B2(keyinput_216), .C1(keyinput_219), .C2(D_REG_4__SCAN_IN), .A(n4297), .ZN(n4298) );
  INV_X1 U4795 ( .A(n4298), .ZN(n4306) );
  XNOR2_X1 U4796 ( .A(D_REG_6__SCAN_IN), .B(keyinput_221), .ZN(n4305) );
  XNOR2_X1 U4797 ( .A(IR_REG_31__SCAN_IN), .B(keyinput_214), .ZN(n4304) );
  INV_X1 U4798 ( .A(keyinput_220), .ZN(n4299) );
  XNOR2_X1 U4799 ( .A(n4299), .B(D_REG_5__SCAN_IN), .ZN(n4302) );
  XNOR2_X1 U4800 ( .A(keyinput_222), .B(D_REG_7__SCAN_IN), .ZN(n4301) );
  XNOR2_X1 U4801 ( .A(keyinput_217), .B(D_REG_2__SCAN_IN), .ZN(n4300) );
  NAND3_X1 U4802 ( .A1(n4302), .A2(n4301), .A3(n4300), .ZN(n4303) );
  NOR4_X1 U4803 ( .A1(n4306), .A2(n4305), .A3(n4304), .A4(n4303), .ZN(n4307)
         );
  NAND3_X1 U4804 ( .A1(n4309), .A2(n4308), .A3(n4307), .ZN(n4324) );
  INV_X1 U4805 ( .A(D_REG_8__SCAN_IN), .ZN(n4316) );
  INV_X1 U4806 ( .A(keyinput_223), .ZN(n4315) );
  INV_X1 U4807 ( .A(D_REG_14__SCAN_IN), .ZN(n4979) );
  INV_X1 U4808 ( .A(D_REG_11__SCAN_IN), .ZN(n4978) );
  AOI22_X1 U4809 ( .A1(n4979), .A2(keyinput_229), .B1(n4978), .B2(keyinput_226), .ZN(n4313) );
  INV_X1 U4810 ( .A(D_REG_9__SCAN_IN), .ZN(n4976) );
  INV_X1 U4811 ( .A(D_REG_10__SCAN_IN), .ZN(n4977) );
  AOI22_X1 U4812 ( .A1(n4976), .A2(keyinput_224), .B1(n4977), .B2(keyinput_225), .ZN(n4312) );
  AOI22_X1 U4813 ( .A1(D_REG_13__SCAN_IN), .A2(keyinput_228), .B1(
        D_REG_8__SCAN_IN), .B2(keyinput_223), .ZN(n4311) );
  AOI22_X1 U4814 ( .A1(D_REG_15__SCAN_IN), .A2(keyinput_230), .B1(
        D_REG_12__SCAN_IN), .B2(keyinput_227), .ZN(n4310) );
  NAND4_X1 U4815 ( .A1(n4313), .A2(n4312), .A3(n4311), .A4(n4310), .ZN(n4314)
         );
  AOI21_X1 U4816 ( .B1(n4316), .B2(n4315), .A(n4314), .ZN(n4317) );
  OAI21_X1 U4817 ( .B1(keyinput_230), .B2(D_REG_15__SCAN_IN), .A(n4317), .ZN(
        n4321) );
  OAI22_X1 U4818 ( .A1(keyinput_224), .A2(n4976), .B1(n4977), .B2(keyinput_225), .ZN(n4320) );
  OAI22_X1 U4819 ( .A1(n4978), .A2(keyinput_226), .B1(keyinput_228), .B2(
        D_REG_13__SCAN_IN), .ZN(n4319) );
  OAI22_X1 U4820 ( .A1(n4979), .A2(keyinput_229), .B1(keyinput_227), .B2(
        D_REG_12__SCAN_IN), .ZN(n4318) );
  NOR4_X1 U4821 ( .A1(n4321), .A2(n4320), .A3(n4319), .A4(n4318), .ZN(n4323)
         );
  XNOR2_X1 U4822 ( .A(D_REG_16__SCAN_IN), .B(keyinput_231), .ZN(n4322) );
  AOI21_X1 U4823 ( .B1(n4324), .B2(n4323), .A(n4322), .ZN(n4328) );
  XNOR2_X1 U4824 ( .A(keyinput_232), .B(D_REG_17__SCAN_IN), .ZN(n4327) );
  XOR2_X1 U4825 ( .A(D_REG_18__SCAN_IN), .B(keyinput_233), .Z(n4326) );
  XOR2_X1 U4826 ( .A(D_REG_19__SCAN_IN), .B(keyinput_234), .Z(n4325) );
  OAI211_X1 U4827 ( .C1(n4328), .C2(n4327), .A(n4326), .B(n4325), .ZN(n4332)
         );
  XNOR2_X1 U4828 ( .A(keyinput_235), .B(D_REG_20__SCAN_IN), .ZN(n4331) );
  XOR2_X1 U4829 ( .A(keyinput_237), .B(D_REG_22__SCAN_IN), .Z(n4330) );
  XNOR2_X1 U4830 ( .A(D_REG_21__SCAN_IN), .B(keyinput_236), .ZN(n4329) );
  AOI211_X1 U4831 ( .C1(n4332), .C2(n4331), .A(n4330), .B(n4329), .ZN(n4349)
         );
  XOR2_X1 U4832 ( .A(D_REG_27__SCAN_IN), .B(keyinput_242), .Z(n4342) );
  INV_X1 U4833 ( .A(keyinput_244), .ZN(n4333) );
  NAND2_X1 U4834 ( .A1(n4333), .A2(D_REG_29__SCAN_IN), .ZN(n4338) );
  INV_X1 U4835 ( .A(D_REG_24__SCAN_IN), .ZN(n4983) );
  INV_X1 U4836 ( .A(D_REG_29__SCAN_IN), .ZN(n4985) );
  AOI22_X1 U4837 ( .A1(n4983), .A2(keyinput_239), .B1(n4985), .B2(keyinput_244), .ZN(n4336) );
  AOI22_X1 U4838 ( .A1(D_REG_23__SCAN_IN), .A2(keyinput_238), .B1(
        D_REG_26__SCAN_IN), .B2(keyinput_241), .ZN(n4335) );
  AOI22_X1 U4839 ( .A1(D_REG_25__SCAN_IN), .A2(keyinput_240), .B1(
        D_REG_28__SCAN_IN), .B2(keyinput_243), .ZN(n4334) );
  AND3_X1 U4840 ( .A1(n4336), .A2(n4335), .A3(n4334), .ZN(n4337) );
  OAI211_X1 U4841 ( .C1(keyinput_238), .C2(D_REG_23__SCAN_IN), .A(n4338), .B(
        n4337), .ZN(n4341) );
  OAI22_X1 U4842 ( .A1(n4983), .A2(keyinput_239), .B1(keyinput_241), .B2(
        D_REG_26__SCAN_IN), .ZN(n4340) );
  OAI22_X1 U4843 ( .A1(keyinput_240), .A2(D_REG_25__SCAN_IN), .B1(keyinput_243), .B2(D_REG_28__SCAN_IN), .ZN(n4339) );
  OR4_X1 U4844 ( .A1(n4342), .A2(n4341), .A3(n4340), .A4(n4339), .ZN(n4348) );
  INV_X1 U4845 ( .A(D_REG_30__SCAN_IN), .ZN(n4986) );
  XNOR2_X1 U4846 ( .A(n4986), .B(keyinput_245), .ZN(n4346) );
  XNOR2_X1 U4847 ( .A(REG0_REG_1__SCAN_IN), .B(keyinput_248), .ZN(n4345) );
  XNOR2_X1 U4848 ( .A(REG0_REG_0__SCAN_IN), .B(keyinput_247), .ZN(n4344) );
  XNOR2_X1 U4849 ( .A(D_REG_31__SCAN_IN), .B(keyinput_246), .ZN(n4343) );
  NOR4_X1 U4850 ( .A1(n4346), .A2(n4345), .A3(n4344), .A4(n4343), .ZN(n4347)
         );
  OAI21_X1 U4851 ( .B1(n4349), .B2(n4348), .A(n4347), .ZN(n4353) );
  XOR2_X1 U4852 ( .A(REG0_REG_3__SCAN_IN), .B(keyinput_250), .Z(n4352) );
  XNOR2_X1 U4853 ( .A(REG0_REG_2__SCAN_IN), .B(keyinput_249), .ZN(n4351) );
  XNOR2_X1 U4854 ( .A(REG0_REG_4__SCAN_IN), .B(keyinput_251), .ZN(n4350) );
  NAND4_X1 U4855 ( .A1(n4353), .A2(n4352), .A3(n4351), .A4(n4350), .ZN(n4357)
         );
  XOR2_X1 U4856 ( .A(REG0_REG_6__SCAN_IN), .B(keyinput_253), .Z(n4356) );
  XOR2_X1 U4857 ( .A(REG0_REG_7__SCAN_IN), .B(keyinput_254), .Z(n4355) );
  XNOR2_X1 U4858 ( .A(REG0_REG_5__SCAN_IN), .B(keyinput_252), .ZN(n4354) );
  AND4_X1 U4859 ( .A1(n4357), .A2(n4356), .A3(n4355), .A4(n4354), .ZN(n4557)
         );
  XNOR2_X1 U4860 ( .A(REG0_REG_8__SCAN_IN), .B(keyinput_255), .ZN(n4556) );
  XOR2_X1 U4861 ( .A(D_REG_23__SCAN_IN), .B(keyinput_110), .Z(n4364) );
  INV_X1 U4862 ( .A(D_REG_26__SCAN_IN), .ZN(n4984) );
  AOI22_X1 U4863 ( .A1(D_REG_25__SCAN_IN), .A2(keyinput_112), .B1(n4984), .B2(
        keyinput_113), .ZN(n4358) );
  OAI221_X1 U4864 ( .B1(D_REG_25__SCAN_IN), .B2(keyinput_112), .C1(n4984), 
        .C2(keyinput_113), .A(n4358), .ZN(n4363) );
  AOI22_X1 U4865 ( .A1(D_REG_28__SCAN_IN), .A2(keyinput_115), .B1(
        D_REG_27__SCAN_IN), .B2(keyinput_114), .ZN(n4359) );
  OAI221_X1 U4866 ( .B1(D_REG_28__SCAN_IN), .B2(keyinput_115), .C1(
        D_REG_27__SCAN_IN), .C2(keyinput_114), .A(n4359), .ZN(n4362) );
  AOI22_X1 U4867 ( .A1(D_REG_24__SCAN_IN), .A2(keyinput_111), .B1(
        D_REG_29__SCAN_IN), .B2(keyinput_116), .ZN(n4360) );
  OAI221_X1 U4868 ( .B1(D_REG_24__SCAN_IN), .B2(keyinput_111), .C1(
        D_REG_29__SCAN_IN), .C2(keyinput_116), .A(n4360), .ZN(n4361) );
  NOR4_X1 U4869 ( .A1(n4364), .A2(n4363), .A3(n4362), .A4(n4361), .ZN(n4548)
         );
  INV_X1 U4870 ( .A(keyinput_104), .ZN(n4536) );
  INV_X1 U4871 ( .A(D_REG_17__SCAN_IN), .ZN(n4980) );
  INV_X1 U4872 ( .A(keyinput_54), .ZN(n4450) );
  OAI22_X1 U4873 ( .A1(n4996), .A2(keyinput_52), .B1(REG3_REG_9__SCAN_IN), 
        .B2(keyinput_51), .ZN(n4365) );
  AOI221_X1 U4874 ( .B1(n4996), .B2(keyinput_52), .C1(keyinput_51), .C2(
        REG3_REG_9__SCAN_IN), .A(n4365), .ZN(n4448) );
  AOI22_X1 U4875 ( .A1(n4368), .A2(keyinput_45), .B1(n4367), .B2(keyinput_46), 
        .ZN(n4366) );
  OAI221_X1 U4876 ( .B1(n4368), .B2(keyinput_45), .C1(n4367), .C2(keyinput_46), 
        .A(n4366), .ZN(n4376) );
  AOI22_X1 U4877 ( .A1(n3956), .A2(keyinput_49), .B1(n4370), .B2(keyinput_47), 
        .ZN(n4369) );
  OAI221_X1 U4878 ( .B1(n3956), .B2(keyinput_49), .C1(n4370), .C2(keyinput_47), 
        .A(n4369), .ZN(n4375) );
  AOI22_X1 U4879 ( .A1(REG3_REG_21__SCAN_IN), .A2(keyinput_43), .B1(
        REG3_REG_17__SCAN_IN), .B2(keyinput_48), .ZN(n4371) );
  OAI221_X1 U4880 ( .B1(REG3_REG_21__SCAN_IN), .B2(keyinput_43), .C1(
        REG3_REG_17__SCAN_IN), .C2(keyinput_48), .A(n4371), .ZN(n4374) );
  AOI22_X1 U4881 ( .A1(REG3_REG_1__SCAN_IN), .A2(keyinput_42), .B1(
        REG3_REG_12__SCAN_IN), .B2(keyinput_44), .ZN(n4372) );
  OAI221_X1 U4882 ( .B1(REG3_REG_1__SCAN_IN), .B2(keyinput_42), .C1(
        REG3_REG_12__SCAN_IN), .C2(keyinput_44), .A(n4372), .ZN(n4373) );
  NOR4_X1 U4883 ( .A1(n4376), .A2(n4375), .A3(n4374), .A4(n4373), .ZN(n4446)
         );
  INV_X1 U4884 ( .A(keyinput_41), .ZN(n4444) );
  INV_X1 U4885 ( .A(keyinput_40), .ZN(n4441) );
  OAI22_X1 U4886 ( .A1(REG3_REG_14__SCAN_IN), .A2(keyinput_35), .B1(
        REG3_REG_19__SCAN_IN), .B2(keyinput_39), .ZN(n4377) );
  AOI221_X1 U4887 ( .B1(REG3_REG_14__SCAN_IN), .B2(keyinput_35), .C1(
        keyinput_39), .C2(REG3_REG_19__SCAN_IN), .A(n4377), .ZN(n4438) );
  OAI22_X1 U4888 ( .A1(n5096), .A2(keyinput_38), .B1(keyinput_37), .B2(
        REG3_REG_10__SCAN_IN), .ZN(n4378) );
  AOI221_X1 U4889 ( .B1(n5096), .B2(keyinput_38), .C1(REG3_REG_10__SCAN_IN), 
        .C2(keyinput_37), .A(n4378), .ZN(n4437) );
  OAI22_X1 U4890 ( .A1(n4381), .A2(keyinput_36), .B1(n4380), .B2(keyinput_34), 
        .ZN(n4379) );
  AOI221_X1 U4891 ( .B1(n4381), .B2(keyinput_36), .C1(keyinput_34), .C2(n4380), 
        .A(n4379), .ZN(n4436) );
  INV_X1 U4892 ( .A(keyinput_33), .ZN(n4433) );
  INV_X1 U4893 ( .A(DATAI_2_), .ZN(n4428) );
  INV_X1 U4894 ( .A(DATAI_4_), .ZN(n5104) );
  AOI22_X1 U4895 ( .A1(DATAI_3_), .A2(keyinput_28), .B1(n5104), .B2(
        keyinput_27), .ZN(n4382) );
  OAI221_X1 U4896 ( .B1(DATAI_3_), .B2(keyinput_28), .C1(n5104), .C2(
        keyinput_27), .A(n4382), .ZN(n4427) );
  INV_X1 U4897 ( .A(DATAI_8_), .ZN(n5133) );
  OAI22_X1 U4898 ( .A1(n5133), .A2(keyinput_23), .B1(DATAI_9_), .B2(
        keyinput_22), .ZN(n4383) );
  AOI221_X1 U4899 ( .B1(n5133), .B2(keyinput_23), .C1(keyinput_22), .C2(
        DATAI_9_), .A(n4383), .ZN(n4426) );
  INV_X1 U4900 ( .A(DATAI_10_), .ZN(n5150) );
  INV_X1 U4901 ( .A(keyinput_21), .ZN(n4420) );
  INV_X1 U4902 ( .A(keyinput_20), .ZN(n4417) );
  INV_X1 U4903 ( .A(DATAI_17_), .ZN(n4410) );
  INV_X1 U4904 ( .A(DATAI_16_), .ZN(n4386) );
  INV_X1 U4905 ( .A(DATAI_15_), .ZN(n4385) );
  OAI22_X1 U4906 ( .A1(n4386), .A2(keyinput_15), .B1(n4385), .B2(keyinput_16), 
        .ZN(n4384) );
  AOI221_X1 U4907 ( .B1(n4386), .B2(keyinput_15), .C1(keyinput_16), .C2(n4385), 
        .A(n4384), .ZN(n4409) );
  INV_X1 U4908 ( .A(DATAI_18_), .ZN(n5228) );
  XOR2_X1 U4909 ( .A(DATAI_23_), .B(keyinput_8), .Z(n4389) );
  XNOR2_X1 U4910 ( .A(DATAI_20_), .B(keyinput_11), .ZN(n4388) );
  XNOR2_X1 U4911 ( .A(DATAI_22_), .B(keyinput_9), .ZN(n4387) );
  NAND3_X1 U4912 ( .A1(n4389), .A2(n4388), .A3(n4387), .ZN(n4393) );
  INV_X1 U4913 ( .A(DATAI_21_), .ZN(n4390) );
  XNOR2_X1 U4914 ( .A(keyinput_10), .B(n4390), .ZN(n4392) );
  XNOR2_X1 U4915 ( .A(DATAI_19_), .B(keyinput_12), .ZN(n4391) );
  NOR3_X1 U4916 ( .A1(n4393), .A2(n4392), .A3(n4391), .ZN(n4408) );
  OAI22_X1 U4917 ( .A1(DATAI_26_), .A2(keyinput_5), .B1(DATAI_25_), .B2(
        keyinput_6), .ZN(n4394) );
  AOI221_X1 U4918 ( .B1(DATAI_26_), .B2(keyinput_5), .C1(keyinput_6), .C2(
        DATAI_25_), .A(n4394), .ZN(n4406) );
  INV_X1 U4919 ( .A(DATAI_27_), .ZN(n4397) );
  INV_X1 U4920 ( .A(DATAI_24_), .ZN(n4396) );
  OAI22_X1 U4921 ( .A1(n4397), .A2(keyinput_4), .B1(n4396), .B2(keyinput_7), 
        .ZN(n4395) );
  AOI221_X1 U4922 ( .B1(n4397), .B2(keyinput_4), .C1(keyinput_7), .C2(n4396), 
        .A(n4395), .ZN(n4405) );
  INV_X1 U4923 ( .A(keyinput_2), .ZN(n4401) );
  INV_X1 U4924 ( .A(DATAI_29_), .ZN(n4400) );
  AOI22_X1 U4925 ( .A1(DATAI_31_), .A2(keyinput_0), .B1(DATAI_30_), .B2(
        keyinput_1), .ZN(n4398) );
  OAI221_X1 U4926 ( .B1(DATAI_31_), .B2(keyinput_0), .C1(DATAI_30_), .C2(
        keyinput_1), .A(n4398), .ZN(n4399) );
  OAI221_X1 U4927 ( .B1(DATAI_29_), .B2(n4401), .C1(n4400), .C2(keyinput_2), 
        .A(n4399), .ZN(n4404) );
  XOR2_X1 U4928 ( .A(n4402), .B(keyinput_3), .Z(n4403) );
  NAND4_X1 U4929 ( .A1(n4406), .A2(n4405), .A3(n4404), .A4(n4403), .ZN(n4407)
         );
  INV_X1 U4930 ( .A(DATAI_14_), .ZN(n4412) );
  AOI22_X1 U4931 ( .A1(DATAI_12_), .A2(keyinput_19), .B1(n4412), .B2(
        keyinput_17), .ZN(n4411) );
  OAI221_X1 U4932 ( .B1(DATAI_12_), .B2(keyinput_19), .C1(n4412), .C2(
        keyinput_17), .A(n4411), .ZN(n4413) );
  AOI211_X1 U4933 ( .C1(DATAI_13_), .C2(keyinput_18), .A(n4414), .B(n4413), 
        .ZN(n4415) );
  OAI21_X1 U4934 ( .B1(DATAI_13_), .B2(keyinput_18), .A(n4415), .ZN(n4416) );
  OAI221_X1 U4935 ( .B1(DATAI_11_), .B2(keyinput_20), .C1(n4418), .C2(n4417), 
        .A(n4416), .ZN(n4419) );
  OAI221_X1 U4936 ( .B1(DATAI_10_), .B2(keyinput_21), .C1(n5150), .C2(n4420), 
        .A(n4419), .ZN(n4425) );
  INV_X1 U4937 ( .A(DATAI_6_), .ZN(n4421) );
  XNOR2_X1 U4938 ( .A(n4421), .B(keyinput_25), .ZN(n4424) );
  AOI22_X1 U4939 ( .A1(DATAI_5_), .A2(keyinput_26), .B1(DATAI_7_), .B2(
        keyinput_24), .ZN(n4422) );
  OAI221_X1 U4940 ( .B1(DATAI_5_), .B2(keyinput_26), .C1(DATAI_7_), .C2(
        keyinput_24), .A(n4422), .ZN(n4423) );
  AOI22_X1 U4941 ( .A1(DATAI_0_), .A2(keyinput_31), .B1(DATAI_1_), .B2(
        keyinput_30), .ZN(n4429) );
  OAI221_X1 U4942 ( .B1(DATAI_0_), .B2(keyinput_31), .C1(DATAI_1_), .C2(
        keyinput_30), .A(n4429), .ZN(n4430) );
  OAI21_X1 U4943 ( .B1(U3149), .B2(keyinput_32), .A(n4431), .ZN(n4432) );
  OAI221_X1 U4944 ( .B1(REG3_REG_7__SCAN_IN), .B2(keyinput_33), .C1(n4434), 
        .C2(n4433), .A(n4432), .ZN(n4435) );
  NAND4_X1 U4945 ( .A1(n4438), .A2(n4437), .A3(n4436), .A4(n4435), .ZN(n4439)
         );
  OAI221_X1 U4946 ( .B1(REG3_REG_28__SCAN_IN), .B2(n4441), .C1(n4440), .C2(
        keyinput_40), .A(n4439), .ZN(n4442) );
  OAI221_X1 U4947 ( .B1(REG3_REG_8__SCAN_IN), .B2(n4444), .C1(n4443), .C2(
        keyinput_41), .A(n4442), .ZN(n4445) );
  OAI221_X1 U4948 ( .B1(REG3_REG_13__SCAN_IN), .B2(keyinput_54), .C1(n4451), 
        .C2(n4450), .A(n4449), .ZN(n4454) );
  INV_X1 U4949 ( .A(keyinput_55), .ZN(n4452) );
  MUX2_X1 U4950 ( .A(n4452), .B(keyinput_55), .S(IR_REG_0__SCAN_IN), .Z(n4453)
         );
  NAND2_X1 U4951 ( .A1(n4454), .A2(n4453), .ZN(n4462) );
  AOI22_X1 U4952 ( .A1(IR_REG_4__SCAN_IN), .A2(keyinput_59), .B1(n4456), .B2(
        keyinput_58), .ZN(n4455) );
  OAI221_X1 U4953 ( .B1(IR_REG_4__SCAN_IN), .B2(keyinput_59), .C1(n4456), .C2(
        keyinput_58), .A(n4455), .ZN(n4460) );
  XNOR2_X1 U4954 ( .A(IR_REG_2__SCAN_IN), .B(keyinput_57), .ZN(n4458) );
  XNOR2_X1 U4955 ( .A(IR_REG_5__SCAN_IN), .B(keyinput_60), .ZN(n4457) );
  NAND2_X1 U4956 ( .A1(n4458), .A2(n4457), .ZN(n4459) );
  AOI211_X1 U4957 ( .C1(n4462), .C2(n4461), .A(n4460), .B(n4459), .ZN(n4465)
         );
  INV_X1 U4958 ( .A(keyinput_61), .ZN(n4463) );
  MUX2_X1 U4959 ( .A(n4463), .B(keyinput_61), .S(IR_REG_6__SCAN_IN), .Z(n4464)
         );
  NOR2_X1 U4960 ( .A1(n4465), .A2(n4464), .ZN(n4468) );
  INV_X1 U4961 ( .A(keyinput_62), .ZN(n4466) );
  MUX2_X1 U4962 ( .A(n4466), .B(keyinput_62), .S(IR_REG_7__SCAN_IN), .Z(n4467)
         );
  INV_X1 U4963 ( .A(keyinput_63), .ZN(n4469) );
  MUX2_X1 U4964 ( .A(keyinput_63), .B(n4469), .S(IR_REG_8__SCAN_IN), .Z(n4475)
         );
  XNOR2_X1 U4965 ( .A(n4470), .B(keyinput_66), .ZN(n4473) );
  XNOR2_X1 U4966 ( .A(IR_REG_10__SCAN_IN), .B(keyinput_65), .ZN(n4472) );
  XNOR2_X1 U4967 ( .A(IR_REG_9__SCAN_IN), .B(keyinput_64), .ZN(n4471) );
  NOR3_X1 U4968 ( .A1(n4473), .A2(n4472), .A3(n4471), .ZN(n4474) );
  INV_X1 U4969 ( .A(keyinput_67), .ZN(n4476) );
  MUX2_X1 U4970 ( .A(n4476), .B(keyinput_67), .S(IR_REG_12__SCAN_IN), .Z(n4477) );
  INV_X1 U4971 ( .A(keyinput_68), .ZN(n4478) );
  MUX2_X1 U4972 ( .A(n4478), .B(keyinput_68), .S(IR_REG_13__SCAN_IN), .Z(n4483) );
  XNOR2_X1 U4973 ( .A(IR_REG_15__SCAN_IN), .B(keyinput_70), .ZN(n4481) );
  XNOR2_X1 U4974 ( .A(IR_REG_16__SCAN_IN), .B(keyinput_71), .ZN(n4480) );
  XNOR2_X1 U4975 ( .A(IR_REG_14__SCAN_IN), .B(keyinput_69), .ZN(n4479) );
  NAND3_X1 U4976 ( .A1(n4481), .A2(n4480), .A3(n4479), .ZN(n4482) );
  AOI22_X1 U4977 ( .A1(IR_REG_17__SCAN_IN), .A2(keyinput_72), .B1(n4485), .B2(
        keyinput_74), .ZN(n4484) );
  OAI221_X1 U4978 ( .B1(IR_REG_17__SCAN_IN), .B2(keyinput_72), .C1(n4485), 
        .C2(keyinput_74), .A(n4484), .ZN(n4489) );
  XOR2_X1 U4979 ( .A(IR_REG_18__SCAN_IN), .B(keyinput_73), .Z(n4488) );
  XNOR2_X1 U4980 ( .A(n4486), .B(keyinput_75), .ZN(n4487) );
  NOR4_X1 U4981 ( .A1(n4490), .A2(n4489), .A3(n4488), .A4(n4487), .ZN(n4493)
         );
  INV_X1 U4982 ( .A(keyinput_76), .ZN(n4491) );
  MUX2_X1 U4983 ( .A(keyinput_76), .B(n4491), .S(IR_REG_21__SCAN_IN), .Z(n4492) );
  NOR2_X1 U4984 ( .A1(n4493), .A2(n4492), .ZN(n4500) );
  INV_X1 U4985 ( .A(keyinput_77), .ZN(n4494) );
  MUX2_X1 U4986 ( .A(keyinput_77), .B(n4494), .S(IR_REG_22__SCAN_IN), .Z(n4499) );
  AOI22_X1 U4987 ( .A1(IR_REG_23__SCAN_IN), .A2(keyinput_78), .B1(n4496), .B2(
        keyinput_79), .ZN(n4495) );
  OAI221_X1 U4988 ( .B1(IR_REG_23__SCAN_IN), .B2(keyinput_78), .C1(n4496), 
        .C2(keyinput_79), .A(n4495), .ZN(n4497) );
  INV_X1 U4989 ( .A(n4497), .ZN(n4498) );
  OAI21_X1 U4990 ( .B1(n4500), .B2(n4499), .A(n4498), .ZN(n4504) );
  XOR2_X1 U4991 ( .A(IR_REG_25__SCAN_IN), .B(keyinput_80), .Z(n4503) );
  INV_X1 U4992 ( .A(keyinput_81), .ZN(n4501) );
  MUX2_X1 U4993 ( .A(keyinput_81), .B(n4501), .S(IR_REG_26__SCAN_IN), .Z(n4502) );
  AOI21_X1 U4994 ( .B1(n4504), .B2(n4503), .A(n4502), .ZN(n4509) );
  XNOR2_X1 U4995 ( .A(n4505), .B(keyinput_82), .ZN(n4508) );
  XNOR2_X1 U4996 ( .A(n4506), .B(keyinput_83), .ZN(n4507) );
  XNOR2_X1 U4997 ( .A(n4510), .B(keyinput_85), .ZN(n4512) );
  XNOR2_X1 U4998 ( .A(IR_REG_29__SCAN_IN), .B(keyinput_84), .ZN(n4511) );
  OAI22_X1 U4999 ( .A1(n4973), .A2(keyinput_90), .B1(n4514), .B2(keyinput_87), 
        .ZN(n4513) );
  AOI221_X1 U5000 ( .B1(n4973), .B2(keyinput_90), .C1(keyinput_87), .C2(n4514), 
        .A(n4513), .ZN(n4524) );
  INV_X1 U5001 ( .A(D_REG_6__SCAN_IN), .ZN(n4974) );
  OAI22_X1 U5002 ( .A1(n4974), .A2(keyinput_93), .B1(keyinput_91), .B2(
        D_REG_4__SCAN_IN), .ZN(n4515) );
  AOI221_X1 U5003 ( .B1(n4974), .B2(keyinput_93), .C1(D_REG_4__SCAN_IN), .C2(
        keyinput_91), .A(n4515), .ZN(n4523) );
  OAI22_X1 U5004 ( .A1(D_REG_1__SCAN_IN), .A2(keyinput_88), .B1(
        D_REG_5__SCAN_IN), .B2(keyinput_92), .ZN(n4516) );
  AOI221_X1 U5005 ( .B1(D_REG_1__SCAN_IN), .B2(keyinput_88), .C1(keyinput_92), 
        .C2(D_REG_5__SCAN_IN), .A(n4516), .ZN(n4522) );
  INV_X1 U5006 ( .A(D_REG_7__SCAN_IN), .ZN(n4975) );
  INV_X1 U5007 ( .A(D_REG_2__SCAN_IN), .ZN(n4972) );
  AOI22_X1 U5008 ( .A1(n4975), .A2(keyinput_94), .B1(n4972), .B2(keyinput_89), 
        .ZN(n4517) );
  OAI221_X1 U5009 ( .B1(n4975), .B2(keyinput_94), .C1(n4972), .C2(keyinput_89), 
        .A(n4517), .ZN(n4520) );
  INV_X1 U5010 ( .A(keyinput_86), .ZN(n4518) );
  XNOR2_X1 U5011 ( .A(n4518), .B(IR_REG_31__SCAN_IN), .ZN(n4519) );
  NOR2_X1 U5012 ( .A1(n4520), .A2(n4519), .ZN(n4521) );
  AOI22_X1 U5013 ( .A1(D_REG_14__SCAN_IN), .A2(keyinput_101), .B1(n4316), .B2(
        keyinput_95), .ZN(n4525) );
  OAI221_X1 U5014 ( .B1(D_REG_14__SCAN_IN), .B2(keyinput_101), .C1(n4316), 
        .C2(keyinput_95), .A(n4525), .ZN(n4532) );
  AOI22_X1 U5015 ( .A1(n4976), .A2(keyinput_96), .B1(n4977), .B2(keyinput_97), 
        .ZN(n4526) );
  OAI221_X1 U5016 ( .B1(n4976), .B2(keyinput_96), .C1(n4977), .C2(keyinput_97), 
        .A(n4526), .ZN(n4531) );
  AOI22_X1 U5017 ( .A1(D_REG_11__SCAN_IN), .A2(keyinput_98), .B1(
        D_REG_12__SCAN_IN), .B2(keyinput_99), .ZN(n4527) );
  OAI221_X1 U5018 ( .B1(D_REG_11__SCAN_IN), .B2(keyinput_98), .C1(
        D_REG_12__SCAN_IN), .C2(keyinput_99), .A(n4527), .ZN(n4530) );
  AOI22_X1 U5019 ( .A1(D_REG_13__SCAN_IN), .A2(keyinput_100), .B1(
        D_REG_15__SCAN_IN), .B2(keyinput_102), .ZN(n4528) );
  OAI221_X1 U5020 ( .B1(D_REG_13__SCAN_IN), .B2(keyinput_100), .C1(
        D_REG_15__SCAN_IN), .C2(keyinput_102), .A(n4528), .ZN(n4529) );
  NOR4_X1 U5021 ( .A1(n4532), .A2(n4531), .A3(n4530), .A4(n4529), .ZN(n4534)
         );
  NOR2_X1 U5022 ( .A1(D_REG_16__SCAN_IN), .A2(keyinput_103), .ZN(n4533) );
  AOI221_X1 U5023 ( .B1(D_REG_17__SCAN_IN), .B2(n4536), .C1(n4980), .C2(
        keyinput_104), .A(n4535), .ZN(n4539) );
  AOI22_X1 U5024 ( .A1(D_REG_18__SCAN_IN), .A2(keyinput_105), .B1(
        D_REG_19__SCAN_IN), .B2(keyinput_106), .ZN(n4537) );
  OAI221_X1 U5025 ( .B1(D_REG_18__SCAN_IN), .B2(keyinput_105), .C1(
        D_REG_19__SCAN_IN), .C2(keyinput_106), .A(n4537), .ZN(n4538) );
  OAI22_X1 U5026 ( .A1(n4539), .A2(n4538), .B1(D_REG_20__SCAN_IN), .B2(
        keyinput_107), .ZN(n4542) );
  INV_X1 U5027 ( .A(D_REG_22__SCAN_IN), .ZN(n4982) );
  OAI22_X1 U5028 ( .A1(n4982), .A2(keyinput_109), .B1(keyinput_108), .B2(
        D_REG_21__SCAN_IN), .ZN(n4540) );
  AOI221_X1 U5029 ( .B1(n4982), .B2(keyinput_109), .C1(D_REG_21__SCAN_IN), 
        .C2(keyinput_108), .A(n4540), .ZN(n4541) );
  OAI221_X1 U5030 ( .B1(n4542), .B2(keyinput_107), .C1(n4542), .C2(
        D_REG_20__SCAN_IN), .A(n4541), .ZN(n4547) );
  INV_X1 U5031 ( .A(REG0_REG_0__SCAN_IN), .ZN(n5053) );
  AOI22_X1 U5032 ( .A1(D_REG_30__SCAN_IN), .A2(keyinput_117), .B1(n5053), .B2(
        keyinput_119), .ZN(n4543) );
  OAI221_X1 U5033 ( .B1(D_REG_30__SCAN_IN), .B2(keyinput_117), .C1(n5053), 
        .C2(keyinput_119), .A(n4543), .ZN(n4546) );
  AOI22_X1 U5034 ( .A1(REG0_REG_1__SCAN_IN), .A2(keyinput_120), .B1(
        D_REG_31__SCAN_IN), .B2(keyinput_118), .ZN(n4544) );
  OAI221_X1 U5035 ( .B1(REG0_REG_1__SCAN_IN), .B2(keyinput_120), .C1(
        D_REG_31__SCAN_IN), .C2(keyinput_118), .A(n4544), .ZN(n4545) );
  INV_X1 U5036 ( .A(REG0_REG_2__SCAN_IN), .ZN(n5072) );
  AOI22_X1 U5037 ( .A1(REG0_REG_4__SCAN_IN), .A2(keyinput_123), .B1(n5072), 
        .B2(keyinput_121), .ZN(n4549) );
  OAI221_X1 U5038 ( .B1(REG0_REG_4__SCAN_IN), .B2(keyinput_123), .C1(n5072), 
        .C2(keyinput_121), .A(n4549), .ZN(n4550) );
  INV_X1 U5039 ( .A(REG0_REG_6__SCAN_IN), .ZN(n5124) );
  OAI22_X1 U5040 ( .A1(n5124), .A2(keyinput_125), .B1(REG0_REG_5__SCAN_IN), 
        .B2(keyinput_124), .ZN(n4551) );
  AOI221_X1 U5041 ( .B1(n5124), .B2(keyinput_125), .C1(keyinput_124), .C2(
        REG0_REG_5__SCAN_IN), .A(n4551), .ZN(n4553) );
  XNOR2_X1 U5042 ( .A(REG0_REG_7__SCAN_IN), .B(keyinput_126), .ZN(n4552) );
  XOR2_X1 U5043 ( .A(REG0_REG_8__SCAN_IN), .B(keyinput_127), .Z(n4554) );
  OAI211_X1 U5044 ( .C1(n4557), .C2(n4556), .A(n4555), .B(n4554), .ZN(n4559)
         );
  MUX2_X1 U5045 ( .A(DATAO_REG_25__SCAN_IN), .B(n4664), .S(U4043), .Z(n4558)
         );
  XNOR2_X1 U5046 ( .A(n4559), .B(n4558), .ZN(U3575) );
  MUX2_X1 U5047 ( .A(n4799), .B(DATAO_REG_24__SCAN_IN), .S(n5017), .Z(U3574)
         );
  MUX2_X1 U5048 ( .A(n4824), .B(DATAO_REG_23__SCAN_IN), .S(n5017), .Z(U3573)
         );
  MUX2_X1 U5049 ( .A(n4840), .B(DATAO_REG_22__SCAN_IN), .S(n5017), .Z(U3572)
         );
  MUX2_X1 U5050 ( .A(n4825), .B(DATAO_REG_21__SCAN_IN), .S(n5017), .Z(U3571)
         );
  MUX2_X1 U5051 ( .A(n4838), .B(DATAO_REG_20__SCAN_IN), .S(n5017), .Z(U3570)
         );
  MUX2_X1 U5052 ( .A(n4865), .B(DATAO_REG_19__SCAN_IN), .S(n5017), .Z(U3569)
         );
  MUX2_X1 U5053 ( .A(DATAO_REG_18__SCAN_IN), .B(n4648), .S(U4043), .Z(U3568)
         );
  MUX2_X1 U5054 ( .A(DATAO_REG_17__SCAN_IN), .B(n4560), .S(U4043), .Z(U3567)
         );
  MUX2_X1 U5055 ( .A(DATAO_REG_16__SCAN_IN), .B(n4561), .S(U4043), .Z(U3566)
         );
  MUX2_X1 U5056 ( .A(DATAO_REG_15__SCAN_IN), .B(n4562), .S(U4043), .Z(U3565)
         );
  MUX2_X1 U5057 ( .A(DATAO_REG_14__SCAN_IN), .B(n4563), .S(U4043), .Z(U3564)
         );
  MUX2_X1 U5058 ( .A(DATAO_REG_13__SCAN_IN), .B(n4564), .S(U4043), .Z(U3563)
         );
  MUX2_X1 U5059 ( .A(DATAO_REG_12__SCAN_IN), .B(n4565), .S(U4043), .Z(U3562)
         );
  MUX2_X1 U5060 ( .A(DATAO_REG_11__SCAN_IN), .B(n4566), .S(U4043), .Z(U3561)
         );
  MUX2_X1 U5061 ( .A(DATAO_REG_10__SCAN_IN), .B(n4567), .S(U4043), .Z(U3560)
         );
  MUX2_X1 U5062 ( .A(n3325), .B(DATAO_REG_9__SCAN_IN), .S(n5017), .Z(U3559) );
  MUX2_X1 U5063 ( .A(n4568), .B(DATAO_REG_8__SCAN_IN), .S(n5017), .Z(U3558) );
  MUX2_X1 U5064 ( .A(DATAO_REG_7__SCAN_IN), .B(n4569), .S(U4043), .Z(U3557) );
  MUX2_X1 U5065 ( .A(n4570), .B(DATAO_REG_6__SCAN_IN), .S(n5017), .Z(U3556) );
  MUX2_X1 U5066 ( .A(DATAO_REG_5__SCAN_IN), .B(n4571), .S(U4043), .Z(U3555) );
  MUX2_X1 U5067 ( .A(DATAO_REG_4__SCAN_IN), .B(n4572), .S(U4043), .Z(U3554) );
  MUX2_X1 U5068 ( .A(n4573), .B(DATAO_REG_3__SCAN_IN), .S(n5017), .Z(U3553) );
  MUX2_X1 U5069 ( .A(n3087), .B(DATAO_REG_2__SCAN_IN), .S(n5017), .Z(U3552) );
  MUX2_X1 U5070 ( .A(DATAO_REG_1__SCAN_IN), .B(n3064), .S(U4043), .Z(U3551) );
  MUX2_X1 U5071 ( .A(n4574), .B(DATAO_REG_0__SCAN_IN), .S(n5017), .Z(U3550) );
  XOR2_X1 U5072 ( .A(REG1_REG_12__SCAN_IN), .B(n4575), .Z(n4583) );
  AOI21_X1 U5073 ( .B1(n5036), .B2(ADDR_REG_12__SCAN_IN), .A(n4576), .ZN(n4577) );
  OAI21_X1 U5074 ( .B1(n2622), .B2(n5042), .A(n4577), .ZN(n4582) );
  AOI211_X1 U5075 ( .C1(n4580), .C2(n4578), .A(n4579), .B(n5031), .ZN(n4581)
         );
  AOI211_X1 U5076 ( .C1(n5038), .C2(n4583), .A(n4582), .B(n4581), .ZN(n4584)
         );
  INV_X1 U5077 ( .A(n4584), .ZN(U3252) );
  INV_X1 U5078 ( .A(n4964), .ZN(n4599) );
  INV_X1 U5079 ( .A(n4585), .ZN(n4589) );
  NAND2_X1 U5080 ( .A1(n4599), .A2(REG1_REG_13__SCAN_IN), .ZN(n4586) );
  OAI211_X1 U5081 ( .C1(REG1_REG_13__SCAN_IN), .C2(n4599), .A(n4587), .B(n4586), .ZN(n4588) );
  NAND3_X1 U5082 ( .A1(n4589), .A2(n5038), .A3(n4588), .ZN(n4598) );
  INV_X1 U5083 ( .A(n4590), .ZN(n4594) );
  INV_X1 U5084 ( .A(n4591), .ZN(n4592) );
  AOI211_X1 U5085 ( .C1(n4594), .C2(n4593), .A(n4592), .B(n5031), .ZN(n4595)
         );
  AOI211_X1 U5086 ( .C1(n5036), .C2(ADDR_REG_13__SCAN_IN), .A(n4596), .B(n4595), .ZN(n4597) );
  OAI211_X1 U5087 ( .C1(n5042), .C2(n4599), .A(n4598), .B(n4597), .ZN(U3253)
         );
  XOR2_X1 U5088 ( .A(REG1_REG_14__SCAN_IN), .B(n4600), .Z(n4608) );
  AOI21_X1 U5089 ( .B1(n5036), .B2(ADDR_REG_14__SCAN_IN), .A(n4601), .ZN(n4602) );
  OAI21_X1 U5090 ( .B1(n2845), .B2(n5042), .A(n4602), .ZN(n4607) );
  AOI211_X1 U5091 ( .C1(n4605), .C2(n4604), .A(n4603), .B(n5031), .ZN(n4606)
         );
  AOI211_X1 U5092 ( .C1(n5038), .C2(n4608), .A(n4607), .B(n4606), .ZN(n4609)
         );
  INV_X1 U5093 ( .A(n4609), .ZN(U3254) );
  INV_X1 U5094 ( .A(n4962), .ZN(n4621) );
  NAND2_X1 U5095 ( .A1(n4621), .A2(REG1_REG_15__SCAN_IN), .ZN(n4610) );
  OAI211_X1 U5096 ( .C1(REG1_REG_15__SCAN_IN), .C2(n4621), .A(n4611), .B(n4610), .ZN(n4612) );
  NAND3_X1 U5097 ( .A1(n2612), .A2(n5038), .A3(n4612), .ZN(n4620) );
  INV_X1 U5098 ( .A(n4613), .ZN(n4614) );
  AOI211_X1 U5099 ( .C1(n4616), .C2(n4615), .A(n4614), .B(n5031), .ZN(n4618)
         );
  AND2_X1 U5100 ( .A1(U3149), .A2(REG3_REG_15__SCAN_IN), .ZN(n4617) );
  AOI211_X1 U5101 ( .C1(n5036), .C2(ADDR_REG_15__SCAN_IN), .A(n4618), .B(n4617), .ZN(n4619) );
  OAI211_X1 U5102 ( .C1(n5042), .C2(n4621), .A(n4620), .B(n4619), .ZN(U3255)
         );
  AOI21_X1 U5103 ( .B1(REG1_REG_16__SCAN_IN), .B2(n4622), .A(n4637), .ZN(n4633) );
  NOR2_X1 U5104 ( .A1(n5042), .A2(n4623), .ZN(n4624) );
  AOI211_X1 U5105 ( .C1(n5003), .C2(ADDR_REG_16__SCAN_IN), .A(n4625), .B(n4624), .ZN(n4631) );
  AOI221_X1 U5106 ( .B1(n4628), .B2(n4626), .C1(n4627), .C2(n4626), .A(n5031), 
        .ZN(n4629) );
  INV_X1 U5107 ( .A(n4629), .ZN(n4630) );
  OAI211_X1 U5108 ( .C1(n4633), .C2(n4632), .A(n4631), .B(n4630), .ZN(U3256)
         );
  INV_X1 U5109 ( .A(n4634), .ZN(n4639) );
  NOR3_X1 U5110 ( .A1(n4637), .A2(n4636), .A3(n4635), .ZN(n4638) );
  OAI21_X1 U5111 ( .B1(n4639), .B2(n4638), .A(n5038), .ZN(n4647) );
  AOI211_X1 U5112 ( .C1(n4642), .C2(n4641), .A(n4640), .B(n5031), .ZN(n4645)
         );
  NOR2_X1 U5113 ( .A1(STATE_REG_SCAN_IN), .A2(n4643), .ZN(n4644) );
  AOI211_X1 U5114 ( .C1(n5036), .C2(ADDR_REG_17__SCAN_IN), .A(n4645), .B(n4644), .ZN(n4646) );
  OAI211_X1 U5115 ( .C1(n2619), .C2(n5042), .A(n4647), .B(n4646), .ZN(U3257)
         );
  AOI22_X1 U5116 ( .A1(n5264), .A2(n5263), .B1(n4651), .B2(n5266), .ZN(n4854)
         );
  NAND2_X1 U5117 ( .A1(n4854), .A2(n4652), .ZN(n4655) );
  NAND2_X1 U5118 ( .A1(n4655), .A2(n4654), .ZN(n4833) );
  NAND2_X1 U5119 ( .A1(n4799), .A2(n4784), .ZN(n4663) );
  NAND2_X1 U5120 ( .A1(n4759), .A2(n4767), .ZN(n4758) );
  NAND2_X1 U5121 ( .A1(n4664), .A2(n4760), .ZN(n4665) );
  NAND2_X1 U5122 ( .A1(n4758), .A2(n4665), .ZN(n4740) );
  NAND2_X1 U5123 ( .A1(n4769), .A2(n4741), .ZN(n4666) );
  NAND2_X1 U5124 ( .A1(n4707), .A2(n4730), .ZN(n4667) );
  INV_X1 U5125 ( .A(n4730), .ZN(n4668) );
  NOR2_X1 U5126 ( .A1(n4722), .A2(n4713), .ZN(n4670) );
  AOI21_X1 U5127 ( .B1(n4706), .B2(n4709), .A(n4670), .ZN(n4671) );
  XNOR2_X1 U5128 ( .A(n4671), .B(n4688), .ZN(n4898) );
  NAND2_X1 U5129 ( .A1(n4898), .A2(n5268), .ZN(n4705) );
  AOI22_X1 U5130 ( .A1(n5301), .A2(REG2_REG_29__SCAN_IN), .B1(n4672), .B2(
        n5097), .ZN(n4704) );
  INV_X1 U5131 ( .A(n4673), .ZN(n4674) );
  INV_X1 U5132 ( .A(n4675), .ZN(n4858) );
  INV_X1 U5133 ( .A(n4681), .ZN(n4682) );
  NOR2_X1 U5134 ( .A1(n4708), .A2(n4686), .ZN(n4687) );
  XOR2_X1 U5135 ( .A(n4688), .B(n4687), .Z(n4694) );
  INV_X1 U5136 ( .A(B_REG_SCAN_IN), .ZN(n4689) );
  NOR2_X1 U5137 ( .A1(n4989), .A2(n4689), .ZN(n4690) );
  NOR2_X1 U5138 ( .A1(n5048), .A2(n4690), .ZN(n5280) );
  OAI22_X1 U5139 ( .A1(n4722), .A2(n4887), .B1(n4698), .B2(n5283), .ZN(n4691)
         );
  AOI21_X1 U5140 ( .B1(n5280), .B2(n4692), .A(n4691), .ZN(n4693) );
  OAI21_X1 U5141 ( .B1(n4694), .B2(n4860), .A(n4693), .ZN(n4900) );
  NAND2_X1 U5142 ( .A1(n4900), .A2(n5258), .ZN(n4703) );
  INV_X1 U5143 ( .A(n4715), .ZN(n4700) );
  AOI21_X1 U5144 ( .B1(n4700), .B2(n4699), .A(n5273), .ZN(n4701) );
  AND2_X1 U5145 ( .A1(n5296), .A2(n4701), .ZN(n4899) );
  NAND2_X1 U5146 ( .A1(n4899), .A2(n4818), .ZN(n4702) );
  NAND4_X1 U5147 ( .A1(n4705), .A2(n4704), .A3(n4703), .A4(n4702), .ZN(U3354)
         );
  XNOR2_X1 U5148 ( .A(n4706), .B(n4709), .ZN(n4911) );
  OAI22_X1 U5149 ( .A1(n4707), .A2(n4887), .B1(n4713), .B2(n5283), .ZN(n4711)
         );
  INV_X1 U5150 ( .A(n4910), .ZN(n4719) );
  OAI21_X1 U5151 ( .B1(n4732), .B2(n4713), .A(n5303), .ZN(n4714) );
  OR2_X1 U5152 ( .A1(n4715), .A2(n4714), .ZN(n4909) );
  AOI22_X1 U5153 ( .A1(n5301), .A2(REG2_REG_28__SCAN_IN), .B1(n4716), .B2(
        n5097), .ZN(n4717) );
  OAI21_X1 U5154 ( .B1(n4909), .B2(n4872), .A(n4717), .ZN(n4718) );
  AOI21_X1 U5155 ( .B1(n4719), .B2(n5258), .A(n4718), .ZN(n4720) );
  OAI21_X1 U5156 ( .B1(n4911), .B2(n4876), .A(n4720), .ZN(U3262) );
  XOR2_X1 U5157 ( .A(n4724), .B(n4721), .Z(n4912) );
  OAI22_X1 U5158 ( .A1(n4722), .A2(n5048), .B1(n5283), .B2(n4730), .ZN(n4728)
         );
  AOI21_X1 U5159 ( .B1(n4725), .B2(n4724), .A(n4723), .ZN(n4726) );
  NOR2_X1 U5160 ( .A1(n4726), .A2(n4860), .ZN(n4727) );
  AOI211_X1 U5161 ( .C1(n4866), .C2(n4769), .A(n4728), .B(n4727), .ZN(n4913)
         );
  NOR2_X1 U5162 ( .A1(n4913), .A2(n5301), .ZN(n4736) );
  NOR2_X1 U5163 ( .A1(n4729), .A2(n4730), .ZN(n4731) );
  OR2_X1 U5164 ( .A1(n4732), .A2(n4731), .ZN(n4915) );
  AOI22_X1 U5165 ( .A1(n5301), .A2(REG2_REG_27__SCAN_IN), .B1(n4733), .B2(
        n5097), .ZN(n4734) );
  OAI21_X1 U5166 ( .B1(n4915), .B2(n4897), .A(n4734), .ZN(n4735) );
  AOI211_X1 U5167 ( .C1(n4912), .C2(n5268), .A(n4736), .B(n4735), .ZN(n4737)
         );
  INV_X1 U5168 ( .A(n4737), .ZN(U3263) );
  OAI21_X1 U5169 ( .B1(n4740), .B2(n4739), .A(n4738), .ZN(n4919) );
  AND2_X1 U5170 ( .A1(n4921), .A2(n4741), .ZN(n4742) );
  NOR2_X1 U5171 ( .A1(n4729), .A2(n4742), .ZN(n4916) );
  INV_X1 U5172 ( .A(REG2_REG_26__SCAN_IN), .ZN(n4744) );
  OAI22_X1 U5173 ( .A1(n5258), .A2(n4744), .B1(n4743), .B2(n5260), .ZN(n4745)
         );
  AOI21_X1 U5174 ( .B1(n4916), .B2(n5298), .A(n4745), .ZN(n4757) );
  INV_X1 U5175 ( .A(n4746), .ZN(n4747) );
  XNOR2_X1 U5176 ( .A(n4750), .B(n4749), .ZN(n4755) );
  INV_X1 U5177 ( .A(n4751), .ZN(n4752) );
  OAI21_X1 U5178 ( .B1(n4753), .B2(n5283), .A(n4752), .ZN(n4754) );
  AOI21_X1 U5179 ( .B1(n4755), .B2(n5256), .A(n4754), .ZN(n4918) );
  OR2_X1 U5180 ( .A1(n4918), .A2(n5301), .ZN(n4756) );
  OAI211_X1 U5181 ( .C1(n4919), .C2(n4876), .A(n4757), .B(n4756), .ZN(U3264)
         );
  OAI21_X1 U5182 ( .B1(n4759), .B2(n4767), .A(n4758), .ZN(n4924) );
  NAND2_X1 U5183 ( .A1(n4785), .A2(n4760), .ZN(n4920) );
  AND2_X1 U5184 ( .A1(n4920), .A2(n5298), .ZN(n4764) );
  INV_X1 U5185 ( .A(REG2_REG_25__SCAN_IN), .ZN(n4762) );
  OAI22_X1 U5186 ( .A1(n5258), .A2(n4762), .B1(n4761), .B2(n5260), .ZN(n4763)
         );
  AOI21_X1 U5187 ( .B1(n4764), .B2(n4921), .A(n4763), .ZN(n4776) );
  NAND2_X1 U5188 ( .A1(n4766), .A2(n4765), .ZN(n4768) );
  XNOR2_X1 U5189 ( .A(n4768), .B(n4767), .ZN(n4774) );
  NAND2_X1 U5190 ( .A1(n4769), .A2(n4839), .ZN(n4771) );
  NAND2_X1 U5191 ( .A1(n4799), .A2(n4866), .ZN(n4770) );
  OAI211_X1 U5192 ( .C1(n5283), .C2(n4772), .A(n4771), .B(n4770), .ZN(n4773)
         );
  AOI21_X1 U5193 ( .B1(n4774), .B2(n5256), .A(n4773), .ZN(n4923) );
  OR2_X1 U5194 ( .A1(n4923), .A2(n5301), .ZN(n4775) );
  OAI211_X1 U5195 ( .C1(n4924), .C2(n4876), .A(n4776), .B(n4775), .ZN(U3265)
         );
  XNOR2_X1 U5196 ( .A(n4777), .B(n4778), .ZN(n4927) );
  XNOR2_X1 U5197 ( .A(n4779), .B(n4778), .ZN(n4783) );
  AOI22_X1 U5198 ( .A1(n4824), .A2(n4866), .B1(n5292), .B2(n4784), .ZN(n4780)
         );
  OAI21_X1 U5199 ( .B1(n4781), .B2(n5048), .A(n4780), .ZN(n4782) );
  AOI21_X1 U5200 ( .B1(n4783), .B2(n5256), .A(n4782), .ZN(n4926) );
  INV_X1 U5201 ( .A(n4926), .ZN(n4790) );
  AOI21_X1 U5202 ( .B1(n4793), .B2(n4784), .A(n5273), .ZN(n4786) );
  NAND2_X1 U5203 ( .A1(n4786), .A2(n4785), .ZN(n4925) );
  AOI22_X1 U5204 ( .A1(n5301), .A2(REG2_REG_24__SCAN_IN), .B1(n4787), .B2(
        n5097), .ZN(n4788) );
  OAI21_X1 U5205 ( .B1(n4925), .B2(n4872), .A(n4788), .ZN(n4789) );
  AOI21_X1 U5206 ( .B1(n4790), .B2(n5258), .A(n4789), .ZN(n4791) );
  OAI21_X1 U5207 ( .B1(n4927), .B2(n4876), .A(n4791), .ZN(U3266) );
  XOR2_X1 U5208 ( .A(n4798), .B(n4792), .Z(n4930) );
  OAI211_X1 U5209 ( .C1(n4812), .C2(n4802), .A(n5303), .B(n4793), .ZN(n4928)
         );
  INV_X1 U5210 ( .A(n4928), .ZN(n4808) );
  NOR2_X1 U5211 ( .A1(n4834), .A2(n4836), .ZN(n4796) );
  INV_X1 U5212 ( .A(n4794), .ZN(n4795) );
  AOI21_X1 U5213 ( .B1(n4862), .B2(n4796), .A(n4795), .ZN(n4821) );
  AND2_X1 U5214 ( .A1(n4821), .A2(n4820), .ZN(n4823) );
  XNOR2_X1 U5215 ( .A(n4798), .B(n2704), .ZN(n4804) );
  NAND2_X1 U5216 ( .A1(n4799), .A2(n4839), .ZN(n4801) );
  NAND2_X1 U5217 ( .A1(n4840), .A2(n4866), .ZN(n4800) );
  OAI211_X1 U5218 ( .C1(n5283), .C2(n4802), .A(n4801), .B(n4800), .ZN(n4803)
         );
  AOI21_X1 U5219 ( .B1(n4804), .B2(n5256), .A(n4803), .ZN(n4929) );
  AOI22_X1 U5220 ( .A1(n5301), .A2(REG2_REG_23__SCAN_IN), .B1(n4805), .B2(
        n5097), .ZN(n4806) );
  OAI21_X1 U5221 ( .B1(n4929), .B2(n5301), .A(n4806), .ZN(n4807) );
  AOI21_X1 U5222 ( .B1(n4808), .B2(n4818), .A(n4807), .ZN(n4809) );
  OAI21_X1 U5223 ( .B1(n4930), .B2(n4876), .A(n4809), .ZN(U3267) );
  OAI21_X1 U5224 ( .B1(n2490), .B2(n4811), .A(n4810), .ZN(n4933) );
  OAI21_X1 U5225 ( .B1(n4845), .B2(n4828), .A(n5303), .ZN(n4813) );
  OR2_X1 U5226 ( .A1(n4813), .A2(n4812), .ZN(n4931) );
  INV_X1 U5227 ( .A(n4931), .ZN(n4819) );
  INV_X1 U5228 ( .A(REG2_REG_22__SCAN_IN), .ZN(n4816) );
  INV_X1 U5229 ( .A(n4814), .ZN(n4815) );
  OAI22_X1 U5230 ( .A1(n5258), .A2(n4816), .B1(n4815), .B2(n5260), .ZN(n4817)
         );
  AOI21_X1 U5231 ( .B1(n4819), .B2(n4818), .A(n4817), .ZN(n4832) );
  NOR2_X1 U5232 ( .A1(n4821), .A2(n4820), .ZN(n4822) );
  OR2_X1 U5233 ( .A1(n4823), .A2(n4822), .ZN(n4830) );
  NAND2_X1 U5234 ( .A1(n4824), .A2(n4839), .ZN(n4827) );
  NAND2_X1 U5235 ( .A1(n4825), .A2(n4866), .ZN(n4826) );
  OAI211_X1 U5236 ( .C1(n5283), .C2(n4828), .A(n4827), .B(n4826), .ZN(n4829)
         );
  AOI21_X1 U5237 ( .B1(n4830), .B2(n5256), .A(n4829), .ZN(n4932) );
  OR2_X1 U5238 ( .A1(n4932), .A2(n5301), .ZN(n4831) );
  OAI211_X1 U5239 ( .C1(n4933), .C2(n4876), .A(n4832), .B(n4831), .ZN(U3268)
         );
  XNOR2_X1 U5240 ( .A(n4833), .B(n4836), .ZN(n4936) );
  INV_X1 U5241 ( .A(n4862), .ZN(n4835) );
  NOR2_X1 U5242 ( .A1(n4835), .A2(n4834), .ZN(n4837) );
  XNOR2_X1 U5243 ( .A(n4837), .B(n4836), .ZN(n4844) );
  NAND2_X1 U5244 ( .A1(n4838), .A2(n4866), .ZN(n4842) );
  NAND2_X1 U5245 ( .A1(n4840), .A2(n4839), .ZN(n4841) );
  OAI211_X1 U5246 ( .C1(n5283), .C2(n4847), .A(n4842), .B(n4841), .ZN(n4843)
         );
  AOI21_X1 U5247 ( .B1(n4844), .B2(n5256), .A(n4843), .ZN(n4935) );
  INV_X1 U5248 ( .A(n4935), .ZN(n4852) );
  INV_X1 U5249 ( .A(n4867), .ZN(n4848) );
  INV_X1 U5250 ( .A(n4845), .ZN(n4846) );
  OAI211_X1 U5251 ( .C1(n4848), .C2(n4847), .A(n4846), .B(n5303), .ZN(n4934)
         );
  AOI22_X1 U5252 ( .A1(n5301), .A2(REG2_REG_21__SCAN_IN), .B1(n4849), .B2(
        n5097), .ZN(n4850) );
  OAI21_X1 U5253 ( .B1(n4934), .B2(n4872), .A(n4850), .ZN(n4851) );
  AOI21_X1 U5254 ( .B1(n4852), .B2(n5258), .A(n4851), .ZN(n4853) );
  OAI21_X1 U5255 ( .B1(n4936), .B2(n4876), .A(n4853), .ZN(U3269) );
  XOR2_X1 U5256 ( .A(n4856), .B(n4854), .Z(n4939) );
  OAI22_X1 U5257 ( .A1(n4855), .A2(n5048), .B1(n5283), .B2(n4868), .ZN(n4864)
         );
  INV_X1 U5258 ( .A(n4856), .ZN(n4857) );
  NAND3_X1 U5259 ( .A1(n4859), .A2(n4858), .A3(n4857), .ZN(n4861) );
  AOI21_X1 U5260 ( .B1(n4862), .B2(n4861), .A(n4860), .ZN(n4863) );
  AOI211_X1 U5261 ( .C1(n4866), .C2(n4865), .A(n4864), .B(n4863), .ZN(n4938)
         );
  INV_X1 U5262 ( .A(n4938), .ZN(n4874) );
  INV_X1 U5263 ( .A(n5265), .ZN(n4869) );
  OAI211_X1 U5264 ( .C1(n4869), .C2(n4868), .A(n5303), .B(n4867), .ZN(n4937)
         );
  AOI22_X1 U5265 ( .A1(n5301), .A2(REG2_REG_20__SCAN_IN), .B1(n4870), .B2(
        n5097), .ZN(n4871) );
  OAI21_X1 U5266 ( .B1(n4937), .B2(n4872), .A(n4871), .ZN(n4873) );
  AOI21_X1 U5267 ( .B1(n4874), .B2(n5258), .A(n4873), .ZN(n4875) );
  OAI21_X1 U5268 ( .B1(n4939), .B2(n4876), .A(n4875), .ZN(U3270) );
  NAND2_X1 U5269 ( .A1(n4877), .A2(n5217), .ZN(n4878) );
  NAND2_X1 U5270 ( .A1(n4879), .A2(n4878), .ZN(n5223) );
  XNOR2_X1 U5271 ( .A(n4880), .B(n4883), .ZN(n5225) );
  NAND2_X1 U5272 ( .A1(n5225), .A2(n5268), .ZN(n4896) );
  NAND2_X1 U5273 ( .A1(n4882), .A2(n4881), .ZN(n4884) );
  XNOR2_X1 U5274 ( .A(n4884), .B(n4883), .ZN(n4892) );
  NOR2_X1 U5275 ( .A1(n4885), .A2(n5283), .ZN(n4891) );
  OR2_X1 U5276 ( .A1(n4886), .A2(n5048), .ZN(n4890) );
  OR2_X1 U5277 ( .A1(n4888), .A2(n4887), .ZN(n4889) );
  NAND2_X1 U5278 ( .A1(n4890), .A2(n4889), .ZN(n5214) );
  AOI211_X1 U5279 ( .C1(n4892), .C2(n5256), .A(n4891), .B(n5214), .ZN(n5222)
         );
  OAI21_X1 U5280 ( .B1(n5221), .B2(n5260), .A(n5222), .ZN(n4894) );
  NOR2_X1 U5281 ( .A1(n5258), .A2(n2853), .ZN(n4893) );
  AOI21_X1 U5282 ( .B1(n4894), .B2(n5258), .A(n4893), .ZN(n4895) );
  OAI211_X1 U5283 ( .C1(n5223), .C2(n4897), .A(n4896), .B(n4895), .ZN(U3273)
         );
  OR2_X1 U5284 ( .A1(n5056), .A2(n2576), .ZN(n5046) );
  NAND2_X1 U5285 ( .A1(n4898), .A2(n5275), .ZN(n4902) );
  NAND2_X1 U5286 ( .A1(n4902), .A2(n4901), .ZN(n4942) );
  NOR2_X1 U5287 ( .A1(n4907), .A2(n4906), .ZN(n4908) );
  AND2_X2 U5288 ( .A1(n4941), .A2(n4908), .ZN(n5307) );
  MUX2_X1 U5289 ( .A(REG1_REG_29__SCAN_IN), .B(n4942), .S(n5307), .Z(U3547) );
  OAI211_X1 U5290 ( .C1(n4911), .C2(n5202), .A(n4910), .B(n4909), .ZN(n4943)
         );
  MUX2_X1 U5291 ( .A(REG1_REG_28__SCAN_IN), .B(n4943), .S(n5307), .Z(U3546) );
  NAND2_X1 U5292 ( .A1(n4912), .A2(n5275), .ZN(n4914) );
  OAI211_X1 U5293 ( .C1(n5273), .C2(n4915), .A(n4914), .B(n4913), .ZN(n4944)
         );
  MUX2_X1 U5294 ( .A(REG1_REG_27__SCAN_IN), .B(n4944), .S(n5307), .Z(U3545) );
  NAND2_X1 U5295 ( .A1(n4916), .A2(n5303), .ZN(n4917) );
  OAI211_X1 U5296 ( .C1(n4919), .C2(n5202), .A(n4918), .B(n4917), .ZN(n4945)
         );
  MUX2_X1 U5297 ( .A(REG1_REG_26__SCAN_IN), .B(n4945), .S(n5307), .Z(U3544) );
  NAND3_X1 U5298 ( .A1(n4921), .A2(n5303), .A3(n4920), .ZN(n4922) );
  OAI211_X1 U5299 ( .C1(n4924), .C2(n5202), .A(n4923), .B(n4922), .ZN(n4946)
         );
  MUX2_X1 U5300 ( .A(REG1_REG_25__SCAN_IN), .B(n4946), .S(n5307), .Z(U3543) );
  OAI211_X1 U5301 ( .C1(n4927), .C2(n5202), .A(n4926), .B(n4925), .ZN(n4947)
         );
  MUX2_X1 U5302 ( .A(REG1_REG_24__SCAN_IN), .B(n4947), .S(n5307), .Z(U3542) );
  OAI211_X1 U5303 ( .C1(n4930), .C2(n5202), .A(n4929), .B(n4928), .ZN(n4948)
         );
  MUX2_X1 U5304 ( .A(REG1_REG_23__SCAN_IN), .B(n4948), .S(n5307), .Z(U3541) );
  OAI211_X1 U5305 ( .C1(n4933), .C2(n5202), .A(n4932), .B(n4931), .ZN(n4949)
         );
  MUX2_X1 U5306 ( .A(REG1_REG_22__SCAN_IN), .B(n4949), .S(n5307), .Z(U3540) );
  OAI211_X1 U5307 ( .C1(n4936), .C2(n5202), .A(n4935), .B(n4934), .ZN(n4950)
         );
  MUX2_X1 U5308 ( .A(REG1_REG_21__SCAN_IN), .B(n4950), .S(n5307), .Z(U3539) );
  OAI211_X1 U5309 ( .C1(n4939), .C2(n5202), .A(n4938), .B(n4937), .ZN(n4951)
         );
  MUX2_X1 U5310 ( .A(REG1_REG_20__SCAN_IN), .B(n4951), .S(n5307), .Z(U3538) );
  AND2_X2 U5311 ( .A1(n4941), .A2(n4940), .ZN(n5311) );
  MUX2_X1 U5312 ( .A(REG0_REG_29__SCAN_IN), .B(n4942), .S(n5311), .Z(U3515) );
  MUX2_X1 U5313 ( .A(REG0_REG_28__SCAN_IN), .B(n4943), .S(n5311), .Z(U3514) );
  MUX2_X1 U5314 ( .A(REG0_REG_27__SCAN_IN), .B(n4944), .S(n5311), .Z(U3513) );
  MUX2_X1 U5315 ( .A(REG0_REG_26__SCAN_IN), .B(n4945), .S(n5311), .Z(U3512) );
  MUX2_X1 U5316 ( .A(REG0_REG_25__SCAN_IN), .B(n4946), .S(n5311), .Z(U3511) );
  MUX2_X1 U5317 ( .A(REG0_REG_24__SCAN_IN), .B(n4947), .S(n5311), .Z(U3510) );
  MUX2_X1 U5318 ( .A(REG0_REG_23__SCAN_IN), .B(n4948), .S(n5311), .Z(U3509) );
  MUX2_X1 U5319 ( .A(REG0_REG_22__SCAN_IN), .B(n4949), .S(n5311), .Z(U3508) );
  MUX2_X1 U5320 ( .A(REG0_REG_21__SCAN_IN), .B(n4950), .S(n5311), .Z(U3507) );
  MUX2_X1 U5321 ( .A(REG0_REG_20__SCAN_IN), .B(n4951), .S(n5311), .Z(U3506) );
  MUX2_X1 U5322 ( .A(n4952), .B(D_REG_1__SCAN_IN), .S(n4988), .Z(U3459) );
  NOR3_X1 U5323 ( .A1(n2921), .A2(IR_REG_30__SCAN_IN), .A3(n2810), .ZN(n4953)
         );
  MUX2_X1 U5324 ( .A(DATAI_31_), .B(n4953), .S(STATE_REG_SCAN_IN), .Z(U3321)
         );
  MUX2_X1 U5325 ( .A(n4954), .B(DATAI_29_), .S(U3149), .Z(U3323) );
  MUX2_X1 U5326 ( .A(n5013), .B(DATAI_27_), .S(U3149), .Z(U3325) );
  MUX2_X1 U5327 ( .A(n4955), .B(DATAI_25_), .S(U3149), .Z(U3327) );
  MUX2_X1 U5328 ( .A(DATAI_24_), .B(n4956), .S(STATE_REG_SCAN_IN), .Z(U3328)
         );
  MUX2_X1 U5329 ( .A(n4957), .B(DATAI_21_), .S(U3149), .Z(U3331) );
  MUX2_X1 U5330 ( .A(n4958), .B(DATAI_20_), .S(U3149), .Z(U3332) );
  MUX2_X1 U5331 ( .A(n4959), .B(DATAI_19_), .S(U3149), .Z(U3333) );
  MUX2_X1 U5332 ( .A(DATAI_17_), .B(n4960), .S(STATE_REG_SCAN_IN), .Z(U3335)
         );
  MUX2_X1 U5333 ( .A(DATAI_16_), .B(n4961), .S(STATE_REG_SCAN_IN), .Z(U3336)
         );
  MUX2_X1 U5334 ( .A(DATAI_15_), .B(n4962), .S(STATE_REG_SCAN_IN), .Z(U3337)
         );
  MUX2_X1 U5335 ( .A(DATAI_14_), .B(n4963), .S(STATE_REG_SCAN_IN), .Z(U3338)
         );
  MUX2_X1 U5336 ( .A(n4964), .B(DATAI_13_), .S(U3149), .Z(U3339) );
  MUX2_X1 U5337 ( .A(DATAI_12_), .B(n4965), .S(STATE_REG_SCAN_IN), .Z(U3340)
         );
  MUX2_X1 U5338 ( .A(n4966), .B(DATAI_11_), .S(U3149), .Z(U3341) );
  MUX2_X1 U5339 ( .A(n4967), .B(DATAI_6_), .S(U3149), .Z(U3346) );
  MUX2_X1 U5340 ( .A(n4968), .B(DATAI_5_), .S(U3149), .Z(U3347) );
  MUX2_X1 U5341 ( .A(n5022), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  MUX2_X1 U5342 ( .A(n2467), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  MUX2_X1 U5343 ( .A(DATAI_0_), .B(IR_REG_0__SCAN_IN), .S(STATE_REG_SCAN_IN), 
        .Z(U3352) );
  OAI21_X1 U5344 ( .B1(STATE_REG_SCAN_IN), .B2(DATAI_23_), .A(n4970), .ZN(
        n4971) );
  INV_X1 U5345 ( .A(n4971), .ZN(U3329) );
  NOR2_X1 U5346 ( .A1(n4987), .A2(n4972), .ZN(U3320) );
  NOR2_X1 U5347 ( .A1(n4987), .A2(n4973), .ZN(U3319) );
  AND2_X1 U5348 ( .A1(n4988), .A2(D_REG_4__SCAN_IN), .ZN(U3318) );
  AND2_X1 U5349 ( .A1(n4988), .A2(D_REG_5__SCAN_IN), .ZN(U3317) );
  NOR2_X1 U5350 ( .A1(n4987), .A2(n4974), .ZN(U3316) );
  NOR2_X1 U5351 ( .A1(n4987), .A2(n4975), .ZN(U3315) );
  NOR2_X1 U5352 ( .A1(n4987), .A2(n4316), .ZN(U3314) );
  NOR2_X1 U5353 ( .A1(n4987), .A2(n4976), .ZN(U3313) );
  NOR2_X1 U5354 ( .A1(n4987), .A2(n4977), .ZN(U3312) );
  NOR2_X1 U5355 ( .A1(n4987), .A2(n4978), .ZN(U3311) );
  AND2_X1 U5356 ( .A1(n4988), .A2(D_REG_12__SCAN_IN), .ZN(U3310) );
  AND2_X1 U5357 ( .A1(n4988), .A2(D_REG_13__SCAN_IN), .ZN(U3309) );
  NOR2_X1 U5358 ( .A1(n4987), .A2(n4979), .ZN(U3308) );
  AND2_X1 U5359 ( .A1(n4988), .A2(D_REG_15__SCAN_IN), .ZN(U3307) );
  AND2_X1 U5360 ( .A1(n4988), .A2(D_REG_16__SCAN_IN), .ZN(U3306) );
  NOR2_X1 U5361 ( .A1(n4987), .A2(n4980), .ZN(U3305) );
  AND2_X1 U5362 ( .A1(n4988), .A2(D_REG_18__SCAN_IN), .ZN(U3304) );
  AND2_X1 U5363 ( .A1(n4988), .A2(D_REG_19__SCAN_IN), .ZN(U3303) );
  INV_X1 U5364 ( .A(D_REG_20__SCAN_IN), .ZN(n4981) );
  NOR2_X1 U5365 ( .A1(n4987), .A2(n4981), .ZN(U3302) );
  AND2_X1 U5366 ( .A1(n4988), .A2(D_REG_21__SCAN_IN), .ZN(U3301) );
  NOR2_X1 U5367 ( .A1(n4987), .A2(n4982), .ZN(U3300) );
  AND2_X1 U5368 ( .A1(n4988), .A2(D_REG_23__SCAN_IN), .ZN(U3299) );
  NOR2_X1 U5369 ( .A1(n4987), .A2(n4983), .ZN(U3298) );
  AND2_X1 U5370 ( .A1(n4988), .A2(D_REG_25__SCAN_IN), .ZN(U3297) );
  NOR2_X1 U5371 ( .A1(n4987), .A2(n4984), .ZN(U3296) );
  AND2_X1 U5372 ( .A1(n4988), .A2(D_REG_27__SCAN_IN), .ZN(U3295) );
  AND2_X1 U5373 ( .A1(n4988), .A2(D_REG_28__SCAN_IN), .ZN(U3294) );
  NOR2_X1 U5374 ( .A1(n4987), .A2(n4985), .ZN(U3293) );
  NOR2_X1 U5375 ( .A1(n4987), .A2(n4986), .ZN(U3292) );
  AND2_X1 U5376 ( .A1(n4988), .A2(D_REG_31__SCAN_IN), .ZN(U3291) );
  NOR2_X1 U5377 ( .A1(n4989), .A2(REG2_REG_0__SCAN_IN), .ZN(n4990) );
  OR2_X1 U5378 ( .A1(n2855), .A2(n4990), .ZN(n5018) );
  INV_X1 U5379 ( .A(n5018), .ZN(n4991) );
  OAI21_X1 U5380 ( .B1(n5013), .B2(REG1_REG_0__SCAN_IN), .A(n4991), .ZN(n4992)
         );
  XNOR2_X1 U5381 ( .A(n4992), .B(IR_REG_0__SCAN_IN), .ZN(n4994) );
  AOI22_X1 U5382 ( .A1(n5003), .A2(ADDR_REG_0__SCAN_IN), .B1(n4994), .B2(n4993), .ZN(n4995) );
  OAI21_X1 U5383 ( .B1(STATE_REG_SCAN_IN), .B2(n4996), .A(n4995), .ZN(U3240)
         );
  AOI21_X1 U5384 ( .B1(REG2_REG_18__SCAN_IN), .B2(n5001), .A(n4997), .ZN(n4999) );
  INV_X1 U5385 ( .A(REG2_REG_19__SCAN_IN), .ZN(n5259) );
  MUX2_X1 U5386 ( .A(REG2_REG_19__SCAN_IN), .B(n5259), .S(n5006), .Z(n4998) );
  XNOR2_X1 U5387 ( .A(n4999), .B(n4998), .ZN(n5010) );
  INV_X1 U5388 ( .A(REG1_REG_19__SCAN_IN), .ZN(n5277) );
  MUX2_X1 U5389 ( .A(REG1_REG_19__SCAN_IN), .B(n5277), .S(n5006), .Z(n5002) );
  NAND2_X1 U5390 ( .A1(n5003), .A2(ADDR_REG_19__SCAN_IN), .ZN(n5005) );
  OAI211_X1 U5391 ( .C1(n5042), .C2(n5006), .A(n5005), .B(n5004), .ZN(n5007)
         );
  AOI21_X1 U5392 ( .B1(n5008), .B2(n5038), .A(n5007), .ZN(n5009) );
  OAI21_X1 U5393 ( .B1(n5010), .B2(n5031), .A(n5009), .ZN(U3259) );
  NOR2_X1 U5394 ( .A1(n5011), .A2(n2855), .ZN(n5015) );
  NOR2_X1 U5395 ( .A1(n2855), .A2(n5012), .ZN(n5014) );
  MUX2_X1 U5396 ( .A(n5015), .B(n5014), .S(n5013), .Z(n5016) );
  AOI211_X1 U5397 ( .C1(n2571), .C2(n5018), .A(n5017), .B(n5016), .ZN(n5045)
         );
  AOI211_X1 U5398 ( .C1(n5021), .C2(n5020), .A(n5019), .B(n5031), .ZN(n5030)
         );
  INV_X1 U5399 ( .A(n5022), .ZN(n5028) );
  AOI22_X1 U5400 ( .A1(n5036), .A2(ADDR_REG_2__SCAN_IN), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n5027) );
  OAI211_X1 U5401 ( .C1(n5025), .C2(n5024), .A(n5038), .B(n5023), .ZN(n5026)
         );
  OAI211_X1 U5402 ( .C1(n5042), .C2(n5028), .A(n5027), .B(n5026), .ZN(n5029)
         );
  OR3_X1 U5403 ( .A1(n5045), .A2(n5030), .A3(n5029), .ZN(U3242) );
  AOI211_X1 U5404 ( .C1(n5034), .C2(n5033), .A(n5032), .B(n5031), .ZN(n5044)
         );
  AOI21_X1 U5405 ( .B1(n5036), .B2(ADDR_REG_4__SCAN_IN), .A(n5035), .ZN(n5041)
         );
  OAI211_X1 U5406 ( .C1(REG1_REG_4__SCAN_IN), .C2(n5039), .A(n5038), .B(n5037), 
        .ZN(n5040) );
  OAI211_X1 U5407 ( .C1(n5042), .C2(n5105), .A(n5041), .B(n5040), .ZN(n5043)
         );
  OR3_X1 U5408 ( .A1(n5045), .A2(n5044), .A3(n5043), .ZN(U3244) );
  INV_X1 U5409 ( .A(n5046), .ZN(n5091) );
  INV_X1 U5410 ( .A(n5051), .ZN(n5058) );
  NOR2_X1 U5411 ( .A1(n2563), .A2(n5047), .ZN(n5057) );
  NOR2_X1 U5412 ( .A1(n5086), .A2(n5256), .ZN(n5050) );
  OAI22_X1 U5413 ( .A1(n5051), .A2(n5050), .B1(n5049), .B2(n5048), .ZN(n5055)
         );
  AOI211_X1 U5414 ( .C1(n5091), .C2(n5058), .A(n5057), .B(n5055), .ZN(n5054)
         );
  AOI22_X1 U5415 ( .A1(n5307), .A2(n5054), .B1(n5052), .B2(n5305), .ZN(U3518)
         );
  AOI22_X1 U5416 ( .A1(n5311), .A2(n5054), .B1(n5053), .B2(n5308), .ZN(U3467)
         );
  AOI21_X1 U5417 ( .B1(n5057), .B2(n5056), .A(n5055), .ZN(n5061) );
  INV_X1 U5418 ( .A(REG2_REG_0__SCAN_IN), .ZN(n5060) );
  AOI22_X1 U5419 ( .A1(n5058), .A2(n5099), .B1(REG3_REG_0__SCAN_IN), .B2(n5097), .ZN(n5059) );
  OAI221_X1 U5420 ( .B1(n5301), .B2(n5061), .C1(n5258), .C2(n5060), .A(n5059), 
        .ZN(U3290) );
  INV_X1 U5421 ( .A(n5062), .ZN(n5065) );
  AOI211_X1 U5422 ( .C1(n5091), .C2(n5065), .A(n5064), .B(n5063), .ZN(n5067)
         );
  AOI22_X1 U5423 ( .A1(n5307), .A2(n5067), .B1(n2990), .B2(n5305), .ZN(U3519)
         );
  INV_X1 U5424 ( .A(REG0_REG_1__SCAN_IN), .ZN(n5066) );
  AOI22_X1 U5425 ( .A1(n5311), .A2(n5067), .B1(n5066), .B2(n5308), .ZN(U3469)
         );
  NOR2_X1 U5426 ( .A1(n5068), .A2(n5273), .ZN(n5070) );
  AOI211_X1 U5427 ( .C1(n5091), .C2(n5071), .A(n5070), .B(n5069), .ZN(n5073)
         );
  AOI22_X1 U5428 ( .A1(n5307), .A2(n5073), .B1(n2755), .B2(n5305), .ZN(U3520)
         );
  AOI22_X1 U5429 ( .A1(n5311), .A2(n5073), .B1(n5072), .B2(n5308), .ZN(U3471)
         );
  INV_X1 U5430 ( .A(DATAI_3_), .ZN(n5074) );
  AOI22_X1 U5431 ( .A1(STATE_REG_SCAN_IN), .A2(n5075), .B1(n5074), .B2(U3149), 
        .ZN(U3349) );
  XOR2_X1 U5432 ( .A(n5079), .B(n5076), .Z(n5100) );
  OAI21_X1 U5433 ( .B1(n5079), .B2(n5078), .A(n5077), .ZN(n5080) );
  NAND2_X1 U5434 ( .A1(n5080), .A2(n5256), .ZN(n5083) );
  INV_X1 U5435 ( .A(n5081), .ZN(n5082) );
  OAI211_X1 U5436 ( .C1(n5283), .C2(n5084), .A(n5083), .B(n5082), .ZN(n5085)
         );
  AOI21_X1 U5437 ( .B1(n5100), .B2(n5086), .A(n5085), .ZN(n5103) );
  INV_X1 U5438 ( .A(n5087), .ZN(n5088) );
  AOI21_X1 U5439 ( .B1(n5090), .B2(n5089), .A(n5088), .ZN(n5098) );
  AOI22_X1 U5440 ( .A1(n5100), .A2(n5091), .B1(n5303), .B2(n5098), .ZN(n5092)
         );
  AND2_X1 U5441 ( .A1(n5103), .A2(n5092), .ZN(n5095) );
  INV_X1 U5442 ( .A(REG1_REG_3__SCAN_IN), .ZN(n5093) );
  AOI22_X1 U5443 ( .A1(n5307), .A2(n5095), .B1(n5093), .B2(n5305), .ZN(U3521)
         );
  INV_X1 U5444 ( .A(REG0_REG_3__SCAN_IN), .ZN(n5094) );
  AOI22_X1 U5445 ( .A1(n5311), .A2(n5095), .B1(n5094), .B2(n5308), .ZN(U3473)
         );
  AOI22_X1 U5446 ( .A1(n5301), .A2(REG2_REG_3__SCAN_IN), .B1(n5097), .B2(n5096), .ZN(n5102) );
  AOI22_X1 U5447 ( .A1(n5100), .A2(n5099), .B1(n5298), .B2(n5098), .ZN(n5101)
         );
  OAI211_X1 U5448 ( .C1(n5301), .C2(n5103), .A(n5102), .B(n5101), .ZN(U3287)
         );
  AOI22_X1 U5449 ( .A1(STATE_REG_SCAN_IN), .A2(n5105), .B1(n5104), .B2(U3149), 
        .ZN(U3348) );
  NAND3_X1 U5450 ( .A1(n3245), .A2(n5106), .A3(n5275), .ZN(n5107) );
  AND3_X1 U5451 ( .A1(n5109), .A2(n5108), .A3(n5107), .ZN(n5112) );
  INV_X1 U5452 ( .A(REG1_REG_4__SCAN_IN), .ZN(n5110) );
  AOI22_X1 U5453 ( .A1(n5307), .A2(n5112), .B1(n5110), .B2(n5305), .ZN(U3522)
         );
  INV_X1 U5454 ( .A(REG0_REG_4__SCAN_IN), .ZN(n5111) );
  AOI22_X1 U5455 ( .A1(n5311), .A2(n5112), .B1(n5111), .B2(n5308), .ZN(U3475)
         );
  NOR2_X1 U5456 ( .A1(n5113), .A2(n5273), .ZN(n5115) );
  AOI211_X1 U5457 ( .C1(n5275), .C2(n5116), .A(n5115), .B(n5114), .ZN(n5119)
         );
  AOI22_X1 U5458 ( .A1(n5307), .A2(n5119), .B1(n5117), .B2(n5305), .ZN(U3523)
         );
  INV_X1 U5459 ( .A(REG0_REG_5__SCAN_IN), .ZN(n5118) );
  AOI22_X1 U5460 ( .A1(n5311), .A2(n5119), .B1(n5118), .B2(n5308), .ZN(U3477)
         );
  NOR2_X1 U5461 ( .A1(n5120), .A2(n5273), .ZN(n5122) );
  AOI211_X1 U5462 ( .C1(n5275), .C2(n5123), .A(n5122), .B(n5121), .ZN(n5125)
         );
  AOI22_X1 U5463 ( .A1(n5307), .A2(n5125), .B1(n2764), .B2(n5305), .ZN(U3524)
         );
  AOI22_X1 U5464 ( .A1(n5311), .A2(n5125), .B1(n5124), .B2(n5308), .ZN(U3479)
         );
  AOI22_X1 U5465 ( .A1(STATE_REG_SCAN_IN), .A2(n5127), .B1(n5126), .B2(U3149), 
        .ZN(U3345) );
  AOI211_X1 U5466 ( .C1(n5130), .C2(n5275), .A(n5129), .B(n5128), .ZN(n5132)
         );
  AOI22_X1 U5467 ( .A1(n5307), .A2(n5132), .B1(n2768), .B2(n5305), .ZN(U3525)
         );
  INV_X1 U5468 ( .A(REG0_REG_7__SCAN_IN), .ZN(n5131) );
  AOI22_X1 U5469 ( .A1(n5311), .A2(n5132), .B1(n5131), .B2(n5308), .ZN(U3481)
         );
  AOI22_X1 U5470 ( .A1(STATE_REG_SCAN_IN), .A2(n5134), .B1(n5133), .B2(U3149), 
        .ZN(U3344) );
  NOR2_X1 U5471 ( .A1(n5135), .A2(n5202), .ZN(n5136) );
  AOI211_X1 U5472 ( .C1(n5303), .C2(n5138), .A(n5137), .B(n5136), .ZN(n5141)
         );
  INV_X1 U5473 ( .A(REG1_REG_8__SCAN_IN), .ZN(n5139) );
  AOI22_X1 U5474 ( .A1(n5307), .A2(n5141), .B1(n5139), .B2(n5305), .ZN(U3526)
         );
  INV_X1 U5475 ( .A(REG0_REG_8__SCAN_IN), .ZN(n5140) );
  AOI22_X1 U5476 ( .A1(n5311), .A2(n5141), .B1(n5140), .B2(n5308), .ZN(U3483)
         );
  INV_X1 U5477 ( .A(DATAI_9_), .ZN(n5142) );
  AOI22_X1 U5478 ( .A1(STATE_REG_SCAN_IN), .A2(n5143), .B1(n5142), .B2(U3149), 
        .ZN(U3343) );
  OAI21_X1 U5479 ( .B1(n5273), .B2(n5145), .A(n5144), .ZN(n5146) );
  AOI21_X1 U5480 ( .B1(n5147), .B2(n5275), .A(n5146), .ZN(n5149) );
  AOI22_X1 U5481 ( .A1(n5307), .A2(n5149), .B1(n2739), .B2(n5305), .ZN(U3527)
         );
  INV_X1 U5482 ( .A(REG0_REG_9__SCAN_IN), .ZN(n5148) );
  AOI22_X1 U5483 ( .A1(n5311), .A2(n5149), .B1(n5148), .B2(n5308), .ZN(U3485)
         );
  AOI22_X1 U5484 ( .A1(STATE_REG_SCAN_IN), .A2(n5151), .B1(n5150), .B2(U3149), 
        .ZN(U3342) );
  NOR2_X1 U5485 ( .A1(n5152), .A2(n5273), .ZN(n5154) );
  AOI211_X1 U5486 ( .C1(n5155), .C2(n5275), .A(n5154), .B(n5153), .ZN(n5158)
         );
  INV_X1 U5487 ( .A(REG1_REG_10__SCAN_IN), .ZN(n5156) );
  AOI22_X1 U5488 ( .A1(n5307), .A2(n5158), .B1(n5156), .B2(n5305), .ZN(U3528)
         );
  INV_X1 U5489 ( .A(REG0_REG_10__SCAN_IN), .ZN(n5157) );
  AOI22_X1 U5490 ( .A1(n5311), .A2(n5158), .B1(n5157), .B2(n5308), .ZN(U3487)
         );
  OAI22_X1 U5491 ( .A1(n5160), .A2(n5202), .B1(n5159), .B2(n5273), .ZN(n5162)
         );
  NOR2_X1 U5492 ( .A1(n5162), .A2(n5161), .ZN(n5165) );
  AOI22_X1 U5493 ( .A1(n5307), .A2(n5165), .B1(n5163), .B2(n5305), .ZN(U3529)
         );
  INV_X1 U5494 ( .A(REG0_REG_11__SCAN_IN), .ZN(n5164) );
  AOI22_X1 U5495 ( .A1(n5311), .A2(n5165), .B1(n5164), .B2(n5308), .ZN(U3489)
         );
  INV_X1 U5496 ( .A(n5166), .ZN(n5167) );
  AOI211_X1 U5497 ( .C1(n5275), .C2(n5169), .A(n5168), .B(n5167), .ZN(n5172)
         );
  INV_X1 U5498 ( .A(REG1_REG_12__SCAN_IN), .ZN(n5170) );
  AOI22_X1 U5499 ( .A1(n5307), .A2(n5172), .B1(n5170), .B2(n5305), .ZN(U3530)
         );
  INV_X1 U5500 ( .A(REG0_REG_12__SCAN_IN), .ZN(n5171) );
  AOI22_X1 U5501 ( .A1(n5311), .A2(n5172), .B1(n5171), .B2(n5308), .ZN(U3491)
         );
  INV_X1 U5502 ( .A(n5173), .ZN(n5176) );
  INV_X1 U5503 ( .A(n5174), .ZN(n5175) );
  AOI21_X1 U5504 ( .B1(n5275), .B2(n5176), .A(n5175), .ZN(n5179) );
  INV_X1 U5505 ( .A(REG1_REG_13__SCAN_IN), .ZN(n5177) );
  AOI22_X1 U5506 ( .A1(n5307), .A2(n5179), .B1(n5177), .B2(n5305), .ZN(U3531)
         );
  INV_X1 U5507 ( .A(REG0_REG_13__SCAN_IN), .ZN(n5178) );
  AOI22_X1 U5508 ( .A1(n5311), .A2(n5179), .B1(n5178), .B2(n5308), .ZN(U3493)
         );
  OAI22_X1 U5509 ( .A1(n5181), .A2(n5202), .B1(n5180), .B2(n5273), .ZN(n5182)
         );
  NOR2_X1 U5510 ( .A1(n5183), .A2(n5182), .ZN(n5186) );
  INV_X1 U5511 ( .A(REG1_REG_14__SCAN_IN), .ZN(n5184) );
  AOI22_X1 U5512 ( .A1(n5307), .A2(n5186), .B1(n5184), .B2(n5305), .ZN(U3532)
         );
  INV_X1 U5513 ( .A(REG0_REG_14__SCAN_IN), .ZN(n5185) );
  AOI22_X1 U5514 ( .A1(n5311), .A2(n5186), .B1(n5185), .B2(n5308), .ZN(U3495)
         );
  AOI22_X1 U5515 ( .A1(n5231), .A2(n5187), .B1(REG3_REG_15__SCAN_IN), .B2(
        U3149), .ZN(n5198) );
  INV_X1 U5516 ( .A(n5188), .ZN(n5189) );
  NOR2_X1 U5517 ( .A1(n5189), .A2(n3598), .ZN(n5191) );
  OAI21_X1 U5518 ( .B1(n5191), .B2(n5193), .A(n5190), .ZN(n5196) );
  AOI21_X1 U5519 ( .B1(n3598), .B2(n5193), .A(n5192), .ZN(n5195) );
  AOI22_X1 U5520 ( .A1(n5196), .A2(n5195), .B1(n5194), .B2(n5237), .ZN(n5197)
         );
  OAI211_X1 U5521 ( .C1(n5244), .C2(n5199), .A(n5198), .B(n5197), .ZN(U3238)
         );
  OAI211_X1 U5522 ( .C1(n5203), .C2(n5202), .A(n5201), .B(n5200), .ZN(n5204)
         );
  INV_X1 U5523 ( .A(n5204), .ZN(n5207) );
  INV_X1 U5524 ( .A(REG1_REG_15__SCAN_IN), .ZN(n5205) );
  AOI22_X1 U5525 ( .A1(n5307), .A2(n5207), .B1(n5205), .B2(n5305), .ZN(U3533)
         );
  INV_X1 U5526 ( .A(REG0_REG_15__SCAN_IN), .ZN(n5206) );
  AOI22_X1 U5527 ( .A1(n5311), .A2(n5207), .B1(n5206), .B2(n5308), .ZN(U3497)
         );
  AOI211_X1 U5528 ( .C1(n5210), .C2(n5275), .A(n5209), .B(n5208), .ZN(n5213)
         );
  INV_X1 U5529 ( .A(REG1_REG_16__SCAN_IN), .ZN(n5211) );
  AOI22_X1 U5530 ( .A1(n5307), .A2(n5213), .B1(n5211), .B2(n5305), .ZN(U3534)
         );
  INV_X1 U5531 ( .A(REG0_REG_16__SCAN_IN), .ZN(n5212) );
  AOI22_X1 U5532 ( .A1(n5311), .A2(n5213), .B1(n5212), .B2(n5308), .ZN(U3499)
         );
  AOI22_X1 U5533 ( .A1(n5231), .A2(n5214), .B1(REG3_REG_17__SCAN_IN), .B2(
        U3149), .ZN(n5220) );
  XNOR2_X1 U5534 ( .A(n5216), .B(n5215), .ZN(n5218) );
  AOI22_X1 U5535 ( .A1(n5218), .A2(n5239), .B1(n5217), .B2(n5237), .ZN(n5219)
         );
  OAI211_X1 U5536 ( .C1(n5244), .C2(n5221), .A(n5220), .B(n5219), .ZN(U3225)
         );
  OAI21_X1 U5537 ( .B1(n5273), .B2(n5223), .A(n5222), .ZN(n5224) );
  AOI21_X1 U5538 ( .B1(n5225), .B2(n5275), .A(n5224), .ZN(n5227) );
  AOI22_X1 U5539 ( .A1(n5307), .A2(n5227), .B1(n2782), .B2(n5305), .ZN(U3535)
         );
  INV_X1 U5540 ( .A(REG0_REG_17__SCAN_IN), .ZN(n5226) );
  AOI22_X1 U5541 ( .A1(n5311), .A2(n5227), .B1(n5226), .B2(n5308), .ZN(U3501)
         );
  AOI22_X1 U5542 ( .A1(STATE_REG_SCAN_IN), .A2(n5229), .B1(n5228), .B2(U3149), 
        .ZN(U3334) );
  AOI22_X1 U5543 ( .A1(n5231), .A2(n5230), .B1(REG3_REG_18__SCAN_IN), .B2(
        U3149), .ZN(n5242) );
  INV_X1 U5544 ( .A(n5232), .ZN(n5234) );
  NAND2_X1 U5545 ( .A1(n5234), .A2(n5233), .ZN(n5235) );
  XNOR2_X1 U5546 ( .A(n5236), .B(n5235), .ZN(n5240) );
  AOI22_X1 U5547 ( .A1(n5240), .A2(n5239), .B1(n5238), .B2(n5237), .ZN(n5241)
         );
  OAI211_X1 U5548 ( .C1(n5244), .C2(n5243), .A(n5242), .B(n5241), .ZN(U3235)
         );
  AOI211_X1 U5549 ( .C1(n5247), .C2(n5275), .A(n5246), .B(n5245), .ZN(n5250)
         );
  AOI22_X1 U5550 ( .A1(n5307), .A2(n5250), .B1(n5248), .B2(n5305), .ZN(U3536)
         );
  INV_X1 U5551 ( .A(REG0_REG_18__SCAN_IN), .ZN(n5249) );
  AOI22_X1 U5552 ( .A1(n5311), .A2(n5250), .B1(n5249), .B2(n5308), .ZN(U3503)
         );
  NAND2_X1 U5553 ( .A1(n5252), .A2(n5251), .ZN(n5253) );
  XNOR2_X1 U5554 ( .A(n5253), .B(n5263), .ZN(n5257) );
  NOR2_X1 U5555 ( .A1(n5266), .A2(n5283), .ZN(n5255) );
  AOI211_X1 U5556 ( .C1(n5257), .C2(n5256), .A(n5255), .B(n5254), .ZN(n5271)
         );
  OAI22_X1 U5557 ( .A1(n5261), .A2(n5260), .B1(n5259), .B2(n5258), .ZN(n5262)
         );
  INV_X1 U5558 ( .A(n5262), .ZN(n5270) );
  XNOR2_X1 U5559 ( .A(n5264), .B(n5263), .ZN(n5276) );
  OAI21_X1 U5560 ( .B1(n4695), .B2(n5266), .A(n5265), .ZN(n5272) );
  INV_X1 U5561 ( .A(n5272), .ZN(n5267) );
  AOI22_X1 U5562 ( .A1(n5276), .A2(n5268), .B1(n5298), .B2(n5267), .ZN(n5269)
         );
  OAI211_X1 U5563 ( .C1(n5301), .C2(n5271), .A(n5270), .B(n5269), .ZN(U3271)
         );
  OAI21_X1 U5564 ( .B1(n5273), .B2(n5272), .A(n5271), .ZN(n5274) );
  AOI21_X1 U5565 ( .B1(n5276), .B2(n5275), .A(n5274), .ZN(n5279) );
  AOI22_X1 U5566 ( .A1(n5307), .A2(n5279), .B1(n5277), .B2(n5305), .ZN(U3537)
         );
  INV_X1 U5567 ( .A(REG0_REG_19__SCAN_IN), .ZN(n5278) );
  AOI22_X1 U5568 ( .A1(n5311), .A2(n5279), .B1(n5278), .B2(n5308), .ZN(U3505)
         );
  INV_X1 U5569 ( .A(n5280), .ZN(n5281) );
  OR2_X1 U5570 ( .A1(n5282), .A2(n5281), .ZN(n5294) );
  OR2_X1 U5571 ( .A1(n5295), .A2(n5283), .ZN(n5284) );
  NAND2_X1 U5572 ( .A1(n5294), .A2(n5284), .ZN(n5287) );
  INV_X1 U5573 ( .A(n5287), .ZN(n5286) );
  XNOR2_X1 U5574 ( .A(n5296), .B(n5295), .ZN(n5288) );
  AOI22_X1 U5575 ( .A1(n5288), .A2(n5298), .B1(REG2_REG_30__SCAN_IN), .B2(
        n5301), .ZN(n5285) );
  OAI21_X1 U5576 ( .B1(n5301), .B2(n5286), .A(n5285), .ZN(U3261) );
  AOI21_X1 U5577 ( .B1(n5288), .B2(n5303), .A(n5287), .ZN(n5291) );
  INV_X1 U5578 ( .A(REG1_REG_30__SCAN_IN), .ZN(n5289) );
  AOI22_X1 U5579 ( .A1(n5307), .A2(n5291), .B1(n5289), .B2(n5305), .ZN(U3548)
         );
  INV_X1 U5580 ( .A(REG0_REG_30__SCAN_IN), .ZN(n5290) );
  AOI22_X1 U5581 ( .A1(n5311), .A2(n5291), .B1(n5290), .B2(n5308), .ZN(U3516)
         );
  NAND2_X1 U5582 ( .A1(n5297), .A2(n5292), .ZN(n5293) );
  NAND2_X1 U5583 ( .A1(n5294), .A2(n5293), .ZN(n5302) );
  INV_X1 U5584 ( .A(n5302), .ZN(n5300) );
  AOI22_X1 U5585 ( .A1(n5304), .A2(n5298), .B1(n5301), .B2(
        REG2_REG_31__SCAN_IN), .ZN(n5299) );
  OAI21_X1 U5586 ( .B1(n5301), .B2(n5300), .A(n5299), .ZN(U3260) );
  AOI21_X1 U5587 ( .B1(n5304), .B2(n5303), .A(n5302), .ZN(n5310) );
  INV_X1 U5588 ( .A(REG1_REG_31__SCAN_IN), .ZN(n5306) );
  AOI22_X1 U5589 ( .A1(n5307), .A2(n5310), .B1(n5306), .B2(n5305), .ZN(U3549)
         );
  INV_X1 U5590 ( .A(REG0_REG_31__SCAN_IN), .ZN(n5309) );
  AOI22_X1 U5591 ( .A1(n5311), .A2(n5310), .B1(n5309), .B2(n5308), .ZN(U3517)
         );
  NAND2_X2 U2941 ( .A1(n2855), .A2(n4989), .ZN(n3025) );
  INV_X1 U2501 ( .A(n2965), .ZN(n3800) );
  INV_X1 U2502 ( .A(n2965), .ZN(n3844) );
  INV_X1 U2519 ( .A(n2935), .ZN(n3044) );
  CLKBUF_X1 U2625 ( .A(n3025), .Z(n4000) );
endmodule

