

module b20_C_gen_AntiSAT_k_128_9 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, keyinput_f0, 
        keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, 
        keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, 
        keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, 
        keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, 
        keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, 
        keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, 
        keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, 
        keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, 
        keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, 
        keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, 
        keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, 
        keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, 
        keyinput_f61, keyinput_f62, keyinput_f63, keyinput_g0, keyinput_g1, 
        keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, 
        keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, 
        keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, 
        keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, 
        keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, 
        keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, 
        keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, 
        keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, 
        keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, 
        keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, 
        keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, 
        keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, 
        keyinput_g62, keyinput_g63, ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, 
        ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, 
        ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, 
        ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, 
        ADD_1068_U5, ADD_1068_U46, U126, U123, P1_U3355, P1_U3354, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3439, P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, 
        P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, 
        P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, 
        P1_U3501, P1_U3504, P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, 
        P1_U3513, P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, 
        P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, 
        P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, 
        P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, 
        P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, 
        P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, 
        P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, 
        P1_U3559, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, 
        P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, 
        P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, 
        P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, 
        P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3086, P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, 
        P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, 
        P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, 
        P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, 
        P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, 
        P2_U3264, P2_U3376, P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, 
        P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, 
        P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, 
        P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, 
        P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, 
        P2_U3396, P2_U3399, P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, 
        P2_U3417, P2_U3420, P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, 
        P2_U3438, P2_U3441, P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, 
        P2_U3450, P2_U3451, P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, 
        P2_U3457, P2_U3458, P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, 
        P2_U3464, P2_U3465, P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, 
        P2_U3471, P2_U3472, P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, 
        P2_U3478, P2_U3479, P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, 
        P2_U3485, P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, 
        P2_U3211, P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, 
        P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, 
        P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, 
        P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, 
        P2_U3183, P2_U3182, P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, 
        P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, 
        P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, 
        P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, 
        P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, 
        P2_U3181, P2_U3180, P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, 
        P2_U3174, P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, 
        P2_U3167, P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, 
        P2_U3160, P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, 
        P2_U3153, P2_U3151, P2_U3150, P2_U3893 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2, keyinput_g3,
         keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, keyinput_g8,
         keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, keyinput_g13,
         keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, keyinput_g18,
         keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, keyinput_g23,
         keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, keyinput_g28,
         keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, keyinput_g33,
         keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, keyinput_g38,
         keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, keyinput_g43,
         keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, keyinput_g48,
         keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, keyinput_g53,
         keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, keyinput_g58,
         keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, keyinput_g63;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4349, n4350, n4351, n4353, n4354, n4355, n4356, n4357, n4358, n4359,
         n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369,
         n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379,
         n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389,
         n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399,
         n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409,
         n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419,
         n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429,
         n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439,
         n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449,
         n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459,
         n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469,
         n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479,
         n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489,
         n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
         n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
         n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
         n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
         n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
         n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549,
         n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559,
         n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
         n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579,
         n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
         n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
         n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
         n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
         n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
         n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
         n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
         n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
         n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
         n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
         n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
         n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
         n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
         n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
         n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
         n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739,
         n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749,
         n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759,
         n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769,
         n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779,
         n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789,
         n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799,
         n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809,
         n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819,
         n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829,
         n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839,
         n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849,
         n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859,
         n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869,
         n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879,
         n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889,
         n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899,
         n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909,
         n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919,
         n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929,
         n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
         n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949,
         n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959,
         n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
         n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979,
         n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989,
         n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999,
         n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009,
         n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019,
         n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029,
         n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039,
         n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049,
         n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059,
         n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069,
         n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079,
         n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089,
         n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099,
         n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109,
         n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119,
         n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129,
         n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139,
         n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149,
         n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159,
         n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169,
         n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179,
         n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189,
         n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199,
         n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209,
         n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219,
         n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229,
         n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239,
         n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249,
         n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259,
         n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269,
         n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279,
         n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289,
         n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299,
         n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309,
         n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319,
         n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329,
         n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339,
         n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349,
         n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359,
         n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369,
         n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379,
         n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389,
         n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399,
         n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409,
         n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419,
         n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429,
         n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439,
         n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449,
         n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459,
         n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469,
         n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479,
         n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489,
         n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499,
         n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509,
         n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519,
         n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529,
         n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539,
         n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549,
         n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559,
         n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569,
         n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579,
         n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589,
         n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599,
         n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609,
         n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619,
         n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629,
         n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639,
         n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649,
         n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659,
         n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669,
         n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679,
         n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689,
         n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699,
         n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709,
         n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719,
         n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729,
         n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739,
         n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749,
         n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759,
         n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769,
         n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779,
         n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789,
         n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799,
         n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809,
         n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819,
         n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829,
         n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839,
         n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849,
         n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859,
         n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869,
         n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879,
         n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889,
         n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899,
         n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909,
         n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919,
         n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929,
         n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939,
         n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949,
         n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959,
         n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969,
         n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979,
         n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989,
         n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999,
         n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009,
         n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019,
         n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029,
         n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039,
         n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049,
         n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059,
         n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069,
         n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079,
         n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089,
         n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099,
         n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109,
         n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119,
         n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129,
         n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139,
         n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149,
         n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159,
         n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169,
         n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179,
         n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189,
         n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199,
         n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209,
         n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219,
         n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229,
         n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239,
         n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249,
         n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259,
         n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269,
         n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279,
         n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289,
         n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299,
         n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309,
         n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319,
         n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329,
         n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339,
         n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349,
         n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359,
         n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369,
         n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379,
         n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389,
         n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399,
         n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409,
         n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419,
         n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429,
         n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439,
         n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449,
         n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459,
         n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469,
         n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479,
         n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489,
         n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499,
         n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509,
         n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519,
         n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529,
         n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539,
         n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549,
         n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559,
         n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569,
         n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579,
         n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589,
         n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599,
         n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609,
         n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619,
         n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629,
         n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639,
         n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649,
         n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659,
         n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669,
         n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679,
         n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689,
         n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699,
         n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709,
         n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719,
         n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729,
         n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739,
         n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749,
         n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759,
         n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769,
         n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779,
         n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789,
         n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799,
         n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809,
         n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819,
         n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829,
         n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839,
         n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849,
         n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859,
         n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869,
         n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879,
         n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889,
         n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899,
         n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909,
         n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919,
         n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929,
         n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939,
         n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949,
         n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959,
         n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969,
         n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979,
         n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989,
         n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999,
         n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009,
         n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019,
         n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029,
         n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039,
         n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049,
         n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059,
         n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069,
         n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079,
         n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089,
         n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099,
         n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109,
         n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119,
         n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129,
         n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139,
         n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149,
         n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159,
         n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169,
         n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179,
         n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189,
         n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199,
         n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209,
         n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219,
         n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229,
         n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239,
         n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249,
         n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259,
         n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269,
         n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279,
         n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289,
         n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299,
         n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309,
         n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319,
         n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329,
         n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339,
         n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349,
         n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359,
         n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369,
         n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379,
         n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389,
         n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399,
         n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409,
         n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419,
         n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429,
         n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439,
         n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449,
         n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459,
         n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469,
         n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479,
         n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489,
         n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499,
         n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509,
         n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519,
         n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529,
         n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539,
         n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549,
         n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559,
         n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569,
         n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579,
         n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589,
         n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599,
         n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609,
         n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619,
         n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629,
         n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639,
         n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649,
         n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659,
         n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669,
         n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679,
         n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689,
         n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699,
         n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709,
         n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719,
         n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729,
         n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739,
         n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749,
         n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759,
         n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769,
         n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779,
         n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789,
         n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799,
         n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809,
         n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819,
         n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829,
         n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839,
         n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849,
         n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859,
         n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869,
         n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879,
         n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889,
         n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899,
         n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909,
         n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919,
         n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929,
         n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939,
         n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949,
         n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959,
         n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969,
         n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979,
         n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989,
         n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999,
         n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009,
         n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019,
         n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029,
         n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039,
         n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049,
         n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059,
         n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069,
         n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079,
         n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089,
         n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099,
         n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109,
         n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119,
         n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129,
         n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139,
         n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149,
         n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159,
         n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169,
         n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179,
         n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189,
         n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199,
         n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209,
         n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219,
         n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229,
         n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239,
         n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249,
         n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259,
         n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269,
         n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279,
         n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289,
         n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299,
         n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309,
         n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319,
         n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329,
         n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339,
         n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349,
         n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359,
         n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369,
         n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379,
         n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389,
         n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399,
         n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409,
         n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419,
         n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429,
         n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439,
         n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449,
         n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459,
         n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469,
         n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479,
         n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489,
         n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499,
         n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509,
         n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519,
         n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529,
         n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539,
         n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549,
         n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559,
         n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569,
         n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579,
         n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589,
         n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599,
         n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609,
         n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619,
         n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629,
         n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639,
         n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649,
         n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659,
         n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669,
         n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679,
         n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689,
         n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699,
         n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709,
         n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719,
         n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729,
         n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739,
         n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749,
         n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759,
         n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769,
         n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779,
         n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789,
         n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799,
         n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809,
         n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819,
         n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829,
         n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839,
         n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849,
         n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859,
         n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869,
         n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879,
         n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889,
         n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899,
         n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909,
         n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919,
         n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929,
         n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939,
         n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949,
         n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959,
         n8960, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970,
         n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980,
         n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990,
         n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000,
         n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010,
         n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020,
         n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030,
         n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040,
         n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050,
         n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060,
         n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070,
         n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080,
         n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090,
         n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100,
         n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110,
         n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120,
         n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130,
         n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140,
         n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150,
         n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160,
         n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170,
         n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180,
         n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190,
         n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200,
         n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210,
         n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220,
         n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230,
         n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240,
         n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250,
         n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260,
         n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270,
         n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280,
         n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290,
         n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300,
         n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310,
         n9311, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321,
         n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331,
         n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341,
         n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351,
         n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361,
         n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371,
         n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381,
         n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391,
         n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401,
         n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411,
         n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421,
         n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431,
         n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441,
         n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451,
         n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461,
         n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471,
         n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481,
         n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491,
         n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501,
         n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511,
         n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521,
         n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531,
         n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541,
         n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551,
         n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561,
         n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571,
         n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733,
         n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743,
         n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753,
         n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763,
         n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773,
         n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783,
         n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793,
         n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803,
         n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813,
         n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823,
         n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833,
         n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843,
         n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853,
         n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863,
         n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873,
         n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883,
         n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893,
         n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903,
         n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913,
         n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923,
         n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933,
         n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943,
         n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953,
         n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963,
         n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973,
         n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983,
         n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993,
         n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002,
         n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010,
         n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018,
         n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026,
         n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034,
         n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042,
         n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050,
         n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058,
         n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066,
         n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074,
         n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082,
         n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090,
         n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098,
         n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106,
         n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114,
         n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122,
         n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130,
         n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138,
         n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146,
         n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154,
         n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162,
         n10165;

  OR2_X1 U4854 ( .A1(n6052), .A2(n9810), .ZN(n4472) );
  OR2_X1 U4855 ( .A1(n8615), .A2(n8614), .ZN(n8617) );
  NOR2_X1 U4856 ( .A1(n6239), .A2(n5989), .ZN(n5990) );
  NAND2_X1 U4857 ( .A1(n7904), .A2(n7908), .ZN(n8064) );
  OR2_X1 U4858 ( .A1(n5932), .A2(n7657), .ZN(n4659) );
  NOR2_X1 U4859 ( .A1(n7406), .A2(n4442), .ZN(n5931) );
  BUF_X2 U4861 ( .A(n5303), .Z(n4357) );
  AND2_X4 U4862 ( .A1(n5016), .A2(n9590), .ZN(n5098) );
  INV_X1 U4864 ( .A(n10165), .ZN(n4349) );
  NOR2_X1 U4865 ( .A1(n7900), .A2(n4638), .ZN(n7971) );
  AND2_X1 U4866 ( .A1(n8449), .A2(n8445), .ZN(n4596) );
  XNOR2_X1 U4867 ( .A(n6804), .B(n4461), .ZN(n6789) );
  OR3_X1 U4868 ( .A1(n7922), .A2(n7976), .A3(n7873), .ZN(n7914) );
  NAND2_X1 U4869 ( .A1(n6364), .A2(n6363), .ZN(n7817) );
  XNOR2_X1 U4870 ( .A(n8129), .B(n8249), .ZN(n7239) );
  INV_X1 U4871 ( .A(n8664), .ZN(n8639) );
  INV_X1 U4872 ( .A(n8446), .ZN(n8454) );
  INV_X1 U4873 ( .A(n8291), .ZN(n6258) );
  AND2_X1 U4874 ( .A1(n8356), .A2(n8353), .ZN(n8477) );
  AND2_X1 U4875 ( .A1(n7987), .A2(n9590), .ZN(n5303) );
  INV_X1 U4876 ( .A(n8064), .ZN(n8058) );
  INV_X1 U4877 ( .A(n7723), .ZN(n4576) );
  NAND2_X2 U4878 ( .A1(n5038), .A2(n7825), .ZN(n5145) );
  INV_X1 U4879 ( .A(n7079), .ZN(n6971) );
  INV_X1 U4880 ( .A(n9139), .ZN(n5741) );
  XNOR2_X1 U4881 ( .A(n7817), .B(n7815), .ZN(n6365) );
  NAND2_X1 U4882 ( .A1(n5509), .A2(n5508), .ZN(n9053) );
  INV_X1 U4883 ( .A(n7841), .ZN(n5712) );
  BUF_X1 U4884 ( .A(n8067), .Z(n4351) );
  NAND2_X1 U4885 ( .A1(n6365), .A2(SI_29_), .ZN(n7819) );
  INV_X1 U4886 ( .A(n6076), .ZN(n6257) );
  NAND4_X1 U4887 ( .A1(n6138), .A2(n6137), .A3(n6136), .A4(n6135), .ZN(n8535)
         );
  INV_X1 U4888 ( .A(n7157), .ZN(n7390) );
  XNOR2_X1 U4889 ( .A(n5245), .B(n5226), .ZN(n6524) );
  INV_X1 U4890 ( .A(n6804), .ZN(n8124) );
  INV_X1 U4891 ( .A(n5097), .ZN(n4354) );
  NAND4_X2 U4892 ( .A1(n4808), .A2(n4813), .A3(n4952), .A4(n4814), .ZN(n4977)
         );
  AND3_X2 U4893 ( .A1(n5482), .A2(n4810), .A3(n4809), .ZN(n4813) );
  AOI21_X2 U4894 ( .B1(n4671), .B2(n4678), .A(n4670), .ZN(n7990) );
  NAND2_X2 U4895 ( .A1(n4679), .A2(n4372), .ZN(n4678) );
  AND2_X2 U4896 ( .A1(n4710), .A2(n4709), .ZN(n5989) );
  AOI22_X2 U4897 ( .A1(n9369), .A2(n5757), .B1(n5799), .B2(n4565), .ZN(n9354)
         );
  AOI21_X2 U4898 ( .B1(n4821), .B2(n4377), .A(n4820), .ZN(n9369) );
  NOR2_X2 U4899 ( .A1(n9764), .A2(n5971), .ZN(n6700) );
  NOR2_X2 U4900 ( .A1(n9876), .A2(n9765), .ZN(n9764) );
  NAND2_X2 U4901 ( .A1(n6426), .A2(n6425), .ZN(n6439) );
  NOR2_X2 U4902 ( .A1(n9788), .A2(n9879), .ZN(n9787) );
  INV_X1 U4903 ( .A(n8124), .ZN(n4350) );
  INV_X1 U4904 ( .A(n8124), .ZN(n8129) );
  OAI21_X2 U4905 ( .B1(n5245), .B2(n5244), .A(n5246), .ZN(n5271) );
  NAND2_X2 U4906 ( .A1(n5222), .A2(n5221), .ZN(n5245) );
  XNOR2_X2 U4907 ( .A(n4667), .B(n6592), .ZN(n7351) );
  OR2_X2 U4908 ( .A1(n7049), .A2(n4668), .ZN(n4667) );
  NAND4_X2 U4909 ( .A1(n6096), .A2(n6095), .A3(n6094), .A4(n6093), .ZN(n6102)
         );
  OAI222_X1 U4910 ( .A1(P2_U3151), .A2(n6065), .B1(n8960), .B2(n8951), .C1(
        n8952), .C2(n8956), .ZN(P2_U3266) );
  XNOR2_X2 U4911 ( .A(n5984), .B(n7481), .ZN(n7476) );
  AND2_X2 U4912 ( .A1(n4713), .A2(n5983), .ZN(n5984) );
  AOI21_X4 U4913 ( .B1(n9069), .B2(n9073), .A(n8972), .ZN(n8971) );
  NAND2_X1 U4914 ( .A1(n6647), .A2(n6649), .ZN(n6648) );
  NAND2_X4 U4915 ( .A1(n4927), .A2(n4926), .ZN(n7825) );
  NAND2_X2 U4916 ( .A1(n4996), .A2(n4995), .ZN(n4927) );
  OAI21_X2 U4917 ( .B1(n4407), .B2(n4597), .A(n4596), .ZN(n8451) );
  XNOR2_X2 U4918 ( .A(n5974), .B(n6013), .ZN(n9788) );
  NOR2_X2 U4919 ( .A1(n6698), .A2(n5973), .ZN(n5974) );
  XNOR2_X2 U4920 ( .A(n5871), .B(n6056), .ZN(n5960) );
  AOI21_X2 U4921 ( .B1(n6648), .B2(n5967), .A(n9773), .ZN(n5971) );
  XNOR2_X2 U4922 ( .A(n5106), .B(n5079), .ZN(n6540) );
  NOR2_X2 U4923 ( .A1(n6695), .A2(n5915), .ZN(n5918) );
  XNOR2_X2 U4924 ( .A(n5005), .B(P1_IR_REG_1__SCAN_IN), .ZN(n9145) );
  NAND2_X1 U4925 ( .A1(n8117), .A2(n8116), .ZN(n8205) );
  NAND2_X1 U4926 ( .A1(n5778), .A2(n5777), .ZN(n8055) );
  NAND2_X1 U4927 ( .A1(n6340), .A2(n6339), .ZN(n8890) );
  AOI21_X1 U4928 ( .B1(n7587), .B2(n6226), .A(n6225), .ZN(n7579) );
  OAI21_X2 U4929 ( .B1(n6939), .B2(n6121), .A(n6120), .ZN(n7034) );
  NAND2_X1 U4930 ( .A1(n8363), .A2(n8364), .ZN(n7129) );
  NAND4_X1 U4931 ( .A1(n6117), .A2(n6116), .A3(n6115), .A4(n6114), .ZN(n8538)
         );
  NAND4_X1 U4932 ( .A1(n6108), .A2(n6107), .A3(n6106), .A4(n6105), .ZN(n8539)
         );
  NAND2_X1 U4933 ( .A1(n7937), .A2(n7941), .ZN(n7092) );
  INV_X1 U4934 ( .A(n6102), .ZN(n4861) );
  CLKBUF_X2 U4935 ( .A(n5093), .Z(n5148) );
  NAND2_X1 U4936 ( .A1(n5741), .A2(n7098), .ZN(n7937) );
  NAND4_X1 U4937 ( .A1(n6085), .A2(n6084), .A3(n6083), .A4(n6082), .ZN(n6382)
         );
  NAND4_X1 U4938 ( .A1(n6150), .A2(n6149), .A3(n6148), .A4(n6147), .ZN(n8536)
         );
  CLKBUF_X2 U4939 ( .A(n6097), .Z(n6369) );
  NAND2_X1 U4940 ( .A1(n5738), .A2(n9140), .ZN(n7936) );
  NAND2_X4 U4941 ( .A1(n6066), .A2(n6063), .ZN(n6211) );
  NAND2_X1 U4942 ( .A1(n5872), .A2(n5858), .ZN(n7692) );
  NAND2_X4 U4944 ( .A1(n5229), .A2(n8031), .ZN(n8036) );
  INV_X1 U4945 ( .A(n7098), .ZN(n5740) );
  INV_X2 U4946 ( .A(n6062), .ZN(n6066) );
  INV_X1 U4947 ( .A(n7142), .ZN(n5738) );
  BUF_X2 U4948 ( .A(n5303), .Z(n4358) );
  INV_X1 U4949 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n4707) );
  INV_X2 U4950 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n6058) );
  AOI21_X1 U4951 ( .B1(n4878), .B2(n4413), .A(n4603), .ZN(n4602) );
  OAI21_X1 U4952 ( .B1(n6457), .B2(n9873), .A(n6448), .ZN(n6449) );
  AND2_X1 U4953 ( .A1(n7918), .A2(n4460), .ZN(n4904) );
  NAND2_X1 U4954 ( .A1(n8205), .A2(n8206), .ZN(n8121) );
  AND2_X1 U4955 ( .A1(n4748), .A2(n4746), .ZN(n9090) );
  NAND2_X1 U4956 ( .A1(n4750), .A2(n4749), .ZN(n4748) );
  OR2_X1 U4957 ( .A1(n8092), .A2(n9516), .ZN(n4645) );
  OR2_X1 U4958 ( .A1(n9203), .A2(n7840), .ZN(n7975) );
  NAND2_X1 U4959 ( .A1(n6371), .A2(n6370), .ZN(n8307) );
  XNOR2_X1 U4960 ( .A(n7824), .B(n7823), .ZN(n8289) );
  NAND2_X1 U4961 ( .A1(n7819), .A2(n7818), .ZN(n7824) );
  NAND2_X1 U4962 ( .A1(n4773), .A2(n4771), .ZN(n8274) );
  NAND2_X1 U4963 ( .A1(n8443), .A2(n8444), .ZN(n8656) );
  NAND2_X1 U4964 ( .A1(n6353), .A2(n6352), .ZN(n8647) );
  OR2_X1 U4965 ( .A1(n8890), .A2(n8639), .ZN(n8443) );
  AND2_X1 U4966 ( .A1(n4694), .A2(n4392), .ZN(n8698) );
  NAND2_X1 U4967 ( .A1(n5667), .A2(n5666), .ZN(n9231) );
  NAND2_X1 U4968 ( .A1(n5773), .A2(n5772), .ZN(n6362) );
  AND2_X1 U4969 ( .A1(n7614), .A2(n7615), .ZN(n7560) );
  AND2_X2 U4970 ( .A1(n5606), .A2(n5605), .ZN(n9548) );
  NAND2_X1 U4971 ( .A1(n5280), .A2(n5279), .ZN(n4743) );
  NAND2_X1 U4972 ( .A1(n5636), .A2(n5635), .ZN(n5660) );
  AOI21_X1 U4973 ( .B1(n4757), .B2(n4382), .A(n4756), .ZN(n4755) );
  AOI21_X1 U4974 ( .B1(P1_REG2_REG_14__SCAN_IN), .B2(n9665), .A(n9657), .ZN(
        n8004) );
  OR2_X1 U4975 ( .A1(n7481), .A2(n5931), .ZN(n5932) );
  NAND2_X1 U4976 ( .A1(n5414), .A2(n5413), .ZN(n9514) );
  NAND2_X1 U4977 ( .A1(n8228), .A2(n8230), .ZN(n8229) );
  NAND4_X2 U4978 ( .A1(n6348), .A2(n6347), .A3(n6346), .A4(n6345), .ZN(n8664)
         );
  AND2_X1 U4979 ( .A1(n8247), .A2(n7237), .ZN(n4807) );
  NAND2_X1 U4980 ( .A1(n5276), .A2(n5275), .ZN(n9629) );
  NAND2_X1 U4981 ( .A1(n4723), .A2(n4722), .ZN(n4721) );
  AND2_X1 U4982 ( .A1(n6302), .A2(n6301), .ZN(n8711) );
  NAND2_X1 U4983 ( .A1(n4619), .A2(n5272), .ZN(n5289) );
  XNOR2_X1 U4984 ( .A(n5271), .B(n4385), .ZN(n6165) );
  AOI21_X1 U4985 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n6925), .A(n6916), .ZN(
        n9605) );
  NOR2_X1 U4986 ( .A1(n6758), .A2(n5977), .ZN(n5978) );
  NOR2_X1 U4987 ( .A1(n6760), .A2(n6759), .ZN(n6758) );
  INV_X1 U4988 ( .A(n6079), .ZN(n4461) );
  AOI21_X1 U4989 ( .B1(P1_REG2_REG_7__SCAN_IN), .B2(n6600), .A(n6599), .ZN(
        n6603) );
  NOR2_X1 U4990 ( .A1(n9787), .A2(n5975), .ZN(n6760) );
  NOR2_X1 U4991 ( .A1(n6756), .A2(n5924), .ZN(n5925) );
  AND4_X1 U4992 ( .A1(n6164), .A2(n6163), .A3(n6162), .A4(n6161), .ZN(n7396)
         );
  AND2_X1 U4993 ( .A1(n6153), .A2(n6152), .ZN(n9850) );
  AND3_X1 U4994 ( .A1(n6100), .A2(n6099), .A3(n6098), .ZN(n9827) );
  INV_X2 U4995 ( .A(n6369), .ZN(n8288) );
  AOI21_X1 U4996 ( .B1(n4935), .B2(n4934), .A(n4420), .ZN(n4933) );
  INV_X1 U4997 ( .A(n8031), .ZN(n5677) );
  NAND2_X1 U4998 ( .A1(n5078), .A2(n5077), .ZN(n9139) );
  CLKBUF_X2 U4999 ( .A(n6091), .Z(n4360) );
  NAND4_X1 U5000 ( .A1(n5033), .A2(n5032), .A3(n5031), .A4(n5030), .ZN(n5736)
         );
  NAND2_X1 U5001 ( .A1(n6062), .A2(n6063), .ZN(n6091) );
  MUX2_X1 U5003 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5857), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n5858) );
  NAND2_X1 U5004 ( .A1(n4450), .A2(n4379), .ZN(n4929) );
  INV_X1 U5005 ( .A(n6065), .ZN(n6063) );
  INV_X2 U5006 ( .A(n8514), .ZN(n6004) );
  INV_X2 U5007 ( .A(n4354), .ZN(n4355) );
  INV_X2 U5008 ( .A(n4354), .ZN(n4356) );
  NAND2_X1 U5009 ( .A1(n8946), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6057) );
  NAND2_X1 U5010 ( .A1(n5853), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5861) );
  NOR2_X1 U5011 ( .A1(n5866), .A2(n4373), .ZN(n6059) );
  OAI21_X1 U5012 ( .B1(n5866), .B2(n4902), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n5871) );
  OR2_X1 U5013 ( .A1(n4932), .A2(n5536), .ZN(n4930) );
  CLKBUF_X2 U5014 ( .A(n5865), .Z(n5866) );
  XNOR2_X1 U5016 ( .A(n5922), .B(n5921), .ZN(n6764) );
  NAND2_X1 U5017 ( .A1(n5485), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4976) );
  XNOR2_X1 U5018 ( .A(n5143), .B(n5118), .ZN(n5141) );
  XNOR2_X1 U5019 ( .A(n5883), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7481) );
  OAI21_X1 U5020 ( .B1(n6053), .B2(n5117), .A(n5116), .ZN(n5143) );
  XNOR2_X1 U5021 ( .A(n4986), .B(n4985), .ZN(n7927) );
  NAND2_X1 U5022 ( .A1(n4964), .A2(n4381), .ZN(n7644) );
  NAND2_X1 U5023 ( .A1(n4418), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4983) );
  OR2_X1 U5024 ( .A1(n4990), .A2(n5010), .ZN(n4991) );
  OR2_X1 U5025 ( .A1(n9581), .A2(n5010), .ZN(n5012) );
  NAND2_X1 U5026 ( .A1(n4984), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4986) );
  NAND2_X2 U5027 ( .A1(n7825), .A2(P1_U3086), .ZN(n9588) );
  OAI21_X1 U5028 ( .B1(n6003), .B2(n5898), .A(n5899), .ZN(n6479) );
  OAI21_X1 U5029 ( .B1(n6003), .B2(n5961), .A(n5963), .ZN(n6476) );
  OR2_X1 U5030 ( .A1(n4902), .A2(P2_IR_REG_28__SCAN_IN), .ZN(n4373) );
  NAND2_X1 U5031 ( .A1(n4998), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n4926) );
  AND2_X1 U5032 ( .A1(n4811), .A2(n4812), .ZN(n4808) );
  AND2_X1 U5033 ( .A1(n4965), .A2(n4859), .ZN(n4858) );
  NAND2_X1 U5034 ( .A1(n9763), .A2(n4707), .ZN(n5897) );
  MUX2_X1 U5035 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5895), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n5896) );
  NAND3_X1 U5036 ( .A1(n4707), .A2(n4708), .A3(n5828), .ZN(n5901) );
  NOR2_X1 U5037 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n4979) );
  INV_X4 U5038 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  INV_X2 U5039 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5837) );
  NOR2_X1 U5040 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .ZN(
        n5854) );
  NOR2_X1 U5041 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n5104) );
  NOR2_X1 U5042 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5053) );
  INV_X1 U5043 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5862) );
  INV_X4 U5044 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U5045 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4997) );
  NOR2_X1 U5046 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n5832) );
  INV_X1 U5047 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n5011) );
  INV_X1 U5048 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n4975) );
  INV_X1 U5049 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5891) );
  NOR2_X1 U5050 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n4812) );
  NOR2_X1 U5051 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n4811) );
  INV_X1 U5052 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5828) );
  OAI21_X1 U5053 ( .B1(n9785), .B2(n4662), .A(n4661), .ZN(n6756) );
  NAND2_X1 U5054 ( .A1(n5900), .A2(P2_IR_REG_2__SCAN_IN), .ZN(n5904) );
  XNOR2_X2 U5055 ( .A(n4983), .B(P1_IR_REG_21__SCAN_IN), .ZN(n7924) );
  AND2_X1 U5056 ( .A1(n5901), .A2(n5902), .ZN(n5903) );
  AOI22_X2 U5057 ( .A1(n9339), .A2(n5759), .B1(n5804), .B2(n9349), .ZN(n9330)
         );
  AOI22_X2 U5058 ( .A1(n9354), .A2(n5758), .B1(n9126), .B2(n9363), .ZN(n9339)
         );
  XNOR2_X2 U5060 ( .A(n4651), .B(P1_IR_REG_27__SCAN_IN), .ZN(n6515) );
  AND2_X1 U5061 ( .A1(n7987), .A2(n5015), .ZN(n5097) );
  NOR2_X2 U5062 ( .A1(n6323), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6330) );
  AOI21_X2 U5063 ( .B1(n8733), .B2(n8738), .A(n6275), .ZN(n8719) );
  OAI22_X2 U5064 ( .A1(n8744), .A2(n6266), .B1(n8764), .B2(n8846), .ZN(n8733)
         );
  NOR2_X2 U5065 ( .A1(n5887), .A2(n5834), .ZN(n5884) );
  AND2_X1 U5066 ( .A1(n5840), .A2(n5885), .ZN(n4862) );
  NOR2_X2 U5067 ( .A1(n6382), .A2(n6645), .ZN(n8316) );
  NOR2_X2 U5068 ( .A1(n5865), .A2(P2_IR_REG_21__SCAN_IN), .ZN(n5863) );
  OAI21_X1 U5069 ( .B1(n6439), .B2(P2_D_REG_0__SCAN_IN), .A(n6617), .ZN(n6780)
         );
  OAI21_X2 U5070 ( .B1(n7034), .B2(n6132), .A(n6131), .ZN(n7123) );
  NAND2_X2 U5071 ( .A1(n8121), .A2(n8120), .ZN(n8179) );
  INV_X1 U5072 ( .A(n6804), .ZN(n4361) );
  OAI21_X2 U5073 ( .B1(n8098), .B2(n8527), .A(n7578), .ZN(n8787) );
  XNOR2_X2 U5074 ( .A(n7557), .B(n7993), .ZN(n7507) );
  OAI21_X2 U5075 ( .B1(n6895), .B2(n4806), .A(n4805), .ZN(n7397) );
  XNOR2_X2 U5076 ( .A(n8113), .B(n8114), .ZN(n8156) );
  XNOR2_X2 U5077 ( .A(n6057), .B(n8947), .ZN(n6062) );
  OAI22_X2 U5078 ( .A1(n8239), .A2(n8238), .B1(n8105), .B2(n8746), .ZN(n8164)
         );
  XNOR2_X2 U5079 ( .A(n4530), .B(P2_IR_REG_27__SCAN_IN), .ZN(n8514) );
  INV_X1 U5080 ( .A(n8514), .ZN(n6002) );
  INV_X1 U5081 ( .A(n8477), .ZN(n6390) );
  AND2_X1 U5082 ( .A1(n5635), .A2(n5623), .ZN(n5633) );
  NAND2_X1 U5083 ( .A1(n4918), .A2(n4400), .ZN(n5481) );
  INV_X1 U5084 ( .A(n5478), .ZN(n4917) );
  OAI21_X1 U5085 ( .B1(n5362), .B2(n5361), .A(n5360), .ZN(n5384) );
  INV_X1 U5086 ( .A(n5358), .ZN(n5359) );
  AND2_X1 U5087 ( .A1(n4766), .A2(n4961), .ZN(n4765) );
  INV_X1 U5088 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n4766) );
  NOR2_X1 U5089 ( .A1(n4857), .A2(P1_IR_REG_28__SCAN_IN), .ZN(n4515) );
  AND2_X1 U5090 ( .A1(n4610), .A2(n8389), .ZN(n4606) );
  AND2_X1 U5091 ( .A1(n4610), .A2(n8392), .ZN(n4607) );
  NOR2_X1 U5092 ( .A1(n4409), .A2(n4593), .ZN(n4592) );
  NAND2_X1 U5093 ( .A1(n8442), .A2(n8441), .ZN(n4597) );
  INV_X1 U5094 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5851) );
  AND2_X1 U5095 ( .A1(n9203), .A2(n9115), .ZN(n4505) );
  NAND2_X1 U5096 ( .A1(n4798), .A2(n4799), .ZN(n4797) );
  INV_X1 U5097 ( .A(n8141), .ZN(n4798) );
  INV_X1 U5098 ( .A(n7426), .ZN(n8512) );
  AND2_X1 U5099 ( .A1(n6764), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5924) );
  NOR2_X1 U5100 ( .A1(n9797), .A2(n5949), .ZN(n8615) );
  OR2_X1 U5101 ( .A1(n6316), .A2(n8700), .ZN(n8460) );
  OR2_X1 U5102 ( .A1(n8727), .A2(n8735), .ZN(n8420) );
  NAND2_X1 U5103 ( .A1(n4697), .A2(n4696), .ZN(n8756) );
  AOI21_X1 U5104 ( .B1(n4698), .B2(n4699), .A(n4425), .ZN(n4696) );
  OR2_X1 U5105 ( .A1(n8857), .A2(n8777), .ZN(n8403) );
  NAND2_X1 U5106 ( .A1(n6405), .A2(n7426), .ZN(n6783) );
  NAND2_X1 U5107 ( .A1(n8516), .A2(n8310), .ZN(n8446) );
  OR2_X1 U5108 ( .A1(n6439), .A2(n6438), .ZN(n6453) );
  NAND2_X1 U5109 ( .A1(n7924), .A2(n7927), .ZN(n5021) );
  INV_X1 U5110 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n4958) );
  INV_X1 U5111 ( .A(n4940), .ZN(n4934) );
  AOI21_X1 U5112 ( .B1(n4940), .B2(n5288), .A(n4939), .ZN(n4938) );
  INV_X1 U5113 ( .A(n5313), .ZN(n4939) );
  OAI21_X1 U5114 ( .B1(n6053), .B2(n5084), .A(n5083), .ZN(n5114) );
  NAND2_X1 U5115 ( .A1(n6053), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n5083) );
  INV_X1 U5116 ( .A(n6211), .ZN(n6308) );
  AND2_X1 U5117 ( .A1(n4880), .A2(n4879), .ZN(n4363) );
  INV_X1 U5118 ( .A(n8458), .ZN(n4879) );
  OAI21_X1 U5119 ( .B1(n8303), .B2(n8302), .A(n4881), .ZN(n4880) );
  INV_X1 U5120 ( .A(n4360), .ZN(n6321) );
  INV_X1 U5121 ( .A(n6090), .ZN(n6373) );
  AND4_X1 U5122 ( .A1(n6174), .A2(n6173), .A3(n6172), .A4(n6171), .ZN(n7258)
         );
  OR2_X1 U5123 ( .A1(n6211), .A2(n6941), .ZN(n6115) );
  CLKBUF_X1 U5124 ( .A(n5887), .Z(n5888) );
  INV_X1 U5125 ( .A(n7042), .ZN(n4722) );
  AND2_X1 U5126 ( .A1(n7048), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n4668) );
  NAND2_X1 U5127 ( .A1(n5860), .A2(n5859), .ZN(n6738) );
  NAND2_X1 U5128 ( .A1(n4716), .A2(n4718), .ZN(n4719) );
  INV_X1 U5129 ( .A(n8611), .ZN(n4718) );
  OAI21_X1 U5130 ( .B1(n9801), .B2(n9802), .A(n4717), .ZN(n4716) );
  AOI21_X1 U5131 ( .B1(n4867), .B2(n4865), .A(n4864), .ZN(n4863) );
  INV_X1 U5132 ( .A(n4867), .ZN(n4866) );
  INV_X1 U5133 ( .A(n8443), .ZN(n4864) );
  NAND2_X1 U5134 ( .A1(n8904), .A2(n8700), .ZN(n6317) );
  AOI21_X1 U5135 ( .B1(n4693), .B2(n4690), .A(n4375), .ZN(n4688) );
  OR2_X1 U5136 ( .A1(n8225), .A2(n8721), .ZN(n8423) );
  NAND2_X1 U5137 ( .A1(n6396), .A2(n8399), .ZN(n8794) );
  AOI21_X1 U5138 ( .B1(n4876), .B2(n4367), .A(n4875), .ZN(n4874) );
  INV_X1 U5139 ( .A(n8364), .ZN(n4893) );
  INV_X1 U5140 ( .A(n7123), .ZN(n4679) );
  INV_X1 U5141 ( .A(n8745), .ZN(n8790) );
  INV_X1 U5142 ( .A(n8763), .ZN(n8788) );
  NAND2_X1 U5143 ( .A1(n6441), .A2(n8304), .ZN(n8759) );
  NAND2_X1 U5144 ( .A1(n5953), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5957) );
  AND2_X1 U5145 ( .A1(n5712), .A2(n7924), .ZN(n6508) );
  AND2_X1 U5146 ( .A1(n5686), .A2(n4967), .ZN(n4968) );
  AND2_X1 U5147 ( .A1(n4978), .A2(n4979), .ZN(n5273) );
  AOI21_X1 U5148 ( .B1(n4636), .B2(n4638), .A(n4635), .ZN(n4634) );
  INV_X1 U5149 ( .A(n7799), .ZN(n4635) );
  OR2_X1 U5150 ( .A1(n9336), .A2(n9124), .ZN(n5760) );
  INV_X1 U5151 ( .A(n4822), .ZN(n4820) );
  OAI21_X1 U5152 ( .B1(n7933), .B2(n4649), .A(n4647), .ZN(n6963) );
  INV_X1 U5153 ( .A(n4648), .ZN(n4647) );
  INV_X1 U5154 ( .A(n7937), .ZN(n4649) );
  INV_X1 U5155 ( .A(n5145), .ZN(n5487) );
  XNOR2_X1 U5156 ( .A(n5014), .B(P1_IR_REG_29__SCAN_IN), .ZN(n5015) );
  NAND2_X1 U5157 ( .A1(n5013), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5014) );
  NAND2_X1 U5158 ( .A1(n4913), .A2(n5620), .ZN(n5634) );
  NAND2_X1 U5159 ( .A1(n5619), .A2(n5618), .ZN(n4913) );
  AOI21_X1 U5160 ( .B1(n4366), .B2(P1_IR_REG_31__SCAN_IN), .A(
        P1_IR_REG_18__SCAN_IN), .ZN(n4762) );
  NAND2_X1 U5161 ( .A1(n4918), .A2(n4919), .ZN(n5479) );
  NOR2_X1 U5162 ( .A1(n4594), .A2(n4404), .ZN(n4589) );
  AOI21_X1 U5163 ( .B1(n4610), .B2(n8401), .A(n4609), .ZN(n4608) );
  NOR2_X1 U5164 ( .A1(n4592), .A2(n4584), .ZN(n4583) );
  NAND2_X1 U5165 ( .A1(n4376), .A2(n8446), .ZN(n4584) );
  INV_X1 U5166 ( .A(n4589), .ZN(n4586) );
  NOR2_X1 U5167 ( .A1(n4590), .A2(n8446), .ZN(n4585) );
  NOR2_X1 U5168 ( .A1(n4594), .A2(n4591), .ZN(n4590) );
  INV_X1 U5169 ( .A(n8779), .ZN(n4591) );
  OAI22_X1 U5170 ( .A1(n4589), .A2(n8446), .B1(n8454), .B2(n4592), .ZN(n4588)
         );
  NOR2_X1 U5171 ( .A1(n4616), .A2(n8446), .ZN(n4615) );
  INV_X1 U5172 ( .A(n8411), .ZN(n4616) );
  NAND2_X1 U5173 ( .A1(n8421), .A2(n4618), .ZN(n4617) );
  AND2_X1 U5174 ( .A1(n8420), .A2(n8446), .ZN(n4618) );
  OR2_X1 U5175 ( .A1(n7778), .A2(n7919), .ZN(n4527) );
  NAND2_X1 U5176 ( .A1(n4511), .A2(n4507), .ZN(n7776) );
  INV_X1 U5177 ( .A(n7775), .ZN(n4511) );
  AOI21_X1 U5178 ( .B1(n4509), .B2(n4508), .A(n4426), .ZN(n4507) );
  NOR2_X1 U5179 ( .A1(n4493), .A2(n4417), .ZN(n4492) );
  INV_X1 U5180 ( .A(n7797), .ZN(n4493) );
  NAND2_X1 U5181 ( .A1(n8062), .A2(n7799), .ZN(n7896) );
  NAND2_X1 U5182 ( .A1(n4432), .A2(n7797), .ZN(n4491) );
  INV_X1 U5183 ( .A(n7881), .ZN(n4489) );
  INV_X1 U5184 ( .A(n7802), .ZN(n4488) );
  OR2_X1 U5185 ( .A1(n7794), .A2(n7793), .ZN(n4494) );
  AOI21_X1 U5186 ( .B1(n4516), .B2(n4517), .A(n4522), .ZN(n7791) );
  NOR2_X1 U5187 ( .A1(n4518), .A2(n4523), .ZN(n4517) );
  INV_X1 U5188 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5875) );
  AND2_X1 U5189 ( .A1(n7975), .A2(n7910), .ZN(n4506) );
  NOR2_X1 U5190 ( .A1(n4632), .A2(n4629), .ZN(n4628) );
  INV_X1 U5191 ( .A(n5798), .ZN(n4632) );
  NAND2_X1 U5192 ( .A1(n7528), .A2(n7760), .ZN(n5797) );
  NAND2_X1 U5193 ( .A1(n5440), .A2(n4384), .ZN(n4923) );
  AND2_X1 U5194 ( .A1(n4786), .A2(n4785), .ZN(n4784) );
  INV_X1 U5195 ( .A(n8221), .ZN(n4785) );
  NOR2_X1 U5196 ( .A1(n4782), .A2(n8221), .ZN(n4781) );
  INV_X1 U5197 ( .A(n4787), .ZN(n4782) );
  INV_X1 U5198 ( .A(n4946), .ZN(n4790) );
  NAND2_X1 U5199 ( .A1(n7504), .A2(n7503), .ZN(n7557) );
  AND2_X1 U5200 ( .A1(n6650), .A2(n5907), .ZN(n5910) );
  NAND2_X1 U5201 ( .A1(n5966), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5907) );
  AND2_X1 U5202 ( .A1(n4666), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n4665) );
  INV_X1 U5203 ( .A(n4538), .ZN(n4537) );
  NOR2_X1 U5204 ( .A1(n5914), .A2(n5913), .ZN(n5915) );
  NAND2_X1 U5205 ( .A1(n4529), .A2(n8596), .ZN(n9806) );
  OR2_X1 U5206 ( .A1(n8598), .A2(n8594), .ZN(n4529) );
  NAND2_X1 U5207 ( .A1(n9806), .A2(n9805), .ZN(n9804) );
  OR2_X1 U5208 ( .A1(n8107), .A2(n8722), .ZN(n8415) );
  AOI21_X1 U5209 ( .B1(n4700), .B2(n6238), .A(n4429), .ZN(n4698) );
  NAND2_X1 U5210 ( .A1(n7197), .A2(n6178), .ZN(n4470) );
  INV_X1 U5211 ( .A(n8315), .ZN(n8310) );
  AND2_X1 U5212 ( .A1(n8493), .A2(n4684), .ZN(n4683) );
  INV_X1 U5213 ( .A(n6349), .ZN(n4681) );
  INV_X1 U5214 ( .A(n4683), .ZN(n4682) );
  INV_X1 U5215 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5850) );
  INV_X1 U5216 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5879) );
  AND2_X1 U5217 ( .A1(n4770), .A2(n5946), .ZN(n4769) );
  NAND2_X1 U5218 ( .A1(n5874), .A2(n5835), .ZN(n5878) );
  INV_X1 U5219 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5829) );
  INV_X1 U5220 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5831) );
  INV_X1 U5221 ( .A(n5356), .ZN(n4760) );
  BUF_X1 U5222 ( .A(n5229), .Z(n5675) );
  NOR2_X1 U5223 ( .A1(n9202), .A2(n7838), .ZN(n4500) );
  AND3_X1 U5224 ( .A1(n7810), .A2(n4954), .A3(n7809), .ZN(n7814) );
  MUX2_X1 U5225 ( .A(n7908), .B(n7904), .S(n7919), .Z(n7813) );
  NOR2_X1 U5226 ( .A1(n7808), .A2(n7807), .ZN(n7809) );
  NAND2_X1 U5227 ( .A1(n4503), .A2(n4502), .ZN(n4501) );
  NAND2_X1 U5228 ( .A1(n4505), .A2(n9202), .ZN(n4502) );
  NAND2_X1 U5229 ( .A1(n4506), .A2(n9532), .ZN(n4503) );
  NAND2_X1 U5230 ( .A1(n4506), .A2(n4498), .ZN(n4497) );
  NOR2_X1 U5231 ( .A1(n9532), .A2(n7919), .ZN(n4498) );
  OR2_X1 U5232 ( .A1(n9231), .A2(n5818), .ZN(n7883) );
  NAND2_X1 U5233 ( .A1(n9231), .A2(n5818), .ZN(n7799) );
  INV_X1 U5234 ( .A(n5764), .ZN(n4849) );
  NOR2_X1 U5235 ( .A1(n7535), .A2(n9066), .ZN(n7536) );
  INV_X1 U5236 ( .A(n5021), .ZN(n7066) );
  NAND2_X1 U5237 ( .A1(n5784), .A2(n7060), .ZN(n4620) );
  OR2_X1 U5238 ( .A1(n9245), .A2(n9249), .ZN(n9246) );
  INV_X1 U5239 ( .A(n9544), .ZN(n9260) );
  INV_X1 U5240 ( .A(n7644), .ZN(n5686) );
  NAND2_X1 U5241 ( .A1(n4910), .A2(n4914), .ZN(n5636) );
  INV_X1 U5242 ( .A(n4915), .ZN(n4914) );
  AND2_X1 U5243 ( .A1(n5661), .A2(n5639), .ZN(n5659) );
  INV_X1 U5244 ( .A(n5292), .ZN(n4941) );
  NAND2_X1 U5245 ( .A1(n5271), .A2(n4385), .ZN(n4619) );
  NAND2_X1 U5246 ( .A1(n5000), .A2(n5001), .ZN(n5057) );
  INV_X1 U5247 ( .A(SI_12_), .ZN(n9989) );
  AND2_X1 U5248 ( .A1(n6440), .A2(n6846), .ZN(n6747) );
  AND2_X1 U5249 ( .A1(n4774), .A2(n4437), .ZN(n4772) );
  INV_X1 U5250 ( .A(n8500), .ZN(n8499) );
  AND2_X1 U5251 ( .A1(n6648), .A2(n5967), .ZN(n5968) );
  NAND2_X1 U5252 ( .A1(n5910), .A2(n9773), .ZN(n4666) );
  OR2_X1 U5253 ( .A1(n6007), .A2(n4536), .ZN(n6691) );
  NAND2_X1 U5254 ( .A1(n6692), .A2(n4537), .ZN(n4536) );
  XNOR2_X1 U5255 ( .A(n5918), .B(n6013), .ZN(n9785) );
  AND2_X1 U5256 ( .A1(n4534), .A2(n4532), .ZN(n9780) );
  NAND2_X1 U5257 ( .A1(n9781), .A2(n4533), .ZN(n4532) );
  OR2_X1 U5258 ( .A1(n6007), .A2(n4535), .ZN(n4534) );
  INV_X1 U5259 ( .A(n6010), .ZN(n4533) );
  NOR2_X1 U5260 ( .A1(n5918), .A2(n6013), .ZN(n5919) );
  NOR2_X1 U5261 ( .A1(n5926), .A2(n6952), .ZN(n7051) );
  OR2_X1 U5262 ( .A1(n7340), .A2(n5982), .ZN(n4715) );
  NAND2_X1 U5263 ( .A1(n4715), .A2(n4714), .ZN(n4713) );
  INV_X1 U5264 ( .A(n7417), .ZN(n4714) );
  NAND2_X1 U5265 ( .A1(n7478), .A2(n7479), .ZN(n7477) );
  OR2_X1 U5266 ( .A1(n7473), .A2(n4658), .ZN(n4657) );
  OR2_X1 U5267 ( .A1(n7657), .A2(n7474), .ZN(n4658) );
  NOR2_X1 U5268 ( .A1(n7653), .A2(n6200), .ZN(n4463) );
  OAI21_X1 U5269 ( .B1(n8577), .B2(n4653), .A(n4652), .ZN(n8602) );
  NAND2_X1 U5270 ( .A1(n4656), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n4653) );
  INV_X1 U5271 ( .A(n8603), .ZN(n4656) );
  OR2_X1 U5272 ( .A1(n8577), .A2(n8578), .ZN(n4655) );
  INV_X1 U5273 ( .A(n8496), .ZN(n6378) );
  NAND2_X1 U5274 ( .A1(n6404), .A2(n6403), .ZN(n8303) );
  NOR2_X1 U5275 ( .A1(n6402), .A2(n4871), .ZN(n4870) );
  INV_X1 U5276 ( .A(n8434), .ZN(n4871) );
  INV_X1 U5277 ( .A(n4898), .ZN(n4897) );
  AND2_X1 U5278 ( .A1(n4899), .A2(n8423), .ZN(n4898) );
  OR2_X1 U5279 ( .A1(n4691), .A2(n4439), .ZN(n4690) );
  INV_X1 U5280 ( .A(n4695), .ZN(n4691) );
  NAND2_X1 U5281 ( .A1(n8712), .A2(n8708), .ZN(n4900) );
  AND2_X1 U5282 ( .A1(n6293), .A2(n6292), .ZN(n8721) );
  NOR2_X1 U5283 ( .A1(n8107), .A2(n6274), .ZN(n6275) );
  NAND2_X1 U5284 ( .A1(n8756), .A2(n8757), .ZN(n8744) );
  NAND2_X1 U5285 ( .A1(n6398), .A2(n8409), .ZN(n8768) );
  AND2_X1 U5286 ( .A1(n8409), .A2(n8407), .ZN(n8779) );
  AND2_X1 U5287 ( .A1(n8403), .A2(n8402), .ZN(n8795) );
  NOR2_X1 U5288 ( .A1(n8787), .A2(n8795), .ZN(n8785) );
  AND2_X1 U5289 ( .A1(n7590), .A2(n8528), .ZN(n6225) );
  NAND2_X1 U5290 ( .A1(n4433), .A2(n8395), .ZN(n4876) );
  NAND2_X1 U5291 ( .A1(n4674), .A2(n4672), .ZN(n6197) );
  INV_X1 U5292 ( .A(n4673), .ZN(n4672) );
  AOI21_X1 U5293 ( .B1(n4892), .B2(n6389), .A(n4890), .ZN(n4889) );
  INV_X1 U5294 ( .A(n8356), .ZN(n4890) );
  AND2_X1 U5295 ( .A1(n6795), .A2(n8454), .ZN(n8745) );
  OR2_X1 U5296 ( .A1(n6097), .A2(n6498), .ZN(n6078) );
  NAND2_X1 U5297 ( .A1(n4669), .A2(n6834), .ZN(n6876) );
  AND2_X1 U5298 ( .A1(n6415), .A2(n8454), .ZN(n8763) );
  NAND2_X1 U5299 ( .A1(n6850), .A2(n6849), .ZN(n6853) );
  CLKBUF_X1 U5300 ( .A(n6780), .Z(n6846) );
  INV_X1 U5301 ( .A(n8753), .ZN(n8846) );
  OR2_X1 U5302 ( .A1(n6851), .A2(n8516), .ZN(n9828) );
  INV_X1 U5303 ( .A(n7692), .ZN(n6425) );
  INV_X1 U5304 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n6060) );
  NAND2_X1 U5305 ( .A1(n5843), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5847) );
  INV_X1 U5306 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5846) );
  INV_X1 U5307 ( .A(n9000), .ZN(n4747) );
  NAND2_X1 U5308 ( .A1(n4752), .A2(n5617), .ZN(n4751) );
  INV_X1 U5309 ( .A(n9040), .ZN(n4752) );
  INV_X1 U5310 ( .A(n4732), .ZN(n4731) );
  OAI21_X1 U5311 ( .B1(n7599), .B2(n4733), .A(n7622), .ZN(n4732) );
  INV_X1 U5312 ( .A(n4738), .ZN(n4737) );
  OAI21_X1 U5313 ( .B1(n8993), .B2(n4739), .A(n5553), .ZN(n4738) );
  NAND2_X1 U5314 ( .A1(n5534), .A2(n5533), .ZN(n4739) );
  INV_X1 U5315 ( .A(n5533), .ZN(n4740) );
  NAND2_X1 U5316 ( .A1(n9071), .A2(n9070), .ZN(n9069) );
  INV_X1 U5317 ( .A(n7981), .ZN(n4909) );
  AND4_X1 U5318 ( .A1(n5307), .A2(n5306), .A3(n5305), .A4(n5304), .ZN(n7460)
         );
  AND4_X1 U5319 ( .A1(n5243), .A2(n5242), .A3(n5241), .A4(n5240), .ZN(n7324)
         );
  AND4_X1 U5320 ( .A1(n5163), .A2(n5162), .A3(n5161), .A4(n5160), .ZN(n7722)
         );
  AND2_X1 U5321 ( .A1(n6507), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6461) );
  AOI21_X1 U5322 ( .B1(n4839), .B2(n4842), .A(n4422), .ZN(n4836) );
  NOR2_X1 U5323 ( .A1(n9246), .A2(n9231), .ZN(n9230) );
  AND2_X1 U5324 ( .A1(n7883), .A2(n7799), .ZN(n9225) );
  OR2_X1 U5325 ( .A1(n9277), .A2(n9002), .ZN(n9253) );
  NAND2_X1 U5326 ( .A1(n4431), .A2(n4855), .ZN(n4850) );
  NOR2_X1 U5327 ( .A1(n5762), .A2(n4852), .ZN(n4851) );
  INV_X1 U5328 ( .A(n4957), .ZN(n4852) );
  AND2_X1 U5329 ( .A1(n7790), .A2(n9270), .ZN(n9288) );
  NAND2_X1 U5330 ( .A1(n9321), .A2(n9320), .ZN(n9319) );
  NAND2_X1 U5331 ( .A1(n4828), .A2(n4826), .ZN(n4825) );
  NAND2_X1 U5332 ( .A1(n4832), .A2(n9107), .ZN(n4831) );
  NAND2_X1 U5333 ( .A1(n9407), .A2(n9409), .ZN(n9408) );
  OAI21_X1 U5334 ( .B1(n7178), .B2(n4819), .A(n7108), .ZN(n4818) );
  INV_X1 U5335 ( .A(n5746), .ZN(n4819) );
  NAND2_X1 U5336 ( .A1(n6463), .A2(n6461), .ZN(n6506) );
  OR2_X1 U5337 ( .A1(n5145), .A2(n6490), .ZN(n5092) );
  AND2_X1 U5338 ( .A1(n5822), .A2(n7927), .ZN(n9477) );
  OR2_X1 U5339 ( .A1(n5145), .A2(n6488), .ZN(n5007) );
  NAND2_X1 U5340 ( .A1(n4424), .A2(n4858), .ZN(n4857) );
  NAND2_X1 U5341 ( .A1(n4562), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4993) );
  NOR2_X1 U5342 ( .A1(n4563), .A2(n4856), .ZN(n4560) );
  INV_X1 U5343 ( .A(n4977), .ZN(n4561) );
  XNOR2_X1 U5344 ( .A(n5771), .B(n5770), .ZN(n7693) );
  XNOR2_X1 U5345 ( .A(n4993), .B(P1_IR_REG_26__SCAN_IN), .ZN(n5700) );
  XNOR2_X1 U5346 ( .A(n5660), .B(n5659), .ZN(n7687) );
  NOR2_X1 U5347 ( .A1(n4977), .A2(n4563), .ZN(n4559) );
  NAND2_X1 U5348 ( .A1(n5273), .A2(n4980), .ZN(n5297) );
  NAND2_X1 U5349 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), 
        .ZN(n4763) );
  NAND2_X1 U5350 ( .A1(n4973), .A2(n4972), .ZN(n5393) );
  INV_X1 U5351 ( .A(n5411), .ZN(n4973) );
  NAND2_X1 U5352 ( .A1(n5192), .A2(n5191), .ZN(n5219) );
  NAND2_X1 U5353 ( .A1(n5141), .A2(n4925), .ZN(n4580) );
  INV_X1 U5354 ( .A(n8908), .ZN(n8160) );
  AND2_X1 U5355 ( .A1(n4796), .A2(n8128), .ZN(n4795) );
  OR2_X1 U5356 ( .A1(n8127), .A2(n8639), .ZN(n8128) );
  NAND2_X1 U5357 ( .A1(n6320), .A2(n6319), .ZN(n8184) );
  INV_X1 U5358 ( .A(n8904), .ZN(n6316) );
  NAND2_X1 U5359 ( .A1(n6286), .A2(n6285), .ZN(n8225) );
  AND4_X1 U5360 ( .A1(n6237), .A2(n6236), .A3(n6235), .A4(n6234), .ZN(n8777)
         );
  NAND2_X1 U5361 ( .A1(n5872), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4530) );
  INV_X1 U5362 ( .A(n7258), .ZN(n8533) );
  INV_X1 U5363 ( .A(n4721), .ZN(n7041) );
  OR2_X1 U5364 ( .A1(n7473), .A2(n7474), .ZN(n4660) );
  XNOR2_X1 U5365 ( .A(n5931), .B(n7481), .ZN(n7473) );
  OR2_X2 U5366 ( .A1(n6738), .A2(n6039), .ZN(n8621) );
  NOR2_X1 U5367 ( .A1(n9800), .A2(n5990), .ZN(n8612) );
  AOI21_X1 U5368 ( .B1(n9796), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n8626), .ZN(
        n4553) );
  INV_X1 U5369 ( .A(n8629), .ZN(n4554) );
  NAND2_X1 U5370 ( .A1(n4719), .A2(n5991), .ZN(n4473) );
  NOR2_X1 U5371 ( .A1(n8613), .A2(n5955), .ZN(n5959) );
  XNOR2_X1 U5372 ( .A(n4469), .B(n8643), .ZN(n4471) );
  INV_X1 U5373 ( .A(n8938), .ZN(n7590) );
  INV_X1 U5374 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n8947) );
  NAND3_X1 U5375 ( .A1(n4801), .A2(n4800), .A3(n4802), .ZN(n6405) );
  OAI22_X1 U5376 ( .A1(n6058), .A2(n4803), .B1(n5837), .B2(
        P2_IR_REG_31__SCAN_IN), .ZN(n4802) );
  XNOR2_X1 U5377 ( .A(n5892), .B(n5891), .ZN(n7048) );
  INV_X1 U5378 ( .A(n9318), .ZN(n9476) );
  NAND2_X1 U5379 ( .A1(n5320), .A2(n5319), .ZN(n7628) );
  INV_X1 U5380 ( .A(n9556), .ZN(n9303) );
  NAND2_X1 U5381 ( .A1(n7917), .A2(n7928), .ZN(n7918) );
  NOR2_X1 U5382 ( .A1(n7916), .A2(n7915), .ZN(n7917) );
  NAND2_X1 U5383 ( .A1(n4909), .A2(n7927), .ZN(n4905) );
  AND2_X1 U5384 ( .A1(n6537), .A2(n6515), .ZN(n9712) );
  NAND2_X1 U5385 ( .A1(n4835), .A2(n5768), .ZN(n9241) );
  OAI22_X1 U5386 ( .A1(n5145), .A2(n6489), .B1(n5038), .B2(n6540), .ZN(n5054)
         );
  NAND2_X1 U5387 ( .A1(n4646), .A2(n4642), .ZN(n6468) );
  NAND2_X1 U5388 ( .A1(n8089), .A2(n9746), .ZN(n4646) );
  NOR2_X1 U5389 ( .A1(n8087), .A2(n4643), .ZN(n4642) );
  AND2_X1 U5390 ( .A1(n5489), .A2(n5488), .ZN(n9566) );
  AOI21_X1 U5391 ( .B1(n4595), .B2(n8373), .A(n8454), .ZN(n8372) );
  NAND2_X1 U5392 ( .A1(n8377), .A2(n8532), .ZN(n4595) );
  INV_X1 U5393 ( .A(n7707), .ZN(n7708) );
  AOI21_X1 U5394 ( .B1(n4612), .B2(n8486), .A(n4611), .ZN(n4610) );
  INV_X1 U5395 ( .A(n8400), .ZN(n4611) );
  INV_X1 U5396 ( .A(n8795), .ZN(n4609) );
  INV_X1 U5397 ( .A(n4588), .ZN(n4587) );
  AOI21_X1 U5398 ( .B1(n4586), .B2(n4585), .A(n4583), .ZN(n4582) );
  NAND2_X1 U5399 ( .A1(n4510), .A2(n7767), .ZN(n4509) );
  OAI21_X1 U5400 ( .B1(n7765), .B2(n4629), .A(n7961), .ZN(n4510) );
  NOR2_X1 U5401 ( .A1(n7965), .A2(n7838), .ZN(n4508) );
  NAND2_X1 U5402 ( .A1(n4613), .A2(n8424), .ZN(n8430) );
  NAND2_X1 U5403 ( .A1(n8412), .A2(n4615), .ZN(n4614) );
  INV_X1 U5404 ( .A(n7783), .ZN(n4526) );
  NAND2_X1 U5405 ( .A1(n4524), .A2(n4519), .ZN(n4518) );
  NAND2_X1 U5406 ( .A1(n4365), .A2(n4449), .ZN(n4519) );
  INV_X1 U5407 ( .A(n4525), .ZN(n4524) );
  OAI211_X1 U5408 ( .C1(n4527), .C2(n7930), .A(n4419), .B(n4526), .ZN(n4525)
         );
  OR2_X1 U5409 ( .A1(n7782), .A2(n4520), .ZN(n4516) );
  NOR2_X1 U5410 ( .A1(n4365), .A2(n4521), .ZN(n4520) );
  INV_X1 U5411 ( .A(n4527), .ZN(n4521) );
  NOR2_X1 U5412 ( .A1(n7786), .A2(n4523), .ZN(n4522) );
  INV_X1 U5413 ( .A(n5620), .ZN(n4916) );
  NOR2_X1 U5414 ( .A1(n8779), .A2(n4701), .ZN(n4700) );
  AND2_X1 U5415 ( .A1(n8795), .A2(n4702), .ZN(n4701) );
  INV_X1 U5416 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5873) );
  AOI21_X1 U5417 ( .B1(n7893), .B2(n7892), .A(n7891), .ZN(n7894) );
  AND2_X1 U5418 ( .A1(n4387), .A2(n7806), .ZN(n7807) );
  AOI21_X1 U5419 ( .B1(n4494), .B2(n4401), .A(n4487), .ZN(n7804) );
  OAI21_X1 U5420 ( .B1(n4491), .B2(n4489), .A(n4488), .ZN(n4487) );
  OR2_X1 U5421 ( .A1(n9275), .A2(n9260), .ZN(n9245) );
  AND2_X1 U5422 ( .A1(n9345), .A2(n4570), .ZN(n9274) );
  NOR2_X1 U5423 ( .A1(n9294), .A2(n4571), .ZN(n4570) );
  INV_X1 U5424 ( .A(n4572), .ZN(n4571) );
  NOR2_X1 U5425 ( .A1(n4573), .A2(n9303), .ZN(n4572) );
  INV_X1 U5426 ( .A(n4574), .ZN(n4573) );
  NOR2_X1 U5427 ( .A1(n9358), .A2(n9363), .ZN(n9344) );
  NOR2_X1 U5428 ( .A1(n9399), .A2(n4567), .ZN(n4566) );
  INV_X1 U5429 ( .A(n4568), .ZN(n4567) );
  NOR2_X1 U5430 ( .A1(n9514), .A2(n9425), .ZN(n4568) );
  NOR2_X1 U5431 ( .A1(n4912), .A2(n4916), .ZN(n4911) );
  INV_X1 U5432 ( .A(n5600), .ZN(n4912) );
  OAI21_X1 U5433 ( .B1(n5618), .B2(n4916), .A(n5633), .ZN(n4915) );
  NAND2_X1 U5434 ( .A1(n5464), .A2(SI_18_), .ZN(n5465) );
  INV_X1 U5435 ( .A(SI_9_), .ZN(n9991) );
  NAND2_X1 U5436 ( .A1(n7507), .A2(n7506), .ZN(n7559) );
  INV_X1 U5437 ( .A(n6453), .ZN(n6445) );
  INV_X1 U5438 ( .A(n8148), .ZN(n4775) );
  NOR2_X1 U5439 ( .A1(n8498), .A2(n4882), .ZN(n4881) );
  INV_X1 U5440 ( .A(n4883), .ZN(n4882) );
  AOI21_X1 U5441 ( .B1(n8805), .B2(n8880), .A(n4884), .ZN(n4883) );
  INV_X1 U5442 ( .A(n8452), .ZN(n4884) );
  NAND2_X1 U5443 ( .A1(n8451), .A2(n8450), .ZN(n8500) );
  NAND2_X1 U5444 ( .A1(n5966), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5967) );
  NAND2_X1 U5445 ( .A1(n6692), .A2(n4394), .ZN(n4535) );
  NOR2_X1 U5446 ( .A1(n5914), .A2(n5972), .ZN(n5973) );
  INV_X1 U5447 ( .A(n6022), .ZN(n4544) );
  INV_X1 U5448 ( .A(n7479), .ZN(n4541) );
  NOR2_X1 U5449 ( .A1(n8602), .A2(n4475), .ZN(n5948) );
  NOR2_X1 U5450 ( .A1(n8599), .A2(n5945), .ZN(n4475) );
  NAND2_X1 U5451 ( .A1(n7019), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n4709) );
  AND2_X1 U5452 ( .A1(n9804), .A2(n4528), .ZN(n6036) );
  NAND2_X1 U5453 ( .A1(n6034), .A2(n6239), .ZN(n4528) );
  NOR2_X1 U5454 ( .A1(n8656), .A2(n4868), .ZN(n4867) );
  INV_X1 U5455 ( .A(n8440), .ZN(n4868) );
  INV_X1 U5456 ( .A(n4870), .ZN(n4865) );
  NAND2_X1 U5457 ( .A1(n4898), .A2(n8713), .ZN(n4896) );
  INV_X1 U5458 ( .A(n4690), .ZN(n4689) );
  NAND2_X1 U5459 ( .A1(n8160), .A2(n8523), .ZN(n4695) );
  NAND2_X1 U5460 ( .A1(n6278), .A2(n10000), .ZN(n6287) );
  INV_X1 U5461 ( .A(n4700), .ZN(n4699) );
  INV_X1 U5462 ( .A(n8398), .ZN(n4875) );
  OR2_X1 U5463 ( .A1(n6218), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6220) );
  OAI21_X1 U5464 ( .B1(n4389), .B2(n7996), .A(n8531), .ZN(n4673) );
  AND2_X1 U5465 ( .A1(n8479), .A2(n4676), .ZN(n4675) );
  INV_X1 U5466 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n6168) );
  NAND2_X1 U5467 ( .A1(n6154), .A2(n8473), .ZN(n7124) );
  INV_X1 U5468 ( .A(n6177), .ZN(n6154) );
  OR2_X1 U5469 ( .A1(n7297), .A2(n6177), .ZN(n7125) );
  NAND2_X1 U5470 ( .A1(n4861), .A2(n4860), .ZN(n8325) );
  NAND2_X1 U5471 ( .A1(n6383), .A2(n6836), .ZN(n6872) );
  NAND2_X1 U5472 ( .A1(n6872), .A2(n8467), .ZN(n6874) );
  INV_X1 U5473 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5951) );
  NOR2_X1 U5474 ( .A1(n5876), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n4770) );
  INV_X1 U5475 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5938) );
  OR2_X1 U5476 ( .A1(n5888), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n5916) );
  INV_X1 U5477 ( .A(n9027), .ZN(n4756) );
  NOR2_X1 U5478 ( .A1(n4838), .A2(n4834), .ZN(n4833) );
  INV_X1 U5479 ( .A(n4843), .ZN(n4834) );
  INV_X1 U5480 ( .A(n4839), .ZN(n4838) );
  NOR2_X1 U5481 ( .A1(n9225), .A2(n4846), .ZN(n4839) );
  AND2_X1 U5482 ( .A1(n9225), .A2(n4637), .ZN(n4636) );
  OR2_X1 U5483 ( .A1(n9242), .A2(n4638), .ZN(n4637) );
  NAND2_X1 U5484 ( .A1(n9253), .A2(n7889), .ZN(n7868) );
  NAND2_X1 U5485 ( .A1(n4625), .A2(n7787), .ZN(n4624) );
  INV_X1 U5486 ( .A(n9320), .ZN(n4625) );
  INV_X1 U5487 ( .A(n7792), .ZN(n4622) );
  NOR2_X1 U5488 ( .A1(n9476), .A2(n9336), .ZN(n4574) );
  OR2_X1 U5489 ( .A1(n9363), .A2(n9375), .ZN(n7967) );
  AOI21_X1 U5490 ( .B1(n4824), .B2(n9385), .A(n4830), .ZN(n4822) );
  AOI21_X1 U5491 ( .B1(n5798), .B2(n9409), .A(n4631), .ZN(n4630) );
  INV_X1 U5492 ( .A(n7762), .ZN(n4631) );
  INV_X1 U5493 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5370) );
  NAND2_X1 U5494 ( .A1(n5797), .A2(n7956), .ZN(n9411) );
  INV_X1 U5495 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5321) );
  NOR2_X1 U5496 ( .A1(n5322), .A2(n5321), .ZN(n5343) );
  OR2_X1 U5497 ( .A1(n5791), .A2(n7107), .ZN(n7950) );
  INV_X1 U5498 ( .A(n9548), .ZN(n9277) );
  AND2_X1 U5499 ( .A1(n9344), .A2(n9349), .ZN(n9345) );
  NAND2_X1 U5500 ( .A1(n7536), .A2(n4566), .ZN(n9397) );
  AND3_X1 U5501 ( .A1(n4371), .A2(n7608), .A3(n7210), .ZN(n7464) );
  OR2_X1 U5502 ( .A1(n7817), .A2(n7816), .ZN(n7818) );
  INV_X1 U5503 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n4859) );
  INV_X1 U5504 ( .A(n4858), .ZN(n4856) );
  AND2_X1 U5505 ( .A1(n5772), .A2(n5665), .ZN(n5770) );
  NAND2_X1 U5506 ( .A1(n4427), .A2(n4979), .ZN(n4563) );
  NOR2_X1 U5507 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n4953) );
  AOI21_X1 U5508 ( .B1(n4921), .B2(n4920), .A(n4448), .ZN(n4919) );
  INV_X1 U5509 ( .A(n4384), .ZN(n4920) );
  NOR2_X1 U5510 ( .A1(n5438), .A2(n5437), .ZN(n5440) );
  INV_X1 U5511 ( .A(n5115), .ZN(n4925) );
  INV_X1 U5512 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4995) );
  INV_X1 U5513 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4994) );
  INV_X1 U5514 ( .A(SI_13_), .ZN(n10110) );
  AOI21_X1 U5515 ( .B1(n4807), .B2(n6898), .A(n4374), .ZN(n4805) );
  INV_X1 U5516 ( .A(n4807), .ZN(n4806) );
  NAND2_X1 U5517 ( .A1(n4428), .A2(n8259), .ZN(n4799) );
  NAND2_X1 U5518 ( .A1(n4775), .A2(n8093), .ZN(n4774) );
  XNOR2_X1 U5519 ( .A(n9827), .B(n4361), .ZN(n6805) );
  XNOR2_X1 U5520 ( .A(n4350), .B(n6993), .ZN(n6817) );
  NOR2_X1 U5521 ( .A1(n4797), .A2(n4793), .ZN(n4792) );
  INV_X1 U5522 ( .A(n8120), .ZN(n4793) );
  OR2_X1 U5523 ( .A1(n4797), .A2(n4390), .ZN(n4796) );
  CLKBUF_X1 U5524 ( .A(n7250), .Z(n7247) );
  NOR2_X1 U5525 ( .A1(n6145), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6159) );
  INV_X1 U5526 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n10098) );
  AND2_X1 U5527 ( .A1(n6159), .A2(n10098), .ZN(n6169) );
  NAND2_X1 U5528 ( .A1(n6787), .A2(n6788), .ZN(n6790) );
  OR2_X1 U5529 ( .A1(n8109), .A2(n6274), .ZN(n4946) );
  NOR2_X1 U5530 ( .A1(n6220), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6230) );
  INV_X1 U5531 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n6123) );
  AOI21_X1 U5532 ( .B1(n4786), .B2(n4781), .A(n4780), .ZN(n4779) );
  NOR2_X1 U5533 ( .A1(n8112), .A2(n8524), .ZN(n4780) );
  NAND2_X1 U5534 ( .A1(n8214), .A2(n8213), .ZN(n8212) );
  AND2_X1 U5535 ( .A1(n6269), .A2(n10064), .ZN(n6278) );
  INV_X1 U5536 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n10064) );
  OR2_X1 U5537 ( .A1(n4790), .A2(n4395), .ZN(n4787) );
  OR2_X1 U5538 ( .A1(n4788), .A2(n4395), .ZN(n4786) );
  INV_X1 U5539 ( .A(n4789), .ZN(n4788) );
  OAI21_X1 U5540 ( .B1(n8213), .B2(n4790), .A(n8172), .ZN(n4789) );
  CLKBUF_X1 U5541 ( .A(n7559), .Z(n7505) );
  NAND2_X1 U5542 ( .A1(n5852), .A2(n4903), .ZN(n4902) );
  NOR2_X1 U5543 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n4903) );
  OAI21_X1 U5544 ( .B1(n5966), .B2(n5906), .A(n5905), .ZN(n6652) );
  INV_X1 U5545 ( .A(n6472), .ZN(n4547) );
  NOR2_X1 U5546 ( .A1(n4551), .A2(n4550), .ZN(n4549) );
  INV_X1 U5547 ( .A(n6499), .ZN(n4550) );
  AND2_X1 U5548 ( .A1(n4664), .A2(n4665), .ZN(n9766) );
  NOR2_X1 U5549 ( .A1(n4539), .A2(n6493), .ZN(n4538) );
  NOR2_X1 U5550 ( .A1(n9785), .A2(n9786), .ZN(n9784) );
  NAND2_X1 U5551 ( .A1(n4663), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n4662) );
  INV_X1 U5552 ( .A(n6757), .ZN(n4663) );
  NAND2_X1 U5553 ( .A1(n7048), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n4720) );
  OAI21_X1 U5554 ( .B1(n7478), .B2(n4542), .A(n4540), .ZN(n8548) );
  INV_X1 U5555 ( .A(n4543), .ZN(n4542) );
  AOI21_X1 U5556 ( .B1(n4541), .B2(n4543), .A(n7649), .ZN(n4540) );
  NOR2_X1 U5557 ( .A1(n7648), .A2(n4544), .ZN(n4543) );
  NAND2_X1 U5558 ( .A1(n4712), .A2(n4711), .ZN(n4710) );
  INV_X1 U5559 ( .A(n8592), .ZN(n4711) );
  AOI21_X1 U5560 ( .B1(n8617), .B2(n8616), .A(n9810), .ZN(n8629) );
  OR2_X1 U5561 ( .A1(n6355), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n7698) );
  AND4_X1 U5562 ( .A1(n6360), .A2(n6359), .A3(n6358), .A4(n6357), .ZN(n8650)
         );
  NOR2_X1 U5563 ( .A1(n6296), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6306) );
  AND2_X1 U5564 ( .A1(n8420), .A2(n8411), .ZN(n8725) );
  OR2_X1 U5565 ( .A1(n6250), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6261) );
  AND2_X1 U5566 ( .A1(n8414), .A2(n8413), .ZN(n8749) );
  NOR2_X1 U5567 ( .A1(n6201), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6209) );
  INV_X1 U5568 ( .A(n8531), .ZN(n7561) );
  OR2_X1 U5569 ( .A1(n6190), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6201) );
  NOR2_X1 U5570 ( .A1(n4891), .A2(n4888), .ZN(n4887) );
  OAI21_X1 U5571 ( .B1(n4889), .B2(n4888), .A(n8357), .ZN(n4886) );
  INV_X1 U5572 ( .A(n8354), .ZN(n4888) );
  INV_X1 U5573 ( .A(n4389), .ZN(n4670) );
  AND2_X1 U5574 ( .A1(n4677), .A2(n8479), .ZN(n4671) );
  NAND2_X1 U5575 ( .A1(n6169), .A2(n6168), .ZN(n6182) );
  OR2_X1 U5576 ( .A1(n6182), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6190) );
  INV_X1 U5577 ( .A(n4470), .ZN(n7199) );
  NAND2_X1 U5578 ( .A1(n4468), .A2(n7129), .ZN(n7197) );
  INV_X1 U5579 ( .A(n7125), .ZN(n4468) );
  OAI21_X1 U5580 ( .B1(n7227), .B2(n6387), .A(n8347), .ZN(n7295) );
  INV_X1 U5581 ( .A(n7301), .ZN(n8475) );
  OR2_X1 U5582 ( .A1(n6143), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6145) );
  INV_X1 U5583 ( .A(n4704), .ZN(n4703) );
  OAI21_X1 U5584 ( .B1(n6103), .B2(n4706), .A(n6112), .ZN(n4704) );
  NAND2_X1 U5585 ( .A1(n8338), .A2(n8332), .ZN(n6987) );
  NAND2_X1 U5586 ( .A1(n6878), .A2(n6103), .ZN(n6988) );
  AND2_X1 U5587 ( .A1(n6427), .A2(n6614), .ZN(n6848) );
  AND2_X1 U5588 ( .A1(n6455), .A2(n6454), .ZN(n6849) );
  XNOR2_X1 U5589 ( .A(n4685), .B(n6378), .ZN(n6381) );
  OAI21_X1 U5590 ( .B1(n6350), .B2(n4682), .A(n4680), .ZN(n4685) );
  AOI21_X1 U5591 ( .B1(n4683), .B2(n4681), .A(n4416), .ZN(n4680) );
  NAND2_X1 U5592 ( .A1(n6268), .A2(n6267), .ZN(n8107) );
  NAND2_X1 U5593 ( .A1(n6055), .A2(n6054), .ZN(n8098) );
  NAND2_X1 U5594 ( .A1(n6207), .A2(n6206), .ZN(n8388) );
  NOR2_X1 U5595 ( .A1(n6441), .A2(n8466), .ZN(n6726) );
  AND2_X1 U5596 ( .A1(n6747), .A2(n6746), .ZN(n6727) );
  AND2_X1 U5597 ( .A1(n6741), .A2(n6746), .ZN(n6732) );
  INV_X1 U5598 ( .A(n6443), .ZN(n6998) );
  INV_X1 U5599 ( .A(n9861), .ZN(n9871) );
  INV_X1 U5600 ( .A(n7003), .ZN(n6645) );
  XNOR2_X1 U5601 ( .A(n5861), .B(n5862), .ZN(n6737) );
  INV_X1 U5602 ( .A(n5865), .ZN(n4531) );
  INV_X1 U5603 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n4901) );
  AND2_X1 U5604 ( .A1(n5956), .A2(n5837), .ZN(n4804) );
  NOR2_X1 U5605 ( .A1(n5956), .A2(n5837), .ZN(n4803) );
  NOR2_X1 U5606 ( .A1(n5834), .A2(P2_IR_REG_10__SCAN_IN), .ZN(n4778) );
  INV_X1 U5607 ( .A(n5888), .ZN(n4777) );
  OR2_X1 U5608 ( .A1(n5893), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n5890) );
  XNOR2_X1 U5609 ( .A(n5894), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6139) );
  NOR2_X1 U5610 ( .A1(n5916), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n5920) );
  INV_X1 U5611 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5921) );
  INV_X1 U5612 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n4708) );
  NAND2_X1 U5613 ( .A1(n6058), .A2(n5828), .ZN(n5902) );
  NAND2_X1 U5614 ( .A1(n5357), .A2(n5356), .ZN(n8963) );
  INV_X1 U5615 ( .A(n5608), .ZN(n5607) );
  AND2_X1 U5616 ( .A1(n5658), .A2(n5657), .ZN(n5681) );
  OR2_X1 U5617 ( .A1(n5182), .A2(n6982), .ZN(n5210) );
  INV_X1 U5618 ( .A(n8971), .ZN(n4750) );
  INV_X1 U5619 ( .A(n4758), .ZN(n4757) );
  OAI21_X1 U5620 ( .B1(n4382), .B2(n4759), .A(n5436), .ZN(n4758) );
  NOR2_X1 U5621 ( .A1(n5432), .A2(n4760), .ZN(n4759) );
  NOR2_X1 U5622 ( .A1(n5238), .A2(n5237), .ZN(n5264) );
  AND2_X1 U5623 ( .A1(n5540), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n5566) );
  NAND2_X1 U5624 ( .A1(n4735), .A2(n4411), .ZN(n9071) );
  INV_X1 U5625 ( .A(n4444), .ZN(n4734) );
  NAND2_X1 U5626 ( .A1(n7597), .A2(n7599), .ZN(n7596) );
  OR2_X1 U5627 ( .A1(n5301), .A2(n7602), .ZN(n5322) );
  INV_X1 U5628 ( .A(n6465), .ZN(n6623) );
  INV_X1 U5629 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n9083) );
  INV_X1 U5630 ( .A(n4745), .ZN(n4744) );
  AOI21_X1 U5631 ( .B1(n4746), .B2(n4753), .A(n5655), .ZN(n4745) );
  NAND2_X1 U5632 ( .A1(n4495), .A2(n4496), .ZN(n7921) );
  AND2_X1 U5633 ( .A1(n4499), .A2(n4497), .ZN(n4496) );
  NOR2_X1 U5634 ( .A1(n4412), .A2(n4504), .ZN(n4499) );
  AND4_X1 U5635 ( .A1(n5674), .A2(n5673), .A3(n5672), .A4(n5671), .ZN(n5818)
         );
  AND4_X1 U5636 ( .A1(n5631), .A2(n5630), .A3(n5629), .A4(n5628), .ZN(n9093)
         );
  AOI21_X1 U5637 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(n9601), .A(n9593), .ZN(
        n9635) );
  AOI21_X1 U5638 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n9653), .A(n9648), .ZN(
        n9659) );
  NOR2_X1 U5639 ( .A1(n8005), .A2(n9673), .ZN(n9689) );
  NOR2_X1 U5640 ( .A1(n8068), .A2(n4351), .ZN(n4558) );
  INV_X1 U5641 ( .A(n4558), .ZN(n9209) );
  NAND2_X1 U5642 ( .A1(n8055), .A2(n8054), .ZN(n8062) );
  OR2_X1 U5643 ( .A1(n8055), .A2(n8054), .ZN(n8060) );
  AND2_X1 U5644 ( .A1(n8060), .A2(n8062), .ZN(n7872) );
  AND2_X1 U5645 ( .A1(n5813), .A2(n5670), .ZN(n9232) );
  AOI21_X1 U5646 ( .B1(n4854), .B2(n4399), .A(n4848), .ZN(n9267) );
  OAI21_X1 U5647 ( .B1(n4850), .B2(n4849), .A(n4402), .ZN(n4848) );
  NAND2_X1 U5648 ( .A1(n4623), .A2(n4621), .ZN(n9285) );
  AOI21_X1 U5649 ( .B1(n4386), .B2(n4626), .A(n4622), .ZN(n4621) );
  NAND2_X1 U5650 ( .A1(n9321), .A2(n4386), .ZN(n4623) );
  INV_X1 U5651 ( .A(n7787), .ZN(n4626) );
  AND4_X1 U5652 ( .A1(n5612), .A2(n5611), .A3(n5610), .A4(n5609), .ZN(n9002)
         );
  NAND2_X1 U5653 ( .A1(n9345), .A2(n4574), .ZN(n9313) );
  NAND2_X1 U5654 ( .A1(n9345), .A2(n9561), .ZN(n9333) );
  OR2_X1 U5655 ( .A1(n5490), .A2(n9083), .ZN(n5492) );
  OR2_X1 U5656 ( .A1(n5492), .A2(n8987), .ZN(n5521) );
  INV_X1 U5657 ( .A(n9124), .ZN(n9343) );
  AND2_X1 U5658 ( .A1(n7967), .A2(n7781), .ZN(n9353) );
  NAND2_X1 U5659 ( .A1(n9031), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n5490) );
  INV_X1 U5660 ( .A(n4831), .ZN(n4829) );
  OR2_X1 U5661 ( .A1(n5371), .A2(n5370), .ZN(n5416) );
  NAND2_X1 U5662 ( .A1(n9411), .A2(n4826), .ZN(n9410) );
  NAND2_X1 U5663 ( .A1(n7536), .A2(n4832), .ZN(n9421) );
  OR2_X1 U5664 ( .A1(n7446), .A2(n9131), .ZN(n5752) );
  OR2_X1 U5665 ( .A1(n7157), .A2(n9133), .ZN(n5749) );
  NAND2_X1 U5666 ( .A1(n7210), .A2(n4362), .ZN(n7332) );
  AOI21_X1 U5667 ( .B1(n4817), .B2(n4819), .A(n4421), .ZN(n4815) );
  NAND2_X1 U5668 ( .A1(n7210), .A2(n7309), .ZN(n7211) );
  NOR2_X1 U5669 ( .A1(n4577), .A2(n7094), .ZN(n7180) );
  NOR2_X1 U5670 ( .A1(n7098), .A2(n7727), .ZN(n4575) );
  OR2_X1 U5671 ( .A1(n9742), .A2(n7924), .ZN(n5825) );
  AND2_X1 U5672 ( .A1(n5726), .A2(n6508), .ZN(n9390) );
  NAND2_X1 U5673 ( .A1(n4578), .A2(n4364), .ZN(n6965) );
  NOR2_X1 U5674 ( .A1(n7094), .A2(n7098), .ZN(n7095) );
  NAND2_X1 U5675 ( .A1(n7933), .A2(n7936), .ZN(n7707) );
  AND4_X1 U5676 ( .A1(n5103), .A2(n5102), .A3(n5101), .A4(n5100), .ZN(n7090)
         );
  NAND2_X1 U5677 ( .A1(n7933), .A2(n4650), .ZN(n7087) );
  NAND2_X1 U5678 ( .A1(n7065), .A2(n5738), .ZN(n5739) );
  NAND2_X1 U5679 ( .A1(n4620), .A2(n5785), .ZN(n6669) );
  INV_X1 U5680 ( .A(n9393), .ZN(n9412) );
  INV_X1 U5681 ( .A(n9390), .ZN(n9414) );
  AND2_X1 U5682 ( .A1(n9205), .A2(n9204), .ZN(n9438) );
  INV_X1 U5683 ( .A(n8082), .ZN(n4644) );
  NAND2_X1 U5684 ( .A1(n5467), .A2(n5466), .ZN(n9491) );
  OR2_X1 U5685 ( .A1(n7919), .A2(n7982), .ZN(n9742) );
  AND2_X1 U5686 ( .A1(n5812), .A2(n5811), .ZN(n9496) );
  INV_X1 U5687 ( .A(n9734), .ZN(n9516) );
  AND2_X1 U5688 ( .A1(n6623), .A2(n6464), .ZN(n7006) );
  INV_X1 U5689 ( .A(n7013), .ZN(n7071) );
  NAND2_X1 U5690 ( .A1(n9741), .A2(n9742), .ZN(n9734) );
  NAND2_X1 U5691 ( .A1(n5700), .A2(n5689), .ZN(n9577) );
  AND2_X1 U5692 ( .A1(n5600), .A2(n5579), .ZN(n5598) );
  XNOR2_X1 U5693 ( .A(n5710), .B(n5709), .ZN(n6507) );
  INV_X1 U5694 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5709) );
  OAI21_X1 U5695 ( .B1(n4977), .B2(n5297), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5707) );
  INV_X1 U5696 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5706) );
  AND2_X1 U5697 ( .A1(n5339), .A2(n5318), .ZN(n8014) );
  NAND2_X1 U5698 ( .A1(n4937), .A2(n4938), .ZN(n5337) );
  NAND2_X1 U5699 ( .A1(n5289), .A2(n4940), .ZN(n4937) );
  OAI21_X1 U5700 ( .B1(n5289), .B2(n5288), .A(n5292), .ZN(n5315) );
  XNOR2_X1 U5701 ( .A(n5289), .B(n5287), .ZN(n6593) );
  NAND2_X1 U5702 ( .A1(n4579), .A2(n5169), .ZN(n5189) );
  NAND2_X1 U5703 ( .A1(n5090), .A2(n5089), .ZN(n5113) );
  XNOR2_X1 U5704 ( .A(n5114), .B(n5085), .ZN(n5112) );
  XNOR2_X1 U5705 ( .A(n5057), .B(n5002), .ZN(n5056) );
  NAND2_X1 U5706 ( .A1(n4794), .A2(n4799), .ZN(n8140) );
  NAND2_X1 U5707 ( .A1(n8179), .A2(n4390), .ZN(n4794) );
  XNOR2_X1 U5708 ( .A(n8127), .B(n8639), .ZN(n8141) );
  AND4_X1 U5709 ( .A1(n6070), .A2(n6069), .A3(n6068), .A4(n6067), .ZN(n8791)
         );
  NAND2_X1 U5710 ( .A1(n4773), .A2(n4774), .ZN(n8150) );
  NAND2_X1 U5711 ( .A1(n8212), .A2(n4946), .ZN(n8173) );
  NAND2_X1 U5712 ( .A1(n6277), .A2(n6276), .ZN(n8727) );
  XNOR2_X1 U5713 ( .A(n8118), .B(n8700), .ZN(n8206) );
  CLKBUF_X1 U5714 ( .A(n6894), .Z(n6825) );
  AND2_X1 U5715 ( .A1(n7370), .A2(n7367), .ZN(n4776) );
  AND2_X1 U5716 ( .A1(n7368), .A2(n7367), .ZN(n7371) );
  AND3_X1 U5717 ( .A1(n6265), .A2(n6264), .A3(n6263), .ZN(n8736) );
  AND4_X1 U5718 ( .A1(n6224), .A2(n6223), .A3(n6222), .A4(n6221), .ZN(n8096)
         );
  OAI21_X1 U5719 ( .B1(n8214), .B2(n4787), .A(n4786), .ZN(n8220) );
  NAND2_X1 U5720 ( .A1(n6249), .A2(n6248), .ZN(n8243) );
  AND2_X1 U5721 ( .A1(n7238), .A2(n7237), .ZN(n8248) );
  INV_X1 U5722 ( .A(n8279), .ZN(n8265) );
  AND2_X1 U5723 ( .A1(n4772), .A2(n8275), .ZN(n4771) );
  AND2_X1 U5724 ( .A1(n4773), .A2(n4772), .ZN(n8276) );
  INV_X1 U5725 ( .A(n8271), .ZN(n8273) );
  INV_X1 U5726 ( .A(n8267), .ZN(n8281) );
  NOR2_X1 U5727 ( .A1(n4363), .A2(n6421), .ZN(n4601) );
  OAI21_X1 U5728 ( .B1(n8513), .B2(n4363), .A(n4413), .ZN(n4598) );
  NOR2_X1 U5729 ( .A1(n4949), .A2(n6421), .ZN(n4603) );
  XNOR2_X1 U5730 ( .A(n5864), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8516) );
  INV_X1 U5731 ( .A(n8711), .ZN(n8523) );
  INV_X1 U5732 ( .A(n8736), .ZN(n8764) );
  AND4_X1 U5733 ( .A1(n6247), .A2(n6246), .A3(n6245), .A4(n6244), .ZN(n8789)
         );
  INV_X1 U5734 ( .A(n7992), .ZN(n8530) );
  OR2_X1 U5735 ( .A1(n4359), .A2(n5972), .ZN(n6116) );
  OR2_X1 U5736 ( .A1(n6091), .A2(n6081), .ZN(n6083) );
  INV_X1 U5737 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n9763) );
  XNOR2_X1 U5738 ( .A(n6005), .B(n6499), .ZN(n6473) );
  NOR2_X1 U5739 ( .A1(n6473), .A2(n6472), .ZN(n6471) );
  OAI21_X1 U5740 ( .B1(n6473), .B2(n4546), .A(n4545), .ZN(n6659) );
  NAND2_X1 U5741 ( .A1(n4549), .A2(n4548), .ZN(n4545) );
  NAND2_X1 U5742 ( .A1(n4548), .A2(n4547), .ZN(n4546) );
  INV_X1 U5743 ( .A(n6661), .ZN(n4548) );
  NOR2_X1 U5744 ( .A1(n6471), .A2(n4549), .ZN(n6660) );
  NAND2_X1 U5745 ( .A1(n4666), .A2(n4664), .ZN(n9767) );
  NAND2_X1 U5746 ( .A1(n6691), .A2(n6010), .ZN(n9782) );
  INV_X1 U5747 ( .A(n4667), .ZN(n5928) );
  INV_X1 U5748 ( .A(n4715), .ZN(n7418) );
  INV_X1 U5749 ( .A(n4713), .ZN(n7416) );
  NOR2_X1 U5750 ( .A1(n5985), .A2(n7475), .ZN(n7647) );
  NAND2_X1 U5751 ( .A1(n7477), .A2(n6022), .ZN(n7650) );
  NAND2_X1 U5752 ( .A1(n4657), .A2(n4659), .ZN(n7656) );
  INV_X1 U5753 ( .A(n8558), .ZN(n4727) );
  INV_X1 U5754 ( .A(n4462), .ZN(n8574) );
  INV_X1 U5755 ( .A(n4655), .ZN(n8576) );
  INV_X1 U5756 ( .A(n4710), .ZN(n8591) );
  INV_X1 U5757 ( .A(n4712), .ZN(n8593) );
  INV_X1 U5758 ( .A(n5944), .ZN(n4654) );
  NOR2_X1 U5759 ( .A1(n4393), .A2(n4467), .ZN(n4466) );
  NAND2_X1 U5760 ( .A1(n9812), .A2(n4454), .ZN(n4467) );
  AND2_X1 U5761 ( .A1(n9801), .A2(n9802), .ZN(n4480) );
  NAND2_X1 U5762 ( .A1(n6401), .A2(n4870), .ZN(n4869) );
  NAND2_X1 U5763 ( .A1(n6401), .A2(n8434), .ZN(n8660) );
  NAND2_X1 U5764 ( .A1(n4900), .A2(n4898), .ZN(n8693) );
  NAND2_X1 U5765 ( .A1(n4687), .A2(n4690), .ZN(n8687) );
  NAND2_X1 U5766 ( .A1(n4686), .A2(n4692), .ZN(n4687) );
  NAND2_X1 U5767 ( .A1(n4686), .A2(n8713), .ZN(n4694) );
  NAND2_X1 U5768 ( .A1(n4900), .A2(n8423), .ZN(n8702) );
  AND2_X1 U5769 ( .A1(n6260), .A2(n6259), .ZN(n8753) );
  NOR2_X1 U5770 ( .A1(n8785), .A2(n6238), .ZN(n8774) );
  NAND2_X1 U5771 ( .A1(n6228), .A2(n6227), .ZN(n8857) );
  NAND2_X1 U5772 ( .A1(n4873), .A2(n4876), .ZN(n7581) );
  OR2_X1 U5773 ( .A1(n7449), .A2(n4367), .ZN(n4873) );
  OR2_X1 U5774 ( .A1(n7449), .A2(n6392), .ZN(n4877) );
  NAND2_X1 U5775 ( .A1(n4885), .A2(n4889), .ZN(n7488) );
  NAND2_X1 U5776 ( .A1(n7122), .A2(n4892), .ZN(n4885) );
  AND2_X1 U5777 ( .A1(n4678), .A2(n4677), .ZN(n7489) );
  NAND2_X1 U5778 ( .A1(n4894), .A2(n8364), .ZN(n7195) );
  NAND2_X1 U5779 ( .A1(n4895), .A2(n8363), .ZN(n4894) );
  INV_X1 U5780 ( .A(n7122), .ZN(n4895) );
  INV_X1 U5781 ( .A(n9819), .ZN(n8798) );
  INV_X1 U5782 ( .A(n8679), .ZN(n9821) );
  INV_X1 U5783 ( .A(n8350), .ZN(n9820) );
  NAND2_X1 U5784 ( .A1(n7693), .A2(n8288), .ZN(n6340) );
  AND2_X1 U5785 ( .A1(n6305), .A2(n6304), .ZN(n8904) );
  INV_X1 U5786 ( .A(n8225), .ZN(n8912) );
  INV_X1 U5787 ( .A(n8243), .ZN(n8925) );
  INV_X1 U5788 ( .A(n8202), .ZN(n8929) );
  AND2_X1 U5789 ( .A1(n6217), .A2(n6216), .ZN(n8938) );
  INV_X1 U5790 ( .A(n8388), .ZN(n8944) );
  NAND2_X1 U5791 ( .A1(n6165), .A2(n8288), .ZN(n6167) );
  OR2_X1 U5792 ( .A1(n9873), .A2(n9861), .ZN(n8943) );
  AND2_X1 U5793 ( .A1(n6737), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6619) );
  NAND2_X1 U5794 ( .A1(n5849), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5845) );
  OR2_X1 U5795 ( .A1(n5847), .A2(n5846), .ZN(n5848) );
  INV_X1 U5796 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7577) );
  NAND2_X1 U5797 ( .A1(n5869), .A2(n5868), .ZN(n8315) );
  XNOR2_X1 U5798 ( .A(n6380), .B(n5841), .ZN(n7426) );
  INV_X1 U5799 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6610) );
  INV_X1 U5800 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6590) );
  CLKBUF_X1 U5801 ( .A(n6003), .Z(n6499) );
  INV_X1 U5802 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n6982) );
  AND4_X1 U5803 ( .A1(n5348), .A2(n5347), .A3(n5346), .A4(n5345), .ZN(n9413)
         );
  NAND2_X1 U5804 ( .A1(n4743), .A2(n5286), .ZN(n9622) );
  NAND2_X1 U5805 ( .A1(n5236), .A2(n4764), .ZN(n7285) );
  INV_X1 U5806 ( .A(n5821), .ZN(n7072) );
  NAND2_X1 U5807 ( .A1(n4736), .A2(n5533), .ZN(n8994) );
  NAND2_X1 U5808 ( .A1(n4742), .A2(n4741), .ZN(n4736) );
  INV_X1 U5809 ( .A(n9053), .ZN(n4742) );
  OAI21_X1 U5810 ( .B1(n5357), .B2(n4382), .A(n4757), .ZN(n9029) );
  OAI21_X1 U5811 ( .B1(n8971), .B2(n9041), .A(n9040), .ZN(n9039) );
  NAND2_X1 U5812 ( .A1(n6706), .A2(n5127), .ZN(n6718) );
  AND4_X1 U5813 ( .A1(n5216), .A2(n5215), .A3(n5214), .A4(n5213), .ZN(n7385)
         );
  INV_X1 U5814 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n9054) );
  AOI21_X1 U5815 ( .B1(n4731), .B2(n4733), .A(n4380), .ZN(n4729) );
  AND4_X1 U5816 ( .A1(n5137), .A2(n5136), .A3(n5135), .A4(n5134), .ZN(n7728)
         );
  INV_X1 U5817 ( .A(n9113), .ZN(n9628) );
  AND2_X1 U5818 ( .A1(n5644), .A2(n5669), .ZN(n9243) );
  AND2_X1 U5819 ( .A1(n5729), .A2(n5714), .ZN(n9102) );
  INV_X1 U5820 ( .A(n9631), .ZN(n9109) );
  INV_X1 U5821 ( .A(n7986), .ZN(n4908) );
  AND4_X1 U5822 ( .A1(n5817), .A2(n5816), .A3(n5815), .A4(n5814), .ZN(n7812)
         );
  INV_X1 U5823 ( .A(n5818), .ZN(n9117) );
  NAND2_X1 U5824 ( .A1(n5099), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5017) );
  OR2_X1 U5825 ( .A1(n6463), .A2(n6462), .ZN(n9141) );
  AOI21_X1 U5826 ( .B1(n9192), .B2(P1_REG2_REG_4__SCAN_IN), .A(n6548), .ZN(
        n6567) );
  AOI21_X1 U5827 ( .B1(n6568), .B2(P1_REG2_REG_5__SCAN_IN), .A(n6565), .ZN(
        n6553) );
  AOI21_X1 U5828 ( .B1(P1_REG2_REG_16__SCAN_IN), .B2(n8012), .A(n9687), .ZN(
        n9695) );
  XNOR2_X1 U5829 ( .A(n4557), .B(n4556), .ZN(n9435) );
  NAND2_X1 U5830 ( .A1(n4558), .A2(n9532), .ZN(n4557) );
  NAND2_X1 U5831 ( .A1(n4840), .A2(n4845), .ZN(n9224) );
  NAND2_X1 U5832 ( .A1(n4835), .A2(n4841), .ZN(n4840) );
  NAND2_X1 U5833 ( .A1(n5641), .A2(n5640), .ZN(n9249) );
  NAND2_X1 U5834 ( .A1(n4847), .A2(n4850), .ZN(n9287) );
  NAND2_X1 U5835 ( .A1(n4854), .A2(n4851), .ZN(n4847) );
  AND2_X1 U5836 ( .A1(n4853), .A2(n4398), .ZN(n9297) );
  NAND2_X1 U5837 ( .A1(n4854), .A2(n4957), .ZN(n4853) );
  NAND2_X1 U5838 ( .A1(n9319), .A2(n7787), .ZN(n9299) );
  AND2_X1 U5839 ( .A1(n5539), .A2(n5538), .ZN(n9318) );
  INV_X1 U5841 ( .A(n9566), .ZN(n9363) );
  NAND2_X1 U5842 ( .A1(n9408), .A2(n4831), .ZN(n7664) );
  NAND2_X1 U5843 ( .A1(n5342), .A2(n5341), .ZN(n9066) );
  OAI21_X1 U5844 ( .B1(n7173), .B2(n4819), .A(n4817), .ZN(n7104) );
  NAND2_X1 U5845 ( .A1(n7174), .A2(n5746), .ZN(n7105) );
  OR2_X1 U5846 ( .A1(n6506), .A2(n5825), .ZN(n7333) );
  NAND2_X1 U5847 ( .A1(n9381), .A2(n7928), .ZN(n9360) );
  NOR2_X2 U5848 ( .A1(n9211), .A2(n7067), .ZN(n9355) );
  INV_X1 U5849 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n4640) );
  OR2_X1 U5850 ( .A1(n6524), .A2(n5111), .ZN(n5228) );
  AND2_X1 U5851 ( .A1(n9757), .A2(n9724), .ZN(n8073) );
  INV_X1 U5852 ( .A(n9757), .ZN(n9754) );
  AOI21_X1 U5853 ( .B1(n9435), .B2(n9477), .A(n9438), .ZN(n9526) );
  INV_X1 U5854 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n4479) );
  AOI211_X1 U5855 ( .C1(n9444), .C2(n9734), .A(n9443), .B(n9442), .ZN(n9533)
         );
  INV_X1 U5856 ( .A(n9249), .ZN(n9540) );
  AND2_X2 U5857 ( .A1(n5625), .A2(n5624), .ZN(n9544) );
  INV_X1 U5858 ( .A(n7628), .ZN(n5753) );
  AND2_X1 U5859 ( .A1(n9749), .A2(n9724), .ZN(n8078) );
  INV_X2 U5860 ( .A(n7292), .ZN(n7309) );
  NAND2_X1 U5861 ( .A1(n4515), .A2(n4514), .ZN(n4513) );
  INV_X1 U5862 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n4514) );
  NAND2_X1 U5863 ( .A1(n4993), .A2(n4992), .ZN(n4651) );
  AND2_X1 U5864 ( .A1(n6491), .A2(P1_U3086), .ZN(n7571) );
  INV_X1 U5865 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7516) );
  XNOR2_X1 U5866 ( .A(n5707), .B(n5706), .ZN(n7841) );
  INV_X1 U5867 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n4985) );
  OAI21_X1 U5868 ( .B1(n5393), .B2(n4366), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5483) );
  OAI21_X1 U5869 ( .B1(n5393), .B2(P1_IR_REG_16__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5442) );
  AND2_X1 U5870 ( .A1(n5367), .A2(n5411), .ZN(n9665) );
  INV_X1 U5871 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6594) );
  INV_X1 U5872 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6522) );
  OR2_X1 U5873 ( .A1(n5164), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n5194) );
  INV_X1 U5874 ( .A(n4723), .ZN(n7043) );
  NAND2_X1 U5875 ( .A1(n9809), .A2(n4464), .ZN(P2_U3199) );
  INV_X1 U5876 ( .A(n4465), .ZN(n4464) );
  OAI21_X1 U5877 ( .B1(n9800), .B2(n4480), .A(n5992), .ZN(n9809) );
  OAI21_X1 U5878 ( .B1(n9811), .B2(n9810), .A(n4466), .ZN(n4465) );
  AOI21_X1 U5879 ( .B1(n4555), .B2(n8627), .A(n4552), .ZN(n8630) );
  OAI21_X1 U5880 ( .B1(n8622), .B2(n8621), .A(n9814), .ZN(n4555) );
  AOI21_X1 U5881 ( .B1(n6050), .B2(n9807), .A(n6049), .ZN(n6051) );
  NAND2_X1 U5882 ( .A1(n4483), .A2(n4481), .ZN(P1_U3262) );
  AOI21_X1 U5883 ( .B1(n8027), .B2(n7928), .A(n4482), .ZN(n4481) );
  NAND2_X1 U5884 ( .A1(n8028), .A2(n7875), .ZN(n4483) );
  OAI21_X1 U5885 ( .B1(n9722), .B2(n7999), .A(n8029), .ZN(n4482) );
  NAND2_X1 U5886 ( .A1(n4641), .A2(n4447), .ZN(P1_U3550) );
  NAND2_X1 U5887 ( .A1(n6468), .A2(n9757), .ZN(n4641) );
  NOR2_X1 U5888 ( .A1(n9757), .A2(n4640), .ZN(n4639) );
  INV_X1 U5889 ( .A(n4477), .ZN(P1_U3518) );
  AOI21_X1 U5890 ( .B1(n6468), .B2(n9749), .A(n4478), .ZN(n4477) );
  NAND2_X1 U5891 ( .A1(n4378), .A2(n4453), .ZN(n4478) );
  NOR2_X1 U5892 ( .A1(n4415), .A2(n4370), .ZN(n6079) );
  AND2_X1 U5893 ( .A1(n7309), .A2(n7390), .ZN(n4362) );
  AND2_X1 U5894 ( .A1(n6971), .A2(n5740), .ZN(n4364) );
  NAND2_X1 U5895 ( .A1(n6383), .A2(n8320), .ZN(n4669) );
  INV_X1 U5896 ( .A(n6013), .ZN(n9795) );
  AND3_X1 U5897 ( .A1(n7966), .A2(n7919), .A3(n7967), .ZN(n4365) );
  NAND2_X1 U5898 ( .A1(n4763), .A2(n4974), .ZN(n4366) );
  NAND2_X1 U5899 ( .A1(n4512), .A2(n4515), .ZN(n5013) );
  OR2_X1 U5900 ( .A1(n6392), .A2(n7586), .ZN(n4367) );
  AND2_X1 U5901 ( .A1(n4414), .A2(n6418), .ZN(n4368) );
  AND2_X1 U5902 ( .A1(n4368), .A2(n9887), .ZN(n4369) );
  INV_X1 U5903 ( .A(n9827), .ZN(n4860) );
  NOR2_X1 U5904 ( .A1(n8291), .A2(n6497), .ZN(n4370) );
  AND2_X1 U5905 ( .A1(n4362), .A2(n5750), .ZN(n4371) );
  INV_X1 U5906 ( .A(n6238), .ZN(n4702) );
  AND2_X1 U5907 ( .A1(n8857), .A2(n8526), .ZN(n6238) );
  INV_X1 U5908 ( .A(n4842), .ZN(n4841) );
  NAND2_X1 U5909 ( .A1(n4403), .A2(n5768), .ZN(n4842) );
  AND2_X1 U5910 ( .A1(n6175), .A2(n6176), .ZN(n4372) );
  NAND2_X1 U5911 ( .A1(n6329), .A2(n6328), .ZN(n8670) );
  AND2_X1 U5912 ( .A1(n7240), .A2(n8536), .ZN(n4374) );
  AND2_X1 U5913 ( .A1(n6316), .A2(n6315), .ZN(n4375) );
  NAND2_X1 U5914 ( .A1(n8463), .A2(n8779), .ZN(n4376) );
  AND2_X1 U5915 ( .A1(n9385), .A2(n4828), .ZN(n4377) );
  INV_X2 U5916 ( .A(n9873), .ZN(n8939) );
  INV_X1 U5917 ( .A(n9409), .ZN(n4826) );
  OR2_X1 U5918 ( .A1(n8085), .A2(n9576), .ZN(n4378) );
  OR2_X1 U5919 ( .A1(n4931), .A2(n5536), .ZN(n4379) );
  AND2_X1 U5920 ( .A1(n5334), .A2(n5333), .ZN(n4380) );
  INV_X1 U5921 ( .A(n9425), .ZN(n4832) );
  INV_X1 U5922 ( .A(n7996), .ZN(n4676) );
  NAND2_X1 U5923 ( .A1(n4768), .A2(n4767), .ZN(n6819) );
  NAND2_X1 U5924 ( .A1(n6790), .A2(n6802), .ZN(n6791) );
  OR2_X1 U5925 ( .A1(P2_U3150), .A2(n6047), .ZN(n8628) );
  INV_X1 U5926 ( .A(n6405), .ZN(n6421) );
  INV_X1 U5927 ( .A(n5098), .ZN(n7837) );
  INV_X1 U5928 ( .A(n7065), .ZN(n9140) );
  AND4_X1 U5929 ( .A1(n5052), .A2(n5051), .A3(n5050), .A4(n5049), .ZN(n7065)
         );
  NAND2_X1 U5930 ( .A1(n6752), .A2(n4461), .ZN(n6383) );
  OR2_X1 U5931 ( .A1(n4962), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n4381) );
  OR2_X1 U5932 ( .A1(n5431), .A2(n5430), .ZN(n4382) );
  OR2_X1 U5933 ( .A1(n6395), .A2(n6394), .ZN(n4383) );
  AND2_X1 U5934 ( .A1(n6141), .A2(n6140), .ZN(n8350) );
  OR2_X1 U5935 ( .A1(n5439), .A2(SI_16_), .ZN(n4384) );
  NOR2_X2 U5936 ( .A1(n8163), .A2(n4956), .ZN(n8214) );
  AND2_X1 U5937 ( .A1(n5272), .A2(n5250), .ZN(n4385) );
  OAI21_X1 U5938 ( .B1(n8951), .B2(n5111), .A(n7811), .ZN(n8067) );
  AND2_X1 U5939 ( .A1(n9298), .A2(n4624), .ZN(n4386) );
  AND3_X1 U5940 ( .A1(n8062), .A2(n7799), .A3(n7919), .ZN(n4387) );
  AND2_X1 U5941 ( .A1(n4837), .A2(n4836), .ZN(n4388) );
  OR2_X1 U5942 ( .A1(n7525), .A2(n8532), .ZN(n4389) );
  INV_X1 U5943 ( .A(n7897), .ZN(n4638) );
  NAND2_X1 U5944 ( .A1(n5064), .A2(n5063), .ZN(n7142) );
  INV_X1 U5945 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5010) );
  AND2_X1 U5946 ( .A1(n8180), .A2(n8259), .ZN(n4390) );
  OR2_X1 U5947 ( .A1(n8583), .A2(n5988), .ZN(n4391) );
  AND3_X1 U5948 ( .A1(n5008), .A2(n5007), .A3(n5006), .ZN(n5821) );
  NAND2_X1 U5949 ( .A1(n4869), .A2(n8440), .ZN(n8655) );
  NAND2_X1 U5950 ( .A1(n8912), .A2(n8721), .ZN(n4392) );
  AND2_X1 U5951 ( .A1(n9808), .A2(n9807), .ZN(n4393) );
  NAND2_X1 U5952 ( .A1(n5444), .A2(n5443), .ZN(n9504) );
  INV_X1 U5953 ( .A(n9504), .ZN(n4565) );
  NAND2_X1 U5954 ( .A1(n7833), .A2(n7832), .ZN(n9203) );
  INV_X1 U5955 ( .A(n9203), .ZN(n4556) );
  INV_X1 U5956 ( .A(n8493), .ZN(n8643) );
  AND2_X1 U5957 ( .A1(n9781), .A2(n4537), .ZN(n4394) );
  NAND2_X1 U5958 ( .A1(n7821), .A2(n7820), .ZN(n9202) );
  AND2_X1 U5959 ( .A1(n8110), .A2(n8735), .ZN(n4395) );
  NOR3_X1 U5960 ( .A1(n7866), .A2(n9329), .A3(n9341), .ZN(n4396) );
  INV_X1 U5961 ( .A(n7788), .ZN(n4523) );
  AND2_X1 U5962 ( .A1(n4775), .A2(n7676), .ZN(n4397) );
  NAND2_X1 U5963 ( .A1(n4559), .A2(n4978), .ZN(n4962) );
  NAND2_X1 U5964 ( .A1(n9318), .A2(n5806), .ZN(n4398) );
  AND2_X1 U5965 ( .A1(n4851), .A2(n5764), .ZN(n4399) );
  NAND2_X1 U5966 ( .A1(n5581), .A2(n5580), .ZN(n9294) );
  AND2_X1 U5967 ( .A1(n4919), .A2(n4917), .ZN(n4400) );
  AND2_X1 U5968 ( .A1(n4492), .A2(n7881), .ZN(n4401) );
  OR2_X1 U5969 ( .A1(n9294), .A2(n9121), .ZN(n4402) );
  INV_X1 U5970 ( .A(n9336), .ZN(n9561) );
  NAND2_X1 U5971 ( .A1(n5520), .A2(n5519), .ZN(n9336) );
  OR2_X1 U5972 ( .A1(n9249), .A2(n9118), .ZN(n4403) );
  AND2_X1 U5973 ( .A1(n8463), .A2(n8407), .ZN(n4404) );
  INV_X1 U5974 ( .A(n4828), .ZN(n4827) );
  NOR2_X1 U5975 ( .A1(n5756), .A2(n4829), .ZN(n4828) );
  AND2_X1 U5976 ( .A1(n5852), .A2(n4901), .ZN(n4405) );
  INV_X1 U5977 ( .A(n9399), .ZN(n9571) );
  NAND2_X1 U5978 ( .A1(n5396), .A2(n5395), .ZN(n9399) );
  NAND2_X1 U5979 ( .A1(n5369), .A2(n5368), .ZN(n9425) );
  INV_X1 U5980 ( .A(n5762), .ZN(n4855) );
  INV_X1 U5981 ( .A(n8401), .ZN(n4612) );
  NOR2_X1 U5982 ( .A1(n8890), .A2(n8664), .ZN(n4406) );
  AND2_X1 U5983 ( .A1(n8438), .A2(n8437), .ZN(n4407) );
  INV_X1 U5984 ( .A(n4753), .ZN(n4749) );
  NAND2_X1 U5985 ( .A1(n5597), .A2(n5617), .ZN(n4753) );
  AND2_X1 U5986 ( .A1(n4490), .A2(n4491), .ZN(n4408) );
  AND2_X1 U5987 ( .A1(n8408), .A2(n8409), .ZN(n4409) );
  AND2_X1 U5988 ( .A1(n4655), .A2(n4654), .ZN(n4410) );
  INV_X1 U5989 ( .A(n4846), .ZN(n4845) );
  INV_X1 U5990 ( .A(n9739), .ZN(n7116) );
  AND3_X1 U5991 ( .A1(n5198), .A2(n5197), .A3(n5196), .ZN(n9739) );
  AND2_X1 U5992 ( .A1(n4737), .A2(n4734), .ZN(n4411) );
  AND2_X1 U5993 ( .A1(n4505), .A2(n4500), .ZN(n4412) );
  AND2_X1 U5994 ( .A1(n4949), .A2(n6421), .ZN(n4413) );
  OR2_X1 U5995 ( .A1(n6420), .A2(n9828), .ZN(n4414) );
  NAND2_X1 U5996 ( .A1(n6078), .A2(n6077), .ZN(n4415) );
  NAND2_X1 U5997 ( .A1(n4531), .A2(n4405), .ZN(n5872) );
  AND2_X1 U5998 ( .A1(n8647), .A2(n8522), .ZN(n4416) );
  NOR2_X1 U5999 ( .A1(n7888), .A2(n7838), .ZN(n4417) );
  OR2_X1 U6000 ( .A1(n5297), .A2(n4982), .ZN(n4418) );
  NAND2_X1 U6001 ( .A1(n7779), .A2(n7919), .ZN(n4419) );
  AND2_X1 U6002 ( .A1(n5336), .A2(SI_12_), .ZN(n4420) );
  AND2_X1 U6003 ( .A1(n9739), .A2(n5747), .ZN(n4421) );
  NOR2_X1 U6004 ( .A1(n9231), .A2(n9117), .ZN(n4422) );
  OR2_X1 U6005 ( .A1(n9114), .A2(n9415), .ZN(n4423) );
  INV_X1 U6006 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5835) );
  INV_X1 U6007 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5009) );
  INV_X1 U6008 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n6056) );
  INV_X1 U6009 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5885) );
  NOR2_X1 U6010 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .ZN(
        n4424) );
  NOR2_X1 U6011 ( .A1(n8243), .A2(n8746), .ZN(n4425) );
  INV_X1 U6012 ( .A(n4936), .ZN(n4935) );
  NAND2_X1 U6013 ( .A1(n4938), .A2(n5335), .ZN(n4936) );
  AND2_X1 U6014 ( .A1(n7763), .A2(n7838), .ZN(n4426) );
  INV_X1 U6015 ( .A(n4693), .ZN(n4692) );
  NAND2_X1 U6016 ( .A1(n4695), .A2(n8713), .ZN(n4693) );
  AND2_X1 U6017 ( .A1(n4953), .A2(n4980), .ZN(n4427) );
  INV_X1 U6018 ( .A(n4824), .ZN(n4823) );
  NAND2_X1 U6019 ( .A1(n4423), .A2(n4825), .ZN(n4824) );
  NAND2_X1 U6020 ( .A1(n8258), .A2(n8260), .ZN(n4428) );
  NOR2_X1 U6021 ( .A1(n8929), .A2(n8789), .ZN(n4429) );
  INV_X1 U6022 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5482) );
  AND2_X1 U6023 ( .A1(n4778), .A2(n4777), .ZN(n4430) );
  NAND2_X1 U6024 ( .A1(n4398), .A2(n5763), .ZN(n4431) );
  INV_X1 U6025 ( .A(n5534), .ZN(n4741) );
  NAND2_X1 U6026 ( .A1(n9269), .A2(n7796), .ZN(n4432) );
  NAND2_X1 U6027 ( .A1(n4383), .A2(n8396), .ZN(n4433) );
  AND4_X1 U6028 ( .A1(n4765), .A2(n5104), .A3(n4960), .A4(n5053), .ZN(n4978)
         );
  AND3_X1 U6029 ( .A1(n8370), .A2(n8369), .A3(n8368), .ZN(n4434) );
  XNOR2_X1 U6030 ( .A(n8303), .B(n6378), .ZN(n6420) );
  AND2_X1 U6031 ( .A1(n4566), .A2(n4565), .ZN(n4435) );
  INV_X1 U6032 ( .A(n8463), .ZN(n4593) );
  NOR2_X1 U6033 ( .A1(n8993), .A2(n4740), .ZN(n4436) );
  INV_X1 U6034 ( .A(n8457), .ZN(n4878) );
  NAND2_X1 U6035 ( .A1(n8097), .A2(n8096), .ZN(n4437) );
  AND2_X1 U6036 ( .A1(n8432), .A2(n4896), .ZN(n4438) );
  AND2_X1 U6037 ( .A1(n8908), .A2(n8523), .ZN(n8462) );
  INV_X1 U6038 ( .A(n8462), .ZN(n4899) );
  INV_X1 U6039 ( .A(n6111), .ZN(n4706) );
  NAND2_X1 U6040 ( .A1(n5300), .A2(n5299), .ZN(n7446) );
  AND2_X1 U6041 ( .A1(n4392), .A2(n6303), .ZN(n4439) );
  INV_X1 U6042 ( .A(n4922), .ZN(n4921) );
  AND2_X1 U6043 ( .A1(n4751), .A2(n4747), .ZN(n4746) );
  INV_X1 U6044 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5946) );
  NAND2_X1 U6045 ( .A1(n5143), .A2(SI_4_), .ZN(n4440) );
  NAND2_X1 U6046 ( .A1(n7677), .A2(n4397), .ZN(n4773) );
  INV_X1 U6047 ( .A(n7956), .ZN(n4629) );
  NAND2_X1 U6048 ( .A1(n6368), .A2(n7819), .ZN(n8951) );
  AND2_X1 U6049 ( .A1(n9345), .A2(n4572), .ZN(n4441) );
  AND4_X1 U6050 ( .A1(n6187), .A2(n6186), .A3(n6185), .A4(n6184), .ZN(n7993)
         );
  NAND2_X1 U6051 ( .A1(n7677), .A2(n7676), .ZN(n8094) );
  AND2_X1 U6052 ( .A1(n6612), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n4442) );
  OR2_X1 U6053 ( .A1(n6459), .A2(n8874), .ZN(n4443) );
  OAI21_X1 U6054 ( .B1(n9407), .B2(n4827), .A(n4823), .ZN(n9383) );
  XOR2_X1 U6055 ( .A(n5571), .B(n5675), .Z(n4444) );
  NAND2_X1 U6056 ( .A1(n4730), .A2(n4729), .ZN(n9059) );
  NAND2_X1 U6057 ( .A1(n7596), .A2(n7598), .ZN(n7621) );
  AND2_X1 U6058 ( .A1(n4877), .A2(n4383), .ZN(n7592) );
  INV_X1 U6059 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5841) );
  NAND2_X1 U6060 ( .A1(n7558), .A2(n7993), .ZN(n7614) );
  OR2_X1 U6061 ( .A1(n6459), .A2(n8943), .ZN(n4445) );
  AND4_X1 U6062 ( .A1(n6336), .A2(n6335), .A3(n6334), .A4(n6333), .ZN(n8678)
         );
  NOR2_X1 U6063 ( .A1(n8540), .A2(n5987), .ZN(n4446) );
  AND4_X1 U6064 ( .A1(n5270), .A2(n5269), .A3(n5268), .A4(n5267), .ZN(n7431)
         );
  NOR2_X1 U6065 ( .A1(n6469), .A2(n4639), .ZN(n4447) );
  NAND2_X1 U6066 ( .A1(n7536), .A2(n4568), .ZN(n4569) );
  AND4_X1 U6067 ( .A1(n5376), .A2(n5375), .A3(n5374), .A4(n5373), .ZN(n9107)
         );
  AND4_X1 U6068 ( .A1(n5327), .A2(n5326), .A3(n5325), .A4(n5324), .ZN(n7531)
         );
  INV_X1 U6069 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n4810) );
  AND2_X1 U6070 ( .A1(n5463), .A2(n10045), .ZN(n4448) );
  NAND2_X1 U6071 ( .A1(n7781), .A2(n7780), .ZN(n4449) );
  OR2_X1 U6072 ( .A1(n4932), .A2(n4931), .ZN(n4450) );
  AND2_X1 U6073 ( .A1(n5874), .A2(n4770), .ZN(n4451) );
  AND2_X1 U6074 ( .A1(n4660), .A2(n5932), .ZN(n4452) );
  INV_X1 U6075 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n4961) );
  OR2_X1 U6076 ( .A1(n9749), .A2(n4479), .ZN(n4453) );
  INV_X1 U6077 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n4809) );
  INV_X1 U6078 ( .A(n7598), .ZN(n4733) );
  XNOR2_X1 U6079 ( .A(n5845), .B(n5844), .ZN(n6424) );
  AND2_X2 U6080 ( .A1(n6456), .A2(n6849), .ZN(n9887) );
  OR2_X1 U6081 ( .A1(n9814), .A2(n9813), .ZN(n4454) );
  NAND2_X1 U6082 ( .A1(n7173), .A2(n7178), .ZN(n7174) );
  NAND2_X1 U6083 ( .A1(n6895), .A2(n6896), .ZN(n7238) );
  AND2_X1 U6084 ( .A1(n6819), .A2(n6818), .ZN(n6824) );
  OR2_X1 U6085 ( .A1(n7653), .A2(n5935), .ZN(n4455) );
  NAND2_X1 U6086 ( .A1(n7238), .A2(n4807), .ZN(n8246) );
  INV_X1 U6087 ( .A(n4892), .ZN(n4891) );
  NOR2_X1 U6088 ( .A1(n6390), .A2(n4893), .ZN(n4892) );
  NAND2_X1 U6089 ( .A1(n4371), .A2(n7210), .ZN(n4564) );
  NOR2_X1 U6090 ( .A1(n6007), .A2(n4538), .ZN(n4456) );
  OR2_X1 U6091 ( .A1(n8624), .A2(n8627), .ZN(n4457) );
  OAI211_X1 U6092 ( .C1(n5038), .C2(n6545), .A(n5092), .B(n5091), .ZN(n7098)
         );
  NAND2_X1 U6093 ( .A1(n7875), .A2(n7841), .ZN(n7919) );
  INV_X1 U6094 ( .A(n8599), .ZN(n7019) );
  INV_X1 U6095 ( .A(n7094), .ZN(n4578) );
  INV_X2 U6096 ( .A(n5111), .ZN(n7830) );
  NAND2_X1 U6097 ( .A1(n5038), .A2(n6491), .ZN(n5111) );
  OR2_X1 U6098 ( .A1(n9887), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n4458) );
  NOR2_X1 U6099 ( .A1(n9784), .A2(n5919), .ZN(n4459) );
  NOR2_X1 U6100 ( .A1(n4962), .A2(n4513), .ZN(n9581) );
  INV_X1 U6101 ( .A(n7928), .ZN(n7875) );
  NOR2_X1 U6102 ( .A1(n5910), .A2(n9773), .ZN(n5911) );
  INV_X1 U6103 ( .A(n5911), .ZN(n4664) );
  AND2_X1 U6104 ( .A1(n4908), .A2(n7982), .ZN(n4460) );
  NAND2_X1 U6105 ( .A1(n5842), .A2(n5841), .ZN(n5865) );
  NAND2_X2 U6106 ( .A1(n6785), .A2(n6784), .ZN(n6804) );
  INV_X1 U6107 ( .A(n6807), .ZN(n4768) );
  NAND2_X2 U6108 ( .A1(n4462), .A2(n4391), .ZN(n4712) );
  OR2_X2 U6109 ( .A1(n8575), .A2(n8864), .ZN(n4462) );
  NOR2_X2 U6110 ( .A1(n7645), .A2(n4463), .ZN(n5986) );
  NOR2_X2 U6111 ( .A1(n7647), .A2(n7646), .ZN(n7645) );
  NAND2_X1 U6112 ( .A1(n7579), .A2(n8394), .ZN(n7578) );
  OAI21_X1 U6113 ( .B1(n6350), .B2(n4406), .A(n6349), .ZN(n4469) );
  OAI21_X1 U6114 ( .B1(n8709), .B2(n4689), .A(n4688), .ZN(n6318) );
  AOI22_X2 U6115 ( .A1(n7450), .A2(n8379), .B1(n8530), .B2(n9870), .ZN(n7542)
         );
  NAND2_X1 U6116 ( .A1(n9859), .A2(n7396), .ZN(n8364) );
  NAND2_X4 U6117 ( .A1(n6076), .A2(n6491), .ZN(n8291) );
  NAND2_X1 U6118 ( .A1(n4470), .A2(n6176), .ZN(n4677) );
  NAND2_X2 U6119 ( .A1(n6002), .A2(n5960), .ZN(n6076) );
  OAI22_X1 U6120 ( .A1(n8719), .A2(n8725), .B1(n8525), .B2(n8727), .ZN(n8709)
         );
  NAND2_X1 U6121 ( .A1(n8663), .A2(n8662), .ZN(n8661) );
  AOI21_X2 U6122 ( .B1(n4471), .B2(n8759), .A(n8640), .ZN(n8809) );
  NAND2_X1 U6123 ( .A1(n4476), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n6477) );
  NOR2_X1 U6124 ( .A1(n8544), .A2(n8543), .ZN(n8542) );
  NOR2_X1 U6125 ( .A1(n8561), .A2(n8560), .ZN(n8559) );
  NAND3_X1 U6126 ( .A1(n4474), .A2(n6051), .A3(n4472), .ZN(P2_U3201) );
  NAND2_X1 U6127 ( .A1(n5944), .A2(n4656), .ZN(n4652) );
  XNOR2_X1 U6128 ( .A(n4473), .B(n5995), .ZN(n5993) );
  NAND2_X1 U6129 ( .A1(n5968), .A2(n9773), .ZN(n5969) );
  OAI21_X2 U6130 ( .B1(n6401), .B2(n4866), .A(n4863), .ZN(n8644) );
  NAND2_X1 U6131 ( .A1(n9238), .A2(n7897), .ZN(n9226) );
  AND2_X2 U6132 ( .A1(n5805), .A2(n7785), .ZN(n9321) );
  NAND2_X2 U6133 ( .A1(n7321), .A2(n5792), .ZN(n7430) );
  OR2_X2 U6134 ( .A1(n9386), .A2(n9385), .ZN(n9388) );
  NAND2_X2 U6135 ( .A1(n9285), .A2(n9288), .ZN(n9284) );
  INV_X1 U6136 ( .A(n6379), .ZN(n5842) );
  NAND2_X1 U6137 ( .A1(n6803), .A2(n6802), .ZN(n8228) );
  OR2_X1 U6138 ( .A1(n5897), .A2(n6081), .ZN(n5963) );
  XNOR2_X2 U6139 ( .A(n5989), .B(n6239), .ZN(n9801) );
  NOR2_X1 U6140 ( .A1(n7342), .A2(n7341), .ZN(n7340) );
  NOR2_X1 U6141 ( .A1(n6947), .A2(n6133), .ZN(n6946) );
  INV_X1 U6142 ( .A(n5986), .ZN(n4728) );
  NAND2_X1 U6143 ( .A1(n5993), .A2(n5992), .ZN(n4474) );
  NOR2_X1 U6144 ( .A1(n6953), .A2(n9826), .ZN(n6952) );
  XNOR2_X1 U6145 ( .A(n5925), .B(n6139), .ZN(n6953) );
  INV_X1 U6146 ( .A(n8617), .ZN(n8613) );
  AND3_X2 U6147 ( .A1(n4657), .A2(n4659), .A3(n4455), .ZN(n5936) );
  NOR2_X1 U6148 ( .A1(n7051), .A2(n7050), .ZN(n7049) );
  OAI211_X1 U6149 ( .C1(n8625), .C2(n4457), .A(n4554), .B(n4553), .ZN(n4552)
         );
  NAND2_X1 U6150 ( .A1(n6477), .A2(n5899), .ZN(n6651) );
  INV_X1 U6151 ( .A(n6479), .ZN(n4476) );
  NAND2_X1 U6152 ( .A1(n4645), .A2(n4644), .ZN(n4643) );
  NAND2_X1 U6153 ( .A1(n5167), .A2(n5166), .ZN(n4579) );
  INV_X1 U6154 ( .A(n4818), .ZN(n4817) );
  INV_X1 U6155 ( .A(n9311), .ZN(n4854) );
  NAND2_X1 U6156 ( .A1(n4816), .A2(n4815), .ZN(n7209) );
  NOR2_X2 U6157 ( .A1(n8557), .A2(n4951), .ZN(n5988) );
  AND3_X2 U6158 ( .A1(n4725), .A2(n4724), .A3(n4727), .ZN(n8557) );
  NAND2_X1 U6159 ( .A1(n5962), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6474) );
  AND2_X2 U6160 ( .A1(n4721), .A2(n4720), .ZN(n5981) );
  NAND3_X1 U6161 ( .A1(n4484), .A2(n4907), .A3(n7985), .ZN(P1_U3242) );
  NAND2_X1 U6162 ( .A1(n4485), .A2(n4904), .ZN(n4484) );
  NAND2_X1 U6163 ( .A1(n4486), .A2(n7875), .ZN(n4485) );
  NAND2_X1 U6164 ( .A1(n7874), .A2(n7914), .ZN(n4486) );
  NAND2_X1 U6165 ( .A1(n4494), .A2(n4492), .ZN(n4490) );
  INV_X1 U6166 ( .A(n7921), .ZN(n7842) );
  NAND2_X1 U6167 ( .A1(n7839), .A2(n4501), .ZN(n4495) );
  INV_X1 U6168 ( .A(n7920), .ZN(n4504) );
  OR2_X2 U6169 ( .A1(n6669), .A2(n5787), .ZN(n7933) );
  INV_X1 U6170 ( .A(n4962), .ZN(n4512) );
  NOR2_X1 U6171 ( .A1(n4962), .A2(n4857), .ZN(n4990) );
  INV_X1 U6172 ( .A(n6008), .ZN(n4539) );
  NOR2_X1 U6173 ( .A1(n8548), .A2(n8547), .ZN(n8546) );
  INV_X1 U6174 ( .A(n6005), .ZN(n4551) );
  NAND3_X1 U6175 ( .A1(n4978), .A2(n4561), .A3(n4560), .ZN(n4562) );
  INV_X1 U6176 ( .A(n4564), .ZN(n7436) );
  NAND2_X1 U6177 ( .A1(n7536), .A2(n4435), .ZN(n9358) );
  INV_X1 U6178 ( .A(n4569), .ZN(n9396) );
  NAND3_X1 U6179 ( .A1(n4576), .A2(n6971), .A3(n4575), .ZN(n4577) );
  NAND3_X1 U6180 ( .A1(n4578), .A2(n4364), .A3(n5744), .ZN(n7181) );
  NAND3_X1 U6181 ( .A1(n4581), .A2(n4580), .A3(n4440), .ZN(n5167) );
  NAND3_X1 U6182 ( .A1(n5141), .A2(n5113), .A3(n5112), .ZN(n4581) );
  OAI21_X1 U6183 ( .B1(n8406), .B2(n4587), .A(n4582), .ZN(n8417) );
  NAND2_X1 U6184 ( .A1(n8414), .A2(n8408), .ZN(n4594) );
  NAND3_X1 U6185 ( .A1(n8359), .A2(n4434), .A3(n8360), .ZN(n8377) );
  NAND3_X1 U6186 ( .A1(n4599), .A2(n4602), .A3(n4598), .ZN(n8520) );
  NAND3_X1 U6187 ( .A1(n4600), .A2(n8457), .A3(n4601), .ZN(n4599) );
  INV_X1 U6188 ( .A(n8513), .ZN(n4600) );
  NAND3_X1 U6189 ( .A1(n4605), .A2(n4604), .A3(n4608), .ZN(n8405) );
  NAND2_X1 U6190 ( .A1(n8393), .A2(n4607), .ZN(n4604) );
  NAND2_X1 U6191 ( .A1(n8390), .A2(n4606), .ZN(n4605) );
  NAND3_X1 U6192 ( .A1(n4617), .A2(n4614), .A3(n8708), .ZN(n4613) );
  INV_X1 U6193 ( .A(n4620), .ZN(n7061) );
  NAND2_X1 U6194 ( .A1(n4627), .A2(n4630), .ZN(n9386) );
  NAND2_X1 U6195 ( .A1(n5797), .A2(n4628), .ZN(n4627) );
  NAND2_X1 U6196 ( .A1(n9239), .A2(n4636), .ZN(n4633) );
  NAND2_X1 U6197 ( .A1(n4633), .A2(n4634), .ZN(n8061) );
  NAND2_X1 U6198 ( .A1(n9239), .A2(n9242), .ZN(n9238) );
  OR2_X2 U6199 ( .A1(n9328), .A2(n9329), .ZN(n5805) );
  OAI21_X2 U6200 ( .B1(n9340), .B2(n9341), .A(n7970), .ZN(n9328) );
  NAND2_X2 U6201 ( .A1(n5803), .A2(n7967), .ZN(n9340) );
  OAI21_X1 U6202 ( .B1(n4650), .B2(n4649), .A(n7711), .ZN(n4648) );
  AND2_X1 U6203 ( .A1(n7849), .A2(n7936), .ZN(n4650) );
  XNOR2_X1 U6204 ( .A(n5943), .B(n8583), .ZN(n8577) );
  INV_X1 U6205 ( .A(n4660), .ZN(n7472) );
  NAND2_X1 U6206 ( .A1(n5919), .A2(n4663), .ZN(n4661) );
  NOR2_X1 U6207 ( .A1(n4665), .A2(n5911), .ZN(n6697) );
  NOR2_X2 U6208 ( .A1(n7351), .A2(n7352), .ZN(n7350) );
  NAND3_X1 U6209 ( .A1(n4678), .A2(n4677), .A3(n4675), .ZN(n4674) );
  NAND2_X1 U6210 ( .A1(n4406), .A2(n6349), .ZN(n4684) );
  CLKBUF_X1 U6211 ( .A(n8709), .Z(n4686) );
  NAND2_X1 U6212 ( .A1(n8787), .A2(n4698), .ZN(n4697) );
  OAI21_X1 U6213 ( .B1(n8787), .B2(n4699), .A(n4698), .ZN(n8761) );
  NAND3_X1 U6215 ( .A1(n6101), .A2(n8321), .A3(n6111), .ZN(n4705) );
  NAND2_X1 U6216 ( .A1(n6101), .A2(n8321), .ZN(n6878) );
  OR2_X1 U6217 ( .A1(n5897), .A2(n6080), .ZN(n5899) );
  AND2_X1 U6218 ( .A1(n5897), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5900) );
  NAND2_X1 U6219 ( .A1(n6419), .A2(n4368), .ZN(n6457) );
  NAND2_X1 U6220 ( .A1(n6419), .A2(n4369), .ZN(n6458) );
  NAND2_X1 U6221 ( .A1(n6419), .A2(n6418), .ZN(n7697) );
  NAND2_X1 U6222 ( .A1(n6474), .A2(n5963), .ZN(n6649) );
  INV_X1 U6223 ( .A(n5990), .ZN(n4717) );
  NOR2_X1 U6224 ( .A1(n9801), .A2(n9802), .ZN(n9800) );
  INV_X1 U6225 ( .A(n4719), .ZN(n8610) );
  OR2_X2 U6226 ( .A1(n6946), .A2(n5979), .ZN(n4723) );
  OR2_X1 U6227 ( .A1(n5987), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n4724) );
  NAND2_X1 U6228 ( .A1(n4726), .A2(n8541), .ZN(n4725) );
  XNOR2_X2 U6229 ( .A(n4728), .B(n6716), .ZN(n8541) );
  INV_X1 U6230 ( .A(n5987), .ZN(n4726) );
  NOR2_X1 U6231 ( .A1(n8541), .A2(n8872), .ZN(n8540) );
  NOR2_X1 U6232 ( .A1(n9883), .A2(n7476), .ZN(n7475) );
  NOR2_X1 U6233 ( .A1(n5929), .A2(n7350), .ZN(n7408) );
  NAND2_X1 U6234 ( .A1(n6651), .A2(n6652), .ZN(n6650) );
  NAND2_X1 U6235 ( .A1(n5896), .A2(n5897), .ZN(n6003) );
  XNOR2_X1 U6236 ( .A(n5988), .B(n8583), .ZN(n8575) );
  OAI21_X1 U6237 ( .B1(n5966), .B2(n5965), .A(n5964), .ZN(n6647) );
  NAND2_X1 U6238 ( .A1(n5970), .A2(n5969), .ZN(n9765) );
  NAND2_X1 U6239 ( .A1(n7597), .A2(n4731), .ZN(n4730) );
  NAND2_X1 U6240 ( .A1(n9053), .A2(n4436), .ZN(n4735) );
  NAND2_X1 U6241 ( .A1(n4735), .A2(n4737), .ZN(n5554) );
  NAND3_X1 U6242 ( .A1(n4743), .A2(n5286), .A3(n5285), .ZN(n9625) );
  NAND2_X1 U6243 ( .A1(n5282), .A2(n5281), .ZN(n5286) );
  AOI21_X1 U6244 ( .B1(n8971), .B2(n4746), .A(n4744), .ZN(n5680) );
  NAND2_X1 U6245 ( .A1(n4748), .A2(n4751), .ZN(n9001) );
  NAND2_X1 U6246 ( .A1(n5357), .A2(n4757), .ZN(n4754) );
  NAND2_X1 U6247 ( .A1(n4754), .A2(n4755), .ZN(n5459) );
  NAND2_X1 U6248 ( .A1(n5393), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4761) );
  NAND2_X1 U6249 ( .A1(n4761), .A2(n4762), .ZN(n5485) );
  NAND3_X1 U6250 ( .A1(n5236), .A2(n4764), .A3(n5235), .ZN(n7283) );
  NAND2_X1 U6251 ( .A1(n5232), .A2(n5231), .ZN(n4764) );
  OR2_X2 U6252 ( .A1(n5232), .A2(n5231), .ZN(n5236) );
  NAND3_X1 U6253 ( .A1(n4960), .A2(n5053), .A3(n5104), .ZN(n5164) );
  NAND3_X1 U6254 ( .A1(n6790), .A2(n6802), .A3(n6792), .ZN(n6803) );
  NAND3_X1 U6255 ( .A1(n6819), .A2(n6818), .A3(n6826), .ZN(n6894) );
  INV_X1 U6256 ( .A(n6809), .ZN(n4767) );
  NAND2_X1 U6257 ( .A1(n5874), .A2(n4769), .ZN(n5950) );
  INV_X1 U6258 ( .A(n5950), .ZN(n5952) );
  NAND2_X1 U6259 ( .A1(n7368), .A2(n4776), .ZN(n7504) );
  INV_X1 U6260 ( .A(n7557), .ZN(n7558) );
  NAND4_X1 U6261 ( .A1(n5833), .A2(n5832), .A3(n5891), .A4(n5831), .ZN(n5834)
         );
  NAND2_X1 U6262 ( .A1(n8214), .A2(n4784), .ZN(n4783) );
  NAND2_X2 U6263 ( .A1(n4783), .A2(n4779), .ZN(n8113) );
  NAND2_X1 U6264 ( .A1(n8121), .A2(n4792), .ZN(n4791) );
  NAND2_X1 U6265 ( .A1(n4791), .A2(n4795), .ZN(n8131) );
  NAND2_X1 U6266 ( .A1(n8179), .A2(n8180), .ZN(n8257) );
  OR3_X1 U6267 ( .A1(n5957), .A2(n5837), .A3(n6058), .ZN(n4801) );
  NAND2_X1 U6268 ( .A1(n5957), .A2(n4804), .ZN(n4800) );
  NAND3_X1 U6269 ( .A1(n4808), .A2(n4814), .A3(n4813), .ZN(n4981) );
  AND2_X1 U6270 ( .A1(n4958), .A2(n4959), .ZN(n4814) );
  NAND2_X1 U6271 ( .A1(n7173), .A2(n4817), .ZN(n4816) );
  INV_X1 U6272 ( .A(n9407), .ZN(n4821) );
  AND2_X1 U6273 ( .A1(n9399), .A2(n9127), .ZN(n4830) );
  NAND2_X1 U6274 ( .A1(n5767), .A2(n4833), .ZN(n4837) );
  NAND2_X1 U6275 ( .A1(n5767), .A2(n4843), .ZN(n4835) );
  NAND2_X1 U6276 ( .A1(n5767), .A2(n5766), .ZN(n9252) );
  NOR2_X1 U6277 ( .A1(n5769), .A2(n4844), .ZN(n4843) );
  INV_X1 U6278 ( .A(n5766), .ZN(n4844) );
  NOR2_X1 U6279 ( .A1(n9540), .A2(n7798), .ZN(n4846) );
  INV_X1 U6280 ( .A(n5901), .ZN(n5830) );
  INV_X1 U6281 ( .A(n8467), .ZN(n8321) );
  AND2_X2 U6282 ( .A1(n8326), .A2(n8325), .ZN(n8467) );
  NAND3_X1 U6283 ( .A1(n6383), .A2(n8320), .A3(n8316), .ZN(n6836) );
  NAND2_X1 U6284 ( .A1(n5884), .A2(n4862), .ZN(n6379) );
  NAND2_X1 U6285 ( .A1(n4872), .A2(n4874), .ZN(n6396) );
  NAND2_X1 U6286 ( .A1(n7449), .A2(n4876), .ZN(n4872) );
  AOI21_X1 U6287 ( .B1(n7122), .B2(n4887), .A(n4886), .ZN(n7989) );
  OAI21_X1 U6288 ( .B1(n8712), .B2(n4897), .A(n4438), .ZN(n6400) );
  INV_X2 U6289 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n7999) );
  NAND2_X1 U6290 ( .A1(n4909), .A2(n7926), .ZN(n4906) );
  NAND3_X1 U6291 ( .A1(n4906), .A2(n4905), .A3(n4908), .ZN(n4907) );
  NAND2_X1 U6292 ( .A1(n5601), .A2(n5600), .ZN(n5619) );
  NAND2_X1 U6293 ( .A1(n5601), .A2(n4911), .ZN(n4910) );
  OR2_X2 U6294 ( .A1(n5441), .A2(n4922), .ZN(n4918) );
  OAI21_X1 U6295 ( .B1(n5441), .B2(n5440), .A(n4384), .ZN(n5461) );
  NAND2_X1 U6296 ( .A1(n4923), .A2(n5460), .ZN(n4922) );
  NAND2_X1 U6297 ( .A1(n4924), .A2(n5115), .ZN(n5142) );
  NAND2_X1 U6298 ( .A1(n5113), .A2(n5112), .ZN(n4924) );
  INV_X2 U6299 ( .A(n7825), .ZN(n4999) );
  NAND3_X1 U6300 ( .A1(n4927), .A2(n4926), .A3(P2_DATAO_REG_1__SCAN_IN), .ZN(
        n5001) );
  NAND2_X1 U6301 ( .A1(n5517), .A2(n4929), .ZN(n4928) );
  NAND2_X1 U6302 ( .A1(n4928), .A2(n4930), .ZN(n5557) );
  NAND2_X1 U6303 ( .A1(n5517), .A2(n5516), .ZN(n5537) );
  INV_X1 U6304 ( .A(n5516), .ZN(n4931) );
  INV_X1 U6305 ( .A(n5535), .ZN(n4932) );
  OAI21_X2 U6306 ( .B1(n5289), .B2(n4936), .A(n4933), .ZN(n5362) );
  NOR2_X2 U6307 ( .A1(n5314), .A2(n4941), .ZN(n4940) );
  AND2_X1 U6308 ( .A1(n5781), .A2(n5021), .ZN(n4987) );
  NOR2_X1 U6309 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n4960) );
  AOI21_X2 U6310 ( .B1(n8652), .B2(n8759), .A(n8651), .ZN(n8813) );
  NAND2_X1 U6311 ( .A1(n8036), .A2(n7072), .ZN(n5023) );
  CLKBUF_X1 U6312 ( .A(n7173), .Z(n7175) );
  NAND4_X2 U6313 ( .A1(n5020), .A2(n5019), .A3(n5018), .A4(n5017), .ZN(n5737)
         );
  MUX2_X1 U6314 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8962), .S(n6076), .Z(n7003) );
  AND2_X2 U6315 ( .A1(n5016), .A2(n5015), .ZN(n5099) );
  INV_X1 U6316 ( .A(n5015), .ZN(n9590) );
  OR2_X1 U6317 ( .A1(n6059), .A2(n6058), .ZN(n6061) );
  OR2_X1 U6318 ( .A1(n8539), .A2(n6993), .ZN(n8338) );
  INV_X1 U6319 ( .A(n8055), .ZN(n8085) );
  NAND2_X1 U6320 ( .A1(n7928), .A2(n7927), .ZN(n5711) );
  NAND2_X1 U6321 ( .A1(n7928), .A2(n5712), .ZN(n5781) );
  INV_X1 U6322 ( .A(n9231), .ZN(n9536) );
  XNOR2_X1 U6323 ( .A(n6362), .B(n6361), .ZN(n6351) );
  OR2_X1 U6324 ( .A1(n6411), .A2(n5906), .ZN(n6093) );
  OR2_X1 U6325 ( .A1(n6411), .A2(n6480), .ZN(n6073) );
  OAI21_X1 U6326 ( .B1(n4999), .B2(n5061), .A(n5060), .ZN(n5088) );
  NAND2_X1 U6327 ( .A1(n4999), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5060) );
  NAND2_X1 U6328 ( .A1(n7825), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5000) );
  NAND2_X2 U6329 ( .A1(n6853), .A2(n8679), .ZN(n9824) );
  AND2_X1 U6330 ( .A1(n6201), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n4942) );
  AND2_X1 U6331 ( .A1(n8103), .A2(n8789), .ZN(n4943) );
  AND2_X1 U6332 ( .A1(n6314), .A2(n6313), .ZN(n8700) );
  INV_X1 U6333 ( .A(n8700), .ZN(n6315) );
  AND3_X1 U6334 ( .A1(n6273), .A2(n6272), .A3(n6271), .ZN(n8722) );
  INV_X1 U6335 ( .A(n8722), .ZN(n6274) );
  NOR2_X1 U6336 ( .A1(n9031), .A2(n5397), .ZN(n4944) );
  OR2_X1 U6337 ( .A1(n9561), .A2(n9343), .ZN(n4945) );
  OR2_X1 U6338 ( .A1(n7072), .A2(n5737), .ZN(n4947) );
  INV_X1 U6339 ( .A(n7653), .ZN(n6688) );
  NAND2_X1 U6340 ( .A1(n9760), .A2(n6004), .ZN(n9803) );
  INV_X1 U6341 ( .A(n9803), .ZN(n5992) );
  AND2_X1 U6342 ( .A1(n7672), .A2(n8530), .ZN(n4948) );
  OR2_X1 U6343 ( .A1(n8805), .A2(n8633), .ZN(n4949) );
  AND2_X1 U6344 ( .A1(n6777), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n4950) );
  INV_X1 U6345 ( .A(n7927), .ZN(n7982) );
  AND2_X1 U6346 ( .A1(n6777), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n4951) );
  INV_X1 U6347 ( .A(n8549), .ZN(n6716) );
  NOR2_X1 U6348 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n4952) );
  INV_X1 U6349 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n5061) );
  INV_X1 U6350 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n5117) );
  INV_X1 U6351 ( .A(n8956), .ZN(n6628) );
  INV_X1 U6352 ( .A(n8107), .ZN(n8920) );
  INV_X1 U6353 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n5972) );
  INV_X1 U6354 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n5906) );
  INV_X1 U6355 ( .A(SI_20_), .ZN(n5536) );
  INV_X1 U6356 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n5084) );
  INV_X1 U6357 ( .A(n9135), .ZN(n5747) );
  OR2_X1 U6358 ( .A1(n7804), .A2(n7803), .ZN(n4954) );
  OR2_X1 U6359 ( .A1(n6804), .A2(n7003), .ZN(n4955) );
  INV_X1 U6360 ( .A(n9629), .ZN(n5750) );
  AND2_X1 U6361 ( .A1(n8106), .A2(n8764), .ZN(n4956) );
  INV_X1 U6362 ( .A(n6001), .ZN(n6694) );
  INV_X1 U6363 ( .A(n6694), .ZN(n5914) );
  INV_X1 U6364 ( .A(n7975), .ZN(n7922) );
  OR2_X1 U6365 ( .A1(n9318), .A2(n5806), .ZN(n4957) );
  INV_X1 U6366 ( .A(n7727), .ZN(n5744) );
  INV_X1 U6367 ( .A(n7728), .ZN(n9137) );
  INV_X1 U6368 ( .A(n7090), .ZN(n9138) );
  INV_X1 U6369 ( .A(n9433), .ZN(n9381) );
  INV_X1 U6370 ( .A(n5217), .ZN(n5066) );
  INV_X1 U6371 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n5965) );
  AND2_X1 U6372 ( .A1(n6783), .A2(n8501), .ZN(n6784) );
  NAND2_X1 U6373 ( .A1(n5966), .A2(n5906), .ZN(n5905) );
  INV_X1 U6374 ( .A(n8036), .ZN(n5093) );
  NAND2_X1 U6375 ( .A1(n5711), .A2(n5021), .ZN(n4988) );
  INV_X1 U6376 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n10000) );
  INV_X1 U6377 ( .A(SI_28_), .ZN(n10062) );
  OR2_X1 U6378 ( .A1(n8115), .A2(n8114), .ZN(n8116) );
  INV_X1 U6379 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n10091) );
  OR2_X1 U6380 ( .A1(n6287), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6296) );
  INV_X1 U6381 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n6208) );
  NAND2_X1 U6382 ( .A1(n6076), .A2(n7825), .ZN(n6097) );
  AND4_X1 U6383 ( .A1(n5854), .A2(n5862), .A3(n5851), .A4(n5850), .ZN(n5852)
         );
  INV_X1 U6384 ( .A(n5933), .ZN(n5874) );
  INV_X1 U6385 ( .A(n5429), .ZN(n5430) );
  OR2_X1 U6386 ( .A1(n9066), .A2(n9129), .ZN(n5755) );
  INV_X1 U6387 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n5209) );
  INV_X1 U6388 ( .A(SI_26_), .ZN(n10071) );
  INV_X1 U6389 ( .A(SI_19_), .ZN(n10095) );
  INV_X1 U6390 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n4972) );
  INV_X1 U6391 ( .A(SI_11_), .ZN(n10014) );
  INV_X1 U6392 ( .A(n7615), .ZN(n7562) );
  NAND2_X1 U6393 ( .A1(n6242), .A2(n10091), .ZN(n6250) );
  AND2_X1 U6394 ( .A1(n6764), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5977) );
  NAND2_X1 U6395 ( .A1(n8184), .A2(n8689), .ZN(n8427) );
  INV_X1 U6396 ( .A(n8713), .ZN(n8708) );
  NAND2_X1 U6397 ( .A1(n8202), .A2(n8789), .ZN(n8407) );
  NOR2_X1 U6398 ( .A1(n9828), .A2(n8310), .ZN(n6733) );
  OR2_X2 U6399 ( .A1(n7369), .A2(n7258), .ZN(n8356) );
  NAND2_X1 U6400 ( .A1(n8345), .A2(n8347), .ZN(n8473) );
  INV_X1 U6401 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5844) );
  NAND2_X1 U6402 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n5895) );
  INV_X1 U6403 ( .A(n7286), .ZN(n5235) );
  INV_X1 U6404 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5131) );
  INV_X1 U6405 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5237) );
  INV_X1 U6406 ( .A(n6639), .ZN(n5047) );
  INV_X1 U6407 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n5415) );
  OR2_X1 U6408 ( .A1(n5210), .A2(n5209), .ZN(n5238) );
  NAND2_X1 U6409 ( .A1(n5750), .A2(n7431), .ZN(n5751) );
  NAND2_X1 U6410 ( .A1(n7309), .A2(n7385), .ZN(n5748) );
  AND2_X1 U6411 ( .A1(n6363), .A2(n5776), .ZN(n6361) );
  INV_X1 U6412 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n4980) );
  INV_X1 U6413 ( .A(SI_17_), .ZN(n10045) );
  INV_X1 U6414 ( .A(SI_14_), .ZN(n5386) );
  NAND2_X1 U6415 ( .A1(n6053), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n5116) );
  AND2_X1 U6416 ( .A1(n6230), .A2(n6229), .ZN(n6242) );
  INV_X1 U6417 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n10048) );
  OR2_X1 U6418 ( .A1(n6211), .A2(n8667), .ZN(n6334) );
  NAND2_X1 U6419 ( .A1(n8615), .A2(n8614), .ZN(n8616) );
  AND2_X1 U6420 ( .A1(n7698), .A2(n6356), .ZN(n8641) );
  NAND2_X1 U6421 ( .A1(n6733), .A2(n6746), .ZN(n8679) );
  OR2_X1 U6422 ( .A1(n6846), .A2(n6444), .ZN(n6455) );
  INV_X1 U6423 ( .A(n8759), .ZN(n8786) );
  AND2_X1 U6424 ( .A1(n6936), .A2(n9828), .ZN(n9866) );
  INV_X1 U6425 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n8987) );
  OR2_X1 U6426 ( .A1(n9088), .A2(n9089), .ZN(n5655) );
  INV_X1 U6427 ( .A(n9392), .ZN(n9415) );
  AND2_X1 U6428 ( .A1(n5418), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9031) );
  INV_X1 U6429 ( .A(n5627), .ZN(n5626) );
  NOR2_X1 U6430 ( .A1(n5521), .A2(n9054), .ZN(n5540) );
  INV_X1 U6431 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n7602) );
  NOR2_X1 U6432 ( .A1(n5416), .A2(n5415), .ZN(n5418) );
  INV_X1 U6433 ( .A(n5718), .ZN(n5729) );
  NAND2_X1 U6434 ( .A1(n5566), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n5583) );
  OR2_X1 U6435 ( .A1(n6554), .A2(n9157), .ZN(n9718) );
  INV_X1 U6436 ( .A(n7868), .ZN(n9269) );
  INV_X1 U6437 ( .A(n7536), .ZN(n9424) );
  AND2_X1 U6438 ( .A1(n9741), .A2(n9406), .ZN(n7067) );
  OR2_X1 U6439 ( .A1(n6506), .A2(n5824), .ZN(n6465) );
  AND2_X1 U6440 ( .A1(n5711), .A2(n5822), .ZN(n9724) );
  INV_X1 U6441 ( .A(n9477), .ZN(n9422) );
  NAND2_X1 U6442 ( .A1(n5704), .A2(n9580), .ZN(n6464) );
  AND2_X1 U6443 ( .A1(n5688), .A2(n5687), .ZN(n5689) );
  AND2_X1 U6444 ( .A1(n5620), .A2(n5604), .ZN(n5618) );
  AND2_X1 U6445 ( .A1(n6749), .A2(n6748), .ZN(n8267) );
  AND2_X1 U6446 ( .A1(n6796), .A2(n6795), .ZN(n8277) );
  NAND2_X1 U6447 ( .A1(n6734), .A2(n8679), .ZN(n8269) );
  OR2_X1 U6448 ( .A1(n6211), .A2(n7698), .ZN(n8299) );
  AND2_X1 U6449 ( .A1(n6284), .A2(n6283), .ZN(n8735) );
  AND4_X1 U6450 ( .A1(n6205), .A2(n6204), .A3(n6203), .A4(n6202), .ZN(n7992)
         );
  INV_X1 U6451 ( .A(n8628), .ZN(n9796) );
  INV_X1 U6452 ( .A(n8673), .ZN(n8801) );
  OR2_X1 U6453 ( .A1(P2_REG0_REG_29__SCAN_IN), .A2(n8939), .ZN(n6448) );
  NAND2_X2 U6454 ( .A1(n6167), .A2(n6166), .ZN(n7369) );
  INV_X1 U6455 ( .A(n9866), .ZN(n9853) );
  AND2_X1 U6456 ( .A1(n6738), .A2(n6619), .ZN(n6746) );
  AND2_X1 U6457 ( .A1(n5941), .A2(n5940), .ZN(n8566) );
  BUF_X4 U6458 ( .A(n6053), .Z(n6491) );
  OAI21_X1 U6459 ( .B1(n9536), .B2(n9113), .A(n5732), .ZN(n5733) );
  AND4_X1 U6460 ( .A1(n5725), .A2(n5724), .A3(n5723), .A4(n5722), .ZN(n8054)
         );
  AND4_X1 U6461 ( .A1(n5496), .A2(n5495), .A3(n5494), .A4(n5493), .ZN(n9375)
         );
  AND4_X1 U6462 ( .A1(n5401), .A2(n5400), .A3(n5399), .A4(n5398), .ZN(n9373)
         );
  INV_X1 U6463 ( .A(n9712), .ZN(n9669) );
  INV_X1 U6464 ( .A(n9718), .ZN(n9699) );
  INV_X1 U6465 ( .A(n9371), .ZN(n9368) );
  INV_X1 U6466 ( .A(n9360), .ZN(n9431) );
  AND2_X1 U6467 ( .A1(n9157), .A2(n6508), .ZN(n9393) );
  INV_X1 U6468 ( .A(n9496), .ZN(n9746) );
  AND3_X1 U6469 ( .A1(n5827), .A2(n5826), .A3(n5825), .ZN(n6467) );
  INV_X1 U6470 ( .A(n6506), .ZN(n9578) );
  INV_X1 U6471 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n4965) );
  XNOR2_X1 U6472 ( .A(n5340), .B(P1_IR_REG_13__SCAN_IN), .ZN(n9653) );
  OR2_X1 U6473 ( .A1(n6725), .A2(n6795), .ZN(n8279) );
  AND2_X1 U6474 ( .A1(n6731), .A2(n6730), .ZN(n8271) );
  AND4_X1 U6475 ( .A1(n8299), .A2(n6377), .A3(n6376), .A4(n6375), .ZN(n8638)
         );
  INV_X1 U6476 ( .A(n8735), .ZN(n8525) );
  INV_X1 U6477 ( .A(n8096), .ZN(n8528) );
  INV_X1 U6478 ( .A(n9772), .ZN(n9814) );
  NAND2_X1 U6479 ( .A1(n9760), .A2(n8514), .ZN(n9810) );
  NAND2_X1 U6480 ( .A1(n9824), .A2(n9815), .ZN(n8673) );
  INV_X1 U6481 ( .A(n8875), .ZN(n8805) );
  NAND2_X1 U6482 ( .A1(n9887), .A2(n9871), .ZN(n8874) );
  INV_X1 U6483 ( .A(n9887), .ZN(n9885) );
  INV_X1 U6484 ( .A(n8184), .ZN(n8900) );
  INV_X1 U6485 ( .A(n8098), .ZN(n8934) );
  AND2_X1 U6486 ( .A1(n6447), .A2(n6446), .ZN(n9873) );
  NAND2_X1 U6487 ( .A1(n6439), .A2(n6746), .ZN(n6613) );
  INV_X1 U6488 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7517) );
  INV_X1 U6489 ( .A(n8566), .ZN(n6777) );
  INV_X1 U6490 ( .A(n9491), .ZN(n9349) );
  NAND2_X1 U6491 ( .A1(n9030), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9631) );
  INV_X1 U6492 ( .A(n9102), .ZN(n9623) );
  AND2_X1 U6493 ( .A1(n5717), .A2(n7333), .ZN(n9113) );
  OR2_X1 U6494 ( .A1(n6554), .A2(n6551), .ZN(n9686) );
  INV_X1 U6495 ( .A(n9364), .ZN(n9429) );
  AND2_X2 U6496 ( .A1(n7007), .A2(n7333), .ZN(n9433) );
  INV_X1 U6497 ( .A(n9355), .ZN(n9404) );
  INV_X1 U6498 ( .A(n9381), .ZN(n9211) );
  INV_X1 U6499 ( .A(n8073), .ZN(n9524) );
  AND2_X2 U6500 ( .A1(n6467), .A2(n6466), .ZN(n9757) );
  INV_X1 U6501 ( .A(n9202), .ZN(n9532) );
  INV_X1 U6502 ( .A(n9294), .ZN(n9552) );
  INV_X1 U6503 ( .A(n8078), .ZN(n9576) );
  NAND2_X1 U6504 ( .A1(n7006), .A2(n6467), .ZN(n9747) );
  INV_X2 U6505 ( .A(n9747), .ZN(n9749) );
  INV_X1 U6506 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7573) );
  INV_X1 U6507 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6631) );
  INV_X1 U6508 ( .A(n8621), .ZN(P2_U3893) );
  INV_X2 U6509 ( .A(n9141), .ZN(P1_U3973) );
  INV_X1 U6510 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n4959) );
  NAND2_X1 U6511 ( .A1(n4962), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4963) );
  MUX2_X1 U6512 ( .A(P1_IR_REG_31__SCAN_IN), .B(n4963), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n4964) );
  NAND2_X1 U6513 ( .A1(n4381), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4966) );
  XNOR2_X2 U6514 ( .A(n4966), .B(n4965), .ZN(n7686) );
  INV_X1 U6515 ( .A(n7686), .ZN(n4967) );
  NAND2_X2 U6516 ( .A1(n5700), .A2(n4968), .ZN(n6463) );
  NOR2_X1 U6517 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n5363) );
  NOR2_X1 U6518 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n4970) );
  INV_X1 U6519 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n4969) );
  AND4_X1 U6520 ( .A1(n4979), .A2(n5363), .A3(n4970), .A4(n4969), .ZN(n4971)
         );
  NAND2_X1 U6521 ( .A1(n4978), .A2(n4971), .ZN(n5411) );
  INV_X1 U6522 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n4974) );
  XNOR2_X2 U6523 ( .A(n4976), .B(n4975), .ZN(n7928) );
  OR2_X1 U6524 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(n4981), .ZN(n4982) );
  OR2_X1 U6525 ( .A1(n5297), .A2(n4981), .ZN(n4984) );
  NAND2_X1 U6526 ( .A1(n6463), .A2(n4987), .ZN(n5229) );
  NAND2_X1 U6527 ( .A1(n4988), .A2(n5781), .ZN(n4989) );
  NAND2_X4 U6528 ( .A1(n4989), .A2(n6463), .ZN(n8031) );
  XNOR2_X2 U6529 ( .A(n4991), .B(n5009), .ZN(n5726) );
  NAND2_X1 U6530 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), 
        .ZN(n4992) );
  NAND2_X1 U6531 ( .A1(n7999), .A2(n4994), .ZN(n4996) );
  NAND2_X1 U6532 ( .A1(n4997), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n4998) );
  BUF_X4 U6533 ( .A(n4999), .Z(n6053) );
  INV_X1 U6534 ( .A(SI_1_), .ZN(n5002) );
  AND2_X1 U6535 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5003) );
  NAND2_X1 U6536 ( .A1(n4999), .A2(n5003), .ZN(n5036) );
  AND2_X1 U6537 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n5004) );
  NAND2_X1 U6538 ( .A1(n7825), .A2(n5004), .ZN(n6088) );
  NAND2_X1 U6539 ( .A1(n5036), .A2(n6088), .ZN(n5055) );
  XNOR2_X1 U6540 ( .A(n5056), .B(n5055), .ZN(n6498) );
  OR2_X1 U6541 ( .A1(n5111), .A2(n6498), .ZN(n5008) );
  INV_X1 U6542 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6488) );
  INV_X2 U6543 ( .A(n5038), .ZN(n5486) );
  NAND2_X1 U6544 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5005) );
  NAND2_X1 U6545 ( .A1(n5486), .A2(n9145), .ZN(n5006) );
  XNOR2_X2 U6546 ( .A(n5012), .B(n5011), .ZN(n7987) );
  NAND2_X1 U6547 ( .A1(n4356), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5020) );
  NAND2_X1 U6548 ( .A1(n5303), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5019) );
  INV_X1 U6549 ( .A(n7987), .ZN(n5016) );
  NAND2_X1 U6550 ( .A1(n5098), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5018) );
  AND2_X2 U6551 ( .A1(n6463), .A2(n7066), .ZN(n5217) );
  NAND2_X1 U6552 ( .A1(n5737), .A2(n5217), .ZN(n5022) );
  NAND2_X1 U6553 ( .A1(n5023), .A2(n5022), .ZN(n5024) );
  INV_X2 U6554 ( .A(n5229), .ZN(n8034) );
  XNOR2_X1 U6555 ( .A(n5024), .B(n8034), .ZN(n5028) );
  INV_X1 U6556 ( .A(n5028), .ZN(n5026) );
  AOI22_X1 U6557 ( .A1(n5737), .A2(n5677), .B1(n7072), .B2(n8030), .ZN(n5027)
         );
  INV_X1 U6558 ( .A(n5027), .ZN(n5025) );
  NAND2_X1 U6559 ( .A1(n5026), .A2(n5025), .ZN(n5029) );
  NAND2_X1 U6560 ( .A1(n5028), .A2(n5027), .ZN(n6675) );
  NAND2_X1 U6561 ( .A1(n5029), .A2(n6675), .ZN(n6638) );
  INV_X1 U6562 ( .A(n6638), .ZN(n5048) );
  INV_X1 U6563 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n5040) );
  NAND2_X1 U6564 ( .A1(n5099), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5033) );
  NAND2_X1 U6565 ( .A1(n4358), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5032) );
  NAND2_X1 U6566 ( .A1(n5098), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5031) );
  NAND2_X1 U6567 ( .A1(n4356), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5030) );
  NAND2_X1 U6568 ( .A1(n5736), .A2(n8030), .ZN(n5039) );
  INV_X1 U6569 ( .A(SI_0_), .ZN(n5035) );
  INV_X1 U6570 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5034) );
  OAI21_X1 U6571 ( .B1(n7825), .B2(n5035), .A(n5034), .ZN(n5037) );
  AND2_X1 U6572 ( .A1(n5037), .A2(n5036), .ZN(n9592) );
  MUX2_X1 U6573 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9592), .S(n5038), .Z(n7013) );
  NAND2_X1 U6574 ( .A1(n7013), .A2(n8036), .ZN(n5044) );
  OAI211_X1 U6575 ( .C1(n5040), .C2(n6463), .A(n5039), .B(n5044), .ZN(n6622)
         );
  NAND2_X1 U6576 ( .A1(n5736), .A2(n5677), .ZN(n5043) );
  INV_X1 U6577 ( .A(n6463), .ZN(n5041) );
  AOI22_X1 U6578 ( .A1(n7013), .A2(n8030), .B1(n5041), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n5042) );
  NAND2_X1 U6579 ( .A1(n5043), .A2(n5042), .ZN(n6621) );
  NAND2_X1 U6580 ( .A1(n6622), .A2(n6621), .ZN(n5046) );
  NAND2_X1 U6581 ( .A1(n5044), .A2(n8034), .ZN(n5045) );
  NAND2_X1 U6582 ( .A1(n5046), .A2(n5045), .ZN(n6639) );
  NAND2_X1 U6583 ( .A1(n5048), .A2(n5047), .ZN(n6636) );
  NAND2_X1 U6584 ( .A1(n6636), .A2(n6675), .ZN(n5072) );
  NAND2_X1 U6585 ( .A1(n5099), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5052) );
  NAND2_X1 U6586 ( .A1(n4355), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5051) );
  NAND2_X1 U6587 ( .A1(n4357), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5050) );
  NAND2_X1 U6588 ( .A1(n5098), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5049) );
  INV_X1 U6589 ( .A(n5217), .ZN(n5173) );
  INV_X1 U6590 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6489) );
  OR2_X1 U6591 ( .A1(n5053), .A2(n5010), .ZN(n5106) );
  INV_X1 U6592 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5079) );
  INV_X1 U6593 ( .A(n5054), .ZN(n5064) );
  NAND2_X1 U6594 ( .A1(n5056), .A2(n5055), .ZN(n5059) );
  NAND2_X1 U6595 ( .A1(n5057), .A2(SI_1_), .ZN(n5058) );
  NAND2_X1 U6596 ( .A1(n5059), .A2(n5058), .ZN(n5087) );
  INV_X1 U6597 ( .A(SI_2_), .ZN(n5062) );
  XNOR2_X1 U6598 ( .A(n5088), .B(n5062), .ZN(n5086) );
  XNOR2_X1 U6599 ( .A(n5087), .B(n5086), .ZN(n6494) );
  OR2_X1 U6600 ( .A1(n5111), .A2(n6494), .ZN(n5063) );
  OAI22_X1 U6601 ( .A1(n7065), .A2(n5173), .B1(n5738), .B2(n5093), .ZN(n5065)
         );
  XNOR2_X1 U6602 ( .A(n5065), .B(n8034), .ZN(n5070) );
  OR2_X1 U6603 ( .A1(n7065), .A2(n8031), .ZN(n5068) );
  INV_X2 U6604 ( .A(n5066), .ZN(n8030) );
  NAND2_X1 U6605 ( .A1(n7142), .A2(n8030), .ZN(n5067) );
  AND2_X1 U6606 ( .A1(n5068), .A2(n5067), .ZN(n5069) );
  NAND2_X1 U6607 ( .A1(n5070), .A2(n5069), .ZN(n5073) );
  OR2_X1 U6608 ( .A1(n5070), .A2(n5069), .ZN(n5071) );
  AND2_X1 U6609 ( .A1(n5073), .A2(n5071), .ZN(n6677) );
  NAND2_X1 U6610 ( .A1(n5072), .A2(n6677), .ZN(n6678) );
  NAND2_X1 U6611 ( .A1(n6678), .A2(n5073), .ZN(n6707) );
  NAND2_X1 U6612 ( .A1(n4355), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5078) );
  INV_X1 U6613 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n7097) );
  NAND2_X1 U6614 ( .A1(n5099), .A2(n7097), .ZN(n5076) );
  NAND2_X1 U6615 ( .A1(n4357), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5075) );
  NAND2_X1 U6616 ( .A1(n5098), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5074) );
  AND3_X1 U6617 ( .A1(n5076), .A2(n5075), .A3(n5074), .ZN(n5077) );
  NAND2_X1 U6618 ( .A1(n5106), .A2(n5079), .ZN(n5080) );
  NAND2_X1 U6619 ( .A1(n5080), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5082) );
  INV_X1 U6620 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5081) );
  XNOR2_X1 U6621 ( .A(n5082), .B(n5081), .ZN(n6545) );
  INV_X1 U6622 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6490) );
  INV_X1 U6623 ( .A(SI_3_), .ZN(n5085) );
  NAND2_X1 U6624 ( .A1(n5087), .A2(n5086), .ZN(n5090) );
  NAND2_X1 U6625 ( .A1(n5088), .A2(SI_2_), .ZN(n5089) );
  XNOR2_X1 U6626 ( .A(n5112), .B(n5113), .ZN(n6492) );
  OR2_X1 U6627 ( .A1(n5111), .A2(n6492), .ZN(n5091) );
  OAI22_X1 U6628 ( .A1(n5741), .A2(n5173), .B1(n5740), .B2(n5148), .ZN(n5094)
         );
  XNOR2_X1 U6629 ( .A(n5094), .B(n8034), .ZN(n5126) );
  OR2_X1 U6630 ( .A1(n5741), .A2(n8031), .ZN(n5096) );
  NAND2_X1 U6631 ( .A1(n7098), .A2(n8030), .ZN(n5095) );
  NAND2_X1 U6632 ( .A1(n5096), .A2(n5095), .ZN(n5124) );
  XNOR2_X1 U6633 ( .A(n5126), .B(n5124), .ZN(n6708) );
  NAND2_X1 U6634 ( .A1(n6707), .A2(n6708), .ZN(n6706) );
  NAND2_X1 U6635 ( .A1(n4356), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5103) );
  NAND2_X1 U6636 ( .A1(n5098), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5102) );
  NAND2_X1 U6637 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5132) );
  OAI21_X1 U6638 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(n5132), .ZN(n6724) );
  INV_X1 U6639 ( .A(n6724), .ZN(n7078) );
  NAND2_X1 U6640 ( .A1(n5099), .A2(n7078), .ZN(n5101) );
  NAND2_X1 U6641 ( .A1(n4358), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5100) );
  OR2_X1 U6642 ( .A1(n5104), .A2(n5010), .ZN(n5105) );
  AND2_X1 U6643 ( .A1(n5106), .A2(n5105), .ZN(n5108) );
  INV_X1 U6644 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5107) );
  NAND2_X1 U6645 ( .A1(n5108), .A2(n5107), .ZN(n5138) );
  INV_X1 U6646 ( .A(n5108), .ZN(n5109) );
  NAND2_X1 U6647 ( .A1(n5109), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n5110) );
  NAND2_X1 U6648 ( .A1(n5138), .A2(n5110), .ZN(n6547) );
  NAND2_X1 U6649 ( .A1(n5114), .A2(SI_3_), .ZN(n5115) );
  INV_X1 U6650 ( .A(SI_4_), .ZN(n5118) );
  XNOR2_X1 U6651 ( .A(n5142), .B(n5141), .ZN(n6496) );
  OR2_X1 U6652 ( .A1(n5111), .A2(n6496), .ZN(n5120) );
  INV_X1 U6653 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6495) );
  OR2_X1 U6654 ( .A1(n5145), .A2(n6495), .ZN(n5119) );
  OAI211_X1 U6655 ( .C1(n5038), .C2(n6547), .A(n5120), .B(n5119), .ZN(n7079)
         );
  OAI22_X1 U6656 ( .A1(n7090), .A2(n5173), .B1(n6971), .B2(n5148), .ZN(n5121)
         );
  XNOR2_X1 U6657 ( .A(n5121), .B(n8034), .ZN(n5128) );
  OR2_X1 U6658 ( .A1(n7090), .A2(n8031), .ZN(n5123) );
  NAND2_X1 U6659 ( .A1(n7079), .A2(n8030), .ZN(n5122) );
  NAND2_X1 U6660 ( .A1(n5123), .A2(n5122), .ZN(n5129) );
  XNOR2_X1 U6661 ( .A(n5128), .B(n5129), .ZN(n6719) );
  INV_X1 U6662 ( .A(n5124), .ZN(n5125) );
  NAND2_X1 U6663 ( .A1(n5126), .A2(n5125), .ZN(n6717) );
  AND2_X1 U6664 ( .A1(n6719), .A2(n6717), .ZN(n5127) );
  INV_X1 U6665 ( .A(n5128), .ZN(n5130) );
  NAND2_X1 U6666 ( .A1(n5130), .A2(n5129), .ZN(n5153) );
  NAND2_X1 U6667 ( .A1(n4355), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5137) );
  NAND2_X1 U6668 ( .A1(n5098), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5136) );
  NOR2_X1 U6669 ( .A1(n5132), .A2(n5131), .ZN(n5158) );
  AND2_X1 U6670 ( .A1(n5132), .A2(n5131), .ZN(n5133) );
  NOR2_X1 U6671 ( .A1(n5158), .A2(n5133), .ZN(n7164) );
  NAND2_X1 U6672 ( .A1(n5099), .A2(n7164), .ZN(n5135) );
  NAND2_X1 U6673 ( .A1(n4358), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5134) );
  NAND2_X1 U6674 ( .A1(n5138), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5140) );
  INV_X1 U6675 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5139) );
  XNOR2_X1 U6676 ( .A(n5140), .B(n5139), .ZN(n6535) );
  MUX2_X1 U6677 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n6053), .Z(n5168) );
  INV_X1 U6678 ( .A(SI_5_), .ZN(n5144) );
  XNOR2_X1 U6679 ( .A(n5168), .B(n5144), .ZN(n5166) );
  XNOR2_X1 U6680 ( .A(n5167), .B(n5166), .ZN(n6501) );
  OR2_X1 U6681 ( .A1(n5111), .A2(n6501), .ZN(n5147) );
  INV_X1 U6682 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6502) );
  OR2_X1 U6683 ( .A1(n5145), .A2(n6502), .ZN(n5146) );
  OAI211_X1 U6684 ( .C1(n5038), .C2(n6535), .A(n5147), .B(n5146), .ZN(n7727)
         );
  OAI22_X1 U6685 ( .A1(n7728), .A2(n5173), .B1(n5744), .B2(n5148), .ZN(n5149)
         );
  XNOR2_X1 U6686 ( .A(n5149), .B(n8034), .ZN(n5154) );
  AND2_X1 U6687 ( .A1(n5153), .A2(n5154), .ZN(n5150) );
  NAND2_X1 U6688 ( .A1(n6718), .A2(n5150), .ZN(n6887) );
  OR2_X1 U6689 ( .A1(n7728), .A2(n8031), .ZN(n5152) );
  NAND2_X1 U6690 ( .A1(n7727), .A2(n8030), .ZN(n5151) );
  NAND2_X1 U6691 ( .A1(n5152), .A2(n5151), .ZN(n6890) );
  NAND2_X1 U6692 ( .A1(n6887), .A2(n6890), .ZN(n5157) );
  NAND2_X1 U6693 ( .A1(n6718), .A2(n5153), .ZN(n5156) );
  INV_X1 U6694 ( .A(n5154), .ZN(n5155) );
  NAND2_X1 U6695 ( .A1(n5156), .A2(n5155), .ZN(n6888) );
  NAND2_X1 U6696 ( .A1(n5157), .A2(n6888), .ZN(n6907) );
  NAND2_X1 U6697 ( .A1(n5098), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5163) );
  NAND2_X1 U6698 ( .A1(n4355), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5162) );
  NAND2_X1 U6699 ( .A1(n5158), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5182) );
  OR2_X1 U6700 ( .A1(n5158), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5159) );
  AND2_X1 U6701 ( .A1(n5182), .A2(n5159), .ZN(n7188) );
  NAND2_X1 U6702 ( .A1(n5099), .A2(n7188), .ZN(n5161) );
  NAND2_X1 U6703 ( .A1(n4357), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5160) );
  NAND2_X1 U6704 ( .A1(n5164), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5165) );
  XNOR2_X1 U6705 ( .A(n5165), .B(n4961), .ZN(n6555) );
  NAND2_X1 U6706 ( .A1(n5168), .A2(SI_5_), .ZN(n5169) );
  MUX2_X1 U6707 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n6053), .Z(n5190) );
  INV_X1 U6708 ( .A(SI_6_), .ZN(n5170) );
  XNOR2_X1 U6709 ( .A(n5190), .B(n5170), .ZN(n5188) );
  XNOR2_X1 U6710 ( .A(n5189), .B(n5188), .ZN(n6504) );
  OR2_X1 U6711 ( .A1(n5111), .A2(n6504), .ZN(n5172) );
  INV_X1 U6712 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6505) );
  OR2_X1 U6713 ( .A1(n5145), .A2(n6505), .ZN(n5171) );
  OAI211_X1 U6714 ( .C1(n5038), .C2(n6555), .A(n5172), .B(n5171), .ZN(n7723)
         );
  OAI22_X1 U6715 ( .A1(n7722), .A2(n5173), .B1(n4576), .B2(n5148), .ZN(n5174)
         );
  XNOR2_X1 U6716 ( .A(n5174), .B(n8034), .ZN(n5177) );
  OR2_X1 U6717 ( .A1(n7722), .A2(n8031), .ZN(n5176) );
  NAND2_X1 U6718 ( .A1(n7723), .A2(n8030), .ZN(n5175) );
  AND2_X1 U6719 ( .A1(n5176), .A2(n5175), .ZN(n5178) );
  NAND2_X1 U6720 ( .A1(n5177), .A2(n5178), .ZN(n6905) );
  NAND2_X1 U6721 ( .A1(n6907), .A2(n6905), .ZN(n5181) );
  INV_X1 U6722 ( .A(n5177), .ZN(n5180) );
  INV_X1 U6723 ( .A(n5178), .ZN(n5179) );
  NAND2_X1 U6724 ( .A1(n5180), .A2(n5179), .ZN(n6906) );
  NAND2_X1 U6725 ( .A1(n5181), .A2(n6906), .ZN(n6978) );
  NAND2_X1 U6726 ( .A1(n4355), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5187) );
  NAND2_X1 U6727 ( .A1(n5098), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5186) );
  NAND2_X1 U6728 ( .A1(n5182), .A2(n6982), .ZN(n5183) );
  AND2_X1 U6729 ( .A1(n5210), .A2(n5183), .ZN(n7113) );
  NAND2_X1 U6730 ( .A1(n5099), .A2(n7113), .ZN(n5185) );
  NAND2_X1 U6731 ( .A1(n4357), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5184) );
  NAND4_X1 U6732 ( .A1(n5187), .A2(n5186), .A3(n5185), .A4(n5184), .ZN(n9135)
         );
  NAND2_X1 U6733 ( .A1(n9135), .A2(n8030), .ZN(n5200) );
  NAND2_X1 U6734 ( .A1(n5189), .A2(n5188), .ZN(n5192) );
  NAND2_X1 U6735 ( .A1(n5190), .A2(SI_6_), .ZN(n5191) );
  MUX2_X1 U6736 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n6053), .Z(n5220) );
  INV_X1 U6737 ( .A(SI_7_), .ZN(n5193) );
  XNOR2_X1 U6738 ( .A(n5220), .B(n5193), .ZN(n5218) );
  XNOR2_X1 U6739 ( .A(n5219), .B(n5218), .ZN(n6513) );
  OR2_X1 U6740 ( .A1(n5111), .A2(n6513), .ZN(n5198) );
  INV_X1 U6741 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6514) );
  OR2_X1 U6742 ( .A1(n5145), .A2(n6514), .ZN(n5197) );
  NAND2_X1 U6743 ( .A1(n5194), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5195) );
  XNOR2_X1 U6744 ( .A(n5195), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6600) );
  NAND2_X1 U6745 ( .A1(n5486), .A2(n6600), .ZN(n5196) );
  NAND2_X1 U6746 ( .A1(n7116), .A2(n8036), .ZN(n5199) );
  NAND2_X1 U6747 ( .A1(n5200), .A2(n5199), .ZN(n5201) );
  XNOR2_X1 U6748 ( .A(n5201), .B(n8034), .ZN(n6976) );
  NAND2_X1 U6749 ( .A1(n9135), .A2(n5677), .ZN(n5203) );
  NAND2_X1 U6750 ( .A1(n7116), .A2(n8030), .ZN(n5202) );
  AND2_X1 U6751 ( .A1(n5203), .A2(n5202), .ZN(n5205) );
  NAND2_X1 U6752 ( .A1(n6976), .A2(n5205), .ZN(n5204) );
  NAND2_X1 U6753 ( .A1(n6978), .A2(n5204), .ZN(n5208) );
  INV_X1 U6754 ( .A(n6976), .ZN(n5206) );
  INV_X1 U6755 ( .A(n5205), .ZN(n6975) );
  NAND2_X1 U6756 ( .A1(n5206), .A2(n6975), .ZN(n5207) );
  NAND2_X1 U6757 ( .A1(n5208), .A2(n5207), .ZN(n5232) );
  NAND2_X1 U6758 ( .A1(n5098), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5216) );
  NAND2_X1 U6759 ( .A1(n4356), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5215) );
  NAND2_X1 U6760 ( .A1(n5210), .A2(n5209), .ZN(n5211) );
  NAND2_X1 U6761 ( .A1(n5238), .A2(n5211), .ZN(n7310) );
  INV_X1 U6762 ( .A(n7310), .ZN(n5212) );
  NAND2_X1 U6763 ( .A1(n5099), .A2(n5212), .ZN(n5214) );
  NAND2_X1 U6764 ( .A1(n4358), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5213) );
  OR2_X1 U6765 ( .A1(n4978), .A2(n5010), .ZN(n5252) );
  INV_X1 U6766 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5251) );
  XNOR2_X1 U6767 ( .A(n5252), .B(n5251), .ZN(n6604) );
  NAND2_X1 U6768 ( .A1(n5219), .A2(n5218), .ZN(n5222) );
  NAND2_X1 U6769 ( .A1(n5220), .A2(SI_7_), .ZN(n5221) );
  INV_X1 U6770 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6523) );
  MUX2_X1 U6771 ( .A(n6523), .B(n6522), .S(n6053), .Z(n5223) );
  INV_X1 U6772 ( .A(SI_8_), .ZN(n10128) );
  NAND2_X1 U6773 ( .A1(n5223), .A2(n10128), .ZN(n5246) );
  INV_X1 U6774 ( .A(n5223), .ZN(n5224) );
  NAND2_X1 U6775 ( .A1(n5224), .A2(SI_8_), .ZN(n5225) );
  NAND2_X1 U6776 ( .A1(n5246), .A2(n5225), .ZN(n5244) );
  INV_X1 U6777 ( .A(n5244), .ZN(n5226) );
  OR2_X1 U6778 ( .A1(n5145), .A2(n6522), .ZN(n5227) );
  OAI211_X1 U6779 ( .C1(n5038), .C2(n6604), .A(n5228), .B(n5227), .ZN(n7292)
         );
  OAI22_X1 U6780 ( .A1(n7385), .A2(n5173), .B1(n7309), .B2(n5148), .ZN(n5230)
         );
  XNOR2_X1 U6781 ( .A(n5230), .B(n5675), .ZN(n5231) );
  OR2_X1 U6782 ( .A1(n7385), .A2(n8031), .ZN(n5234) );
  NAND2_X1 U6783 ( .A1(n7292), .A2(n8030), .ZN(n5233) );
  NAND2_X1 U6784 ( .A1(n5234), .A2(n5233), .ZN(n7286) );
  NAND2_X1 U6785 ( .A1(n7283), .A2(n5236), .ZN(n7381) );
  NAND2_X1 U6786 ( .A1(n4355), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5243) );
  NAND2_X1 U6787 ( .A1(n5098), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5242) );
  AND2_X1 U6788 ( .A1(n5238), .A2(n5237), .ZN(n5239) );
  NOR2_X1 U6789 ( .A1(n5264), .A2(n5239), .ZN(n7387) );
  NAND2_X1 U6790 ( .A1(n5099), .A2(n7387), .ZN(n5241) );
  NAND2_X1 U6791 ( .A1(n4357), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5240) );
  INV_X1 U6792 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n5247) );
  MUX2_X1 U6793 ( .A(n6590), .B(n5247), .S(n6053), .Z(n5248) );
  NAND2_X1 U6794 ( .A1(n5248), .A2(n9991), .ZN(n5272) );
  INV_X1 U6795 ( .A(n5248), .ZN(n5249) );
  NAND2_X1 U6796 ( .A1(n5249), .A2(SI_9_), .ZN(n5250) );
  NAND2_X1 U6797 ( .A1(n6165), .A2(n7830), .ZN(n5256) );
  NAND2_X1 U6798 ( .A1(n5252), .A2(n5251), .ZN(n5253) );
  NAND2_X1 U6799 ( .A1(n5253), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5254) );
  XNOR2_X1 U6800 ( .A(n5254), .B(P1_IR_REG_9__SCAN_IN), .ZN(n9611) );
  AOI22_X1 U6801 ( .A1(n5487), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5486), .B2(
        n9611), .ZN(n5255) );
  NAND2_X1 U6802 ( .A1(n5256), .A2(n5255), .ZN(n7157) );
  OAI22_X1 U6803 ( .A1(n7324), .A2(n5173), .B1(n7390), .B2(n5148), .ZN(n5257)
         );
  XNOR2_X1 U6804 ( .A(n5257), .B(n8034), .ZN(n5262) );
  OR2_X1 U6805 ( .A1(n7324), .A2(n8031), .ZN(n5259) );
  NAND2_X1 U6806 ( .A1(n7157), .A2(n8030), .ZN(n5258) );
  NAND2_X1 U6807 ( .A1(n5259), .A2(n5258), .ZN(n5260) );
  XNOR2_X1 U6808 ( .A(n5262), .B(n5260), .ZN(n7382) );
  NAND2_X1 U6809 ( .A1(n7381), .A2(n7382), .ZN(n7380) );
  INV_X1 U6810 ( .A(n5260), .ZN(n5261) );
  NAND2_X1 U6811 ( .A1(n5262), .A2(n5261), .ZN(n5263) );
  NAND2_X1 U6812 ( .A1(n7380), .A2(n5263), .ZN(n5282) );
  INV_X1 U6813 ( .A(n5282), .ZN(n5280) );
  NAND2_X1 U6814 ( .A1(n5097), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5270) );
  NAND2_X1 U6815 ( .A1(n5264), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5301) );
  OR2_X1 U6816 ( .A1(n5264), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5265) );
  NAND2_X1 U6817 ( .A1(n5301), .A2(n5265), .ZN(n9632) );
  INV_X1 U6818 ( .A(n9632), .ZN(n5266) );
  NAND2_X1 U6819 ( .A1(n5099), .A2(n5266), .ZN(n5269) );
  NAND2_X1 U6820 ( .A1(n4358), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5268) );
  NAND2_X1 U6821 ( .A1(n5098), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5267) );
  MUX2_X1 U6822 ( .A(n6610), .B(n6594), .S(n6491), .Z(n5290) );
  XNOR2_X1 U6823 ( .A(n5290), .B(SI_10_), .ZN(n5287) );
  NAND2_X1 U6824 ( .A1(n6593), .A2(n7830), .ZN(n5276) );
  OR2_X1 U6825 ( .A1(n5273), .A2(n5010), .ZN(n5274) );
  XNOR2_X1 U6826 ( .A(n5274), .B(P1_IR_REG_10__SCAN_IN), .ZN(n9601) );
  AOI22_X1 U6827 ( .A1(n5487), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5486), .B2(
        n9601), .ZN(n5275) );
  NAND2_X1 U6828 ( .A1(n9629), .A2(n8036), .ZN(n5277) );
  OAI21_X1 U6829 ( .B1(n7431), .B2(n5173), .A(n5277), .ZN(n5278) );
  XNOR2_X1 U6830 ( .A(n5278), .B(n8034), .ZN(n5281) );
  INV_X1 U6831 ( .A(n5281), .ZN(n5279) );
  OR2_X1 U6832 ( .A1(n7431), .A2(n8031), .ZN(n5284) );
  NAND2_X1 U6833 ( .A1(n9629), .A2(n8030), .ZN(n5283) );
  NAND2_X1 U6834 ( .A1(n5284), .A2(n5283), .ZN(n9621) );
  INV_X1 U6835 ( .A(n9621), .ZN(n5285) );
  NAND2_X1 U6836 ( .A1(n9625), .A2(n5286), .ZN(n7597) );
  INV_X1 U6837 ( .A(n5287), .ZN(n5288) );
  INV_X1 U6838 ( .A(n5290), .ZN(n5291) );
  NAND2_X1 U6839 ( .A1(n5291), .A2(SI_10_), .ZN(n5292) );
  INV_X1 U6840 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n5293) );
  MUX2_X1 U6841 ( .A(n5293), .B(n6631), .S(n6491), .Z(n5294) );
  NAND2_X1 U6842 ( .A1(n5294), .A2(n10014), .ZN(n5313) );
  INV_X1 U6843 ( .A(n5294), .ZN(n5295) );
  NAND2_X1 U6844 ( .A1(n5295), .A2(SI_11_), .ZN(n5296) );
  NAND2_X1 U6845 ( .A1(n5313), .A2(n5296), .ZN(n5314) );
  XNOR2_X1 U6846 ( .A(n5315), .B(n5314), .ZN(n6627) );
  NAND2_X1 U6847 ( .A1(n6627), .A2(n7830), .ZN(n5300) );
  INV_X1 U6848 ( .A(n5297), .ZN(n5316) );
  OR2_X1 U6849 ( .A1(n5316), .A2(n5010), .ZN(n5298) );
  XNOR2_X1 U6850 ( .A(n5298), .B(P1_IR_REG_11__SCAN_IN), .ZN(n9641) );
  AOI22_X1 U6851 ( .A1(n5487), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5486), .B2(
        n9641), .ZN(n5299) );
  NAND2_X1 U6852 ( .A1(n7446), .A2(n8036), .ZN(n5309) );
  NAND2_X1 U6853 ( .A1(n4356), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5307) );
  NAND2_X1 U6854 ( .A1(n5301), .A2(n7602), .ZN(n5302) );
  AND2_X1 U6855 ( .A1(n5322), .A2(n5302), .ZN(n7605) );
  NAND2_X1 U6856 ( .A1(n5099), .A2(n7605), .ZN(n5306) );
  NAND2_X1 U6857 ( .A1(n4358), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5305) );
  NAND2_X1 U6858 ( .A1(n5098), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5304) );
  OR2_X1 U6859 ( .A1(n7460), .A2(n5173), .ZN(n5308) );
  NAND2_X1 U6860 ( .A1(n5309), .A2(n5308), .ZN(n5310) );
  XNOR2_X1 U6861 ( .A(n5310), .B(n8034), .ZN(n5312) );
  INV_X1 U6862 ( .A(n7460), .ZN(n9131) );
  AOI22_X1 U6863 ( .A1(n7446), .A2(n8030), .B1(n5677), .B2(n9131), .ZN(n5311)
         );
  OR2_X1 U6864 ( .A1(n5312), .A2(n5311), .ZN(n7599) );
  NAND2_X1 U6865 ( .A1(n5312), .A2(n5311), .ZN(n7598) );
  MUX2_X1 U6866 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n6491), .Z(n5336) );
  XNOR2_X1 U6867 ( .A(n5336), .B(n9989), .ZN(n5335) );
  XNOR2_X1 U6868 ( .A(n5337), .B(n5335), .ZN(n6673) );
  NAND2_X1 U6869 ( .A1(n6673), .A2(n7830), .ZN(n5320) );
  NAND2_X1 U6870 ( .A1(n5316), .A2(n4810), .ZN(n5365) );
  NAND2_X1 U6871 ( .A1(n5365), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5317) );
  NAND2_X1 U6872 ( .A1(n5317), .A2(n4809), .ZN(n5339) );
  OR2_X1 U6873 ( .A1(n5317), .A2(n4809), .ZN(n5318) );
  AOI22_X1 U6874 ( .A1(n5487), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5486), .B2(
        n8014), .ZN(n5319) );
  NAND2_X1 U6875 ( .A1(n7628), .A2(n8036), .ZN(n5329) );
  NAND2_X1 U6876 ( .A1(n5098), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5327) );
  NAND2_X1 U6877 ( .A1(n4355), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5326) );
  AND2_X1 U6878 ( .A1(n5322), .A2(n5321), .ZN(n5323) );
  NOR2_X1 U6879 ( .A1(n5343), .A2(n5323), .ZN(n7623) );
  NAND2_X1 U6880 ( .A1(n5099), .A2(n7623), .ZN(n5325) );
  NAND2_X1 U6881 ( .A1(n4358), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5324) );
  OR2_X1 U6882 ( .A1(n7531), .A2(n5173), .ZN(n5328) );
  NAND2_X1 U6883 ( .A1(n5329), .A2(n5328), .ZN(n5330) );
  XNOR2_X1 U6884 ( .A(n5330), .B(n5675), .ZN(n5332) );
  NOR2_X1 U6885 ( .A1(n7531), .A2(n8031), .ZN(n5331) );
  AOI21_X1 U6886 ( .B1(n7628), .B2(n8030), .A(n5331), .ZN(n5333) );
  XNOR2_X1 U6887 ( .A(n5332), .B(n5333), .ZN(n7622) );
  INV_X1 U6888 ( .A(n5332), .ZN(n5334) );
  MUX2_X1 U6889 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n6491), .Z(n5358) );
  XNOR2_X1 U6890 ( .A(n5358), .B(SI_13_), .ZN(n5338) );
  XNOR2_X1 U6891 ( .A(n5362), .B(n5338), .ZN(n6689) );
  NAND2_X1 U6892 ( .A1(n6689), .A2(n7830), .ZN(n5342) );
  NAND2_X1 U6893 ( .A1(n5339), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5340) );
  AOI22_X1 U6894 ( .A1(n5487), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n5486), .B2(
        n9653), .ZN(n5341) );
  NAND2_X1 U6895 ( .A1(n9066), .A2(n8036), .ZN(n5350) );
  NAND2_X1 U6896 ( .A1(n4355), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5348) );
  NAND2_X1 U6897 ( .A1(n4357), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5347) );
  NAND2_X1 U6898 ( .A1(n5343), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n5371) );
  OR2_X1 U6899 ( .A1(n5343), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n5344) );
  AND2_X1 U6900 ( .A1(n5371), .A2(n5344), .ZN(n9061) );
  NAND2_X1 U6901 ( .A1(n5099), .A2(n9061), .ZN(n5346) );
  NAND2_X1 U6902 ( .A1(n5098), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5345) );
  OR2_X1 U6903 ( .A1(n9413), .A2(n5173), .ZN(n5349) );
  NAND2_X1 U6904 ( .A1(n5350), .A2(n5349), .ZN(n5351) );
  XNOR2_X1 U6905 ( .A(n5351), .B(n5675), .ZN(n5353) );
  NOR2_X1 U6906 ( .A1(n9413), .A2(n8031), .ZN(n5352) );
  AOI21_X1 U6907 ( .B1(n9066), .B2(n8030), .A(n5352), .ZN(n5354) );
  XNOR2_X1 U6908 ( .A(n5353), .B(n5354), .ZN(n9060) );
  NAND2_X1 U6909 ( .A1(n9059), .A2(n9060), .ZN(n5357) );
  INV_X1 U6910 ( .A(n5353), .ZN(n5355) );
  NAND2_X1 U6911 ( .A1(n5355), .A2(n5354), .ZN(n5356) );
  NOR2_X1 U6912 ( .A1(n5359), .A2(n10110), .ZN(n5361) );
  NAND2_X1 U6913 ( .A1(n5359), .A2(n10110), .ZN(n5360) );
  MUX2_X1 U6914 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n6491), .Z(n5385) );
  XNOR2_X1 U6915 ( .A(n5385), .B(n5386), .ZN(n5383) );
  XNOR2_X1 U6916 ( .A(n5384), .B(n5383), .ZN(n6773) );
  NAND2_X1 U6917 ( .A1(n6773), .A2(n7830), .ZN(n5369) );
  INV_X1 U6918 ( .A(n5363), .ZN(n5364) );
  OAI21_X1 U6919 ( .B1(n5365), .B2(n5364), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5366) );
  MUX2_X1 U6920 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5366), .S(
        P1_IR_REG_14__SCAN_IN), .Z(n5367) );
  AOI22_X1 U6921 ( .A1(n5487), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5486), .B2(
        n9665), .ZN(n5368) );
  NAND2_X1 U6922 ( .A1(n9425), .A2(n8036), .ZN(n5378) );
  NAND2_X1 U6923 ( .A1(n4356), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5376) );
  NAND2_X1 U6924 ( .A1(n5098), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5375) );
  NAND2_X1 U6925 ( .A1(n5371), .A2(n5370), .ZN(n5372) );
  AND2_X1 U6926 ( .A1(n5416), .A2(n5372), .ZN(n9427) );
  NAND2_X1 U6927 ( .A1(n5099), .A2(n9427), .ZN(n5374) );
  NAND2_X1 U6928 ( .A1(n4357), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5373) );
  OR2_X1 U6929 ( .A1(n9107), .A2(n5173), .ZN(n5377) );
  NAND2_X1 U6930 ( .A1(n5378), .A2(n5377), .ZN(n5379) );
  XNOR2_X1 U6931 ( .A(n5379), .B(n5675), .ZN(n5428) );
  INV_X1 U6932 ( .A(n5428), .ZN(n9011) );
  NAND2_X1 U6933 ( .A1(n9425), .A2(n8030), .ZN(n5381) );
  OR2_X1 U6934 ( .A1(n9107), .A2(n8031), .ZN(n5380) );
  NAND2_X1 U6935 ( .A1(n5381), .A2(n5380), .ZN(n8964) );
  INV_X1 U6936 ( .A(n8964), .ZN(n5382) );
  AND2_X1 U6937 ( .A1(n9011), .A2(n5382), .ZN(n5432) );
  NAND2_X1 U6938 ( .A1(n5384), .A2(n5383), .ZN(n5389) );
  INV_X1 U6939 ( .A(n5385), .ZN(n5387) );
  NAND2_X1 U6940 ( .A1(n5387), .A2(n5386), .ZN(n5388) );
  NAND2_X1 U6941 ( .A1(n5389), .A2(n5388), .ZN(n5407) );
  MUX2_X1 U6942 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n6491), .Z(n5409) );
  NOR2_X1 U6943 ( .A1(n5409), .A2(SI_15_), .ZN(n5391) );
  NAND2_X1 U6944 ( .A1(n5409), .A2(SI_15_), .ZN(n5390) );
  OAI21_X2 U6945 ( .B1(n5407), .B2(n5391), .A(n5390), .ZN(n5441) );
  MUX2_X1 U6946 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .S(n6491), .Z(n5439) );
  XNOR2_X1 U6947 ( .A(n5439), .B(SI_16_), .ZN(n5392) );
  XNOR2_X1 U6948 ( .A(n5441), .B(n5392), .ZN(n7017) );
  NAND2_X1 U6949 ( .A1(n7017), .A2(n7830), .ZN(n5396) );
  NAND2_X1 U6950 ( .A1(n5393), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5394) );
  XNOR2_X1 U6951 ( .A(n5394), .B(P1_IR_REG_16__SCAN_IN), .ZN(n8012) );
  AOI22_X1 U6952 ( .A1(n5487), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n5486), .B2(
        n8012), .ZN(n5395) );
  NAND2_X1 U6953 ( .A1(n9399), .A2(n8036), .ZN(n5403) );
  NAND2_X1 U6954 ( .A1(n5098), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5401) );
  NAND2_X1 U6955 ( .A1(n4355), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n5400) );
  NOR2_X1 U6956 ( .A1(n5418), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5397) );
  NAND2_X1 U6957 ( .A1(n5099), .A2(n4944), .ZN(n5399) );
  NAND2_X1 U6958 ( .A1(n4358), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5398) );
  OR2_X1 U6959 ( .A1(n9373), .A2(n5173), .ZN(n5402) );
  NAND2_X1 U6960 ( .A1(n5403), .A2(n5402), .ZN(n5404) );
  XNOR2_X1 U6961 ( .A(n5404), .B(n5675), .ZN(n9017) );
  NAND2_X1 U6962 ( .A1(n9399), .A2(n8030), .ZN(n5406) );
  OR2_X1 U6963 ( .A1(n9373), .A2(n8031), .ZN(n5405) );
  NAND2_X1 U6964 ( .A1(n5406), .A2(n5405), .ZN(n9018) );
  NAND2_X1 U6965 ( .A1(n9017), .A2(n9018), .ZN(n9016) );
  INV_X1 U6966 ( .A(n9016), .ZN(n5431) );
  INV_X1 U6967 ( .A(SI_15_), .ZN(n5408) );
  XNOR2_X1 U6968 ( .A(n5409), .B(n5408), .ZN(n5410) );
  XNOR2_X1 U6969 ( .A(n5407), .B(n5410), .ZN(n6778) );
  NAND2_X1 U6970 ( .A1(n6778), .A2(n7830), .ZN(n5414) );
  NAND2_X1 U6971 ( .A1(n5411), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5412) );
  XNOR2_X1 U6972 ( .A(n5412), .B(P1_IR_REG_15__SCAN_IN), .ZN(n9678) );
  AOI22_X1 U6973 ( .A1(n5487), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n5486), .B2(
        n9678), .ZN(n5413) );
  NAND2_X1 U6974 ( .A1(n9514), .A2(n8036), .ZN(n5424) );
  NAND2_X1 U6975 ( .A1(n5098), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5422) );
  NAND2_X1 U6976 ( .A1(n4355), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5421) );
  AND2_X1 U6977 ( .A1(n5416), .A2(n5415), .ZN(n5417) );
  NOR2_X1 U6978 ( .A1(n5418), .A2(n5417), .ZN(n9110) );
  NAND2_X1 U6979 ( .A1(n5099), .A2(n9110), .ZN(n5420) );
  NAND2_X1 U6980 ( .A1(n4357), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5419) );
  NAND4_X1 U6981 ( .A1(n5422), .A2(n5421), .A3(n5420), .A4(n5419), .ZN(n9392)
         );
  NAND2_X1 U6982 ( .A1(n9392), .A2(n8030), .ZN(n5423) );
  NAND2_X1 U6983 ( .A1(n5424), .A2(n5423), .ZN(n5425) );
  XNOR2_X1 U6984 ( .A(n5425), .B(n5675), .ZN(n9014) );
  NAND2_X1 U6985 ( .A1(n9514), .A2(n8030), .ZN(n5427) );
  NAND2_X1 U6986 ( .A1(n9392), .A2(n5677), .ZN(n5426) );
  NAND2_X1 U6987 ( .A1(n5427), .A2(n5426), .ZN(n9013) );
  AOI22_X1 U6988 ( .A1(n9014), .A2(n9013), .B1(n5428), .B2(n8964), .ZN(n5429)
         );
  INV_X1 U6989 ( .A(n9017), .ZN(n5435) );
  OAI21_X1 U6990 ( .B1(n9014), .B2(n9013), .A(n9018), .ZN(n5434) );
  NOR2_X1 U6991 ( .A1(n9018), .A2(n9013), .ZN(n5433) );
  INV_X1 U6992 ( .A(n9014), .ZN(n9012) );
  AOI22_X1 U6993 ( .A1(n5435), .A2(n5434), .B1(n5433), .B2(n9012), .ZN(n5436)
         );
  INV_X1 U6994 ( .A(n5439), .ZN(n5438) );
  INV_X1 U6995 ( .A(SI_16_), .ZN(n5437) );
  MUX2_X1 U6996 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .S(n6491), .Z(n5462) );
  XNOR2_X1 U6997 ( .A(n5462), .B(n10045), .ZN(n5460) );
  XNOR2_X1 U6998 ( .A(n5461), .B(n5460), .ZN(n7026) );
  NAND2_X1 U6999 ( .A1(n7026), .A2(n7830), .ZN(n5444) );
  XNOR2_X1 U7000 ( .A(n5442), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9700) );
  AOI22_X1 U7001 ( .A1(n5487), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n5486), .B2(
        n9700), .ZN(n5443) );
  NAND2_X1 U7002 ( .A1(n9504), .A2(n8036), .ZN(n5451) );
  NAND2_X1 U7003 ( .A1(n5098), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5449) );
  NAND2_X1 U7004 ( .A1(n4356), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n5448) );
  OR2_X1 U7005 ( .A1(n9031), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n5445) );
  AND2_X1 U7006 ( .A1(n5490), .A2(n5445), .ZN(n9377) );
  NAND2_X1 U7007 ( .A1(n5099), .A2(n9377), .ZN(n5447) );
  NAND2_X1 U7008 ( .A1(n4357), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5446) );
  NAND4_X1 U7009 ( .A1(n5449), .A2(n5448), .A3(n5447), .A4(n5446), .ZN(n9391)
         );
  NAND2_X1 U7010 ( .A1(n9391), .A2(n8030), .ZN(n5450) );
  NAND2_X1 U7011 ( .A1(n5451), .A2(n5450), .ZN(n5452) );
  XNOR2_X1 U7012 ( .A(n5452), .B(n5675), .ZN(n5455) );
  NAND2_X1 U7013 ( .A1(n9504), .A2(n8030), .ZN(n5454) );
  NAND2_X1 U7014 ( .A1(n9391), .A2(n5677), .ZN(n5453) );
  NAND2_X1 U7015 ( .A1(n5454), .A2(n5453), .ZN(n5456) );
  NAND2_X1 U7016 ( .A1(n5455), .A2(n5456), .ZN(n9027) );
  INV_X1 U7017 ( .A(n5455), .ZN(n5458) );
  INV_X1 U7018 ( .A(n5456), .ZN(n5457) );
  NAND2_X1 U7019 ( .A1(n5458), .A2(n5457), .ZN(n9026) );
  NAND2_X1 U7020 ( .A1(n5459), .A2(n9026), .ZN(n8980) );
  INV_X1 U7021 ( .A(n5462), .ZN(n5463) );
  MUX2_X1 U7022 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n6491), .Z(n5464) );
  OAI21_X1 U7023 ( .B1(n5464), .B2(SI_18_), .A(n5465), .ZN(n5478) );
  NAND2_X1 U7024 ( .A1(n5481), .A2(n5465), .ZN(n5510) );
  MUX2_X1 U7025 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(P2_DATAO_REG_19__SCAN_IN), 
        .S(n6491), .Z(n5514) );
  XNOR2_X1 U7026 ( .A(n5514), .B(SI_19_), .ZN(n5511) );
  XNOR2_X1 U7027 ( .A(n5510), .B(n5511), .ZN(n7305) );
  NAND2_X1 U7028 ( .A1(n7305), .A2(n7830), .ZN(n5467) );
  AOI22_X1 U7029 ( .A1(n5487), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n7875), .B2(
        n5486), .ZN(n5466) );
  NAND2_X1 U7030 ( .A1(n9491), .A2(n8036), .ZN(n5474) );
  NAND2_X1 U7031 ( .A1(n5097), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n5472) );
  NAND2_X1 U7032 ( .A1(n5098), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n5471) );
  NAND2_X1 U7033 ( .A1(n5492), .A2(n8987), .ZN(n5468) );
  AND2_X1 U7034 ( .A1(n5521), .A2(n5468), .ZN(n9346) );
  NAND2_X1 U7035 ( .A1(n5099), .A2(n9346), .ZN(n5470) );
  NAND2_X1 U7036 ( .A1(n4357), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5469) );
  NAND4_X1 U7037 ( .A1(n5472), .A2(n5471), .A3(n5470), .A4(n5469), .ZN(n9125)
         );
  NAND2_X1 U7038 ( .A1(n9125), .A2(n8030), .ZN(n5473) );
  NAND2_X1 U7039 ( .A1(n5474), .A2(n5473), .ZN(n5475) );
  XNOR2_X1 U7040 ( .A(n5475), .B(n5675), .ZN(n8983) );
  NAND2_X1 U7041 ( .A1(n9491), .A2(n5217), .ZN(n5477) );
  NAND2_X1 U7042 ( .A1(n9125), .A2(n5677), .ZN(n5476) );
  NAND2_X1 U7043 ( .A1(n5477), .A2(n5476), .ZN(n8982) );
  NAND2_X1 U7044 ( .A1(n5479), .A2(n5478), .ZN(n5480) );
  AND2_X1 U7045 ( .A1(n5481), .A2(n5480), .ZN(n7120) );
  NAND2_X1 U7046 ( .A1(n7120), .A2(n7830), .ZN(n5489) );
  OR2_X1 U7047 ( .A1(n5483), .A2(n5482), .ZN(n5484) );
  AND2_X1 U7048 ( .A1(n5485), .A2(n5484), .ZN(n9706) );
  AOI22_X1 U7049 ( .A1(n5487), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n5486), .B2(
        n9706), .ZN(n5488) );
  NAND2_X1 U7050 ( .A1(n4355), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n5496) );
  NAND2_X1 U7051 ( .A1(n5098), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n5495) );
  NAND2_X1 U7052 ( .A1(n5490), .A2(n9083), .ZN(n5491) );
  AND2_X1 U7053 ( .A1(n5492), .A2(n5491), .ZN(n9356) );
  NAND2_X1 U7054 ( .A1(n5099), .A2(n9356), .ZN(n5494) );
  NAND2_X1 U7055 ( .A1(n4358), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n5493) );
  OAI22_X1 U7056 ( .A1(n9566), .A2(n5148), .B1(n9375), .B2(n5173), .ZN(n5497)
         );
  XNOR2_X1 U7057 ( .A(n5497), .B(n5675), .ZN(n5501) );
  OR2_X1 U7058 ( .A1(n9566), .A2(n5173), .ZN(n5499) );
  OR2_X1 U7059 ( .A1(n9375), .A2(n8031), .ZN(n5498) );
  NAND2_X1 U7060 ( .A1(n5499), .A2(n5498), .ZN(n9081) );
  AOI22_X1 U7061 ( .A1(n8983), .A2(n8982), .B1(n5501), .B2(n9081), .ZN(n5500)
         );
  NAND2_X1 U7062 ( .A1(n8980), .A2(n5500), .ZN(n5509) );
  INV_X1 U7063 ( .A(n8983), .ZN(n5507) );
  INV_X1 U7064 ( .A(n5501), .ZN(n8981) );
  INV_X1 U7065 ( .A(n9081), .ZN(n5502) );
  NAND2_X1 U7066 ( .A1(n8981), .A2(n5502), .ZN(n5503) );
  NAND2_X1 U7067 ( .A1(n5503), .A2(n8982), .ZN(n5506) );
  INV_X1 U7068 ( .A(n5503), .ZN(n5505) );
  INV_X1 U7069 ( .A(n8982), .ZN(n5504) );
  AOI22_X1 U7070 ( .A1(n5507), .A2(n5506), .B1(n5505), .B2(n5504), .ZN(n5508)
         );
  INV_X1 U7071 ( .A(n5510), .ZN(n5513) );
  INV_X1 U7072 ( .A(n5511), .ZN(n5512) );
  NAND2_X1 U7073 ( .A1(n5513), .A2(n5512), .ZN(n5517) );
  INV_X1 U7074 ( .A(n5514), .ZN(n5515) );
  NAND2_X1 U7075 ( .A1(n5515), .A2(n10095), .ZN(n5516) );
  MUX2_X1 U7076 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(P2_DATAO_REG_20__SCAN_IN), 
        .S(n6491), .Z(n5535) );
  XNOR2_X1 U7077 ( .A(n5535), .B(n5536), .ZN(n5518) );
  XNOR2_X1 U7078 ( .A(n5537), .B(n5518), .ZN(n7404) );
  NAND2_X1 U7079 ( .A1(n7404), .A2(n7830), .ZN(n5520) );
  INV_X1 U7080 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7405) );
  OR2_X1 U7081 ( .A1(n5145), .A2(n7405), .ZN(n5519) );
  NAND2_X1 U7082 ( .A1(n9336), .A2(n8036), .ZN(n5528) );
  AND2_X1 U7083 ( .A1(n5521), .A2(n9054), .ZN(n5522) );
  NOR2_X1 U7084 ( .A1(n5540), .A2(n5522), .ZN(n9331) );
  NAND2_X1 U7085 ( .A1(n9331), .A2(n5099), .ZN(n5526) );
  NAND2_X1 U7086 ( .A1(n4355), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n5525) );
  NAND2_X1 U7087 ( .A1(n5098), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n5524) );
  NAND2_X1 U7088 ( .A1(n4358), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n5523) );
  NAND4_X1 U7089 ( .A1(n5526), .A2(n5525), .A3(n5524), .A4(n5523), .ZN(n9124)
         );
  NAND2_X1 U7090 ( .A1(n9124), .A2(n8030), .ZN(n5527) );
  NAND2_X1 U7091 ( .A1(n5528), .A2(n5527), .ZN(n5529) );
  XNOR2_X1 U7092 ( .A(n5529), .B(n8034), .ZN(n9051) );
  AND2_X1 U7093 ( .A1(n9124), .A2(n5677), .ZN(n5530) );
  AOI21_X1 U7094 ( .B1(n9336), .B2(n8030), .A(n5530), .ZN(n9050) );
  AND2_X1 U7095 ( .A1(n9051), .A2(n9050), .ZN(n5534) );
  INV_X1 U7096 ( .A(n9051), .ZN(n5532) );
  INV_X1 U7097 ( .A(n9050), .ZN(n5531) );
  NAND2_X1 U7098 ( .A1(n5532), .A2(n5531), .ZN(n5533) );
  MUX2_X1 U7099 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n6491), .Z(n5558) );
  XNOR2_X1 U7100 ( .A(n5558), .B(SI_21_), .ZN(n5555) );
  XNOR2_X1 U7101 ( .A(n5557), .B(n5555), .ZN(n7497) );
  NAND2_X1 U7102 ( .A1(n7497), .A2(n7830), .ZN(n5539) );
  INV_X1 U7103 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7498) );
  OR2_X1 U7104 ( .A1(n5145), .A2(n7498), .ZN(n5538) );
  NOR2_X1 U7105 ( .A1(n5540), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n5541) );
  OR2_X1 U7106 ( .A1(n5566), .A2(n5541), .ZN(n9315) );
  INV_X1 U7107 ( .A(n5099), .ZN(n5570) );
  NAND2_X1 U7108 ( .A1(n5098), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n5543) );
  NAND2_X1 U7109 ( .A1(n4356), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n5542) );
  AND2_X1 U7110 ( .A1(n5543), .A2(n5542), .ZN(n5545) );
  NAND2_X1 U7111 ( .A1(n4357), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5544) );
  OAI211_X1 U7112 ( .C1(n9315), .C2(n5570), .A(n5545), .B(n5544), .ZN(n9123)
         );
  INV_X1 U7113 ( .A(n9123), .ZN(n5806) );
  OAI22_X1 U7114 ( .A1(n9318), .A2(n5148), .B1(n5806), .B2(n5173), .ZN(n5546)
         );
  XNOR2_X1 U7115 ( .A(n5546), .B(n5675), .ZN(n5549) );
  OR2_X1 U7116 ( .A1(n9318), .A2(n5173), .ZN(n5548) );
  NAND2_X1 U7117 ( .A1(n9123), .A2(n5677), .ZN(n5547) );
  NAND2_X1 U7118 ( .A1(n5548), .A2(n5547), .ZN(n5550) );
  XNOR2_X1 U7119 ( .A(n5549), .B(n5550), .ZN(n8993) );
  INV_X1 U7120 ( .A(n5549), .ZN(n5552) );
  INV_X1 U7121 ( .A(n5550), .ZN(n5551) );
  NAND2_X1 U7122 ( .A1(n5552), .A2(n5551), .ZN(n5553) );
  INV_X1 U7123 ( .A(n5555), .ZN(n5556) );
  NAND2_X1 U7124 ( .A1(n5557), .A2(n5556), .ZN(n5560) );
  NAND2_X1 U7125 ( .A1(n5558), .A2(SI_21_), .ZN(n5559) );
  NAND2_X1 U7126 ( .A1(n5560), .A2(n5559), .ZN(n5576) );
  MUX2_X1 U7127 ( .A(n7517), .B(n7516), .S(n6491), .Z(n5561) );
  NAND2_X1 U7128 ( .A1(n5561), .A2(n10061), .ZN(n5574) );
  INV_X1 U7129 ( .A(n5561), .ZN(n5562) );
  NAND2_X1 U7130 ( .A1(n5562), .A2(SI_22_), .ZN(n5563) );
  NAND2_X1 U7131 ( .A1(n5574), .A2(n5563), .ZN(n5575) );
  XNOR2_X1 U7132 ( .A(n5576), .B(n5575), .ZN(n7515) );
  NAND2_X1 U7133 ( .A1(n7515), .A2(n7830), .ZN(n5565) );
  OR2_X1 U7134 ( .A1(n5145), .A2(n7516), .ZN(n5564) );
  AND2_X2 U7135 ( .A1(n5565), .A2(n5564), .ZN(n9556) );
  OR2_X1 U7136 ( .A1(n5566), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n5567) );
  NAND2_X1 U7137 ( .A1(n5567), .A2(n5583), .ZN(n9304) );
  AOI22_X1 U7138 ( .A1(n5098), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n5097), .B2(
        P1_REG1_REG_22__SCAN_IN), .ZN(n5569) );
  NAND2_X1 U7139 ( .A1(n4357), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5568) );
  OAI211_X1 U7140 ( .C1(n9304), .C2(n5570), .A(n5569), .B(n5568), .ZN(n9122)
         );
  INV_X1 U7141 ( .A(n9122), .ZN(n8995) );
  OAI22_X1 U7142 ( .A1(n9556), .A2(n5148), .B1(n8995), .B2(n5173), .ZN(n5571)
         );
  OR2_X1 U7143 ( .A1(n9556), .A2(n5173), .ZN(n5573) );
  NAND2_X1 U7144 ( .A1(n9122), .A2(n5677), .ZN(n5572) );
  AND2_X1 U7145 ( .A1(n5573), .A2(n5572), .ZN(n9070) );
  NAND2_X1 U7146 ( .A1(n5554), .A2(n4444), .ZN(n9073) );
  OAI21_X2 U7147 ( .B1(n5576), .B2(n5575), .A(n5574), .ZN(n5599) );
  MUX2_X1 U7148 ( .A(n7577), .B(n7573), .S(n6491), .Z(n5577) );
  NAND2_X1 U7149 ( .A1(n5577), .A2(n10106), .ZN(n5600) );
  INV_X1 U7150 ( .A(n5577), .ZN(n5578) );
  NAND2_X1 U7151 ( .A1(n5578), .A2(SI_23_), .ZN(n5579) );
  XNOR2_X1 U7152 ( .A(n5599), .B(n5598), .ZN(n7574) );
  NAND2_X1 U7153 ( .A1(n7574), .A2(n7830), .ZN(n5581) );
  OR2_X1 U7154 ( .A1(n5145), .A2(n7573), .ZN(n5580) );
  NAND2_X1 U7155 ( .A1(n9294), .A2(n8036), .ZN(n5589) );
  NAND2_X1 U7156 ( .A1(n5098), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n5587) );
  NAND2_X1 U7157 ( .A1(n4356), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n5586) );
  INV_X1 U7158 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n8976) );
  INV_X1 U7159 ( .A(n5583), .ZN(n5582) );
  NAND2_X1 U7160 ( .A1(n5582), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5608) );
  AOI21_X1 U7161 ( .B1(n8976), .B2(n5583), .A(n5607), .ZN(n9289) );
  NAND2_X1 U7162 ( .A1(n5099), .A2(n9289), .ZN(n5585) );
  NAND2_X1 U7163 ( .A1(n4358), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5584) );
  NAND4_X1 U7164 ( .A1(n5587), .A2(n5586), .A3(n5585), .A4(n5584), .ZN(n9121)
         );
  NAND2_X1 U7165 ( .A1(n9121), .A2(n5217), .ZN(n5588) );
  NAND2_X1 U7166 ( .A1(n5589), .A2(n5588), .ZN(n5590) );
  XNOR2_X1 U7167 ( .A(n5590), .B(n8034), .ZN(n5592) );
  AND2_X1 U7168 ( .A1(n9121), .A2(n5677), .ZN(n5591) );
  AOI21_X1 U7169 ( .B1(n9294), .B2(n8030), .A(n5591), .ZN(n5593) );
  NAND2_X1 U7170 ( .A1(n5592), .A2(n5593), .ZN(n5597) );
  INV_X1 U7171 ( .A(n5592), .ZN(n5595) );
  INV_X1 U7172 ( .A(n5593), .ZN(n5594) );
  NAND2_X1 U7173 ( .A1(n5595), .A2(n5594), .ZN(n5596) );
  NAND2_X1 U7174 ( .A1(n5597), .A2(n5596), .ZN(n8972) );
  INV_X1 U7175 ( .A(n5597), .ZN(n9041) );
  NAND2_X1 U7176 ( .A1(n5599), .A2(n5598), .ZN(n5601) );
  INV_X1 U7177 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n8137) );
  INV_X1 U7178 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7643) );
  MUX2_X1 U7179 ( .A(n8137), .B(n7643), .S(n6491), .Z(n5602) );
  INV_X1 U7180 ( .A(SI_24_), .ZN(n10074) );
  NAND2_X1 U7181 ( .A1(n5602), .A2(n10074), .ZN(n5620) );
  INV_X1 U7182 ( .A(n5602), .ZN(n5603) );
  NAND2_X1 U7183 ( .A1(n5603), .A2(SI_24_), .ZN(n5604) );
  XNOR2_X1 U7184 ( .A(n5619), .B(n5618), .ZN(n7642) );
  NAND2_X1 U7185 ( .A1(n7642), .A2(n7830), .ZN(n5606) );
  OR2_X1 U7186 ( .A1(n5145), .A2(n7643), .ZN(n5605) );
  NAND2_X1 U7187 ( .A1(n5098), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5612) );
  NAND2_X1 U7188 ( .A1(n4355), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n5611) );
  INV_X1 U7189 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9046) );
  NAND2_X1 U7190 ( .A1(n5607), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n5627) );
  AOI21_X1 U7191 ( .B1(n9046), .B2(n5608), .A(n5626), .ZN(n9278) );
  NAND2_X1 U7192 ( .A1(n5099), .A2(n9278), .ZN(n5610) );
  NAND2_X1 U7193 ( .A1(n4358), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5609) );
  OAI22_X1 U7194 ( .A1(n9548), .A2(n5148), .B1(n9002), .B2(n5173), .ZN(n5613)
         );
  XNOR2_X1 U7195 ( .A(n5613), .B(n5675), .ZN(n5615) );
  OAI22_X1 U7196 ( .A1(n9548), .A2(n5173), .B1(n9002), .B2(n8031), .ZN(n5614)
         );
  OR2_X1 U7197 ( .A1(n5615), .A2(n5614), .ZN(n5617) );
  NAND2_X1 U7198 ( .A1(n5615), .A2(n5614), .ZN(n5616) );
  AND2_X1 U7199 ( .A1(n5617), .A2(n5616), .ZN(n9040) );
  INV_X1 U7200 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n8052) );
  INV_X1 U7201 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7685) );
  MUX2_X1 U7202 ( .A(n8052), .B(n7685), .S(n6491), .Z(n5621) );
  NAND2_X1 U7203 ( .A1(n5621), .A2(n10009), .ZN(n5635) );
  INV_X1 U7204 ( .A(n5621), .ZN(n5622) );
  NAND2_X1 U7205 ( .A1(n5622), .A2(SI_25_), .ZN(n5623) );
  XNOR2_X1 U7206 ( .A(n5634), .B(n5633), .ZN(n7684) );
  NAND2_X1 U7207 ( .A1(n7684), .A2(n7830), .ZN(n5625) );
  OR2_X1 U7208 ( .A1(n5145), .A2(n7685), .ZN(n5624) );
  NAND2_X1 U7209 ( .A1(n5098), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5631) );
  NAND2_X1 U7210 ( .A1(n5097), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n5630) );
  INV_X1 U7211 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n9005) );
  NAND2_X1 U7212 ( .A1(n5626), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n5642) );
  INV_X1 U7213 ( .A(n5642), .ZN(n5643) );
  AOI21_X1 U7214 ( .B1(n9005), .B2(n5627), .A(n5643), .ZN(n9261) );
  NAND2_X1 U7215 ( .A1(n5099), .A2(n9261), .ZN(n5629) );
  NAND2_X1 U7216 ( .A1(n4357), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5628) );
  OAI22_X1 U7217 ( .A1(n9544), .A2(n5148), .B1(n9093), .B2(n5173), .ZN(n5632)
         );
  XNOR2_X1 U7218 ( .A(n5632), .B(n5675), .ZN(n5654) );
  OAI22_X1 U7219 ( .A1(n9544), .A2(n5173), .B1(n9093), .B2(n8031), .ZN(n5653)
         );
  XNOR2_X1 U7220 ( .A(n5654), .B(n5653), .ZN(n9000) );
  INV_X1 U7221 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7690) );
  INV_X1 U7222 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7688) );
  MUX2_X1 U7223 ( .A(n7690), .B(n7688), .S(n6491), .Z(n5637) );
  NAND2_X1 U7224 ( .A1(n5637), .A2(n10071), .ZN(n5661) );
  INV_X1 U7225 ( .A(n5637), .ZN(n5638) );
  NAND2_X1 U7226 ( .A1(n5638), .A2(SI_26_), .ZN(n5639) );
  NAND2_X1 U7227 ( .A1(n7687), .A2(n7830), .ZN(n5641) );
  OR2_X1 U7228 ( .A1(n5145), .A2(n7688), .ZN(n5640) );
  NAND2_X1 U7229 ( .A1(n5098), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n5648) );
  NAND2_X1 U7230 ( .A1(n4356), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n5647) );
  INV_X1 U7231 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9094) );
  NAND2_X1 U7232 ( .A1(n9094), .A2(n5642), .ZN(n5644) );
  NAND2_X1 U7233 ( .A1(P1_REG3_REG_26__SCAN_IN), .A2(n5643), .ZN(n5669) );
  NAND2_X1 U7234 ( .A1(n5099), .A2(n9243), .ZN(n5646) );
  NAND2_X1 U7235 ( .A1(n4358), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5645) );
  NAND4_X1 U7236 ( .A1(n5648), .A2(n5647), .A3(n5646), .A4(n5645), .ZN(n9118)
         );
  AND2_X1 U7237 ( .A1(n9118), .A2(n5677), .ZN(n5649) );
  AOI21_X1 U7238 ( .B1(n9249), .B2(n8030), .A(n5649), .ZN(n5656) );
  NAND2_X1 U7239 ( .A1(n9249), .A2(n8036), .ZN(n5651) );
  NAND2_X1 U7240 ( .A1(n9118), .A2(n5217), .ZN(n5650) );
  NAND2_X1 U7241 ( .A1(n5651), .A2(n5650), .ZN(n5652) );
  XNOR2_X1 U7242 ( .A(n5652), .B(n5675), .ZN(n5658) );
  XOR2_X1 U7243 ( .A(n5656), .B(n5658), .Z(n9088) );
  NOR2_X1 U7244 ( .A1(n5654), .A2(n5653), .ZN(n9089) );
  INV_X1 U7245 ( .A(n5656), .ZN(n5657) );
  NAND2_X1 U7246 ( .A1(n5660), .A2(n5659), .ZN(n5662) );
  NAND2_X1 U7247 ( .A1(n5662), .A2(n5661), .ZN(n5771) );
  INV_X1 U7248 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n8958) );
  INV_X1 U7249 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n7694) );
  MUX2_X1 U7250 ( .A(n8958), .B(n7694), .S(n6491), .Z(n5663) );
  INV_X1 U7251 ( .A(SI_27_), .ZN(n9959) );
  NAND2_X1 U7252 ( .A1(n5663), .A2(n9959), .ZN(n5772) );
  INV_X1 U7253 ( .A(n5663), .ZN(n5664) );
  NAND2_X1 U7254 ( .A1(n5664), .A2(SI_27_), .ZN(n5665) );
  NAND2_X1 U7255 ( .A1(n7693), .A2(n7830), .ZN(n5667) );
  OR2_X1 U7256 ( .A1(n5145), .A2(n7694), .ZN(n5666) );
  NAND2_X1 U7257 ( .A1(n5098), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n5674) );
  NAND2_X1 U7258 ( .A1(n4355), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n5673) );
  INV_X1 U7259 ( .A(n5669), .ZN(n5668) );
  NAND2_X1 U7260 ( .A1(n5668), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n5813) );
  INV_X1 U7261 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n5730) );
  NAND2_X1 U7262 ( .A1(n5669), .A2(n5730), .ZN(n5670) );
  NAND2_X1 U7263 ( .A1(n5099), .A2(n9232), .ZN(n5672) );
  NAND2_X1 U7264 ( .A1(n4357), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5671) );
  AOI22_X1 U7265 ( .A1(n9231), .A2(n8036), .B1(n8030), .B2(n9117), .ZN(n5676)
         );
  XNOR2_X1 U7266 ( .A(n5676), .B(n5675), .ZN(n5679) );
  AOI22_X1 U7267 ( .A1(n9231), .A2(n5217), .B1(n5677), .B2(n9117), .ZN(n5678)
         );
  NAND2_X1 U7268 ( .A1(n5679), .A2(n5678), .ZN(n8044) );
  OAI21_X1 U7269 ( .B1(n5679), .B2(n5678), .A(n8044), .ZN(n5682) );
  NOR3_X2 U7270 ( .A1(n5680), .A2(n5681), .A3(n5682), .ZN(n8051) );
  INV_X1 U7271 ( .A(n5680), .ZN(n9092) );
  INV_X1 U7272 ( .A(n5681), .ZN(n5684) );
  INV_X1 U7273 ( .A(n5682), .ZN(n5683) );
  AOI21_X1 U7274 ( .B1(n9092), .B2(n5684), .A(n5683), .ZN(n5715) );
  INV_X1 U7275 ( .A(P1_B_REG_SCAN_IN), .ZN(n5685) );
  NAND2_X1 U7276 ( .A1(n5686), .A2(n5685), .ZN(n5688) );
  NAND3_X1 U7277 ( .A1(n7686), .A2(P1_B_REG_SCAN_IN), .A3(n7644), .ZN(n5687)
         );
  INV_X1 U7278 ( .A(n9577), .ZN(n5703) );
  NOR4_X1 U7279 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n5698) );
  NOR4_X1 U7280 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n5697) );
  OR4_X1 U7281 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n5695) );
  NOR4_X1 U7282 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n5693) );
  NOR4_X1 U7283 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n5692) );
  NOR4_X1 U7284 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5691) );
  NOR4_X1 U7285 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n5690) );
  NAND4_X1 U7286 ( .A1(n5693), .A2(n5692), .A3(n5691), .A4(n5690), .ZN(n5694)
         );
  NOR4_X1 U7287 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n5695), .A4(n5694), .ZN(n5696) );
  NAND3_X1 U7288 ( .A1(n5698), .A2(n5697), .A3(n5696), .ZN(n5699) );
  NAND2_X1 U7289 ( .A1(n5703), .A2(n5699), .ZN(n5826) );
  INV_X1 U7290 ( .A(n5826), .ZN(n5701) );
  INV_X1 U7291 ( .A(n5700), .ZN(n7689) );
  NAND2_X1 U7292 ( .A1(n7689), .A2(n7686), .ZN(n9579) );
  OAI21_X1 U7293 ( .B1(n9577), .B2(P1_D_REG_1__SCAN_IN), .A(n9579), .ZN(n5827)
         );
  NOR2_X1 U7294 ( .A1(n5701), .A2(n5827), .ZN(n7005) );
  INV_X1 U7295 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n5702) );
  NAND2_X1 U7296 ( .A1(n5703), .A2(n5702), .ZN(n5704) );
  NAND2_X1 U7297 ( .A1(n7689), .A2(n7644), .ZN(n9580) );
  INV_X1 U7298 ( .A(n6464), .ZN(n5705) );
  NAND2_X1 U7299 ( .A1(n7005), .A2(n5705), .ZN(n5718) );
  NAND2_X1 U7300 ( .A1(n5707), .A2(n5706), .ZN(n5708) );
  NAND2_X1 U7301 ( .A1(n5708), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5710) );
  INV_X1 U7302 ( .A(n7924), .ZN(n7931) );
  AND2_X1 U7303 ( .A1(n7841), .A2(n7931), .ZN(n5822) );
  OR2_X1 U7304 ( .A1(n9724), .A2(n6508), .ZN(n5713) );
  NOR2_X1 U7305 ( .A1(n6506), .A2(n5713), .ZN(n5714) );
  OAI21_X1 U7306 ( .B1(n8051), .B2(n5715), .A(n9102), .ZN(n5735) );
  NAND2_X1 U7307 ( .A1(n5822), .A2(n7982), .ZN(n7012) );
  INV_X1 U7308 ( .A(n7012), .ZN(n5716) );
  NAND3_X1 U7309 ( .A1(n5729), .A2(n9578), .A3(n5716), .ZN(n5717) );
  NAND2_X1 U7310 ( .A1(n5718), .A2(n5825), .ZN(n6624) );
  AND2_X1 U7311 ( .A1(n5711), .A2(n6508), .ZN(n5824) );
  INV_X1 U7312 ( .A(n6507), .ZN(n5719) );
  NOR2_X1 U7313 ( .A1(n5824), .A2(n5719), .ZN(n5720) );
  AND2_X1 U7314 ( .A1(n6463), .A2(n5720), .ZN(n5721) );
  NAND2_X1 U7315 ( .A1(n6624), .A2(n5721), .ZN(n9030) );
  NAND2_X1 U7316 ( .A1(n5097), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n5725) );
  NAND2_X1 U7317 ( .A1(n4358), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5724) );
  XNOR2_X1 U7318 ( .A(n5813), .B(P1_REG3_REG_28__SCAN_IN), .ZN(n8081) );
  NAND2_X1 U7319 ( .A1(n5099), .A2(n8081), .ZN(n5723) );
  NAND2_X1 U7320 ( .A1(n5098), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n5722) );
  OR2_X1 U7321 ( .A1(n8054), .A2(n9414), .ZN(n5728) );
  INV_X1 U7322 ( .A(n5726), .ZN(n9157) );
  NAND2_X1 U7323 ( .A1(n9118), .A2(n9393), .ZN(n5727) );
  AND2_X1 U7324 ( .A1(n5728), .A2(n5727), .ZN(n9228) );
  NOR2_X1 U7325 ( .A1(n6506), .A2(n5711), .ZN(n7983) );
  NAND2_X1 U7326 ( .A1(n5729), .A2(n7983), .ZN(n9095) );
  OAI22_X1 U7327 ( .A1(n9228), .A2(n9095), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n5730), .ZN(n5731) );
  AOI21_X1 U7328 ( .B1(n9232), .B2(n9109), .A(n5731), .ZN(n5732) );
  INV_X1 U7329 ( .A(n5733), .ZN(n5734) );
  NAND2_X1 U7330 ( .A1(n5735), .A2(n5734), .ZN(P1_U3214) );
  INV_X1 U7331 ( .A(n9107), .ZN(n9128) );
  XNOR2_X1 U7332 ( .A(n5737), .B(n5821), .ZN(n5783) );
  NAND2_X1 U7333 ( .A1(n5736), .A2(n7013), .ZN(n7069) );
  NAND2_X1 U7334 ( .A1(n5783), .A2(n7069), .ZN(n7068) );
  NAND2_X1 U7335 ( .A1(n7068), .A2(n4947), .ZN(n6667) );
  NAND2_X1 U7336 ( .A1(n7065), .A2(n7142), .ZN(n5786) );
  NAND2_X1 U7337 ( .A1(n7936), .A2(n5786), .ZN(n6665) );
  NAND2_X1 U7338 ( .A1(n6667), .A2(n6665), .ZN(n6666) );
  NAND2_X1 U7339 ( .A1(n6666), .A2(n5739), .ZN(n7093) );
  NAND2_X1 U7340 ( .A1(n9139), .A2(n5740), .ZN(n7941) );
  NAND2_X1 U7341 ( .A1(n7093), .A2(n7092), .ZN(n7091) );
  NAND2_X1 U7342 ( .A1(n5741), .A2(n5740), .ZN(n5742) );
  NAND2_X1 U7343 ( .A1(n7091), .A2(n5742), .ZN(n6960) );
  NAND2_X1 U7344 ( .A1(n7090), .A2(n7079), .ZN(n7714) );
  NAND2_X1 U7345 ( .A1(n9138), .A2(n6971), .ZN(n7940) );
  NAND2_X1 U7346 ( .A1(n7714), .A2(n7940), .ZN(n7847) );
  NAND2_X1 U7347 ( .A1(n6960), .A2(n7847), .ZN(n6961) );
  NAND2_X1 U7348 ( .A1(n7090), .A2(n6971), .ZN(n5743) );
  NAND2_X1 U7349 ( .A1(n6961), .A2(n5743), .ZN(n6860) );
  NAND2_X1 U7350 ( .A1(n7728), .A2(n7727), .ZN(n7713) );
  NAND2_X1 U7351 ( .A1(n9137), .A2(n5744), .ZN(n7944) );
  NAND2_X1 U7352 ( .A1(n7713), .A2(n7944), .ZN(n6859) );
  NAND2_X1 U7353 ( .A1(n6860), .A2(n6859), .ZN(n6858) );
  NAND2_X1 U7354 ( .A1(n7728), .A2(n5744), .ZN(n5745) );
  NAND2_X1 U7355 ( .A1(n6858), .A2(n5745), .ZN(n7173) );
  NAND2_X1 U7356 ( .A1(n7722), .A2(n4576), .ZN(n5746) );
  OAI21_X1 U7357 ( .B1(n7722), .B2(n4576), .A(n5746), .ZN(n7716) );
  INV_X1 U7358 ( .A(n7716), .ZN(n7178) );
  XNOR2_X1 U7359 ( .A(n9135), .B(n9739), .ZN(n7108) );
  NAND2_X1 U7360 ( .A1(n7385), .A2(n7292), .ZN(n7740) );
  INV_X1 U7361 ( .A(n7385), .ZN(n9134) );
  NAND2_X1 U7362 ( .A1(n9134), .A2(n7309), .ZN(n7150) );
  NAND2_X1 U7363 ( .A1(n7740), .A2(n7150), .ZN(n7216) );
  NAND2_X1 U7364 ( .A1(n7209), .A2(n7216), .ZN(n7208) );
  NAND2_X1 U7365 ( .A1(n7208), .A2(n5748), .ZN(n7160) );
  INV_X1 U7366 ( .A(n7324), .ZN(n9133) );
  NAND2_X1 U7367 ( .A1(n9133), .A2(n7390), .ZN(n7750) );
  NAND2_X1 U7368 ( .A1(n7324), .A2(n7157), .ZN(n7745) );
  NAND2_X1 U7369 ( .A1(n7750), .A2(n7745), .ZN(n7159) );
  NAND2_X1 U7370 ( .A1(n7160), .A2(n7159), .ZN(n7158) );
  NAND2_X1 U7371 ( .A1(n7158), .A2(n5749), .ZN(n7331) );
  OR2_X1 U7372 ( .A1(n7431), .A2(n9629), .ZN(n7949) );
  NAND2_X1 U7373 ( .A1(n9629), .A2(n7431), .ZN(n7746) );
  NAND2_X1 U7374 ( .A1(n7949), .A2(n7746), .ZN(n7330) );
  NAND2_X1 U7375 ( .A1(n7331), .A2(n7330), .ZN(n7329) );
  INV_X1 U7376 ( .A(n7431), .ZN(n9132) );
  NAND2_X1 U7377 ( .A1(n7329), .A2(n5751), .ZN(n7428) );
  OR2_X1 U7378 ( .A1(n7446), .A2(n7460), .ZN(n7752) );
  NAND2_X1 U7379 ( .A1(n7446), .A2(n7460), .ZN(n7753) );
  NAND2_X1 U7380 ( .A1(n7752), .A2(n7753), .ZN(n7858) );
  NAND2_X1 U7381 ( .A1(n7428), .A2(n7858), .ZN(n7427) );
  NAND2_X1 U7382 ( .A1(n7427), .A2(n5752), .ZN(n7456) );
  OR2_X1 U7383 ( .A1(n7628), .A2(n7531), .ZN(n7756) );
  NAND2_X1 U7384 ( .A1(n7628), .A2(n7531), .ZN(n7955) );
  NAND2_X1 U7385 ( .A1(n7756), .A2(n7955), .ZN(n7859) );
  NAND2_X1 U7386 ( .A1(n7456), .A2(n7859), .ZN(n7455) );
  INV_X1 U7387 ( .A(n7531), .ZN(n9130) );
  NAND2_X1 U7388 ( .A1(n5753), .A2(n7531), .ZN(n5754) );
  NAND2_X1 U7389 ( .A1(n7455), .A2(n5754), .ZN(n7529) );
  OR2_X1 U7390 ( .A1(n9066), .A2(n9413), .ZN(n7760) );
  NAND2_X1 U7391 ( .A1(n9066), .A2(n9413), .ZN(n7956) );
  NAND2_X1 U7392 ( .A1(n7760), .A2(n7956), .ZN(n7845) );
  NAND2_X1 U7393 ( .A1(n7529), .A2(n7845), .ZN(n7530) );
  INV_X1 U7394 ( .A(n9413), .ZN(n9129) );
  NAND2_X1 U7395 ( .A1(n7530), .A2(n5755), .ZN(n9407) );
  OR2_X1 U7396 ( .A1(n9425), .A2(n9107), .ZN(n7761) );
  NAND2_X1 U7397 ( .A1(n9425), .A2(n9107), .ZN(n7767) );
  NAND2_X1 U7398 ( .A1(n7761), .A2(n7767), .ZN(n9409) );
  NOR2_X1 U7399 ( .A1(n9514), .A2(n9392), .ZN(n5756) );
  INV_X1 U7400 ( .A(n9514), .ZN(n9114) );
  OR2_X1 U7401 ( .A1(n9399), .A2(n9373), .ZN(n7770) );
  NAND2_X1 U7402 ( .A1(n9399), .A2(n9373), .ZN(n9370) );
  NAND2_X1 U7403 ( .A1(n7770), .A2(n9370), .ZN(n9385) );
  INV_X1 U7404 ( .A(n9373), .ZN(n9127) );
  NAND2_X1 U7405 ( .A1(n9504), .A2(n9391), .ZN(n5757) );
  INV_X1 U7406 ( .A(n9391), .ZN(n5799) );
  NAND2_X1 U7407 ( .A1(n9566), .A2(n9375), .ZN(n5758) );
  INV_X1 U7408 ( .A(n9375), .ZN(n9126) );
  NAND2_X1 U7409 ( .A1(n9491), .A2(n9125), .ZN(n5759) );
  INV_X1 U7410 ( .A(n9125), .ZN(n5804) );
  NAND2_X1 U7411 ( .A1(n9330), .A2(n5760), .ZN(n5761) );
  NAND2_X1 U7412 ( .A1(n5761), .A2(n4945), .ZN(n9311) );
  NAND2_X1 U7413 ( .A1(n9556), .A2(n8995), .ZN(n5763) );
  NOR2_X1 U7414 ( .A1(n9556), .A2(n8995), .ZN(n5762) );
  NAND2_X1 U7415 ( .A1(n9294), .A2(n9121), .ZN(n5764) );
  NAND2_X1 U7416 ( .A1(n9548), .A2(n9002), .ZN(n5765) );
  NAND2_X1 U7417 ( .A1(n9267), .A2(n5765), .ZN(n5767) );
  INV_X1 U7418 ( .A(n9002), .ZN(n9120) );
  NAND2_X1 U7419 ( .A1(n9277), .A2(n9120), .ZN(n5766) );
  NOR2_X1 U7420 ( .A1(n9544), .A2(n9093), .ZN(n5769) );
  NAND2_X1 U7421 ( .A1(n9544), .A2(n9093), .ZN(n5768) );
  INV_X1 U7422 ( .A(n9118), .ZN(n7798) );
  NAND2_X1 U7423 ( .A1(n5771), .A2(n5770), .ZN(n5773) );
  INV_X1 U7424 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8957) );
  INV_X1 U7425 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n7705) );
  MUX2_X1 U7426 ( .A(n8957), .B(n7705), .S(n6491), .Z(n5774) );
  NAND2_X1 U7427 ( .A1(n5774), .A2(n10062), .ZN(n6363) );
  INV_X1 U7428 ( .A(n5774), .ZN(n5775) );
  NAND2_X1 U7429 ( .A1(n5775), .A2(SI_28_), .ZN(n5776) );
  NAND2_X1 U7430 ( .A1(n6351), .A2(n7830), .ZN(n5778) );
  OR2_X1 U7431 ( .A1(n5145), .A2(n7705), .ZN(n5777) );
  INV_X1 U7432 ( .A(n7872), .ZN(n5779) );
  NAND2_X1 U7433 ( .A1(n4388), .A2(n5779), .ZN(n8057) );
  OAI21_X1 U7434 ( .B1(n4388), .B2(n5779), .A(n8057), .ZN(n8092) );
  INV_X1 U7435 ( .A(n6508), .ZN(n7912) );
  OR2_X1 U7436 ( .A1(n5711), .A2(n7912), .ZN(n5780) );
  INV_X1 U7437 ( .A(n5822), .ZN(n6633) );
  NAND2_X1 U7438 ( .A1(n5780), .A2(n6633), .ZN(n7008) );
  AND2_X1 U7439 ( .A1(n5711), .A2(n5781), .ZN(n5782) );
  OR2_X1 U7440 ( .A1(n7008), .A2(n5782), .ZN(n9741) );
  BUF_X1 U7441 ( .A(n5783), .Z(n7852) );
  INV_X1 U7442 ( .A(n7852), .ZN(n5784) );
  NOR2_X1 U7443 ( .A1(n5736), .A2(n7071), .ZN(n7060) );
  INV_X1 U7444 ( .A(n5737), .ZN(n6670) );
  NAND2_X1 U7445 ( .A1(n6670), .A2(n7072), .ZN(n5785) );
  INV_X1 U7446 ( .A(n5786), .ZN(n5787) );
  INV_X1 U7447 ( .A(n7092), .ZN(n7849) );
  INV_X1 U7448 ( .A(n7847), .ZN(n7711) );
  NAND2_X1 U7449 ( .A1(n6963), .A2(n7714), .ZN(n6857) );
  INV_X1 U7450 ( .A(n6859), .ZN(n7848) );
  NAND2_X1 U7451 ( .A1(n6857), .A2(n7848), .ZN(n5788) );
  NAND2_X1 U7452 ( .A1(n5788), .A2(n7713), .ZN(n7177) );
  NAND2_X1 U7453 ( .A1(n5747), .A2(n7116), .ZN(n7214) );
  NAND2_X1 U7454 ( .A1(n7740), .A2(n7214), .ZN(n7734) );
  AND2_X1 U7455 ( .A1(n7750), .A2(n7150), .ZN(n7742) );
  NAND2_X1 U7456 ( .A1(n7734), .A2(n7742), .ZN(n5789) );
  NAND2_X1 U7457 ( .A1(n5789), .A2(n7745), .ZN(n5791) );
  NAND2_X1 U7458 ( .A1(n7722), .A2(n7723), .ZN(n7721) );
  INV_X1 U7459 ( .A(n7721), .ZN(n7107) );
  OR2_X1 U7460 ( .A1(n7177), .A2(n7950), .ZN(n7321) );
  NAND2_X1 U7461 ( .A1(n9135), .A2(n9739), .ZN(n5790) );
  AND2_X1 U7462 ( .A1(n7150), .A2(n5790), .ZN(n7736) );
  INV_X1 U7463 ( .A(n7722), .ZN(n9136) );
  NAND2_X1 U7464 ( .A1(n9136), .A2(n4576), .ZN(n7729) );
  AND3_X1 U7465 ( .A1(n7736), .A2(n7750), .A3(n7729), .ZN(n7854) );
  OR2_X1 U7466 ( .A1(n7854), .A2(n5791), .ZN(n7948) );
  INV_X1 U7467 ( .A(n7330), .ZN(n7855) );
  AND2_X1 U7468 ( .A1(n7948), .A2(n7855), .ZN(n5792) );
  INV_X1 U7469 ( .A(n7746), .ZN(n7749) );
  NOR2_X1 U7470 ( .A1(n7858), .A2(n7749), .ZN(n5793) );
  NAND2_X1 U7471 ( .A1(n7430), .A2(n5793), .ZN(n7457) );
  INV_X1 U7472 ( .A(n7752), .ZN(n5794) );
  NOR2_X1 U7473 ( .A1(n7859), .A2(n5794), .ZN(n5795) );
  NAND2_X1 U7474 ( .A1(n7457), .A2(n5795), .ZN(n5796) );
  NAND2_X1 U7475 ( .A1(n5796), .A2(n7955), .ZN(n7528) );
  OR2_X1 U7476 ( .A1(n9514), .A2(n9415), .ZN(n7762) );
  NAND2_X1 U7477 ( .A1(n9514), .A2(n9415), .ZN(n7766) );
  NAND2_X1 U7478 ( .A1(n7762), .A2(n7766), .ZN(n7863) );
  INV_X1 U7479 ( .A(n7767), .ZN(n7960) );
  NOR2_X1 U7480 ( .A1(n7863), .A2(n7960), .ZN(n5798) );
  OR2_X1 U7481 ( .A1(n9504), .A2(n5799), .ZN(n7777) );
  NAND2_X1 U7482 ( .A1(n9504), .A2(n5799), .ZN(n7780) );
  NAND2_X1 U7483 ( .A1(n7777), .A2(n7780), .ZN(n9371) );
  INV_X1 U7484 ( .A(n9370), .ZN(n5800) );
  NOR2_X1 U7485 ( .A1(n9371), .A2(n5800), .ZN(n5801) );
  NAND2_X1 U7486 ( .A1(n9388), .A2(n5801), .ZN(n5802) );
  NAND2_X1 U7487 ( .A1(n5802), .A2(n7777), .ZN(n9352) );
  NAND2_X1 U7488 ( .A1(n9363), .A2(n9375), .ZN(n7781) );
  NAND2_X1 U7489 ( .A1(n9352), .A2(n9353), .ZN(n5803) );
  OR2_X1 U7490 ( .A1(n9491), .A2(n5804), .ZN(n7966) );
  NAND2_X1 U7491 ( .A1(n9491), .A2(n5804), .ZN(n7970) );
  NAND2_X1 U7492 ( .A1(n7966), .A2(n7970), .ZN(n9341) );
  XNOR2_X1 U7493 ( .A(n9336), .B(n9343), .ZN(n9329) );
  OR2_X1 U7494 ( .A1(n9336), .A2(n9343), .ZN(n7785) );
  XNOR2_X1 U7495 ( .A(n9476), .B(n9123), .ZN(n9320) );
  NAND2_X1 U7496 ( .A1(n9476), .A2(n5806), .ZN(n7787) );
  XNOR2_X1 U7497 ( .A(n9303), .B(n9122), .ZN(n9298) );
  NAND2_X1 U7498 ( .A1(n9303), .A2(n8995), .ZN(n7792) );
  INV_X1 U7499 ( .A(n9121), .ZN(n7795) );
  OR2_X1 U7500 ( .A1(n9294), .A2(n7795), .ZN(n7790) );
  NAND2_X1 U7501 ( .A1(n9294), .A2(n7795), .ZN(n9270) );
  NAND2_X1 U7502 ( .A1(n9277), .A2(n9002), .ZN(n7889) );
  INV_X1 U7503 ( .A(n9270), .ZN(n7793) );
  NOR2_X1 U7504 ( .A1(n7868), .A2(n7793), .ZN(n5807) );
  NAND2_X1 U7505 ( .A1(n9284), .A2(n5807), .ZN(n9268) );
  OR2_X1 U7506 ( .A1(n9260), .A2(n9093), .ZN(n7881) );
  NAND2_X1 U7507 ( .A1(n9260), .A2(n9093), .ZN(n7890) );
  NAND2_X1 U7508 ( .A1(n7881), .A2(n7890), .ZN(n9254) );
  INV_X1 U7509 ( .A(n9253), .ZN(n5808) );
  NOR2_X1 U7510 ( .A1(n9254), .A2(n5808), .ZN(n5809) );
  NAND2_X1 U7511 ( .A1(n9268), .A2(n5809), .ZN(n5810) );
  NAND2_X1 U7512 ( .A1(n5810), .A2(n7890), .ZN(n9239) );
  XNOR2_X1 U7513 ( .A(n9249), .B(n9118), .ZN(n9242) );
  NAND2_X1 U7514 ( .A1(n9249), .A2(n7798), .ZN(n7897) );
  XNOR2_X1 U7515 ( .A(n8061), .B(n7872), .ZN(n8089) );
  NAND2_X1 U7516 ( .A1(n7875), .A2(n5712), .ZN(n5812) );
  NAND2_X1 U7517 ( .A1(n7924), .A2(n7982), .ZN(n5811) );
  NAND2_X1 U7518 ( .A1(n5098), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n5817) );
  NAND2_X1 U7519 ( .A1(n4356), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n5816) );
  INV_X1 U7520 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n8043) );
  NOR2_X1 U7521 ( .A1(n5813), .A2(n8043), .ZN(n9215) );
  NAND2_X1 U7522 ( .A1(n5099), .A2(n9215), .ZN(n5815) );
  NAND2_X1 U7523 ( .A1(n4357), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n5814) );
  OR2_X1 U7524 ( .A1(n7812), .A2(n9414), .ZN(n5820) );
  OR2_X1 U7525 ( .A1(n5818), .A2(n9412), .ZN(n5819) );
  NAND2_X1 U7526 ( .A1(n5820), .A2(n5819), .ZN(n8082) );
  NAND2_X1 U7527 ( .A1(n5821), .A2(n7071), .ZN(n7070) );
  OR2_X1 U7528 ( .A1(n7070), .A2(n7142), .ZN(n7094) );
  AND2_X1 U7529 ( .A1(n7180), .A2(n9739), .ZN(n7210) );
  INV_X1 U7530 ( .A(n7446), .ZN(n7608) );
  NAND2_X1 U7531 ( .A1(n7464), .A2(n5753), .ZN(n7535) );
  NAND2_X1 U7532 ( .A1(n9274), .A2(n9548), .ZN(n9275) );
  INV_X1 U7533 ( .A(n9230), .ZN(n5823) );
  NAND2_X1 U7534 ( .A1(n9230), .A2(n8085), .ZN(n8068) );
  INV_X1 U7535 ( .A(n8068), .ZN(n8069) );
  AOI211_X1 U7536 ( .C1(n8055), .C2(n5823), .A(n9422), .B(n8069), .ZN(n8087)
         );
  NAND2_X1 U7537 ( .A1(n5830), .A2(n5829), .ZN(n5887) );
  NOR2_X1 U7538 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n5833) );
  NOR2_X1 U7539 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n5836) );
  NAND4_X1 U7540 ( .A1(n5836), .A2(n5879), .A3(n5951), .A4(n5835), .ZN(n5839)
         );
  NAND4_X1 U7541 ( .A1(n5875), .A2(n5873), .A3(n5946), .A4(n5837), .ZN(n5838)
         );
  NOR2_X1 U7542 ( .A1(n5839), .A2(n5838), .ZN(n5840) );
  NAND2_X1 U7543 ( .A1(n5863), .A2(n5851), .ZN(n5853) );
  NAND2_X1 U7544 ( .A1(n5861), .A2(n5862), .ZN(n5843) );
  NAND2_X1 U7545 ( .A1(n5847), .A2(n5846), .ZN(n5849) );
  INV_X1 U7546 ( .A(n6424), .ZN(n5860) );
  NAND2_X1 U7547 ( .A1(n5849), .A2(n5848), .ZN(n6422) );
  INV_X1 U7548 ( .A(n5853), .ZN(n5855) );
  NAND3_X1 U7549 ( .A1(n5855), .A2(n5854), .A3(n5862), .ZN(n5856) );
  NAND2_X1 U7550 ( .A1(n5856), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5857) );
  NOR2_X1 U7551 ( .A1(n6422), .A2(n7692), .ZN(n5859) );
  INV_X1 U7552 ( .A(n6737), .ZN(n7575) );
  OR2_X1 U7553 ( .A1(n6738), .A2(n7575), .ZN(n6043) );
  INV_X1 U7554 ( .A(n5863), .ZN(n5868) );
  NAND2_X1 U7555 ( .A1(n5868), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5864) );
  NAND2_X1 U7556 ( .A1(n5866), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5867) );
  MUX2_X1 U7557 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5867), .S(
        P2_IR_REG_21__SCAN_IN), .Z(n5869) );
  NAND2_X1 U7558 ( .A1(n6737), .A2(n8454), .ZN(n5870) );
  NAND2_X1 U7559 ( .A1(n6043), .A2(n5870), .ZN(n6042) );
  OAI21_X1 U7560 ( .B1(n6042), .B2(n6257), .A(P2_STATE_REG_SCAN_IN), .ZN(
        P2_U3150) );
  NAND2_X1 U7561 ( .A1(n4430), .A2(n5873), .ZN(n5933) );
  NAND3_X1 U7562 ( .A1(n5879), .A2(n5938), .A3(n5875), .ZN(n5876) );
  OR2_X1 U7563 ( .A1(n4451), .A2(n6058), .ZN(n5877) );
  XNOR2_X1 U7564 ( .A(n5877), .B(P2_IR_REG_16__SCAN_IN), .ZN(n8599) );
  NAND2_X1 U7565 ( .A1(n5878), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5882) );
  NAND2_X1 U7566 ( .A1(n5882), .A2(n5879), .ZN(n5880) );
  NAND2_X1 U7567 ( .A1(n5880), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5939) );
  NAND2_X1 U7568 ( .A1(n5939), .A2(n5938), .ZN(n5941) );
  NAND2_X1 U7569 ( .A1(n5941), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5881) );
  XNOR2_X1 U7570 ( .A(n5881), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8583) );
  XNOR2_X1 U7571 ( .A(n5882), .B(P2_IR_REG_13__SCAN_IN), .ZN(n8549) );
  OR2_X1 U7572 ( .A1(n4430), .A2(n6058), .ZN(n5883) );
  OR2_X1 U7573 ( .A1(n5884), .A2(n6058), .ZN(n5886) );
  XNOR2_X1 U7574 ( .A(n5886), .B(n5885), .ZN(n6612) );
  NAND2_X1 U7575 ( .A1(n5920), .A2(n5921), .ZN(n5893) );
  OAI21_X1 U7576 ( .B1(n5890), .B2(P2_IR_REG_8__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5889) );
  XNOR2_X1 U7577 ( .A(n5889), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7343) );
  NAND2_X1 U7578 ( .A1(n5890), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5892) );
  NAND2_X1 U7579 ( .A1(n5893), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5894) );
  INV_X1 U7580 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6080) );
  NOR2_X1 U7581 ( .A1(n6080), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n5898) );
  INV_X1 U7582 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6480) );
  NAND2_X2 U7583 ( .A1(n5904), .A2(n5903), .ZN(n5966) );
  NAND2_X1 U7584 ( .A1(n5901), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5908) );
  MUX2_X1 U7585 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5908), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n5909) );
  AND2_X1 U7586 ( .A1(n5909), .A2(n5888), .ZN(n9773) );
  NAND2_X1 U7587 ( .A1(n5888), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5912) );
  XNOR2_X1 U7588 ( .A(n5912), .B(P2_IR_REG_4__SCAN_IN), .ZN(n6001) );
  INV_X1 U7589 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n5913) );
  AOI22_X1 U7590 ( .A1(P2_REG2_REG_4__SCAN_IN), .A2(n6001), .B1(n6694), .B2(
        n5913), .ZN(n6696) );
  NOR2_X1 U7591 ( .A1(n6697), .A2(n6696), .ZN(n6695) );
  NAND2_X1 U7592 ( .A1(n5916), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5917) );
  XNOR2_X1 U7593 ( .A(n5917), .B(P2_IR_REG_5__SCAN_IN), .ZN(n6013) );
  INV_X1 U7594 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n9786) );
  OR2_X1 U7595 ( .A1(n5920), .A2(n6058), .ZN(n5922) );
  NAND2_X1 U7596 ( .A1(P2_REG2_REG_6__SCAN_IN), .A2(n6764), .ZN(n5923) );
  OAI21_X1 U7597 ( .B1(P2_REG2_REG_6__SCAN_IN), .B2(n6764), .A(n5923), .ZN(
        n6757) );
  NOR2_X1 U7598 ( .A1(n6139), .A2(n5925), .ZN(n5926) );
  INV_X1 U7599 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n9826) );
  NAND2_X1 U7600 ( .A1(P2_REG2_REG_8__SCAN_IN), .A2(n7048), .ZN(n5927) );
  OAI21_X1 U7601 ( .B1(P2_REG2_REG_8__SCAN_IN), .B2(n7048), .A(n5927), .ZN(
        n7050) );
  NOR2_X1 U7602 ( .A1(n7343), .A2(n5928), .ZN(n5929) );
  INV_X1 U7603 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7352) );
  INV_X1 U7604 ( .A(n7343), .ZN(n6592) );
  NAND2_X1 U7605 ( .A1(P2_REG2_REG_10__SCAN_IN), .A2(n6612), .ZN(n5930) );
  OAI21_X1 U7606 ( .B1(P2_REG2_REG_10__SCAN_IN), .B2(n6612), .A(n5930), .ZN(
        n7407) );
  NOR2_X1 U7607 ( .A1(n7408), .A2(n7407), .ZN(n7406) );
  INV_X1 U7608 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7474) );
  NAND2_X1 U7609 ( .A1(n5933), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5934) );
  XNOR2_X1 U7610 ( .A(n5934), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7653) );
  INV_X1 U7611 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n5935) );
  AOI22_X1 U7612 ( .A1(P2_REG2_REG_12__SCAN_IN), .A2(n7653), .B1(n6688), .B2(
        n5935), .ZN(n7657) );
  NOR2_X1 U7613 ( .A1(n8549), .A2(n5936), .ZN(n5937) );
  INV_X1 U7614 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n8544) );
  XNOR2_X1 U7615 ( .A(n5936), .B(n8549), .ZN(n8543) );
  NOR2_X1 U7616 ( .A1(n5937), .A2(n8542), .ZN(n8561) );
  OR2_X1 U7617 ( .A1(n5939), .A2(n5938), .ZN(n5940) );
  INV_X1 U7618 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n5942) );
  AOI22_X1 U7619 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n8566), .B1(n6777), .B2(
        n5942), .ZN(n8560) );
  NOR2_X1 U7620 ( .A1(n8559), .A2(n4950), .ZN(n5943) );
  NOR2_X1 U7621 ( .A1(n8583), .A2(n5943), .ZN(n5944) );
  INV_X1 U7622 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8578) );
  INV_X1 U7623 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n5945) );
  AOI22_X1 U7624 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n8599), .B1(n7019), .B2(
        n5945), .ZN(n8603) );
  NAND2_X1 U7625 ( .A1(n5950), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5947) );
  XNOR2_X1 U7626 ( .A(n5947), .B(P2_IR_REG_17__SCAN_IN), .ZN(n6239) );
  XNOR2_X1 U7627 ( .A(n5948), .B(n6239), .ZN(n9798) );
  INV_X1 U7628 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n9799) );
  NOR2_X1 U7629 ( .A1(n9798), .A2(n9799), .ZN(n9797) );
  NOR2_X1 U7630 ( .A1(n6239), .A2(n5948), .ZN(n5949) );
  NAND2_X1 U7631 ( .A1(n5952), .A2(n5951), .ZN(n5953) );
  XNOR2_X1 U7632 ( .A(n5957), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8627) );
  INV_X1 U7633 ( .A(n8627), .ZN(n7138) );
  NAND2_X1 U7634 ( .A1(n7138), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n5954) );
  OAI21_X1 U7635 ( .B1(n7138), .B2(P2_REG2_REG_18__SCAN_IN), .A(n5954), .ZN(
        n8614) );
  INV_X1 U7636 ( .A(n5954), .ZN(n5955) );
  INV_X1 U7637 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n5958) );
  INV_X1 U7638 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5956) );
  MUX2_X1 U7639 ( .A(n5958), .B(P2_REG2_REG_19__SCAN_IN), .S(n6421), .Z(n5994)
         );
  XNOR2_X1 U7640 ( .A(n5959), .B(n5994), .ZN(n6052) );
  OR2_X1 U7641 ( .A1(n5960), .A2(P2_U3151), .ZN(n8954) );
  NOR2_X1 U7642 ( .A1(n6042), .A2(n8954), .ZN(n9760) );
  INV_X1 U7643 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n9876) );
  INV_X1 U7644 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n6081) );
  NOR2_X1 U7645 ( .A1(n6081), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n5961) );
  INV_X1 U7646 ( .A(n6476), .ZN(n5962) );
  INV_X1 U7647 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6845) );
  NAND2_X1 U7648 ( .A1(n5966), .A2(n5965), .ZN(n5964) );
  INV_X1 U7649 ( .A(n5971), .ZN(n5970) );
  AOI22_X1 U7650 ( .A1(P2_REG1_REG_4__SCAN_IN), .A2(n6001), .B1(n6694), .B2(
        n5972), .ZN(n6699) );
  NOR2_X1 U7651 ( .A1(n6700), .A2(n6699), .ZN(n6698) );
  INV_X1 U7652 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n9879) );
  NOR2_X1 U7653 ( .A1(n6013), .A2(n5974), .ZN(n5975) );
  NAND2_X1 U7654 ( .A1(P2_REG1_REG_6__SCAN_IN), .A2(n6764), .ZN(n5976) );
  OAI21_X1 U7655 ( .B1(P2_REG1_REG_6__SCAN_IN), .B2(n6764), .A(n5976), .ZN(
        n6759) );
  NOR2_X1 U7656 ( .A1(n6139), .A2(n5978), .ZN(n5979) );
  XNOR2_X1 U7657 ( .A(n5978), .B(n6139), .ZN(n6947) );
  NAND2_X1 U7658 ( .A1(P2_REG1_REG_8__SCAN_IN), .A2(n7048), .ZN(n5980) );
  OAI21_X1 U7659 ( .B1(P2_REG1_REG_8__SCAN_IN), .B2(n7048), .A(n5980), .ZN(
        n7042) );
  NOR2_X1 U7660 ( .A1(n7343), .A2(n5981), .ZN(n5982) );
  INV_X1 U7661 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n7341) );
  NAND2_X1 U7662 ( .A1(P2_REG1_REG_10__SCAN_IN), .A2(n6612), .ZN(n5983) );
  OAI21_X1 U7663 ( .B1(n6612), .B2(P2_REG1_REG_10__SCAN_IN), .A(n5983), .ZN(
        n7417) );
  NOR2_X1 U7664 ( .A1(n7481), .A2(n5984), .ZN(n5985) );
  INV_X1 U7665 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n9883) );
  INV_X1 U7666 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n6200) );
  MUX2_X1 U7667 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n6200), .S(n7653), .Z(n7646)
         );
  NOR2_X1 U7668 ( .A1(n8549), .A2(n5986), .ZN(n5987) );
  INV_X1 U7669 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n8872) );
  INV_X1 U7670 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8868) );
  AOI22_X1 U7671 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n8566), .B1(n6777), .B2(
        n8868), .ZN(n8558) );
  INV_X1 U7672 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8864) );
  XNOR2_X1 U7673 ( .A(n7019), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n8592) );
  INV_X1 U7674 ( .A(n6239), .ZN(n9813) );
  INV_X1 U7675 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n9802) );
  NAND2_X1 U7676 ( .A1(n7138), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n5991) );
  OAI21_X1 U7677 ( .B1(n7138), .B2(P2_REG1_REG_18__SCAN_IN), .A(n5991), .ZN(
        n8611) );
  XNOR2_X1 U7678 ( .A(n6421), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n5995) );
  MUX2_X1 U7679 ( .A(n5995), .B(n5994), .S(n8514), .Z(n6038) );
  MUX2_X1 U7680 ( .A(n9799), .B(n9802), .S(n6004), .Z(n6034) );
  XNOR2_X1 U7681 ( .A(n6034), .B(n9813), .ZN(n9805) );
  MUX2_X1 U7682 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n6004), .Z(n5996) );
  AND2_X1 U7683 ( .A1(n5996), .A2(n7019), .ZN(n8594) );
  MUX2_X1 U7684 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n6004), .Z(n6030) );
  INV_X1 U7685 ( .A(n8583), .ZN(n6816) );
  NOR2_X1 U7686 ( .A1(n6030), .A2(n6816), .ZN(n6032) );
  MUX2_X1 U7687 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n6004), .Z(n6027) );
  NOR2_X1 U7688 ( .A1(n6027), .A2(n6777), .ZN(n6029) );
  MUX2_X1 U7689 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n6004), .Z(n6024) );
  NOR2_X1 U7690 ( .A1(n6024), .A2(n6716), .ZN(n6026) );
  MUX2_X1 U7691 ( .A(P2_REG2_REG_12__SCAN_IN), .B(P2_REG1_REG_12__SCAN_IN), 
        .S(n6004), .Z(n6023) );
  NOR2_X1 U7692 ( .A1(n6023), .A2(n6688), .ZN(n7648) );
  MUX2_X1 U7693 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n6004), .Z(n5998) );
  INV_X1 U7694 ( .A(n5998), .ZN(n5997) );
  NAND2_X1 U7695 ( .A1(n5997), .A2(n7481), .ZN(n6022) );
  XNOR2_X1 U7696 ( .A(n5998), .B(n7481), .ZN(n7479) );
  MUX2_X1 U7697 ( .A(P2_REG2_REG_10__SCAN_IN), .B(P2_REG1_REG_10__SCAN_IN), 
        .S(n6004), .Z(n5999) );
  OR2_X1 U7698 ( .A1(n5999), .A2(n6612), .ZN(n6021) );
  INV_X1 U7699 ( .A(n6612), .ZN(n7409) );
  XNOR2_X1 U7700 ( .A(n5999), .B(n7409), .ZN(n7412) );
  MUX2_X1 U7701 ( .A(P2_REG2_REG_9__SCAN_IN), .B(P2_REG1_REG_9__SCAN_IN), .S(
        n6004), .Z(n6000) );
  OR2_X1 U7702 ( .A1(n6000), .A2(n6592), .ZN(n6020) );
  XNOR2_X1 U7703 ( .A(n6000), .B(n7343), .ZN(n7346) );
  MUX2_X1 U7704 ( .A(P2_REG2_REG_8__SCAN_IN), .B(P2_REG1_REG_8__SCAN_IN), .S(
        n6004), .Z(n6018) );
  OR2_X1 U7705 ( .A1(n6018), .A2(n7048), .ZN(n6019) );
  INV_X1 U7706 ( .A(n6764), .ZN(n6151) );
  MUX2_X1 U7707 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n6004), .Z(n6014) );
  INV_X1 U7708 ( .A(n6014), .ZN(n6015) );
  MUX2_X1 U7709 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n6004), .Z(n6011) );
  INV_X1 U7710 ( .A(n6011), .ZN(n6012) );
  MUX2_X1 U7711 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n6004), .Z(n6009) );
  XNOR2_X1 U7712 ( .A(n6009), .B(n6001), .ZN(n6692) );
  INV_X1 U7713 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6104) );
  MUX2_X1 U7714 ( .A(n6104), .B(n9876), .S(n6004), .Z(n6008) );
  INV_X1 U7715 ( .A(n9773), .ZN(n6493) );
  XNOR2_X1 U7716 ( .A(n6008), .B(n6493), .ZN(n9775) );
  MUX2_X1 U7717 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n6004), .Z(n6006) );
  MUX2_X1 U7718 ( .A(P2_REG2_REG_1__SCAN_IN), .B(P2_REG1_REG_1__SCAN_IN), .S(
        n6004), .Z(n6005) );
  MUX2_X1 U7719 ( .A(P2_REG2_REG_0__SCAN_IN), .B(P2_REG1_REG_0__SCAN_IN), .S(
        n6004), .Z(n9758) );
  NOR2_X1 U7720 ( .A1(n9758), .A2(n9763), .ZN(n6472) );
  XNOR2_X1 U7721 ( .A(n6006), .B(n5966), .ZN(n6661) );
  AOI21_X1 U7722 ( .B1(n6006), .B2(n5966), .A(n6659), .ZN(n9776) );
  NAND2_X1 U7723 ( .A1(n9775), .A2(n9776), .ZN(n9774) );
  INV_X1 U7724 ( .A(n9774), .ZN(n6007) );
  NAND2_X1 U7725 ( .A1(n6009), .A2(n6694), .ZN(n6010) );
  XNOR2_X1 U7726 ( .A(n6011), .B(n6013), .ZN(n9781) );
  OAI21_X1 U7727 ( .B1(n6013), .B2(n6012), .A(n9780), .ZN(n6754) );
  XNOR2_X1 U7728 ( .A(n6014), .B(n6764), .ZN(n6755) );
  NOR2_X1 U7729 ( .A1(n6754), .A2(n6755), .ZN(n6753) );
  AOI21_X1 U7730 ( .B1(n6151), .B2(n6015), .A(n6753), .ZN(n6949) );
  INV_X1 U7731 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6133) );
  MUX2_X1 U7732 ( .A(n9826), .B(n6133), .S(n6004), .Z(n6016) );
  XNOR2_X1 U7733 ( .A(n6016), .B(n6139), .ZN(n6948) );
  INV_X1 U7734 ( .A(n6016), .ZN(n6017) );
  INV_X1 U7735 ( .A(n6139), .ZN(n6951) );
  OAI22_X1 U7736 ( .A1(n6949), .A2(n6948), .B1(n6017), .B2(n6951), .ZN(n7046)
         );
  INV_X1 U7737 ( .A(n7048), .ZN(n6155) );
  XNOR2_X1 U7738 ( .A(n6018), .B(n6155), .ZN(n7045) );
  NAND2_X1 U7739 ( .A1(n7046), .A2(n7045), .ZN(n7044) );
  NAND2_X1 U7740 ( .A1(n6019), .A2(n7044), .ZN(n7345) );
  NAND2_X1 U7741 ( .A1(n7346), .A2(n7345), .ZN(n7344) );
  NAND2_X1 U7742 ( .A1(n6020), .A2(n7344), .ZN(n7411) );
  NAND2_X1 U7743 ( .A1(n7412), .A2(n7411), .ZN(n7410) );
  NAND2_X1 U7744 ( .A1(n6021), .A2(n7410), .ZN(n7478) );
  AND2_X1 U7745 ( .A1(n6023), .A2(n6688), .ZN(n7649) );
  AOI21_X1 U7746 ( .B1(n6024), .B2(n6716), .A(n6026), .ZN(n6025) );
  INV_X1 U7747 ( .A(n6025), .ZN(n8547) );
  NOR2_X1 U7748 ( .A1(n6026), .A2(n8546), .ZN(n8564) );
  AOI21_X1 U7749 ( .B1(n6027), .B2(n6777), .A(n6029), .ZN(n6028) );
  INV_X1 U7750 ( .A(n6028), .ZN(n8565) );
  NOR2_X1 U7751 ( .A1(n8564), .A2(n8565), .ZN(n8563) );
  NOR2_X1 U7752 ( .A1(n6029), .A2(n8563), .ZN(n8581) );
  AOI21_X1 U7753 ( .B1(n6030), .B2(n6816), .A(n6032), .ZN(n6031) );
  INV_X1 U7754 ( .A(n6031), .ZN(n8582) );
  NOR2_X1 U7755 ( .A1(n8581), .A2(n8582), .ZN(n8580) );
  NOR2_X1 U7756 ( .A1(n6032), .A2(n8580), .ZN(n8598) );
  INV_X1 U7757 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n6233) );
  MUX2_X1 U7758 ( .A(n5945), .B(n6233), .S(n6004), .Z(n6033) );
  NAND2_X1 U7759 ( .A1(n6033), .A2(n8599), .ZN(n8596) );
  MUX2_X1 U7760 ( .A(P2_REG2_REG_18__SCAN_IN), .B(P2_REG1_REG_18__SCAN_IN), 
        .S(n6004), .Z(n6035) );
  NOR2_X1 U7761 ( .A1(n6036), .A2(n6035), .ZN(n8620) );
  NAND2_X1 U7762 ( .A1(n6036), .A2(n6035), .ZN(n8618) );
  OAI21_X1 U7763 ( .B1(n8620), .B2(n8627), .A(n8618), .ZN(n6037) );
  XOR2_X1 U7764 ( .A(n6038), .B(n6037), .Z(n6050) );
  INV_X1 U7765 ( .A(n6619), .ZN(n6039) );
  INV_X1 U7766 ( .A(n5960), .ZN(n6407) );
  NOR2_X2 U7767 ( .A1(n8621), .A2(n6407), .ZN(n9807) );
  NOR2_X1 U7768 ( .A1(n6004), .A2(P2_U3151), .ZN(n6040) );
  NAND2_X1 U7769 ( .A1(n6040), .A2(n5960), .ZN(n6041) );
  OR2_X1 U7770 ( .A1(n6042), .A2(n6041), .ZN(n6046) );
  INV_X1 U7771 ( .A(n6043), .ZN(n6047) );
  INV_X1 U7772 ( .A(n8954), .ZN(n6044) );
  NAND2_X1 U7773 ( .A1(n6047), .A2(n6044), .ZN(n6045) );
  NAND2_X1 U7774 ( .A1(n6046), .A2(n6045), .ZN(n9772) );
  NAND2_X1 U7775 ( .A1(n9796), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n6048) );
  NAND2_X1 U7776 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8167) );
  OAI211_X1 U7777 ( .C1(n9814), .C2(n6405), .A(n6048), .B(n8167), .ZN(n6049)
         );
  NAND2_X1 U7778 ( .A1(n6778), .A2(n8288), .ZN(n6055) );
  AOI22_X1 U7779 ( .A1(n6258), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n6257), .B2(
        n8583), .ZN(n6054) );
  NAND2_X1 U7780 ( .A1(n6059), .A2(n6060), .ZN(n8946) );
  XNOR2_X2 U7781 ( .A(n6061), .B(n6060), .ZN(n6065) );
  AND2_X4 U7782 ( .A1(n6062), .A2(n6065), .ZN(n6090) );
  NAND2_X1 U7783 ( .A1(n6090), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n6070) );
  OR2_X1 U7784 ( .A1(n4359), .A2(n8864), .ZN(n6069) );
  NOR2_X1 U7785 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n6122) );
  NAND2_X1 U7786 ( .A1(n6122), .A2(n6123), .ZN(n6143) );
  NAND2_X1 U7787 ( .A1(n6209), .A2(n6208), .ZN(n6218) );
  AND2_X1 U7788 ( .A1(n6220), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6064) );
  NOR2_X1 U7789 ( .A1(n6230), .A2(n6064), .ZN(n7582) );
  OR2_X1 U7790 ( .A1(n6211), .A2(n7582), .ZN(n6068) );
  NAND2_X4 U7791 ( .A1(n6066), .A2(n6065), .ZN(n6411) );
  OR2_X1 U7792 ( .A1(n6411), .A2(n8578), .ZN(n6067) );
  INV_X1 U7793 ( .A(n8791), .ZN(n8527) );
  INV_X1 U7794 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n6470) );
  OR2_X1 U7795 ( .A1(n6211), .A2(n6470), .ZN(n6072) );
  NAND2_X1 U7796 ( .A1(n6090), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n6071) );
  AND2_X1 U7797 ( .A1(n6072), .A2(n6071), .ZN(n6075) );
  OR2_X1 U7798 ( .A1(n4360), .A2(n6845), .ZN(n6074) );
  NAND3_X2 U7799 ( .A1(n6075), .A2(n6074), .A3(n6073), .ZN(n6788) );
  INV_X1 U7800 ( .A(n6788), .ZN(n6752) );
  INV_X1 U7801 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6497) );
  OR2_X1 U7802 ( .A1(n6076), .A2(n6499), .ZN(n6077) );
  NAND2_X1 U7803 ( .A1(n6788), .A2(n6079), .ZN(n8320) );
  OR2_X1 U7804 ( .A1(n6411), .A2(n6080), .ZN(n6085) );
  NAND2_X1 U7805 ( .A1(n6090), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n6084) );
  INV_X1 U7806 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n10111) );
  OR2_X1 U7807 ( .A1(n6211), .A2(n10111), .ZN(n6082) );
  NAND2_X1 U7808 ( .A1(n7825), .A2(SI_0_), .ZN(n6087) );
  INV_X1 U7809 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n6086) );
  NAND2_X1 U7810 ( .A1(n6087), .A2(n6086), .ZN(n6089) );
  AND2_X1 U7811 ( .A1(n6089), .A2(n6088), .ZN(n8962) );
  NAND2_X1 U7812 ( .A1(n6382), .A2(n7003), .ZN(n6834) );
  OR2_X1 U7813 ( .A1(n6788), .A2(n4461), .ZN(n6875) );
  NAND2_X1 U7814 ( .A1(n6876), .A2(n6875), .ZN(n6101) );
  NAND2_X1 U7815 ( .A1(n6090), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n6096) );
  OR2_X1 U7816 ( .A1(n4359), .A2(n5965), .ZN(n6095) );
  INV_X1 U7817 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n6092) );
  OR2_X1 U7818 ( .A1(n6211), .A2(n6092), .ZN(n6094) );
  OR2_X1 U7819 ( .A1(n6076), .A2(n5966), .ZN(n6100) );
  OR2_X1 U7820 ( .A1(n8291), .A2(n5061), .ZN(n6099) );
  OR2_X1 U7821 ( .A1(n6369), .A2(n6494), .ZN(n6098) );
  NAND2_X1 U7822 ( .A1(n6102), .A2(n9827), .ZN(n8326) );
  OR2_X1 U7823 ( .A1(n6102), .A2(n4860), .ZN(n6103) );
  NAND2_X1 U7824 ( .A1(n6090), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n6108) );
  OR2_X1 U7825 ( .A1(n4360), .A2(n9876), .ZN(n6107) );
  OR2_X1 U7826 ( .A1(n6211), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n6106) );
  OR2_X1 U7827 ( .A1(n6411), .A2(n6104), .ZN(n6105) );
  OR2_X1 U7828 ( .A1(n6097), .A2(n6492), .ZN(n6110) );
  OR2_X1 U7829 ( .A1(n8291), .A2(n5084), .ZN(n6109) );
  OAI211_X1 U7830 ( .C1(n6076), .C2(n6493), .A(n6110), .B(n6109), .ZN(n9834)
         );
  NAND2_X1 U7831 ( .A1(n8539), .A2(n9834), .ZN(n6111) );
  OR2_X1 U7832 ( .A1(n8539), .A2(n9834), .ZN(n6112) );
  NAND2_X1 U7833 ( .A1(n6090), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n6117) );
  AND2_X1 U7834 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n6113) );
  NOR2_X1 U7835 ( .A1(n6122), .A2(n6113), .ZN(n6941) );
  OR2_X1 U7836 ( .A1(n6411), .A2(n5913), .ZN(n6114) );
  OR2_X1 U7837 ( .A1(n6369), .A2(n6496), .ZN(n6119) );
  OR2_X1 U7838 ( .A1(n8291), .A2(n5117), .ZN(n6118) );
  OAI211_X1 U7839 ( .C1(n6076), .C2(n6694), .A(n6119), .B(n6118), .ZN(n6943)
         );
  NOR2_X1 U7840 ( .A1(n8538), .A2(n6943), .ZN(n6121) );
  NAND2_X1 U7841 ( .A1(n8538), .A2(n6943), .ZN(n6120) );
  NAND2_X1 U7842 ( .A1(n6090), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n6128) );
  OR2_X1 U7843 ( .A1(n4360), .A2(n9879), .ZN(n6127) );
  OR2_X1 U7844 ( .A1(n6123), .A2(n6122), .ZN(n6124) );
  AND2_X1 U7845 ( .A1(n6143), .A2(n6124), .ZN(n7036) );
  OR2_X1 U7846 ( .A1(n6211), .A2(n7036), .ZN(n6126) );
  OR2_X1 U7847 ( .A1(n6411), .A2(n9786), .ZN(n6125) );
  NAND4_X1 U7848 ( .A1(n6128), .A2(n6127), .A3(n6126), .A4(n6125), .ZN(n8537)
         );
  OR2_X1 U7849 ( .A1(n6369), .A2(n6501), .ZN(n6130) );
  INV_X1 U7850 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6500) );
  OR2_X1 U7851 ( .A1(n8291), .A2(n6500), .ZN(n6129) );
  OAI211_X1 U7852 ( .C1(n6076), .C2(n9795), .A(n6130), .B(n6129), .ZN(n9845)
         );
  AND2_X1 U7853 ( .A1(n8537), .A2(n9845), .ZN(n6132) );
  OR2_X1 U7854 ( .A1(n8537), .A2(n9845), .ZN(n6131) );
  NAND2_X1 U7855 ( .A1(n6090), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n6138) );
  OR2_X1 U7856 ( .A1(n4360), .A2(n6133), .ZN(n6137) );
  AND2_X1 U7857 ( .A1(n6145), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6134) );
  NOR2_X1 U7858 ( .A1(n6159), .A2(n6134), .ZN(n7393) );
  OR2_X1 U7859 ( .A1(n6211), .A2(n7393), .ZN(n6136) );
  OR2_X1 U7860 ( .A1(n6411), .A2(n9826), .ZN(n6135) );
  INV_X1 U7861 ( .A(n8535), .ZN(n7241) );
  OR2_X1 U7862 ( .A1(n6513), .A2(n6369), .ZN(n6141) );
  AOI22_X1 U7863 ( .A1(n6258), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6257), .B2(
        n6139), .ZN(n6140) );
  AND2_X1 U7864 ( .A1(n7241), .A2(n8350), .ZN(n6177) );
  NAND2_X1 U7865 ( .A1(n6090), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n6150) );
  INV_X1 U7866 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6142) );
  OR2_X1 U7867 ( .A1(n4359), .A2(n6142), .ZN(n6149) );
  NAND2_X1 U7868 ( .A1(n6143), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6144) );
  AND2_X1 U7869 ( .A1(n6145), .A2(n6144), .ZN(n8251) );
  OR2_X1 U7870 ( .A1(n6211), .A2(n8251), .ZN(n6148) );
  INV_X1 U7871 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6146) );
  OR2_X1 U7872 ( .A1(n6411), .A2(n6146), .ZN(n6147) );
  AOI22_X1 U7873 ( .A1(n6258), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n6257), .B2(
        n6151), .ZN(n6153) );
  OR2_X1 U7874 ( .A1(n6504), .A2(n6369), .ZN(n6152) );
  OR2_X1 U7875 ( .A1(n8536), .A2(n9850), .ZN(n8345) );
  NAND2_X1 U7876 ( .A1(n8536), .A2(n9850), .ZN(n8347) );
  OR2_X1 U7877 ( .A1(n6524), .A2(n6369), .ZN(n6157) );
  AOI22_X1 U7878 ( .A1(n6258), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6257), .B2(
        n6155), .ZN(n6156) );
  NAND2_X2 U7879 ( .A1(n6157), .A2(n6156), .ZN(n9859) );
  NAND2_X1 U7880 ( .A1(n6090), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n6164) );
  INV_X1 U7881 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6158) );
  OR2_X1 U7882 ( .A1(n4360), .A2(n6158), .ZN(n6163) );
  INV_X1 U7883 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7134) );
  OR2_X1 U7884 ( .A1(n6411), .A2(n7134), .ZN(n6162) );
  NOR2_X1 U7885 ( .A1(n6159), .A2(n10098), .ZN(n6160) );
  OR2_X1 U7886 ( .A1(n6169), .A2(n6160), .ZN(n7260) );
  INV_X1 U7887 ( .A(n7260), .ZN(n7133) );
  OR2_X1 U7888 ( .A1(n6211), .A2(n7133), .ZN(n6161) );
  OR2_X2 U7889 ( .A1(n9859), .A2(n7396), .ZN(n8363) );
  INV_X1 U7890 ( .A(n7129), .ZN(n8476) );
  OR2_X1 U7891 ( .A1(n7124), .A2(n8476), .ZN(n7127) );
  INV_X1 U7892 ( .A(n7127), .ZN(n6175) );
  AOI22_X1 U7893 ( .A1(n6258), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6257), .B2(
        n7343), .ZN(n6166) );
  NAND2_X1 U7894 ( .A1(n6090), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n6174) );
  OR2_X1 U7895 ( .A1(n4359), .A2(n7341), .ZN(n6173) );
  OR2_X1 U7896 ( .A1(n6169), .A2(n6168), .ZN(n6170) );
  AND2_X1 U7897 ( .A1(n6182), .A2(n6170), .ZN(n7374) );
  OR2_X1 U7898 ( .A1(n6211), .A2(n7374), .ZN(n6172) );
  OR2_X1 U7899 ( .A1(n6411), .A2(n7352), .ZN(n6171) );
  OR2_X1 U7900 ( .A1(n7369), .A2(n8533), .ZN(n6176) );
  XNOR2_X1 U7901 ( .A(n8350), .B(n8535), .ZN(n7301) );
  INV_X1 U7902 ( .A(n9850), .ZN(n8249) );
  NAND2_X1 U7903 ( .A1(n8536), .A2(n8249), .ZN(n7296) );
  AND2_X1 U7904 ( .A1(n7301), .A2(n7296), .ZN(n7297) );
  NAND2_X1 U7905 ( .A1(n7369), .A2(n7258), .ZN(n8353) );
  INV_X1 U7906 ( .A(n7396), .ZN(n8534) );
  NAND2_X1 U7907 ( .A1(n9859), .A2(n8534), .ZN(n7196) );
  AND2_X1 U7908 ( .A1(n6390), .A2(n7196), .ZN(n6178) );
  NAND2_X1 U7909 ( .A1(n6593), .A2(n8288), .ZN(n6180) );
  AOI22_X1 U7910 ( .A1(n6258), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6257), .B2(
        n7409), .ZN(n6179) );
  NAND2_X1 U7911 ( .A1(n6180), .A2(n6179), .ZN(n7525) );
  NAND2_X1 U7912 ( .A1(n6090), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n6187) );
  INV_X1 U7913 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n6181) );
  OR2_X1 U7914 ( .A1(n4360), .A2(n6181), .ZN(n6186) );
  INV_X1 U7915 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7521) );
  OR2_X1 U7916 ( .A1(n6411), .A2(n7521), .ZN(n6185) );
  NAND2_X1 U7917 ( .A1(n6182), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6183) );
  AND2_X1 U7918 ( .A1(n6190), .A2(n6183), .ZN(n7520) );
  OR2_X1 U7919 ( .A1(n6211), .A2(n7520), .ZN(n6184) );
  OR2_X1 U7920 ( .A1(n7525), .A2(n7993), .ZN(n8357) );
  NAND2_X1 U7921 ( .A1(n7525), .A2(n7993), .ZN(n8354) );
  NAND2_X1 U7922 ( .A1(n8357), .A2(n8354), .ZN(n8479) );
  INV_X1 U7923 ( .A(n7993), .ZN(n8532) );
  NAND2_X1 U7924 ( .A1(n6627), .A2(n8288), .ZN(n6189) );
  AOI22_X1 U7925 ( .A1(n6258), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6257), .B2(
        n7481), .ZN(n6188) );
  NAND2_X1 U7926 ( .A1(n6189), .A2(n6188), .ZN(n7996) );
  NAND2_X1 U7927 ( .A1(n6090), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n6195) );
  OR2_X1 U7928 ( .A1(n4359), .A2(n9883), .ZN(n6194) );
  OR2_X1 U7929 ( .A1(n6411), .A2(n7474), .ZN(n6193) );
  NAND2_X1 U7930 ( .A1(n6190), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6191) );
  AND2_X1 U7931 ( .A1(n6201), .A2(n6191), .ZN(n7994) );
  OR2_X1 U7932 ( .A1(n6211), .A2(n7994), .ZN(n6192) );
  NAND4_X1 U7933 ( .A1(n6195), .A2(n6194), .A3(n6193), .A4(n6192), .ZN(n8531)
         );
  NAND2_X1 U7934 ( .A1(n7990), .A2(n7996), .ZN(n6196) );
  NAND2_X1 U7935 ( .A1(n6197), .A2(n6196), .ZN(n7450) );
  NAND2_X1 U7936 ( .A1(n6673), .A2(n8288), .ZN(n6199) );
  AOI22_X1 U7937 ( .A1(n6258), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6257), .B2(
        n7653), .ZN(n6198) );
  NAND2_X1 U7938 ( .A1(n6199), .A2(n6198), .ZN(n9870) );
  NAND2_X1 U7939 ( .A1(n6090), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n6205) );
  OR2_X1 U7940 ( .A1(n4360), .A2(n6200), .ZN(n6204) );
  NOR2_X1 U7941 ( .A1(n6209), .A2(n4942), .ZN(n7567) );
  OR2_X1 U7942 ( .A1(n6211), .A2(n7567), .ZN(n6203) );
  OR2_X1 U7943 ( .A1(n6411), .A2(n5935), .ZN(n6202) );
  OR2_X1 U7944 ( .A1(n9870), .A2(n7992), .ZN(n8383) );
  NAND2_X1 U7945 ( .A1(n9870), .A2(n7992), .ZN(n8382) );
  NAND2_X1 U7946 ( .A1(n8383), .A2(n8382), .ZN(n8379) );
  NAND2_X1 U7947 ( .A1(n6689), .A2(n8288), .ZN(n6207) );
  AOI22_X1 U7948 ( .A1(n6258), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6257), .B2(
        n8549), .ZN(n6206) );
  NAND2_X1 U7949 ( .A1(n6090), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n6215) );
  OR2_X1 U7950 ( .A1(n4359), .A2(n8872), .ZN(n6214) );
  OR2_X1 U7951 ( .A1(n6209), .A2(n6208), .ZN(n6210) );
  AND2_X1 U7952 ( .A1(n6210), .A2(n6218), .ZN(n7679) );
  OR2_X1 U7953 ( .A1(n6211), .A2(n7679), .ZN(n6213) );
  OR2_X1 U7954 ( .A1(n6411), .A2(n8544), .ZN(n6212) );
  NAND4_X1 U7955 ( .A1(n6215), .A2(n6214), .A3(n6213), .A4(n6212), .ZN(n8529)
         );
  NOR2_X1 U7956 ( .A1(n8388), .A2(n8529), .ZN(n8392) );
  NAND2_X1 U7957 ( .A1(n8388), .A2(n8529), .ZN(n8386) );
  OAI21_X2 U7958 ( .B1(n7542), .B2(n8392), .A(n8386), .ZN(n7587) );
  NAND2_X1 U7959 ( .A1(n6773), .A2(n8288), .ZN(n6217) );
  AOI22_X1 U7960 ( .A1(n6258), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6257), .B2(
        n8566), .ZN(n6216) );
  NAND2_X1 U7961 ( .A1(n6090), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n6224) );
  OR2_X1 U7962 ( .A1(n4360), .A2(n8868), .ZN(n6223) );
  NAND2_X1 U7963 ( .A1(n6218), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6219) );
  AND2_X1 U7964 ( .A1(n6220), .A2(n6219), .ZN(n8151) );
  OR2_X1 U7965 ( .A1(n6211), .A2(n8151), .ZN(n6222) );
  OR2_X1 U7966 ( .A1(n6411), .A2(n5942), .ZN(n6221) );
  NAND2_X1 U7967 ( .A1(n8938), .A2(n8096), .ZN(n6226) );
  OR2_X1 U7968 ( .A1(n8098), .A2(n8791), .ZN(n8399) );
  NAND2_X1 U7969 ( .A1(n8098), .A2(n8791), .ZN(n8398) );
  NAND2_X1 U7970 ( .A1(n8399), .A2(n8398), .ZN(n8394) );
  NAND2_X1 U7971 ( .A1(n7017), .A2(n8288), .ZN(n6228) );
  AOI22_X1 U7972 ( .A1(n6258), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6257), .B2(
        n8599), .ZN(n6227) );
  INV_X1 U7973 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n6229) );
  NOR2_X1 U7974 ( .A1(n6230), .A2(n6229), .ZN(n6231) );
  OR2_X1 U7975 ( .A1(n6242), .A2(n6231), .ZN(n8796) );
  NAND2_X1 U7976 ( .A1(n6308), .A2(n8796), .ZN(n6237) );
  INV_X1 U7977 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n6232) );
  OR2_X1 U7978 ( .A1(n6373), .A2(n6232), .ZN(n6236) );
  OR2_X1 U7979 ( .A1(n4359), .A2(n6233), .ZN(n6235) );
  OR2_X1 U7980 ( .A1(n6411), .A2(n5945), .ZN(n6234) );
  NAND2_X1 U7981 ( .A1(n8857), .A2(n8777), .ZN(n8402) );
  INV_X1 U7982 ( .A(n8777), .ZN(n8526) );
  NAND2_X1 U7983 ( .A1(n7026), .A2(n8288), .ZN(n6241) );
  AOI22_X1 U7984 ( .A1(n6258), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6257), .B2(
        n6239), .ZN(n6240) );
  NAND2_X1 U7985 ( .A1(n6241), .A2(n6240), .ZN(n8202) );
  OR2_X1 U7986 ( .A1(n6242), .A2(n10091), .ZN(n6243) );
  NAND2_X1 U7987 ( .A1(n6250), .A2(n6243), .ZN(n8780) );
  NAND2_X1 U7988 ( .A1(n6308), .A2(n8780), .ZN(n6247) );
  OR2_X1 U7989 ( .A1(n4359), .A2(n9802), .ZN(n6246) );
  OR2_X1 U7990 ( .A1(n6411), .A2(n9799), .ZN(n6245) );
  INV_X1 U7991 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n8927) );
  OR2_X1 U7992 ( .A1(n6373), .A2(n8927), .ZN(n6244) );
  OR2_X1 U7993 ( .A1(n8202), .A2(n8789), .ZN(n8409) );
  NAND2_X1 U7994 ( .A1(n7120), .A2(n8288), .ZN(n6249) );
  AOI22_X1 U7995 ( .A1(n6258), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6257), .B2(
        n8627), .ZN(n6248) );
  NAND2_X1 U7996 ( .A1(n6250), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6251) );
  NAND2_X1 U7997 ( .A1(n6261), .A2(n6251), .ZN(n8769) );
  NAND2_X1 U7998 ( .A1(n8769), .A2(n6308), .ZN(n6256) );
  NAND2_X1 U7999 ( .A1(n6090), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n6255) );
  NAND2_X1 U8000 ( .A1(n6321), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n6254) );
  INV_X1 U8001 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n6252) );
  OR2_X1 U8002 ( .A1(n6411), .A2(n6252), .ZN(n6253) );
  NAND4_X1 U8003 ( .A1(n6256), .A2(n6255), .A3(n6254), .A4(n6253), .ZN(n8746)
         );
  NAND2_X1 U8004 ( .A1(n8243), .A2(n8746), .ZN(n8757) );
  NAND2_X1 U8005 ( .A1(n7305), .A2(n8288), .ZN(n6260) );
  AOI22_X1 U8006 ( .A1(n6258), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n6421), .B2(
        n6257), .ZN(n6259) );
  AND2_X1 U8007 ( .A1(n6261), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6262) );
  NOR2_X2 U8008 ( .A1(n6261), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6269) );
  OR2_X1 U8009 ( .A1(n6262), .A2(n6269), .ZN(n8751) );
  NAND2_X1 U8010 ( .A1(n8751), .A2(n6308), .ZN(n6265) );
  AOI22_X1 U8011 ( .A1(n6090), .A2(P2_REG0_REG_19__SCAN_IN), .B1(n6321), .B2(
        P2_REG1_REG_19__SCAN_IN), .ZN(n6264) );
  OR2_X1 U8012 ( .A1(n6411), .A2(n5958), .ZN(n6263) );
  NOR2_X1 U8013 ( .A1(n8753), .A2(n8736), .ZN(n6266) );
  NAND2_X1 U8014 ( .A1(n7404), .A2(n8288), .ZN(n6268) );
  INV_X1 U8015 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7424) );
  OR2_X1 U8016 ( .A1(n8291), .A2(n7424), .ZN(n6267) );
  NOR2_X1 U8017 ( .A1(n6269), .A2(n10064), .ZN(n6270) );
  OR2_X1 U8018 ( .A1(n6278), .A2(n6270), .ZN(n8739) );
  NAND2_X1 U8019 ( .A1(n8739), .A2(n6308), .ZN(n6273) );
  AOI22_X1 U8020 ( .A1(n6090), .A2(P2_REG0_REG_20__SCAN_IN), .B1(n6321), .B2(
        P2_REG1_REG_20__SCAN_IN), .ZN(n6272) );
  INV_X1 U8021 ( .A(n6411), .ZN(n6309) );
  NAND2_X1 U8022 ( .A1(n6309), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n6271) );
  NAND2_X1 U8023 ( .A1(n8107), .A2(n8722), .ZN(n8723) );
  NAND2_X1 U8024 ( .A1(n8415), .A2(n8723), .ZN(n8738) );
  NAND2_X1 U8025 ( .A1(n7497), .A2(n8288), .ZN(n6277) );
  INV_X1 U8026 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7499) );
  OR2_X1 U8027 ( .A1(n8291), .A2(n7499), .ZN(n6276) );
  OR2_X1 U8028 ( .A1(n6278), .A2(n10000), .ZN(n6279) );
  NAND2_X1 U8029 ( .A1(n6287), .A2(n6279), .ZN(n8728) );
  NAND2_X1 U8030 ( .A1(n8728), .A2(n6308), .ZN(n6284) );
  INV_X1 U8031 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8914) );
  NAND2_X1 U8032 ( .A1(n6321), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n6281) );
  NAND2_X1 U8033 ( .A1(n6309), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n6280) );
  OAI211_X1 U8034 ( .C1(n6373), .C2(n8914), .A(n6281), .B(n6280), .ZN(n6282)
         );
  INV_X1 U8035 ( .A(n6282), .ZN(n6283) );
  NAND2_X1 U8036 ( .A1(n8727), .A2(n8735), .ZN(n8411) );
  NAND2_X1 U8037 ( .A1(n7515), .A2(n8288), .ZN(n6286) );
  OR2_X1 U8038 ( .A1(n8291), .A2(n7517), .ZN(n6285) );
  NAND2_X1 U8039 ( .A1(n6287), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6288) );
  NAND2_X1 U8040 ( .A1(n6296), .A2(n6288), .ZN(n8714) );
  NAND2_X1 U8041 ( .A1(n8714), .A2(n6308), .ZN(n6293) );
  INV_X1 U8042 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n8910) );
  NAND2_X1 U8043 ( .A1(n6309), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n6290) );
  NAND2_X1 U8044 ( .A1(n6321), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n6289) );
  OAI211_X1 U8045 ( .C1(n6373), .C2(n8910), .A(n6290), .B(n6289), .ZN(n6291)
         );
  INV_X1 U8046 ( .A(n6291), .ZN(n6292) );
  NAND2_X1 U8047 ( .A1(n8225), .A2(n8721), .ZN(n8422) );
  NAND2_X1 U8048 ( .A1(n8423), .A2(n8422), .ZN(n8713) );
  NAND2_X1 U8049 ( .A1(n7574), .A2(n8288), .ZN(n6295) );
  OR2_X1 U8050 ( .A1(n8291), .A2(n7577), .ZN(n6294) );
  AND2_X2 U8051 ( .A1(n6295), .A2(n6294), .ZN(n8908) );
  AND2_X1 U8052 ( .A1(n6296), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6297) );
  OR2_X1 U8053 ( .A1(n6306), .A2(n6297), .ZN(n8703) );
  NAND2_X1 U8054 ( .A1(n8703), .A2(n6308), .ZN(n6302) );
  INV_X1 U8055 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n8906) );
  NAND2_X1 U8056 ( .A1(n6309), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n6299) );
  NAND2_X1 U8057 ( .A1(n6321), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n6298) );
  OAI211_X1 U8058 ( .C1(n6373), .C2(n8906), .A(n6299), .B(n6298), .ZN(n6300)
         );
  INV_X1 U8059 ( .A(n6300), .ZN(n6301) );
  NAND2_X1 U8060 ( .A1(n8908), .A2(n8711), .ZN(n6303) );
  NAND2_X1 U8061 ( .A1(n7642), .A2(n8288), .ZN(n6305) );
  OR2_X1 U8062 ( .A1(n8291), .A2(n8137), .ZN(n6304) );
  OR2_X1 U8063 ( .A1(n6306), .A2(n10048), .ZN(n6307) );
  NAND2_X1 U8064 ( .A1(n10048), .A2(n6306), .ZN(n6323) );
  NAND2_X1 U8065 ( .A1(n6307), .A2(n6323), .ZN(n8691) );
  NAND2_X1 U8066 ( .A1(n8691), .A2(n6308), .ZN(n6314) );
  INV_X1 U8067 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n8902) );
  NAND2_X1 U8068 ( .A1(n6321), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n6311) );
  NAND2_X1 U8069 ( .A1(n6309), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n6310) );
  OAI211_X1 U8070 ( .C1(n6373), .C2(n8902), .A(n6311), .B(n6310), .ZN(n6312)
         );
  INV_X1 U8071 ( .A(n6312), .ZN(n6313) );
  NAND2_X1 U8072 ( .A1(n6318), .A2(n6317), .ZN(n8676) );
  NAND2_X1 U8073 ( .A1(n7684), .A2(n8288), .ZN(n6320) );
  OR2_X1 U8074 ( .A1(n8291), .A2(n8052), .ZN(n6319) );
  NAND2_X1 U8075 ( .A1(n6321), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n6327) );
  INV_X1 U8076 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n6322) );
  OR2_X1 U8077 ( .A1(n6411), .A2(n6322), .ZN(n6326) );
  AOI21_X1 U8078 ( .B1(P2_REG3_REG_25__SCAN_IN), .B2(n6323), .A(n6330), .ZN(
        n8680) );
  OR2_X1 U8079 ( .A1(n6211), .A2(n8680), .ZN(n6325) );
  INV_X1 U8080 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n8898) );
  OR2_X1 U8081 ( .A1(n6373), .A2(n8898), .ZN(n6324) );
  AND4_X2 U8082 ( .A1(n6327), .A2(n6326), .A3(n6325), .A4(n6324), .ZN(n8689)
         );
  OR2_X1 U8083 ( .A1(n8184), .A2(n8689), .ZN(n8434) );
  NAND2_X1 U8084 ( .A1(n8434), .A2(n8427), .ZN(n8683) );
  AOI22_X1 U8085 ( .A1(n8676), .A2(n8683), .B1(n8689), .B2(n8900), .ZN(n8663)
         );
  NAND2_X1 U8086 ( .A1(n7687), .A2(n8288), .ZN(n6329) );
  OR2_X1 U8087 ( .A1(n8291), .A2(n7690), .ZN(n6328) );
  NAND2_X1 U8088 ( .A1(n6090), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6336) );
  INV_X1 U8089 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8820) );
  OR2_X1 U8090 ( .A1(n4359), .A2(n8820), .ZN(n6335) );
  INV_X1 U8091 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n10108) );
  NAND2_X1 U8092 ( .A1(n10108), .A2(n6330), .ZN(n6343) );
  INV_X1 U8093 ( .A(n6330), .ZN(n6331) );
  NAND2_X1 U8094 ( .A1(P2_REG3_REG_26__SCAN_IN), .A2(n6331), .ZN(n6332) );
  AND2_X1 U8095 ( .A1(n6343), .A2(n6332), .ZN(n8667) );
  INV_X1 U8096 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8668) );
  OR2_X1 U8097 ( .A1(n6411), .A2(n8668), .ZN(n6333) );
  OR2_X1 U8098 ( .A1(n8670), .A2(n8678), .ZN(n8439) );
  NAND2_X1 U8099 ( .A1(n8670), .A2(n8678), .ZN(n8440) );
  NAND2_X1 U8100 ( .A1(n8439), .A2(n8440), .ZN(n8662) );
  INV_X1 U8101 ( .A(n8670), .ZN(n8896) );
  INV_X1 U8102 ( .A(n8678), .ZN(n6337) );
  NAND2_X1 U8103 ( .A1(n8670), .A2(n6337), .ZN(n6338) );
  NAND2_X1 U8104 ( .A1(n8661), .A2(n6338), .ZN(n8649) );
  INV_X1 U8105 ( .A(n8649), .ZN(n6350) );
  OR2_X1 U8106 ( .A1(n8291), .A2(n8958), .ZN(n6339) );
  NAND2_X1 U8107 ( .A1(n6090), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6348) );
  INV_X1 U8108 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n6341) );
  OR2_X1 U8109 ( .A1(n4360), .A2(n6341), .ZN(n6347) );
  INV_X1 U8110 ( .A(n6343), .ZN(n6342) );
  INV_X1 U8111 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n10090) );
  NAND2_X1 U8112 ( .A1(n6342), .A2(n10090), .ZN(n6355) );
  NAND2_X1 U8113 ( .A1(n6343), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6344) );
  AND2_X1 U8114 ( .A1(n6355), .A2(n6344), .ZN(n8653) );
  OR2_X1 U8115 ( .A1(n6211), .A2(n8653), .ZN(n6346) );
  INV_X1 U8116 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n8654) );
  OR2_X1 U8117 ( .A1(n6411), .A2(n8654), .ZN(n6345) );
  NAND2_X1 U8118 ( .A1(n8890), .A2(n8664), .ZN(n6349) );
  NAND2_X1 U8119 ( .A1(n6351), .A2(n8288), .ZN(n6353) );
  OR2_X1 U8120 ( .A1(n8291), .A2(n8957), .ZN(n6352) );
  NAND2_X1 U8121 ( .A1(n6090), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6360) );
  INV_X1 U8122 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n6354) );
  OR2_X1 U8123 ( .A1(n4360), .A2(n6354), .ZN(n6359) );
  NAND2_X1 U8124 ( .A1(n6355), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n6356) );
  OR2_X1 U8125 ( .A1(n6211), .A2(n8641), .ZN(n6358) );
  INV_X1 U8126 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n8642) );
  OR2_X1 U8127 ( .A1(n6411), .A2(n8642), .ZN(n6357) );
  XNOR2_X1 U8128 ( .A(n8647), .B(n8650), .ZN(n8493) );
  INV_X1 U8129 ( .A(n8650), .ZN(n8522) );
  NAND2_X1 U8130 ( .A1(n6362), .A2(n6361), .ZN(n6364) );
  MUX2_X1 U8131 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .S(n6491), .Z(n7815) );
  INV_X1 U8132 ( .A(n6365), .ZN(n6367) );
  INV_X1 U8133 ( .A(SI_29_), .ZN(n6366) );
  NAND2_X1 U8134 ( .A1(n6367), .A2(n6366), .ZN(n6368) );
  OR2_X1 U8135 ( .A1(n8951), .A2(n6369), .ZN(n6371) );
  INV_X1 U8136 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8952) );
  OR2_X1 U8137 ( .A1(n8291), .A2(n8952), .ZN(n6370) );
  INV_X1 U8138 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n6372) );
  OR2_X1 U8139 ( .A1(n6373), .A2(n6372), .ZN(n6377) );
  INV_X1 U8140 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6374) );
  OR2_X1 U8141 ( .A1(n4359), .A2(n6374), .ZN(n6376) );
  INV_X1 U8142 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n7700) );
  OR2_X1 U8143 ( .A1(n6411), .A2(n7700), .ZN(n6375) );
  OR2_X2 U8144 ( .A1(n8307), .A2(n8638), .ZN(n8502) );
  NAND2_X1 U8145 ( .A1(n8307), .A2(n8638), .ZN(n8452) );
  NAND2_X1 U8146 ( .A1(n8502), .A2(n8452), .ZN(n8496) );
  NAND2_X1 U8147 ( .A1(n6421), .A2(n8516), .ZN(n6441) );
  NAND2_X1 U8148 ( .A1(n6379), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6380) );
  NAND2_X1 U8149 ( .A1(n8310), .A2(n8512), .ZN(n8304) );
  NAND2_X1 U8150 ( .A1(n6381), .A2(n8759), .ZN(n6419) );
  NAND2_X1 U8151 ( .A1(n6874), .A2(n8325), .ZN(n6992) );
  INV_X1 U8152 ( .A(n9834), .ZN(n6993) );
  NAND2_X1 U8153 ( .A1(n8539), .A2(n6993), .ZN(n8332) );
  INV_X1 U8154 ( .A(n6987), .ZN(n8469) );
  NAND2_X1 U8155 ( .A1(n6992), .A2(n8469), .ZN(n6384) );
  NAND2_X1 U8156 ( .A1(n6384), .A2(n8338), .ZN(n6938) );
  INV_X1 U8157 ( .A(n6943), .ZN(n9841) );
  OR2_X1 U8158 ( .A1(n8538), .A2(n9841), .ZN(n8333) );
  NAND2_X1 U8159 ( .A1(n8538), .A2(n9841), .ZN(n8341) );
  NAND2_X1 U8160 ( .A1(n8333), .A2(n8341), .ZN(n8471) );
  INV_X1 U8161 ( .A(n8471), .ZN(n8339) );
  NAND2_X1 U8162 ( .A1(n6938), .A2(n8339), .ZN(n6385) );
  NAND2_X1 U8163 ( .A1(n6385), .A2(n8333), .ZN(n7032) );
  INV_X1 U8164 ( .A(n9845), .ZN(n6386) );
  OR2_X1 U8165 ( .A1(n8537), .A2(n6386), .ZN(n8344) );
  NAND2_X1 U8166 ( .A1(n8537), .A2(n6386), .ZN(n8342) );
  NAND2_X1 U8167 ( .A1(n8344), .A2(n8342), .ZN(n8472) );
  INV_X1 U8168 ( .A(n8472), .ZN(n7033) );
  NAND2_X1 U8169 ( .A1(n7032), .A2(n7033), .ZN(n7031) );
  NAND2_X1 U8170 ( .A1(n7031), .A2(n8344), .ZN(n7227) );
  INV_X1 U8171 ( .A(n8345), .ZN(n6387) );
  NAND2_X1 U8172 ( .A1(n7295), .A2(n8475), .ZN(n6388) );
  NAND2_X1 U8173 ( .A1(n8350), .A2(n8535), .ZN(n8362) );
  NAND2_X1 U8174 ( .A1(n6388), .A2(n8362), .ZN(n7122) );
  INV_X1 U8175 ( .A(n8363), .ZN(n6389) );
  OR2_X1 U8176 ( .A1(n7996), .A2(n7561), .ZN(n8373) );
  NAND2_X1 U8177 ( .A1(n7989), .A2(n8373), .ZN(n6391) );
  NAND2_X1 U8178 ( .A1(n7996), .A2(n7561), .ZN(n8371) );
  NAND2_X1 U8179 ( .A1(n6391), .A2(n8371), .ZN(n7449) );
  INV_X1 U8180 ( .A(n8529), .ZN(n7589) );
  AND2_X1 U8181 ( .A1(n8388), .A2(n7589), .ZN(n6395) );
  OR2_X1 U8182 ( .A1(n8379), .A2(n6395), .ZN(n6392) );
  OR2_X1 U8183 ( .A1(n8388), .A2(n7589), .ZN(n6393) );
  AND2_X1 U8184 ( .A1(n6393), .A2(n8383), .ZN(n6394) );
  OR2_X1 U8185 ( .A1(n7590), .A2(n8096), .ZN(n8396) );
  AND2_X1 U8186 ( .A1(n7590), .A2(n8096), .ZN(n7586) );
  NAND2_X1 U8187 ( .A1(n8794), .A2(n8402), .ZN(n6397) );
  NAND2_X1 U8188 ( .A1(n6397), .A2(n8403), .ZN(n8778) );
  NAND2_X1 U8189 ( .A1(n8778), .A2(n8407), .ZN(n6398) );
  AND2_X1 U8190 ( .A1(n8925), .A2(n8746), .ZN(n8464) );
  INV_X1 U8191 ( .A(n8746), .ZN(n8776) );
  NAND2_X1 U8192 ( .A1(n8243), .A2(n8776), .ZN(n8463) );
  OAI21_X1 U8193 ( .B1(n8768), .B2(n8464), .A(n8463), .ZN(n8750) );
  OR2_X1 U8194 ( .A1(n8846), .A2(n8736), .ZN(n8414) );
  NAND2_X1 U8195 ( .A1(n8846), .A2(n8736), .ZN(n8413) );
  NAND2_X1 U8196 ( .A1(n8750), .A2(n8749), .ZN(n8748) );
  NAND2_X1 U8197 ( .A1(n8748), .A2(n8413), .ZN(n8737) );
  NAND2_X1 U8198 ( .A1(n8737), .A2(n8415), .ZN(n8724) );
  AND2_X1 U8199 ( .A1(n8411), .A2(n8723), .ZN(n8418) );
  NAND2_X1 U8200 ( .A1(n8724), .A2(n8418), .ZN(n6399) );
  NAND2_X1 U8201 ( .A1(n6399), .A2(n8420), .ZN(n8712) );
  NAND2_X1 U8202 ( .A1(n6316), .A2(n8700), .ZN(n8459) );
  NAND2_X1 U8203 ( .A1(n8160), .A2(n8711), .ZN(n8692) );
  AND2_X1 U8204 ( .A1(n8459), .A2(n8692), .ZN(n8432) );
  NAND2_X1 U8205 ( .A1(n6400), .A2(n8460), .ZN(n8682) );
  NAND2_X1 U8206 ( .A1(n8682), .A2(n8427), .ZN(n6401) );
  INV_X1 U8207 ( .A(n8439), .ZN(n6402) );
  NAND2_X1 U8208 ( .A1(n8890), .A2(n8639), .ZN(n8444) );
  NAND2_X1 U8209 ( .A1(n8644), .A2(n8643), .ZN(n6404) );
  OR2_X1 U8210 ( .A1(n8647), .A2(n8650), .ZN(n6403) );
  NAND2_X1 U8211 ( .A1(n6405), .A2(n8516), .ZN(n6450) );
  NAND2_X1 U8212 ( .A1(n8310), .A2(n7426), .ZN(n8501) );
  OR2_X1 U8213 ( .A1(n6450), .A2(n8501), .ZN(n6443) );
  INV_X1 U8214 ( .A(n8516), .ZN(n7519) );
  NAND2_X1 U8215 ( .A1(n7519), .A2(n8315), .ZN(n9861) );
  NAND2_X1 U8216 ( .A1(n6783), .A2(n6450), .ZN(n6406) );
  NAND3_X1 U8217 ( .A1(n6443), .A2(n9861), .A3(n6406), .ZN(n6936) );
  XNOR2_X1 U8218 ( .A(n8514), .B(n6407), .ZN(n6415) );
  NAND2_X1 U8219 ( .A1(n6076), .A2(P2_B_REG_SCAN_IN), .ZN(n6408) );
  AND2_X1 U8220 ( .A1(n8763), .A2(n6408), .ZN(n8632) );
  NAND2_X1 U8221 ( .A1(n6090), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n6414) );
  INV_X1 U8222 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n6409) );
  OR2_X1 U8223 ( .A1(n4360), .A2(n6409), .ZN(n6413) );
  INV_X1 U8224 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n6410) );
  OR2_X1 U8225 ( .A1(n6411), .A2(n6410), .ZN(n6412) );
  NAND4_X1 U8226 ( .A1(n8299), .A2(n6414), .A3(n6413), .A4(n6412), .ZN(n8521)
         );
  INV_X1 U8227 ( .A(n6415), .ZN(n6795) );
  AOI22_X1 U8228 ( .A1(n8632), .A2(n8521), .B1(n8522), .B2(n8745), .ZN(n6416)
         );
  OAI21_X1 U8229 ( .B1(n6420), .B2(n6936), .A(n6416), .ZN(n6417) );
  INV_X1 U8230 ( .A(n6417), .ZN(n6418) );
  NAND2_X1 U8231 ( .A1(n6421), .A2(n7426), .ZN(n6851) );
  XNOR2_X1 U8232 ( .A(n6422), .B(P2_B_REG_SCAN_IN), .ZN(n6423) );
  NAND2_X1 U8233 ( .A1(n6424), .A2(n6423), .ZN(n6426) );
  OR2_X1 U8234 ( .A1(n6439), .A2(P2_D_REG_1__SCAN_IN), .ZN(n6427) );
  NAND2_X1 U8235 ( .A1(n6424), .A2(n7692), .ZN(n6614) );
  NOR2_X1 U8236 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .ZN(
        n6431) );
  NOR4_X1 U8237 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n6430) );
  NOR4_X1 U8238 ( .A1(P2_D_REG_12__SCAN_IN), .A2(P2_D_REG_25__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_23__SCAN_IN), .ZN(n6429) );
  NOR4_X1 U8239 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_28__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_26__SCAN_IN), .ZN(n6428) );
  NAND4_X1 U8240 ( .A1(n6431), .A2(n6430), .A3(n6429), .A4(n6428), .ZN(n6437)
         );
  NOR4_X1 U8241 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n6435) );
  NOR4_X1 U8242 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_15__SCAN_IN), .ZN(n6434) );
  NOR4_X1 U8243 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6433) );
  NOR4_X1 U8244 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n6432) );
  NAND4_X1 U8245 ( .A1(n6435), .A2(n6434), .A3(n6433), .A4(n6432), .ZN(n6436)
         );
  NOR2_X1 U8246 ( .A1(n6437), .A2(n6436), .ZN(n6438) );
  NOR2_X1 U8247 ( .A1(n6848), .A2(n6445), .ZN(n6440) );
  NAND2_X1 U8248 ( .A1(n6422), .A2(n7692), .ZN(n6617) );
  NAND2_X1 U8249 ( .A1(n8315), .A2(n8512), .ZN(n8466) );
  INV_X1 U8250 ( .A(n6726), .ZN(n6744) );
  AND2_X1 U8251 ( .A1(n8446), .A2(n9861), .ZN(n6442) );
  NAND2_X1 U8252 ( .A1(n6744), .A2(n6442), .ZN(n6728) );
  NAND2_X1 U8253 ( .A1(n6851), .A2(n9871), .ZN(n8686) );
  NAND2_X1 U8254 ( .A1(n6728), .A2(n8686), .ZN(n6739) );
  NAND2_X1 U8255 ( .A1(n6727), .A2(n6739), .ZN(n6447) );
  INV_X1 U8256 ( .A(n6848), .ZN(n6444) );
  NOR2_X1 U8257 ( .A1(n6455), .A2(n6445), .ZN(n6741) );
  OAI21_X1 U8258 ( .B1(n6726), .B2(n6998), .A(n6732), .ZN(n6446) );
  INV_X1 U8259 ( .A(n8307), .ZN(n6459) );
  NAND2_X1 U8260 ( .A1(n6449), .A2(n4445), .ZN(P2_U3456) );
  NOR2_X1 U8261 ( .A1(n6846), .A2(n6733), .ZN(n6452) );
  OR2_X1 U8262 ( .A1(n6450), .A2(n7426), .ZN(n6451) );
  AND2_X1 U8263 ( .A1(n6451), .A2(n8446), .ZN(n6847) );
  MUX2_X1 U8264 ( .A(n6848), .B(n6452), .S(n6847), .Z(n6456) );
  NAND2_X1 U8265 ( .A1(n6783), .A2(n8454), .ZN(n6736) );
  AND3_X1 U8266 ( .A1(n6453), .A2(n6746), .A3(n6736), .ZN(n6454) );
  NAND2_X1 U8267 ( .A1(n6458), .A2(n4458), .ZN(n6460) );
  NAND2_X1 U8268 ( .A1(n6460), .A2(n4443), .ZN(P2_U3488) );
  INV_X1 U8269 ( .A(n6461), .ZN(n6462) );
  NOR2_X1 U8270 ( .A1(n6465), .A2(n6464), .ZN(n6466) );
  NOR2_X1 U8271 ( .A1(n8085), .A2(n9524), .ZN(n6469) );
  OAI22_X1 U8272 ( .A1(n9814), .A2(n6499), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6470), .ZN(n6486) );
  INV_X1 U8273 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n9891) );
  NOR2_X1 U8274 ( .A1(n8628), .A2(n9891), .ZN(n6485) );
  INV_X1 U8275 ( .A(n9807), .ZN(n8624) );
  AOI211_X1 U8276 ( .C1(n6473), .C2(n6472), .A(n6471), .B(n8624), .ZN(n6484)
         );
  INV_X1 U8277 ( .A(n6474), .ZN(n6475) );
  AOI21_X1 U8278 ( .B1(n6845), .B2(n6476), .A(n6475), .ZN(n6482) );
  INV_X1 U8279 ( .A(n6477), .ZN(n6478) );
  AOI21_X1 U8280 ( .B1(n6480), .B2(n6479), .A(n6478), .ZN(n6481) );
  OAI22_X1 U8281 ( .A1(n6482), .A2(n9803), .B1(n9810), .B2(n6481), .ZN(n6483)
         );
  OR4_X1 U8282 ( .A1(n6486), .A2(n6485), .A3(n6484), .A4(n6483), .ZN(P2_U3183)
         );
  INV_X2 U8283 ( .A(n7571), .ZN(n9591) );
  INV_X1 U8284 ( .A(n9145), .ZN(n6487) );
  OAI222_X1 U8285 ( .A1(n9588), .A2(n6488), .B1(n9591), .B2(n6498), .C1(
        P1_U3086), .C2(n6487), .ZN(P1_U3354) );
  OAI222_X1 U8286 ( .A1(n9588), .A2(n6489), .B1(n9591), .B2(n6494), .C1(
        P1_U3086), .C2(n6540), .ZN(P1_U3353) );
  OAI222_X1 U8287 ( .A1(n9588), .A2(n6490), .B1(n9591), .B2(n6492), .C1(
        P1_U3086), .C2(n6545), .ZN(P1_U3352) );
  AND2_X1 U8288 ( .A1(n7825), .A2(P2_U3151), .ZN(n8953) );
  INV_X2 U8289 ( .A(n8953), .ZN(n8960) );
  NAND2_X2 U8290 ( .A1(n6491), .A2(P2_U3151), .ZN(n8956) );
  OAI222_X1 U8291 ( .A1(n6493), .A2(P2_U3151), .B1(n8960), .B2(n6492), .C1(
        n5084), .C2(n8956), .ZN(P2_U3292) );
  OAI222_X1 U8292 ( .A1(n5966), .A2(P2_U3151), .B1(n8960), .B2(n6494), .C1(
        n5061), .C2(n8956), .ZN(P2_U3293) );
  OAI222_X1 U8293 ( .A1(n9588), .A2(n6495), .B1(n9591), .B2(n6496), .C1(
        P1_U3086), .C2(n6547), .ZN(P1_U3351) );
  OAI222_X1 U8294 ( .A1(n6694), .A2(P2_U3151), .B1(n8960), .B2(n6496), .C1(
        n5117), .C2(n8956), .ZN(P2_U3291) );
  OAI222_X1 U8295 ( .A1(n6499), .A2(P2_U3151), .B1(n8960), .B2(n6498), .C1(
        n6497), .C2(n8956), .ZN(P2_U3294) );
  OAI222_X1 U8296 ( .A1(n9795), .A2(P2_U3151), .B1(n8960), .B2(n6501), .C1(
        n6500), .C2(n8956), .ZN(P2_U3290) );
  OAI222_X1 U8297 ( .A1(n9588), .A2(n6502), .B1(n9591), .B2(n6501), .C1(
        P1_U3086), .C2(n6535), .ZN(P1_U3350) );
  INV_X1 U8298 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6503) );
  OAI222_X1 U8299 ( .A1(n6764), .A2(P2_U3151), .B1(n8960), .B2(n6504), .C1(
        n6503), .C2(n8956), .ZN(P2_U3289) );
  OAI222_X1 U8300 ( .A1(n9588), .A2(n6505), .B1(n9591), .B2(n6504), .C1(
        P1_U3086), .C2(n6555), .ZN(P1_U3349) );
  OR2_X1 U8301 ( .A1(n6507), .A2(P1_U3086), .ZN(n7986) );
  NAND2_X1 U8302 ( .A1(n6506), .A2(n7986), .ZN(n6518) );
  INV_X1 U8303 ( .A(n6518), .ZN(n6510) );
  NAND2_X1 U8304 ( .A1(n6508), .A2(n6507), .ZN(n6509) );
  AND2_X1 U8305 ( .A1(n5038), .A2(n6509), .ZN(n6519) );
  OR2_X1 U8306 ( .A1(n6510), .A2(n6519), .ZN(n9722) );
  INV_X1 U8307 ( .A(n9722), .ZN(n9188) );
  NOR2_X1 U8308 ( .A1(n9188), .A2(P1_U3973), .ZN(P1_U3085) );
  INV_X1 U8309 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6511) );
  OAI222_X1 U8310 ( .A1(n6951), .A2(P2_U3151), .B1(n8960), .B2(n6513), .C1(
        n6511), .C2(n8956), .ZN(P2_U3288) );
  INV_X1 U8311 ( .A(n6600), .ZN(n6512) );
  OAI222_X1 U8312 ( .A1(n9588), .A2(n6514), .B1(n9591), .B2(n6513), .C1(
        P1_U3086), .C2(n6512), .ZN(P1_U3348) );
  INV_X1 U8313 ( .A(n6515), .ZN(n9154) );
  INV_X1 U8314 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n6516) );
  AOI21_X1 U8315 ( .B1(n9154), .B2(n6516), .A(n5726), .ZN(n9160) );
  OAI21_X1 U8316 ( .B1(P1_REG1_REG_0__SCAN_IN), .B2(n9154), .A(n9160), .ZN(
        n6517) );
  XOR2_X1 U8317 ( .A(P1_IR_REG_0__SCAN_IN), .B(n6517), .Z(n6521) );
  NAND2_X1 U8318 ( .A1(n6519), .A2(n6518), .ZN(n6554) );
  AOI22_X1 U8319 ( .A1(n9188), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n6520) );
  OAI21_X1 U8320 ( .B1(n6521), .B2(n6554), .A(n6520), .ZN(P1_U3243) );
  AND2_X1 U8321 ( .A1(n6613), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U8322 ( .A1(n6613), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U8323 ( .A1(n6613), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U8324 ( .A1(n6613), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U8325 ( .A1(n6613), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U8326 ( .A1(n6613), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U8327 ( .A1(n6613), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U8328 ( .A1(n6613), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U8329 ( .A1(n6613), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U8330 ( .A1(n6613), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U8331 ( .A1(n6613), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U8332 ( .A1(n6613), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U8333 ( .A1(n6613), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  OAI222_X1 U8334 ( .A1(n9588), .A2(n6522), .B1(n9591), .B2(n6524), .C1(
        P1_U3086), .C2(n6604), .ZN(P1_U3347) );
  OAI222_X1 U8335 ( .A1(n7048), .A2(P2_U3151), .B1(n8960), .B2(n6524), .C1(
        n6523), .C2(n8956), .ZN(P2_U3287) );
  INV_X1 U8336 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6529) );
  NAND2_X1 U8337 ( .A1(n5097), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6527) );
  NAND2_X1 U8338 ( .A1(n5098), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6526) );
  NAND2_X1 U8339 ( .A1(n4358), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6525) );
  AND3_X1 U8340 ( .A1(n6527), .A2(n6526), .A3(n6525), .ZN(n7840) );
  INV_X1 U8341 ( .A(n7840), .ZN(n9205) );
  NAND2_X1 U8342 ( .A1(n9205), .A2(P1_U3973), .ZN(n6528) );
  OAI21_X1 U8343 ( .B1(P1_U3973), .B2(n6529), .A(n6528), .ZN(P1_U3585) );
  INV_X1 U8344 ( .A(n6535), .ZN(n6568) );
  INV_X1 U8345 ( .A(n6547), .ZN(n9192) );
  INV_X1 U8346 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6530) );
  MUX2_X1 U8347 ( .A(n6530), .B(P1_REG1_REG_2__SCAN_IN), .S(n6540), .Z(n9170)
         );
  INV_X1 U8348 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n9750) );
  MUX2_X1 U8349 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n9750), .S(n9145), .Z(n9148)
         );
  AND2_X1 U8350 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n9147) );
  NAND2_X1 U8351 ( .A1(n9148), .A2(n9147), .ZN(n9146) );
  NAND2_X1 U8352 ( .A1(n9145), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6531) );
  NAND2_X1 U8353 ( .A1(n9146), .A2(n6531), .ZN(n9169) );
  NAND2_X1 U8354 ( .A1(n9170), .A2(n9169), .ZN(n9168) );
  INV_X1 U8355 ( .A(n6540), .ZN(n9164) );
  NAND2_X1 U8356 ( .A1(n9164), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6532) );
  NAND2_X1 U8357 ( .A1(n9168), .A2(n6532), .ZN(n9182) );
  XNOR2_X1 U8358 ( .A(n6545), .B(P1_REG1_REG_3__SCAN_IN), .ZN(n9183) );
  NAND2_X1 U8359 ( .A1(n9182), .A2(n9183), .ZN(n9181) );
  INV_X1 U8360 ( .A(n6545), .ZN(n9177) );
  NAND2_X1 U8361 ( .A1(n9177), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6533) );
  NAND2_X1 U8362 ( .A1(n9181), .A2(n6533), .ZN(n9190) );
  XNOR2_X1 U8363 ( .A(n6547), .B(P1_REG1_REG_4__SCAN_IN), .ZN(n9191) );
  NAND2_X1 U8364 ( .A1(n9190), .A2(n9191), .ZN(n9189) );
  INV_X1 U8365 ( .A(n9189), .ZN(n6534) );
  AOI21_X1 U8366 ( .B1(n9192), .B2(P1_REG1_REG_4__SCAN_IN), .A(n6534), .ZN(
        n6564) );
  XOR2_X1 U8367 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n6535), .Z(n6563) );
  NOR2_X1 U8368 ( .A1(n6564), .A2(n6563), .ZN(n6562) );
  AOI21_X1 U8369 ( .B1(n6568), .B2(P1_REG1_REG_5__SCAN_IN), .A(n6562), .ZN(
        n6539) );
  INV_X1 U8370 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6536) );
  MUX2_X1 U8371 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n6536), .S(n6555), .Z(n6538)
         );
  NOR2_X1 U8372 ( .A1(n6539), .A2(n6538), .ZN(n6578) );
  INV_X1 U8373 ( .A(n6554), .ZN(n6537) );
  AOI211_X1 U8374 ( .C1(n6539), .C2(n6538), .A(n6578), .B(n9669), .ZN(n6561)
         );
  INV_X1 U8375 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6541) );
  MUX2_X1 U8376 ( .A(n6541), .B(P1_REG2_REG_2__SCAN_IN), .S(n6540), .Z(n9167)
         );
  INV_X1 U8377 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6542) );
  MUX2_X1 U8378 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n6542), .S(n9145), .Z(n9150)
         );
  AND2_X1 U8379 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n9155) );
  NAND2_X1 U8380 ( .A1(n9150), .A2(n9155), .ZN(n9149) );
  NAND2_X1 U8381 ( .A1(n9145), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6543) );
  NAND2_X1 U8382 ( .A1(n9149), .A2(n6543), .ZN(n9166) );
  NAND2_X1 U8383 ( .A1(n9167), .A2(n9166), .ZN(n9165) );
  NAND2_X1 U8384 ( .A1(n9164), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6544) );
  NAND2_X1 U8385 ( .A1(n9165), .A2(n6544), .ZN(n9179) );
  XNOR2_X1 U8386 ( .A(n6545), .B(P1_REG2_REG_3__SCAN_IN), .ZN(n9180) );
  NAND2_X1 U8387 ( .A1(n9179), .A2(n9180), .ZN(n9178) );
  NAND2_X1 U8388 ( .A1(n9177), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6546) );
  NAND2_X1 U8389 ( .A1(n9178), .A2(n6546), .ZN(n9196) );
  XNOR2_X1 U8390 ( .A(n6547), .B(P1_REG2_REG_4__SCAN_IN), .ZN(n9197) );
  NAND2_X1 U8391 ( .A1(n9196), .A2(n9197), .ZN(n9195) );
  INV_X1 U8392 ( .A(n9195), .ZN(n6548) );
  XNOR2_X1 U8393 ( .A(n6568), .B(P1_REG2_REG_5__SCAN_IN), .ZN(n6566) );
  NOR2_X1 U8394 ( .A1(n6567), .A2(n6566), .ZN(n6565) );
  INV_X1 U8395 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6549) );
  MUX2_X1 U8396 ( .A(n6549), .B(P1_REG2_REG_6__SCAN_IN), .S(n6555), .Z(n6550)
         );
  INV_X1 U8397 ( .A(n6550), .ZN(n6552) );
  NOR2_X1 U8398 ( .A1(n6553), .A2(n6552), .ZN(n6575) );
  OR2_X1 U8399 ( .A1(n5726), .A2(n6515), .ZN(n6551) );
  AOI211_X1 U8400 ( .C1(n6553), .C2(n6552), .A(n6575), .B(n9686), .ZN(n6560)
         );
  INV_X1 U8401 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n6558) );
  INV_X1 U8402 ( .A(n6555), .ZN(n6579) );
  NAND2_X1 U8403 ( .A1(n9699), .A2(n6579), .ZN(n6557) );
  NAND2_X1 U8404 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3086), .ZN(n6556) );
  OAI211_X1 U8405 ( .C1(n6558), .C2(n9722), .A(n6557), .B(n6556), .ZN(n6559)
         );
  OR3_X1 U8406 ( .A1(n6561), .A2(n6560), .A3(n6559), .ZN(P1_U3249) );
  AOI211_X1 U8407 ( .C1(n6564), .C2(n6563), .A(n6562), .B(n9669), .ZN(n6574)
         );
  AOI211_X1 U8408 ( .C1(n6567), .C2(n6566), .A(n6565), .B(n9686), .ZN(n6573)
         );
  INV_X1 U8409 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n6571) );
  NAND2_X1 U8410 ( .A1(n9699), .A2(n6568), .ZN(n6570) );
  NAND2_X1 U8411 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n6569) );
  OAI211_X1 U8412 ( .C1(n6571), .C2(n9722), .A(n6570), .B(n6569), .ZN(n6572)
         );
  OR3_X1 U8413 ( .A1(n6574), .A2(n6573), .A3(n6572), .ZN(P1_U3248) );
  AOI21_X1 U8414 ( .B1(n6579), .B2(P1_REG2_REG_6__SCAN_IN), .A(n6575), .ZN(
        n6577) );
  XNOR2_X1 U8415 ( .A(n6600), .B(P1_REG2_REG_7__SCAN_IN), .ZN(n6576) );
  NOR2_X1 U8416 ( .A1(n6577), .A2(n6576), .ZN(n6599) );
  AOI211_X1 U8417 ( .C1(n6577), .C2(n6576), .A(n9686), .B(n6599), .ZN(n6587)
         );
  AOI21_X1 U8418 ( .B1(n6579), .B2(P1_REG1_REG_6__SCAN_IN), .A(n6578), .ZN(
        n6581) );
  XNOR2_X1 U8419 ( .A(n6600), .B(P1_REG1_REG_7__SCAN_IN), .ZN(n6580) );
  NOR2_X1 U8420 ( .A1(n6581), .A2(n6580), .ZN(n6595) );
  AOI211_X1 U8421 ( .C1(n6581), .C2(n6580), .A(n9669), .B(n6595), .ZN(n6586)
         );
  INV_X1 U8422 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n6584) );
  NAND2_X1 U8423 ( .A1(n9699), .A2(n6600), .ZN(n6583) );
  NAND2_X1 U8424 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n6582) );
  OAI211_X1 U8425 ( .C1(n6584), .C2(n9722), .A(n6583), .B(n6582), .ZN(n6585)
         );
  OR3_X1 U8426 ( .A1(n6587), .A2(n6586), .A3(n6585), .ZN(P1_U3250) );
  INV_X1 U8427 ( .A(n6165), .ZN(n6591) );
  INV_X1 U8428 ( .A(n9588), .ZN(n9585) );
  AOI22_X1 U8429 ( .A1(n9611), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n9585), .ZN(n6588) );
  OAI21_X1 U8430 ( .B1(n6591), .B2(n9591), .A(n6588), .ZN(P1_U3346) );
  NAND2_X1 U8431 ( .A1(n8621), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n6589) );
  OAI21_X1 U8432 ( .B1(n8789), .B2(n8621), .A(n6589), .ZN(P2_U3508) );
  OAI222_X1 U8433 ( .A1(P2_U3151), .A2(n6592), .B1(n8960), .B2(n6591), .C1(
        n6590), .C2(n8956), .ZN(P2_U3286) );
  INV_X1 U8434 ( .A(n6593), .ZN(n6611) );
  INV_X1 U8435 ( .A(n9601), .ZN(n6915) );
  OAI222_X1 U8436 ( .A1(n9591), .A2(n6611), .B1(n6915), .B2(P1_U3086), .C1(
        n6594), .C2(n9588), .ZN(P1_U3345) );
  AOI21_X1 U8437 ( .B1(P1_REG1_REG_7__SCAN_IN), .B2(n6600), .A(n6595), .ZN(
        n6598) );
  INV_X1 U8438 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6596) );
  MUX2_X1 U8439 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n6596), .S(n6604), .Z(n6597)
         );
  NOR2_X1 U8440 ( .A1(n6598), .A2(n6597), .ZN(n6924) );
  AOI211_X1 U8441 ( .C1(n6598), .C2(n6597), .A(n9669), .B(n6924), .ZN(n6609)
         );
  INV_X1 U8442 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n6601) );
  MUX2_X1 U8443 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n6601), .S(n6604), .Z(n6602)
         );
  NOR2_X1 U8444 ( .A1(n6603), .A2(n6602), .ZN(n6916) );
  AOI211_X1 U8445 ( .C1(n6603), .C2(n6602), .A(n9686), .B(n6916), .ZN(n6608)
         );
  INV_X1 U8446 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n6606) );
  INV_X1 U8447 ( .A(n6604), .ZN(n6925) );
  NAND2_X1 U8448 ( .A1(n9699), .A2(n6925), .ZN(n6605) );
  NAND2_X1 U8449 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n7287) );
  OAI211_X1 U8450 ( .C1(n6606), .C2(n9722), .A(n6605), .B(n7287), .ZN(n6607)
         );
  OR3_X1 U8451 ( .A1(n6609), .A2(n6608), .A3(n6607), .ZN(P1_U3251) );
  OAI222_X1 U8452 ( .A1(P2_U3151), .A2(n6612), .B1(n8960), .B2(n6611), .C1(
        n6610), .C2(n8956), .ZN(P2_U3285) );
  INV_X1 U8453 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n6616) );
  INV_X1 U8454 ( .A(n6614), .ZN(n6615) );
  AOI22_X1 U8455 ( .A1(n6613), .A2(n6616), .B1(n6619), .B2(n6615), .ZN(
        P2_U3377) );
  INV_X1 U8456 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n6620) );
  INV_X1 U8457 ( .A(n6617), .ZN(n6618) );
  AOI22_X1 U8458 ( .A1(n6613), .A2(n6620), .B1(n6619), .B2(n6618), .ZN(
        P2_U3376) );
  XNOR2_X1 U8459 ( .A(n6622), .B(n6621), .ZN(n9156) );
  NAND2_X1 U8460 ( .A1(n6624), .A2(n6623), .ZN(n6681) );
  AOI22_X1 U8461 ( .A1(n9628), .A2(n7013), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        n6681), .ZN(n6626) );
  OR2_X1 U8462 ( .A1(n9095), .A2(n9414), .ZN(n8988) );
  INV_X1 U8463 ( .A(n8988), .ZN(n9104) );
  NAND2_X1 U8464 ( .A1(n9104), .A2(n5737), .ZN(n6625) );
  OAI211_X1 U8465 ( .C1(n9156), .C2(n9623), .A(n6626), .B(n6625), .ZN(P1_U3232) );
  AND2_X1 U8466 ( .A1(n6613), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U8467 ( .A1(n6613), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U8468 ( .A1(n6613), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  AND2_X1 U8469 ( .A1(n6613), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U8470 ( .A1(n6613), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U8471 ( .A1(n6613), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U8472 ( .A1(n6613), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U8473 ( .A1(n6613), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U8474 ( .A1(n6613), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U8475 ( .A1(n6613), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U8476 ( .A1(n6613), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U8477 ( .A1(n6613), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U8478 ( .A1(n6613), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U8479 ( .A1(n6613), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U8480 ( .A1(n6613), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U8481 ( .A1(n6613), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U8482 ( .A1(n6613), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  INV_X1 U8483 ( .A(n6627), .ZN(n6630) );
  AOI22_X1 U8484 ( .A1(n7481), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n6628), .ZN(n6629) );
  OAI21_X1 U8485 ( .B1(n6630), .B2(n8960), .A(n6629), .ZN(P2_U3284) );
  INV_X1 U8486 ( .A(n9641), .ZN(n6918) );
  OAI222_X1 U8487 ( .A1(n9588), .A2(n6631), .B1(n9591), .B2(n6630), .C1(
        P1_U3086), .C2(n6918), .ZN(P1_U3344) );
  INV_X1 U8488 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6635) );
  AND2_X1 U8489 ( .A1(n5736), .A2(n7071), .ZN(n7932) );
  OR2_X1 U8490 ( .A1(n7932), .A2(n7060), .ZN(n7846) );
  OAI21_X1 U8491 ( .B1(n9734), .B2(n9746), .A(n7846), .ZN(n6632) );
  NAND2_X1 U8492 ( .A1(n5737), .A2(n9390), .ZN(n7009) );
  OAI211_X1 U8493 ( .C1(n6633), .C2(n7071), .A(n6632), .B(n7009), .ZN(n9525)
         );
  NAND2_X1 U8494 ( .A1(n9525), .A2(n9749), .ZN(n6634) );
  OAI21_X1 U8495 ( .B1(n9749), .B2(n6635), .A(n6634), .ZN(P1_U3453) );
  INV_X1 U8496 ( .A(n6636), .ZN(n6637) );
  AOI21_X1 U8497 ( .B1(n6639), .B2(n6638), .A(n6637), .ZN(n6642) );
  AOI22_X1 U8498 ( .A1(n9628), .A2(n7072), .B1(P1_REG3_REG_1__SCAN_IN), .B2(
        n6681), .ZN(n6641) );
  OR2_X1 U8499 ( .A1(n9095), .A2(n9412), .ZN(n9106) );
  INV_X1 U8500 ( .A(n9106), .ZN(n6682) );
  AOI22_X1 U8501 ( .A1(n6682), .A2(n5736), .B1(n9104), .B2(n9140), .ZN(n6640)
         );
  OAI211_X1 U8502 ( .C1(n6642), .C2(n9623), .A(n6641), .B(n6640), .ZN(P1_U3222) );
  NAND2_X1 U8503 ( .A1(n6382), .A2(n6645), .ZN(n8312) );
  INV_X1 U8504 ( .A(n8312), .ZN(n6643) );
  NOR2_X1 U8505 ( .A1(n8316), .A2(n6643), .ZN(n8470) );
  INV_X1 U8506 ( .A(n8470), .ZN(n6735) );
  OAI21_X1 U8507 ( .B1(n8759), .B2(n9853), .A(n6735), .ZN(n6644) );
  NAND2_X1 U8508 ( .A1(n6788), .A2(n8763), .ZN(n6999) );
  OAI211_X1 U8509 ( .C1(n6645), .C2(n9861), .A(n6644), .B(n6999), .ZN(n7023)
         );
  NAND2_X1 U8510 ( .A1(n7023), .A2(n9887), .ZN(n6646) );
  OAI21_X1 U8511 ( .B1(n9887), .B2(n6081), .A(n6646), .ZN(P2_U3459) );
  OAI21_X1 U8512 ( .B1(n6647), .B2(n6649), .A(n6648), .ZN(n6655) );
  INV_X1 U8513 ( .A(n9810), .ZN(n6654) );
  OAI21_X1 U8514 ( .B1(n6652), .B2(n6651), .A(n6650), .ZN(n6653) );
  AOI22_X1 U8515 ( .A1(n5992), .A2(n6655), .B1(n6654), .B2(n6653), .ZN(n6658)
         );
  INV_X1 U8516 ( .A(n5966), .ZN(n6656) );
  NAND2_X1 U8517 ( .A1(n9772), .A2(n6656), .ZN(n6657) );
  OAI211_X1 U8518 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n6092), .A(n6658), .B(n6657), .ZN(n6663) );
  AOI211_X1 U8519 ( .C1(n6661), .C2(n6660), .A(n8624), .B(n6659), .ZN(n6662)
         );
  AOI211_X1 U8520 ( .C1(n9796), .C2(P2_ADDR_REG_2__SCAN_IN), .A(n6663), .B(
        n6662), .ZN(n6664) );
  INV_X1 U8521 ( .A(n6664), .ZN(P2_U3184) );
  OAI21_X1 U8522 ( .B1(n6667), .B2(n6665), .A(n6666), .ZN(n7148) );
  AOI21_X1 U8523 ( .B1(n7070), .B2(n7142), .A(n9422), .ZN(n6668) );
  AND2_X1 U8524 ( .A1(n7094), .A2(n6668), .ZN(n7141) );
  XNOR2_X1 U8525 ( .A(n6665), .B(n6669), .ZN(n6671) );
  OAI222_X1 U8526 ( .A1(n9414), .A2(n5741), .B1(n6671), .B2(n9496), .C1(n9412), 
        .C2(n6670), .ZN(n7145) );
  AOI211_X1 U8527 ( .C1(n9734), .C2(n7148), .A(n7141), .B(n7145), .ZN(n6772)
         );
  AOI22_X1 U8528 ( .A1(n8073), .A2(n7142), .B1(n9754), .B2(
        P1_REG1_REG_2__SCAN_IN), .ZN(n6672) );
  OAI21_X1 U8529 ( .B1(n6772), .B2(n9754), .A(n6672), .ZN(P1_U3524) );
  INV_X1 U8530 ( .A(n6673), .ZN(n6687) );
  INV_X1 U8531 ( .A(n8014), .ZN(n6930) );
  INV_X1 U8532 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6674) );
  OAI222_X1 U8533 ( .A1(n9591), .A2(n6687), .B1(n6930), .B2(P1_U3086), .C1(
        n6674), .C2(n9588), .ZN(P1_U3343) );
  INV_X1 U8534 ( .A(n6675), .ZN(n6676) );
  NOR2_X1 U8535 ( .A1(n6677), .A2(n6676), .ZN(n6680) );
  INV_X1 U8536 ( .A(n6678), .ZN(n6679) );
  AOI21_X1 U8537 ( .B1(n6680), .B2(n6636), .A(n6679), .ZN(n6685) );
  AOI22_X1 U8538 ( .A1(n9628), .A2(n7142), .B1(P1_REG3_REG_2__SCAN_IN), .B2(
        n6681), .ZN(n6684) );
  AOI22_X1 U8539 ( .A1(n6682), .A2(n5737), .B1(n9104), .B2(n9139), .ZN(n6683)
         );
  OAI211_X1 U8540 ( .C1(n6685), .C2(n9623), .A(n6684), .B(n6683), .ZN(P1_U3237) );
  INV_X1 U8541 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6686) );
  OAI222_X1 U8542 ( .A1(P2_U3151), .A2(n6688), .B1(n8960), .B2(n6687), .C1(
        n6686), .C2(n8956), .ZN(P2_U3283) );
  INV_X1 U8543 ( .A(n6689), .ZN(n6715) );
  AOI22_X1 U8544 ( .A1(n9653), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n9585), .ZN(n6690) );
  OAI21_X1 U8545 ( .B1(n6715), .B2(n9591), .A(n6690), .ZN(P1_U3342) );
  NAND2_X1 U8546 ( .A1(P2_U3151), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n6827) );
  OAI211_X1 U8547 ( .C1(n4456), .C2(n6692), .A(n9807), .B(n6691), .ZN(n6693)
         );
  OAI211_X1 U8548 ( .C1(n9814), .C2(n6694), .A(n6827), .B(n6693), .ZN(n6704)
         );
  AOI21_X1 U8549 ( .B1(n6697), .B2(n6696), .A(n6695), .ZN(n6702) );
  AOI21_X1 U8550 ( .B1(n6700), .B2(n6699), .A(n6698), .ZN(n6701) );
  OAI22_X1 U8551 ( .A1(n6702), .A2(n9810), .B1(n9803), .B2(n6701), .ZN(n6703)
         );
  AOI211_X1 U8552 ( .C1(n9796), .C2(P2_ADDR_REG_4__SCAN_IN), .A(n6704), .B(
        n6703), .ZN(n6705) );
  INV_X1 U8553 ( .A(n6705), .ZN(P2_U3186) );
  OAI21_X1 U8554 ( .B1(n6708), .B2(n6707), .A(n6706), .ZN(n6712) );
  AOI22_X1 U8555 ( .A1(n9104), .A2(n9138), .B1(n9628), .B2(n7098), .ZN(n6710)
         );
  MUX2_X1 U8556 ( .A(n9631), .B(P1_STATE_REG_SCAN_IN), .S(
        P1_REG3_REG_3__SCAN_IN), .Z(n6709) );
  OAI211_X1 U8557 ( .C1(n7065), .C2(n9106), .A(n6710), .B(n6709), .ZN(n6711)
         );
  AOI21_X1 U8558 ( .B1(n6712), .B2(n9102), .A(n6711), .ZN(n6713) );
  INV_X1 U8559 ( .A(n6713), .ZN(P1_U3218) );
  INV_X1 U8560 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6714) );
  OAI222_X1 U8561 ( .A1(n6716), .A2(P2_U3151), .B1(n8960), .B2(n6715), .C1(
        n6714), .C2(n8956), .ZN(P2_U3282) );
  AND2_X1 U8562 ( .A1(n6706), .A2(n6717), .ZN(n6720) );
  OAI211_X1 U8563 ( .C1(n6720), .C2(n6719), .A(n9102), .B(n6718), .ZN(n6723)
         );
  AND2_X1 U8564 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n9187) );
  OAI22_X1 U8565 ( .A1(n7728), .A2(n8988), .B1(n9106), .B2(n5741), .ZN(n6721)
         );
  AOI211_X1 U8566 ( .C1(n7079), .C2(n9628), .A(n9187), .B(n6721), .ZN(n6722)
         );
  OAI211_X1 U8567 ( .C1(n9631), .C2(n6724), .A(n6723), .B(n6722), .ZN(P1_U3230) );
  AND2_X1 U8568 ( .A1(n6727), .A2(n6998), .ZN(n6796) );
  INV_X1 U8569 ( .A(n6796), .ZN(n6725) );
  NAND2_X1 U8570 ( .A1(n6727), .A2(n6726), .ZN(n6731) );
  INV_X1 U8571 ( .A(n6728), .ZN(n6729) );
  NAND2_X1 U8572 ( .A1(n6732), .A2(n6729), .ZN(n6730) );
  NAND2_X1 U8573 ( .A1(n6732), .A2(n9871), .ZN(n6734) );
  AOI22_X1 U8574 ( .A1(n8273), .A2(n6735), .B1(n7003), .B2(n8269), .ZN(n6751)
         );
  AND3_X1 U8575 ( .A1(n6738), .A2(n6737), .A3(n6736), .ZN(n6743) );
  INV_X1 U8576 ( .A(n6739), .ZN(n6740) );
  OR2_X1 U8577 ( .A1(n6741), .A2(n6740), .ZN(n6742) );
  OAI211_X1 U8578 ( .C1(n6747), .C2(n6744), .A(n6743), .B(n6742), .ZN(n6745)
         );
  NAND2_X1 U8579 ( .A1(n6745), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6749) );
  NAND2_X1 U8580 ( .A1(n6746), .A2(n6998), .ZN(n8515) );
  OR2_X1 U8581 ( .A1(n6747), .A2(n8515), .ZN(n6748) );
  NAND2_X1 U8582 ( .A1(n8267), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8232) );
  NAND2_X1 U8583 ( .A1(n8232), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n6750) );
  OAI211_X1 U8584 ( .C1(n6752), .C2(n8279), .A(n6751), .B(n6750), .ZN(P2_U3172) );
  AOI21_X1 U8585 ( .B1(n6755), .B2(n6754), .A(n6753), .ZN(n6768) );
  AOI21_X1 U8586 ( .B1(n4459), .B2(n6757), .A(n6756), .ZN(n6762) );
  AOI21_X1 U8587 ( .B1(n6760), .B2(n6759), .A(n6758), .ZN(n6761) );
  OAI22_X1 U8588 ( .A1(n6762), .A2(n9810), .B1(n6761), .B2(n9803), .ZN(n6763)
         );
  INV_X1 U8589 ( .A(n6763), .ZN(n6767) );
  NAND2_X1 U8590 ( .A1(P2_U3151), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n8250) );
  OAI21_X1 U8591 ( .B1(n9814), .B2(n6764), .A(n8250), .ZN(n6765) );
  AOI21_X1 U8592 ( .B1(n9796), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n6765), .ZN(
        n6766) );
  OAI211_X1 U8593 ( .C1(n6768), .C2(n8624), .A(n6767), .B(n6766), .ZN(P2_U3188) );
  INV_X1 U8594 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n6769) );
  OAI22_X1 U8595 ( .A1(n9576), .A2(n5738), .B1(n9749), .B2(n6769), .ZN(n6770)
         );
  INV_X1 U8596 ( .A(n6770), .ZN(n6771) );
  OAI21_X1 U8597 ( .B1(n6772), .B2(n9747), .A(n6771), .ZN(P1_U3459) );
  INV_X1 U8598 ( .A(n6773), .ZN(n6776) );
  AOI22_X1 U8599 ( .A1(n9665), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n9585), .ZN(n6774) );
  OAI21_X1 U8600 ( .B1(n6776), .B2(n9591), .A(n6774), .ZN(P1_U3341) );
  INV_X1 U8601 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6775) );
  OAI222_X1 U8602 ( .A1(P2_U3151), .A2(n6777), .B1(n8960), .B2(n6776), .C1(
        n6775), .C2(n8956), .ZN(P2_U3281) );
  INV_X1 U8603 ( .A(n6778), .ZN(n6815) );
  INV_X1 U8604 ( .A(n9678), .ZN(n8016) );
  INV_X1 U8605 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6779) );
  OAI222_X1 U8606 ( .A1(n9591), .A2(n6815), .B1(n8016), .B2(P1_U3086), .C1(
        n6779), .C2(n9588), .ZN(P1_U3340) );
  INV_X1 U8607 ( .A(n8316), .ZN(n6786) );
  INV_X1 U8608 ( .A(n6780), .ZN(n6782) );
  INV_X1 U8609 ( .A(n8466), .ZN(n6781) );
  NAND2_X1 U8610 ( .A1(n6782), .A2(n6781), .ZN(n6785) );
  NAND2_X1 U8611 ( .A1(n6786), .A2(n4955), .ZN(n6792) );
  INV_X1 U8612 ( .A(n6792), .ZN(n6794) );
  INV_X1 U8613 ( .A(n6789), .ZN(n6787) );
  NAND2_X1 U8614 ( .A1(n6789), .A2(n6752), .ZN(n6802) );
  INV_X1 U8615 ( .A(n6803), .ZN(n6793) );
  AOI21_X1 U8616 ( .B1(n6794), .B2(n6791), .A(n6793), .ZN(n6800) );
  AOI22_X1 U8617 ( .A1(n8277), .A2(n6382), .B1(n4461), .B2(n8269), .ZN(n6797)
         );
  OAI21_X1 U8618 ( .B1(n4861), .B2(n8279), .A(n6797), .ZN(n6798) );
  AOI21_X1 U8619 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(n8232), .A(n6798), .ZN(
        n6799) );
  OAI21_X1 U8620 ( .B1(n8271), .B2(n6800), .A(n6799), .ZN(P2_U3162) );
  NAND2_X1 U8621 ( .A1(n8621), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n6801) );
  OAI21_X1 U8622 ( .B1(n8689), .B2(n8621), .A(n6801), .ZN(P2_U3516) );
  XNOR2_X1 U8623 ( .A(n6817), .B(n8539), .ZN(n6809) );
  XNOR2_X1 U8624 ( .A(n6805), .B(n6102), .ZN(n8230) );
  NAND2_X1 U8625 ( .A1(n6805), .A2(n4861), .ZN(n6806) );
  NAND2_X1 U8626 ( .A1(n8229), .A2(n6806), .ZN(n6807) );
  INV_X1 U8627 ( .A(n6819), .ZN(n6808) );
  AOI211_X1 U8628 ( .C1(n6809), .C2(n6807), .A(n8271), .B(n6808), .ZN(n6813)
         );
  AOI22_X1 U8629 ( .A1(n8265), .A2(n8538), .B1(n8277), .B2(n6102), .ZN(n6811)
         );
  INV_X1 U8630 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n10011) );
  NOR2_X1 U8631 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10011), .ZN(n9771) );
  AOI21_X1 U8632 ( .B1(n8269), .B2(n9834), .A(n9771), .ZN(n6810) );
  OAI211_X1 U8633 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n8267), .A(n6811), .B(
        n6810), .ZN(n6812) );
  OR2_X1 U8634 ( .A1(n6813), .A2(n6812), .ZN(P2_U3158) );
  INV_X1 U8635 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6814) );
  OAI222_X1 U8636 ( .A1(P2_U3151), .A2(n6816), .B1(n8960), .B2(n6815), .C1(
        n6814), .C2(n8956), .ZN(P2_U3280) );
  NAND2_X1 U8637 ( .A1(n6817), .A2(n8539), .ZN(n6818) );
  XNOR2_X1 U8638 ( .A(n8129), .B(n6943), .ZN(n6821) );
  INV_X1 U8639 ( .A(n8538), .ZN(n6820) );
  NAND2_X1 U8640 ( .A1(n6821), .A2(n6820), .ZN(n6897) );
  INV_X1 U8641 ( .A(n6821), .ZN(n6822) );
  NAND2_X1 U8642 ( .A1(n6822), .A2(n8538), .ZN(n6823) );
  AND2_X1 U8643 ( .A1(n6897), .A2(n6823), .ZN(n6826) );
  OAI21_X1 U8644 ( .B1(n6824), .B2(n6826), .A(n6825), .ZN(n6832) );
  AOI22_X1 U8645 ( .A1(n8265), .A2(n8537), .B1(n8277), .B2(n8539), .ZN(n6830)
         );
  INV_X1 U8646 ( .A(n6827), .ZN(n6828) );
  AOI21_X1 U8647 ( .B1(n8269), .B2(n6943), .A(n6828), .ZN(n6829) );
  OAI211_X1 U8648 ( .C1(n6941), .C2(n8267), .A(n6830), .B(n6829), .ZN(n6831)
         );
  AOI21_X1 U8649 ( .B1(n6832), .B2(n8273), .A(n6831), .ZN(n6833) );
  INV_X1 U8650 ( .A(n6833), .ZN(P2_U3170) );
  OAI21_X1 U8651 ( .B1(n6834), .B2(n4669), .A(n6876), .ZN(n6840) );
  INV_X1 U8652 ( .A(n6382), .ZN(n6835) );
  OAI22_X1 U8653 ( .A1(n6835), .A2(n8790), .B1(n4861), .B2(n8788), .ZN(n6839)
         );
  INV_X1 U8654 ( .A(n6836), .ZN(n6837) );
  AOI21_X1 U8655 ( .B1(n6786), .B2(n4669), .A(n6837), .ZN(n6856) );
  NOR2_X1 U8656 ( .A1(n6856), .A2(n6936), .ZN(n6838) );
  AOI211_X1 U8657 ( .C1(n8759), .C2(n6840), .A(n6839), .B(n6838), .ZN(n6852)
         );
  INV_X1 U8658 ( .A(n6856), .ZN(n6842) );
  INV_X1 U8659 ( .A(n9828), .ZN(n6841) );
  AOI22_X1 U8660 ( .A1(n6842), .A2(n6841), .B1(n9871), .B2(n4461), .ZN(n6843)
         );
  NAND2_X1 U8661 ( .A1(n6852), .A2(n6843), .ZN(n7028) );
  NAND2_X1 U8662 ( .A1(n7028), .A2(n9887), .ZN(n6844) );
  OAI21_X1 U8663 ( .B1(n9887), .B2(n6845), .A(n6844), .ZN(P2_U3460) );
  MUX2_X1 U8664 ( .A(n6782), .B(n6848), .S(n6847), .Z(n6850) );
  NOR2_X1 U8665 ( .A1(n6851), .A2(n8315), .ZN(n6935) );
  NAND2_X1 U8666 ( .A1(n9824), .A2(n6935), .ZN(n7704) );
  MUX2_X1 U8667 ( .A(n6480), .B(n6852), .S(n9824), .Z(n6855) );
  NOR2_X2 U8668 ( .A1(n6853), .A2(n8686), .ZN(n9819) );
  AOI22_X1 U8669 ( .A1(n9819), .A2(n4461), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n9821), .ZN(n6854) );
  OAI211_X1 U8670 ( .C1(n6856), .C2(n7704), .A(n6855), .B(n6854), .ZN(P2_U3232) );
  XNOR2_X1 U8671 ( .A(n6857), .B(n6859), .ZN(n7172) );
  OAI21_X1 U8672 ( .B1(n6860), .B2(n6859), .A(n6858), .ZN(n7163) );
  AOI21_X1 U8673 ( .B1(n6965), .B2(n7727), .A(n9422), .ZN(n6861) );
  AND2_X1 U8674 ( .A1(n6861), .A2(n7181), .ZN(n7169) );
  OR2_X1 U8675 ( .A1(n7090), .A2(n9412), .ZN(n6863) );
  OR2_X1 U8676 ( .A1(n7722), .A2(n9414), .ZN(n6862) );
  NAND2_X1 U8677 ( .A1(n6863), .A2(n6862), .ZN(n7165) );
  AOI211_X1 U8678 ( .C1(n7163), .C2(n9734), .A(n7169), .B(n7165), .ZN(n6864)
         );
  OAI21_X1 U8679 ( .B1(n9496), .B2(n7172), .A(n6864), .ZN(n6870) );
  INV_X1 U8680 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6865) );
  OAI22_X1 U8681 ( .A1(n9524), .A2(n5744), .B1(n9757), .B2(n6865), .ZN(n6866)
         );
  AOI21_X1 U8682 ( .B1(n6870), .B2(n9757), .A(n6866), .ZN(n6867) );
  INV_X1 U8683 ( .A(n6867), .ZN(P1_U3527) );
  INV_X1 U8684 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n6868) );
  OAI22_X1 U8685 ( .A1(n9576), .A2(n5744), .B1(n9749), .B2(n6868), .ZN(n6869)
         );
  AOI21_X1 U8686 ( .B1(n6870), .B2(n9749), .A(n6869), .ZN(n6871) );
  INV_X1 U8687 ( .A(n6871), .ZN(P1_U3468) );
  OR2_X1 U8688 ( .A1(n6872), .A2(n8467), .ZN(n6873) );
  NAND2_X1 U8689 ( .A1(n6874), .A2(n6873), .ZN(n6880) );
  INV_X1 U8690 ( .A(n6880), .ZN(n9829) );
  NAND3_X1 U8691 ( .A1(n6876), .A2(n8467), .A3(n6875), .ZN(n6877) );
  AND2_X1 U8692 ( .A1(n6878), .A2(n6877), .ZN(n6883) );
  INV_X1 U8693 ( .A(n6936), .ZN(n6879) );
  NAND2_X1 U8694 ( .A1(n6880), .A2(n6879), .ZN(n6882) );
  AOI22_X1 U8695 ( .A1(n8745), .A2(n6788), .B1(n8539), .B2(n8763), .ZN(n6881)
         );
  OAI211_X1 U8696 ( .C1(n8786), .C2(n6883), .A(n6882), .B(n6881), .ZN(n9831)
         );
  OAI22_X1 U8697 ( .A1(n8679), .A2(n6092), .B1(n9827), .B2(n8686), .ZN(n6884)
         );
  NOR2_X1 U8698 ( .A1(n9831), .A2(n6884), .ZN(n6885) );
  INV_X2 U8699 ( .A(n9824), .ZN(n8803) );
  MUX2_X1 U8700 ( .A(n6885), .B(n5906), .S(n8803), .Z(n6886) );
  OAI21_X1 U8701 ( .B1(n9829), .B2(n7704), .A(n6886), .ZN(P2_U3231) );
  NAND2_X1 U8702 ( .A1(n6888), .A2(n6887), .ZN(n6889) );
  XOR2_X1 U8703 ( .A(n6890), .B(n6889), .Z(n6893) );
  AOI22_X1 U8704 ( .A1(n9628), .A2(n7727), .B1(P1_REG3_REG_5__SCAN_IN), .B2(
        P1_U3086), .ZN(n6892) );
  INV_X1 U8705 ( .A(n9095), .ZN(n9618) );
  AOI22_X1 U8706 ( .A1(n7164), .A2(n9109), .B1(n7165), .B2(n9618), .ZN(n6891)
         );
  OAI211_X1 U8707 ( .C1(n6893), .C2(n9623), .A(n6892), .B(n6891), .ZN(P1_U3227) );
  NAND2_X1 U8708 ( .A1(n6894), .A2(n6897), .ZN(n6895) );
  XNOR2_X1 U8709 ( .A(n8129), .B(n9845), .ZN(n7236) );
  XNOR2_X1 U8710 ( .A(n7236), .B(n8537), .ZN(n6896) );
  INV_X1 U8711 ( .A(n6896), .ZN(n6898) );
  NAND3_X1 U8712 ( .A1(n6825), .A2(n6898), .A3(n6897), .ZN(n6899) );
  AOI21_X1 U8713 ( .B1(n7238), .B2(n6899), .A(n8271), .ZN(n6904) );
  AOI22_X1 U8714 ( .A1(n8265), .A2(n8536), .B1(n8277), .B2(n8538), .ZN(n6902)
         );
  NAND2_X1 U8715 ( .A1(P2_U3151), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n9793) );
  INV_X1 U8716 ( .A(n9793), .ZN(n6900) );
  AOI21_X1 U8717 ( .B1(n8269), .B2(n9845), .A(n6900), .ZN(n6901) );
  OAI211_X1 U8718 ( .C1(n7036), .C2(n8267), .A(n6902), .B(n6901), .ZN(n6903)
         );
  OR2_X1 U8719 ( .A1(n6904), .A2(n6903), .ZN(P2_U3167) );
  NAND2_X1 U8720 ( .A1(n6906), .A2(n6905), .ZN(n6908) );
  XOR2_X1 U8721 ( .A(n6908), .B(n6907), .Z(n6913) );
  AOI22_X1 U8722 ( .A1(n9104), .A2(n9135), .B1(P1_REG3_REG_6__SCAN_IN), .B2(
        P1_U3086), .ZN(n6910) );
  NAND2_X1 U8723 ( .A1(n9109), .A2(n7188), .ZN(n6909) );
  OAI211_X1 U8724 ( .C1(n7728), .C2(n9106), .A(n6910), .B(n6909), .ZN(n6911)
         );
  AOI21_X1 U8725 ( .B1(n7723), .B2(n9628), .A(n6911), .ZN(n6912) );
  OAI21_X1 U8726 ( .B1(n6913), .B2(n9623), .A(n6912), .ZN(P1_U3239) );
  NOR2_X1 U8727 ( .A1(n8014), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n6914) );
  AOI21_X1 U8728 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n8014), .A(n6914), .ZN(
        n6921) );
  INV_X1 U8729 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7334) );
  AOI22_X1 U8730 ( .A1(n9601), .A2(n7334), .B1(P1_REG2_REG_10__SCAN_IN), .B2(
        n6915), .ZN(n9594) );
  NOR2_X1 U8731 ( .A1(n9611), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6917) );
  AOI21_X1 U8732 ( .B1(n9611), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6917), .ZN(
        n9606) );
  NAND2_X1 U8733 ( .A1(n9605), .A2(n9606), .ZN(n9604) );
  OAI21_X1 U8734 ( .B1(n9611), .B2(P1_REG2_REG_9__SCAN_IN), .A(n9604), .ZN(
        n9595) );
  NOR2_X1 U8735 ( .A1(n9594), .A2(n9595), .ZN(n9593) );
  INV_X1 U8736 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n6919) );
  AOI22_X1 U8737 ( .A1(n9641), .A2(n6919), .B1(P1_REG2_REG_11__SCAN_IN), .B2(
        n6918), .ZN(n9634) );
  NOR2_X1 U8738 ( .A1(n9635), .A2(n9634), .ZN(n9633) );
  AOI21_X1 U8739 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n9641), .A(n9633), .ZN(
        n6920) );
  NAND2_X1 U8740 ( .A1(n6921), .A2(n6920), .ZN(n8002) );
  OAI21_X1 U8741 ( .B1(n6921), .B2(n6920), .A(n8002), .ZN(n6922) );
  INV_X1 U8742 ( .A(n6922), .ZN(n6934) );
  INV_X1 U8743 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6923) );
  MUX2_X1 U8744 ( .A(n6923), .B(P1_REG1_REG_10__SCAN_IN), .S(n9601), .Z(n9597)
         );
  AOI21_X1 U8745 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(n6925), .A(n6924), .ZN(
        n9608) );
  NOR2_X1 U8746 ( .A1(n9611), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6926) );
  AOI21_X1 U8747 ( .B1(n9611), .B2(P1_REG1_REG_9__SCAN_IN), .A(n6926), .ZN(
        n9609) );
  NAND2_X1 U8748 ( .A1(n9608), .A2(n9609), .ZN(n9607) );
  OAI21_X1 U8749 ( .B1(n9611), .B2(P1_REG1_REG_9__SCAN_IN), .A(n9607), .ZN(
        n9598) );
  NOR2_X1 U8750 ( .A1(n9597), .A2(n9598), .ZN(n9596) );
  AOI21_X1 U8751 ( .B1(n9601), .B2(P1_REG1_REG_10__SCAN_IN), .A(n9596), .ZN(
        n9638) );
  XNOR2_X1 U8752 ( .A(n9641), .B(P1_REG1_REG_11__SCAN_IN), .ZN(n9637) );
  NOR2_X1 U8753 ( .A1(n9638), .A2(n9637), .ZN(n9636) );
  AOI21_X1 U8754 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(n9641), .A(n9636), .ZN(
        n6928) );
  INV_X1 U8755 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n7552) );
  AOI22_X1 U8756 ( .A1(n8014), .A2(P1_REG1_REG_12__SCAN_IN), .B1(n7552), .B2(
        n6930), .ZN(n6927) );
  NAND2_X1 U8757 ( .A1(n6928), .A2(n6927), .ZN(n8013) );
  OAI21_X1 U8758 ( .B1(n6928), .B2(n6927), .A(n8013), .ZN(n6932) );
  NAND2_X1 U8759 ( .A1(n9188), .A2(P1_ADDR_REG_12__SCAN_IN), .ZN(n6929) );
  NAND2_X1 U8760 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7625) );
  OAI211_X1 U8761 ( .C1(n6930), .C2(n9718), .A(n6929), .B(n7625), .ZN(n6931)
         );
  AOI21_X1 U8762 ( .B1(n6932), .B2(n9712), .A(n6931), .ZN(n6933) );
  OAI21_X1 U8763 ( .B1(n6934), .B2(n9686), .A(n6933), .ZN(P1_U3255) );
  INV_X1 U8764 ( .A(n6935), .ZN(n6937) );
  NAND2_X1 U8765 ( .A1(n6937), .A2(n6936), .ZN(n9815) );
  XNOR2_X1 U8766 ( .A(n6938), .B(n8471), .ZN(n9839) );
  XNOR2_X1 U8767 ( .A(n6939), .B(n8471), .ZN(n6940) );
  AOI222_X1 U8768 ( .A1(n8759), .A2(n6940), .B1(n8537), .B2(n8763), .C1(n8539), 
        .C2(n8745), .ZN(n9840) );
  MUX2_X1 U8769 ( .A(n5913), .B(n9840), .S(n9824), .Z(n6945) );
  INV_X1 U8770 ( .A(n6941), .ZN(n6942) );
  AOI22_X1 U8771 ( .A1(n9819), .A2(n6943), .B1(n9821), .B2(n6942), .ZN(n6944)
         );
  OAI211_X1 U8772 ( .C1(n8673), .C2(n9839), .A(n6945), .B(n6944), .ZN(P2_U3229) );
  AOI21_X1 U8773 ( .B1(n6133), .B2(n6947), .A(n6946), .ZN(n6959) );
  XNOR2_X1 U8774 ( .A(n6949), .B(n6948), .ZN(n6957) );
  NAND2_X1 U8775 ( .A1(n9796), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n6950) );
  NAND2_X1 U8776 ( .A1(P2_U3151), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7391) );
  OAI211_X1 U8777 ( .C1(n9814), .C2(n6951), .A(n6950), .B(n7391), .ZN(n6956)
         );
  AOI21_X1 U8778 ( .B1(n9826), .B2(n6953), .A(n6952), .ZN(n6954) );
  NOR2_X1 U8779 ( .A1(n6954), .A2(n9810), .ZN(n6955) );
  AOI211_X1 U8780 ( .C1(n9807), .C2(n6957), .A(n6956), .B(n6955), .ZN(n6958)
         );
  OAI21_X1 U8781 ( .B1(n6959), .B2(n9803), .A(n6958), .ZN(P2_U3189) );
  OAI21_X1 U8782 ( .B1(n6960), .B2(n7847), .A(n6961), .ZN(n7084) );
  INV_X1 U8783 ( .A(n7084), .ZN(n6966) );
  NAND3_X1 U8784 ( .A1(n7087), .A2(n7937), .A3(n7847), .ZN(n6962) );
  NAND2_X1 U8785 ( .A1(n6963), .A2(n6962), .ZN(n6964) );
  AOI222_X1 U8786 ( .A1(n9746), .A2(n6964), .B1(n9137), .B2(n9390), .C1(n9139), 
        .C2(n9393), .ZN(n7086) );
  OAI211_X1 U8787 ( .C1(n7095), .C2(n6971), .A(n6965), .B(n9477), .ZN(n7082)
         );
  OAI211_X1 U8788 ( .C1(n9516), .C2(n6966), .A(n7086), .B(n7082), .ZN(n6973)
         );
  INV_X1 U8789 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6967) );
  OAI22_X1 U8790 ( .A1(n9524), .A2(n6971), .B1(n9757), .B2(n6967), .ZN(n6968)
         );
  AOI21_X1 U8791 ( .B1(n6973), .B2(n9757), .A(n6968), .ZN(n6969) );
  INV_X1 U8792 ( .A(n6969), .ZN(P1_U3526) );
  INV_X1 U8793 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n6970) );
  OAI22_X1 U8794 ( .A1(n9576), .A2(n6971), .B1(n9749), .B2(n6970), .ZN(n6972)
         );
  AOI21_X1 U8795 ( .B1(n6973), .B2(n9749), .A(n6972), .ZN(n6974) );
  INV_X1 U8796 ( .A(n6974), .ZN(P1_U3465) );
  XNOR2_X1 U8797 ( .A(n6976), .B(n6975), .ZN(n6977) );
  XNOR2_X1 U8798 ( .A(n6978), .B(n6977), .ZN(n6986) );
  NOR2_X1 U8799 ( .A1(n9113), .A2(n9739), .ZN(n6984) );
  OR2_X1 U8800 ( .A1(n7722), .A2(n9412), .ZN(n6980) );
  OR2_X1 U8801 ( .A1(n7385), .A2(n9414), .ZN(n6979) );
  NAND2_X1 U8802 ( .A1(n6980), .A2(n6979), .ZN(n7112) );
  NAND2_X1 U8803 ( .A1(n7112), .A2(n9618), .ZN(n6981) );
  OAI21_X1 U8804 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n6982), .A(n6981), .ZN(n6983) );
  AOI211_X1 U8805 ( .C1(n9109), .C2(n7113), .A(n6984), .B(n6983), .ZN(n6985)
         );
  OAI21_X1 U8806 ( .B1(n6986), .B2(n9623), .A(n6985), .ZN(P1_U3213) );
  XNOR2_X1 U8807 ( .A(n6988), .B(n6987), .ZN(n6989) );
  NAND2_X1 U8808 ( .A1(n6989), .A2(n8759), .ZN(n6991) );
  AOI22_X1 U8809 ( .A1(n8745), .A2(n6102), .B1(n8538), .B2(n8763), .ZN(n6990)
         );
  AND2_X1 U8810 ( .A1(n6991), .A2(n6990), .ZN(n9836) );
  XNOR2_X1 U8811 ( .A(n8469), .B(n6992), .ZN(n9833) );
  NOR2_X1 U8812 ( .A1(n9824), .A2(n6104), .ZN(n6995) );
  OAI22_X1 U8813 ( .A1(n8798), .A2(n6993), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n8679), .ZN(n6994) );
  AOI211_X1 U8814 ( .C1(n9833), .C2(n8801), .A(n6995), .B(n6994), .ZN(n6996)
         );
  OAI21_X1 U8815 ( .B1(n8803), .B2(n9836), .A(n6996), .ZN(P2_U3230) );
  NAND2_X1 U8816 ( .A1(n9141), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n6997) );
  OAI21_X1 U8817 ( .B1(n7812), .B2(n9141), .A(n6997), .ZN(P1_U3583) );
  OR3_X1 U8818 ( .A1(n8470), .A2(n9871), .A3(n6998), .ZN(n7000) );
  OAI211_X1 U8819 ( .C1(n8679), .C2(n10111), .A(n7000), .B(n6999), .ZN(n7001)
         );
  MUX2_X1 U8820 ( .A(n7001), .B(P2_REG2_REG_0__SCAN_IN), .S(n8803), .Z(n7002)
         );
  AOI21_X1 U8821 ( .B1(n9819), .B2(n7003), .A(n7002), .ZN(n7004) );
  INV_X1 U8822 ( .A(n7004), .ZN(P2_U3233) );
  NAND2_X1 U8823 ( .A1(n7006), .A2(n7005), .ZN(n7007) );
  INV_X1 U8824 ( .A(n7008), .ZN(n7011) );
  INV_X1 U8825 ( .A(n7009), .ZN(n7010) );
  AOI21_X1 U8826 ( .B1(n7846), .B2(n7011), .A(n7010), .ZN(n7016) );
  NOR2_X1 U8827 ( .A1(n9360), .A2(n9422), .ZN(n9326) );
  NOR2_X2 U8828 ( .A1(n9433), .A2(n7012), .ZN(n9364) );
  OAI21_X1 U8829 ( .B1(n9326), .B2(n9364), .A(n7013), .ZN(n7015) );
  INV_X2 U8830 ( .A(n7333), .ZN(n9426) );
  AOI22_X1 U8831 ( .A1(n9211), .A2(P1_REG2_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(n9426), .ZN(n7014) );
  OAI211_X1 U8832 ( .C1(n9211), .C2(n7016), .A(n7015), .B(n7014), .ZN(P1_U3293) );
  INV_X1 U8833 ( .A(n7017), .ZN(n7020) );
  INV_X1 U8834 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7018) );
  OAI222_X1 U8835 ( .A1(n7019), .A2(P2_U3151), .B1(n8960), .B2(n7020), .C1(
        n7018), .C2(n8956), .ZN(P2_U3279) );
  INV_X1 U8836 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n7021) );
  INV_X1 U8837 ( .A(n8012), .ZN(n9685) );
  OAI222_X1 U8838 ( .A1(n9588), .A2(n7021), .B1(n9591), .B2(n7020), .C1(
        P1_U3086), .C2(n9685), .ZN(P1_U3339) );
  NAND2_X1 U8839 ( .A1(n8621), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n7022) );
  OAI21_X1 U8840 ( .B1(n8638), .B2(n8621), .A(n7022), .ZN(P2_U3520) );
  INV_X1 U8841 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n7025) );
  NAND2_X1 U8842 ( .A1(n7023), .A2(n8939), .ZN(n7024) );
  OAI21_X1 U8843 ( .B1(n8939), .B2(n7025), .A(n7024), .ZN(P2_U3390) );
  INV_X1 U8844 ( .A(n7026), .ZN(n7059) );
  AOI22_X1 U8845 ( .A1(n9700), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n9585), .ZN(n7027) );
  OAI21_X1 U8846 ( .B1(n7059), .B2(n9591), .A(n7027), .ZN(P1_U3338) );
  INV_X1 U8847 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n7030) );
  NAND2_X1 U8848 ( .A1(n7028), .A2(n8939), .ZN(n7029) );
  OAI21_X1 U8849 ( .B1(n7030), .B2(n8939), .A(n7029), .ZN(P2_U3393) );
  OAI21_X1 U8850 ( .B1(n7032), .B2(n7033), .A(n7031), .ZN(n9846) );
  INV_X1 U8851 ( .A(n9846), .ZN(n7040) );
  XNOR2_X1 U8852 ( .A(n7034), .B(n7033), .ZN(n7035) );
  AOI222_X1 U8853 ( .A1(n8759), .A2(n7035), .B1(n8536), .B2(n8763), .C1(n8538), 
        .C2(n8745), .ZN(n9848) );
  MUX2_X1 U8854 ( .A(n9786), .B(n9848), .S(n9824), .Z(n7039) );
  INV_X1 U8855 ( .A(n7036), .ZN(n7037) );
  AOI22_X1 U8856 ( .A1(n9819), .A2(n9845), .B1(n9821), .B2(n7037), .ZN(n7038)
         );
  OAI211_X1 U8857 ( .C1(n8673), .C2(n7040), .A(n7039), .B(n7038), .ZN(P2_U3228) );
  AOI21_X1 U8858 ( .B1(n7043), .B2(n7042), .A(n7041), .ZN(n7057) );
  OAI21_X1 U8859 ( .B1(n7046), .B2(n7045), .A(n7044), .ZN(n7055) );
  NAND2_X1 U8860 ( .A1(n9796), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n7047) );
  NAND2_X1 U8861 ( .A1(P2_U3151), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n7255) );
  OAI211_X1 U8862 ( .C1(n9814), .C2(n7048), .A(n7047), .B(n7255), .ZN(n7054)
         );
  AOI21_X1 U8863 ( .B1(n7051), .B2(n7050), .A(n7049), .ZN(n7052) );
  NOR2_X1 U8864 ( .A1(n7052), .A2(n9810), .ZN(n7053) );
  AOI211_X1 U8865 ( .C1(n9807), .C2(n7055), .A(n7054), .B(n7053), .ZN(n7056)
         );
  OAI21_X1 U8866 ( .B1(n7057), .B2(n9803), .A(n7056), .ZN(P2_U3190) );
  INV_X1 U8867 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7058) );
  OAI222_X1 U8868 ( .A1(P2_U3151), .A2(n9813), .B1(n8960), .B2(n7059), .C1(
        n7058), .C2(n8956), .ZN(P2_U3278) );
  INV_X1 U8869 ( .A(n5736), .ZN(n7064) );
  INV_X1 U8870 ( .A(n7060), .ZN(n7062) );
  AOI21_X1 U8871 ( .B1(n7852), .B2(n7062), .A(n7061), .ZN(n7063) );
  OAI222_X1 U8872 ( .A1(n9414), .A2(n7065), .B1(n9412), .B2(n7064), .C1(n9496), 
        .C2(n7063), .ZN(n9726) );
  INV_X1 U8873 ( .A(n9726), .ZN(n7077) );
  NAND2_X1 U8874 ( .A1(n7875), .A2(n7066), .ZN(n9406) );
  OAI21_X1 U8875 ( .B1(n7852), .B2(n7069), .A(n7068), .ZN(n9728) );
  OAI211_X1 U8876 ( .C1(n7071), .C2(n5821), .A(n9477), .B(n7070), .ZN(n9725)
         );
  NAND2_X1 U8877 ( .A1(n9364), .A2(n7072), .ZN(n7074) );
  AOI22_X1 U8878 ( .A1(n9426), .A2(P1_REG3_REG_1__SCAN_IN), .B1(
        P1_REG2_REG_1__SCAN_IN), .B2(n9211), .ZN(n7073) );
  OAI211_X1 U8879 ( .C1(n9360), .C2(n9725), .A(n7074), .B(n7073), .ZN(n7075)
         );
  AOI21_X1 U8880 ( .B1(n9355), .B2(n9728), .A(n7075), .ZN(n7076) );
  OAI21_X1 U8881 ( .B1(n7077), .B2(n9433), .A(n7076), .ZN(P1_U3292) );
  AOI22_X1 U8882 ( .A1(n9433), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n7078), .B2(
        n9426), .ZN(n7081) );
  NAND2_X1 U8883 ( .A1(n9364), .A2(n7079), .ZN(n7080) );
  OAI211_X1 U8884 ( .C1(n7082), .C2(n9360), .A(n7081), .B(n7080), .ZN(n7083)
         );
  AOI21_X1 U8885 ( .B1(n7084), .B2(n9355), .A(n7083), .ZN(n7085) );
  OAI21_X1 U8886 ( .B1(n7086), .B2(n9433), .A(n7085), .ZN(P1_U3289) );
  INV_X1 U8887 ( .A(n7087), .ZN(n7088) );
  AOI21_X1 U8888 ( .B1(n7707), .B2(n7092), .A(n7088), .ZN(n7089) );
  OAI222_X1 U8889 ( .A1(n9414), .A2(n7090), .B1(n9412), .B2(n7065), .C1(n9496), 
        .C2(n7089), .ZN(n9731) );
  INV_X1 U8890 ( .A(n9731), .ZN(n7103) );
  OAI21_X1 U8891 ( .B1(n7093), .B2(n7092), .A(n7091), .ZN(n9733) );
  INV_X1 U8892 ( .A(n7095), .ZN(n7096) );
  OAI211_X1 U8893 ( .C1(n5740), .C2(n4578), .A(n7096), .B(n9477), .ZN(n9730)
         );
  AOI22_X1 U8894 ( .A1(n9211), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n9426), .B2(
        n7097), .ZN(n7100) );
  NAND2_X1 U8895 ( .A1(n9364), .A2(n7098), .ZN(n7099) );
  OAI211_X1 U8896 ( .C1(n9730), .C2(n9360), .A(n7100), .B(n7099), .ZN(n7101)
         );
  AOI21_X1 U8897 ( .B1(n9733), .B2(n9355), .A(n7101), .ZN(n7102) );
  OAI21_X1 U8898 ( .B1(n7103), .B2(n9433), .A(n7102), .ZN(P1_U3290) );
  OAI21_X1 U8899 ( .B1(n7105), .B2(n7108), .A(n7104), .ZN(n7106) );
  INV_X1 U8900 ( .A(n7106), .ZN(n9740) );
  AOI21_X1 U8901 ( .B1(n7177), .B2(n7729), .A(n7107), .ZN(n7109) );
  INV_X1 U8902 ( .A(n7109), .ZN(n7110) );
  INV_X1 U8903 ( .A(n7108), .ZN(n7733) );
  NOR2_X1 U8904 ( .A1(n7109), .A2(n7108), .ZN(n7151) );
  INV_X1 U8905 ( .A(n7151), .ZN(n7215) );
  OAI21_X1 U8906 ( .B1(n7110), .B2(n7733), .A(n7215), .ZN(n9745) );
  NAND2_X1 U8907 ( .A1(n9381), .A2(n9746), .ZN(n9367) );
  INV_X1 U8908 ( .A(n9367), .ZN(n8088) );
  OAI21_X1 U8909 ( .B1(n7180), .B2(n9739), .A(n9477), .ZN(n7111) );
  OR2_X1 U8910 ( .A1(n7111), .A2(n7210), .ZN(n9737) );
  INV_X1 U8911 ( .A(n7112), .ZN(n9736) );
  AOI22_X1 U8912 ( .A1(n9211), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n7113), .B2(
        n9426), .ZN(n7114) );
  OAI21_X1 U8913 ( .B1(n9736), .B2(n9433), .A(n7114), .ZN(n7115) );
  AOI21_X1 U8914 ( .B1(n9364), .B2(n7116), .A(n7115), .ZN(n7117) );
  OAI21_X1 U8915 ( .B1(n9737), .B2(n9360), .A(n7117), .ZN(n7118) );
  AOI21_X1 U8916 ( .B1(n9745), .B2(n8088), .A(n7118), .ZN(n7119) );
  OAI21_X1 U8917 ( .B1(n9740), .B2(n9404), .A(n7119), .ZN(P1_U3286) );
  INV_X1 U8918 ( .A(n7120), .ZN(n7139) );
  AOI22_X1 U8919 ( .A1(n9706), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n9585), .ZN(n7121) );
  OAI21_X1 U8920 ( .B1(n7139), .B2(n9591), .A(n7121), .ZN(P1_U3337) );
  XNOR2_X1 U8921 ( .A(n7122), .B(n8476), .ZN(n9856) );
  OR2_X1 U8922 ( .A1(n7123), .A2(n7124), .ZN(n7126) );
  NAND2_X1 U8923 ( .A1(n7126), .A2(n7125), .ZN(n7130) );
  OR2_X1 U8924 ( .A1(n7123), .A2(n7127), .ZN(n7200) );
  AND2_X1 U8925 ( .A1(n7200), .A2(n7197), .ZN(n7128) );
  OAI211_X1 U8926 ( .C1(n7130), .C2(n7129), .A(n7128), .B(n8759), .ZN(n7132)
         );
  AOI22_X1 U8927 ( .A1(n8533), .A2(n8763), .B1(n8745), .B2(n8535), .ZN(n7131)
         );
  NAND2_X1 U8928 ( .A1(n7132), .A2(n7131), .ZN(n9857) );
  NAND2_X1 U8929 ( .A1(n9857), .A2(n9824), .ZN(n7137) );
  OAI22_X1 U8930 ( .A1(n9824), .A2(n7134), .B1(n7133), .B2(n8679), .ZN(n7135)
         );
  AOI21_X1 U8931 ( .B1(n9819), .B2(n9859), .A(n7135), .ZN(n7136) );
  OAI211_X1 U8932 ( .C1(n9856), .C2(n8673), .A(n7137), .B(n7136), .ZN(P2_U3225) );
  INV_X1 U8933 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7140) );
  OAI222_X1 U8934 ( .A1(n8956), .A2(n7140), .B1(n8960), .B2(n7139), .C1(
        P2_U3151), .C2(n7138), .ZN(P2_U3277) );
  INV_X1 U8935 ( .A(n7141), .ZN(n7144) );
  AOI22_X1 U8936 ( .A1(n9364), .A2(n7142), .B1(n9426), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n7143) );
  OAI21_X1 U8937 ( .B1(n9360), .B2(n7144), .A(n7143), .ZN(n7147) );
  MUX2_X1 U8938 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n7145), .S(n9381), .Z(n7146)
         );
  AOI211_X1 U8939 ( .C1(n9355), .C2(n7148), .A(n7147), .B(n7146), .ZN(n7149)
         );
  INV_X1 U8940 ( .A(n7149), .ZN(P1_U3291) );
  OAI21_X1 U8941 ( .B1(n7151), .B2(n7734), .A(n7150), .ZN(n7152) );
  XOR2_X1 U8942 ( .A(n7159), .B(n7152), .Z(n7273) );
  OR2_X1 U8943 ( .A1(n7385), .A2(n9412), .ZN(n7271) );
  AOI22_X1 U8944 ( .A1(n9211), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n7387), .B2(
        n9426), .ZN(n7153) );
  OAI21_X1 U8945 ( .B1(n7271), .B2(n9433), .A(n7153), .ZN(n7156) );
  AOI21_X1 U8946 ( .B1(n7211), .B2(n7157), .A(n9422), .ZN(n7154) );
  AOI22_X1 U8947 ( .A1(n7154), .A2(n7332), .B1(n9390), .B2(n9132), .ZN(n7272)
         );
  NOR2_X1 U8948 ( .A1(n7272), .A2(n9360), .ZN(n7155) );
  AOI211_X1 U8949 ( .C1(n9364), .C2(n7157), .A(n7156), .B(n7155), .ZN(n7162)
         );
  OAI21_X1 U8950 ( .B1(n7160), .B2(n7159), .A(n7158), .ZN(n7275) );
  NAND2_X1 U8951 ( .A1(n7275), .A2(n9355), .ZN(n7161) );
  OAI211_X1 U8952 ( .C1(n7273), .C2(n9367), .A(n7162), .B(n7161), .ZN(P1_U3284) );
  NAND2_X1 U8953 ( .A1(n7163), .A2(n9355), .ZN(n7171) );
  AOI22_X1 U8954 ( .A1(n9433), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n7164), .B2(
        n9426), .ZN(n7167) );
  NAND2_X1 U8955 ( .A1(n7165), .A2(n9381), .ZN(n7166) );
  OAI211_X1 U8956 ( .C1(n9429), .C2(n5744), .A(n7167), .B(n7166), .ZN(n7168)
         );
  AOI21_X1 U8957 ( .B1(n7169), .B2(n9431), .A(n7168), .ZN(n7170) );
  OAI211_X1 U8958 ( .C1(n7172), .C2(n9367), .A(n7171), .B(n7170), .ZN(P1_U3288) );
  OAI21_X1 U8959 ( .B1(n7175), .B2(n7178), .A(n7174), .ZN(n7176) );
  INV_X1 U8960 ( .A(n7176), .ZN(n7194) );
  XOR2_X1 U8961 ( .A(n7178), .B(n7177), .Z(n7179) );
  AOI222_X1 U8962 ( .A1(n9137), .A2(n9393), .B1(n9135), .B2(n9390), .C1(n9746), 
        .C2(n7179), .ZN(n7187) );
  AOI21_X1 U8963 ( .B1(n7723), .B2(n7181), .A(n7180), .ZN(n7191) );
  AOI22_X1 U8964 ( .A1(n7191), .A2(n9477), .B1(n9724), .B2(n7723), .ZN(n7182)
         );
  OAI211_X1 U8965 ( .C1(n9516), .C2(n7194), .A(n7187), .B(n7182), .ZN(n7184)
         );
  NAND2_X1 U8966 ( .A1(n7184), .A2(n9757), .ZN(n7183) );
  OAI21_X1 U8967 ( .B1(n9757), .B2(n6536), .A(n7183), .ZN(P1_U3528) );
  INV_X1 U8968 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n7186) );
  NAND2_X1 U8969 ( .A1(n7184), .A2(n9749), .ZN(n7185) );
  OAI21_X1 U8970 ( .B1(n9749), .B2(n7186), .A(n7185), .ZN(P1_U3471) );
  MUX2_X1 U8971 ( .A(n6549), .B(n7187), .S(n9381), .Z(n7193) );
  INV_X1 U8972 ( .A(n7188), .ZN(n7189) );
  OAI22_X1 U8973 ( .A1(n9429), .A2(n4576), .B1(n7189), .B2(n7333), .ZN(n7190)
         );
  AOI21_X1 U8974 ( .B1(n7191), .B2(n9326), .A(n7190), .ZN(n7192) );
  OAI211_X1 U8975 ( .C1(n7194), .C2(n9404), .A(n7193), .B(n7192), .ZN(P1_U3287) );
  XNOR2_X1 U8976 ( .A(n7195), .B(n8477), .ZN(n7265) );
  INV_X1 U8977 ( .A(n7265), .ZN(n7207) );
  AND2_X1 U8978 ( .A1(n7197), .A2(n7196), .ZN(n7198) );
  NAND2_X1 U8979 ( .A1(n7200), .A2(n7198), .ZN(n7202) );
  AND2_X1 U8980 ( .A1(n7200), .A2(n7199), .ZN(n7201) );
  AOI21_X1 U8981 ( .B1(n8477), .B2(n7202), .A(n7201), .ZN(n7203) );
  OAI222_X1 U8982 ( .A1(n8788), .A2(n7993), .B1(n8790), .B2(n7396), .C1(n8786), 
        .C2(n7203), .ZN(n7264) );
  NAND2_X1 U8983 ( .A1(n7264), .A2(n9824), .ZN(n7206) );
  OAI22_X1 U8984 ( .A1(n9824), .A2(n7352), .B1(n7374), .B2(n8679), .ZN(n7204)
         );
  AOI21_X1 U8985 ( .B1(n9819), .B2(n7369), .A(n7204), .ZN(n7205) );
  OAI211_X1 U8986 ( .C1(n8673), .C2(n7207), .A(n7206), .B(n7205), .ZN(P2_U3224) );
  OAI21_X1 U8987 ( .B1(n7209), .B2(n7216), .A(n7208), .ZN(n7307) );
  INV_X1 U8988 ( .A(n7210), .ZN(n7213) );
  INV_X1 U8989 ( .A(n7211), .ZN(n7212) );
  AOI211_X1 U8990 ( .C1(n7292), .C2(n7213), .A(n9422), .B(n7212), .ZN(n7313)
         );
  NAND2_X1 U8991 ( .A1(n7215), .A2(n7214), .ZN(n7217) );
  XNOR2_X1 U8992 ( .A(n7217), .B(n7216), .ZN(n7221) );
  OR2_X1 U8993 ( .A1(n7324), .A2(n9414), .ZN(n7219) );
  NAND2_X1 U8994 ( .A1(n9135), .A2(n9393), .ZN(n7218) );
  NAND2_X1 U8995 ( .A1(n7219), .A2(n7218), .ZN(n7289) );
  INV_X1 U8996 ( .A(n7289), .ZN(n7220) );
  OAI21_X1 U8997 ( .B1(n7221), .B2(n9496), .A(n7220), .ZN(n7308) );
  AOI211_X1 U8998 ( .C1(n9734), .C2(n7307), .A(n7313), .B(n7308), .ZN(n7226)
         );
  AOI22_X1 U8999 ( .A1(n8073), .A2(n7292), .B1(n9754), .B2(
        P1_REG1_REG_8__SCAN_IN), .ZN(n7222) );
  OAI21_X1 U9000 ( .B1(n7226), .B2(n9754), .A(n7222), .ZN(P1_U3530) );
  INV_X1 U9001 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n7223) );
  OAI22_X1 U9002 ( .A1(n9576), .A2(n7309), .B1(n9749), .B2(n7223), .ZN(n7224)
         );
  INV_X1 U9003 ( .A(n7224), .ZN(n7225) );
  OAI21_X1 U9004 ( .B1(n7226), .B2(n9747), .A(n7225), .ZN(P1_U3477) );
  INV_X1 U9005 ( .A(n8473), .ZN(n7228) );
  XNOR2_X1 U9006 ( .A(n7227), .B(n7228), .ZN(n9854) );
  OAI22_X1 U9007 ( .A1(n8798), .A2(n9850), .B1(n8251), .B2(n8679), .ZN(n7233)
         );
  OR2_X1 U9008 ( .A1(n7123), .A2(n7228), .ZN(n7298) );
  NAND2_X1 U9009 ( .A1(n7123), .A2(n7228), .ZN(n7229) );
  NAND3_X1 U9010 ( .A1(n7298), .A2(n8759), .A3(n7229), .ZN(n7231) );
  AOI22_X1 U9011 ( .A1(n8745), .A2(n8537), .B1(n8535), .B2(n8763), .ZN(n7230)
         );
  NAND2_X1 U9012 ( .A1(n7231), .A2(n7230), .ZN(n9851) );
  MUX2_X1 U9013 ( .A(n9851), .B(P2_REG2_REG_6__SCAN_IN), .S(n8803), .Z(n7232)
         );
  AOI211_X1 U9014 ( .C1(n8801), .C2(n9854), .A(n7233), .B(n7232), .ZN(n7234)
         );
  INV_X1 U9015 ( .A(n7234), .ZN(P2_U3227) );
  INV_X1 U9016 ( .A(n9859), .ZN(n7263) );
  INV_X1 U9017 ( .A(n8269), .ZN(n8285) );
  INV_X1 U9018 ( .A(n8537), .ZN(n7235) );
  NAND2_X1 U9019 ( .A1(n7236), .A2(n7235), .ZN(n7237) );
  XNOR2_X1 U9020 ( .A(n7239), .B(n8536), .ZN(n8247) );
  INV_X1 U9021 ( .A(n7239), .ZN(n7240) );
  INV_X1 U9022 ( .A(n7397), .ZN(n7246) );
  XNOR2_X1 U9023 ( .A(n9820), .B(n4353), .ZN(n7242) );
  NAND2_X1 U9024 ( .A1(n7242), .A2(n7241), .ZN(n7249) );
  INV_X1 U9025 ( .A(n7242), .ZN(n7243) );
  NAND2_X1 U9026 ( .A1(n7243), .A2(n8535), .ZN(n7244) );
  NAND2_X1 U9027 ( .A1(n7249), .A2(n7244), .ZN(n7399) );
  INV_X1 U9028 ( .A(n7399), .ZN(n7245) );
  NAND2_X1 U9029 ( .A1(n7246), .A2(n7245), .ZN(n7250) );
  INV_X1 U9030 ( .A(n7247), .ZN(n7398) );
  INV_X1 U9031 ( .A(n7249), .ZN(n7248) );
  XNOR2_X1 U9032 ( .A(n9859), .B(n4353), .ZN(n7366) );
  XNOR2_X1 U9033 ( .A(n7366), .B(n8534), .ZN(n7251) );
  NOR3_X1 U9034 ( .A1(n7398), .A2(n7248), .A3(n7251), .ZN(n7254) );
  NAND2_X1 U9035 ( .A1(n7250), .A2(n7249), .ZN(n7252) );
  NAND2_X1 U9036 ( .A1(n7252), .A2(n7251), .ZN(n7368) );
  INV_X1 U9037 ( .A(n7368), .ZN(n7253) );
  OAI21_X1 U9038 ( .B1(n7254), .B2(n7253), .A(n8273), .ZN(n7262) );
  INV_X1 U9039 ( .A(n7255), .ZN(n7256) );
  AOI21_X1 U9040 ( .B1(n8277), .B2(n8535), .A(n7256), .ZN(n7257) );
  OAI21_X1 U9041 ( .B1(n7258), .B2(n8279), .A(n7257), .ZN(n7259) );
  AOI21_X1 U9042 ( .B1(n7260), .B2(n8281), .A(n7259), .ZN(n7261) );
  OAI211_X1 U9043 ( .C1(n7263), .C2(n8285), .A(n7262), .B(n7261), .ZN(P2_U3161) );
  AOI21_X1 U9044 ( .B1(n7265), .B2(n9853), .A(n7264), .ZN(n7270) );
  INV_X1 U9045 ( .A(n8874), .ZN(n8816) );
  AOI22_X1 U9046 ( .A1(n8816), .A2(n7369), .B1(n9885), .B2(
        P2_REG1_REG_9__SCAN_IN), .ZN(n7266) );
  OAI21_X1 U9047 ( .B1(n7270), .B2(n9885), .A(n7266), .ZN(P2_U3468) );
  INV_X1 U9048 ( .A(n8943), .ZN(n8891) );
  INV_X1 U9049 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n7267) );
  NOR2_X1 U9050 ( .A1(n8939), .A2(n7267), .ZN(n7268) );
  AOI21_X1 U9051 ( .B1(n8891), .B2(n7369), .A(n7268), .ZN(n7269) );
  OAI21_X1 U9052 ( .B1(n7270), .B2(n9873), .A(n7269), .ZN(P2_U3417) );
  OAI211_X1 U9053 ( .C1(n7273), .C2(n9496), .A(n7272), .B(n7271), .ZN(n7274)
         );
  AOI21_X1 U9054 ( .B1(n9734), .B2(n7275), .A(n7274), .ZN(n7282) );
  INV_X1 U9055 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n7276) );
  OAI22_X1 U9056 ( .A1(n9524), .A2(n7390), .B1(n9757), .B2(n7276), .ZN(n7277)
         );
  INV_X1 U9057 ( .A(n7277), .ZN(n7278) );
  OAI21_X1 U9058 ( .B1(n7282), .B2(n9754), .A(n7278), .ZN(P1_U3531) );
  INV_X1 U9059 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n7279) );
  OAI22_X1 U9060 ( .A1(n9576), .A2(n7390), .B1(n9749), .B2(n7279), .ZN(n7280)
         );
  INV_X1 U9061 ( .A(n7280), .ZN(n7281) );
  OAI21_X1 U9062 ( .B1(n7282), .B2(n9747), .A(n7281), .ZN(P1_U3480) );
  INV_X1 U9063 ( .A(n7283), .ZN(n7284) );
  AOI21_X1 U9064 ( .B1(n7286), .B2(n7285), .A(n7284), .ZN(n7294) );
  INV_X1 U9065 ( .A(n7287), .ZN(n7288) );
  AOI21_X1 U9066 ( .B1(n7289), .B2(n9618), .A(n7288), .ZN(n7290) );
  OAI21_X1 U9067 ( .B1(n7310), .B2(n9631), .A(n7290), .ZN(n7291) );
  AOI21_X1 U9068 ( .B1(n7292), .B2(n9628), .A(n7291), .ZN(n7293) );
  OAI21_X1 U9069 ( .B1(n7294), .B2(n9623), .A(n7293), .ZN(P1_U3221) );
  XNOR2_X1 U9070 ( .A(n7295), .B(n8475), .ZN(n9817) );
  AND2_X1 U9071 ( .A1(n7298), .A2(n7296), .ZN(n7300) );
  NAND2_X1 U9072 ( .A1(n7298), .A2(n7297), .ZN(n7299) );
  OAI21_X1 U9073 ( .B1(n7301), .B2(n7300), .A(n7299), .ZN(n7302) );
  AOI222_X1 U9074 ( .A1(n8759), .A2(n7302), .B1(n8534), .B2(n8763), .C1(n8536), 
        .C2(n8745), .ZN(n9816) );
  OAI21_X1 U9075 ( .B1(n9866), .B2(n9817), .A(n9816), .ZN(n7319) );
  INV_X1 U9076 ( .A(n7319), .ZN(n7304) );
  AOI22_X1 U9077 ( .A1(n8816), .A2(n9820), .B1(n9885), .B2(
        P2_REG1_REG_7__SCAN_IN), .ZN(n7303) );
  OAI21_X1 U9078 ( .B1(n7304), .B2(n9885), .A(n7303), .ZN(P2_U3466) );
  INV_X1 U9079 ( .A(n7305), .ZN(n7695) );
  INV_X1 U9080 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7306) );
  OAI222_X1 U9081 ( .A1(n6405), .A2(P2_U3151), .B1(n8960), .B2(n7695), .C1(
        n7306), .C2(n8956), .ZN(P2_U3276) );
  INV_X1 U9082 ( .A(n7307), .ZN(n7316) );
  NAND2_X1 U9083 ( .A1(n7308), .A2(n9381), .ZN(n7315) );
  NOR2_X1 U9084 ( .A1(n9429), .A2(n7309), .ZN(n7312) );
  OAI22_X1 U9085 ( .A1(n9381), .A2(n6601), .B1(n7310), .B2(n7333), .ZN(n7311)
         );
  AOI211_X1 U9086 ( .C1(n7313), .C2(n9431), .A(n7312), .B(n7311), .ZN(n7314)
         );
  OAI211_X1 U9087 ( .C1(n7316), .C2(n9404), .A(n7315), .B(n7314), .ZN(P1_U3285) );
  INV_X1 U9088 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n7317) );
  OAI22_X1 U9089 ( .A1(n8350), .A2(n8943), .B1(n8939), .B2(n7317), .ZN(n7318)
         );
  AOI21_X1 U9090 ( .B1(n7319), .B2(n8939), .A(n7318), .ZN(n7320) );
  INV_X1 U9091 ( .A(n7320), .ZN(P2_U3411) );
  INV_X1 U9092 ( .A(n7430), .ZN(n7323) );
  AOI21_X1 U9093 ( .B1(n7321), .B2(n7948), .A(n7855), .ZN(n7322) );
  OAI21_X1 U9094 ( .B1(n7323), .B2(n7322), .A(n9746), .ZN(n7328) );
  OR2_X1 U9095 ( .A1(n7324), .A2(n9412), .ZN(n7326) );
  OR2_X1 U9096 ( .A1(n7460), .A2(n9414), .ZN(n7325) );
  NAND2_X1 U9097 ( .A1(n7326), .A2(n7325), .ZN(n9619) );
  INV_X1 U9098 ( .A(n9619), .ZN(n7327) );
  NAND2_X1 U9099 ( .A1(n7328), .A2(n7327), .ZN(n7358) );
  INV_X1 U9100 ( .A(n7358), .ZN(n7339) );
  OAI21_X1 U9101 ( .B1(n7331), .B2(n7330), .A(n7329), .ZN(n7360) );
  NAND2_X1 U9102 ( .A1(n7360), .A2(n9355), .ZN(n7338) );
  AOI211_X1 U9103 ( .C1(n9629), .C2(n7332), .A(n9422), .B(n7436), .ZN(n7359)
         );
  NOR2_X1 U9104 ( .A1(n9429), .A2(n5750), .ZN(n7336) );
  OAI22_X1 U9105 ( .A1(n9381), .A2(n7334), .B1(n9632), .B2(n7333), .ZN(n7335)
         );
  AOI211_X1 U9106 ( .C1(n7359), .C2(n9431), .A(n7336), .B(n7335), .ZN(n7337)
         );
  OAI211_X1 U9107 ( .C1(n9211), .C2(n7339), .A(n7338), .B(n7337), .ZN(P1_U3283) );
  AOI21_X1 U9108 ( .B1(n7342), .B2(n7341), .A(n7340), .ZN(n7357) );
  NAND2_X1 U9109 ( .A1(n9772), .A2(n7343), .ZN(n7349) );
  NAND2_X1 U9110 ( .A1(P2_U3151), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n7372) );
  OAI21_X1 U9111 ( .B1(n7346), .B2(n7345), .A(n7344), .ZN(n7347) );
  NAND2_X1 U9112 ( .A1(n9807), .A2(n7347), .ZN(n7348) );
  NAND3_X1 U9113 ( .A1(n7349), .A2(n7372), .A3(n7348), .ZN(n7355) );
  AOI21_X1 U9114 ( .B1(n7352), .B2(n7351), .A(n7350), .ZN(n7353) );
  NOR2_X1 U9115 ( .A1(n7353), .A2(n9810), .ZN(n7354) );
  AOI211_X1 U9116 ( .C1(n9796), .C2(P2_ADDR_REG_9__SCAN_IN), .A(n7355), .B(
        n7354), .ZN(n7356) );
  OAI21_X1 U9117 ( .B1(n7357), .B2(n9803), .A(n7356), .ZN(P2_U3191) );
  AOI211_X1 U9118 ( .C1(n7360), .C2(n9734), .A(n7359), .B(n7358), .ZN(n7365)
         );
  AOI22_X1 U9119 ( .A1(n9629), .A2(n8073), .B1(n9754), .B2(
        P1_REG1_REG_10__SCAN_IN), .ZN(n7361) );
  OAI21_X1 U9120 ( .B1(n7365), .B2(n9754), .A(n7361), .ZN(P1_U3532) );
  INV_X1 U9121 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n7362) );
  NOR2_X1 U9122 ( .A1(n9749), .A2(n7362), .ZN(n7363) );
  AOI21_X1 U9123 ( .B1(n8078), .B2(n9629), .A(n7363), .ZN(n7364) );
  OAI21_X1 U9124 ( .B1(n7365), .B2(n9747), .A(n7364), .ZN(P1_U3483) );
  INV_X1 U9125 ( .A(n7369), .ZN(n7379) );
  NAND2_X1 U9126 ( .A1(n7366), .A2(n7396), .ZN(n7367) );
  XNOR2_X1 U9127 ( .A(n7369), .B(n4353), .ZN(n7501) );
  XNOR2_X1 U9128 ( .A(n7501), .B(n8533), .ZN(n7370) );
  OAI211_X1 U9129 ( .C1(n7371), .C2(n7370), .A(n7504), .B(n8273), .ZN(n7378)
         );
  NAND2_X1 U9130 ( .A1(n8277), .A2(n8534), .ZN(n7373) );
  OAI211_X1 U9131 ( .C1(n7993), .C2(n8279), .A(n7373), .B(n7372), .ZN(n7376)
         );
  NOR2_X1 U9132 ( .A1(n8267), .A2(n7374), .ZN(n7375) );
  NOR2_X1 U9133 ( .A1(n7376), .A2(n7375), .ZN(n7377) );
  OAI211_X1 U9134 ( .C1(n7379), .C2(n8285), .A(n7378), .B(n7377), .ZN(P2_U3171) );
  OAI21_X1 U9135 ( .B1(n7382), .B2(n7381), .A(n7380), .ZN(n7383) );
  NAND2_X1 U9136 ( .A1(n7383), .A2(n9102), .ZN(n7389) );
  NAND2_X1 U9137 ( .A1(n9104), .A2(n9132), .ZN(n7384) );
  NAND2_X1 U9138 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n9613) );
  OAI211_X1 U9139 ( .C1(n7385), .C2(n9106), .A(n7384), .B(n9613), .ZN(n7386)
         );
  AOI21_X1 U9140 ( .B1(n7387), .B2(n9109), .A(n7386), .ZN(n7388) );
  OAI211_X1 U9141 ( .C1(n7390), .C2(n9113), .A(n7389), .B(n7388), .ZN(P1_U3231) );
  INV_X1 U9142 ( .A(n7391), .ZN(n7392) );
  AOI21_X1 U9143 ( .B1(n8277), .B2(n8536), .A(n7392), .ZN(n7395) );
  INV_X1 U9144 ( .A(n7393), .ZN(n9822) );
  NAND2_X1 U9145 ( .A1(n8281), .A2(n9822), .ZN(n7394) );
  OAI211_X1 U9146 ( .C1(n7396), .C2(n8279), .A(n7395), .B(n7394), .ZN(n7402)
         );
  AOI21_X1 U9147 ( .B1(n7397), .B2(n7399), .A(n7398), .ZN(n7400) );
  NOR2_X1 U9148 ( .A1(n7400), .A2(n8271), .ZN(n7401) );
  AOI211_X1 U9149 ( .C1(n9820), .C2(n8269), .A(n7402), .B(n7401), .ZN(n7403)
         );
  INV_X1 U9150 ( .A(n7403), .ZN(P2_U3153) );
  INV_X1 U9151 ( .A(n7404), .ZN(n7425) );
  OAI222_X1 U9152 ( .A1(n9591), .A2(n7425), .B1(n7927), .B2(P1_U3086), .C1(
        n7405), .C2(n9588), .ZN(P1_U3335) );
  AOI21_X1 U9153 ( .B1(n7408), .B2(n7407), .A(n7406), .ZN(n7423) );
  NAND2_X1 U9154 ( .A1(n9772), .A2(n7409), .ZN(n7415) );
  INV_X1 U9155 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n10093) );
  OR2_X1 U9156 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10093), .ZN(n7509) );
  OAI21_X1 U9157 ( .B1(n7412), .B2(n7411), .A(n7410), .ZN(n7413) );
  NAND2_X1 U9158 ( .A1(n9807), .A2(n7413), .ZN(n7414) );
  NAND3_X1 U9159 ( .A1(n7415), .A2(n7509), .A3(n7414), .ZN(n7421) );
  AOI21_X1 U9160 ( .B1(n7418), .B2(n7417), .A(n7416), .ZN(n7419) );
  NOR2_X1 U9161 ( .A1(n7419), .A2(n9803), .ZN(n7420) );
  AOI211_X1 U9162 ( .C1(n9796), .C2(P2_ADDR_REG_10__SCAN_IN), .A(n7421), .B(
        n7420), .ZN(n7422) );
  OAI21_X1 U9163 ( .B1(n7423), .B2(n9810), .A(n7422), .ZN(P2_U3192) );
  OAI222_X1 U9164 ( .A1(P2_U3151), .A2(n7426), .B1(n8960), .B2(n7425), .C1(
        n7424), .C2(n8956), .ZN(P2_U3275) );
  OAI21_X1 U9165 ( .B1(n7428), .B2(n7858), .A(n7427), .ZN(n7444) );
  INV_X1 U9166 ( .A(n7444), .ZN(n7441) );
  NAND2_X1 U9167 ( .A1(n7457), .A2(n9746), .ZN(n7435) );
  INV_X1 U9168 ( .A(n7858), .ZN(n7429) );
  AOI21_X1 U9169 ( .B1(n7430), .B2(n7746), .A(n7429), .ZN(n7434) );
  OR2_X1 U9170 ( .A1(n7531), .A2(n9414), .ZN(n7433) );
  OR2_X1 U9171 ( .A1(n7431), .A2(n9412), .ZN(n7432) );
  AND2_X1 U9172 ( .A1(n7433), .A2(n7432), .ZN(n7603) );
  OAI21_X1 U9173 ( .B1(n7435), .B2(n7434), .A(n7603), .ZN(n7442) );
  AOI211_X1 U9174 ( .C1(n7446), .C2(n4564), .A(n9422), .B(n7464), .ZN(n7443)
         );
  NAND2_X1 U9175 ( .A1(n7443), .A2(n9431), .ZN(n7438) );
  AOI22_X1 U9176 ( .A1(n9433), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n7605), .B2(
        n9426), .ZN(n7437) );
  OAI211_X1 U9177 ( .C1(n7608), .C2(n9429), .A(n7438), .B(n7437), .ZN(n7439)
         );
  AOI21_X1 U9178 ( .B1(n9381), .B2(n7442), .A(n7439), .ZN(n7440) );
  OAI21_X1 U9179 ( .B1(n7441), .B2(n9404), .A(n7440), .ZN(P1_U3282) );
  AOI211_X1 U9180 ( .C1(n7444), .C2(n9734), .A(n7443), .B(n7442), .ZN(n7448)
         );
  AOI22_X1 U9181 ( .A1(n7446), .A2(n8073), .B1(P1_REG1_REG_11__SCAN_IN), .B2(
        n9754), .ZN(n7445) );
  OAI21_X1 U9182 ( .B1(n7448), .B2(n9754), .A(n7445), .ZN(P1_U3533) );
  AOI22_X1 U9183 ( .A1(n7446), .A2(n8078), .B1(P1_REG0_REG_11__SCAN_IN), .B2(
        n9747), .ZN(n7447) );
  OAI21_X1 U9184 ( .B1(n7448), .B2(n9747), .A(n7447), .ZN(P1_U3486) );
  XNOR2_X1 U9185 ( .A(n7449), .B(n8379), .ZN(n9867) );
  XNOR2_X1 U9186 ( .A(n7450), .B(n8379), .ZN(n7451) );
  OAI222_X1 U9187 ( .A1(n8788), .A2(n7589), .B1(n8790), .B2(n7561), .C1(n7451), 
        .C2(n8786), .ZN(n9868) );
  NAND2_X1 U9188 ( .A1(n9868), .A2(n9824), .ZN(n7454) );
  OAI22_X1 U9189 ( .A1(n9824), .A2(n5935), .B1(n7567), .B2(n8679), .ZN(n7452)
         );
  AOI21_X1 U9190 ( .B1(n9870), .B2(n9819), .A(n7452), .ZN(n7453) );
  OAI211_X1 U9191 ( .C1(n8673), .C2(n9867), .A(n7454), .B(n7453), .ZN(P2_U3221) );
  OAI21_X1 U9192 ( .B1(n7456), .B2(n7859), .A(n7455), .ZN(n7551) );
  INV_X1 U9193 ( .A(n7551), .ZN(n7471) );
  NAND2_X1 U9194 ( .A1(n7457), .A2(n7752), .ZN(n7458) );
  XNOR2_X1 U9195 ( .A(n7458), .B(n7859), .ZN(n7459) );
  NAND2_X1 U9196 ( .A1(n7459), .A2(n9746), .ZN(n7463) );
  OR2_X1 U9197 ( .A1(n9413), .A2(n9414), .ZN(n7462) );
  OR2_X1 U9198 ( .A1(n7460), .A2(n9412), .ZN(n7461) );
  AND2_X1 U9199 ( .A1(n7462), .A2(n7461), .ZN(n7626) );
  NAND2_X1 U9200 ( .A1(n7463), .A2(n7626), .ZN(n7549) );
  INV_X1 U9201 ( .A(n7464), .ZN(n7466) );
  INV_X1 U9202 ( .A(n7535), .ZN(n7465) );
  AOI211_X1 U9203 ( .C1(n7628), .C2(n7466), .A(n9422), .B(n7465), .ZN(n7550)
         );
  NAND2_X1 U9204 ( .A1(n7550), .A2(n9431), .ZN(n7468) );
  AOI22_X1 U9205 ( .A1(n9433), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n7623), .B2(
        n9426), .ZN(n7467) );
  OAI211_X1 U9206 ( .C1(n5753), .C2(n9429), .A(n7468), .B(n7467), .ZN(n7469)
         );
  AOI21_X1 U9207 ( .B1(n9381), .B2(n7549), .A(n7469), .ZN(n7470) );
  OAI21_X1 U9208 ( .B1(n7471), .B2(n9404), .A(n7470), .ZN(P1_U3281) );
  AOI21_X1 U9209 ( .B1(n7474), .B2(n7473), .A(n7472), .ZN(n7487) );
  AOI21_X1 U9210 ( .B1(n7476), .B2(n9883), .A(n7475), .ZN(n7484) );
  OAI21_X1 U9211 ( .B1(n7479), .B2(n7478), .A(n7477), .ZN(n7480) );
  AOI22_X1 U9212 ( .A1(n9796), .A2(P2_ADDR_REG_11__SCAN_IN), .B1(n9807), .B2(
        n7480), .ZN(n7483) );
  INV_X1 U9213 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n10070) );
  NOR2_X1 U9214 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10070), .ZN(n7609) );
  AOI21_X1 U9215 ( .B1(n9772), .B2(n7481), .A(n7609), .ZN(n7482) );
  OAI211_X1 U9216 ( .C1(n7484), .C2(n9803), .A(n7483), .B(n7482), .ZN(n7485)
         );
  INV_X1 U9217 ( .A(n7485), .ZN(n7486) );
  OAI21_X1 U9218 ( .B1(n7487), .B2(n9810), .A(n7486), .ZN(P2_U3193) );
  XOR2_X1 U9219 ( .A(n7488), .B(n8479), .Z(n7522) );
  XNOR2_X1 U9220 ( .A(n7489), .B(n8479), .ZN(n7490) );
  AOI222_X1 U9221 ( .A1(n8759), .A2(n7490), .B1(n8531), .B2(n8763), .C1(n8533), 
        .C2(n8745), .ZN(n7527) );
  OAI21_X1 U9222 ( .B1(n9866), .B2(n7522), .A(n7527), .ZN(n7495) );
  INV_X1 U9223 ( .A(n7525), .ZN(n8374) );
  OAI22_X1 U9224 ( .A1(n8374), .A2(n8874), .B1(n9887), .B2(n6181), .ZN(n7491)
         );
  AOI21_X1 U9225 ( .B1(n7495), .B2(n9887), .A(n7491), .ZN(n7492) );
  INV_X1 U9226 ( .A(n7492), .ZN(P2_U3469) );
  INV_X1 U9227 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n7493) );
  OAI22_X1 U9228 ( .A1(n8374), .A2(n8943), .B1(n8939), .B2(n7493), .ZN(n7494)
         );
  AOI21_X1 U9229 ( .B1(n7495), .B2(n8939), .A(n7494), .ZN(n7496) );
  INV_X1 U9230 ( .A(n7496), .ZN(P2_U3420) );
  INV_X1 U9231 ( .A(n7497), .ZN(n7500) );
  OAI222_X1 U9232 ( .A1(n9588), .A2(n7498), .B1(n9591), .B2(n7500), .C1(
        P1_U3086), .C2(n7931), .ZN(P1_U3334) );
  OAI222_X1 U9233 ( .A1(n8315), .A2(P2_U3151), .B1(n8960), .B2(n7500), .C1(
        n7499), .C2(n8956), .ZN(P2_U3274) );
  INV_X1 U9234 ( .A(n7501), .ZN(n7502) );
  NAND2_X1 U9235 ( .A1(n7502), .A2(n8533), .ZN(n7503) );
  XNOR2_X1 U9236 ( .A(n7525), .B(n4353), .ZN(n7506) );
  OAI21_X1 U9237 ( .B1(n7507), .B2(n7506), .A(n7505), .ZN(n7508) );
  NAND2_X1 U9238 ( .A1(n7508), .A2(n8273), .ZN(n7514) );
  NAND2_X1 U9239 ( .A1(n8277), .A2(n8533), .ZN(n7510) );
  OAI211_X1 U9240 ( .C1(n7561), .C2(n8279), .A(n7510), .B(n7509), .ZN(n7512)
         );
  NOR2_X1 U9241 ( .A1(n8267), .A2(n7520), .ZN(n7511) );
  NOR2_X1 U9242 ( .A1(n7512), .A2(n7511), .ZN(n7513) );
  OAI211_X1 U9243 ( .C1(n8374), .C2(n8285), .A(n7514), .B(n7513), .ZN(P2_U3157) );
  INV_X1 U9244 ( .A(n7515), .ZN(n7518) );
  OAI222_X1 U9245 ( .A1(n9588), .A2(n7516), .B1(n9591), .B2(n7518), .C1(
        P1_U3086), .C2(n7841), .ZN(P1_U3333) );
  OAI222_X1 U9246 ( .A1(n7519), .A2(P2_U3151), .B1(n8960), .B2(n7518), .C1(
        n7517), .C2(n8956), .ZN(P2_U3273) );
  OAI22_X1 U9247 ( .A1(n9824), .A2(n7521), .B1(n7520), .B2(n8679), .ZN(n7524)
         );
  NOR2_X1 U9248 ( .A1(n7522), .A2(n8673), .ZN(n7523) );
  AOI211_X1 U9249 ( .C1(n9819), .C2(n7525), .A(n7524), .B(n7523), .ZN(n7526)
         );
  OAI21_X1 U9250 ( .B1(n8803), .B2(n7527), .A(n7526), .ZN(P2_U3223) );
  XNOR2_X1 U9251 ( .A(n7528), .B(n7845), .ZN(n7633) );
  OAI21_X1 U9252 ( .B1(n7529), .B2(n7845), .A(n7530), .ZN(n7635) );
  NAND2_X1 U9253 ( .A1(n7635), .A2(n9355), .ZN(n7541) );
  OR2_X1 U9254 ( .A1(n7531), .A2(n9412), .ZN(n7533) );
  OR2_X1 U9255 ( .A1(n9107), .A2(n9414), .ZN(n7532) );
  NAND2_X1 U9256 ( .A1(n7533), .A2(n7532), .ZN(n9062) );
  INV_X1 U9257 ( .A(n9062), .ZN(n7632) );
  AOI22_X1 U9258 ( .A1(n9433), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n9061), .B2(
        n9426), .ZN(n7534) );
  OAI21_X1 U9259 ( .B1(n7632), .B2(n9433), .A(n7534), .ZN(n7539) );
  AOI21_X1 U9260 ( .B1(n7535), .B2(n9066), .A(n9422), .ZN(n7537) );
  NAND2_X1 U9261 ( .A1(n7537), .A2(n9424), .ZN(n7631) );
  NOR2_X1 U9262 ( .A1(n7631), .A2(n9360), .ZN(n7538) );
  AOI211_X1 U9263 ( .C1(n9364), .C2(n9066), .A(n7539), .B(n7538), .ZN(n7540)
         );
  OAI211_X1 U9264 ( .C1(n7633), .C2(n9367), .A(n7541), .B(n7540), .ZN(P1_U3280) );
  XNOR2_X1 U9265 ( .A(n8388), .B(n7589), .ZN(n8485) );
  XOR2_X1 U9266 ( .A(n7542), .B(n8485), .Z(n7543) );
  OAI222_X1 U9267 ( .A1(n8788), .A2(n8096), .B1(n8790), .B2(n7992), .C1(n8786), 
        .C2(n7543), .ZN(n8870) );
  OAI22_X1 U9268 ( .A1(n8944), .A2(n8686), .B1(n7679), .B2(n8679), .ZN(n7544)
         );
  OAI21_X1 U9269 ( .B1(n8870), .B2(n7544), .A(n9824), .ZN(n7548) );
  OR2_X1 U9270 ( .A1(n7449), .A2(n8379), .ZN(n7545) );
  NAND2_X1 U9271 ( .A1(n7545), .A2(n8383), .ZN(n7546) );
  XNOR2_X1 U9272 ( .A(n7546), .B(n8485), .ZN(n8871) );
  AOI22_X1 U9273 ( .A1(n8871), .A2(n8801), .B1(P2_REG2_REG_13__SCAN_IN), .B2(
        n8803), .ZN(n7547) );
  NAND2_X1 U9274 ( .A1(n7548), .A2(n7547), .ZN(P2_U3220) );
  AOI211_X1 U9275 ( .C1(n7551), .C2(n9734), .A(n7550), .B(n7549), .ZN(n7554)
         );
  MUX2_X1 U9276 ( .A(n7552), .B(n7554), .S(n9757), .Z(n7553) );
  OAI21_X1 U9277 ( .B1(n5753), .B2(n9524), .A(n7553), .ZN(P1_U3534) );
  INV_X1 U9278 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n7555) );
  MUX2_X1 U9279 ( .A(n7555), .B(n7554), .S(n9749), .Z(n7556) );
  OAI21_X1 U9280 ( .B1(n5753), .B2(n9576), .A(n7556), .ZN(P1_U3489) );
  NAND2_X1 U9281 ( .A1(n8373), .A2(n8371), .ZN(n8465) );
  XNOR2_X1 U9282 ( .A(n8465), .B(n8124), .ZN(n7615) );
  NAND2_X1 U9283 ( .A1(n7560), .A2(n7559), .ZN(n7613) );
  NAND2_X1 U9284 ( .A1(n7562), .A2(n8531), .ZN(n7563) );
  NAND2_X1 U9285 ( .A1(n7613), .A2(n7563), .ZN(n7674) );
  XNOR2_X1 U9286 ( .A(n9870), .B(n4353), .ZN(n7671) );
  XNOR2_X1 U9287 ( .A(n7671), .B(n8530), .ZN(n7673) );
  XNOR2_X1 U9288 ( .A(n7674), .B(n7673), .ZN(n7570) );
  INV_X1 U9289 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7564) );
  NOR2_X1 U9290 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7564), .ZN(n7652) );
  NOR2_X1 U9291 ( .A1(n8279), .A2(n7589), .ZN(n7565) );
  AOI211_X1 U9292 ( .C1(n8277), .C2(n8531), .A(n7652), .B(n7565), .ZN(n7566)
         );
  OAI21_X1 U9293 ( .B1(n7567), .B2(n8267), .A(n7566), .ZN(n7568) );
  AOI21_X1 U9294 ( .B1(n9870), .B2(n8269), .A(n7568), .ZN(n7569) );
  OAI21_X1 U9295 ( .B1(n7570), .B2(n8271), .A(n7569), .ZN(P2_U3164) );
  NAND2_X1 U9296 ( .A1(n7574), .A2(n7571), .ZN(n7572) );
  OAI211_X1 U9297 ( .C1(n7573), .C2(n9588), .A(n7572), .B(n7986), .ZN(P1_U3332) );
  NAND2_X1 U9298 ( .A1(n7574), .A2(n8953), .ZN(n7576) );
  NAND2_X1 U9299 ( .A1(n7575), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8519) );
  OAI211_X1 U9300 ( .C1(n7577), .C2(n8956), .A(n7576), .B(n8519), .ZN(P2_U3272) );
  OAI21_X1 U9301 ( .B1(n7579), .B2(n8394), .A(n7578), .ZN(n7580) );
  AOI222_X1 U9302 ( .A1(n8759), .A2(n7580), .B1(n8526), .B2(n8763), .C1(n8528), 
        .C2(n8745), .ZN(n8861) );
  XNOR2_X1 U9303 ( .A(n7581), .B(n8394), .ZN(n8863) );
  INV_X1 U9304 ( .A(n7582), .ZN(n8282) );
  AOI22_X1 U9305 ( .A1(n8803), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n9821), .B2(
        n8282), .ZN(n7583) );
  OAI21_X1 U9306 ( .B1(n8934), .B2(n8798), .A(n7583), .ZN(n7584) );
  AOI21_X1 U9307 ( .B1(n8863), .B2(n8801), .A(n7584), .ZN(n7585) );
  OAI21_X1 U9308 ( .B1(n8861), .B2(n8803), .A(n7585), .ZN(P2_U3218) );
  INV_X1 U9309 ( .A(n8686), .ZN(n7591) );
  INV_X1 U9310 ( .A(n7586), .ZN(n8395) );
  NAND2_X1 U9311 ( .A1(n8395), .A2(n8396), .ZN(n8486) );
  XNOR2_X1 U9312 ( .A(n7587), .B(n8486), .ZN(n7588) );
  OAI222_X1 U9313 ( .A1(n8788), .A2(n8791), .B1(n8790), .B2(n7589), .C1(n7588), 
        .C2(n8786), .ZN(n8866) );
  AOI21_X1 U9314 ( .B1(n7591), .B2(n7590), .A(n8866), .ZN(n7595) );
  XOR2_X1 U9315 ( .A(n7592), .B(n8486), .Z(n8867) );
  OAI22_X1 U9316 ( .A1(n9824), .A2(n5942), .B1(n8151), .B2(n8679), .ZN(n7593)
         );
  AOI21_X1 U9317 ( .B1(n8867), .B2(n8801), .A(n7593), .ZN(n7594) );
  OAI21_X1 U9318 ( .B1(n7595), .B2(n8803), .A(n7594), .ZN(P2_U3219) );
  NOR2_X1 U9319 ( .A1(n7596), .A2(n4733), .ZN(n7601) );
  AOI21_X1 U9320 ( .B1(n7599), .B2(n7598), .A(n7597), .ZN(n7600) );
  OAI21_X1 U9321 ( .B1(n7601), .B2(n7600), .A(n9102), .ZN(n7607) );
  OAI22_X1 U9322 ( .A1(n7603), .A2(n9095), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7602), .ZN(n7604) );
  AOI21_X1 U9323 ( .B1(n7605), .B2(n9109), .A(n7604), .ZN(n7606) );
  OAI211_X1 U9324 ( .C1(n7608), .C2(n9113), .A(n7607), .B(n7606), .ZN(P1_U3236) );
  AOI21_X1 U9325 ( .B1(n8277), .B2(n8532), .A(n7609), .ZN(n7612) );
  INV_X1 U9326 ( .A(n7994), .ZN(n7610) );
  NAND2_X1 U9327 ( .A1(n8281), .A2(n7610), .ZN(n7611) );
  OAI211_X1 U9328 ( .C1(n7992), .C2(n8279), .A(n7612), .B(n7611), .ZN(n7619)
         );
  INV_X1 U9329 ( .A(n7613), .ZN(n7617) );
  AOI21_X1 U9330 ( .B1(n7505), .B2(n7614), .A(n7615), .ZN(n7616) );
  NOR3_X1 U9331 ( .A1(n7617), .A2(n7616), .A3(n8271), .ZN(n7618) );
  AOI211_X1 U9332 ( .C1(n7996), .C2(n8269), .A(n7619), .B(n7618), .ZN(n7620)
         );
  INV_X1 U9333 ( .A(n7620), .ZN(P2_U3176) );
  XOR2_X1 U9334 ( .A(n7621), .B(n7622), .Z(n7630) );
  NAND2_X1 U9335 ( .A1(n9109), .A2(n7623), .ZN(n7624) );
  OAI211_X1 U9336 ( .C1(n7626), .C2(n9095), .A(n7625), .B(n7624), .ZN(n7627)
         );
  AOI21_X1 U9337 ( .B1(n7628), .B2(n9628), .A(n7627), .ZN(n7629) );
  OAI21_X1 U9338 ( .B1(n7630), .B2(n9623), .A(n7629), .ZN(P1_U3224) );
  INV_X1 U9339 ( .A(n9066), .ZN(n7641) );
  INV_X1 U9340 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n7636) );
  OAI211_X1 U9341 ( .C1(n7633), .C2(n9496), .A(n7632), .B(n7631), .ZN(n7634)
         );
  AOI21_X1 U9342 ( .B1(n7635), .B2(n9734), .A(n7634), .ZN(n7638) );
  MUX2_X1 U9343 ( .A(n7636), .B(n7638), .S(n9757), .Z(n7637) );
  OAI21_X1 U9344 ( .B1(n7641), .B2(n9524), .A(n7637), .ZN(P1_U3535) );
  INV_X1 U9345 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n7639) );
  MUX2_X1 U9346 ( .A(n7639), .B(n7638), .S(n9749), .Z(n7640) );
  OAI21_X1 U9347 ( .B1(n7641), .B2(n9576), .A(n7640), .ZN(P1_U3492) );
  INV_X1 U9348 ( .A(n7642), .ZN(n8138) );
  OAI222_X1 U9349 ( .A1(n9591), .A2(n8138), .B1(P1_U3086), .B2(n7644), .C1(
        n7643), .C2(n9588), .ZN(P1_U3331) );
  AOI21_X1 U9350 ( .B1(n7647), .B2(n7646), .A(n7645), .ZN(n7663) );
  NOR2_X1 U9351 ( .A1(n7649), .A2(n7648), .ZN(n7651) );
  XNOR2_X1 U9352 ( .A(n7651), .B(n7650), .ZN(n7661) );
  INV_X1 U9353 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7655) );
  AOI21_X1 U9354 ( .B1(n9772), .B2(n7653), .A(n7652), .ZN(n7654) );
  OAI21_X1 U9355 ( .B1(n8628), .B2(n7655), .A(n7654), .ZN(n7660) );
  AOI21_X1 U9356 ( .B1(n4452), .B2(n7657), .A(n7656), .ZN(n7658) );
  NOR2_X1 U9357 ( .A1(n7658), .A2(n9810), .ZN(n7659) );
  AOI211_X1 U9358 ( .C1(n9807), .C2(n7661), .A(n7660), .B(n7659), .ZN(n7662)
         );
  OAI21_X1 U9359 ( .B1(n7663), .B2(n9803), .A(n7662), .ZN(P2_U3194) );
  XOR2_X1 U9360 ( .A(n7863), .B(n7664), .Z(n9517) );
  NAND2_X1 U9361 ( .A1(n9410), .A2(n7767), .ZN(n7665) );
  XNOR2_X1 U9362 ( .A(n7665), .B(n7863), .ZN(n7666) );
  OAI222_X1 U9363 ( .A1(n9414), .A2(n9373), .B1(n7666), .B2(n9496), .C1(n9412), 
        .C2(n9107), .ZN(n9512) );
  AOI211_X1 U9364 ( .C1(n9514), .C2(n9421), .A(n9422), .B(n9396), .ZN(n9513)
         );
  NAND2_X1 U9365 ( .A1(n9513), .A2(n9431), .ZN(n7668) );
  AOI22_X1 U9366 ( .A1(n9433), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n9110), .B2(
        n9426), .ZN(n7667) );
  OAI211_X1 U9367 ( .C1(n9114), .C2(n9429), .A(n7668), .B(n7667), .ZN(n7669)
         );
  AOI21_X1 U9368 ( .B1(n9381), .B2(n9512), .A(n7669), .ZN(n7670) );
  OAI21_X1 U9369 ( .B1(n9517), .B2(n9404), .A(n7670), .ZN(P1_U3278) );
  INV_X1 U9370 ( .A(n7671), .ZN(n7672) );
  AOI21_X2 U9371 ( .B1(n7674), .B2(n7673), .A(n4948), .ZN(n7677) );
  XNOR2_X1 U9372 ( .A(n8388), .B(n8124), .ZN(n7675) );
  NOR2_X1 U9373 ( .A1(n7675), .A2(n8529), .ZN(n8093) );
  AOI21_X1 U9374 ( .B1(n7675), .B2(n8529), .A(n8093), .ZN(n7676) );
  OAI21_X1 U9375 ( .B1(n7677), .B2(n7676), .A(n8094), .ZN(n7678) );
  NAND2_X1 U9376 ( .A1(n7678), .A2(n8273), .ZN(n7683) );
  OR2_X1 U9377 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6208), .ZN(n8550) );
  OAI21_X1 U9378 ( .B1(n8279), .B2(n8096), .A(n8550), .ZN(n7681) );
  NOR2_X1 U9379 ( .A1(n8267), .A2(n7679), .ZN(n7680) );
  AOI211_X1 U9380 ( .C1(n8277), .C2(n8530), .A(n7681), .B(n7680), .ZN(n7682)
         );
  OAI211_X1 U9381 ( .C1(n8944), .C2(n8285), .A(n7683), .B(n7682), .ZN(P2_U3174) );
  INV_X1 U9382 ( .A(n7684), .ZN(n8053) );
  OAI222_X1 U9383 ( .A1(n9591), .A2(n8053), .B1(P1_U3086), .B2(n7686), .C1(
        n7685), .C2(n9588), .ZN(P1_U3330) );
  INV_X1 U9384 ( .A(n7687), .ZN(n7691) );
  OAI222_X1 U9385 ( .A1(n9591), .A2(n7691), .B1(P1_U3086), .B2(n7689), .C1(
        n7688), .C2(n9588), .ZN(P1_U3329) );
  OAI222_X1 U9386 ( .A1(n7692), .A2(P2_U3151), .B1(n8960), .B2(n7691), .C1(
        n7690), .C2(n8956), .ZN(P2_U3269) );
  INV_X1 U9387 ( .A(n7693), .ZN(n8959) );
  OAI222_X1 U9388 ( .A1(n9591), .A2(n8959), .B1(P1_U3086), .B2(n6515), .C1(
        n7694), .C2(n9588), .ZN(P1_U3328) );
  INV_X1 U9389 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7696) );
  OAI222_X1 U9390 ( .A1(n9588), .A2(n7696), .B1(n9591), .B2(n7695), .C1(
        P1_U3086), .C2(n7928), .ZN(P1_U3336) );
  NAND2_X1 U9391 ( .A1(n7697), .A2(n9824), .ZN(n7703) );
  INV_X1 U9392 ( .A(n7698), .ZN(n7699) );
  NAND2_X1 U9393 ( .A1(n9821), .A2(n7699), .ZN(n8634) );
  OAI21_X1 U9394 ( .B1(n9824), .B2(n7700), .A(n8634), .ZN(n7701) );
  AOI21_X1 U9395 ( .B1(n8307), .B2(n9819), .A(n7701), .ZN(n7702) );
  OAI211_X1 U9396 ( .C1(n6420), .C2(n7704), .A(n7703), .B(n7702), .ZN(P2_U3204) );
  INV_X1 U9397 ( .A(n6351), .ZN(n7706) );
  OAI222_X1 U9398 ( .A1(n9591), .A2(n7706), .B1(n5726), .B2(P1_U3086), .C1(
        n7705), .C2(n9588), .ZN(P1_U3327) );
  MUX2_X1 U9399 ( .A(n9253), .B(n7889), .S(n7919), .Z(n7797) );
  INV_X1 U9400 ( .A(n7770), .ZN(n7763) );
  NAND2_X1 U9401 ( .A1(n7707), .A2(n7937), .ZN(n7710) );
  NAND2_X1 U9402 ( .A1(n7708), .A2(n7941), .ZN(n7709) );
  INV_X1 U9403 ( .A(n7919), .ZN(n7838) );
  MUX2_X1 U9404 ( .A(n7710), .B(n7709), .S(n7838), .Z(n7720) );
  MUX2_X1 U9405 ( .A(n7937), .B(n7941), .S(n7919), .Z(n7712) );
  AND2_X1 U9406 ( .A1(n7712), .A2(n7711), .ZN(n7719) );
  NAND2_X1 U9407 ( .A1(n7714), .A2(n7713), .ZN(n7943) );
  NAND2_X1 U9408 ( .A1(n7943), .A2(n7919), .ZN(n7717) );
  OR2_X1 U9409 ( .A1(n7940), .A2(n7919), .ZN(n7715) );
  NAND4_X1 U9410 ( .A1(n7717), .A2(n7716), .A3(n7944), .A4(n7715), .ZN(n7718)
         );
  AOI21_X1 U9411 ( .B1(n7720), .B2(n7719), .A(n7718), .ZN(n7739) );
  NAND4_X1 U9412 ( .A1(n7721), .A2(n9137), .A3(n5744), .A4(n7919), .ZN(n7732)
         );
  OAI21_X1 U9413 ( .B1(n7722), .B2(n7838), .A(n4576), .ZN(n7726) );
  NAND2_X1 U9414 ( .A1(n7722), .A2(n7838), .ZN(n7724) );
  NAND2_X1 U9415 ( .A1(n7724), .A2(n7723), .ZN(n7725) );
  NAND2_X1 U9416 ( .A1(n7726), .A2(n7725), .ZN(n7731) );
  NAND4_X1 U9417 ( .A1(n7729), .A2(n7728), .A3(n7838), .A4(n7727), .ZN(n7730)
         );
  NAND4_X1 U9418 ( .A1(n7733), .A2(n7732), .A3(n7731), .A4(n7730), .ZN(n7738)
         );
  INV_X1 U9419 ( .A(n7734), .ZN(n7735) );
  MUX2_X1 U9420 ( .A(n7736), .B(n7735), .S(n7919), .Z(n7737) );
  OAI21_X1 U9421 ( .B1(n7739), .B2(n7738), .A(n7737), .ZN(n7744) );
  AND2_X1 U9422 ( .A1(n7745), .A2(n7740), .ZN(n7741) );
  MUX2_X1 U9423 ( .A(n7742), .B(n7741), .S(n7838), .Z(n7743) );
  NAND2_X1 U9424 ( .A1(n7744), .A2(n7743), .ZN(n7751) );
  NAND2_X1 U9425 ( .A1(n7751), .A2(n7745), .ZN(n7747) );
  NAND2_X1 U9426 ( .A1(n7753), .A2(n7746), .ZN(n7952) );
  AOI21_X1 U9427 ( .B1(n7747), .B2(n7949), .A(n7952), .ZN(n7748) );
  NAND2_X1 U9428 ( .A1(n7756), .A2(n7752), .ZN(n7957) );
  OAI21_X1 U9429 ( .B1(n7748), .B2(n7957), .A(n7955), .ZN(n7759) );
  AOI21_X1 U9430 ( .B1(n7751), .B2(n7750), .A(n7749), .ZN(n7755) );
  NAND2_X1 U9431 ( .A1(n7752), .A2(n7949), .ZN(n7754) );
  OAI211_X1 U9432 ( .C1(n7755), .C2(n7754), .A(n7955), .B(n7753), .ZN(n7757)
         );
  NAND2_X1 U9433 ( .A1(n7757), .A2(n7756), .ZN(n7758) );
  MUX2_X1 U9434 ( .A(n7759), .B(n7758), .S(n7838), .Z(n7765) );
  AND2_X1 U9435 ( .A1(n7761), .A2(n7760), .ZN(n7961) );
  NAND2_X1 U9436 ( .A1(n7770), .A2(n7762), .ZN(n7965) );
  INV_X1 U9437 ( .A(n7961), .ZN(n7764) );
  AOI21_X1 U9438 ( .B1(n7765), .B2(n7956), .A(n7764), .ZN(n7774) );
  NAND2_X1 U9439 ( .A1(n9370), .A2(n7766), .ZN(n7959) );
  NAND2_X1 U9440 ( .A1(n7767), .A2(n7838), .ZN(n7768) );
  OR2_X1 U9441 ( .A1(n7959), .A2(n7768), .ZN(n7773) );
  NOR2_X1 U9442 ( .A1(n9514), .A2(n7919), .ZN(n7769) );
  AOI21_X1 U9443 ( .B1(n7959), .B2(n7770), .A(n7769), .ZN(n7772) );
  AOI21_X1 U9444 ( .B1(n9370), .B2(n9392), .A(n7919), .ZN(n7771) );
  OAI22_X1 U9445 ( .A1(n7774), .A2(n7773), .B1(n7772), .B2(n7771), .ZN(n7775)
         );
  NAND2_X1 U9446 ( .A1(n7776), .A2(n9368), .ZN(n7782) );
  AND2_X1 U9447 ( .A1(n7967), .A2(n7777), .ZN(n7930) );
  NAND2_X1 U9448 ( .A1(n7970), .A2(n7781), .ZN(n7778) );
  NAND2_X1 U9449 ( .A1(n9336), .A2(n9343), .ZN(n7784) );
  NAND2_X1 U9450 ( .A1(n7784), .A2(n7970), .ZN(n7779) );
  AOI21_X1 U9451 ( .B1(n7785), .B2(n7966), .A(n7919), .ZN(n7783) );
  AND2_X1 U9452 ( .A1(n7787), .A2(n7784), .ZN(n7884) );
  NAND2_X1 U9453 ( .A1(n9318), .A2(n9123), .ZN(n7885) );
  AND2_X1 U9454 ( .A1(n7885), .A2(n7785), .ZN(n7876) );
  MUX2_X1 U9455 ( .A(n7884), .B(n7876), .S(n7919), .Z(n7786) );
  MUX2_X1 U9456 ( .A(n7787), .B(n7885), .S(n7838), .Z(n7788) );
  NAND2_X1 U9457 ( .A1(n9556), .A2(n9122), .ZN(n7789) );
  NAND2_X1 U9458 ( .A1(n7790), .A2(n7789), .ZN(n7877) );
  AOI22_X1 U9459 ( .A1(n7791), .A2(n9298), .B1(n7838), .B2(n7877), .ZN(n7794)
         );
  AND2_X1 U9460 ( .A1(n9270), .A2(n7792), .ZN(n7888) );
  OR3_X1 U9461 ( .A1(n9294), .A2(n7838), .A3(n7795), .ZN(n7796) );
  NAND2_X1 U9462 ( .A1(n7897), .A2(n7890), .ZN(n7802) );
  AOI21_X1 U9463 ( .B1(n4408), .B2(n7881), .A(n7802), .ZN(n7801) );
  OR2_X1 U9464 ( .A1(n9249), .A2(n7798), .ZN(n7882) );
  INV_X1 U9465 ( .A(n7882), .ZN(n7800) );
  OAI21_X1 U9466 ( .B1(n7801), .B2(n7800), .A(n4387), .ZN(n7810) );
  NAND4_X1 U9467 ( .A1(n8060), .A2(n7838), .A3(n7882), .A4(n7883), .ZN(n7803)
         );
  NAND3_X1 U9468 ( .A1(n7896), .A2(n7838), .A3(n8060), .ZN(n7805) );
  OAI21_X1 U9469 ( .B1(n7838), .B2(n8060), .A(n7805), .ZN(n7808) );
  INV_X1 U9470 ( .A(n7883), .ZN(n7806) );
  INV_X1 U9471 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n9589) );
  OR2_X1 U9472 ( .A1(n5145), .A2(n9589), .ZN(n7811) );
  OR2_X2 U9473 ( .A1(n4351), .A2(n7812), .ZN(n7904) );
  NAND2_X1 U9474 ( .A1(n4351), .A2(n7812), .ZN(n7908) );
  OAI21_X1 U9475 ( .B1(n7814), .B2(n8064), .A(n7813), .ZN(n7839) );
  INV_X1 U9476 ( .A(n7815), .ZN(n7816) );
  MUX2_X1 U9477 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n7825), .Z(n7822) );
  XNOR2_X1 U9478 ( .A(n7822), .B(SI_30_), .ZN(n7823) );
  NAND2_X1 U9479 ( .A1(n8289), .A2(n7830), .ZN(n7821) );
  INV_X1 U9480 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n7988) );
  OR2_X1 U9481 ( .A1(n5145), .A2(n7988), .ZN(n7820) );
  OAI22_X1 U9482 ( .A1(n7824), .A2(n7823), .B1(SI_30_), .B2(n7822), .ZN(n7829)
         );
  MUX2_X1 U9483 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n7825), .Z(n7827) );
  INV_X1 U9484 ( .A(SI_31_), .ZN(n7826) );
  XNOR2_X1 U9485 ( .A(n7827), .B(n7826), .ZN(n7828) );
  XNOR2_X1 U9486 ( .A(n7829), .B(n7828), .ZN(n8945) );
  NAND2_X1 U9487 ( .A1(n8945), .A2(n7830), .ZN(n7833) );
  INV_X1 U9488 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n7831) );
  OR2_X1 U9489 ( .A1(n5145), .A2(n7831), .ZN(n7832) );
  INV_X1 U9490 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n7836) );
  NAND2_X1 U9491 ( .A1(n4355), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n7835) );
  NAND2_X1 U9492 ( .A1(n4357), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n7834) );
  OAI211_X1 U9493 ( .C1(n7837), .C2(n7836), .A(n7835), .B(n7834), .ZN(n9115)
         );
  NAND2_X1 U9494 ( .A1(n9205), .A2(n9115), .ZN(n7910) );
  NAND2_X1 U9495 ( .A1(n9203), .A2(n7840), .ZN(n7920) );
  OAI21_X1 U9496 ( .B1(n7842), .B2(n7841), .A(n7924), .ZN(n7874) );
  INV_X1 U9497 ( .A(n9115), .ZN(n7844) );
  OR2_X1 U9498 ( .A1(n9202), .A2(n7844), .ZN(n7843) );
  NAND2_X1 U9499 ( .A1(n7920), .A2(n7843), .ZN(n7976) );
  NAND2_X1 U9500 ( .A1(n9202), .A2(n7844), .ZN(n7909) );
  INV_X1 U9501 ( .A(n9254), .ZN(n7870) );
  INV_X1 U9502 ( .A(n9385), .ZN(n9384) );
  INV_X1 U9503 ( .A(n7845), .ZN(n7862) );
  NOR2_X1 U9504 ( .A1(n7846), .A2(n7924), .ZN(n7851) );
  NOR2_X1 U9505 ( .A1(n7847), .A2(n6665), .ZN(n7850) );
  NAND4_X1 U9506 ( .A1(n7851), .A2(n7850), .A3(n7849), .A4(n7848), .ZN(n7853)
         );
  NOR2_X1 U9507 ( .A1(n7853), .A2(n7852), .ZN(n7857) );
  INV_X1 U9508 ( .A(n7950), .ZN(n7856) );
  NAND4_X1 U9509 ( .A1(n7857), .A2(n7856), .A3(n7855), .A4(n7854), .ZN(n7860)
         );
  NOR3_X1 U9510 ( .A1(n7860), .A2(n7859), .A3(n7858), .ZN(n7861) );
  NAND3_X1 U9511 ( .A1(n4826), .A2(n7862), .A3(n7861), .ZN(n7864) );
  NOR2_X1 U9512 ( .A1(n7864), .A2(n7863), .ZN(n7865) );
  NAND4_X1 U9513 ( .A1(n9353), .A2(n9368), .A3(n9384), .A4(n7865), .ZN(n7866)
         );
  NAND4_X1 U9514 ( .A1(n9288), .A2(n4396), .A3(n9298), .A4(n9320), .ZN(n7867)
         );
  NOR2_X1 U9515 ( .A1(n7868), .A2(n7867), .ZN(n7869) );
  AND4_X1 U9516 ( .A1(n9225), .A2(n7870), .A3(n7869), .A4(n9242), .ZN(n7871)
         );
  NAND4_X1 U9517 ( .A1(n7909), .A2(n8058), .A3(n7872), .A4(n7871), .ZN(n7873)
         );
  INV_X1 U9518 ( .A(n7876), .ZN(n7899) );
  NAND2_X1 U9519 ( .A1(n7877), .A2(n9270), .ZN(n7878) );
  NAND2_X1 U9520 ( .A1(n9253), .A2(n7878), .ZN(n7879) );
  NAND2_X1 U9521 ( .A1(n7879), .A2(n7889), .ZN(n7880) );
  AND2_X1 U9522 ( .A1(n7881), .A2(n7880), .ZN(n7893) );
  INV_X1 U9523 ( .A(n7893), .ZN(n7898) );
  NAND2_X1 U9524 ( .A1(n7883), .A2(n7882), .ZN(n7901) );
  INV_X1 U9525 ( .A(n7884), .ZN(n7886) );
  NAND2_X1 U9526 ( .A1(n7886), .A2(n7885), .ZN(n7887) );
  NAND3_X1 U9527 ( .A1(n7889), .A2(n7888), .A3(n7887), .ZN(n7892) );
  INV_X1 U9528 ( .A(n7890), .ZN(n7891) );
  NOR2_X1 U9529 ( .A1(n7901), .A2(n7894), .ZN(n7895) );
  OR2_X1 U9530 ( .A1(n7896), .A2(n7895), .ZN(n7900) );
  OAI21_X1 U9531 ( .B1(n7899), .B2(n7898), .A(n7971), .ZN(n7905) );
  INV_X1 U9532 ( .A(n7900), .ZN(n7902) );
  NAND2_X1 U9533 ( .A1(n7902), .A2(n7901), .ZN(n7903) );
  NAND4_X1 U9534 ( .A1(n7905), .A2(n7904), .A3(n8060), .A4(n7903), .ZN(n7929)
         );
  INV_X1 U9535 ( .A(n7971), .ZN(n7906) );
  NOR2_X1 U9536 ( .A1(n7906), .A2(n9328), .ZN(n7907) );
  OAI22_X1 U9537 ( .A1(n7929), .A2(n7907), .B1(n9532), .B2(n9205), .ZN(n7911)
         );
  NAND2_X1 U9538 ( .A1(n7909), .A2(n7908), .ZN(n7972) );
  OAI22_X1 U9539 ( .A1(n7911), .A2(n7972), .B1(n9202), .B2(n7910), .ZN(n7913)
         );
  AOI211_X1 U9540 ( .C1(n7913), .C2(n7975), .A(n7912), .B(n4504), .ZN(n7916)
         );
  INV_X1 U9541 ( .A(n7914), .ZN(n7915) );
  OAI22_X1 U9542 ( .A1(n7921), .A2(n5712), .B1(n7920), .B2(n7919), .ZN(n7925)
         );
  NAND2_X1 U9543 ( .A1(n7922), .A2(n7875), .ZN(n7923) );
  NAND3_X1 U9544 ( .A1(n7925), .A2(n7924), .A3(n7923), .ZN(n7926) );
  NOR2_X1 U9545 ( .A1(n7928), .A2(n7982), .ZN(n7980) );
  INV_X1 U9546 ( .A(n5711), .ZN(n7979) );
  INV_X1 U9547 ( .A(n7929), .ZN(n7974) );
  INV_X1 U9548 ( .A(n7930), .ZN(n7964) );
  AOI21_X1 U9549 ( .B1(n5737), .B2(n5821), .A(n7931), .ZN(n7935) );
  INV_X1 U9550 ( .A(n7932), .ZN(n7934) );
  AOI21_X1 U9551 ( .B1(n7935), .B2(n7934), .A(n7933), .ZN(n7939) );
  INV_X1 U9552 ( .A(n7936), .ZN(n7938) );
  OAI21_X1 U9553 ( .B1(n7939), .B2(n7938), .A(n7937), .ZN(n7942) );
  NAND3_X1 U9554 ( .A1(n7942), .A2(n7941), .A3(n7940), .ZN(n7947) );
  INV_X1 U9555 ( .A(n7943), .ZN(n7946) );
  INV_X1 U9556 ( .A(n7944), .ZN(n7945) );
  AOI21_X1 U9557 ( .B1(n7947), .B2(n7946), .A(n7945), .ZN(n7951) );
  OAI211_X1 U9558 ( .C1(n7951), .C2(n7950), .A(n7949), .B(n7948), .ZN(n7954)
         );
  INV_X1 U9559 ( .A(n7952), .ZN(n7953) );
  AND2_X1 U9560 ( .A1(n7954), .A2(n7953), .ZN(n7958) );
  OAI211_X1 U9561 ( .C1(n7958), .C2(n7957), .A(n7956), .B(n7955), .ZN(n7962)
         );
  AOI211_X1 U9562 ( .C1(n7962), .C2(n7961), .A(n7960), .B(n7959), .ZN(n7963)
         );
  AOI211_X1 U9563 ( .C1(n7965), .C2(n9370), .A(n7964), .B(n7963), .ZN(n7968)
         );
  OAI211_X1 U9564 ( .C1(n7968), .C2(n4449), .A(n7967), .B(n7966), .ZN(n7969)
         );
  NAND3_X1 U9565 ( .A1(n7971), .A2(n7970), .A3(n7969), .ZN(n7973) );
  AOI21_X1 U9566 ( .B1(n7974), .B2(n7973), .A(n7972), .ZN(n7977) );
  OAI21_X1 U9567 ( .B1(n7977), .B2(n7976), .A(n7975), .ZN(n7978) );
  MUX2_X1 U9568 ( .A(n7980), .B(n7979), .S(n7978), .Z(n7981) );
  NAND3_X1 U9569 ( .A1(n7983), .A2(n9393), .A3(n9154), .ZN(n7984) );
  OAI211_X1 U9570 ( .C1(n5712), .C2(n7986), .A(n7984), .B(P1_B_REG_SCAN_IN), 
        .ZN(n7985) );
  INV_X1 U9571 ( .A(n8289), .ZN(n8139) );
  OAI222_X1 U9572 ( .A1(n9588), .A2(n7988), .B1(n9591), .B2(n8139), .C1(
        P1_U3086), .C2(n7987), .ZN(P1_U3325) );
  XNOR2_X1 U9573 ( .A(n7989), .B(n8465), .ZN(n9862) );
  XNOR2_X1 U9574 ( .A(n7990), .B(n8465), .ZN(n7991) );
  OAI222_X1 U9575 ( .A1(n8790), .A2(n7993), .B1(n8788), .B2(n7992), .C1(n8786), 
        .C2(n7991), .ZN(n9864) );
  NAND2_X1 U9576 ( .A1(n9864), .A2(n9824), .ZN(n7998) );
  OAI22_X1 U9577 ( .A1(n9824), .A2(n7474), .B1(n7994), .B2(n8679), .ZN(n7995)
         );
  AOI21_X1 U9578 ( .B1(n7996), .B2(n9819), .A(n7995), .ZN(n7997) );
  OAI211_X1 U9579 ( .C1(n9862), .C2(n8673), .A(n7998), .B(n7997), .ZN(P2_U3222) );
  INV_X1 U9580 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n8000) );
  XNOR2_X1 U9581 ( .A(n9700), .B(n8000), .ZN(n9696) );
  NAND2_X1 U9582 ( .A1(n9653), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n8001) );
  OAI21_X1 U9583 ( .B1(n9653), .B2(P1_REG2_REG_13__SCAN_IN), .A(n8001), .ZN(
        n9649) );
  OAI21_X1 U9584 ( .B1(n8014), .B2(P1_REG2_REG_12__SCAN_IN), .A(n8002), .ZN(
        n9650) );
  NOR2_X1 U9585 ( .A1(n9649), .A2(n9650), .ZN(n9648) );
  NAND2_X1 U9586 ( .A1(n9665), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n8003) );
  OAI21_X1 U9587 ( .B1(n9665), .B2(P1_REG2_REG_14__SCAN_IN), .A(n8003), .ZN(
        n9658) );
  NOR2_X1 U9588 ( .A1(n9659), .A2(n9658), .ZN(n9657) );
  NOR2_X1 U9589 ( .A1(n8004), .A2(n8016), .ZN(n8005) );
  INV_X1 U9590 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9674) );
  XOR2_X1 U9591 ( .A(n8004), .B(n9678), .Z(n9675) );
  NOR2_X1 U9592 ( .A1(n9674), .A2(n9675), .ZN(n9673) );
  NAND2_X1 U9593 ( .A1(n8012), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n8006) );
  OAI21_X1 U9594 ( .B1(n8012), .B2(P1_REG2_REG_16__SCAN_IN), .A(n8006), .ZN(
        n9688) );
  NOR2_X1 U9595 ( .A1(n9689), .A2(n9688), .ZN(n9687) );
  NOR2_X1 U9596 ( .A1(n9700), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n8007) );
  AOI21_X1 U9597 ( .B1(n9696), .B2(n9695), .A(n8007), .ZN(n9709) );
  OR2_X1 U9598 ( .A1(n9706), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n8008) );
  NAND2_X1 U9599 ( .A1(n9706), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n8009) );
  AND2_X1 U9600 ( .A1(n8008), .A2(n8009), .ZN(n9710) );
  NAND2_X1 U9601 ( .A1(n9709), .A2(n9710), .ZN(n9707) );
  NAND2_X1 U9602 ( .A1(n9707), .A2(n8009), .ZN(n8010) );
  XNOR2_X1 U9603 ( .A(n8010), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n8025) );
  INV_X1 U9604 ( .A(n8025), .ZN(n8024) );
  INV_X1 U9605 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n8011) );
  XNOR2_X1 U9606 ( .A(n9700), .B(n8011), .ZN(n9698) );
  OR2_X1 U9607 ( .A1(n8012), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n8018) );
  INV_X1 U9608 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9510) );
  XNOR2_X1 U9609 ( .A(n8012), .B(n9510), .ZN(n9683) );
  XNOR2_X1 U9610 ( .A(n9653), .B(P1_REG1_REG_13__SCAN_IN), .ZN(n9646) );
  OAI21_X1 U9611 ( .B1(P1_REG1_REG_12__SCAN_IN), .B2(n8014), .A(n8013), .ZN(
        n9647) );
  NOR2_X1 U9612 ( .A1(n9646), .A2(n9647), .ZN(n9645) );
  AOI21_X1 U9613 ( .B1(n9653), .B2(P1_REG1_REG_13__SCAN_IN), .A(n9645), .ZN(
        n9662) );
  XNOR2_X1 U9614 ( .A(n9665), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n9661) );
  NOR2_X1 U9615 ( .A1(n9662), .A2(n9661), .ZN(n9660) );
  AOI21_X1 U9616 ( .B1(P1_REG1_REG_14__SCAN_IN), .B2(n9665), .A(n9660), .ZN(
        n8015) );
  NOR2_X1 U9617 ( .A1(n8015), .A2(n8016), .ZN(n8017) );
  INV_X1 U9618 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9671) );
  XNOR2_X1 U9619 ( .A(n8016), .B(n8015), .ZN(n9672) );
  NOR2_X1 U9620 ( .A1(n9671), .A2(n9672), .ZN(n9670) );
  NOR2_X1 U9621 ( .A1(n8017), .A2(n9670), .ZN(n9684) );
  NAND2_X1 U9622 ( .A1(n9683), .A2(n9684), .ZN(n9682) );
  NAND2_X1 U9623 ( .A1(n8018), .A2(n9682), .ZN(n9697) );
  NOR2_X1 U9624 ( .A1(n9700), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n8019) );
  AOI21_X1 U9625 ( .B1(n9698), .B2(n9697), .A(n8019), .ZN(n9714) );
  OR2_X1 U9626 ( .A1(n9706), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n8020) );
  NAND2_X1 U9627 ( .A1(n9706), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n8021) );
  AND2_X1 U9628 ( .A1(n8020), .A2(n8021), .ZN(n9713) );
  NAND2_X1 U9629 ( .A1(n9714), .A2(n9713), .ZN(n9711) );
  NAND2_X1 U9630 ( .A1(n9711), .A2(n8021), .ZN(n8022) );
  XNOR2_X1 U9631 ( .A(n8022), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n8026) );
  NAND2_X1 U9632 ( .A1(n9712), .A2(n8026), .ZN(n8023) );
  OAI211_X1 U9633 ( .C1(n9686), .C2(n8024), .A(n8023), .B(n9718), .ZN(n8028)
         );
  OAI22_X1 U9634 ( .A1(n9669), .A2(n8026), .B1(n8025), .B2(n9686), .ZN(n8027)
         );
  NAND2_X1 U9635 ( .A1(P1_REG3_REG_19__SCAN_IN), .A2(P1_U3086), .ZN(n8029) );
  NAND2_X1 U9636 ( .A1(n8055), .A2(n8030), .ZN(n8033) );
  OR2_X1 U9637 ( .A1(n8054), .A2(n8031), .ZN(n8032) );
  NAND2_X1 U9638 ( .A1(n8033), .A2(n8032), .ZN(n8035) );
  XNOR2_X1 U9639 ( .A(n8035), .B(n8034), .ZN(n8039) );
  NAND2_X1 U9640 ( .A1(n8055), .A2(n8036), .ZN(n8037) );
  OAI21_X1 U9641 ( .B1(n8054), .B2(n5173), .A(n8037), .ZN(n8038) );
  XNOR2_X1 U9642 ( .A(n8039), .B(n8038), .ZN(n8040) );
  INV_X1 U9643 ( .A(n8040), .ZN(n8045) );
  NAND3_X1 U9644 ( .A1(n8045), .A2(n9102), .A3(n8044), .ZN(n8050) );
  NAND3_X1 U9645 ( .A1(n8051), .A2(n9102), .A3(n8040), .ZN(n8049) );
  NAND2_X1 U9646 ( .A1(n9109), .A2(n8081), .ZN(n8042) );
  NAND2_X1 U9647 ( .A1(n8082), .A2(n9618), .ZN(n8041) );
  OAI211_X1 U9648 ( .C1(P1_STATE_REG_SCAN_IN), .C2(n8043), .A(n8042), .B(n8041), .ZN(n8047) );
  NOR3_X1 U9649 ( .A1(n8045), .A2(n9623), .A3(n8044), .ZN(n8046) );
  AOI211_X1 U9650 ( .C1(n8055), .C2(n9628), .A(n8047), .B(n8046), .ZN(n8048)
         );
  OAI211_X1 U9651 ( .C1(n8051), .C2(n8050), .A(n8049), .B(n8048), .ZN(P1_U3220) );
  OAI222_X1 U9652 ( .A1(n6424), .A2(P2_U3151), .B1(n8960), .B2(n8053), .C1(
        n8052), .C2(n8956), .ZN(P2_U3270) );
  INV_X1 U9653 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n8072) );
  INV_X1 U9654 ( .A(n8054), .ZN(n9116) );
  NAND2_X1 U9655 ( .A1(n8055), .A2(n9116), .ZN(n8056) );
  NAND2_X1 U9656 ( .A1(n8057), .A2(n8056), .ZN(n8059) );
  XNOR2_X2 U9657 ( .A(n8059), .B(n8058), .ZN(n9214) );
  NAND2_X1 U9658 ( .A1(n8061), .A2(n8060), .ZN(n8063) );
  NAND2_X1 U9659 ( .A1(n8063), .A2(n8062), .ZN(n8065) );
  XNOR2_X1 U9660 ( .A(n8065), .B(n8064), .ZN(n9223) );
  NAND2_X1 U9661 ( .A1(n9154), .A2(P1_B_REG_SCAN_IN), .ZN(n8066) );
  AND2_X1 U9662 ( .A1(n9390), .A2(n8066), .ZN(n9204) );
  AOI22_X1 U9663 ( .A1(n9116), .A2(n9393), .B1(n9115), .B2(n9204), .ZN(n9217)
         );
  INV_X1 U9664 ( .A(n4351), .ZN(n8070) );
  OAI211_X1 U9665 ( .C1(n8070), .C2(n8069), .A(n9477), .B(n9209), .ZN(n9218)
         );
  OAI211_X1 U9666 ( .C1(n9223), .C2(n9496), .A(n9217), .B(n9218), .ZN(n8071)
         );
  AOI21_X1 U9667 ( .B1(n9214), .B2(n9734), .A(n8071), .ZN(n8076) );
  MUX2_X1 U9668 ( .A(n8072), .B(n8076), .S(n9757), .Z(n8075) );
  NAND2_X1 U9669 ( .A1(n4351), .A2(n8073), .ZN(n8074) );
  NAND2_X1 U9670 ( .A1(n8075), .A2(n8074), .ZN(P1_U3551) );
  INV_X1 U9671 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n8077) );
  MUX2_X1 U9672 ( .A(n8077), .B(n8076), .S(n9749), .Z(n8080) );
  NAND2_X1 U9673 ( .A1(n4351), .A2(n8078), .ZN(n8079) );
  NAND2_X1 U9674 ( .A1(n8080), .A2(n8079), .ZN(P1_U3519) );
  AOI22_X1 U9675 ( .A1(n9433), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n8081), .B2(
        n9426), .ZN(n8084) );
  NAND2_X1 U9676 ( .A1(n8082), .A2(n9381), .ZN(n8083) );
  OAI211_X1 U9677 ( .C1(n8085), .C2(n9429), .A(n8084), .B(n8083), .ZN(n8086)
         );
  AOI21_X1 U9678 ( .B1(n8087), .B2(n9431), .A(n8086), .ZN(n8091) );
  NAND2_X1 U9679 ( .A1(n8089), .A2(n8088), .ZN(n8090) );
  OAI211_X1 U9680 ( .C1(n8092), .C2(n9404), .A(n8091), .B(n8090), .ZN(P1_U3265) );
  INV_X1 U9681 ( .A(n8093), .ZN(n8147) );
  XNOR2_X1 U9682 ( .A(n8938), .B(n4353), .ZN(n8095) );
  XNOR2_X1 U9683 ( .A(n8095), .B(n8528), .ZN(n8148) );
  INV_X1 U9684 ( .A(n8095), .ZN(n8097) );
  XNOR2_X1 U9685 ( .A(n8098), .B(n4353), .ZN(n8099) );
  XNOR2_X1 U9686 ( .A(n8099), .B(n8527), .ZN(n8275) );
  OR2_X1 U9687 ( .A1(n8099), .A2(n8791), .ZN(n8100) );
  NAND2_X1 U9688 ( .A1(n8274), .A2(n8100), .ZN(n8191) );
  XNOR2_X1 U9689 ( .A(n8857), .B(n4353), .ZN(n8101) );
  NAND2_X1 U9690 ( .A1(n8101), .A2(n8777), .ZN(n8187) );
  NOR2_X1 U9691 ( .A1(n8101), .A2(n8777), .ZN(n8189) );
  AOI21_X2 U9692 ( .B1(n8191), .B2(n8187), .A(n8189), .ZN(n8198) );
  XNOR2_X1 U9693 ( .A(n8929), .B(n4353), .ZN(n8102) );
  XNOR2_X1 U9694 ( .A(n8102), .B(n8789), .ZN(n8197) );
  INV_X1 U9695 ( .A(n8102), .ZN(n8103) );
  AOI21_X1 U9696 ( .B1(n8198), .B2(n8197), .A(n4943), .ZN(n8239) );
  XNOR2_X1 U9697 ( .A(n8243), .B(n4353), .ZN(n8104) );
  XNOR2_X1 U9698 ( .A(n8104), .B(n8776), .ZN(n8238) );
  INV_X1 U9699 ( .A(n8104), .ZN(n8105) );
  XNOR2_X1 U9700 ( .A(n8753), .B(n4353), .ZN(n8106) );
  XNOR2_X1 U9701 ( .A(n8106), .B(n8764), .ZN(n8165) );
  NOR2_X1 U9702 ( .A1(n8164), .A2(n8165), .ZN(n8163) );
  XNOR2_X1 U9703 ( .A(n8107), .B(n4353), .ZN(n8108) );
  XOR2_X1 U9704 ( .A(n8722), .B(n8108), .Z(n8213) );
  INV_X1 U9705 ( .A(n8108), .ZN(n8109) );
  XNOR2_X1 U9706 ( .A(n8727), .B(n4353), .ZN(n8110) );
  XNOR2_X1 U9707 ( .A(n8110), .B(n8525), .ZN(n8172) );
  XNOR2_X1 U9708 ( .A(n8225), .B(n4353), .ZN(n8111) );
  XNOR2_X1 U9709 ( .A(n8111), .B(n8721), .ZN(n8221) );
  INV_X1 U9710 ( .A(n8111), .ZN(n8112) );
  INV_X1 U9711 ( .A(n8721), .ZN(n8524) );
  XNOR2_X1 U9712 ( .A(n8908), .B(n4353), .ZN(n8114) );
  NAND2_X1 U9713 ( .A1(n8156), .A2(n8711), .ZN(n8117) );
  INV_X1 U9714 ( .A(n8113), .ZN(n8115) );
  XNOR2_X1 U9715 ( .A(n8904), .B(n4353), .ZN(n8118) );
  INV_X1 U9716 ( .A(n8118), .ZN(n8119) );
  NAND2_X1 U9717 ( .A1(n8119), .A2(n8700), .ZN(n8120) );
  XNOR2_X1 U9718 ( .A(n8900), .B(n4353), .ZN(n8122) );
  XNOR2_X1 U9719 ( .A(n8122), .B(n8689), .ZN(n8180) );
  INV_X1 U9720 ( .A(n8122), .ZN(n8123) );
  NAND2_X1 U9721 ( .A1(n8123), .A2(n8689), .ZN(n8258) );
  XNOR2_X1 U9722 ( .A(n8670), .B(n8124), .ZN(n8126) );
  INV_X1 U9723 ( .A(n8126), .ZN(n8125) );
  NAND2_X1 U9724 ( .A1(n8125), .A2(n8678), .ZN(n8260) );
  NAND2_X1 U9725 ( .A1(n8126), .A2(n6337), .ZN(n8259) );
  XNOR2_X1 U9726 ( .A(n8890), .B(n4353), .ZN(n8127) );
  XNOR2_X1 U9727 ( .A(n8643), .B(n4353), .ZN(n8130) );
  XNOR2_X1 U9728 ( .A(n8131), .B(n8130), .ZN(n8136) );
  NOR2_X1 U9729 ( .A1(n8267), .A2(n8641), .ZN(n8134) );
  AOI22_X1 U9730 ( .A1(n8277), .A2(n8664), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n8132) );
  OAI21_X1 U9731 ( .B1(n8638), .B2(n8279), .A(n8132), .ZN(n8133) );
  AOI211_X1 U9732 ( .C1(n8647), .C2(n8269), .A(n8134), .B(n8133), .ZN(n8135)
         );
  OAI21_X1 U9733 ( .B1(n8136), .B2(n8271), .A(n8135), .ZN(P2_U3160) );
  OAI222_X1 U9734 ( .A1(n6422), .A2(P2_U3151), .B1(n8960), .B2(n8138), .C1(
        n8137), .C2(n8956), .ZN(P2_U3271) );
  INV_X1 U9735 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8290) );
  OAI222_X1 U9736 ( .A1(n6062), .A2(P2_U3151), .B1(n8960), .B2(n8139), .C1(
        n8290), .C2(n8956), .ZN(P2_U3265) );
  XNOR2_X1 U9737 ( .A(n8140), .B(n8141), .ZN(n8146) );
  NOR2_X1 U9738 ( .A1(n8267), .A2(n8653), .ZN(n8144) );
  AOI22_X1 U9739 ( .A1(n8277), .A2(n6337), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n8142) );
  OAI21_X1 U9740 ( .B1(n8650), .B2(n8279), .A(n8142), .ZN(n8143) );
  AOI211_X1 U9741 ( .C1(n8890), .C2(n8269), .A(n8144), .B(n8143), .ZN(n8145)
         );
  OAI21_X1 U9742 ( .B1(n8146), .B2(n8271), .A(n8145), .ZN(P2_U3154) );
  AND3_X1 U9743 ( .A1(n8094), .A2(n8148), .A3(n8147), .ZN(n8149) );
  OAI21_X1 U9744 ( .B1(n8150), .B2(n8149), .A(n8273), .ZN(n8155) );
  NAND2_X1 U9745 ( .A1(P2_U3151), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8567) );
  OAI21_X1 U9746 ( .B1(n8279), .B2(n8791), .A(n8567), .ZN(n8153) );
  NOR2_X1 U9747 ( .A1(n8267), .A2(n8151), .ZN(n8152) );
  AOI211_X1 U9748 ( .C1(n8277), .C2(n8529), .A(n8153), .B(n8152), .ZN(n8154)
         );
  OAI211_X1 U9749 ( .C1(n8938), .C2(n8285), .A(n8155), .B(n8154), .ZN(P2_U3155) );
  XNOR2_X1 U9750 ( .A(n8156), .B(n8523), .ZN(n8162) );
  AOI22_X1 U9751 ( .A1(n8277), .A2(n8524), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n8158) );
  NAND2_X1 U9752 ( .A1(n8281), .A2(n8703), .ZN(n8157) );
  OAI211_X1 U9753 ( .C1(n8700), .C2(n8279), .A(n8158), .B(n8157), .ZN(n8159)
         );
  AOI21_X1 U9754 ( .B1(n8160), .B2(n8269), .A(n8159), .ZN(n8161) );
  OAI21_X1 U9755 ( .B1(n8162), .B2(n8271), .A(n8161), .ZN(P2_U3156) );
  AOI211_X1 U9756 ( .C1(n8165), .C2(n8164), .A(n8271), .B(n8163), .ZN(n8166)
         );
  INV_X1 U9757 ( .A(n8166), .ZN(n8171) );
  NAND2_X1 U9758 ( .A1(n8277), .A2(n8746), .ZN(n8168) );
  OAI211_X1 U9759 ( .C1(n8722), .C2(n8279), .A(n8168), .B(n8167), .ZN(n8169)
         );
  AOI21_X1 U9760 ( .B1(n8751), .B2(n8281), .A(n8169), .ZN(n8170) );
  OAI211_X1 U9761 ( .C1(n8753), .C2(n8285), .A(n8171), .B(n8170), .ZN(P2_U3159) );
  XOR2_X1 U9762 ( .A(n8173), .B(n8172), .Z(n8178) );
  INV_X1 U9763 ( .A(n8277), .ZN(n8263) );
  AOI22_X1 U9764 ( .A1(n8265), .A2(n8524), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n8175) );
  NAND2_X1 U9765 ( .A1(n8281), .A2(n8728), .ZN(n8174) );
  OAI211_X1 U9766 ( .C1(n8263), .C2(n8722), .A(n8175), .B(n8174), .ZN(n8176)
         );
  AOI21_X1 U9767 ( .B1(n8727), .B2(n8269), .A(n8176), .ZN(n8177) );
  OAI21_X1 U9768 ( .B1(n8178), .B2(n8271), .A(n8177), .ZN(P2_U3163) );
  XOR2_X1 U9769 ( .A(n8180), .B(n8179), .Z(n8186) );
  INV_X1 U9770 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n10016) );
  OAI22_X1 U9771 ( .A1(n8279), .A2(n8678), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10016), .ZN(n8181) );
  AOI21_X1 U9772 ( .B1(n6315), .B2(n8277), .A(n8181), .ZN(n8182) );
  OAI21_X1 U9773 ( .B1(n8680), .B2(n8267), .A(n8182), .ZN(n8183) );
  AOI21_X1 U9774 ( .B1(n8184), .B2(n8269), .A(n8183), .ZN(n8185) );
  OAI21_X1 U9775 ( .B1(n8186), .B2(n8271), .A(n8185), .ZN(P2_U3165) );
  INV_X1 U9776 ( .A(n8187), .ZN(n8188) );
  NOR2_X1 U9777 ( .A1(n8189), .A2(n8188), .ZN(n8190) );
  XNOR2_X1 U9778 ( .A(n8191), .B(n8190), .ZN(n8196) );
  NAND2_X1 U9779 ( .A1(n8277), .A2(n8527), .ZN(n8192) );
  NAND2_X1 U9780 ( .A1(P2_U3151), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8601) );
  OAI211_X1 U9781 ( .C1(n8789), .C2(n8279), .A(n8192), .B(n8601), .ZN(n8193)
         );
  AOI21_X1 U9782 ( .B1(n8796), .B2(n8281), .A(n8193), .ZN(n8195) );
  NAND2_X1 U9783 ( .A1(n8857), .A2(n8269), .ZN(n8194) );
  OAI211_X1 U9784 ( .C1(n8196), .C2(n8271), .A(n8195), .B(n8194), .ZN(P2_U3166) );
  XOR2_X1 U9785 ( .A(n8198), .B(n8197), .Z(n8204) );
  AOI22_X1 U9786 ( .A1(n8265), .A2(n8746), .B1(P2_REG3_REG_17__SCAN_IN), .B2(
        P2_U3151), .ZN(n8200) );
  NAND2_X1 U9787 ( .A1(n8281), .A2(n8780), .ZN(n8199) );
  OAI211_X1 U9788 ( .C1(n8263), .C2(n8777), .A(n8200), .B(n8199), .ZN(n8201)
         );
  AOI21_X1 U9789 ( .B1(n8202), .B2(n8269), .A(n8201), .ZN(n8203) );
  OAI21_X1 U9790 ( .B1(n8204), .B2(n8271), .A(n8203), .ZN(P2_U3168) );
  XOR2_X1 U9791 ( .A(n8206), .B(n8205), .Z(n8211) );
  OAI22_X1 U9792 ( .A1(n8279), .A2(n8689), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10048), .ZN(n8208) );
  NOR2_X1 U9793 ( .A1(n8263), .A2(n8711), .ZN(n8207) );
  AOI211_X1 U9794 ( .C1(n8691), .C2(n8281), .A(n8208), .B(n8207), .ZN(n8210)
         );
  NAND2_X1 U9795 ( .A1(n6316), .A2(n8269), .ZN(n8209) );
  OAI211_X1 U9796 ( .C1(n8211), .C2(n8271), .A(n8210), .B(n8209), .ZN(P2_U3169) );
  OAI21_X1 U9797 ( .B1(n8214), .B2(n8213), .A(n8212), .ZN(n8215) );
  NAND2_X1 U9798 ( .A1(n8215), .A2(n8273), .ZN(n8219) );
  AOI22_X1 U9799 ( .A1(n8265), .A2(n8525), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8216) );
  OAI21_X1 U9800 ( .B1(n8736), .B2(n8263), .A(n8216), .ZN(n8217) );
  AOI21_X1 U9801 ( .B1(n8739), .B2(n8281), .A(n8217), .ZN(n8218) );
  OAI211_X1 U9802 ( .C1(n8920), .C2(n8285), .A(n8219), .B(n8218), .ZN(P2_U3173) );
  XOR2_X1 U9803 ( .A(n8221), .B(n8220), .Z(n8227) );
  AOI22_X1 U9804 ( .A1(n8277), .A2(n8525), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8223) );
  NAND2_X1 U9805 ( .A1(n8281), .A2(n8714), .ZN(n8222) );
  OAI211_X1 U9806 ( .C1(n8711), .C2(n8279), .A(n8223), .B(n8222), .ZN(n8224)
         );
  AOI21_X1 U9807 ( .B1(n8225), .B2(n8269), .A(n8224), .ZN(n8226) );
  OAI21_X1 U9808 ( .B1(n8227), .B2(n8271), .A(n8226), .ZN(P2_U3175) );
  OAI21_X1 U9809 ( .B1(n8230), .B2(n8228), .A(n8229), .ZN(n8231) );
  NAND2_X1 U9810 ( .A1(n8231), .A2(n8273), .ZN(n8237) );
  AOI22_X1 U9811 ( .A1(n8277), .A2(n6788), .B1(n4860), .B2(n8269), .ZN(n8236)
         );
  NAND2_X1 U9812 ( .A1(n8232), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n8235) );
  INV_X1 U9813 ( .A(n8539), .ZN(n8233) );
  OR2_X1 U9814 ( .A1(n8279), .A2(n8233), .ZN(n8234) );
  NAND4_X1 U9815 ( .A1(n8237), .A2(n8236), .A3(n8235), .A4(n8234), .ZN(
        P2_U3177) );
  XOR2_X1 U9816 ( .A(n8239), .B(n8238), .Z(n8245) );
  AOI22_X1 U9817 ( .A1(n8265), .A2(n8764), .B1(P2_REG3_REG_18__SCAN_IN), .B2(
        P2_U3151), .ZN(n8241) );
  NAND2_X1 U9818 ( .A1(n8281), .A2(n8769), .ZN(n8240) );
  OAI211_X1 U9819 ( .C1(n8263), .C2(n8789), .A(n8241), .B(n8240), .ZN(n8242)
         );
  AOI21_X1 U9820 ( .B1(n8243), .B2(n8269), .A(n8242), .ZN(n8244) );
  OAI21_X1 U9821 ( .B1(n8245), .B2(n8271), .A(n8244), .ZN(P2_U3178) );
  OAI211_X1 U9822 ( .C1(n8248), .C2(n8247), .A(n8246), .B(n8273), .ZN(n8256)
         );
  AOI22_X1 U9823 ( .A1(n8265), .A2(n8535), .B1(n8249), .B2(n8269), .ZN(n8255)
         );
  INV_X1 U9824 ( .A(n8250), .ZN(n8253) );
  NOR2_X1 U9825 ( .A1(n8267), .A2(n8251), .ZN(n8252) );
  AOI211_X1 U9826 ( .C1(n8277), .C2(n8537), .A(n8253), .B(n8252), .ZN(n8254)
         );
  NAND3_X1 U9827 ( .A1(n8256), .A2(n8255), .A3(n8254), .ZN(P2_U3179) );
  NAND2_X1 U9828 ( .A1(n8257), .A2(n8258), .ZN(n8262) );
  NAND2_X1 U9829 ( .A1(n8260), .A2(n8259), .ZN(n8261) );
  XNOR2_X1 U9830 ( .A(n8262), .B(n8261), .ZN(n8272) );
  OAI22_X1 U9831 ( .A1(n8263), .A2(n8689), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10108), .ZN(n8264) );
  AOI21_X1 U9832 ( .B1(n8265), .B2(n8664), .A(n8264), .ZN(n8266) );
  OAI21_X1 U9833 ( .B1(n8667), .B2(n8267), .A(n8266), .ZN(n8268) );
  AOI21_X1 U9834 ( .B1(n8670), .B2(n8269), .A(n8268), .ZN(n8270) );
  OAI21_X1 U9835 ( .B1(n8272), .B2(n8271), .A(n8270), .ZN(P2_U3180) );
  OAI211_X1 U9836 ( .C1(n8276), .C2(n8275), .A(n8274), .B(n8273), .ZN(n8284)
         );
  NAND2_X1 U9837 ( .A1(n8277), .A2(n8528), .ZN(n8278) );
  NAND2_X1 U9838 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8584) );
  OAI211_X1 U9839 ( .C1(n8777), .C2(n8279), .A(n8278), .B(n8584), .ZN(n8280)
         );
  AOI21_X1 U9840 ( .B1(n8282), .B2(n8281), .A(n8280), .ZN(n8283) );
  OAI211_X1 U9841 ( .C1(n8934), .C2(n8285), .A(n8284), .B(n8283), .ZN(P2_U3181) );
  NAND2_X1 U9842 ( .A1(n8945), .A2(n8288), .ZN(n8287) );
  OR2_X1 U9843 ( .A1(n8291), .A2(n6529), .ZN(n8286) );
  NAND2_X1 U9844 ( .A1(n8287), .A2(n8286), .ZN(n8875) );
  NAND2_X1 U9845 ( .A1(n8289), .A2(n8288), .ZN(n8293) );
  OR2_X1 U9846 ( .A1(n8291), .A2(n8290), .ZN(n8292) );
  NAND2_X1 U9847 ( .A1(n8293), .A2(n8292), .ZN(n8880) );
  NAND2_X1 U9848 ( .A1(n6090), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n8298) );
  INV_X1 U9849 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n8294) );
  OR2_X1 U9850 ( .A1(n4359), .A2(n8294), .ZN(n8297) );
  INV_X1 U9851 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n8295) );
  OR2_X1 U9852 ( .A1(n6411), .A2(n8295), .ZN(n8296) );
  NAND4_X1 U9853 ( .A1(n8299), .A2(n8298), .A3(n8297), .A4(n8296), .ZN(n8633)
         );
  INV_X1 U9854 ( .A(n8633), .ZN(n8300) );
  OR2_X1 U9855 ( .A1(n8875), .A2(n8300), .ZN(n8511) );
  INV_X1 U9856 ( .A(n8521), .ZN(n8301) );
  NAND2_X1 U9857 ( .A1(n8880), .A2(n8301), .ZN(n8453) );
  NAND2_X1 U9858 ( .A1(n8511), .A2(n8453), .ZN(n8498) );
  INV_X1 U9859 ( .A(n8502), .ZN(n8302) );
  INV_X1 U9860 ( .A(n8880), .ZN(n8808) );
  AND2_X1 U9861 ( .A1(n8808), .A2(n8521), .ZN(n8497) );
  INV_X1 U9862 ( .A(n8497), .ZN(n8504) );
  INV_X1 U9863 ( .A(n8304), .ZN(n8305) );
  OAI21_X1 U9864 ( .B1(n8805), .B2(n8504), .A(n8305), .ZN(n8458) );
  NAND2_X1 U9865 ( .A1(n8638), .A2(n8454), .ZN(n8306) );
  NAND2_X1 U9866 ( .A1(n8502), .A2(n8306), .ZN(n8309) );
  OR2_X1 U9867 ( .A1(n8307), .A2(n8446), .ZN(n8308) );
  NAND2_X1 U9868 ( .A1(n8309), .A2(n8308), .ZN(n8449) );
  NAND2_X1 U9869 ( .A1(n8312), .A2(n8310), .ZN(n8311) );
  NAND2_X1 U9870 ( .A1(n8311), .A2(n8446), .ZN(n8314) );
  NAND3_X1 U9871 ( .A1(n8320), .A2(n8312), .A3(n8516), .ZN(n8313) );
  NAND2_X1 U9872 ( .A1(n8314), .A2(n8313), .ZN(n8318) );
  NAND2_X1 U9873 ( .A1(n8316), .A2(n8315), .ZN(n8317) );
  NAND2_X1 U9874 ( .A1(n8318), .A2(n8317), .ZN(n8319) );
  MUX2_X1 U9875 ( .A(n8446), .B(n8319), .S(n6383), .Z(n8324) );
  NOR2_X1 U9876 ( .A1(n8320), .A2(n8454), .ZN(n8322) );
  NOR2_X1 U9877 ( .A1(n8322), .A2(n8321), .ZN(n8323) );
  NAND2_X1 U9878 ( .A1(n8324), .A2(n8323), .ZN(n8331) );
  NAND2_X1 U9879 ( .A1(n8338), .A2(n8325), .ZN(n8328) );
  NAND2_X1 U9880 ( .A1(n8332), .A2(n8326), .ZN(n8327) );
  MUX2_X1 U9881 ( .A(n8328), .B(n8327), .S(n8454), .Z(n8329) );
  INV_X1 U9882 ( .A(n8329), .ZN(n8330) );
  NAND2_X1 U9883 ( .A1(n8331), .A2(n8330), .ZN(n8340) );
  NAND3_X1 U9884 ( .A1(n8340), .A2(n8339), .A3(n8332), .ZN(n8334) );
  NAND3_X1 U9885 ( .A1(n8334), .A2(n8344), .A3(n8333), .ZN(n8335) );
  NAND3_X1 U9886 ( .A1(n8335), .A2(n8347), .A3(n8342), .ZN(n8337) );
  AND2_X1 U9887 ( .A1(n8353), .A2(n8446), .ZN(n8361) );
  AND2_X1 U9888 ( .A1(n8364), .A2(n8345), .ZN(n8336) );
  NAND4_X1 U9889 ( .A1(n8337), .A2(n8361), .A3(n8336), .A4(n8475), .ZN(n8370)
         );
  NAND3_X1 U9890 ( .A1(n8340), .A2(n8339), .A3(n8338), .ZN(n8343) );
  NAND3_X1 U9891 ( .A1(n8343), .A2(n8342), .A3(n8341), .ZN(n8346) );
  NAND3_X1 U9892 ( .A1(n8346), .A2(n8345), .A3(n8344), .ZN(n8349) );
  AND3_X1 U9893 ( .A1(n8363), .A2(n8454), .A3(n8347), .ZN(n8348) );
  NAND4_X1 U9894 ( .A1(n8349), .A2(n8348), .A3(n8356), .A4(n8475), .ZN(n8369)
         );
  OAI21_X1 U9895 ( .B1(n8350), .B2(n8535), .A(n8364), .ZN(n8351) );
  NAND3_X1 U9896 ( .A1(n8356), .A2(n8363), .A3(n8351), .ZN(n8352) );
  NAND3_X1 U9897 ( .A1(n8354), .A2(n8353), .A3(n8352), .ZN(n8355) );
  NAND2_X1 U9898 ( .A1(n8355), .A2(n8454), .ZN(n8360) );
  NAND2_X1 U9899 ( .A1(n8357), .A2(n8356), .ZN(n8358) );
  NAND2_X1 U9900 ( .A1(n8358), .A2(n8446), .ZN(n8359) );
  INV_X1 U9901 ( .A(n8361), .ZN(n8367) );
  NAND2_X1 U9902 ( .A1(n8363), .A2(n8362), .ZN(n8365) );
  NAND2_X1 U9903 ( .A1(n8365), .A2(n8364), .ZN(n8366) );
  OR2_X1 U9904 ( .A1(n8367), .A2(n8366), .ZN(n8368) );
  MUX2_X1 U9905 ( .A(n8454), .B(n8372), .S(n8371), .Z(n8381) );
  AND2_X1 U9906 ( .A1(n8373), .A2(n8454), .ZN(n8376) );
  NOR2_X1 U9907 ( .A1(n8465), .A2(n8532), .ZN(n8375) );
  MUX2_X1 U9908 ( .A(n8376), .B(n8375), .S(n8374), .Z(n8378) );
  AND2_X1 U9909 ( .A1(n8378), .A2(n8377), .ZN(n8380) );
  INV_X1 U9910 ( .A(n8379), .ZN(n8483) );
  OAI21_X1 U9911 ( .B1(n8381), .B2(n8380), .A(n8483), .ZN(n8385) );
  MUX2_X1 U9912 ( .A(n8383), .B(n8382), .S(n8454), .Z(n8384) );
  NAND2_X1 U9913 ( .A1(n8385), .A2(n8384), .ZN(n8391) );
  INV_X1 U9914 ( .A(n8386), .ZN(n8387) );
  NAND2_X1 U9915 ( .A1(n8391), .A2(n8387), .ZN(n8390) );
  MUX2_X1 U9916 ( .A(n8529), .B(n8388), .S(n8446), .Z(n8389) );
  INV_X1 U9917 ( .A(n8391), .ZN(n8393) );
  INV_X1 U9918 ( .A(n8394), .ZN(n8488) );
  MUX2_X1 U9919 ( .A(n8396), .B(n8395), .S(n8446), .Z(n8397) );
  NAND2_X1 U9920 ( .A1(n8488), .A2(n8397), .ZN(n8401) );
  MUX2_X1 U9921 ( .A(n8399), .B(n8398), .S(n8454), .Z(n8400) );
  MUX2_X1 U9922 ( .A(n8403), .B(n8402), .S(n8454), .Z(n8404) );
  NAND2_X1 U9923 ( .A1(n8405), .A2(n8404), .ZN(n8406) );
  INV_X1 U9924 ( .A(n8464), .ZN(n8408) );
  NAND3_X1 U9925 ( .A1(n8417), .A2(n8723), .A3(n8413), .ZN(n8410) );
  NAND3_X1 U9926 ( .A1(n8410), .A2(n8420), .A3(n8415), .ZN(n8412) );
  INV_X1 U9927 ( .A(n8413), .ZN(n8416) );
  OAI211_X1 U9928 ( .C1(n8417), .C2(n8416), .A(n8415), .B(n8414), .ZN(n8419)
         );
  NAND2_X1 U9929 ( .A1(n8419), .A2(n8418), .ZN(n8421) );
  MUX2_X1 U9930 ( .A(n8423), .B(n8422), .S(n8454), .Z(n8424) );
  NAND2_X1 U9931 ( .A1(n8430), .A2(n8692), .ZN(n8425) );
  NAND3_X1 U9932 ( .A1(n8425), .A2(n8460), .A3(n4899), .ZN(n8426) );
  NAND3_X1 U9933 ( .A1(n8426), .A2(n8446), .A3(n8459), .ZN(n8429) );
  INV_X1 U9934 ( .A(n8683), .ZN(n8675) );
  NOR2_X1 U9935 ( .A1(n8427), .A2(n8454), .ZN(n8428) );
  AOI21_X1 U9936 ( .B1(n8429), .B2(n8675), .A(n8428), .ZN(n8436) );
  NAND2_X1 U9937 ( .A1(n8430), .A2(n4899), .ZN(n8433) );
  NAND2_X1 U9938 ( .A1(n8460), .A2(n8454), .ZN(n8431) );
  AOI21_X1 U9939 ( .B1(n8433), .B2(n8432), .A(n8431), .ZN(n8435) );
  OAI22_X1 U9940 ( .A1(n8436), .A2(n8435), .B1(n8446), .B2(n8434), .ZN(n8438)
         );
  INV_X1 U9941 ( .A(n8662), .ZN(n8437) );
  INV_X1 U9942 ( .A(n8656), .ZN(n8442) );
  MUX2_X1 U9943 ( .A(n8440), .B(n8439), .S(n8454), .Z(n8441) );
  MUX2_X1 U9944 ( .A(n8444), .B(n8443), .S(n8446), .Z(n8445) );
  MUX2_X1 U9945 ( .A(n8522), .B(n8647), .S(n8446), .Z(n8448) );
  INV_X1 U9946 ( .A(n8448), .ZN(n8447) );
  NOR2_X1 U9947 ( .A1(n8451), .A2(n8447), .ZN(n8505) );
  NAND2_X1 U9948 ( .A1(n8449), .A2(n8448), .ZN(n8450) );
  OAI211_X1 U9949 ( .C1(n8499), .C2(n8522), .A(n8452), .B(n8453), .ZN(n8456)
         );
  AOI211_X1 U9950 ( .C1(n8454), .C2(n8453), .A(n8512), .B(n8497), .ZN(n8455)
         );
  OAI21_X1 U9951 ( .B1(n8505), .B2(n8456), .A(n8455), .ZN(n8457) );
  NAND2_X1 U9952 ( .A1(n8460), .A2(n8459), .ZN(n8695) );
  INV_X1 U9953 ( .A(n8692), .ZN(n8461) );
  NOR2_X1 U9954 ( .A1(n8462), .A2(n8461), .ZN(n8701) );
  NOR2_X1 U9955 ( .A1(n8464), .A2(n4593), .ZN(n8767) );
  INV_X1 U9956 ( .A(n8465), .ZN(n8482) );
  NOR2_X1 U9957 ( .A1(n4669), .A2(n8466), .ZN(n8468) );
  NAND4_X1 U9958 ( .A1(n8470), .A2(n8469), .A3(n8468), .A4(n8467), .ZN(n8474)
         );
  NOR4_X1 U9959 ( .A1(n8474), .A2(n8473), .A3(n8472), .A4(n8471), .ZN(n8478)
         );
  NAND4_X1 U9960 ( .A1(n8476), .A2(n8477), .A3(n8478), .A4(n8475), .ZN(n8480)
         );
  NOR2_X1 U9961 ( .A1(n8480), .A2(n8479), .ZN(n8481) );
  NAND3_X1 U9962 ( .A1(n8483), .A2(n8482), .A3(n8481), .ZN(n8484) );
  NOR3_X1 U9963 ( .A1(n8486), .A2(n8485), .A3(n8484), .ZN(n8487) );
  AND3_X1 U9964 ( .A1(n8795), .A2(n8488), .A3(n8487), .ZN(n8489) );
  NAND4_X1 U9965 ( .A1(n8749), .A2(n8779), .A3(n8767), .A4(n8489), .ZN(n8490)
         );
  NOR2_X1 U9966 ( .A1(n8738), .A2(n8490), .ZN(n8491) );
  NAND4_X1 U9967 ( .A1(n8701), .A2(n8708), .A3(n8725), .A4(n8491), .ZN(n8492)
         );
  OR3_X1 U9968 ( .A1(n8683), .A2(n8695), .A3(n8492), .ZN(n8494) );
  OR4_X1 U9969 ( .A1(n8494), .A2(n8493), .A3(n8656), .A4(n8662), .ZN(n8495) );
  OR4_X1 U9970 ( .A1(n8498), .A2(n8497), .A3(n8496), .A4(n8495), .ZN(n8510) );
  INV_X1 U9971 ( .A(n8647), .ZN(n8887) );
  NAND2_X1 U9972 ( .A1(n8500), .A2(n8887), .ZN(n8508) );
  INV_X1 U9973 ( .A(n8501), .ZN(n8503) );
  AND4_X1 U9974 ( .A1(n8504), .A2(n8503), .A3(n8516), .A4(n8502), .ZN(n8507)
         );
  INV_X1 U9975 ( .A(n8505), .ZN(n8506) );
  NAND3_X1 U9976 ( .A1(n8508), .A2(n8507), .A3(n8506), .ZN(n8509) );
  OAI211_X1 U9977 ( .C1(n8512), .C2(n8511), .A(n8510), .B(n8509), .ZN(n8513)
         );
  NOR3_X1 U9978 ( .A1(n8515), .A2(n8514), .A3(n5960), .ZN(n8518) );
  OAI21_X1 U9979 ( .B1(n8519), .B2(n8516), .A(P2_B_REG_SCAN_IN), .ZN(n8517) );
  OAI22_X1 U9980 ( .A1(n8520), .A2(n8519), .B1(n8518), .B2(n8517), .ZN(
        P2_U3296) );
  MUX2_X1 U9981 ( .A(n8633), .B(P2_DATAO_REG_31__SCAN_IN), .S(n8621), .Z(
        P2_U3522) );
  MUX2_X1 U9982 ( .A(n8521), .B(P2_DATAO_REG_30__SCAN_IN), .S(n8621), .Z(
        P2_U3521) );
  MUX2_X1 U9983 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n8522), .S(P2_U3893), .Z(
        P2_U3519) );
  MUX2_X1 U9984 ( .A(n8664), .B(P2_DATAO_REG_27__SCAN_IN), .S(n8621), .Z(
        P2_U3518) );
  MUX2_X1 U9985 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n6337), .S(P2_U3893), .Z(
        P2_U3517) );
  MUX2_X1 U9986 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n6315), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U9987 ( .A(n8523), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8621), .Z(
        P2_U3514) );
  MUX2_X1 U9988 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8524), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U9989 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8525), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U9990 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n6274), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U9991 ( .A(n8764), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8621), .Z(
        P2_U3510) );
  MUX2_X1 U9992 ( .A(n8746), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8621), .Z(
        P2_U3509) );
  MUX2_X1 U9993 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8526), .S(P2_U3893), .Z(
        P2_U3507) );
  MUX2_X1 U9994 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8527), .S(P2_U3893), .Z(
        P2_U3506) );
  MUX2_X1 U9995 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8528), .S(P2_U3893), .Z(
        P2_U3505) );
  MUX2_X1 U9996 ( .A(n8529), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8621), .Z(
        P2_U3504) );
  MUX2_X1 U9997 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n8530), .S(P2_U3893), .Z(
        P2_U3503) );
  MUX2_X1 U9998 ( .A(n8531), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8621), .Z(
        P2_U3502) );
  MUX2_X1 U9999 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n8532), .S(P2_U3893), .Z(
        P2_U3501) );
  MUX2_X1 U10000 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n8533), .S(P2_U3893), .Z(
        P2_U3500) );
  MUX2_X1 U10001 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n8534), .S(P2_U3893), .Z(
        P2_U3499) );
  MUX2_X1 U10002 ( .A(n8535), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8621), .Z(
        P2_U3498) );
  MUX2_X1 U10003 ( .A(n8536), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8621), .Z(
        P2_U3497) );
  MUX2_X1 U10004 ( .A(n8537), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8621), .Z(
        P2_U3496) );
  MUX2_X1 U10005 ( .A(n8538), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8621), .Z(
        P2_U3495) );
  MUX2_X1 U10006 ( .A(n8539), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8621), .Z(
        P2_U3494) );
  MUX2_X1 U10007 ( .A(n6102), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8621), .Z(
        P2_U3493) );
  MUX2_X1 U10008 ( .A(n6788), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8621), .Z(
        P2_U3492) );
  MUX2_X1 U10009 ( .A(n6382), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8621), .Z(
        P2_U3491) );
  AOI21_X1 U10010 ( .B1(n8872), .B2(n8541), .A(n8540), .ZN(n8556) );
  AOI21_X1 U10011 ( .B1(n8544), .B2(n8543), .A(n8542), .ZN(n8545) );
  NOR2_X1 U10012 ( .A1(n8545), .A2(n9810), .ZN(n8554) );
  AOI21_X1 U10013 ( .B1(n8548), .B2(n8547), .A(n8546), .ZN(n8552) );
  AOI22_X1 U10014 ( .A1(n9772), .A2(n8549), .B1(n9796), .B2(
        P2_ADDR_REG_13__SCAN_IN), .ZN(n8551) );
  OAI211_X1 U10015 ( .C1(n8552), .C2(n8624), .A(n8551), .B(n8550), .ZN(n8553)
         );
  NOR2_X1 U10016 ( .A1(n8554), .A2(n8553), .ZN(n8555) );
  OAI21_X1 U10017 ( .B1(n8556), .B2(n9803), .A(n8555), .ZN(P2_U3195) );
  AOI21_X1 U10018 ( .B1(n4446), .B2(n8558), .A(n8557), .ZN(n8573) );
  AOI21_X1 U10019 ( .B1(n8561), .B2(n8560), .A(n8559), .ZN(n8562) );
  NOR2_X1 U10020 ( .A1(n8562), .A2(n9810), .ZN(n8571) );
  AOI21_X1 U10021 ( .B1(n8565), .B2(n8564), .A(n8563), .ZN(n8569) );
  AOI22_X1 U10022 ( .A1(n9772), .A2(n8566), .B1(n9796), .B2(
        P2_ADDR_REG_14__SCAN_IN), .ZN(n8568) );
  OAI211_X1 U10023 ( .C1(n8569), .C2(n8624), .A(n8568), .B(n8567), .ZN(n8570)
         );
  NOR2_X1 U10024 ( .A1(n8571), .A2(n8570), .ZN(n8572) );
  OAI21_X1 U10025 ( .B1(n8573), .B2(n9803), .A(n8572), .ZN(P2_U3196) );
  AOI21_X1 U10026 ( .B1(n8864), .B2(n8575), .A(n8574), .ZN(n8590) );
  AOI21_X1 U10027 ( .B1(n8578), .B2(n8577), .A(n8576), .ZN(n8579) );
  NOR2_X1 U10028 ( .A1(n8579), .A2(n9810), .ZN(n8588) );
  AOI21_X1 U10029 ( .B1(n8582), .B2(n8581), .A(n8580), .ZN(n8586) );
  AOI22_X1 U10030 ( .A1(n9772), .A2(n8583), .B1(n9796), .B2(
        P2_ADDR_REG_15__SCAN_IN), .ZN(n8585) );
  OAI211_X1 U10031 ( .C1(n8586), .C2(n8624), .A(n8585), .B(n8584), .ZN(n8587)
         );
  NOR2_X1 U10032 ( .A1(n8588), .A2(n8587), .ZN(n8589) );
  OAI21_X1 U10033 ( .B1(n8590), .B2(n9803), .A(n8589), .ZN(P2_U3197) );
  AOI21_X1 U10034 ( .B1(n8593), .B2(n8592), .A(n8591), .ZN(n8609) );
  INV_X1 U10035 ( .A(n8594), .ZN(n8595) );
  NAND2_X1 U10036 ( .A1(n8596), .A2(n8595), .ZN(n8597) );
  XNOR2_X1 U10037 ( .A(n8598), .B(n8597), .ZN(n8607) );
  INV_X1 U10038 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n9893) );
  NAND2_X1 U10039 ( .A1(n9772), .A2(n8599), .ZN(n8600) );
  OAI211_X1 U10040 ( .C1(n8628), .C2(n9893), .A(n8601), .B(n8600), .ZN(n8606)
         );
  AOI21_X1 U10041 ( .B1(n4410), .B2(n8603), .A(n8602), .ZN(n8604) );
  NOR2_X1 U10042 ( .A1(n8604), .A2(n9810), .ZN(n8605) );
  AOI211_X1 U10043 ( .C1(n9807), .C2(n8607), .A(n8606), .B(n8605), .ZN(n8608)
         );
  OAI21_X1 U10044 ( .B1(n8609), .B2(n9803), .A(n8608), .ZN(P2_U3198) );
  AOI21_X1 U10045 ( .B1(n8612), .B2(n8611), .A(n8610), .ZN(n8631) );
  INV_X1 U10046 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n9911) );
  INV_X1 U10047 ( .A(n8618), .ZN(n8619) );
  NOR2_X1 U10048 ( .A1(n8620), .A2(n8619), .ZN(n8625) );
  INV_X1 U10049 ( .A(n8625), .ZN(n8622) );
  INV_X1 U10050 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n8623) );
  NOR2_X1 U10051 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8623), .ZN(n8626) );
  OAI21_X1 U10052 ( .B1(n8631), .B2(n9803), .A(n8630), .ZN(P2_U3200) );
  NAND2_X1 U10053 ( .A1(n8633), .A2(n8632), .ZN(n8876) );
  AOI21_X1 U10054 ( .B1(n8634), .B2(n8876), .A(n8803), .ZN(n8636) );
  AOI21_X1 U10055 ( .B1(n8803), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8636), .ZN(
        n8635) );
  OAI21_X1 U10056 ( .B1(n8805), .B2(n8798), .A(n8635), .ZN(P2_U3202) );
  AOI21_X1 U10057 ( .B1(n8803), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8636), .ZN(
        n8637) );
  OAI21_X1 U10058 ( .B1(n8808), .B2(n8798), .A(n8637), .ZN(P2_U3203) );
  OAI22_X1 U10059 ( .A1(n8639), .A2(n8790), .B1(n8638), .B2(n8788), .ZN(n8640)
         );
  OAI22_X1 U10060 ( .A1(n9824), .A2(n8642), .B1(n8641), .B2(n8679), .ZN(n8646)
         );
  XNOR2_X1 U10061 ( .A(n8644), .B(n8643), .ZN(n8810) );
  NOR2_X1 U10062 ( .A1(n8810), .A2(n8673), .ZN(n8645) );
  AOI211_X1 U10063 ( .C1(n9819), .C2(n8647), .A(n8646), .B(n8645), .ZN(n8648)
         );
  OAI21_X1 U10064 ( .B1(n8809), .B2(n8803), .A(n8648), .ZN(P2_U3205) );
  XOR2_X1 U10065 ( .A(n8649), .B(n8656), .Z(n8652) );
  OAI22_X1 U10066 ( .A1(n8650), .A2(n8788), .B1(n8678), .B2(n8790), .ZN(n8651)
         );
  OAI22_X1 U10067 ( .A1(n9824), .A2(n8654), .B1(n8653), .B2(n8679), .ZN(n8658)
         );
  XNOR2_X1 U10068 ( .A(n8655), .B(n8656), .ZN(n8814) );
  NOR2_X1 U10069 ( .A1(n8814), .A2(n8673), .ZN(n8657) );
  AOI211_X1 U10070 ( .C1(n9819), .C2(n8890), .A(n8658), .B(n8657), .ZN(n8659)
         );
  OAI21_X1 U10071 ( .B1(n8813), .B2(n8803), .A(n8659), .ZN(P2_U3206) );
  XNOR2_X1 U10072 ( .A(n8660), .B(n8662), .ZN(n8819) );
  INV_X1 U10073 ( .A(n8819), .ZN(n8674) );
  OAI211_X1 U10074 ( .C1(n8663), .C2(n8662), .A(n8661), .B(n8759), .ZN(n8666)
         );
  NAND2_X1 U10075 ( .A1(n8664), .A2(n8763), .ZN(n8665) );
  OAI211_X1 U10076 ( .C1(n8689), .C2(n8790), .A(n8666), .B(n8665), .ZN(n8818)
         );
  NAND2_X1 U10077 ( .A1(n8818), .A2(n9824), .ZN(n8672) );
  OAI22_X1 U10078 ( .A1(n9824), .A2(n8668), .B1(n8667), .B2(n8679), .ZN(n8669)
         );
  AOI21_X1 U10079 ( .B1(n8670), .B2(n9819), .A(n8669), .ZN(n8671) );
  OAI211_X1 U10080 ( .C1(n8674), .C2(n8673), .A(n8672), .B(n8671), .ZN(
        P2_U3207) );
  XNOR2_X1 U10081 ( .A(n8676), .B(n8675), .ZN(n8677) );
  OAI222_X1 U10082 ( .A1(n8788), .A2(n8678), .B1(n8790), .B2(n8700), .C1(n8786), .C2(n8677), .ZN(n8822) );
  OAI22_X1 U10083 ( .A1(n8900), .A2(n8686), .B1(n8680), .B2(n8679), .ZN(n8681)
         );
  OAI21_X1 U10084 ( .B1(n8822), .B2(n8681), .A(n9824), .ZN(n8685) );
  XNOR2_X1 U10085 ( .A(n8682), .B(n8683), .ZN(n8823) );
  AOI22_X1 U10086 ( .A1(n8823), .A2(n8801), .B1(P2_REG2_REG_25__SCAN_IN), .B2(
        n8803), .ZN(n8684) );
  NAND2_X1 U10087 ( .A1(n8685), .A2(n8684), .ZN(P2_U3208) );
  NOR2_X1 U10088 ( .A1(n8904), .A2(n8686), .ZN(n8690) );
  XOR2_X1 U10089 ( .A(n8695), .B(n8687), .Z(n8688) );
  OAI222_X1 U10090 ( .A1(n8790), .A2(n8711), .B1(n8788), .B2(n8689), .C1(n8688), .C2(n8786), .ZN(n8826) );
  AOI211_X1 U10091 ( .C1(n9821), .C2(n8691), .A(n8690), .B(n8826), .ZN(n8697)
         );
  NAND2_X1 U10092 ( .A1(n8693), .A2(n8692), .ZN(n8694) );
  XOR2_X1 U10093 ( .A(n8695), .B(n8694), .Z(n8827) );
  AOI22_X1 U10094 ( .A1(n8827), .A2(n8801), .B1(P2_REG2_REG_24__SCAN_IN), .B2(
        n8803), .ZN(n8696) );
  OAI21_X1 U10095 ( .B1(n8697), .B2(n8803), .A(n8696), .ZN(P2_U3209) );
  XOR2_X1 U10096 ( .A(n8701), .B(n8698), .Z(n8699) );
  OAI222_X1 U10097 ( .A1(n8790), .A2(n8721), .B1(n8788), .B2(n8700), .C1(n8786), .C2(n8699), .ZN(n8830) );
  INV_X1 U10098 ( .A(n8830), .ZN(n8707) );
  XOR2_X1 U10099 ( .A(n8702), .B(n8701), .Z(n8831) );
  AOI22_X1 U10100 ( .A1(n8703), .A2(n9821), .B1(n8803), .B2(
        P2_REG2_REG_23__SCAN_IN), .ZN(n8704) );
  OAI21_X1 U10101 ( .B1(n8908), .B2(n8798), .A(n8704), .ZN(n8705) );
  AOI21_X1 U10102 ( .B1(n8831), .B2(n8801), .A(n8705), .ZN(n8706) );
  OAI21_X1 U10103 ( .B1(n8707), .B2(n8803), .A(n8706), .ZN(P2_U3210) );
  XNOR2_X1 U10104 ( .A(n4686), .B(n8708), .ZN(n8710) );
  OAI222_X1 U10105 ( .A1(n8788), .A2(n8711), .B1(n8790), .B2(n8735), .C1(n8786), .C2(n8710), .ZN(n8834) );
  INV_X1 U10106 ( .A(n8834), .ZN(n8718) );
  XNOR2_X1 U10107 ( .A(n8712), .B(n8713), .ZN(n8835) );
  AOI22_X1 U10108 ( .A1(n8803), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n9821), .B2(
        n8714), .ZN(n8715) );
  OAI21_X1 U10109 ( .B1(n8912), .B2(n8798), .A(n8715), .ZN(n8716) );
  AOI21_X1 U10110 ( .B1(n8835), .B2(n8801), .A(n8716), .ZN(n8717) );
  OAI21_X1 U10111 ( .B1(n8718), .B2(n8803), .A(n8717), .ZN(P2_U3211) );
  XOR2_X1 U10112 ( .A(n8725), .B(n8719), .Z(n8720) );
  OAI222_X1 U10113 ( .A1(n8790), .A2(n8722), .B1(n8788), .B2(n8721), .C1(n8786), .C2(n8720), .ZN(n8838) );
  INV_X1 U10114 ( .A(n8838), .ZN(n8732) );
  NAND2_X1 U10115 ( .A1(n8724), .A2(n8723), .ZN(n8726) );
  XNOR2_X1 U10116 ( .A(n8726), .B(n8725), .ZN(n8839) );
  INV_X1 U10117 ( .A(n8727), .ZN(n8916) );
  AOI22_X1 U10118 ( .A1(n8803), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n9821), .B2(
        n8728), .ZN(n8729) );
  OAI21_X1 U10119 ( .B1(n8916), .B2(n8798), .A(n8729), .ZN(n8730) );
  AOI21_X1 U10120 ( .B1(n8839), .B2(n8801), .A(n8730), .ZN(n8731) );
  OAI21_X1 U10121 ( .B1(n8732), .B2(n8803), .A(n8731), .ZN(P2_U3212) );
  XOR2_X1 U10122 ( .A(n8733), .B(n8738), .Z(n8734) );
  OAI222_X1 U10123 ( .A1(n8790), .A2(n8736), .B1(n8788), .B2(n8735), .C1(n8786), .C2(n8734), .ZN(n8842) );
  INV_X1 U10124 ( .A(n8842), .ZN(n8743) );
  XOR2_X1 U10125 ( .A(n8737), .B(n8738), .Z(n8843) );
  AOI22_X1 U10126 ( .A1(n8803), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n9821), .B2(
        n8739), .ZN(n8740) );
  OAI21_X1 U10127 ( .B1(n8920), .B2(n8798), .A(n8740), .ZN(n8741) );
  AOI21_X1 U10128 ( .B1(n8843), .B2(n8801), .A(n8741), .ZN(n8742) );
  OAI21_X1 U10129 ( .B1(n8743), .B2(n8803), .A(n8742), .ZN(P2_U3213) );
  XNOR2_X1 U10130 ( .A(n8744), .B(n8749), .ZN(n8747) );
  AOI222_X1 U10131 ( .A1(n8759), .A2(n8747), .B1(n6274), .B2(n8763), .C1(n8746), .C2(n8745), .ZN(n8849) );
  OAI21_X1 U10132 ( .B1(n8750), .B2(n8749), .A(n8748), .ZN(n8847) );
  AOI22_X1 U10133 ( .A1(n8803), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n9821), .B2(
        n8751), .ZN(n8752) );
  OAI21_X1 U10134 ( .B1(n8753), .B2(n8798), .A(n8752), .ZN(n8754) );
  AOI21_X1 U10135 ( .B1(n8847), .B2(n8801), .A(n8754), .ZN(n8755) );
  OAI21_X1 U10136 ( .B1(n8849), .B2(n8803), .A(n8755), .ZN(P2_U3214) );
  INV_X1 U10137 ( .A(n8767), .ZN(n8762) );
  INV_X1 U10138 ( .A(n8756), .ZN(n8758) );
  NAND2_X1 U10139 ( .A1(n8758), .A2(n8757), .ZN(n8760) );
  OAI211_X1 U10140 ( .C1(n8762), .C2(n8761), .A(n8760), .B(n8759), .ZN(n8766)
         );
  NAND2_X1 U10141 ( .A1(n8764), .A2(n8763), .ZN(n8765) );
  OAI211_X1 U10142 ( .C1(n8789), .C2(n8790), .A(n8766), .B(n8765), .ZN(n8850)
         );
  INV_X1 U10143 ( .A(n8850), .ZN(n8773) );
  XOR2_X1 U10144 ( .A(n8768), .B(n8767), .Z(n8851) );
  AOI22_X1 U10145 ( .A1(n8803), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n9821), .B2(
        n8769), .ZN(n8770) );
  OAI21_X1 U10146 ( .B1(n8925), .B2(n8798), .A(n8770), .ZN(n8771) );
  AOI21_X1 U10147 ( .B1(n8851), .B2(n8801), .A(n8771), .ZN(n8772) );
  OAI21_X1 U10148 ( .B1(n8773), .B2(n8803), .A(n8772), .ZN(P2_U3215) );
  XNOR2_X1 U10149 ( .A(n8774), .B(n8779), .ZN(n8775) );
  OAI222_X1 U10150 ( .A1(n8790), .A2(n8777), .B1(n8788), .B2(n8776), .C1(n8775), .C2(n8786), .ZN(n8854) );
  INV_X1 U10151 ( .A(n8854), .ZN(n8784) );
  XOR2_X1 U10152 ( .A(n8778), .B(n8779), .Z(n8855) );
  AOI22_X1 U10153 ( .A1(n8803), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n9821), .B2(
        n8780), .ZN(n8781) );
  OAI21_X1 U10154 ( .B1(n8929), .B2(n8798), .A(n8781), .ZN(n8782) );
  AOI21_X1 U10155 ( .B1(n8855), .B2(n8801), .A(n8782), .ZN(n8783) );
  OAI21_X1 U10156 ( .B1(n8784), .B2(n8803), .A(n8783), .ZN(P2_U3216) );
  AOI211_X1 U10157 ( .C1(n8795), .C2(n8787), .A(n8786), .B(n8785), .ZN(n8793)
         );
  OAI22_X1 U10158 ( .A1(n8791), .A2(n8790), .B1(n8789), .B2(n8788), .ZN(n8792)
         );
  NOR2_X1 U10159 ( .A1(n8793), .A2(n8792), .ZN(n8860) );
  XOR2_X1 U10160 ( .A(n8794), .B(n8795), .Z(n8858) );
  INV_X1 U10161 ( .A(n8857), .ZN(n8799) );
  AOI22_X1 U10162 ( .A1(n8803), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n9821), .B2(
        n8796), .ZN(n8797) );
  OAI21_X1 U10163 ( .B1(n8799), .B2(n8798), .A(n8797), .ZN(n8800) );
  AOI21_X1 U10164 ( .B1(n8858), .B2(n8801), .A(n8800), .ZN(n8802) );
  OAI21_X1 U10165 ( .B1(n8860), .B2(n8803), .A(n8802), .ZN(P2_U3217) );
  NOR2_X1 U10166 ( .A1(n9885), .A2(n8876), .ZN(n8806) );
  AOI21_X1 U10167 ( .B1(P2_REG1_REG_31__SCAN_IN), .B2(n9885), .A(n8806), .ZN(
        n8804) );
  OAI21_X1 U10168 ( .B1(n8805), .B2(n8874), .A(n8804), .ZN(P2_U3490) );
  AOI21_X1 U10169 ( .B1(P2_REG1_REG_30__SCAN_IN), .B2(n9885), .A(n8806), .ZN(
        n8807) );
  OAI21_X1 U10170 ( .B1(n8808), .B2(n8874), .A(n8807), .ZN(P2_U3489) );
  OAI21_X1 U10171 ( .B1(n9866), .B2(n8810), .A(n8809), .ZN(n8884) );
  MUX2_X1 U10172 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n8884), .S(n9887), .Z(n8811) );
  INV_X1 U10173 ( .A(n8811), .ZN(n8812) );
  OAI21_X1 U10174 ( .B1(n8887), .B2(n8874), .A(n8812), .ZN(P2_U3487) );
  OAI21_X1 U10175 ( .B1(n9866), .B2(n8814), .A(n8813), .ZN(n8888) );
  MUX2_X1 U10176 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8888), .S(n9887), .Z(n8815) );
  AOI21_X1 U10177 ( .B1(n8816), .B2(n8890), .A(n8815), .ZN(n8817) );
  INV_X1 U10178 ( .A(n8817), .ZN(P2_U3486) );
  AOI21_X1 U10179 ( .B1(n9853), .B2(n8819), .A(n8818), .ZN(n8893) );
  MUX2_X1 U10180 ( .A(n8820), .B(n8893), .S(n9887), .Z(n8821) );
  OAI21_X1 U10181 ( .B1(n8896), .B2(n8874), .A(n8821), .ZN(P2_U3485) );
  INV_X1 U10182 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n8824) );
  AOI21_X1 U10183 ( .B1(n9853), .B2(n8823), .A(n8822), .ZN(n8897) );
  MUX2_X1 U10184 ( .A(n8824), .B(n8897), .S(n9887), .Z(n8825) );
  OAI21_X1 U10185 ( .B1(n8900), .B2(n8874), .A(n8825), .ZN(P2_U3484) );
  INV_X1 U10186 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n8828) );
  AOI21_X1 U10187 ( .B1(n8827), .B2(n9853), .A(n8826), .ZN(n8901) );
  MUX2_X1 U10188 ( .A(n8828), .B(n8901), .S(n9887), .Z(n8829) );
  OAI21_X1 U10189 ( .B1(n8904), .B2(n8874), .A(n8829), .ZN(P2_U3483) );
  INV_X1 U10190 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8832) );
  AOI21_X1 U10191 ( .B1(n9853), .B2(n8831), .A(n8830), .ZN(n8905) );
  MUX2_X1 U10192 ( .A(n8832), .B(n8905), .S(n9887), .Z(n8833) );
  OAI21_X1 U10193 ( .B1(n8908), .B2(n8874), .A(n8833), .ZN(P2_U3482) );
  INV_X1 U10194 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8836) );
  AOI21_X1 U10195 ( .B1(n9853), .B2(n8835), .A(n8834), .ZN(n8909) );
  MUX2_X1 U10196 ( .A(n8836), .B(n8909), .S(n9887), .Z(n8837) );
  OAI21_X1 U10197 ( .B1(n8912), .B2(n8874), .A(n8837), .ZN(P2_U3481) );
  INV_X1 U10198 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8840) );
  AOI21_X1 U10199 ( .B1(n8839), .B2(n9853), .A(n8838), .ZN(n8913) );
  MUX2_X1 U10200 ( .A(n8840), .B(n8913), .S(n9887), .Z(n8841) );
  OAI21_X1 U10201 ( .B1(n8916), .B2(n8874), .A(n8841), .ZN(P2_U3480) );
  INV_X1 U10202 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8844) );
  AOI21_X1 U10203 ( .B1(n8843), .B2(n9853), .A(n8842), .ZN(n8917) );
  MUX2_X1 U10204 ( .A(n8844), .B(n8917), .S(n9887), .Z(n8845) );
  OAI21_X1 U10205 ( .B1(n8920), .B2(n8874), .A(n8845), .ZN(P2_U3479) );
  AOI22_X1 U10206 ( .A1(n8847), .A2(n9853), .B1(n9871), .B2(n8846), .ZN(n8848)
         );
  NAND2_X1 U10207 ( .A1(n8849), .A2(n8848), .ZN(n8921) );
  MUX2_X1 U10208 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8921), .S(n9887), .Z(
        P2_U3478) );
  INV_X1 U10209 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8852) );
  AOI21_X1 U10210 ( .B1(n9853), .B2(n8851), .A(n8850), .ZN(n8922) );
  MUX2_X1 U10211 ( .A(n8852), .B(n8922), .S(n9887), .Z(n8853) );
  OAI21_X1 U10212 ( .B1(n8925), .B2(n8874), .A(n8853), .ZN(P2_U3477) );
  AOI21_X1 U10213 ( .B1(n9853), .B2(n8855), .A(n8854), .ZN(n8926) );
  MUX2_X1 U10214 ( .A(n9802), .B(n8926), .S(n9887), .Z(n8856) );
  OAI21_X1 U10215 ( .B1(n8929), .B2(n8874), .A(n8856), .ZN(P2_U3476) );
  AOI22_X1 U10216 ( .A1(n8858), .A2(n9853), .B1(n9871), .B2(n8857), .ZN(n8859)
         );
  NAND2_X1 U10217 ( .A1(n8860), .A2(n8859), .ZN(n8930) );
  MUX2_X1 U10218 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8930), .S(n9887), .Z(
        P2_U3475) );
  INV_X1 U10219 ( .A(n8861), .ZN(n8862) );
  AOI21_X1 U10220 ( .B1(n8863), .B2(n9853), .A(n8862), .ZN(n8931) );
  MUX2_X1 U10221 ( .A(n8864), .B(n8931), .S(n9887), .Z(n8865) );
  OAI21_X1 U10222 ( .B1(n8934), .B2(n8874), .A(n8865), .ZN(P2_U3474) );
  AOI21_X1 U10223 ( .B1(n8867), .B2(n9853), .A(n8866), .ZN(n8935) );
  MUX2_X1 U10224 ( .A(n8868), .B(n8935), .S(n9887), .Z(n8869) );
  OAI21_X1 U10225 ( .B1(n8938), .B2(n8874), .A(n8869), .ZN(P2_U3473) );
  AOI21_X1 U10226 ( .B1(n8871), .B2(n9853), .A(n8870), .ZN(n8940) );
  MUX2_X1 U10227 ( .A(n8872), .B(n8940), .S(n9887), .Z(n8873) );
  OAI21_X1 U10228 ( .B1(n8944), .B2(n8874), .A(n8873), .ZN(P2_U3472) );
  INV_X1 U10229 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n8879) );
  NAND2_X1 U10230 ( .A1(n8875), .A2(n8891), .ZN(n8878) );
  INV_X1 U10231 ( .A(n8876), .ZN(n8877) );
  NAND2_X1 U10232 ( .A1(n8939), .A2(n8877), .ZN(n8881) );
  OAI211_X1 U10233 ( .C1(n8879), .C2(n8939), .A(n8878), .B(n8881), .ZN(
        P2_U3458) );
  INV_X1 U10234 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n8883) );
  NAND2_X1 U10235 ( .A1(n8880), .A2(n8891), .ZN(n8882) );
  OAI211_X1 U10236 ( .C1(n8883), .C2(n8939), .A(n8882), .B(n8881), .ZN(
        P2_U3457) );
  MUX2_X1 U10237 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n8884), .S(n8939), .Z(n8885) );
  INV_X1 U10238 ( .A(n8885), .ZN(n8886) );
  OAI21_X1 U10239 ( .B1(n8887), .B2(n8943), .A(n8886), .ZN(P2_U3455) );
  MUX2_X1 U10240 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8888), .S(n8939), .Z(n8889) );
  AOI21_X1 U10241 ( .B1(n8891), .B2(n8890), .A(n8889), .ZN(n8892) );
  INV_X1 U10242 ( .A(n8892), .ZN(P2_U3454) );
  INV_X1 U10243 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8894) );
  MUX2_X1 U10244 ( .A(n8894), .B(n8893), .S(n8939), .Z(n8895) );
  OAI21_X1 U10245 ( .B1(n8896), .B2(n8943), .A(n8895), .ZN(P2_U3453) );
  MUX2_X1 U10246 ( .A(n8898), .B(n8897), .S(n8939), .Z(n8899) );
  OAI21_X1 U10247 ( .B1(n8900), .B2(n8943), .A(n8899), .ZN(P2_U3452) );
  MUX2_X1 U10248 ( .A(n8902), .B(n8901), .S(n8939), .Z(n8903) );
  OAI21_X1 U10249 ( .B1(n8904), .B2(n8943), .A(n8903), .ZN(P2_U3451) );
  MUX2_X1 U10250 ( .A(n8906), .B(n8905), .S(n8939), .Z(n8907) );
  OAI21_X1 U10251 ( .B1(n8908), .B2(n8943), .A(n8907), .ZN(P2_U3450) );
  MUX2_X1 U10252 ( .A(n8910), .B(n8909), .S(n8939), .Z(n8911) );
  OAI21_X1 U10253 ( .B1(n8912), .B2(n8943), .A(n8911), .ZN(P2_U3449) );
  MUX2_X1 U10254 ( .A(n8914), .B(n8913), .S(n8939), .Z(n8915) );
  OAI21_X1 U10255 ( .B1(n8916), .B2(n8943), .A(n8915), .ZN(P2_U3448) );
  INV_X1 U10256 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n8918) );
  MUX2_X1 U10257 ( .A(n8918), .B(n8917), .S(n8939), .Z(n8919) );
  OAI21_X1 U10258 ( .B1(n8920), .B2(n8943), .A(n8919), .ZN(P2_U3447) );
  MUX2_X1 U10259 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n8921), .S(n8939), .Z(
        P2_U3446) );
  INV_X1 U10260 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n8923) );
  MUX2_X1 U10261 ( .A(n8923), .B(n8922), .S(n8939), .Z(n8924) );
  OAI21_X1 U10262 ( .B1(n8925), .B2(n8943), .A(n8924), .ZN(P2_U3444) );
  MUX2_X1 U10263 ( .A(n8927), .B(n8926), .S(n8939), .Z(n8928) );
  OAI21_X1 U10264 ( .B1(n8929), .B2(n8943), .A(n8928), .ZN(P2_U3441) );
  MUX2_X1 U10265 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n8930), .S(n8939), .Z(
        P2_U3438) );
  INV_X1 U10266 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n8932) );
  MUX2_X1 U10267 ( .A(n8932), .B(n8931), .S(n8939), .Z(n8933) );
  OAI21_X1 U10268 ( .B1(n8934), .B2(n8943), .A(n8933), .ZN(P2_U3435) );
  INV_X1 U10269 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n8936) );
  MUX2_X1 U10270 ( .A(n8936), .B(n8935), .S(n8939), .Z(n8937) );
  OAI21_X1 U10271 ( .B1(n8938), .B2(n8943), .A(n8937), .ZN(P2_U3432) );
  INV_X1 U10272 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n8941) );
  MUX2_X1 U10273 ( .A(n8941), .B(n8940), .S(n8939), .Z(n8942) );
  OAI21_X1 U10274 ( .B1(n8944), .B2(n8943), .A(n8942), .ZN(P2_U3429) );
  INV_X1 U10275 ( .A(n8945), .ZN(n9587) );
  NAND3_X1 U10276 ( .A1(n8947), .A2(P2_STATE_REG_SCAN_IN), .A3(
        P2_IR_REG_31__SCAN_IN), .ZN(n8948) );
  OAI22_X1 U10277 ( .A1(n8946), .A2(n8948), .B1(n6529), .B2(n8956), .ZN(n8949)
         );
  INV_X1 U10278 ( .A(n8949), .ZN(n8950) );
  OAI21_X1 U10279 ( .B1(n9587), .B2(n8960), .A(n8950), .ZN(P2_U3264) );
  NAND2_X1 U10280 ( .A1(n6351), .A2(n8953), .ZN(n8955) );
  OAI211_X1 U10281 ( .C1(n8957), .C2(n8956), .A(n8955), .B(n8954), .ZN(
        P2_U3267) );
  OAI222_X1 U10282 ( .A1(P2_U3151), .A2(n6004), .B1(n8960), .B2(n8959), .C1(
        n8958), .C2(n8956), .ZN(P2_U3268) );
  MUX2_X1 U10283 ( .A(n8962), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  XNOR2_X1 U10284 ( .A(n8963), .B(n9011), .ZN(n8965) );
  NOR2_X1 U10285 ( .A1(n8965), .A2(n8964), .ZN(n9010) );
  AOI21_X1 U10286 ( .B1(n8965), .B2(n8964), .A(n9010), .ZN(n8970) );
  AOI22_X1 U10287 ( .A1(n9104), .A2(n9392), .B1(P1_REG3_REG_14__SCAN_IN), .B2(
        P1_U3086), .ZN(n8967) );
  NAND2_X1 U10288 ( .A1(n9109), .A2(n9427), .ZN(n8966) );
  OAI211_X1 U10289 ( .C1(n9413), .C2(n9106), .A(n8967), .B(n8966), .ZN(n8968)
         );
  AOI21_X1 U10290 ( .B1(n9425), .B2(n9628), .A(n8968), .ZN(n8969) );
  OAI21_X1 U10291 ( .B1(n8970), .B2(n9623), .A(n8969), .ZN(P1_U3215) );
  AND3_X1 U10292 ( .A1(n9069), .A2(n9073), .A3(n8972), .ZN(n8973) );
  OAI21_X1 U10293 ( .B1(n8971), .B2(n8973), .A(n9102), .ZN(n8979) );
  NAND2_X1 U10294 ( .A1(n9122), .A2(n9393), .ZN(n8975) );
  OR2_X1 U10295 ( .A1(n9002), .A2(n9414), .ZN(n8974) );
  AND2_X1 U10296 ( .A1(n8975), .A2(n8974), .ZN(n9465) );
  OAI22_X1 U10297 ( .A1(n9465), .A2(n9095), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8976), .ZN(n8977) );
  AOI21_X1 U10298 ( .B1(n9289), .B2(n9109), .A(n8977), .ZN(n8978) );
  OAI211_X1 U10299 ( .C1(n9552), .C2(n9113), .A(n8979), .B(n8978), .ZN(
        P1_U3216) );
  XNOR2_X1 U10300 ( .A(n8980), .B(n8981), .ZN(n9082) );
  NOR2_X1 U10301 ( .A1(n9082), .A2(n9081), .ZN(n9080) );
  AOI21_X1 U10302 ( .B1(n8981), .B2(n8980), .A(n9080), .ZN(n8985) );
  XNOR2_X1 U10303 ( .A(n8983), .B(n8982), .ZN(n8984) );
  XNOR2_X1 U10304 ( .A(n8985), .B(n8984), .ZN(n8986) );
  NAND2_X1 U10305 ( .A1(n8986), .A2(n9102), .ZN(n8992) );
  NOR2_X1 U10306 ( .A1(n9106), .A2(n9375), .ZN(n8990) );
  OAI22_X1 U10307 ( .A1(n8988), .A2(n9343), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8987), .ZN(n8989) );
  AOI211_X1 U10308 ( .C1(n9109), .C2(n9346), .A(n8990), .B(n8989), .ZN(n8991)
         );
  OAI211_X1 U10309 ( .C1(n9349), .C2(n9113), .A(n8992), .B(n8991), .ZN(
        P1_U3219) );
  XOR2_X1 U10310 ( .A(n8994), .B(n8993), .Z(n8999) );
  OAI22_X1 U10311 ( .A1(n8995), .A2(n9414), .B1(n9343), .B2(n9412), .ZN(n9322)
         );
  AOI22_X1 U10312 ( .A1(n9322), .A2(n9618), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3086), .ZN(n8996) );
  OAI21_X1 U10313 ( .B1(n9315), .B2(n9631), .A(n8996), .ZN(n8997) );
  AOI21_X1 U10314 ( .B1(n9476), .B2(n9628), .A(n8997), .ZN(n8998) );
  OAI21_X1 U10315 ( .B1(n8999), .B2(n9623), .A(n8998), .ZN(P1_U3223) );
  AOI21_X1 U10316 ( .B1(n9001), .B2(n9000), .A(n9090), .ZN(n9009) );
  OR2_X1 U10317 ( .A1(n9002), .A2(n9412), .ZN(n9004) );
  NAND2_X1 U10318 ( .A1(n9118), .A2(n9390), .ZN(n9003) );
  AND2_X1 U10319 ( .A1(n9004), .A2(n9003), .ZN(n9257) );
  OAI22_X1 U10320 ( .A1(n9257), .A2(n9095), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9005), .ZN(n9007) );
  NOR2_X1 U10321 ( .A1(n9544), .A2(n9113), .ZN(n9006) );
  AOI211_X1 U10322 ( .C1(n9109), .C2(n9261), .A(n9007), .B(n9006), .ZN(n9008)
         );
  OAI21_X1 U10323 ( .B1(n9009), .B2(n9623), .A(n9008), .ZN(P1_U3225) );
  AOI21_X1 U10324 ( .B1(n9011), .B2(n8963), .A(n9010), .ZN(n9015) );
  XNOR2_X1 U10325 ( .A(n9015), .B(n9012), .ZN(n9100) );
  INV_X1 U10326 ( .A(n9013), .ZN(n9101) );
  NAND2_X1 U10327 ( .A1(n9100), .A2(n9101), .ZN(n9099) );
  OAI21_X1 U10328 ( .B1(n9015), .B2(n9014), .A(n9099), .ZN(n9020) );
  OAI21_X1 U10329 ( .B1(n9018), .B2(n9017), .A(n9016), .ZN(n9019) );
  XNOR2_X1 U10330 ( .A(n9020), .B(n9019), .ZN(n9025) );
  AOI22_X1 U10331 ( .A1(n9104), .A2(n9391), .B1(P1_REG3_REG_16__SCAN_IN), .B2(
        P1_U3086), .ZN(n9022) );
  NAND2_X1 U10332 ( .A1(n9109), .A2(n4944), .ZN(n9021) );
  OAI211_X1 U10333 ( .C1(n9415), .C2(n9106), .A(n9022), .B(n9021), .ZN(n9023)
         );
  AOI21_X1 U10334 ( .B1(n9399), .B2(n9628), .A(n9023), .ZN(n9024) );
  OAI21_X1 U10335 ( .B1(n9025), .B2(n9623), .A(n9024), .ZN(P1_U3226) );
  NAND2_X1 U10336 ( .A1(n9027), .A2(n9026), .ZN(n9028) );
  XNOR2_X1 U10337 ( .A(n9029), .B(n9028), .ZN(n9038) );
  AND2_X1 U10338 ( .A1(n9030), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9033) );
  NOR2_X1 U10339 ( .A1(n9631), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9032) );
  MUX2_X1 U10340 ( .A(n9033), .B(n9032), .S(n9031), .Z(n9036) );
  NAND2_X1 U10341 ( .A1(n9104), .A2(n9126), .ZN(n9034) );
  NAND2_X1 U10342 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9703) );
  OAI211_X1 U10343 ( .C1(n9373), .C2(n9106), .A(n9034), .B(n9703), .ZN(n9035)
         );
  AOI211_X1 U10344 ( .C1(n9504), .C2(n9628), .A(n9036), .B(n9035), .ZN(n9037)
         );
  OAI21_X1 U10345 ( .B1(n9038), .B2(n9623), .A(n9037), .ZN(P1_U3228) );
  INV_X1 U10346 ( .A(n9039), .ZN(n9043) );
  NOR3_X1 U10347 ( .A1(n8971), .A2(n9041), .A3(n9040), .ZN(n9042) );
  OAI21_X1 U10348 ( .B1(n9043), .B2(n9042), .A(n9102), .ZN(n9049) );
  OR2_X1 U10349 ( .A1(n9093), .A2(n9414), .ZN(n9045) );
  NAND2_X1 U10350 ( .A1(n9121), .A2(n9393), .ZN(n9044) );
  AND2_X1 U10351 ( .A1(n9045), .A2(n9044), .ZN(n9271) );
  OAI22_X1 U10352 ( .A1(n9271), .A2(n9095), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9046), .ZN(n9047) );
  AOI21_X1 U10353 ( .B1(n9278), .B2(n9109), .A(n9047), .ZN(n9048) );
  OAI211_X1 U10354 ( .C1(n9548), .C2(n9113), .A(n9049), .B(n9048), .ZN(
        P1_U3229) );
  XNOR2_X1 U10355 ( .A(n9051), .B(n9050), .ZN(n9052) );
  XNOR2_X1 U10356 ( .A(n9053), .B(n9052), .ZN(n9058) );
  AOI22_X1 U10357 ( .A1(n9123), .A2(n9390), .B1(n9125), .B2(n9393), .ZN(n9483)
         );
  OAI22_X1 U10358 ( .A1(n9483), .A2(n9095), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9054), .ZN(n9056) );
  NOR2_X1 U10359 ( .A1(n9561), .A2(n9113), .ZN(n9055) );
  AOI211_X1 U10360 ( .C1(n9109), .C2(n9331), .A(n9056), .B(n9055), .ZN(n9057)
         );
  OAI21_X1 U10361 ( .B1(n9058), .B2(n9623), .A(n9057), .ZN(P1_U3233) );
  XOR2_X1 U10362 ( .A(n9059), .B(n9060), .Z(n9068) );
  INV_X1 U10363 ( .A(n9061), .ZN(n9064) );
  AOI22_X1 U10364 ( .A1(n9062), .A2(n9618), .B1(P1_REG3_REG_13__SCAN_IN), .B2(
        P1_U3086), .ZN(n9063) );
  OAI21_X1 U10365 ( .B1(n9064), .B2(n9631), .A(n9063), .ZN(n9065) );
  AOI21_X1 U10366 ( .B1(n9066), .B2(n9628), .A(n9065), .ZN(n9067) );
  OAI21_X1 U10367 ( .B1(n9068), .B2(n9623), .A(n9067), .ZN(P1_U3234) );
  INV_X1 U10368 ( .A(n9069), .ZN(n9074) );
  AOI21_X1 U10369 ( .B1(n9071), .B2(n9073), .A(n9070), .ZN(n9072) );
  AOI21_X1 U10370 ( .B1(n9074), .B2(n9073), .A(n9072), .ZN(n9079) );
  NOR2_X1 U10371 ( .A1(n9631), .A2(n9304), .ZN(n9077) );
  AOI22_X1 U10372 ( .A1(n9123), .A2(n9393), .B1(n9121), .B2(n9390), .ZN(n9301)
         );
  INV_X1 U10373 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9075) );
  OAI22_X1 U10374 ( .A1(n9301), .A2(n9095), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9075), .ZN(n9076) );
  AOI211_X1 U10375 ( .C1(n9303), .C2(n9628), .A(n9077), .B(n9076), .ZN(n9078)
         );
  OAI21_X1 U10376 ( .B1(n9079), .B2(n9623), .A(n9078), .ZN(P1_U3235) );
  AOI21_X1 U10377 ( .B1(n9082), .B2(n9081), .A(n9080), .ZN(n9087) );
  AOI22_X1 U10378 ( .A1(n9393), .A2(n9391), .B1(n9125), .B2(n9390), .ZN(n9495)
         );
  OAI22_X1 U10379 ( .A1(n9495), .A2(n9095), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9083), .ZN(n9085) );
  NOR2_X1 U10380 ( .A1(n9566), .A2(n9113), .ZN(n9084) );
  AOI211_X1 U10381 ( .C1(n9109), .C2(n9356), .A(n9085), .B(n9084), .ZN(n9086)
         );
  OAI21_X1 U10382 ( .B1(n9087), .B2(n9623), .A(n9086), .ZN(P1_U3238) );
  OAI21_X1 U10383 ( .B1(n9090), .B2(n9089), .A(n9088), .ZN(n9091) );
  NAND3_X1 U10384 ( .A1(n9092), .A2(n9102), .A3(n9091), .ZN(n9098) );
  INV_X1 U10385 ( .A(n9093), .ZN(n9119) );
  AOI22_X1 U10386 ( .A1(n9393), .A2(n9119), .B1(n9117), .B2(n9390), .ZN(n9448)
         );
  OAI22_X1 U10387 ( .A1(n9448), .A2(n9095), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9094), .ZN(n9096) );
  AOI21_X1 U10388 ( .B1(n9243), .B2(n9109), .A(n9096), .ZN(n9097) );
  OAI211_X1 U10389 ( .C1(n9540), .C2(n9113), .A(n9098), .B(n9097), .ZN(
        P1_U3240) );
  OAI21_X1 U10390 ( .B1(n9101), .B2(n9100), .A(n9099), .ZN(n9103) );
  NAND2_X1 U10391 ( .A1(n9103), .A2(n9102), .ZN(n9112) );
  AOI22_X1 U10392 ( .A1(n9104), .A2(n9127), .B1(P1_REG3_REG_15__SCAN_IN), .B2(
        P1_U3086), .ZN(n9105) );
  OAI21_X1 U10393 ( .B1(n9107), .B2(n9106), .A(n9105), .ZN(n9108) );
  AOI21_X1 U10394 ( .B1(n9110), .B2(n9109), .A(n9108), .ZN(n9111) );
  OAI211_X1 U10395 ( .C1(n9114), .C2(n9113), .A(n9112), .B(n9111), .ZN(
        P1_U3241) );
  MUX2_X1 U10396 ( .A(n9115), .B(P1_DATAO_REG_30__SCAN_IN), .S(n9141), .Z(
        P1_U3584) );
  MUX2_X1 U10397 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9116), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U10398 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9117), .S(P1_U3973), .Z(
        P1_U3581) );
  MUX2_X1 U10399 ( .A(n9118), .B(P1_DATAO_REG_26__SCAN_IN), .S(n9141), .Z(
        P1_U3580) );
  MUX2_X1 U10400 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9119), .S(P1_U3973), .Z(
        P1_U3579) );
  MUX2_X1 U10401 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9120), .S(P1_U3973), .Z(
        P1_U3578) );
  MUX2_X1 U10402 ( .A(n9121), .B(P1_DATAO_REG_23__SCAN_IN), .S(n9141), .Z(
        P1_U3577) );
  MUX2_X1 U10403 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9122), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10404 ( .A(n9123), .B(P1_DATAO_REG_21__SCAN_IN), .S(n9141), .Z(
        P1_U3575) );
  MUX2_X1 U10405 ( .A(n9124), .B(P1_DATAO_REG_20__SCAN_IN), .S(n9141), .Z(
        P1_U3574) );
  MUX2_X1 U10406 ( .A(n9125), .B(P1_DATAO_REG_19__SCAN_IN), .S(n9141), .Z(
        P1_U3573) );
  MUX2_X1 U10407 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9126), .S(P1_U3973), .Z(
        P1_U3572) );
  MUX2_X1 U10408 ( .A(n9391), .B(P1_DATAO_REG_17__SCAN_IN), .S(n9141), .Z(
        P1_U3571) );
  MUX2_X1 U10409 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9127), .S(P1_U3973), .Z(
        P1_U3570) );
  MUX2_X1 U10410 ( .A(n9392), .B(P1_DATAO_REG_15__SCAN_IN), .S(n9141), .Z(
        P1_U3569) );
  MUX2_X1 U10411 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9128), .S(P1_U3973), .Z(
        P1_U3568) );
  MUX2_X1 U10412 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9129), .S(P1_U3973), .Z(
        P1_U3567) );
  MUX2_X1 U10413 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9130), .S(P1_U3973), .Z(
        P1_U3566) );
  MUX2_X1 U10414 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9131), .S(P1_U3973), .Z(
        P1_U3565) );
  MUX2_X1 U10415 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9132), .S(P1_U3973), .Z(
        P1_U3564) );
  MUX2_X1 U10416 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9133), .S(P1_U3973), .Z(
        P1_U3563) );
  MUX2_X1 U10417 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9134), .S(P1_U3973), .Z(
        P1_U3562) );
  MUX2_X1 U10418 ( .A(n9135), .B(P1_DATAO_REG_7__SCAN_IN), .S(n9141), .Z(
        P1_U3561) );
  MUX2_X1 U10419 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9136), .S(P1_U3973), .Z(
        P1_U3560) );
  MUX2_X1 U10420 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9137), .S(P1_U3973), .Z(
        P1_U3559) );
  MUX2_X1 U10421 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9138), .S(P1_U3973), .Z(
        P1_U3558) );
  MUX2_X1 U10422 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9139), .S(P1_U3973), .Z(
        P1_U3557) );
  MUX2_X1 U10423 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n9140), .S(P1_U3973), .Z(
        P1_U3556) );
  MUX2_X1 U10424 ( .A(n5737), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9141), .Z(
        P1_U3555) );
  MUX2_X1 U10425 ( .A(n5736), .B(P1_DATAO_REG_0__SCAN_IN), .S(n9141), .Z(
        P1_U3554) );
  INV_X1 U10426 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9143) );
  INV_X1 U10427 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n9142) );
  OAI22_X1 U10428 ( .A1(n9722), .A2(n9143), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9142), .ZN(n9144) );
  AOI21_X1 U10429 ( .B1(n9145), .B2(n9699), .A(n9144), .ZN(n9153) );
  OAI211_X1 U10430 ( .C1(n9148), .C2(n9147), .A(n9712), .B(n9146), .ZN(n9152)
         );
  INV_X1 U10431 ( .A(n9686), .ZN(n9708) );
  OAI211_X1 U10432 ( .C1(n9155), .C2(n9150), .A(n9708), .B(n9149), .ZN(n9151)
         );
  NAND3_X1 U10433 ( .A1(n9153), .A2(n9152), .A3(n9151), .ZN(P1_U3244) );
  MUX2_X1 U10434 ( .A(n9156), .B(n9155), .S(n9154), .Z(n9158) );
  NAND2_X1 U10435 ( .A1(n9158), .A2(n9157), .ZN(n9159) );
  OAI211_X1 U10436 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n9160), .A(n9159), .B(
        P1_U3973), .ZN(n9201) );
  INV_X1 U10437 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n9162) );
  INV_X1 U10438 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n9161) );
  OAI22_X1 U10439 ( .A1(n9722), .A2(n9162), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9161), .ZN(n9163) );
  AOI21_X1 U10440 ( .B1(n9164), .B2(n9699), .A(n9163), .ZN(n9173) );
  OAI211_X1 U10441 ( .C1(n9167), .C2(n9166), .A(n9708), .B(n9165), .ZN(n9172)
         );
  OAI211_X1 U10442 ( .C1(n9170), .C2(n9169), .A(n9712), .B(n9168), .ZN(n9171)
         );
  NAND4_X1 U10443 ( .A1(n9201), .A2(n9173), .A3(n9172), .A4(n9171), .ZN(
        P1_U3245) );
  INV_X1 U10444 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n9175) );
  NAND2_X1 U10445 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_U3086), .ZN(n9174) );
  OAI21_X1 U10446 ( .B1(n9722), .B2(n9175), .A(n9174), .ZN(n9176) );
  AOI21_X1 U10447 ( .B1(n9177), .B2(n9699), .A(n9176), .ZN(n9186) );
  OAI211_X1 U10448 ( .C1(n9180), .C2(n9179), .A(n9708), .B(n9178), .ZN(n9185)
         );
  OAI211_X1 U10449 ( .C1(n9183), .C2(n9182), .A(n9712), .B(n9181), .ZN(n9184)
         );
  NAND3_X1 U10450 ( .A1(n9186), .A2(n9185), .A3(n9184), .ZN(P1_U3246) );
  AOI21_X1 U10451 ( .B1(n9188), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n9187), .ZN(
        n9200) );
  OAI211_X1 U10452 ( .C1(n9191), .C2(n9190), .A(n9712), .B(n9189), .ZN(n9194)
         );
  NAND2_X1 U10453 ( .A1(n9699), .A2(n9192), .ZN(n9193) );
  AND2_X1 U10454 ( .A1(n9194), .A2(n9193), .ZN(n9199) );
  OAI211_X1 U10455 ( .C1(n9197), .C2(n9196), .A(n9708), .B(n9195), .ZN(n9198)
         );
  NAND4_X1 U10456 ( .A1(n9201), .A2(n9200), .A3(n9199), .A4(n9198), .ZN(
        P1_U3247) );
  NAND2_X1 U10457 ( .A1(n9435), .A2(n9326), .ZN(n9208) );
  INV_X1 U10458 ( .A(n9438), .ZN(n9206) );
  NOR2_X1 U10459 ( .A1(n9206), .A2(n9433), .ZN(n9210) );
  AOI21_X1 U10460 ( .B1(n9211), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9210), .ZN(
        n9207) );
  OAI211_X1 U10461 ( .C1(n4556), .C2(n9429), .A(n9208), .B(n9207), .ZN(
        P1_U3263) );
  XNOR2_X1 U10462 ( .A(n9532), .B(n9209), .ZN(n9439) );
  NAND2_X1 U10463 ( .A1(n9439), .A2(n9326), .ZN(n9213) );
  AOI21_X1 U10464 ( .B1(n9211), .B2(P1_REG2_REG_30__SCAN_IN), .A(n9210), .ZN(
        n9212) );
  OAI211_X1 U10465 ( .C1(n9532), .C2(n9429), .A(n9213), .B(n9212), .ZN(
        P1_U3264) );
  NAND2_X1 U10466 ( .A1(n9214), .A2(n9355), .ZN(n9222) );
  AOI22_X1 U10467 ( .A1(n9433), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n9215), .B2(
        n9426), .ZN(n9216) );
  OAI21_X1 U10468 ( .B1(n9217), .B2(n9433), .A(n9216), .ZN(n9220) );
  NOR2_X1 U10469 ( .A1(n9218), .A2(n9360), .ZN(n9219) );
  AOI211_X1 U10470 ( .C1(n9364), .C2(n4351), .A(n9220), .B(n9219), .ZN(n9221)
         );
  OAI211_X1 U10471 ( .C1(n9223), .C2(n9367), .A(n9222), .B(n9221), .ZN(
        P1_U3356) );
  XNOR2_X1 U10472 ( .A(n9224), .B(n9225), .ZN(n9444) );
  INV_X1 U10473 ( .A(n9444), .ZN(n9237) );
  XNOR2_X1 U10474 ( .A(n9226), .B(n9225), .ZN(n9227) );
  NAND2_X1 U10475 ( .A1(n9227), .A2(n9746), .ZN(n9229) );
  NAND2_X1 U10476 ( .A1(n9229), .A2(n9228), .ZN(n9442) );
  AOI211_X1 U10477 ( .C1(n9231), .C2(n9246), .A(n9422), .B(n9230), .ZN(n9443)
         );
  NAND2_X1 U10478 ( .A1(n9443), .A2(n9431), .ZN(n9234) );
  AOI22_X1 U10479 ( .A1(n9433), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n9232), .B2(
        n9426), .ZN(n9233) );
  OAI211_X1 U10480 ( .C1(n9536), .C2(n9429), .A(n9234), .B(n9233), .ZN(n9235)
         );
  AOI21_X1 U10481 ( .B1(n9442), .B2(n9381), .A(n9235), .ZN(n9236) );
  OAI21_X1 U10482 ( .B1(n9237), .B2(n9404), .A(n9236), .ZN(P1_U3266) );
  OAI21_X1 U10483 ( .B1(n9239), .B2(n9242), .A(n9238), .ZN(n9240) );
  INV_X1 U10484 ( .A(n9240), .ZN(n9449) );
  XOR2_X1 U10485 ( .A(n9242), .B(n9241), .Z(n9451) );
  NAND2_X1 U10486 ( .A1(n9451), .A2(n9355), .ZN(n9251) );
  AOI22_X1 U10487 ( .A1(n9433), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n9243), .B2(
        n9426), .ZN(n9244) );
  OAI21_X1 U10488 ( .B1(n9448), .B2(n9433), .A(n9244), .ZN(n9248) );
  INV_X1 U10489 ( .A(n9245), .ZN(n9259) );
  OAI211_X1 U10490 ( .C1(n9540), .C2(n9259), .A(n9246), .B(n9477), .ZN(n9447)
         );
  NOR2_X1 U10491 ( .A1(n9447), .A2(n9360), .ZN(n9247) );
  AOI211_X1 U10492 ( .C1(n9364), .C2(n9249), .A(n9248), .B(n9247), .ZN(n9250)
         );
  OAI211_X1 U10493 ( .C1(n9449), .C2(n9367), .A(n9251), .B(n9250), .ZN(
        P1_U3267) );
  XOR2_X1 U10494 ( .A(n9252), .B(n9254), .Z(n9456) );
  INV_X1 U10495 ( .A(n9456), .ZN(n9266) );
  NAND2_X1 U10496 ( .A1(n9268), .A2(n9253), .ZN(n9255) );
  XNOR2_X1 U10497 ( .A(n9255), .B(n9254), .ZN(n9256) );
  NAND2_X1 U10498 ( .A1(n9256), .A2(n9746), .ZN(n9258) );
  NAND2_X1 U10499 ( .A1(n9258), .A2(n9257), .ZN(n9454) );
  AOI211_X1 U10500 ( .C1(n9260), .C2(n9275), .A(n9422), .B(n9259), .ZN(n9455)
         );
  NAND2_X1 U10501 ( .A1(n9455), .A2(n9431), .ZN(n9263) );
  AOI22_X1 U10502 ( .A1(n9433), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n9261), .B2(
        n9426), .ZN(n9262) );
  OAI211_X1 U10503 ( .C1(n9544), .C2(n9429), .A(n9263), .B(n9262), .ZN(n9264)
         );
  AOI21_X1 U10504 ( .B1(n9381), .B2(n9454), .A(n9264), .ZN(n9265) );
  OAI21_X1 U10505 ( .B1(n9266), .B2(n9404), .A(n9265), .ZN(P1_U3268) );
  XNOR2_X1 U10506 ( .A(n9267), .B(n9269), .ZN(n9461) );
  INV_X1 U10507 ( .A(n9461), .ZN(n9283) );
  NAND2_X1 U10508 ( .A1(n9268), .A2(n9746), .ZN(n9273) );
  AOI21_X1 U10509 ( .B1(n9284), .B2(n9270), .A(n9269), .ZN(n9272) );
  OAI21_X1 U10510 ( .B1(n9273), .B2(n9272), .A(n9271), .ZN(n9459) );
  INV_X1 U10511 ( .A(n9274), .ZN(n9291) );
  INV_X1 U10512 ( .A(n9275), .ZN(n9276) );
  AOI211_X1 U10513 ( .C1(n9277), .C2(n9291), .A(n9422), .B(n9276), .ZN(n9460)
         );
  NAND2_X1 U10514 ( .A1(n9460), .A2(n9431), .ZN(n9280) );
  AOI22_X1 U10515 ( .A1(n9433), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n9278), .B2(
        n9426), .ZN(n9279) );
  OAI211_X1 U10516 ( .C1(n9548), .C2(n9429), .A(n9280), .B(n9279), .ZN(n9281)
         );
  AOI21_X1 U10517 ( .B1(n9381), .B2(n9459), .A(n9281), .ZN(n9282) );
  OAI21_X1 U10518 ( .B1(n9283), .B2(n9404), .A(n9282), .ZN(P1_U3269) );
  OAI21_X1 U10519 ( .B1(n9285), .B2(n9288), .A(n9284), .ZN(n9286) );
  INV_X1 U10520 ( .A(n9286), .ZN(n9466) );
  XOR2_X1 U10521 ( .A(n9288), .B(n9287), .Z(n9468) );
  NAND2_X1 U10522 ( .A1(n9468), .A2(n9355), .ZN(n9296) );
  AOI22_X1 U10523 ( .A1(n9211), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n9289), .B2(
        n9426), .ZN(n9290) );
  OAI21_X1 U10524 ( .B1(n9465), .B2(n9433), .A(n9290), .ZN(n9293) );
  OAI211_X1 U10525 ( .C1(n9552), .C2(n4441), .A(n9291), .B(n9477), .ZN(n9464)
         );
  NOR2_X1 U10526 ( .A1(n9464), .A2(n9360), .ZN(n9292) );
  AOI211_X1 U10527 ( .C1(n9364), .C2(n9294), .A(n9293), .B(n9292), .ZN(n9295)
         );
  OAI211_X1 U10528 ( .C1(n9466), .C2(n9367), .A(n9296), .B(n9295), .ZN(
        P1_U3270) );
  XNOR2_X1 U10529 ( .A(n9297), .B(n9298), .ZN(n9473) );
  INV_X1 U10530 ( .A(n9473), .ZN(n9310) );
  XNOR2_X1 U10531 ( .A(n9299), .B(n9298), .ZN(n9300) );
  NAND2_X1 U10532 ( .A1(n9300), .A2(n9746), .ZN(n9302) );
  NAND2_X1 U10533 ( .A1(n9302), .A2(n9301), .ZN(n9471) );
  AOI211_X1 U10534 ( .C1(n9303), .C2(n9313), .A(n9422), .B(n4441), .ZN(n9472)
         );
  NAND2_X1 U10535 ( .A1(n9472), .A2(n9431), .ZN(n9307) );
  INV_X1 U10536 ( .A(n9304), .ZN(n9305) );
  AOI22_X1 U10537 ( .A1(n9433), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n9305), .B2(
        n9426), .ZN(n9306) );
  OAI211_X1 U10538 ( .C1(n9556), .C2(n9429), .A(n9307), .B(n9306), .ZN(n9308)
         );
  AOI21_X1 U10539 ( .B1(n9381), .B2(n9471), .A(n9308), .ZN(n9309) );
  OAI21_X1 U10540 ( .B1(n9310), .B2(n9404), .A(n9309), .ZN(P1_U3271) );
  XOR2_X1 U10541 ( .A(n9311), .B(n9320), .Z(n9481) );
  INV_X1 U10542 ( .A(n9313), .ZN(n9314) );
  AOI21_X1 U10543 ( .B1(n9476), .B2(n9333), .A(n9314), .ZN(n9478) );
  INV_X1 U10544 ( .A(n9315), .ZN(n9316) );
  AOI22_X1 U10545 ( .A1(n9211), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n9316), .B2(
        n9426), .ZN(n9317) );
  OAI21_X1 U10546 ( .B1(n9318), .B2(n9429), .A(n9317), .ZN(n9325) );
  OAI21_X1 U10547 ( .B1(n9321), .B2(n9320), .A(n9319), .ZN(n9323) );
  AOI21_X1 U10548 ( .B1(n9323), .B2(n9746), .A(n9322), .ZN(n9480) );
  NOR2_X1 U10549 ( .A1(n9480), .A2(n9433), .ZN(n9324) );
  AOI211_X1 U10550 ( .C1(n9478), .C2(n9326), .A(n9325), .B(n9324), .ZN(n9327)
         );
  OAI21_X1 U10551 ( .B1(n9481), .B2(n9404), .A(n9327), .ZN(P1_U3272) );
  XNOR2_X1 U10552 ( .A(n9328), .B(n9329), .ZN(n9484) );
  XOR2_X1 U10553 ( .A(n9330), .B(n9329), .Z(n9486) );
  NAND2_X1 U10554 ( .A1(n9486), .A2(n9355), .ZN(n9338) );
  AOI22_X1 U10555 ( .A1(n9433), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9331), .B2(
        n9426), .ZN(n9332) );
  OAI21_X1 U10556 ( .B1(n9483), .B2(n9433), .A(n9332), .ZN(n9335) );
  OAI211_X1 U10557 ( .C1(n9345), .C2(n9561), .A(n9477), .B(n9333), .ZN(n9482)
         );
  NOR2_X1 U10558 ( .A1(n9482), .A2(n9360), .ZN(n9334) );
  AOI211_X1 U10559 ( .C1(n9364), .C2(n9336), .A(n9335), .B(n9334), .ZN(n9337)
         );
  OAI211_X1 U10560 ( .C1(n9484), .C2(n9367), .A(n9338), .B(n9337), .ZN(
        P1_U3273) );
  XOR2_X1 U10561 ( .A(n9339), .B(n9341), .Z(n9493) );
  XOR2_X1 U10562 ( .A(n9340), .B(n9341), .Z(n9342) );
  OAI222_X1 U10563 ( .A1(n9414), .A2(n9343), .B1(n9412), .B2(n9375), .C1(n9496), .C2(n9342), .ZN(n9489) );
  INV_X1 U10564 ( .A(n9344), .ZN(n9359) );
  AOI211_X1 U10565 ( .C1(n9491), .C2(n9359), .A(n9422), .B(n9345), .ZN(n9490)
         );
  NAND2_X1 U10566 ( .A1(n9490), .A2(n9431), .ZN(n9348) );
  AOI22_X1 U10567 ( .A1(n9433), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9346), .B2(
        n9426), .ZN(n9347) );
  OAI211_X1 U10568 ( .C1(n9349), .C2(n9429), .A(n9348), .B(n9347), .ZN(n9350)
         );
  AOI21_X1 U10569 ( .B1(n9489), .B2(n9381), .A(n9350), .ZN(n9351) );
  OAI21_X1 U10570 ( .B1(n9493), .B2(n9404), .A(n9351), .ZN(P1_U3274) );
  XNOR2_X1 U10571 ( .A(n9352), .B(n9353), .ZN(n9497) );
  XNOR2_X1 U10572 ( .A(n9354), .B(n9353), .ZN(n9499) );
  NAND2_X1 U10573 ( .A1(n9499), .A2(n9355), .ZN(n9366) );
  AOI22_X1 U10574 ( .A1(n9433), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9356), .B2(
        n9426), .ZN(n9357) );
  OAI21_X1 U10575 ( .B1(n9495), .B2(n9433), .A(n9357), .ZN(n9362) );
  INV_X1 U10576 ( .A(n9358), .ZN(n9376) );
  OAI211_X1 U10577 ( .C1(n9566), .C2(n9376), .A(n9359), .B(n9477), .ZN(n9494)
         );
  NOR2_X1 U10578 ( .A1(n9494), .A2(n9360), .ZN(n9361) );
  AOI211_X1 U10579 ( .C1(n9364), .C2(n9363), .A(n9362), .B(n9361), .ZN(n9365)
         );
  OAI211_X1 U10580 ( .C1(n9497), .C2(n9367), .A(n9366), .B(n9365), .ZN(
        P1_U3275) );
  XNOR2_X1 U10581 ( .A(n9369), .B(n9368), .ZN(n9506) );
  NAND2_X1 U10582 ( .A1(n9388), .A2(n9370), .ZN(n9372) );
  XNOR2_X1 U10583 ( .A(n9372), .B(n9371), .ZN(n9374) );
  OAI222_X1 U10584 ( .A1(n9414), .A2(n9375), .B1(n9374), .B2(n9496), .C1(n9412), .C2(n9373), .ZN(n9502) );
  AOI211_X1 U10585 ( .C1(n9504), .C2(n9397), .A(n9422), .B(n9376), .ZN(n9503)
         );
  NAND2_X1 U10586 ( .A1(n9503), .A2(n9431), .ZN(n9379) );
  AOI22_X1 U10587 ( .A1(n9433), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9377), .B2(
        n9426), .ZN(n9378) );
  OAI211_X1 U10588 ( .C1(n4565), .C2(n9429), .A(n9379), .B(n9378), .ZN(n9380)
         );
  AOI21_X1 U10589 ( .B1(n9381), .B2(n9502), .A(n9380), .ZN(n9382) );
  OAI21_X1 U10590 ( .B1(n9506), .B2(n9404), .A(n9382), .ZN(P1_U3276) );
  XNOR2_X1 U10591 ( .A(n9383), .B(n9384), .ZN(n9509) );
  INV_X1 U10592 ( .A(n9509), .ZN(n9405) );
  NAND2_X1 U10593 ( .A1(n9386), .A2(n9385), .ZN(n9387) );
  NAND2_X1 U10594 ( .A1(n9388), .A2(n9387), .ZN(n9389) );
  NAND2_X1 U10595 ( .A1(n9389), .A2(n9746), .ZN(n9395) );
  AOI22_X1 U10596 ( .A1(n9393), .A2(n9392), .B1(n9391), .B2(n9390), .ZN(n9394)
         );
  NAND2_X1 U10597 ( .A1(n9395), .A2(n9394), .ZN(n9507) );
  INV_X1 U10598 ( .A(n9397), .ZN(n9398) );
  AOI211_X1 U10599 ( .C1(n9399), .C2(n4569), .A(n9422), .B(n9398), .ZN(n9508)
         );
  NAND2_X1 U10600 ( .A1(n9508), .A2(n9431), .ZN(n9401) );
  AOI22_X1 U10601 ( .A1(n9433), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n4944), .B2(
        n9426), .ZN(n9400) );
  OAI211_X1 U10602 ( .C1(n9571), .C2(n9429), .A(n9401), .B(n9400), .ZN(n9402)
         );
  AOI21_X1 U10603 ( .B1(n9381), .B2(n9507), .A(n9402), .ZN(n9403) );
  OAI21_X1 U10604 ( .B1(n9405), .B2(n9404), .A(n9403), .ZN(P1_U3277) );
  INV_X1 U10605 ( .A(n9406), .ZN(n9420) );
  OAI21_X1 U10606 ( .B1(n9407), .B2(n9409), .A(n9408), .ZN(n9520) );
  INV_X1 U10607 ( .A(n9520), .ZN(n9419) );
  OAI21_X1 U10608 ( .B1(n4826), .B2(n9411), .A(n9410), .ZN(n9417) );
  OAI22_X1 U10609 ( .A1(n9415), .A2(n9414), .B1(n9413), .B2(n9412), .ZN(n9416)
         );
  AOI21_X1 U10610 ( .B1(n9417), .B2(n9746), .A(n9416), .ZN(n9418) );
  OAI21_X1 U10611 ( .B1(n9419), .B2(n9741), .A(n9418), .ZN(n9518) );
  AOI21_X1 U10612 ( .B1(n9420), .B2(n9520), .A(n9518), .ZN(n9434) );
  INV_X1 U10613 ( .A(n9421), .ZN(n9423) );
  AOI211_X1 U10614 ( .C1(n9425), .C2(n9424), .A(n9423), .B(n9422), .ZN(n9519)
         );
  AOI22_X1 U10615 ( .A1(n9433), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n9427), .B2(
        n9426), .ZN(n9428) );
  OAI21_X1 U10616 ( .B1(n4832), .B2(n9429), .A(n9428), .ZN(n9430) );
  AOI21_X1 U10617 ( .B1(n9519), .B2(n9431), .A(n9430), .ZN(n9432) );
  OAI21_X1 U10618 ( .B1(n9434), .B2(n9433), .A(n9432), .ZN(P1_U3279) );
  INV_X1 U10619 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9436) );
  MUX2_X1 U10620 ( .A(n9436), .B(n9526), .S(n9757), .Z(n9437) );
  OAI21_X1 U10621 ( .B1(n4556), .B2(n9524), .A(n9437), .ZN(P1_U3553) );
  INV_X1 U10622 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9440) );
  AOI21_X1 U10623 ( .B1(n9439), .B2(n9477), .A(n9438), .ZN(n9529) );
  MUX2_X1 U10624 ( .A(n9440), .B(n9529), .S(n9757), .Z(n9441) );
  OAI21_X1 U10625 ( .B1(n9532), .B2(n9524), .A(n9441), .ZN(P1_U3552) );
  INV_X1 U10626 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n9445) );
  MUX2_X1 U10627 ( .A(n9445), .B(n9533), .S(n9757), .Z(n9446) );
  OAI21_X1 U10628 ( .B1(n9536), .B2(n9524), .A(n9446), .ZN(P1_U3549) );
  INV_X1 U10629 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n9452) );
  OAI211_X1 U10630 ( .C1(n9449), .C2(n9496), .A(n9448), .B(n9447), .ZN(n9450)
         );
  AOI21_X1 U10631 ( .B1(n9451), .B2(n9734), .A(n9450), .ZN(n9537) );
  MUX2_X1 U10632 ( .A(n9452), .B(n9537), .S(n9757), .Z(n9453) );
  OAI21_X1 U10633 ( .B1(n9540), .B2(n9524), .A(n9453), .ZN(P1_U3548) );
  INV_X1 U10634 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n9457) );
  AOI211_X1 U10635 ( .C1(n9456), .C2(n9734), .A(n9455), .B(n9454), .ZN(n9541)
         );
  MUX2_X1 U10636 ( .A(n9457), .B(n9541), .S(n9757), .Z(n9458) );
  OAI21_X1 U10637 ( .B1(n9544), .B2(n9524), .A(n9458), .ZN(P1_U3547) );
  INV_X1 U10638 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n9462) );
  AOI211_X1 U10639 ( .C1(n9461), .C2(n9734), .A(n9460), .B(n9459), .ZN(n9545)
         );
  MUX2_X1 U10640 ( .A(n9462), .B(n9545), .S(n9757), .Z(n9463) );
  OAI21_X1 U10641 ( .B1(n9548), .B2(n9524), .A(n9463), .ZN(P1_U3546) );
  INV_X1 U10642 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n9469) );
  OAI211_X1 U10643 ( .C1(n9466), .C2(n9496), .A(n9465), .B(n9464), .ZN(n9467)
         );
  AOI21_X1 U10644 ( .B1(n9468), .B2(n9734), .A(n9467), .ZN(n9549) );
  MUX2_X1 U10645 ( .A(n9469), .B(n9549), .S(n9757), .Z(n9470) );
  OAI21_X1 U10646 ( .B1(n9552), .B2(n9524), .A(n9470), .ZN(P1_U3545) );
  INV_X1 U10647 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n9474) );
  AOI211_X1 U10648 ( .C1(n9473), .C2(n9734), .A(n9472), .B(n9471), .ZN(n9553)
         );
  MUX2_X1 U10649 ( .A(n9474), .B(n9553), .S(n9757), .Z(n9475) );
  OAI21_X1 U10650 ( .B1(n9556), .B2(n9524), .A(n9475), .ZN(P1_U3544) );
  AOI22_X1 U10651 ( .A1(n9478), .A2(n9477), .B1(n9724), .B2(n9476), .ZN(n9479)
         );
  OAI211_X1 U10652 ( .C1(n9481), .C2(n9516), .A(n9480), .B(n9479), .ZN(n9557)
         );
  MUX2_X1 U10653 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9557), .S(n9757), .Z(
        P1_U3543) );
  INV_X1 U10654 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n9487) );
  OAI211_X1 U10655 ( .C1(n9484), .C2(n9496), .A(n9483), .B(n9482), .ZN(n9485)
         );
  AOI21_X1 U10656 ( .B1(n9486), .B2(n9734), .A(n9485), .ZN(n9558) );
  MUX2_X1 U10657 ( .A(n9487), .B(n9558), .S(n9757), .Z(n9488) );
  OAI21_X1 U10658 ( .B1(n9561), .B2(n9524), .A(n9488), .ZN(P1_U3542) );
  AOI211_X1 U10659 ( .C1(n9724), .C2(n9491), .A(n9490), .B(n9489), .ZN(n9492)
         );
  OAI21_X1 U10660 ( .B1(n9493), .B2(n9516), .A(n9492), .ZN(n9562) );
  MUX2_X1 U10661 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9562), .S(n9757), .Z(
        P1_U3541) );
  INV_X1 U10662 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9500) );
  OAI211_X1 U10663 ( .C1(n9497), .C2(n9496), .A(n9495), .B(n9494), .ZN(n9498)
         );
  AOI21_X1 U10664 ( .B1(n9499), .B2(n9734), .A(n9498), .ZN(n9563) );
  MUX2_X1 U10665 ( .A(n9500), .B(n9563), .S(n9757), .Z(n9501) );
  OAI21_X1 U10666 ( .B1(n9566), .B2(n9524), .A(n9501), .ZN(P1_U3540) );
  AOI211_X1 U10667 ( .C1(n9724), .C2(n9504), .A(n9503), .B(n9502), .ZN(n9505)
         );
  OAI21_X1 U10668 ( .B1(n9506), .B2(n9516), .A(n9505), .ZN(n9567) );
  MUX2_X1 U10669 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9567), .S(n9757), .Z(
        P1_U3539) );
  AOI211_X1 U10670 ( .C1(n9509), .C2(n9734), .A(n9508), .B(n9507), .ZN(n9568)
         );
  MUX2_X1 U10671 ( .A(n9510), .B(n9568), .S(n9757), .Z(n9511) );
  OAI21_X1 U10672 ( .B1(n9571), .B2(n9524), .A(n9511), .ZN(P1_U3538) );
  AOI211_X1 U10673 ( .C1(n9724), .C2(n9514), .A(n9513), .B(n9512), .ZN(n9515)
         );
  OAI21_X1 U10674 ( .B1(n9517), .B2(n9516), .A(n9515), .ZN(n9572) );
  MUX2_X1 U10675 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9572), .S(n9757), .Z(
        P1_U3537) );
  INV_X1 U10676 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9522) );
  INV_X1 U10677 ( .A(n9742), .ZN(n9521) );
  AOI211_X1 U10678 ( .C1(n9521), .C2(n9520), .A(n9519), .B(n9518), .ZN(n9573)
         );
  MUX2_X1 U10679 ( .A(n9522), .B(n9573), .S(n9757), .Z(n9523) );
  OAI21_X1 U10680 ( .B1(n4832), .B2(n9524), .A(n9523), .ZN(P1_U3536) );
  MUX2_X1 U10681 ( .A(n9525), .B(P1_REG1_REG_0__SCAN_IN), .S(n9754), .Z(
        P1_U3522) );
  INV_X1 U10682 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n9527) );
  MUX2_X1 U10683 ( .A(n9527), .B(n9526), .S(n9749), .Z(n9528) );
  OAI21_X1 U10684 ( .B1(n4556), .B2(n9576), .A(n9528), .ZN(P1_U3521) );
  INV_X1 U10685 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9530) );
  MUX2_X1 U10686 ( .A(n9530), .B(n9529), .S(n9749), .Z(n9531) );
  OAI21_X1 U10687 ( .B1(n9532), .B2(n9576), .A(n9531), .ZN(P1_U3520) );
  INV_X1 U10688 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n9534) );
  MUX2_X1 U10689 ( .A(n9534), .B(n9533), .S(n9749), .Z(n9535) );
  OAI21_X1 U10690 ( .B1(n9536), .B2(n9576), .A(n9535), .ZN(P1_U3517) );
  INV_X1 U10691 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n9538) );
  MUX2_X1 U10692 ( .A(n9538), .B(n9537), .S(n9749), .Z(n9539) );
  OAI21_X1 U10693 ( .B1(n9540), .B2(n9576), .A(n9539), .ZN(P1_U3516) );
  INV_X1 U10694 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n9542) );
  MUX2_X1 U10695 ( .A(n9542), .B(n9541), .S(n9749), .Z(n9543) );
  OAI21_X1 U10696 ( .B1(n9544), .B2(n9576), .A(n9543), .ZN(P1_U3515) );
  INV_X1 U10697 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n9546) );
  MUX2_X1 U10698 ( .A(n9546), .B(n9545), .S(n9749), .Z(n9547) );
  OAI21_X1 U10699 ( .B1(n9548), .B2(n9576), .A(n9547), .ZN(P1_U3514) );
  INV_X1 U10700 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n9550) );
  MUX2_X1 U10701 ( .A(n9550), .B(n9549), .S(n9749), .Z(n9551) );
  OAI21_X1 U10702 ( .B1(n9552), .B2(n9576), .A(n9551), .ZN(P1_U3513) );
  INV_X1 U10703 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n9554) );
  MUX2_X1 U10704 ( .A(n9554), .B(n9553), .S(n9749), .Z(n9555) );
  OAI21_X1 U10705 ( .B1(n9556), .B2(n9576), .A(n9555), .ZN(P1_U3512) );
  MUX2_X1 U10706 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9557), .S(n9749), .Z(
        P1_U3511) );
  INV_X1 U10707 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n9559) );
  MUX2_X1 U10708 ( .A(n9559), .B(n9558), .S(n9749), .Z(n9560) );
  OAI21_X1 U10709 ( .B1(n9561), .B2(n9576), .A(n9560), .ZN(P1_U3510) );
  MUX2_X1 U10710 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9562), .S(n9749), .Z(
        P1_U3509) );
  INV_X1 U10711 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n9564) );
  MUX2_X1 U10712 ( .A(n9564), .B(n9563), .S(n9749), .Z(n9565) );
  OAI21_X1 U10713 ( .B1(n9566), .B2(n9576), .A(n9565), .ZN(P1_U3507) );
  MUX2_X1 U10714 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9567), .S(n9749), .Z(
        P1_U3504) );
  INV_X1 U10715 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n9569) );
  MUX2_X1 U10716 ( .A(n9569), .B(n9568), .S(n9749), .Z(n9570) );
  OAI21_X1 U10717 ( .B1(n9571), .B2(n9576), .A(n9570), .ZN(P1_U3501) );
  MUX2_X1 U10718 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n9572), .S(n9749), .Z(
        P1_U3498) );
  INV_X1 U10719 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n9574) );
  MUX2_X1 U10720 ( .A(n9574), .B(n9573), .S(n9749), .Z(n9575) );
  OAI21_X1 U10721 ( .B1(n4832), .B2(n9576), .A(n9575), .ZN(P1_U3495) );
  MUX2_X1 U10722 ( .A(n9579), .B(P1_D_REG_1__SCAN_IN), .S(n4349), .Z(P1_U3440)
         );
  MUX2_X1 U10723 ( .A(n9580), .B(P1_D_REG_0__SCAN_IN), .S(n4349), .Z(P1_U3439)
         );
  INV_X1 U10724 ( .A(n9581), .ZN(n9583) );
  NOR4_X1 U10725 ( .A1(n9583), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3086), .A4(
        n5010), .ZN(n9584) );
  AOI21_X1 U10726 ( .B1(n9585), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9584), .ZN(
        n9586) );
  OAI21_X1 U10727 ( .B1(n9587), .B2(n9591), .A(n9586), .ZN(P1_U3324) );
  OAI222_X1 U10728 ( .A1(n9591), .A2(n8951), .B1(n9590), .B2(P1_U3086), .C1(
        n9589), .C2(n9588), .ZN(P1_U3326) );
  MUX2_X1 U10729 ( .A(n9592), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U10730 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n9603) );
  AOI211_X1 U10731 ( .C1(n9595), .C2(n9594), .A(n9593), .B(n9686), .ZN(n9600)
         );
  AOI211_X1 U10732 ( .C1(n9598), .C2(n9597), .A(n9596), .B(n9669), .ZN(n9599)
         );
  AOI211_X1 U10733 ( .C1(n9699), .C2(n9601), .A(n9600), .B(n9599), .ZN(n9602)
         );
  NAND2_X1 U10734 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n9616) );
  OAI211_X1 U10735 ( .C1(n9722), .C2(n9603), .A(n9602), .B(n9616), .ZN(
        P1_U3253) );
  INV_X1 U10736 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n9615) );
  OAI21_X1 U10737 ( .B1(n9606), .B2(n9605), .A(n9604), .ZN(n9612) );
  OAI21_X1 U10738 ( .B1(n9609), .B2(n9608), .A(n9607), .ZN(n9610) );
  AOI222_X1 U10739 ( .A1(n9612), .A2(n9708), .B1(n9611), .B2(n9699), .C1(n9610), .C2(n9712), .ZN(n9614) );
  OAI211_X1 U10740 ( .C1(n9722), .C2(n9615), .A(n9614), .B(n9613), .ZN(
        P1_U3252) );
  INV_X1 U10741 ( .A(n9616), .ZN(n9617) );
  AOI21_X1 U10742 ( .B1(n9619), .B2(n9618), .A(n9617), .ZN(n9620) );
  INV_X1 U10743 ( .A(n9620), .ZN(n9627) );
  NAND2_X1 U10744 ( .A1(n9622), .A2(n9621), .ZN(n9624) );
  AOI21_X1 U10745 ( .B1(n9625), .B2(n9624), .A(n9623), .ZN(n9626) );
  AOI211_X1 U10746 ( .C1(n9629), .C2(n9628), .A(n9627), .B(n9626), .ZN(n9630)
         );
  OAI21_X1 U10747 ( .B1(n9632), .B2(n9631), .A(n9630), .ZN(P1_U3217) );
  XNOR2_X1 U10748 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  INV_X1 U10749 ( .A(P2_RD_REG_SCAN_IN), .ZN(n10096) );
  XOR2_X1 U10750 ( .A(P1_RD_REG_SCAN_IN), .B(n10096), .Z(U126) );
  INV_X1 U10751 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n9644) );
  AOI211_X1 U10752 ( .C1(n9635), .C2(n9634), .A(n9633), .B(n9686), .ZN(n9640)
         );
  AOI211_X1 U10753 ( .C1(n9638), .C2(n9637), .A(n9636), .B(n9669), .ZN(n9639)
         );
  AOI211_X1 U10754 ( .C1(n9699), .C2(n9641), .A(n9640), .B(n9639), .ZN(n9643)
         );
  NAND2_X1 U10755 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n9642) );
  OAI211_X1 U10756 ( .C1(n9722), .C2(n9644), .A(n9643), .B(n9642), .ZN(
        P1_U3254) );
  INV_X1 U10757 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n9656) );
  AOI211_X1 U10758 ( .C1(n9647), .C2(n9646), .A(n9645), .B(n9669), .ZN(n9652)
         );
  AOI211_X1 U10759 ( .C1(n9650), .C2(n9649), .A(n9648), .B(n9686), .ZN(n9651)
         );
  AOI211_X1 U10760 ( .C1(n9699), .C2(n9653), .A(n9652), .B(n9651), .ZN(n9655)
         );
  NAND2_X1 U10761 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n9654) );
  OAI211_X1 U10762 ( .C1(n9722), .C2(n9656), .A(n9655), .B(n9654), .ZN(
        P1_U3256) );
  INV_X1 U10763 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n9668) );
  AOI211_X1 U10764 ( .C1(n9659), .C2(n9658), .A(n9657), .B(n9686), .ZN(n9664)
         );
  AOI211_X1 U10765 ( .C1(n9662), .C2(n9661), .A(n9660), .B(n9669), .ZN(n9663)
         );
  AOI211_X1 U10766 ( .C1(n9699), .C2(n9665), .A(n9664), .B(n9663), .ZN(n9667)
         );
  NAND2_X1 U10767 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n9666) );
  OAI211_X1 U10768 ( .C1(n9722), .C2(n9668), .A(n9667), .B(n9666), .ZN(
        P1_U3257) );
  INV_X1 U10769 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n9681) );
  AOI211_X1 U10770 ( .C1(n9672), .C2(n9671), .A(n9670), .B(n9669), .ZN(n9677)
         );
  AOI211_X1 U10771 ( .C1(n9675), .C2(n9674), .A(n9673), .B(n9686), .ZN(n9676)
         );
  AOI211_X1 U10772 ( .C1(n9699), .C2(n9678), .A(n9677), .B(n9676), .ZN(n9680)
         );
  NAND2_X1 U10773 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_U3086), .ZN(n9679) );
  OAI211_X1 U10774 ( .C1(n9722), .C2(n9681), .A(n9680), .B(n9679), .ZN(
        P1_U3258) );
  INV_X1 U10775 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n9894) );
  OAI21_X1 U10776 ( .B1(n9684), .B2(n9683), .A(n9682), .ZN(n9692) );
  NOR2_X1 U10777 ( .A1(n9718), .A2(n9685), .ZN(n9691) );
  AOI211_X1 U10778 ( .C1(n9689), .C2(n9688), .A(n9687), .B(n9686), .ZN(n9690)
         );
  AOI211_X1 U10779 ( .C1(n9712), .C2(n9692), .A(n9691), .B(n9690), .ZN(n9694)
         );
  NAND2_X1 U10780 ( .A1(P1_REG3_REG_16__SCAN_IN), .A2(P1_U3086), .ZN(n9693) );
  OAI211_X1 U10781 ( .C1(n9722), .C2(n9894), .A(n9694), .B(n9693), .ZN(
        P1_U3259) );
  INV_X1 U10782 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9705) );
  XNOR2_X1 U10783 ( .A(n9696), .B(n9695), .ZN(n9702) );
  XNOR2_X1 U10784 ( .A(n9698), .B(n9697), .ZN(n9701) );
  AOI222_X1 U10785 ( .A1(n9702), .A2(n9708), .B1(n9712), .B2(n9701), .C1(n9700), .C2(n9699), .ZN(n9704) );
  OAI211_X1 U10786 ( .C1(n9722), .C2(n9705), .A(n9704), .B(n9703), .ZN(
        P1_U3260) );
  INV_X1 U10787 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n9938) );
  INV_X1 U10788 ( .A(n9706), .ZN(n9717) );
  OAI211_X1 U10789 ( .C1(n9710), .C2(n9709), .A(n9708), .B(n9707), .ZN(n9716)
         );
  OAI211_X1 U10790 ( .C1(n9714), .C2(n9713), .A(n9712), .B(n9711), .ZN(n9715)
         );
  OAI211_X1 U10791 ( .C1(n9718), .C2(n9717), .A(n9716), .B(n9715), .ZN(n9719)
         );
  INV_X1 U10792 ( .A(n9719), .ZN(n9721) );
  NAND2_X1 U10793 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_U3086), .ZN(n9720) );
  OAI211_X1 U10794 ( .C1(n9722), .C2(n9938), .A(n9721), .B(n9720), .ZN(
        P1_U3261) );
  AND2_X1 U10795 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n4349), .ZN(P1_U3294) );
  AND2_X1 U10796 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n4349), .ZN(P1_U3295) );
  AND2_X1 U10797 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n4349), .ZN(P1_U3296) );
  AND2_X1 U10798 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n4349), .ZN(P1_U3297) );
  AND2_X1 U10799 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n4349), .ZN(P1_U3298) );
  AND2_X1 U10800 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n4349), .ZN(P1_U3299) );
  AND2_X1 U10801 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n4349), .ZN(P1_U3300) );
  AND2_X1 U10802 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n4349), .ZN(P1_U3301) );
  AND2_X1 U10803 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n4349), .ZN(P1_U3302) );
  AND2_X1 U10804 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n4349), .ZN(P1_U3303) );
  AND2_X1 U10805 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n4349), .ZN(P1_U3304) );
  AND2_X1 U10806 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n4349), .ZN(P1_U3305) );
  AND2_X1 U10807 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n4349), .ZN(P1_U3306) );
  AND2_X1 U10808 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n4349), .ZN(P1_U3307) );
  AND2_X1 U10809 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n4349), .ZN(P1_U3308) );
  AND2_X1 U10810 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n4349), .ZN(P1_U3309) );
  AND2_X1 U10811 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n4349), .ZN(P1_U3310) );
  AND2_X1 U10812 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n4349), .ZN(P1_U3311) );
  AND2_X1 U10813 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n4349), .ZN(P1_U3312) );
  AND2_X1 U10814 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n4349), .ZN(P1_U3313) );
  AND2_X1 U10815 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n4349), .ZN(P1_U3314) );
  AND2_X1 U10816 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n4349), .ZN(P1_U3315) );
  AND2_X1 U10817 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n4349), .ZN(P1_U3316) );
  AND2_X1 U10818 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n4349), .ZN(P1_U3317) );
  AND2_X1 U10819 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n4349), .ZN(P1_U3318) );
  AND2_X1 U10820 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n4349), .ZN(P1_U3319) );
  AND2_X1 U10821 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n4349), .ZN(P1_U3320) );
  AND2_X1 U10822 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n4349), .ZN(P1_U3321) );
  AND2_X1 U10823 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n4349), .ZN(P1_U3322) );
  AND2_X1 U10824 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n4349), .ZN(P1_U3323) );
  INV_X1 U10825 ( .A(n9724), .ZN(n9738) );
  OAI21_X1 U10826 ( .B1(n5821), .B2(n9738), .A(n9725), .ZN(n9727) );
  AOI211_X1 U10827 ( .C1(n9734), .C2(n9728), .A(n9727), .B(n9726), .ZN(n9751)
         );
  INV_X1 U10828 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9729) );
  AOI22_X1 U10829 ( .A1(n9749), .A2(n9751), .B1(n9729), .B2(n9747), .ZN(
        P1_U3456) );
  OAI21_X1 U10830 ( .B1(n5740), .B2(n9738), .A(n9730), .ZN(n9732) );
  AOI211_X1 U10831 ( .C1(n9734), .C2(n9733), .A(n9732), .B(n9731), .ZN(n9753)
         );
  INV_X1 U10832 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n9735) );
  AOI22_X1 U10833 ( .A1(n9749), .A2(n9753), .B1(n9735), .B2(n9747), .ZN(
        P1_U3462) );
  OAI211_X1 U10834 ( .C1(n9739), .C2(n9738), .A(n9737), .B(n9736), .ZN(n9744)
         );
  AOI21_X1 U10835 ( .B1(n9742), .B2(n9741), .A(n9740), .ZN(n9743) );
  AOI211_X1 U10836 ( .C1(n9746), .C2(n9745), .A(n9744), .B(n9743), .ZN(n9756)
         );
  INV_X1 U10837 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9748) );
  AOI22_X1 U10838 ( .A1(n9749), .A2(n9756), .B1(n9748), .B2(n9747), .ZN(
        P1_U3474) );
  AOI22_X1 U10839 ( .A1(n9757), .A2(n9751), .B1(n9750), .B2(n9754), .ZN(
        P1_U3523) );
  INV_X1 U10840 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n9752) );
  AOI22_X1 U10841 ( .A1(n9757), .A2(n9753), .B1(n9752), .B2(n9754), .ZN(
        P1_U3525) );
  INV_X1 U10842 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n9755) );
  AOI22_X1 U10843 ( .A1(n9757), .A2(n9756), .B1(n9755), .B2(n9754), .ZN(
        P1_U3529) );
  AOI22_X1 U10844 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(n9796), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3151), .ZN(n9762) );
  XOR2_X1 U10845 ( .A(P2_IR_REG_0__SCAN_IN), .B(n9758), .Z(n9759) );
  OAI21_X1 U10846 ( .B1(n9760), .B2(n9807), .A(n9759), .ZN(n9761) );
  OAI211_X1 U10847 ( .C1(n9814), .C2(n9763), .A(n9762), .B(n9761), .ZN(
        P2_U3182) );
  AOI21_X1 U10848 ( .B1(n9765), .B2(n9876), .A(n9764), .ZN(n9769) );
  AOI21_X1 U10849 ( .B1(n9767), .B2(n6104), .A(n9766), .ZN(n9768) );
  OAI22_X1 U10850 ( .A1(n9769), .A2(n9803), .B1(n9810), .B2(n9768), .ZN(n9770)
         );
  AOI211_X1 U10851 ( .C1(n9773), .C2(n9772), .A(n9771), .B(n9770), .ZN(n9779)
         );
  OAI21_X1 U10852 ( .B1(n9776), .B2(n9775), .A(n9774), .ZN(n9777) );
  AOI22_X1 U10853 ( .A1(n9777), .A2(n9807), .B1(n9796), .B2(
        P2_ADDR_REG_3__SCAN_IN), .ZN(n9778) );
  NAND2_X1 U10854 ( .A1(n9779), .A2(n9778), .ZN(P2_U3185) );
  OAI211_X1 U10855 ( .C1(n9782), .C2(n9781), .A(n9780), .B(n9807), .ZN(n9783)
         );
  INV_X1 U10856 ( .A(n9783), .ZN(n9792) );
  AOI21_X1 U10857 ( .B1(n9786), .B2(n9785), .A(n9784), .ZN(n9790) );
  AOI21_X1 U10858 ( .B1(n9879), .B2(n9788), .A(n9787), .ZN(n9789) );
  OAI22_X1 U10859 ( .A1(n9790), .A2(n9810), .B1(n9789), .B2(n9803), .ZN(n9791)
         );
  AOI211_X1 U10860 ( .C1(P2_ADDR_REG_5__SCAN_IN), .C2(n9796), .A(n9792), .B(
        n9791), .ZN(n9794) );
  OAI211_X1 U10861 ( .C1(n9814), .C2(n9795), .A(n9794), .B(n9793), .ZN(
        P2_U3187) );
  AOI22_X1 U10862 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(n9796), .B1(
        P2_REG3_REG_17__SCAN_IN), .B2(P2_U3151), .ZN(n9812) );
  AOI21_X1 U10863 ( .B1(n9799), .B2(n9798), .A(n9797), .ZN(n9811) );
  OAI21_X1 U10864 ( .B1(n9806), .B2(n9805), .A(n9804), .ZN(n9808) );
  INV_X1 U10865 ( .A(n9815), .ZN(n9818) );
  OAI21_X1 U10866 ( .B1(n9818), .B2(n9817), .A(n9816), .ZN(n9823) );
  AOI222_X1 U10867 ( .A1(n9824), .A2(n9823), .B1(n9822), .B2(n9821), .C1(n9820), .C2(n9819), .ZN(n9825) );
  OAI21_X1 U10868 ( .B1(n9824), .B2(n9826), .A(n9825), .ZN(P2_U3226) );
  OAI22_X1 U10869 ( .A1(n9829), .A2(n9828), .B1(n9827), .B2(n9861), .ZN(n9830)
         );
  OR2_X1 U10870 ( .A1(n9831), .A2(n9830), .ZN(n9874) );
  OAI22_X1 U10871 ( .A1(n8939), .A2(P2_REG0_REG_2__SCAN_IN), .B1(n9874), .B2(
        n9873), .ZN(n9832) );
  INV_X1 U10872 ( .A(n9832), .ZN(P2_U3396) );
  INV_X1 U10873 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n9838) );
  NAND2_X1 U10874 ( .A1(n9833), .A2(n9853), .ZN(n9837) );
  NAND2_X1 U10875 ( .A1(n9834), .A2(n9871), .ZN(n9835) );
  AND3_X1 U10876 ( .A1(n9837), .A2(n9836), .A3(n9835), .ZN(n9877) );
  AOI22_X1 U10877 ( .A1(n9873), .A2(n9838), .B1(n9877), .B2(n8939), .ZN(
        P2_U3399) );
  INV_X1 U10878 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n9844) );
  INV_X1 U10879 ( .A(n9839), .ZN(n9843) );
  OAI21_X1 U10880 ( .B1(n9841), .B2(n9861), .A(n9840), .ZN(n9842) );
  AOI21_X1 U10881 ( .B1(n9843), .B2(n9853), .A(n9842), .ZN(n9878) );
  AOI22_X1 U10882 ( .A1(n9873), .A2(n9844), .B1(n9878), .B2(n8939), .ZN(
        P2_U3402) );
  INV_X1 U10883 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n9849) );
  AOI22_X1 U10884 ( .A1(n9846), .A2(n9853), .B1(n9871), .B2(n9845), .ZN(n9847)
         );
  AND2_X1 U10885 ( .A1(n9848), .A2(n9847), .ZN(n9880) );
  AOI22_X1 U10886 ( .A1(n9873), .A2(n9849), .B1(n9880), .B2(n8939), .ZN(
        P2_U3405) );
  INV_X1 U10887 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n9855) );
  NOR2_X1 U10888 ( .A1(n9850), .A2(n9861), .ZN(n9852) );
  AOI211_X1 U10889 ( .C1(n9854), .C2(n9853), .A(n9852), .B(n9851), .ZN(n9881)
         );
  AOI22_X1 U10890 ( .A1(n9873), .A2(n9855), .B1(n9881), .B2(n8939), .ZN(
        P2_U3408) );
  INV_X1 U10891 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n9860) );
  NOR2_X1 U10892 ( .A1(n9856), .A2(n9866), .ZN(n9858) );
  AOI211_X1 U10893 ( .C1(n9871), .C2(n9859), .A(n9858), .B(n9857), .ZN(n9882)
         );
  AOI22_X1 U10894 ( .A1(n9873), .A2(n9860), .B1(n9882), .B2(n8939), .ZN(
        P2_U3414) );
  INV_X1 U10895 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n9865) );
  OAI22_X1 U10896 ( .A1(n9862), .A2(n9866), .B1(n4676), .B2(n9861), .ZN(n9863)
         );
  NOR2_X1 U10897 ( .A1(n9864), .A2(n9863), .ZN(n9884) );
  AOI22_X1 U10898 ( .A1(n9873), .A2(n9865), .B1(n9884), .B2(n8939), .ZN(
        P2_U3423) );
  INV_X1 U10899 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n9872) );
  NOR2_X1 U10900 ( .A1(n9867), .A2(n9866), .ZN(n9869) );
  AOI211_X1 U10901 ( .C1(n9871), .C2(n9870), .A(n9869), .B(n9868), .ZN(n9886)
         );
  AOI22_X1 U10902 ( .A1(n9873), .A2(n9872), .B1(n9886), .B2(n8939), .ZN(
        P2_U3426) );
  OAI22_X1 U10903 ( .A1(n9885), .A2(n9874), .B1(P2_REG1_REG_2__SCAN_IN), .B2(
        n9887), .ZN(n9875) );
  INV_X1 U10904 ( .A(n9875), .ZN(P2_U3461) );
  AOI22_X1 U10905 ( .A1(n9887), .A2(n9877), .B1(n9876), .B2(n9885), .ZN(
        P2_U3462) );
  AOI22_X1 U10906 ( .A1(n9887), .A2(n9878), .B1(n5972), .B2(n9885), .ZN(
        P2_U3463) );
  AOI22_X1 U10907 ( .A1(n9887), .A2(n9880), .B1(n9879), .B2(n9885), .ZN(
        P2_U3464) );
  AOI22_X1 U10908 ( .A1(n9887), .A2(n9881), .B1(n6142), .B2(n9885), .ZN(
        P2_U3465) );
  AOI22_X1 U10909 ( .A1(n9887), .A2(n9882), .B1(n6158), .B2(n9885), .ZN(
        P2_U3467) );
  AOI22_X1 U10910 ( .A1(n9887), .A2(n9884), .B1(n9883), .B2(n9885), .ZN(
        P2_U3470) );
  AOI22_X1 U10911 ( .A1(n9887), .A2(n9886), .B1(n6200), .B2(n9885), .ZN(
        P2_U3471) );
  NAND3_X1 U10912 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .A3(P2_ADDR_REG_0__SCAN_IN), .ZN(n9890) );
  AND2_X1 U10913 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n9888) );
  NOR2_X1 U10914 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n9888), .ZN(n9889) );
  INV_X1 U10915 ( .A(n9889), .ZN(n9907) );
  NAND2_X1 U10916 ( .A1(n9891), .A2(n9890), .ZN(n9906) );
  OAI222_X1 U10917 ( .A1(n9891), .A2(n9890), .B1(n9891), .B2(n9907), .C1(n9889), .C2(n9906), .ZN(ADD_1068_U5) );
  XOR2_X1 U10918 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  NOR2_X1 U10919 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n9892) );
  AOI21_X1 U10920 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n9892), .ZN(n9915) );
  AOI22_X1 U10921 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .B1(n9894), .B2(n9893), .ZN(n9918) );
  NOR2_X1 U10922 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n9895) );
  AOI21_X1 U10923 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n9895), .ZN(n9921) );
  NOR2_X1 U10924 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n9896) );
  AOI21_X1 U10925 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n9896), .ZN(n9924) );
  NOR2_X1 U10926 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n9897) );
  AOI21_X1 U10927 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n9897), .ZN(n9927) );
  NOR2_X1 U10928 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n9898) );
  AOI21_X1 U10929 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n9898), .ZN(n9930) );
  NOR2_X1 U10930 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n9899) );
  AOI21_X1 U10931 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n9899), .ZN(n9933) );
  NOR2_X1 U10932 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n9900) );
  AOI21_X1 U10933 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n9900), .ZN(n9936) );
  NOR2_X1 U10934 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n9901) );
  AOI21_X1 U10935 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(P2_ADDR_REG_9__SCAN_IN), 
        .A(n9901), .ZN(n10144) );
  NOR2_X1 U10936 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n9902) );
  AOI21_X1 U10937 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(P2_ADDR_REG_8__SCAN_IN), 
        .A(n9902), .ZN(n10147) );
  NOR2_X1 U10938 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n9903) );
  AOI21_X1 U10939 ( .B1(P1_ADDR_REG_7__SCAN_IN), .B2(P2_ADDR_REG_7__SCAN_IN), 
        .A(n9903), .ZN(n10150) );
  NOR2_X1 U10940 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n9904) );
  AOI21_X1 U10941 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(P2_ADDR_REG_6__SCAN_IN), 
        .A(n9904), .ZN(n10153) );
  NOR2_X1 U10942 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(P2_ADDR_REG_5__SCAN_IN), 
        .ZN(n9905) );
  AOI21_X1 U10943 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(P1_ADDR_REG_5__SCAN_IN), 
        .A(n9905), .ZN(n10156) );
  NAND2_X1 U10944 ( .A1(n9907), .A2(n9906), .ZN(n10141) );
  NAND2_X1 U10945 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n9908) );
  OAI21_X1 U10946 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(P2_ADDR_REG_2__SCAN_IN), 
        .A(n9908), .ZN(n10140) );
  NOR2_X1 U10947 ( .A1(n10141), .A2(n10140), .ZN(n10139) );
  AOI21_X1 U10948 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(P1_ADDR_REG_2__SCAN_IN), 
        .A(n10139), .ZN(n10159) );
  NAND2_X1 U10949 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n9909) );
  OAI21_X1 U10950 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n9909), .ZN(n10158) );
  NOR2_X1 U10951 ( .A1(n10159), .A2(n10158), .ZN(n10157) );
  AOI21_X1 U10952 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(P1_ADDR_REG_3__SCAN_IN), 
        .A(n10157), .ZN(n10162) );
  NOR2_X1 U10953 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n9910) );
  AOI21_X1 U10954 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(P1_ADDR_REG_4__SCAN_IN), 
        .A(n9910), .ZN(n10161) );
  NAND2_X1 U10955 ( .A1(n10162), .A2(n10161), .ZN(n10160) );
  OAI21_X1 U10956 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(P2_ADDR_REG_4__SCAN_IN), 
        .A(n10160), .ZN(n10155) );
  NAND2_X1 U10957 ( .A1(n10156), .A2(n10155), .ZN(n10154) );
  OAI21_X1 U10958 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(P2_ADDR_REG_5__SCAN_IN), 
        .A(n10154), .ZN(n10152) );
  NAND2_X1 U10959 ( .A1(n10153), .A2(n10152), .ZN(n10151) );
  OAI21_X1 U10960 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(P1_ADDR_REG_6__SCAN_IN), 
        .A(n10151), .ZN(n10149) );
  NAND2_X1 U10961 ( .A1(n10150), .A2(n10149), .ZN(n10148) );
  OAI21_X1 U10962 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(P1_ADDR_REG_7__SCAN_IN), 
        .A(n10148), .ZN(n10146) );
  NAND2_X1 U10963 ( .A1(n10147), .A2(n10146), .ZN(n10145) );
  OAI21_X1 U10964 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(P1_ADDR_REG_8__SCAN_IN), 
        .A(n10145), .ZN(n10143) );
  NAND2_X1 U10965 ( .A1(n10144), .A2(n10143), .ZN(n10142) );
  OAI21_X1 U10966 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(P1_ADDR_REG_9__SCAN_IN), 
        .A(n10142), .ZN(n9935) );
  NAND2_X1 U10967 ( .A1(n9936), .A2(n9935), .ZN(n9934) );
  OAI21_X1 U10968 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n9934), .ZN(n9932) );
  NAND2_X1 U10969 ( .A1(n9933), .A2(n9932), .ZN(n9931) );
  OAI21_X1 U10970 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n9931), .ZN(n9929) );
  NAND2_X1 U10971 ( .A1(n9930), .A2(n9929), .ZN(n9928) );
  OAI21_X1 U10972 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n9928), .ZN(n9926) );
  NAND2_X1 U10973 ( .A1(n9927), .A2(n9926), .ZN(n9925) );
  OAI21_X1 U10974 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n9925), .ZN(n9923) );
  NAND2_X1 U10975 ( .A1(n9924), .A2(n9923), .ZN(n9922) );
  OAI21_X1 U10976 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n9922), .ZN(n9920) );
  NAND2_X1 U10977 ( .A1(n9921), .A2(n9920), .ZN(n9919) );
  OAI21_X1 U10978 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n9919), .ZN(n9917) );
  NAND2_X1 U10979 ( .A1(n9918), .A2(n9917), .ZN(n9916) );
  OAI21_X1 U10980 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n9916), .ZN(n9914) );
  NAND2_X1 U10981 ( .A1(n9915), .A2(n9914), .ZN(n9913) );
  OAI21_X1 U10982 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n9913), .ZN(n9937) );
  NAND2_X1 U10983 ( .A1(n9938), .A2(n9937), .ZN(n9939) );
  OAI21_X1 U10984 ( .B1(n9937), .B2(n9938), .A(n9939), .ZN(n9912) );
  XOR2_X1 U10985 ( .A(n9912), .B(n9911), .Z(ADD_1068_U55) );
  OAI21_X1 U10986 ( .B1(n9915), .B2(n9914), .A(n9913), .ZN(ADD_1068_U56) );
  OAI21_X1 U10987 ( .B1(n9918), .B2(n9917), .A(n9916), .ZN(ADD_1068_U57) );
  OAI21_X1 U10988 ( .B1(n9921), .B2(n9920), .A(n9919), .ZN(ADD_1068_U58) );
  OAI21_X1 U10989 ( .B1(n9924), .B2(n9923), .A(n9922), .ZN(ADD_1068_U59) );
  OAI21_X1 U10990 ( .B1(n9927), .B2(n9926), .A(n9925), .ZN(ADD_1068_U60) );
  OAI21_X1 U10991 ( .B1(n9930), .B2(n9929), .A(n9928), .ZN(ADD_1068_U61) );
  OAI21_X1 U10992 ( .B1(n9933), .B2(n9932), .A(n9931), .ZN(ADD_1068_U62) );
  OAI21_X1 U10993 ( .B1(n9936), .B2(n9935), .A(n9934), .ZN(ADD_1068_U63) );
  NOR2_X1 U10994 ( .A1(n9938), .A2(n9937), .ZN(n9940) );
  OAI21_X1 U10995 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n9940), .A(n9939), .ZN(
        n10138) );
  AOI22_X1 U10996 ( .A1(SI_3_), .A2(keyinput_g29), .B1(P2_REG3_REG_28__SCAN_IN), .B2(keyinput_g42), .ZN(n9941) );
  OAI221_X1 U10997 ( .B1(SI_3_), .B2(keyinput_g29), .C1(
        P2_REG3_REG_28__SCAN_IN), .C2(keyinput_g42), .A(n9941), .ZN(n9948) );
  AOI22_X1 U10998 ( .A1(SI_17_), .A2(keyinput_g15), .B1(SI_24_), .B2(
        keyinput_g8), .ZN(n9942) );
  OAI221_X1 U10999 ( .B1(SI_17_), .B2(keyinput_g15), .C1(SI_24_), .C2(
        keyinput_g8), .A(n9942), .ZN(n9947) );
  AOI22_X1 U11000 ( .A1(SI_19_), .A2(keyinput_g13), .B1(SI_22_), .B2(
        keyinput_g10), .ZN(n9943) );
  OAI221_X1 U11001 ( .B1(SI_19_), .B2(keyinput_g13), .C1(SI_22_), .C2(
        keyinput_g10), .A(n9943), .ZN(n9946) );
  AOI22_X1 U11002 ( .A1(SI_29_), .A2(keyinput_g3), .B1(P2_REG3_REG_15__SCAN_IN), .B2(keyinput_g63), .ZN(n9944) );
  OAI221_X1 U11003 ( .B1(SI_29_), .B2(keyinput_g3), .C1(
        P2_REG3_REG_15__SCAN_IN), .C2(keyinput_g63), .A(n9944), .ZN(n9945) );
  NOR4_X1 U11004 ( .A1(n9948), .A2(n9947), .A3(n9946), .A4(n9945), .ZN(n9976)
         );
  XOR2_X1 U11005 ( .A(SI_31_), .B(keyinput_g1), .Z(n9955) );
  AOI22_X1 U11006 ( .A1(SI_16_), .A2(keyinput_g16), .B1(
        P2_REG3_REG_19__SCAN_IN), .B2(keyinput_g41), .ZN(n9949) );
  OAI221_X1 U11007 ( .B1(SI_16_), .B2(keyinput_g16), .C1(
        P2_REG3_REG_19__SCAN_IN), .C2(keyinput_g41), .A(n9949), .ZN(n9954) );
  AOI22_X1 U11008 ( .A1(SI_14_), .A2(keyinput_g18), .B1(P2_REG3_REG_9__SCAN_IN), .B2(keyinput_g53), .ZN(n9950) );
  OAI221_X1 U11009 ( .B1(SI_14_), .B2(keyinput_g18), .C1(
        P2_REG3_REG_9__SCAN_IN), .C2(keyinput_g53), .A(n9950), .ZN(n9953) );
  AOI22_X1 U11010 ( .A1(P2_REG3_REG_2__SCAN_IN), .A2(keyinput_g59), .B1(SI_0_), 
        .B2(keyinput_g32), .ZN(n9951) );
  OAI221_X1 U11011 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(keyinput_g59), .C1(SI_0_), .C2(keyinput_g32), .A(n9951), .ZN(n9952) );
  NOR4_X1 U11012 ( .A1(n9955), .A2(n9954), .A3(n9953), .A4(n9952), .ZN(n9975)
         );
  AOI22_X1 U11013 ( .A1(SI_2_), .A2(keyinput_g30), .B1(SI_15_), .B2(
        keyinput_g17), .ZN(n9956) );
  OAI221_X1 U11014 ( .B1(SI_2_), .B2(keyinput_g30), .C1(SI_15_), .C2(
        keyinput_g17), .A(n9956), .ZN(n9964) );
  AOI22_X1 U11015 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(keyinput_g37), .B1(
        P2_REG3_REG_27__SCAN_IN), .B2(keyinput_g36), .ZN(n9957) );
  OAI221_X1 U11016 ( .B1(P2_REG3_REG_14__SCAN_IN), .B2(keyinput_g37), .C1(
        P2_REG3_REG_27__SCAN_IN), .C2(keyinput_g36), .A(n9957), .ZN(n9963) );
  AOI22_X1 U11017 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(keyinput_g60), .B1(n9959), .B2(keyinput_g5), .ZN(n9958) );
  OAI221_X1 U11018 ( .B1(P2_REG3_REG_18__SCAN_IN), .B2(keyinput_g60), .C1(
        n9959), .C2(keyinput_g5), .A(n9958), .ZN(n9962) );
  AOI22_X1 U11019 ( .A1(SI_6_), .A2(keyinput_g26), .B1(P2_REG3_REG_12__SCAN_IN), .B2(keyinput_g46), .ZN(n9960) );
  OAI221_X1 U11020 ( .B1(SI_6_), .B2(keyinput_g26), .C1(
        P2_REG3_REG_12__SCAN_IN), .C2(keyinput_g46), .A(n9960), .ZN(n9961) );
  NOR4_X1 U11021 ( .A1(n9964), .A2(n9963), .A3(n9962), .A4(n9961), .ZN(n9974)
         );
  AOI22_X1 U11022 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(keyinput_g48), .B1(
        P2_REG3_REG_26__SCAN_IN), .B2(keyinput_g62), .ZN(n9965) );
  OAI221_X1 U11023 ( .B1(P2_REG3_REG_16__SCAN_IN), .B2(keyinput_g48), .C1(
        P2_REG3_REG_26__SCAN_IN), .C2(keyinput_g62), .A(n9965), .ZN(n9972) );
  AOI22_X1 U11024 ( .A1(P2_WR_REG_SCAN_IN), .A2(keyinput_g0), .B1(SI_7_), .B2(
        keyinput_g25), .ZN(n9966) );
  OAI221_X1 U11025 ( .B1(P2_WR_REG_SCAN_IN), .B2(keyinput_g0), .C1(SI_7_), 
        .C2(keyinput_g25), .A(n9966), .ZN(n9971) );
  AOI22_X1 U11026 ( .A1(SI_30_), .A2(keyinput_g2), .B1(P2_REG3_REG_10__SCAN_IN), .B2(keyinput_g39), .ZN(n9967) );
  OAI221_X1 U11027 ( .B1(SI_30_), .B2(keyinput_g2), .C1(
        P2_REG3_REG_10__SCAN_IN), .C2(keyinput_g39), .A(n9967), .ZN(n9970) );
  AOI22_X1 U11028 ( .A1(SI_23_), .A2(keyinput_g9), .B1(SI_26_), .B2(
        keyinput_g6), .ZN(n9968) );
  OAI221_X1 U11029 ( .B1(SI_23_), .B2(keyinput_g9), .C1(SI_26_), .C2(
        keyinput_g6), .A(n9968), .ZN(n9969) );
  NOR4_X1 U11030 ( .A1(n9972), .A2(n9971), .A3(n9970), .A4(n9969), .ZN(n9973)
         );
  NAND4_X1 U11031 ( .A1(n9976), .A2(n9975), .A3(n9974), .A4(n9973), .ZN(n10134) );
  INV_X1 U11032 ( .A(SI_10_), .ZN(n10105) );
  AOI22_X1 U11033 ( .A1(n10096), .A2(keyinput_g33), .B1(keyinput_g22), .B2(
        n10105), .ZN(n9977) );
  OAI221_X1 U11034 ( .B1(n10096), .B2(keyinput_g33), .C1(n10105), .C2(
        keyinput_g22), .A(n9977), .ZN(n9986) );
  INV_X1 U11035 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n10051) );
  AOI22_X1 U11036 ( .A1(n10051), .A2(keyinput_g35), .B1(P2_U3151), .B2(
        keyinput_g34), .ZN(n9978) );
  OAI221_X1 U11037 ( .B1(n10051), .B2(keyinput_g35), .C1(P2_U3151), .C2(
        keyinput_g34), .A(n9978), .ZN(n9985) );
  INV_X1 U11038 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n9980) );
  AOI22_X1 U11039 ( .A1(n9980), .A2(keyinput_g38), .B1(keyinput_g19), .B2(
        n10110), .ZN(n9979) );
  OAI221_X1 U11040 ( .B1(n9980), .B2(keyinput_g38), .C1(n10110), .C2(
        keyinput_g19), .A(n9979), .ZN(n9984) );
  XNOR2_X1 U11041 ( .A(P2_REG3_REG_17__SCAN_IN), .B(keyinput_g50), .ZN(n9982)
         );
  XNOR2_X1 U11042 ( .A(SI_4_), .B(keyinput_g28), .ZN(n9981) );
  NAND2_X1 U11043 ( .A1(n9982), .A2(n9981), .ZN(n9983) );
  NOR4_X1 U11044 ( .A1(n9986), .A2(n9985), .A3(n9984), .A4(n9983), .ZN(n10024)
         );
  AOI22_X1 U11045 ( .A1(n10064), .A2(keyinput_g55), .B1(keyinput_g56), .B2(
        n6208), .ZN(n9987) );
  OAI221_X1 U11046 ( .B1(n10064), .B2(keyinput_g55), .C1(n6208), .C2(
        keyinput_g56), .A(n9987), .ZN(n9997) );
  AOI22_X1 U11047 ( .A1(n10070), .A2(keyinput_g58), .B1(keyinput_g20), .B2(
        n9989), .ZN(n9988) );
  OAI221_X1 U11048 ( .B1(n10070), .B2(keyinput_g58), .C1(n9989), .C2(
        keyinput_g20), .A(n9988), .ZN(n9996) );
  AOI22_X1 U11049 ( .A1(n9991), .A2(keyinput_g23), .B1(n10048), .B2(
        keyinput_g51), .ZN(n9990) );
  OAI221_X1 U11050 ( .B1(n9991), .B2(keyinput_g23), .C1(n10048), .C2(
        keyinput_g51), .A(n9990), .ZN(n9995) );
  XNOR2_X1 U11051 ( .A(P2_REG3_REG_4__SCAN_IN), .B(keyinput_g52), .ZN(n9993)
         );
  XNOR2_X1 U11052 ( .A(SI_5_), .B(keyinput_g27), .ZN(n9992) );
  NAND2_X1 U11053 ( .A1(n9993), .A2(n9992), .ZN(n9994) );
  NOR4_X1 U11054 ( .A1(n9997), .A2(n9996), .A3(n9995), .A4(n9994), .ZN(n10023)
         );
  INV_X1 U11055 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n10047) );
  AOI22_X1 U11056 ( .A1(n10047), .A2(keyinput_g61), .B1(keyinput_g4), .B2(
        n10062), .ZN(n9998) );
  OAI221_X1 U11057 ( .B1(n10047), .B2(keyinput_g61), .C1(n10062), .C2(
        keyinput_g4), .A(n9998), .ZN(n10007) );
  AOI22_X1 U11058 ( .A1(n6123), .A2(keyinput_g49), .B1(n10000), .B2(
        keyinput_g45), .ZN(n9999) );
  OAI221_X1 U11059 ( .B1(n6123), .B2(keyinput_g49), .C1(n10000), .C2(
        keyinput_g45), .A(n9999), .ZN(n10006) );
  INV_X1 U11060 ( .A(SI_18_), .ZN(n10041) );
  AOI22_X1 U11061 ( .A1(n10098), .A2(keyinput_g43), .B1(keyinput_g14), .B2(
        n10041), .ZN(n10001) );
  OAI221_X1 U11062 ( .B1(n10098), .B2(keyinput_g43), .C1(n10041), .C2(
        keyinput_g14), .A(n10001), .ZN(n10005) );
  XNOR2_X1 U11063 ( .A(P2_REG3_REG_22__SCAN_IN), .B(keyinput_g57), .ZN(n10003)
         );
  XNOR2_X1 U11064 ( .A(SI_1_), .B(keyinput_g31), .ZN(n10002) );
  NAND2_X1 U11065 ( .A1(n10003), .A2(n10002), .ZN(n10004) );
  NOR4_X1 U11066 ( .A1(n10007), .A2(n10006), .A3(n10005), .A4(n10004), .ZN(
        n10022) );
  INV_X1 U11067 ( .A(SI_25_), .ZN(n10009) );
  AOI22_X1 U11068 ( .A1(n6470), .A2(keyinput_g44), .B1(n10009), .B2(
        keyinput_g7), .ZN(n10008) );
  OAI221_X1 U11069 ( .B1(n6470), .B2(keyinput_g44), .C1(n10009), .C2(
        keyinput_g7), .A(n10008), .ZN(n10020) );
  INV_X1 U11070 ( .A(SI_21_), .ZN(n10012) );
  AOI22_X1 U11071 ( .A1(n10012), .A2(keyinput_g11), .B1(n10011), .B2(
        keyinput_g40), .ZN(n10010) );
  OAI221_X1 U11072 ( .B1(n10012), .B2(keyinput_g11), .C1(n10011), .C2(
        keyinput_g40), .A(n10010), .ZN(n10019) );
  AOI22_X1 U11073 ( .A1(n5536), .A2(keyinput_g12), .B1(keyinput_g21), .B2(
        n10014), .ZN(n10013) );
  OAI221_X1 U11074 ( .B1(n5536), .B2(keyinput_g12), .C1(n10014), .C2(
        keyinput_g21), .A(n10013), .ZN(n10018) );
  AOI22_X1 U11075 ( .A1(n10016), .A2(keyinput_g47), .B1(keyinput_g54), .B2(
        n10111), .ZN(n10015) );
  OAI221_X1 U11076 ( .B1(n10016), .B2(keyinput_g47), .C1(n10111), .C2(
        keyinput_g54), .A(n10015), .ZN(n10017) );
  NOR4_X1 U11077 ( .A1(n10020), .A2(n10019), .A3(n10018), .A4(n10017), .ZN(
        n10021) );
  NAND4_X1 U11078 ( .A1(n10024), .A2(n10023), .A3(n10022), .A4(n10021), .ZN(
        n10133) );
  INV_X1 U11079 ( .A(keyinput_f24), .ZN(n10126) );
  OAI22_X1 U11080 ( .A1(P2_REG3_REG_2__SCAN_IN), .A2(keyinput_f59), .B1(
        keyinput_f1), .B2(SI_31_), .ZN(n10025) );
  AOI221_X1 U11081 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(keyinput_f59), .C1(
        SI_31_), .C2(keyinput_f1), .A(n10025), .ZN(n10032) );
  OAI22_X1 U11082 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(keyinput_f60), .B1(SI_2_), .B2(keyinput_f30), .ZN(n10026) );
  AOI221_X1 U11083 ( .B1(P2_REG3_REG_18__SCAN_IN), .B2(keyinput_f60), .C1(
        keyinput_f30), .C2(SI_2_), .A(n10026), .ZN(n10031) );
  OAI22_X1 U11084 ( .A1(SI_21_), .A2(keyinput_f11), .B1(keyinput_f12), .B2(
        SI_20_), .ZN(n10027) );
  AOI221_X1 U11085 ( .B1(SI_21_), .B2(keyinput_f11), .C1(SI_20_), .C2(
        keyinput_f12), .A(n10027), .ZN(n10030) );
  OAI22_X1 U11086 ( .A1(SI_12_), .A2(keyinput_f20), .B1(SI_6_), .B2(
        keyinput_f26), .ZN(n10028) );
  AOI221_X1 U11087 ( .B1(SI_12_), .B2(keyinput_f20), .C1(keyinput_f26), .C2(
        SI_6_), .A(n10028), .ZN(n10029) );
  NAND4_X1 U11088 ( .A1(n10032), .A2(n10031), .A3(n10030), .A4(n10029), .ZN(
        n10125) );
  OAI22_X1 U11089 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(keyinput_f40), .B1(SI_7_), 
        .B2(keyinput_f25), .ZN(n10033) );
  AOI221_X1 U11090 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(keyinput_f40), .C1(
        keyinput_f25), .C2(SI_7_), .A(n10033), .ZN(n10039) );
  OAI22_X1 U11091 ( .A1(SI_27_), .A2(keyinput_f5), .B1(keyinput_f7), .B2(
        SI_25_), .ZN(n10034) );
  AOI221_X1 U11092 ( .B1(SI_27_), .B2(keyinput_f5), .C1(SI_25_), .C2(
        keyinput_f7), .A(n10034), .ZN(n10038) );
  OAI22_X1 U11093 ( .A1(P2_REG3_REG_21__SCAN_IN), .A2(keyinput_f45), .B1(
        keyinput_f32), .B2(SI_0_), .ZN(n10035) );
  AOI221_X1 U11094 ( .B1(P2_REG3_REG_21__SCAN_IN), .B2(keyinput_f45), .C1(
        SI_0_), .C2(keyinput_f32), .A(n10035), .ZN(n10037) );
  XNOR2_X1 U11095 ( .A(SI_29_), .B(keyinput_f3), .ZN(n10036) );
  NAND4_X1 U11096 ( .A1(n10039), .A2(n10038), .A3(n10037), .A4(n10036), .ZN(
        n10124) );
  XOR2_X1 U11097 ( .A(keyinput_f0), .B(P2_WR_REG_SCAN_IN), .Z(n10043) );
  AOI22_X1 U11098 ( .A1(n10041), .A2(keyinput_f14), .B1(n6208), .B2(
        keyinput_f56), .ZN(n10040) );
  OAI221_X1 U11099 ( .B1(n10041), .B2(keyinput_f14), .C1(n6208), .C2(
        keyinput_f56), .A(n10040), .ZN(n10042) );
  AOI211_X1 U11100 ( .C1(n10045), .C2(keyinput_f15), .A(n10043), .B(n10042), 
        .ZN(n10044) );
  OAI21_X1 U11101 ( .B1(n10045), .B2(keyinput_f15), .A(n10044), .ZN(n10059) );
  OAI22_X1 U11102 ( .A1(n10048), .A2(keyinput_f51), .B1(n10047), .B2(
        keyinput_f61), .ZN(n10046) );
  AOI221_X1 U11103 ( .B1(n10048), .B2(keyinput_f51), .C1(keyinput_f61), .C2(
        n10047), .A(n10046), .ZN(n10049) );
  INV_X1 U11104 ( .A(n10049), .ZN(n10058) );
  AOI22_X1 U11105 ( .A1(n6470), .A2(keyinput_f44), .B1(n10051), .B2(
        keyinput_f35), .ZN(n10050) );
  OAI221_X1 U11106 ( .B1(n6470), .B2(keyinput_f44), .C1(n10051), .C2(
        keyinput_f35), .A(n10050), .ZN(n10057) );
  XNOR2_X1 U11107 ( .A(SI_4_), .B(keyinput_f28), .ZN(n10055) );
  XNOR2_X1 U11108 ( .A(SI_5_), .B(keyinput_f27), .ZN(n10054) );
  XNOR2_X1 U11109 ( .A(P2_REG3_REG_15__SCAN_IN), .B(keyinput_f63), .ZN(n10053)
         );
  XNOR2_X1 U11110 ( .A(P2_REG3_REG_16__SCAN_IN), .B(keyinput_f48), .ZN(n10052)
         );
  NAND4_X1 U11111 ( .A1(n10055), .A2(n10054), .A3(n10053), .A4(n10052), .ZN(
        n10056) );
  NOR4_X1 U11112 ( .A1(n10059), .A2(n10058), .A3(n10057), .A4(n10056), .ZN(
        n10068) );
  INV_X1 U11113 ( .A(SI_22_), .ZN(n10061) );
  OAI22_X1 U11114 ( .A1(n10062), .A2(keyinput_f4), .B1(n10061), .B2(
        keyinput_f10), .ZN(n10060) );
  AOI221_X1 U11115 ( .B1(n10062), .B2(keyinput_f4), .C1(keyinput_f10), .C2(
        n10061), .A(n10060), .ZN(n10067) );
  INV_X1 U11116 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n10065) );
  OAI22_X1 U11117 ( .A1(n10065), .A2(keyinput_f57), .B1(n10064), .B2(
        keyinput_f55), .ZN(n10063) );
  AOI221_X1 U11118 ( .B1(n10065), .B2(keyinput_f57), .C1(keyinput_f55), .C2(
        n10064), .A(n10063), .ZN(n10066) );
  NAND3_X1 U11119 ( .A1(n10068), .A2(n10067), .A3(n10066), .ZN(n10123) );
  AOI22_X1 U11120 ( .A1(n10071), .A2(keyinput_f6), .B1(n10070), .B2(
        keyinput_f58), .ZN(n10069) );
  OAI221_X1 U11121 ( .B1(n10071), .B2(keyinput_f6), .C1(n10070), .C2(
        keyinput_f58), .A(n10069), .ZN(n10080) );
  AOI22_X1 U11122 ( .A1(SI_9_), .A2(keyinput_f23), .B1(P2_REG3_REG_4__SCAN_IN), 
        .B2(keyinput_f52), .ZN(n10072) );
  OAI221_X1 U11123 ( .B1(SI_9_), .B2(keyinput_f23), .C1(P2_REG3_REG_4__SCAN_IN), .C2(keyinput_f52), .A(n10072), .ZN(n10079) );
  AOI22_X1 U11124 ( .A1(SI_11_), .A2(keyinput_f21), .B1(SI_16_), .B2(
        keyinput_f16), .ZN(n10073) );
  OAI221_X1 U11125 ( .B1(SI_11_), .B2(keyinput_f21), .C1(SI_16_), .C2(
        keyinput_f16), .A(n10073), .ZN(n10078) );
  XNOR2_X1 U11126 ( .A(n10074), .B(keyinput_f8), .ZN(n10076) );
  XNOR2_X1 U11127 ( .A(SI_1_), .B(keyinput_f31), .ZN(n10075) );
  NAND2_X1 U11128 ( .A1(n10076), .A2(n10075), .ZN(n10077) );
  NOR4_X1 U11129 ( .A1(n10080), .A2(n10079), .A3(n10078), .A4(n10077), .ZN(
        n10121) );
  AOI22_X1 U11130 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(keyinput_f46), .B1(
        P2_REG3_REG_14__SCAN_IN), .B2(keyinput_f37), .ZN(n10081) );
  OAI221_X1 U11131 ( .B1(P2_REG3_REG_12__SCAN_IN), .B2(keyinput_f46), .C1(
        P2_REG3_REG_14__SCAN_IN), .C2(keyinput_f37), .A(n10081), .ZN(n10088)
         );
  AOI22_X1 U11132 ( .A1(SI_30_), .A2(keyinput_f2), .B1(P2_REG3_REG_23__SCAN_IN), .B2(keyinput_f38), .ZN(n10082) );
  OAI221_X1 U11133 ( .B1(SI_30_), .B2(keyinput_f2), .C1(
        P2_REG3_REG_23__SCAN_IN), .C2(keyinput_f38), .A(n10082), .ZN(n10087)
         );
  AOI22_X1 U11134 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(keyinput_f53), .B1(
        P2_STATE_REG_SCAN_IN), .B2(keyinput_f34), .ZN(n10083) );
  OAI221_X1 U11135 ( .B1(P2_REG3_REG_9__SCAN_IN), .B2(keyinput_f53), .C1(
        P2_STATE_REG_SCAN_IN), .C2(keyinput_f34), .A(n10083), .ZN(n10086) );
  AOI22_X1 U11136 ( .A1(SI_14_), .A2(keyinput_f18), .B1(
        P2_REG3_REG_28__SCAN_IN), .B2(keyinput_f42), .ZN(n10084) );
  OAI221_X1 U11137 ( .B1(SI_14_), .B2(keyinput_f18), .C1(
        P2_REG3_REG_28__SCAN_IN), .C2(keyinput_f42), .A(n10084), .ZN(n10085)
         );
  NOR4_X1 U11138 ( .A1(n10088), .A2(n10087), .A3(n10086), .A4(n10085), .ZN(
        n10120) );
  AOI22_X1 U11139 ( .A1(n10091), .A2(keyinput_f50), .B1(n10090), .B2(
        keyinput_f36), .ZN(n10089) );
  OAI221_X1 U11140 ( .B1(n10091), .B2(keyinput_f50), .C1(n10090), .C2(
        keyinput_f36), .A(n10089), .ZN(n10103) );
  AOI22_X1 U11141 ( .A1(n6123), .A2(keyinput_f49), .B1(n10093), .B2(
        keyinput_f39), .ZN(n10092) );
  OAI221_X1 U11142 ( .B1(n6123), .B2(keyinput_f49), .C1(n10093), .C2(
        keyinput_f39), .A(n10092), .ZN(n10102) );
  AOI22_X1 U11143 ( .A1(n10096), .A2(keyinput_f33), .B1(keyinput_f13), .B2(
        n10095), .ZN(n10094) );
  OAI221_X1 U11144 ( .B1(n10096), .B2(keyinput_f33), .C1(n10095), .C2(
        keyinput_f13), .A(n10094), .ZN(n10101) );
  INV_X1 U11145 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n10099) );
  AOI22_X1 U11146 ( .A1(n10099), .A2(keyinput_f41), .B1(keyinput_f43), .B2(
        n10098), .ZN(n10097) );
  OAI221_X1 U11147 ( .B1(n10099), .B2(keyinput_f41), .C1(n10098), .C2(
        keyinput_f43), .A(n10097), .ZN(n10100) );
  NOR4_X1 U11148 ( .A1(n10103), .A2(n10102), .A3(n10101), .A4(n10100), .ZN(
        n10119) );
  INV_X1 U11149 ( .A(SI_23_), .ZN(n10106) );
  AOI22_X1 U11150 ( .A1(n10106), .A2(keyinput_f9), .B1(keyinput_f22), .B2(
        n10105), .ZN(n10104) );
  OAI221_X1 U11151 ( .B1(n10106), .B2(keyinput_f9), .C1(n10105), .C2(
        keyinput_f22), .A(n10104), .ZN(n10117) );
  AOI22_X1 U11152 ( .A1(n5408), .A2(keyinput_f17), .B1(n10108), .B2(
        keyinput_f62), .ZN(n10107) );
  OAI221_X1 U11153 ( .B1(n5408), .B2(keyinput_f17), .C1(n10108), .C2(
        keyinput_f62), .A(n10107), .ZN(n10116) );
  AOI22_X1 U11154 ( .A1(n10111), .A2(keyinput_f54), .B1(n10110), .B2(
        keyinput_f19), .ZN(n10109) );
  OAI221_X1 U11155 ( .B1(n10111), .B2(keyinput_f54), .C1(n10110), .C2(
        keyinput_f19), .A(n10109), .ZN(n10115) );
  XNOR2_X1 U11156 ( .A(P2_REG3_REG_25__SCAN_IN), .B(keyinput_f47), .ZN(n10113)
         );
  XNOR2_X1 U11157 ( .A(SI_3_), .B(keyinput_f29), .ZN(n10112) );
  NAND2_X1 U11158 ( .A1(n10113), .A2(n10112), .ZN(n10114) );
  NOR4_X1 U11159 ( .A1(n10117), .A2(n10116), .A3(n10115), .A4(n10114), .ZN(
        n10118) );
  NAND4_X1 U11160 ( .A1(n10121), .A2(n10120), .A3(n10119), .A4(n10118), .ZN(
        n10122) );
  NOR4_X1 U11161 ( .A1(n10125), .A2(n10124), .A3(n10123), .A4(n10122), .ZN(
        n10129) );
  OAI211_X1 U11162 ( .C1(n10126), .C2(n10129), .A(SI_8_), .B(keyinput_g24), 
        .ZN(n10131) );
  INV_X1 U11163 ( .A(keyinput_g24), .ZN(n10127) );
  OAI211_X1 U11164 ( .C1(n10129), .C2(keyinput_f24), .A(n10128), .B(n10127), 
        .ZN(n10130) );
  NAND2_X1 U11165 ( .A1(n10131), .A2(n10130), .ZN(n10132) );
  OAI21_X1 U11166 ( .B1(n10134), .B2(n10133), .A(n10132), .ZN(n10136) );
  XNOR2_X1 U11167 ( .A(n7999), .B(P2_ADDR_REG_19__SCAN_IN), .ZN(n10135) );
  XNOR2_X1 U11168 ( .A(n10136), .B(n10135), .ZN(n10137) );
  XNOR2_X1 U11169 ( .A(n10138), .B(n10137), .ZN(ADD_1068_U4) );
  AOI21_X1 U11170 ( .B1(n10141), .B2(n10140), .A(n10139), .ZN(ADD_1068_U54) );
  OAI21_X1 U11171 ( .B1(n10144), .B2(n10143), .A(n10142), .ZN(ADD_1068_U47) );
  OAI21_X1 U11172 ( .B1(n10147), .B2(n10146), .A(n10145), .ZN(ADD_1068_U48) );
  OAI21_X1 U11173 ( .B1(n10150), .B2(n10149), .A(n10148), .ZN(ADD_1068_U49) );
  OAI21_X1 U11174 ( .B1(n10153), .B2(n10152), .A(n10151), .ZN(ADD_1068_U50) );
  OAI21_X1 U11175 ( .B1(n10156), .B2(n10155), .A(n10154), .ZN(ADD_1068_U51) );
  AOI21_X1 U11176 ( .B1(n10159), .B2(n10158), .A(n10157), .ZN(ADD_1068_U53) );
  OAI21_X1 U11177 ( .B1(n10162), .B2(n10161), .A(n10160), .ZN(ADD_1068_U52) );
  NAND2_X1 U4860 ( .A1(n4705), .A2(n4703), .ZN(n6939) );
  CLKBUF_X2 U4863 ( .A(n4350), .Z(n4353) );
  CLKBUF_X2 U4943 ( .A(n6091), .Z(n4359) );
  NAND2_X2 U5002 ( .A1(n5726), .A2(n6515), .ZN(n5038) );
  XNOR2_X1 U5015 ( .A(n5981), .B(n7343), .ZN(n7342) );
  AND2_X1 U5059 ( .A1(n9578), .A2(n9577), .ZN(n10165) );
endmodule

