

module b22_C_gen_AntiSAT_k_256_2 ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput_f0, 
        keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, 
        keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, 
        keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, 
        keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, 
        keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, 
        keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, 
        keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, 
        keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, 
        keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, 
        keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, 
        keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, 
        keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, 
        keyinput_f61, keyinput_f62, keyinput_f63, keyinput_f64, keyinput_f65, 
        keyinput_f66, keyinput_f67, keyinput_f68, keyinput_f69, keyinput_f70, 
        keyinput_f71, keyinput_f72, keyinput_f73, keyinput_f74, keyinput_f75, 
        keyinput_f76, keyinput_f77, keyinput_f78, keyinput_f79, keyinput_f80, 
        keyinput_f81, keyinput_f82, keyinput_f83, keyinput_f84, keyinput_f85, 
        keyinput_f86, keyinput_f87, keyinput_f88, keyinput_f89, keyinput_f90, 
        keyinput_f91, keyinput_f92, keyinput_f93, keyinput_f94, keyinput_f95, 
        keyinput_f96, keyinput_f97, keyinput_f98, keyinput_f99, keyinput_f100, 
        keyinput_f101, keyinput_f102, keyinput_f103, keyinput_f104, 
        keyinput_f105, keyinput_f106, keyinput_f107, keyinput_f108, 
        keyinput_f109, keyinput_f110, keyinput_f111, keyinput_f112, 
        keyinput_f113, keyinput_f114, keyinput_f115, keyinput_f116, 
        keyinput_f117, keyinput_f118, keyinput_f119, keyinput_f120, 
        keyinput_f121, keyinput_f122, keyinput_f123, keyinput_f124, 
        keyinput_f125, keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, 
        keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, 
        keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, 
        keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, 
        keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, 
        keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, 
        keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, 
        keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, 
        keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, 
        keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, 
        keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, 
        keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, 
        keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, 
        keyinput_g62, keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, 
        keyinput_g67, keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, 
        keyinput_g72, keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, 
        keyinput_g77, keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, 
        keyinput_g82, keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, 
        keyinput_g87, keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, 
        keyinput_g92, keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, 
        keyinput_g97, keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101, 
        keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105, 
        keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109, 
        keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113, 
        keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117, 
        keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121, 
        keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125, 
        keyinput_g126, keyinput_g127, SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, 
        SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, 
        SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, 
        SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, 
        SUB_1596_U5, SUB_1596_U53, U29, U28, P1_U3355, P1_U3354, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3445, P1_U3446, P1_U3323, P1_U3322, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3459, P1_U3462, 
        P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, 
        P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, 
        P1_U3507, P1_U3510, P1_U3513, P1_U3515, P1_U3516, P1_U3517, P1_U3518, 
        P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, 
        P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, 
        P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, 
        P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, 
        P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, 
        P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3293, 
        P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, 
        P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, 
        P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, 
        P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, 
        P1_U3586, P1_U3587, P1_U3588, P1_U3589, P1_U3590, P1_U3591, P1_U3242, 
        P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3086, P1_U3085, P1_U4016, P2_U3327, P2_U3326, P2_U3325, 
        P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, 
        P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, 
        P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, 
        P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, 
        P2_U3296, P2_U3416, P2_U3417, P2_U3295, P2_U3294, P2_U3293, P2_U3292, 
        P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, 
        P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, 
        P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, 
        P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3430, P2_U3433, 
        P2_U3436, P2_U3439, P2_U3442, P2_U3445, P2_U3448, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3486, P2_U3487, P2_U3488, P2_U3489, 
        P2_U3490, P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, 
        P2_U3497, P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, 
        P2_U3504, P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3265, 
        P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, 
        P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, 
        P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3214, P2_U3531, P2_U3532, P2_U3533, P2_U3534, P2_U3535, 
        P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, P2_U3542, 
        P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, P2_U3549, 
        P2_U3550, P2_U3551, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3328, 
        P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, P2_U3207, 
        P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, 
        P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, 
        P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, 
        P2_U3185, P2_U3088, P2_U3087, P2_U3947, P3_U3295, P3_U3294, P3_U3293, 
        P3_U3292, P3_U3291, P3_U3290, P3_U3289, P3_U3288, P3_U3287, P3_U3286, 
        P3_U3285, P3_U3284, P3_U3283, P3_U3282, P3_U3281, P3_U3280, P3_U3279, 
        P3_U3278, P3_U3277, P3_U3276, P3_U3275, P3_U3274, P3_U3273, P3_U3272, 
        P3_U3271, P3_U3270, P3_U3269, P3_U3268, P3_U3267, P3_U3266, P3_U3265, 
        P3_U3264, P3_U3376, P3_U3377, P3_U3263, P3_U3262, P3_U3261, P3_U3260, 
        P3_U3259, P3_U3258, P3_U3257, P3_U3256, P3_U3255, P3_U3254, P3_U3253, 
        P3_U3252, P3_U3251, P3_U3250, P3_U3249, P3_U3248, P3_U3247, P3_U3246, 
        P3_U3245, P3_U3244, P3_U3243, P3_U3242, P3_U3241, P3_U3240, P3_U3239, 
        P3_U3238, P3_U3237, P3_U3236, P3_U3235, P3_U3234, P3_U3390, P3_U3393, 
        P3_U3396, P3_U3399, P3_U3402, P3_U3405, P3_U3408, P3_U3411, P3_U3414, 
        P3_U3417, P3_U3420, P3_U3423, P3_U3426, P3_U3429, P3_U3432, P3_U3435, 
        P3_U3438, P3_U3441, P3_U3444, P3_U3446, P3_U3447, P3_U3448, P3_U3449, 
        P3_U3450, P3_U3451, P3_U3452, P3_U3453, P3_U3454, P3_U3455, P3_U3456, 
        P3_U3457, P3_U3458, P3_U3459, P3_U3460, P3_U3461, P3_U3462, P3_U3463, 
        P3_U3464, P3_U3465, P3_U3466, P3_U3467, P3_U3468, P3_U3469, P3_U3470, 
        P3_U3471, P3_U3472, P3_U3473, P3_U3474, P3_U3475, P3_U3476, P3_U3477, 
        P3_U3478, P3_U3479, P3_U3480, P3_U3481, P3_U3482, P3_U3483, P3_U3484, 
        P3_U3485, P3_U3486, P3_U3487, P3_U3488, P3_U3489, P3_U3490, P3_U3233, 
        P3_U3232, P3_U3231, P3_U3230, P3_U3229, P3_U3228, P3_U3227, P3_U3226, 
        P3_U3225, P3_U3224, P3_U3223, P3_U3222, P3_U3221, P3_U3220, P3_U3219, 
        P3_U3218, P3_U3217, P3_U3216, P3_U3215, P3_U3214, P3_U3213, P3_U3212, 
        P3_U3211, P3_U3210, P3_U3209, P3_U3208, P3_U3207, P3_U3206, P3_U3205, 
        P3_U3204, P3_U3203, P3_U3202, P3_U3201, P3_U3200, P3_U3199, P3_U3198, 
        P3_U3197, P3_U3196, P3_U3195, P3_U3194, P3_U3193, P3_U3192, P3_U3191, 
        P3_U3190, P3_U3189, P3_U3188, P3_U3187, P3_U3186, P3_U3185, P3_U3184, 
        P3_U3183, P3_U3182, P3_U3491, P3_U3492, P3_U3493, P3_U3494, P3_U3495, 
        P3_U3496, P3_U3497, P3_U3498, P3_U3499, P3_U3500, P3_U3501, P3_U3502, 
        P3_U3503, P3_U3504, P3_U3505, P3_U3506, P3_U3507, P3_U3508, P3_U3509, 
        P3_U3510, P3_U3511, P3_U3512, P3_U3513, P3_U3514, P3_U3515, P3_U3516, 
        P3_U3517, P3_U3518, P3_U3519, P3_U3520, P3_U3521, P3_U3522, P3_U3296, 
        P3_U3181, P3_U3180, P3_U3179, P3_U3178, P3_U3177, P3_U3176, P3_U3175, 
        P3_U3174, P3_U3173, P3_U3172, P3_U3171, P3_U3170, P3_U3169, P3_U3168, 
        P3_U3167, P3_U3166, P3_U3165, P3_U3164, P3_U3163, P3_U3162, P3_U3161, 
        P3_U3160, P3_U3159, P3_U3158, P3_U3157, P3_U3156, P3_U3155, P3_U3154, 
        P3_U3153, P3_U3151, P3_U3150, P3_U3897 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput_f0,
         keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5,
         keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10,
         keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15,
         keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20,
         keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25,
         keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30,
         keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35,
         keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40,
         keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45,
         keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50,
         keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55,
         keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60,
         keyinput_f61, keyinput_f62, keyinput_f63, keyinput_f64, keyinput_f65,
         keyinput_f66, keyinput_f67, keyinput_f68, keyinput_f69, keyinput_f70,
         keyinput_f71, keyinput_f72, keyinput_f73, keyinput_f74, keyinput_f75,
         keyinput_f76, keyinput_f77, keyinput_f78, keyinput_f79, keyinput_f80,
         keyinput_f81, keyinput_f82, keyinput_f83, keyinput_f84, keyinput_f85,
         keyinput_f86, keyinput_f87, keyinput_f88, keyinput_f89, keyinput_f90,
         keyinput_f91, keyinput_f92, keyinput_f93, keyinput_f94, keyinput_f95,
         keyinput_f96, keyinput_f97, keyinput_f98, keyinput_f99, keyinput_f100,
         keyinput_f101, keyinput_f102, keyinput_f103, keyinput_f104,
         keyinput_f105, keyinput_f106, keyinput_f107, keyinput_f108,
         keyinput_f109, keyinput_f110, keyinput_f111, keyinput_f112,
         keyinput_f113, keyinput_f114, keyinput_f115, keyinput_f116,
         keyinput_f117, keyinput_f118, keyinput_f119, keyinput_f120,
         keyinput_f121, keyinput_f122, keyinput_f123, keyinput_f124,
         keyinput_f125, keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1,
         keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6,
         keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11,
         keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16,
         keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21,
         keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26,
         keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31,
         keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36,
         keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41,
         keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46,
         keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51,
         keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56,
         keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61,
         keyinput_g62, keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66,
         keyinput_g67, keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71,
         keyinput_g72, keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76,
         keyinput_g77, keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81,
         keyinput_g82, keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86,
         keyinput_g87, keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91,
         keyinput_g92, keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96,
         keyinput_g97, keyinput_g98, keyinput_g99, keyinput_g100,
         keyinput_g101, keyinput_g102, keyinput_g103, keyinput_g104,
         keyinput_g105, keyinput_g106, keyinput_g107, keyinput_g108,
         keyinput_g109, keyinput_g110, keyinput_g111, keyinput_g112,
         keyinput_g113, keyinput_g114, keyinput_g115, keyinput_g116,
         keyinput_g117, keyinput_g118, keyinput_g119, keyinput_g120,
         keyinput_g121, keyinput_g122, keyinput_g123, keyinput_g124,
         keyinput_g125, keyinput_g126, keyinput_g127;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6669, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679,
         n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689,
         n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699,
         n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709,
         n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719,
         n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729,
         n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739,
         n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749,
         n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759,
         n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769,
         n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779,
         n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789,
         n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799,
         n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809,
         n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819,
         n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829,
         n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839,
         n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849,
         n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859,
         n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869,
         n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879,
         n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889,
         n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899,
         n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909,
         n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919,
         n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929,
         n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939,
         n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949,
         n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959,
         n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969,
         n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979,
         n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989,
         n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999,
         n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009,
         n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019,
         n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029,
         n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039,
         n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049,
         n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059,
         n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069,
         n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079,
         n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089,
         n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099,
         n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109,
         n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119,
         n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129,
         n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139,
         n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149,
         n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159,
         n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169,
         n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179,
         n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189,
         n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199,
         n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209,
         n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219,
         n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229,
         n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239,
         n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249,
         n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259,
         n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269,
         n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279,
         n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289,
         n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299,
         n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309,
         n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319,
         n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329,
         n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339,
         n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349,
         n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359,
         n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369,
         n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379,
         n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389,
         n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399,
         n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409,
         n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419,
         n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429,
         n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439,
         n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449,
         n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459,
         n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469,
         n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479,
         n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489,
         n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499,
         n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509,
         n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519,
         n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529,
         n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539,
         n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549,
         n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559,
         n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569,
         n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579,
         n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589,
         n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599,
         n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609,
         n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619,
         n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629,
         n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639,
         n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649,
         n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659,
         n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669,
         n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679,
         n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689,
         n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699,
         n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709,
         n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719,
         n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729,
         n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739,
         n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749,
         n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759,
         n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769,
         n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779,
         n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789,
         n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799,
         n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809,
         n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819,
         n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829,
         n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839,
         n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849,
         n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859,
         n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869,
         n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879,
         n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889,
         n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899,
         n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909,
         n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919,
         n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929,
         n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939,
         n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949,
         n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959,
         n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969,
         n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979,
         n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989,
         n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999,
         n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009,
         n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019,
         n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029,
         n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039,
         n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049,
         n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059,
         n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069,
         n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079,
         n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089,
         n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099,
         n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109,
         n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119,
         n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129,
         n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139,
         n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149,
         n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159,
         n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169,
         n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179,
         n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189,
         n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199,
         n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209,
         n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219,
         n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229,
         n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239,
         n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249,
         n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259,
         n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269,
         n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279,
         n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289,
         n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299,
         n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309,
         n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319,
         n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329,
         n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339,
         n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349,
         n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359,
         n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369,
         n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379,
         n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389,
         n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399,
         n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409,
         n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419,
         n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429,
         n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439,
         n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449,
         n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459,
         n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469,
         n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479,
         n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489,
         n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499,
         n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509,
         n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519,
         n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529,
         n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539,
         n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549,
         n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559,
         n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569,
         n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579,
         n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589,
         n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599,
         n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609,
         n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619,
         n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629,
         n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639,
         n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649,
         n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659,
         n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669,
         n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679,
         n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689,
         n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699,
         n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709,
         n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719,
         n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729,
         n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739,
         n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749,
         n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759,
         n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769,
         n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779,
         n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789,
         n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799,
         n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809,
         n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819,
         n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829,
         n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839,
         n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849,
         n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859,
         n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869,
         n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879,
         n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889,
         n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899,
         n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909,
         n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919,
         n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929,
         n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939,
         n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949,
         n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959,
         n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969,
         n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979,
         n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989,
         n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999,
         n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009,
         n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019,
         n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029,
         n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039,
         n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049,
         n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059,
         n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069,
         n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079,
         n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089,
         n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099,
         n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109,
         n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119,
         n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129,
         n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139,
         n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149,
         n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159,
         n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169,
         n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179,
         n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189,
         n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199,
         n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209,
         n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219,
         n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229,
         n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239,
         n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249,
         n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259,
         n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269,
         n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279,
         n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289,
         n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299,
         n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309,
         n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319,
         n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329,
         n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339,
         n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349,
         n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359,
         n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369,
         n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379,
         n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389,
         n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399,
         n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409,
         n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419,
         n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429,
         n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439,
         n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449,
         n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459,
         n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469,
         n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479,
         n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489,
         n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499,
         n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509,
         n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519,
         n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529,
         n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539,
         n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549,
         n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559,
         n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569,
         n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579,
         n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589,
         n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599,
         n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609,
         n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619,
         n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629,
         n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639,
         n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649,
         n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659,
         n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669,
         n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679,
         n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689,
         n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699,
         n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709,
         n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719,
         n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729,
         n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739,
         n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749,
         n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759,
         n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769,
         n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779,
         n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789,
         n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799,
         n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809,
         n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819,
         n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829,
         n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839,
         n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849,
         n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859,
         n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869,
         n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879,
         n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889,
         n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899,
         n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909,
         n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919,
         n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929,
         n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939,
         n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949,
         n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959,
         n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969,
         n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979,
         n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989,
         n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999,
         n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
         n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
         n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
         n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703,
         n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
         n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
         n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
         n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
         n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751,
         n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
         n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
         n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
         n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
         n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791,
         n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
         n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807,
         n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
         n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
         n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
         n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
         n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847,
         n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
         n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863,
         n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
         n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
         n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
         n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895,
         n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
         n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911,
         n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919,
         n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
         n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935,
         n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
         n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951,
         n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959,
         n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967,
         n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
         n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983,
         n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991,
         n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
         n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007,
         n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
         n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
         n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031,
         n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039,
         n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047,
         n11048, n11049, n11050, n11052, n11053, n11054, n11055, n11056,
         n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064,
         n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072,
         n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080,
         n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088,
         n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096,
         n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104,
         n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112,
         n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120,
         n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128,
         n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136,
         n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144,
         n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152,
         n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160,
         n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168,
         n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176,
         n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184,
         n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192,
         n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200,
         n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208,
         n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216,
         n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224,
         n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232,
         n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240,
         n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248,
         n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256,
         n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264,
         n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272,
         n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280,
         n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288,
         n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296,
         n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304,
         n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312,
         n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320,
         n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328,
         n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336,
         n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344,
         n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352,
         n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360,
         n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368,
         n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376,
         n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384,
         n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392,
         n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400,
         n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408,
         n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416,
         n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424,
         n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432,
         n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440,
         n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448,
         n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456,
         n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464,
         n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472,
         n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480,
         n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488,
         n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496,
         n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504,
         n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512,
         n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520,
         n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528,
         n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536,
         n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544,
         n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552,
         n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560,
         n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568,
         n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576,
         n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584,
         n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592,
         n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600,
         n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608,
         n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616,
         n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624,
         n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632,
         n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640,
         n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648,
         n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656,
         n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664,
         n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672,
         n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680,
         n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688,
         n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696,
         n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704,
         n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712,
         n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720,
         n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728,
         n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736,
         n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744,
         n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752,
         n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760,
         n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768,
         n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776,
         n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784,
         n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792,
         n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800,
         n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808,
         n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816,
         n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824,
         n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832,
         n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840,
         n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848,
         n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856,
         n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864,
         n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872,
         n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880,
         n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888,
         n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896,
         n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904,
         n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912,
         n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920,
         n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928,
         n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936,
         n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944,
         n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952,
         n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960,
         n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968,
         n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976,
         n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984,
         n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992,
         n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000,
         n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008,
         n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016,
         n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024,
         n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032,
         n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040,
         n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048,
         n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056,
         n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064,
         n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072,
         n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080,
         n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088,
         n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096,
         n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104,
         n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112,
         n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120,
         n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128,
         n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136,
         n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144,
         n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152,
         n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160,
         n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168,
         n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176,
         n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184,
         n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192,
         n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200,
         n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208,
         n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216,
         n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224,
         n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232,
         n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240,
         n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248,
         n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256,
         n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264,
         n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272,
         n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280,
         n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288,
         n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296,
         n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304,
         n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312,
         n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320,
         n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328,
         n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336,
         n12337, n12338, n12339, n12340, n12341, n12342, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13429, n13430, n13431, n13432, n13433, n13434,
         n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442,
         n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450,
         n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458,
         n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466,
         n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474,
         n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482,
         n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490,
         n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498,
         n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506,
         n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514,
         n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522,
         n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530,
         n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538,
         n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546,
         n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554,
         n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562,
         n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570,
         n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578,
         n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586,
         n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594,
         n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602,
         n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610,
         n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618,
         n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626,
         n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634,
         n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642,
         n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650,
         n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658,
         n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666,
         n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674,
         n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682,
         n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690,
         n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698,
         n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706,
         n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714,
         n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722,
         n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730,
         n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738,
         n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746,
         n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754,
         n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762,
         n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770,
         n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778,
         n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786,
         n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794,
         n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802,
         n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810,
         n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818,
         n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826,
         n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834,
         n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842,
         n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850,
         n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858,
         n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866,
         n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874,
         n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882,
         n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890,
         n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898,
         n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906,
         n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914,
         n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922,
         n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930,
         n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938,
         n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946,
         n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954,
         n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962,
         n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970,
         n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978,
         n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986,
         n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994,
         n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002,
         n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010,
         n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018,
         n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026,
         n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034,
         n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042,
         n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050,
         n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058,
         n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066,
         n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074,
         n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082,
         n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090,
         n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098,
         n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106,
         n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114,
         n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122,
         n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130,
         n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138,
         n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146,
         n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154,
         n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162,
         n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170,
         n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178,
         n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186,
         n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194,
         n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202,
         n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210,
         n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218,
         n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226,
         n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14234,
         n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242,
         n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250,
         n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258,
         n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266,
         n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274,
         n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282,
         n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290,
         n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298,
         n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306,
         n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314,
         n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322,
         n14323, n14324, n14325, n14326, n14327, n14328, n14329, n14330,
         n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338,
         n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346,
         n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354,
         n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362,
         n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370,
         n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378,
         n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386,
         n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394,
         n14395, n14396, n14397, n14398, n14399, n14400, n14401, n14402,
         n14403, n14404, n14405, n14406, n14407, n14408, n14409, n14410,
         n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418,
         n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426,
         n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434,
         n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442,
         n14443, n14444, n14445, n14446, n14447, n14448, n14449, n14450,
         n14451, n14452, n14453, n14454, n14455, n14456, n14457, n14458,
         n14459, n14460, n14461, n14462, n14463, n14464, n14465, n14466,
         n14467, n14468, n14469, n14470, n14471, n14472, n14473, n14474,
         n14475, n14476, n14477, n14478, n14479, n14480, n14481, n14482,
         n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490,
         n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498,
         n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506,
         n14507, n14508, n14509, n14510, n14511, n14512, n14513, n14514,
         n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522,
         n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530,
         n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538,
         n14539, n14540, n14541, n14542, n14543, n14544, n14545, n14546,
         n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554,
         n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562,
         n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570,
         n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578,
         n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586,
         n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594,
         n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602,
         n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14610,
         n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618,
         n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626,
         n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634,
         n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642,
         n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650,
         n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658,
         n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666,
         n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674,
         n14675, n14676, n14677, n14678, n14679, n14680, n14681, n14682,
         n14683, n14684, n14685, n14686, n14687, n14688, n14689, n14690,
         n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698,
         n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706,
         n14707, n14708, n14709, n14710, n14711, n14712, n14713, n14714,
         n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722,
         n14723, n14724, n14725, n14726, n14727, n14728, n14729, n14730,
         n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738,
         n14739, n14740, n14741, n14742, n14743, n14744, n14745, n14746,
         n14747, n14748, n14749, n14750, n14751, n14752, n14753, n14754,
         n14755, n14756, n14757, n14758, n14759, n14760, n14761, n14762,
         n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770,
         n14771, n14772, n14773, n14774, n14775, n14776, n14777, n14778,
         n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786,
         n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794,
         n14795, n14796, n14797, n14798, n14799, n14800, n14801, n14802,
         n14803, n14804, n14805, n14806, n14807, n14808, n14809, n14810,
         n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818,
         n14819, n14820, n14821, n14822, n14823, n14824, n14825, n14826,
         n14827, n14828, n14829, n14830, n14831, n14832, n14833, n14834,
         n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14842,
         n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850,
         n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858,
         n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866,
         n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874,
         n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882,
         n14883, n14884, n14885, n14886, n14888, n14889, n14890, n14891,
         n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899,
         n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907,
         n14908, n14909, n14910, n14911, n14912, n14913, n14914, n14915,
         n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923,
         n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931,
         n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939,
         n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947,
         n14948, n14949, n14950, n14951, n14952, n14953, n14954, n14955,
         n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963,
         n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971,
         n14972, n14973, n14974, n14975, n14976, n14977, n14978, n14979,
         n14980, n14981, n14982, n14983, n14984, n14985, n14986, n14987,
         n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995,
         n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003,
         n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011,
         n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019,
         n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027,
         n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15035,
         n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043,
         n15044, n15045, n15046, n15047, n15048, n15049, n15050, n15051,
         n15052, n15053, n15054, n15055, n15056, n15057, n15058, n15059,
         n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067,
         n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075,
         n15076, n15077, n15078, n15079, n15080, n15081, n15082, n15083,
         n15084, n15085, n15086, n15087, n15088, n15089, n15090, n15091,
         n15092, n15093, n15094, n15095, n15096, n15097, n15098, n15099,
         n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107,
         n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115,
         n15116, n15117, n15118, n15119, n15120, n15121, n15122, n15123,
         n15124, n15125, n15126, n15127, n15128, n15129, n15130, n15131,
         n15132, n15133, n15134, n15135, n15136, n15137, n15138, n15139,
         n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147,
         n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155,
         n15156, n15157, n15158, n15159, n15160, n15161, n15162, n15163,
         n15164, n15165, n15166, n15167, n15168, n15169, n15170, n15171,
         n15172, n15173, n15174, n15175, n15176, n15177, n15178, n15179,
         n15180, n15181, n15182, n15183, n15184, n15185, n15186, n15187,
         n15188, n15189, n15190, n15191, n15192, n15193, n15194, n15195,
         n15196, n15197, n15198, n15199, n15200, n15201, n15202, n15203,
         n15204, n15205, n15206, n15207, n15208, n15209, n15210, n15211,
         n15212, n15213, n15214, n15215, n15216, n15217, n15218, n15219,
         n15220, n15221, n15222, n15223, n15224, n15225, n15226, n15227,
         n15228, n15229, n15230, n15231, n15232, n15233, n15234, n15235,
         n15236, n15237, n15238, n15239, n15240, n15241, n15242, n15243,
         n15244, n15245, n15246, n15247, n15248, n15249, n15250, n15251,
         n15252, n15253, n15254, n15255, n15256, n15257, n15258, n15259,
         n15260, n15261, n15262, n15263, n15264, n15265, n15266, n15267,
         n15268, n15269, n15270, n15271, n15272, n15273, n15274, n15275,
         n15276, n15277, n15278, n15279, n15280, n15281, n15282, n15283,
         n15284, n15285, n15286, n15287, n15288, n15289, n15290, n15291,
         n15292, n15293, n15294, n15295, n15296, n15297, n15298, n15299,
         n15300, n15301, n15302, n15303, n15304, n15305, n15306, n15307,
         n15308, n15309, n15310, n15311, n15312, n15313, n15314, n15315,
         n15316, n15317, n15318, n15319, n15320, n15321, n15322, n15323,
         n15324, n15325, n15326, n15327, n15328, n15329, n15330, n15331,
         n15332, n15333, n15334, n15335, n15336, n15337, n15338, n15339,
         n15340, n15341, n15342, n15343, n15344, n15345, n15346, n15347,
         n15348, n15349, n15350, n15351, n15352, n15353, n15354, n15355,
         n15356, n15357, n15358, n15359, n15360, n15361, n15362, n15363,
         n15364, n15365, n15366, n15367, n15368, n15369, n15370, n15371,
         n15372, n15373, n15374, n15375, n15376, n15377, n15378, n15379,
         n15380, n15381, n15382, n15383, n15384, n15385, n15386, n15387,
         n15388, n15389, n15390, n15391, n15392, n15393, n15394, n15395,
         n15396, n15397, n15398, n15399, n15400, n15401, n15402, n15403,
         n15404, n15405, n15406, n15407, n15408, n15409, n15410, n15411,
         n15412, n15413, n15414, n15415, n15416, n15417, n15418, n15419,
         n15420, n15421, n15422, n15423, n15424, n15425, n15426, n15427,
         n15428, n15429, n15430, n15431, n15432, n15433, n15434, n15436,
         n15437, n15438, n15439, n15440, n15441, n15442, n15443, n15444,
         n15445, n15446, n15447, n15448, n15449, n15450, n15451, n15452,
         n15453, n15454, n15455, n15456, n15457, n15458, n15459, n15460,
         n15461, n15462, n15463, n15464, n15465, n15466, n15467, n15468,
         n15469, n15470, n15471, n15472, n15473, n15474, n15475, n15476,
         n15477, n15478, n15479, n15480, n15481, n15482, n15483, n15484,
         n15485, n15486, n15487, n15488, n15489, n15490, n15491, n15492,
         n15493, n15494, n15495, n15496, n15497, n15498, n15499, n15500,
         n15501, n15502, n15503, n15504, n15505, n15506, n15507, n15508,
         n15509, n15510, n15511, n15512, n15513, n15514, n15515, n15516,
         n15517, n15518, n15519, n15520, n15521, n15522, n15523, n15524,
         n15525, n15526, n15527, n15528, n15529, n15530, n15531, n15532,
         n15533, n15534, n15535, n15536, n15537, n15538, n15539, n15540,
         n15541, n15542, n15543, n15544, n15545, n15546, n15547, n15548,
         n15549, n15550, n15551, n15552, n15553, n15554, n15555, n15556,
         n15557, n15558, n15559, n15560, n15561, n15562, n15563, n15564,
         n15565, n15566, n15567, n15568, n15569, n15570, n15571, n15572,
         n15573, n15574, n15575, n15576, n15577, n15578, n15579, n15580,
         n15581, n15582, n15583, n15584, n15585, n15586, n15587, n15588,
         n15589, n15590, n15591, n15592, n15593, n15594, n15595, n15596,
         n15597, n15598, n15599, n15600, n15601, n15602, n15603, n15604,
         n15605, n15606, n15607, n15608, n15609, n15610, n15611, n15612,
         n15613, n15614, n15615, n15616, n15617, n15618, n15619, n15620,
         n15621, n15622, n15623, n15624, n15625, n15626, n15627, n15628,
         n15629, n15630, n15631, n15632, n15633, n15634, n15635, n15636,
         n15637, n15638, n15639, n15640, n15641, n15642, n15643, n15644,
         n15645, n15646, n15647, n15648, n15649, n15650, n15651, n15652,
         n15653, n15654, n15655, n15656, n15657, n15658, n15659, n15660,
         n15661, n15662, n15663, n15664, n15665, n15666, n15667, n15668,
         n15669, n15670, n15671, n15672, n15673, n15674, n15675, n15676,
         n15677, n15678, n15679, n15680, n15681, n15682, n15683, n15684,
         n15685, n15686, n15687, n15688, n15689, n15690, n15691, n15692,
         n15693, n15694, n15695, n15696, n15697, n15698, n15699, n15700,
         n15701, n15702, n15703, n15704, n15705, n15706, n15707, n15708,
         n15709, n15710, n15711, n15712, n15713, n15714, n15715, n15716,
         n15717, n15718, n15719, n15720, n15721, n15722, n15723, n15724,
         n15725, n15726, n15727, n15728, n15729, n15730, n15731, n15732,
         n15733, n15734, n15735, n15736, n15737, n15738, n15739, n15740,
         n15741, n15742, n15743, n15744, n15745, n15746, n15747, n15748,
         n15749, n15750, n15751, n15752, n15753, n15754, n15755, n15756,
         n15757, n15758, n15759, n15760, n15761, n15762, n15763, n15764,
         n15765, n15766, n15767, n15768;

  AND2_X1 U7417 ( .A1(n13939), .A2(n13942), .ZN(n14023) );
  NAND2_X2 U7418 ( .A1(n6671), .A2(P3_U3151), .ZN(n13440) );
  AND2_X1 U7419 ( .A1(n8261), .A2(n8260), .ZN(n14032) );
  OAI21_X1 U7420 ( .B1(n15210), .B2(n15211), .A(n7205), .ZN(n7204) );
  NAND2_X1 U7421 ( .A1(n6878), .A2(n7560), .ZN(n13512) );
  INV_X1 U7422 ( .A(n12648), .ZN(n12635) );
  NAND2_X2 U7423 ( .A1(n10727), .A2(n14212), .ZN(n12646) );
  OR2_X1 U7424 ( .A1(n15682), .A2(n15695), .ZN(n12845) );
  CLKBUF_X2 U7425 ( .A(n7777), .Z(n9223) );
  CLKBUF_X2 U7426 ( .A(n8480), .Z(n11989) );
  NAND2_X2 U7427 ( .A1(n8280), .A2(n8286), .ZN(n9029) );
  NAND2_X1 U7428 ( .A1(n13431), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8450) );
  CLKBUF_X1 U7429 ( .A(n8286), .Z(n12137) );
  INV_X1 U7430 ( .A(n14390), .ZN(n14411) );
  INV_X1 U7431 ( .A(n11986), .ZN(n8960) );
  AND2_X1 U7433 ( .A1(n8332), .A2(n12531), .ZN(n11490) );
  OAI21_X1 U7434 ( .B1(n11480), .B2(n9725), .A(n9726), .ZN(n11620) );
  INV_X1 U7435 ( .A(n8480), .ZN(n8798) );
  AND2_X1 U7436 ( .A1(n12990), .A2(n12848), .ZN(n12963) );
  NAND2_X1 U7437 ( .A1(n11761), .A2(n11760), .ZN(n11875) );
  INV_X2 U7438 ( .A(n11777), .ZN(n13912) );
  NOR2_X2 U7440 ( .A1(n11958), .A2(n14019), .ZN(n7173) );
  NAND2_X1 U7441 ( .A1(n7714), .A2(n7326), .ZN(n7913) );
  AND3_X1 U7442 ( .A1(n6677), .A2(n6692), .A3(n7567), .ZN(n8097) );
  BUF_X1 U7443 ( .A(n14376), .Z(n9633) );
  NAND2_X1 U7444 ( .A1(n8224), .A2(n8223), .ZN(n8240) );
  INV_X1 U7445 ( .A(n8855), .ZN(n10432) );
  OAI21_X1 U7446 ( .B1(n9813), .B2(n7352), .A(n7350), .ZN(n11830) );
  NAND2_X1 U7447 ( .A1(n7953), .A2(n7952), .ZN(n14019) );
  NAND2_X1 U7448 ( .A1(n8191), .A2(n8190), .ZN(n13965) );
  INV_X1 U7449 ( .A(n8253), .ZN(n8338) );
  INV_X2 U7450 ( .A(n8410), .ZN(n11777) );
  NAND2_X1 U7451 ( .A1(n9642), .A2(n9641), .ZN(n14812) );
  NAND2_X1 U7452 ( .A1(n9578), .A2(n9577), .ZN(n14851) );
  OAI211_X1 U7453 ( .C1(n9370), .C2(n10466), .A(n7510), .B(n7509), .ZN(n11189)
         );
  NAND2_X1 U7454 ( .A1(n8891), .A2(n8890), .ZN(n13127) );
  INV_X2 U7455 ( .A(n6669), .ZN(n9049) );
  XNOR2_X1 U7456 ( .A(n9337), .B(n9336), .ZN(n14883) );
  INV_X2 U7457 ( .A(n14381), .ZN(n9753) );
  OR2_X1 U7458 ( .A1(n11712), .A2(n11713), .ZN(n7521) );
  NOR2_X2 U7459 ( .A1(n15219), .A2(n15218), .ZN(n15217) );
  XNOR2_X2 U7460 ( .A(n12997), .B(n13015), .ZN(n15568) );
  OAI21_X2 U7461 ( .B1(n14658), .B2(n7477), .A(n7475), .ZN(n14634) );
  AOI21_X2 U7462 ( .B1(n14191), .B2(n14674), .A(n14662), .ZN(n14658) );
  XNOR2_X2 U7463 ( .A(n13477), .B(n13475), .ZN(n13503) );
  OAI21_X2 U7464 ( .B1(n13141), .B2(n13126), .A(n7122), .ZN(n13109) );
  NAND2_X1 U7465 ( .A1(n9724), .A2(n9723), .ZN(n11480) );
  NAND2_X2 U7466 ( .A1(n13588), .A2(n13474), .ZN(n13477) );
  AOI22_X2 U7467 ( .A1(n14293), .A2(n14292), .B1(n14291), .B2(n14290), .ZN(
        n14296) );
  BUF_X4 U7468 ( .A(n9086), .Z(n6669) );
  NAND2_X1 U7469 ( .A1(n11493), .A2(n12531), .ZN(n9086) );
  XNOR2_X2 U7470 ( .A(n8450), .B(n6968), .ZN(n12684) );
  OAI22_X2 U7471 ( .A1(n14756), .A2(n7604), .B1(n7605), .B2(n7603), .ZN(n14728) );
  XNOR2_X2 U7472 ( .A(n12465), .B(n12463), .ZN(n12462) );
  NOR2_X2 U7473 ( .A1(n9983), .A2(n9982), .ZN(n15205) );
  NAND2_X2 U7474 ( .A1(n12305), .A2(n12304), .ZN(n12465) );
  AOI21_X2 U7475 ( .B1(n9932), .B2(n9926), .A(n9930), .ZN(n9927) );
  NAND2_X2 U7476 ( .A1(n15757), .A2(n15756), .ZN(n15755) );
  XNOR2_X2 U7477 ( .A(n9959), .B(n6871), .ZN(n15757) );
  BUF_X8 U7479 ( .A(n10432), .Z(n6671) );
  NAND2_X2 U7480 ( .A1(n15752), .A2(n9957), .ZN(n9959) );
  NAND2_X2 U7481 ( .A1(n12667), .A2(n6675), .ZN(n8465) );
  OAI21_X2 U7482 ( .B1(n12503), .B2(n7109), .A(n7106), .ZN(n12556) );
  NOR2_X2 U7484 ( .A1(n12996), .A2(n6823), .ZN(n12997) );
  NAND2_X2 U7485 ( .A1(n15759), .A2(n9968), .ZN(n9970) );
  XNOR2_X1 U7486 ( .A(n9963), .B(n7231), .ZN(n14904) );
  INV_X2 U7487 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n7029) );
  NAND2_X2 U7488 ( .A1(n15755), .A2(n9960), .ZN(n9963) );
  XNOR2_X2 U7489 ( .A(n14507), .B(P3_ADDR_REG_1__SCAN_IN), .ZN(n9949) );
  INV_X2 U7490 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n14507) );
  AOI21_X2 U7491 ( .B1(P3_ADDR_REG_12__SCAN_IN), .B2(n15256), .A(n9922), .ZN(
        n9981) );
  NAND2_X1 U7492 ( .A1(n14123), .A2(n12628), .ZN(n14188) );
  NOR2_X1 U7493 ( .A1(n9190), .A2(n9189), .ZN(n9192) );
  INV_X2 U7494 ( .A(n14032), .ZN(n13541) );
  OAI21_X1 U7495 ( .B1(n13223), .B2(n7399), .A(n12940), .ZN(n13209) );
  NAND2_X1 U7496 ( .A1(n7204), .A2(n15209), .ZN(n15214) );
  OR2_X1 U7497 ( .A1(n9111), .A2(n9110), .ZN(n9116) );
  AND2_X1 U7498 ( .A1(n7179), .A2(n15200), .ZN(n9983) );
  NAND2_X1 U7499 ( .A1(n7173), .A2(n7172), .ZN(n12204) );
  OAI21_X1 U7500 ( .B1(n11740), .B2(n7517), .A(n7516), .ZN(n7515) );
  INV_X1 U7501 ( .A(n9870), .ZN(n7125) );
  INV_X1 U7502 ( .A(n14228), .ZN(n6672) );
  NAND2_X2 U7503 ( .A1(n12864), .A2(n12861), .ZN(n11373) );
  INV_X4 U7504 ( .A(n12645), .ZN(n12621) );
  INV_X1 U7505 ( .A(n14498), .ZN(n11445) );
  NAND2_X1 U7506 ( .A1(n9382), .A2(n9381), .ZN(n14224) );
  CLKBUF_X2 U7507 ( .A(n9226), .Z(n9241) );
  CLKBUF_X3 U7508 ( .A(n9049), .Z(n9226) );
  INV_X2 U7509 ( .A(n9049), .ZN(n9239) );
  NAND2_X1 U7510 ( .A1(n12854), .A2(n12859), .ZN(n12857) );
  INV_X1 U7511 ( .A(n14337), .ZN(n14390) );
  NAND2_X1 U7512 ( .A1(n12850), .A2(n12845), .ZN(n15702) );
  NOR2_X1 U7513 ( .A1(n11368), .A2(n15699), .ZN(n15696) );
  INV_X4 U7514 ( .A(n12963), .ZN(n12975) );
  NAND2_X1 U7515 ( .A1(n15682), .A2(n15695), .ZN(n12850) );
  INV_X1 U7516 ( .A(n12531), .ZN(n7564) );
  CLKBUF_X2 U7517 ( .A(n8623), .Z(n12806) );
  INV_X2 U7518 ( .A(n13037), .ZN(n7356) );
  INV_X4 U7519 ( .A(n9370), .ZN(n14407) );
  XNOR2_X1 U7520 ( .A(n9905), .B(P3_ADDR_REG_4__SCAN_IN), .ZN(n9943) );
  NAND3_X1 U7521 ( .A1(n7722), .A2(n6885), .A3(n7739), .ZN(n7743) );
  INV_X2 U7522 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  OAI21_X1 U7523 ( .B1(n14030), .B2(n15523), .A(n7097), .ZN(n14031) );
  OAI21_X1 U7524 ( .B1(n9207), .B2(n7003), .A(n7002), .ZN(n9294) );
  NAND2_X1 U7525 ( .A1(n14188), .A2(n14189), .ZN(n14187) );
  AOI21_X1 U7526 ( .B1(n9198), .B2(n9197), .A(n6974), .ZN(n9200) );
  AOI21_X1 U7527 ( .B1(n8909), .B2(n12842), .A(n13085), .ZN(n8969) );
  NOR4_X1 U7528 ( .A1(n9288), .A2(n9287), .A3(n9286), .A4(n9285), .ZN(n9290)
         );
  NAND2_X1 U7529 ( .A1(n8238), .A2(n7489), .ZN(n13947) );
  NAND2_X1 U7530 ( .A1(n13479), .A2(n13478), .ZN(n13570) );
  OAI21_X1 U7531 ( .B1(n9192), .B2(n9191), .A(n6977), .ZN(n6976) );
  AND2_X1 U7532 ( .A1(n8400), .A2(n8271), .ZN(n9284) );
  XNOR2_X1 U7533 ( .A(n13744), .B(n9225), .ZN(n9286) );
  NAND2_X1 U7534 ( .A1(n14896), .A2(n14895), .ZN(n14894) );
  OAI21_X1 U7535 ( .B1(n14896), .B2(n14895), .A(n7230), .ZN(n7229) );
  NAND2_X1 U7536 ( .A1(n14682), .A2(n7613), .ZN(n14797) );
  AND2_X1 U7537 ( .A1(n9236), .A2(n9235), .ZN(n14029) );
  XNOR2_X1 U7538 ( .A(n9209), .B(n9208), .ZN(n14071) );
  NAND2_X1 U7539 ( .A1(n9651), .A2(n14694), .ZN(n14814) );
  NAND2_X1 U7540 ( .A1(n9739), .A2(n9677), .ZN(n14657) );
  NAND2_X1 U7541 ( .A1(n13156), .A2(n8953), .ZN(n13145) );
  AOI21_X2 U7542 ( .B1(n14079), .B2(n9234), .A(n6795), .ZN(n13766) );
  NAND2_X1 U7543 ( .A1(n8227), .A2(n8226), .ZN(n13778) );
  OR2_X1 U7544 ( .A1(n8256), .A2(n8255), .ZN(n8259) );
  NOR2_X1 U7545 ( .A1(n14967), .A2(n13003), .ZN(n14986) );
  OR2_X1 U7546 ( .A1(n12469), .A2(n6893), .ZN(n6887) );
  NAND2_X1 U7547 ( .A1(n7128), .A2(n6731), .ZN(n13347) );
  NAND2_X1 U7548 ( .A1(n9617), .A2(n9616), .ZN(n14827) );
  OAI21_X1 U7549 ( .B1(n8202), .B2(n7223), .A(n8205), .ZN(n8222) );
  NAND2_X1 U7550 ( .A1(n9355), .A2(n9354), .ZN(n14758) );
  XNOR2_X1 U7551 ( .A(n8204), .B(SI_24_), .ZN(n8202) );
  NAND2_X1 U7552 ( .A1(n8101), .A2(n8100), .ZN(n13893) );
  NAND2_X1 U7553 ( .A1(n8189), .A2(n8188), .ZN(n8204) );
  NAND2_X1 U7554 ( .A1(n8126), .A2(n8125), .ZN(n13986) );
  NAND2_X1 U7555 ( .A1(n8083), .A2(n8082), .ZN(n14053) );
  OR2_X1 U7556 ( .A1(n12232), .A2(n14438), .ZN(n15163) );
  NAND2_X1 U7557 ( .A1(n8182), .A2(n8181), .ZN(n8189) );
  NOR2_X1 U7558 ( .A1(n15599), .A2(n13001), .ZN(n15618) );
  OAI21_X2 U7559 ( .B1(n8137), .B2(n7018), .A(n7016), .ZN(n8182) );
  OR2_X1 U7560 ( .A1(n9107), .A2(n9106), .ZN(n9111) );
  NAND2_X1 U7561 ( .A1(n8124), .A2(n8123), .ZN(n8137) );
  NAND2_X1 U7562 ( .A1(n12241), .A2(n12240), .ZN(n12246) );
  NAND2_X1 U7563 ( .A1(n12086), .A2(n12109), .ZN(n12241) );
  NAND2_X1 U7564 ( .A1(n8055), .A2(n8054), .ZN(n13443) );
  XNOR2_X1 U7565 ( .A(n13000), .B(n13020), .ZN(n15600) );
  OAI21_X1 U7566 ( .B1(n15568), .B2(n7291), .A(n7290), .ZN(n15583) );
  NAND2_X1 U7567 ( .A1(n7171), .A2(n12205), .ZN(n12263) );
  NAND2_X1 U7568 ( .A1(n15643), .A2(n12895), .ZN(n15048) );
  INV_X1 U7569 ( .A(n12204), .ZN(n7171) );
  NAND2_X1 U7570 ( .A1(n7397), .A2(n6735), .ZN(n15643) );
  NAND2_X1 U7571 ( .A1(n7998), .A2(n7997), .ZN(n12277) );
  OAI211_X1 U7572 ( .C1(n6973), .C2(n6970), .A(n6971), .B(n6969), .ZN(n7660)
         );
  NAND2_X1 U7573 ( .A1(n11830), .A2(n9820), .ZN(n12046) );
  NAND2_X1 U7574 ( .A1(n12187), .A2(n12893), .ZN(n7397) );
  OR2_X1 U7575 ( .A1(n14911), .A2(n14910), .ZN(n7178) );
  AND2_X1 U7576 ( .A1(n11739), .A2(n11738), .ZN(n11740) );
  INV_X1 U7577 ( .A(n13220), .ZN(n6673) );
  CLKBUF_X2 U7578 ( .A(n13220), .Z(n6674) );
  NAND2_X1 U7579 ( .A1(n7160), .A2(n7159), .ZN(n11636) );
  NAND2_X1 U7580 ( .A1(n7935), .A2(n7934), .ZN(n12068) );
  OR2_X1 U7581 ( .A1(n7993), .A2(SI_14_), .ZN(n8008) );
  NAND2_X1 U7582 ( .A1(n7919), .A2(n7918), .ZN(n15507) );
  NAND2_X1 U7583 ( .A1(n11676), .A2(n7638), .ZN(n11792) );
  AND2_X1 U7584 ( .A1(n15577), .A2(n15576), .ZN(n15578) );
  OAI21_X1 U7585 ( .B1(n7992), .B2(n7678), .A(n7991), .ZN(n7993) );
  CLKBUF_X1 U7586 ( .A(n13303), .Z(n15714) );
  NOR2_X1 U7587 ( .A1(n11047), .A2(n11045), .ZN(n13605) );
  NAND2_X1 U7588 ( .A1(n11593), .A2(n15488), .ZN(n11635) );
  NAND2_X1 U7589 ( .A1(n7911), .A2(n7910), .ZN(n7931) );
  NAND2_X1 U7590 ( .A1(n11363), .A2(n15675), .ZN(n15693) );
  NOR2_X1 U7591 ( .A1(n14904), .A2(n14905), .ZN(n14903) );
  NOR2_X1 U7592 ( .A1(n7514), .A2(n6763), .ZN(n10814) );
  NAND2_X1 U7593 ( .A1(n7835), .A2(n7836), .ZN(n11429) );
  AND2_X1 U7594 ( .A1(n9042), .A2(n9041), .ZN(n9046) );
  NOR2_X1 U7595 ( .A1(n9910), .A2(n6827), .ZN(n9912) );
  BUF_X1 U7596 ( .A(n14505), .Z(n6808) );
  INV_X2 U7597 ( .A(n11014), .ZN(n10728) );
  OR2_X1 U7598 ( .A1(n8738), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n8755) );
  NAND2_X1 U7599 ( .A1(n7773), .A2(n7772), .ZN(n13515) );
  OR2_X2 U7600 ( .A1(n12648), .A2(n15122), .ZN(n11014) );
  NAND2_X1 U7601 ( .A1(n7830), .A2(n7829), .ZN(n7848) );
  NAND2_X1 U7602 ( .A1(n7723), .A2(n7724), .ZN(n11129) );
  NAND4_X1 U7603 ( .A1(n7781), .A2(n7780), .A3(n7779), .A4(n7778), .ZN(n13655)
         );
  NAND4_X1 U7604 ( .A1(n9422), .A2(n9421), .A3(n9420), .A4(n9419), .ZN(n14498)
         );
  NAND2_X1 U7605 ( .A1(n7746), .A2(n7745), .ZN(n13932) );
  AND2_X1 U7606 ( .A1(n10734), .A2(n14218), .ZN(n11192) );
  NAND4_X1 U7607 ( .A1(n7751), .A2(n7750), .A3(n7749), .A4(n7748), .ZN(n13658)
         );
  AND2_X2 U7608 ( .A1(n6681), .A2(n14381), .ZN(n15122) );
  AND2_X1 U7609 ( .A1(n8468), .A2(n7396), .ZN(n11368) );
  BUF_X2 U7610 ( .A(n9582), .Z(n6841) );
  AND2_X1 U7611 ( .A1(n9753), .A2(n14387), .ZN(n14218) );
  NAND4_X1 U7612 ( .A1(n8498), .A2(n8497), .A3(n8496), .A4(n8495), .ZN(n15681)
         );
  NAND4_X1 U7613 ( .A1(n8458), .A2(n8457), .A3(n8456), .A4(n8455), .ZN(n15699)
         );
  CLKBUF_X3 U7614 ( .A(n9418), .Z(n14376) );
  BUF_X2 U7615 ( .A(n7774), .Z(n9219) );
  CLKBUF_X2 U7616 ( .A(n7818), .Z(n9234) );
  XNOR2_X1 U7617 ( .A(n7564), .B(n9029), .ZN(n7563) );
  AND2_X1 U7618 ( .A1(n14878), .A2(n9325), .ZN(n9582) );
  NAND2_X1 U7619 ( .A1(n9742), .A2(n14619), .ZN(n14212) );
  AOI21_X1 U7620 ( .B1(n9943), .B2(n15239), .A(n9906), .ZN(n9907) );
  XNOR2_X1 U7621 ( .A(n8912), .B(n8911), .ZN(n11681) );
  INV_X2 U7622 ( .A(n13039), .ZN(n13027) );
  NAND2_X1 U7623 ( .A1(n10483), .A2(n6671), .ZN(n9371) );
  AND2_X2 U7624 ( .A1(n7734), .A2(n7733), .ZN(n8253) );
  XNOR2_X1 U7625 ( .A(n7731), .B(P2_IR_REG_30__SCAN_IN), .ZN(n7734) );
  MUX2_X1 U7626 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9705), .S(
        P1_IR_REG_21__SCAN_IN), .Z(n9707) );
  MUX2_X1 U7627 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9702), .S(
        P1_IR_REG_22__SCAN_IN), .Z(n9703) );
  XNOR2_X1 U7628 ( .A(n9710), .B(n9709), .ZN(n14387) );
  NAND2_X1 U7629 ( .A1(n9353), .A2(n9708), .ZN(n14619) );
  MUX2_X1 U7630 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8281), .S(
        P2_IR_REG_22__SCAN_IN), .Z(n8285) );
  NAND2_X1 U7631 ( .A1(n8284), .A2(n8283), .ZN(n8381) );
  NAND2_X1 U7632 ( .A1(n7729), .A2(n7730), .ZN(n14074) );
  NAND2_X1 U7633 ( .A1(n14872), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7403) );
  NAND2_X1 U7634 ( .A1(n7827), .A2(SI_6_), .ZN(n7847) );
  XNOR2_X1 U7635 ( .A(n8463), .B(n8462), .ZN(n13029) );
  INV_X1 U7636 ( .A(n10929), .ZN(n7299) );
  NAND2_X1 U7637 ( .A1(n6867), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n11303) );
  NAND2_X1 U7638 ( .A1(n9323), .A2(n9322), .ZN(n14872) );
  MUX2_X1 U7639 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8275), .S(
        P2_IR_REG_21__SCAN_IN), .Z(n8276) );
  NAND2_X1 U7640 ( .A1(n7591), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9337) );
  AND2_X2 U7641 ( .A1(n9332), .A2(n9321), .ZN(n9323) );
  NOR2_X1 U7642 ( .A1(n6960), .A2(n6959), .ZN(n8451) );
  AOI21_X1 U7643 ( .B1(n6875), .B2(n6874), .A(n7226), .ZN(n9948) );
  NAND2_X2 U7644 ( .A1(n7073), .A2(n7072), .ZN(n10433) );
  AND2_X1 U7645 ( .A1(n7134), .A2(n7683), .ZN(n9319) );
  NAND4_X2 U7646 ( .A1(n7026), .A2(n7028), .A3(n7025), .A4(n7024), .ZN(n10967)
         );
  NAND2_X1 U7647 ( .A1(n8533), .A2(n7635), .ZN(n7634) );
  AND2_X1 U7648 ( .A1(n7030), .A2(n7029), .ZN(n7289) );
  AND2_X1 U7649 ( .A1(n8534), .A2(n8447), .ZN(n7635) );
  CLKBUF_X1 U7650 ( .A(n9515), .Z(n10050) );
  INV_X1 U7651 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n7791) );
  NOR2_X1 U7652 ( .A1(P3_IR_REG_4__SCAN_IN), .A2(P3_IR_REG_2__SCAN_IN), .ZN(
        n7348) );
  INV_X1 U7653 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n8426) );
  INV_X1 U7654 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n7030) );
  NOR2_X1 U7655 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .ZN(
        n7347) );
  INV_X1 U7656 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n9489) );
  INV_X1 U7657 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n7694) );
  INV_X1 U7658 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n9411) );
  INV_X4 U7659 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  INV_X1 U7660 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n7854) );
  INV_X1 U7661 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n9436) );
  NOR2_X1 U7662 ( .A1(P3_IR_REG_25__SCAN_IN), .A2(P3_IR_REG_26__SCAN_IN), .ZN(
        n7395) );
  INV_X4 U7663 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U7664 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n9515) );
  INV_X1 U7665 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n8697) );
  NOR2_X1 U7666 ( .A1(P3_IR_REG_9__SCAN_IN), .A2(P3_IR_REG_11__SCAN_IN), .ZN(
        n8428) );
  NOR2_X1 U7667 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n9307) );
  CLKBUF_X1 U7668 ( .A(P1_IR_REG_7__SCAN_IN), .Z(n10312) );
  INV_X1 U7669 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n9545) );
  NOR2_X2 U7670 ( .A1(n14742), .A2(n14827), .ZN(n14729) );
  NAND2_X4 U7671 ( .A1(n7713), .A2(n7714), .ZN(n7821) );
  NAND2_X2 U7672 ( .A1(n8831), .A2(n8830), .ZN(n13159) );
  XNOR2_X1 U7673 ( .A(n11736), .B(n11737), .ZN(n11712) );
  AND4_X2 U7674 ( .A1(n9385), .A2(n9384), .A3(n9387), .A4(n9386), .ZN(n11203)
         );
  NOR2_X1 U7675 ( .A1(n11018), .A2(n6752), .ZN(n11197) );
  NOR2_X2 U7676 ( .A1(n14918), .A2(n14917), .ZN(n14957) );
  XNOR2_X1 U7677 ( .A(n8463), .B(n8462), .ZN(n6675) );
  CLKBUF_X1 U7678 ( .A(n14883), .Z(n6676) );
  AOI21_X1 U7679 ( .B1(n7594), .B2(n7597), .A(n7593), .ZN(n7592) );
  INV_X1 U7680 ( .A(n14074), .ZN(n7733) );
  NOR2_X1 U7681 ( .A1(n7728), .A2(n7686), .ZN(n7713) );
  NOR2_X1 U7682 ( .A1(n14065), .A2(n7001), .ZN(n7000) );
  INV_X1 U7683 ( .A(n7707), .ZN(n7001) );
  INV_X1 U7684 ( .A(n14881), .ZN(n9325) );
  XNOR2_X1 U7685 ( .A(n14786), .B(n14481), .ZN(n14446) );
  AND2_X1 U7686 ( .A1(n7479), .A2(n14446), .ZN(n7478) );
  NAND2_X1 U7687 ( .A1(n9739), .A2(n14657), .ZN(n7479) );
  AND3_X2 U7688 ( .A1(n9320), .A2(n9336), .A3(n9319), .ZN(n9332) );
  NAND2_X1 U7689 ( .A1(n8242), .A2(n8241), .ZN(n8256) );
  OAI21_X1 U7690 ( .B1(n8240), .B2(n12290), .A(n8239), .ZN(n8242) );
  INV_X1 U7691 ( .A(n12806), .ZN(n12799) );
  OR2_X1 U7693 ( .A1(n8336), .A2(n8335), .ZN(n8401) );
  INV_X1 U7694 ( .A(n7913), .ZN(n7818) );
  AOI21_X1 U7695 ( .B1(n7538), .B2(n7541), .A(n7536), .ZN(n7535) );
  INV_X1 U7696 ( .A(n14152), .ZN(n7536) );
  AOI21_X1 U7697 ( .B1(n7592), .B2(n7140), .A(n6745), .ZN(n7139) );
  INV_X1 U7698 ( .A(n7594), .ZN(n7140) );
  OR2_X1 U7699 ( .A1(n9233), .A2(n7197), .ZN(n7194) );
  NAND2_X1 U7700 ( .A1(n9232), .A2(n9217), .ZN(n7197) );
  NAND2_X1 U7701 ( .A1(n15210), .A2(n15211), .ZN(n15209) );
  AOI22_X1 U7702 ( .A1(n6669), .A2(n13932), .B1(n9049), .B2(n13658), .ZN(n9037) );
  INV_X1 U7703 ( .A(n9119), .ZN(n7669) );
  INV_X1 U7704 ( .A(n14355), .ZN(n7433) );
  NAND2_X1 U7705 ( .A1(n7421), .A2(n14353), .ZN(n7426) );
  NAND2_X1 U7706 ( .A1(n7430), .A2(n7427), .ZN(n7423) );
  NAND2_X1 U7707 ( .A1(n7431), .A2(n7433), .ZN(n7430) );
  INV_X1 U7708 ( .A(n7432), .ZN(n7431) );
  OR2_X1 U7709 ( .A1(n9742), .A2(n14619), .ZN(n14211) );
  OR2_X1 U7710 ( .A1(n8945), .A2(n13193), .ZN(n7064) );
  INV_X1 U7711 ( .A(n7887), .ZN(n7221) );
  OR2_X1 U7712 ( .A1(n13095), .A2(n10366), .ZN(n12970) );
  OR2_X1 U7713 ( .A1(n13181), .A2(n13195), .ZN(n12950) );
  OR2_X1 U7714 ( .A1(n13225), .A2(n13207), .ZN(n12939) );
  OR2_X1 U7715 ( .A1(n15698), .A2(n15687), .ZN(n12854) );
  INV_X1 U7716 ( .A(n11681), .ZN(n12848) );
  NAND2_X1 U7717 ( .A1(n8676), .A2(n8675), .ZN(n8677) );
  NAND2_X1 U7718 ( .A1(n7272), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n7271) );
  NAND2_X1 U7719 ( .A1(n10472), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n8606) );
  AOI21_X1 U7720 ( .B1(n9196), .B2(n9195), .A(n9194), .ZN(n6974) );
  NAND2_X1 U7721 ( .A1(n14074), .A2(n14069), .ZN(n7775) );
  AND2_X1 U7722 ( .A1(n8245), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n8262) );
  INV_X1 U7723 ( .A(n13785), .ZN(n7323) );
  INV_X1 U7724 ( .A(n8328), .ZN(n7324) );
  OR2_X1 U7725 ( .A1(n13859), .A2(n13637), .ZN(n7506) );
  AND2_X1 U7726 ( .A1(n7334), .A2(n6903), .ZN(n6902) );
  INV_X1 U7727 ( .A(n12389), .ZN(n6903) );
  INV_X1 U7728 ( .A(n7334), .ZN(n6904) );
  NOR2_X1 U7729 ( .A1(n7963), .A2(n7095), .ZN(n7094) );
  INV_X1 U7730 ( .A(n7945), .ZN(n7095) );
  OR2_X1 U7731 ( .A1(n13778), .A2(n7161), .ZN(n6835) );
  INV_X1 U7732 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n7340) );
  NAND2_X1 U7733 ( .A1(n7552), .A2(n7550), .ZN(n7549) );
  INV_X1 U7734 ( .A(n7555), .ZN(n7550) );
  INV_X1 U7735 ( .A(n12646), .ZN(n12618) );
  AOI21_X1 U7736 ( .B1(n14366), .B2(n14367), .A(n6839), .ZN(n6845) );
  INV_X1 U7737 ( .A(n14365), .ZN(n6839) );
  NAND2_X1 U7738 ( .A1(n11208), .A2(n11189), .ZN(n14222) );
  AOI21_X1 U7739 ( .B1(n14071), .B2(n14407), .A(n9691), .ZN(n14391) );
  INV_X1 U7740 ( .A(n7458), .ZN(n7457) );
  OR2_X1 U7741 ( .A1(n8222), .A2(n8221), .ZN(n8224) );
  OR2_X1 U7742 ( .A1(n8136), .A2(n11515), .ZN(n7021) );
  AND2_X1 U7743 ( .A1(n9318), .A2(n7558), .ZN(n7557) );
  INV_X1 U7744 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n7558) );
  OR2_X1 U7745 ( .A1(n9547), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n9503) );
  XNOR2_X1 U7746 ( .A(n7946), .B(SI_11_), .ZN(n7949) );
  NAND2_X1 U7747 ( .A1(n10433), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n7071) );
  AOI21_X1 U7748 ( .B1(n7373), .B2(n12219), .A(n6756), .ZN(n7371) );
  INV_X1 U7749 ( .A(n6956), .ZN(n6955) );
  AOI21_X1 U7750 ( .B1(n6956), .B2(n6954), .A(n9872), .ZN(n6953) );
  INV_X1 U7751 ( .A(n9869), .ZN(n6954) );
  AND2_X1 U7752 ( .A1(n7365), .A2(n6796), .ZN(n7364) );
  OR2_X1 U7753 ( .A1(n7367), .A2(n7370), .ZN(n7365) );
  AND2_X1 U7754 ( .A1(n12720), .A2(n9865), .ZN(n12748) );
  NAND2_X1 U7755 ( .A1(n9849), .A2(n7358), .ZN(n12758) );
  NOR2_X1 U7756 ( .A1(n12761), .A2(n7359), .ZN(n7358) );
  INV_X1 U7757 ( .A(n9848), .ZN(n7359) );
  NAND2_X1 U7758 ( .A1(n12702), .A2(n12701), .ZN(n9849) );
  AND2_X1 U7759 ( .A1(n12787), .A2(n12717), .ZN(n6956) );
  NAND2_X1 U7760 ( .A1(n11330), .A2(n11331), .ZN(n11846) );
  XNOR2_X1 U7761 ( .A(n11848), .B(n11857), .ZN(n15562) );
  INV_X1 U7762 ( .A(n15016), .ZN(n13060) );
  AOI21_X1 U7763 ( .B1(n13109), .B2(n12839), .A(n12837), .ZN(n8909) );
  NAND2_X1 U7764 ( .A1(n8870), .A2(n8869), .ZN(n8885) );
  INV_X1 U7765 ( .A(n12912), .ZN(n7133) );
  INV_X1 U7766 ( .A(n13278), .ZN(n15697) );
  INV_X1 U7767 ( .A(n8811), .ZN(n12805) );
  OAI21_X1 U7768 ( .B1(n10343), .B2(n10342), .A(n10344), .ZN(n10349) );
  NAND2_X1 U7769 ( .A1(n8836), .A2(n8835), .ZN(n8847) );
  NAND2_X1 U7770 ( .A1(n8822), .A2(n7282), .ZN(n8836) );
  NOR2_X1 U7771 ( .A1(n8833), .A2(n7283), .ZN(n7282) );
  INV_X1 U7772 ( .A(n7255), .ZN(n7254) );
  OAI21_X1 U7773 ( .B1(n8712), .B2(n7256), .A(n8730), .ZN(n7255) );
  INV_X1 U7774 ( .A(n7052), .ZN(n7051) );
  OAI21_X1 U7775 ( .B1(n8627), .B2(n7053), .A(n8640), .ZN(n7052) );
  AOI21_X1 U7776 ( .B1(n8536), .B2(n7046), .A(n7045), .ZN(n7044) );
  INV_X1 U7777 ( .A(n8518), .ZN(n7046) );
  INV_X1 U7778 ( .A(n8538), .ZN(n7045) );
  INV_X1 U7779 ( .A(n8536), .ZN(n7047) );
  NAND2_X1 U7780 ( .A1(n10410), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n8518) );
  NAND2_X1 U7781 ( .A1(n7184), .A2(n9253), .ZN(n7183) );
  NAND2_X1 U7782 ( .A1(n7186), .A2(n7185), .ZN(n7184) );
  NAND2_X1 U7783 ( .A1(n9230), .A2(n7662), .ZN(n7185) );
  NAND2_X1 U7784 ( .A1(n9247), .A2(n9248), .ZN(n7186) );
  AOI21_X1 U7785 ( .B1(n13764), .B2(n8253), .A(n8252), .ZN(n13616) );
  OR2_X1 U7786 ( .A1(n7775), .A2(n7732), .ZN(n7737) );
  AND2_X1 U7787 ( .A1(n7733), .A2(n14069), .ZN(n7774) );
  NOR2_X1 U7788 ( .A1(n13707), .A2(n13706), .ZN(n13708) );
  NAND2_X1 U7789 ( .A1(n13847), .A2(n8159), .ZN(n13821) );
  NAND2_X1 U7790 ( .A1(n7487), .A2(n7485), .ZN(n8113) );
  INV_X1 U7791 ( .A(n7486), .ZN(n7485) );
  OAI21_X1 U7792 ( .B1(n13904), .B2(n7488), .A(n6760), .ZN(n7486) );
  NAND2_X1 U7793 ( .A1(n6944), .A2(n6943), .ZN(n8319) );
  NOR2_X1 U7794 ( .A1(n6947), .A2(n8316), .ZN(n6943) );
  NAND2_X1 U7795 ( .A1(n12210), .A2(n8006), .ZN(n7498) );
  NAND2_X1 U7796 ( .A1(n8301), .A2(n8300), .ZN(n11646) );
  AND2_X1 U7797 ( .A1(n9272), .A2(n11599), .ZN(n7077) );
  AND2_X1 U7798 ( .A1(n8398), .A2(n8397), .ZN(n9224) );
  BUF_X1 U7799 ( .A(n6717), .Z(n8396) );
  INV_X1 U7800 ( .A(n7713), .ZN(n7327) );
  NAND2_X1 U7801 ( .A1(n7730), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7731) );
  INV_X1 U7802 ( .A(n8282), .ZN(n8284) );
  OR2_X1 U7803 ( .A1(n9341), .A2(n9305), .ZN(n9681) );
  NAND2_X1 U7804 ( .A1(n14111), .A2(n14169), .ZN(n12598) );
  AND2_X1 U7805 ( .A1(n9698), .A2(n9697), .ZN(n14392) );
  AND2_X1 U7806 ( .A1(n9688), .A2(n9687), .ZN(n14368) );
  XNOR2_X1 U7807 ( .A(n14393), .B(n14392), .ZN(n14449) );
  INV_X1 U7808 ( .A(n7478), .ZN(n7477) );
  AOI21_X1 U7809 ( .B1(n7478), .B2(n7476), .A(n6757), .ZN(n7475) );
  AND2_X1 U7810 ( .A1(n9663), .A2(n9662), .ZN(n14665) );
  AND2_X1 U7811 ( .A1(n14680), .A2(n7441), .ZN(n14662) );
  NOR2_X1 U7812 ( .A1(n14669), .A2(n7442), .ZN(n7441) );
  INV_X1 U7813 ( .A(n7445), .ZN(n7442) );
  OR2_X1 U7814 ( .A1(n12552), .A2(n15132), .ZN(n14303) );
  NAND2_X1 U7815 ( .A1(n12313), .A2(n9557), .ZN(n15120) );
  BUF_X1 U7816 ( .A(n9371), .Z(n14408) );
  AND2_X1 U7817 ( .A1(n7595), .A2(n9502), .ZN(n7594) );
  NAND2_X1 U7818 ( .A1(n14433), .A2(n7596), .ZN(n7595) );
  INV_X1 U7819 ( .A(n9486), .ZN(n7596) );
  NAND2_X1 U7820 ( .A1(n11805), .A2(n14432), .ZN(n9487) );
  INV_X1 U7821 ( .A(n11911), .ZN(n7464) );
  INV_X2 U7822 ( .A(n10483), .ZN(n9590) );
  INV_X1 U7823 ( .A(n9742), .ZN(n14210) );
  NAND2_X1 U7824 ( .A1(n9213), .A2(n9212), .ZN(n9233) );
  OAI21_X1 U7825 ( .B1(n8259), .B2(n7235), .A(n7233), .ZN(n9213) );
  INV_X1 U7826 ( .A(n9323), .ZN(n9334) );
  OR2_X1 U7827 ( .A1(n9975), .A2(n9920), .ZN(n9937) );
  AOI21_X1 U7828 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(n9925), .A(n9924), .ZN(
        n9932) );
  NOR2_X1 U7829 ( .A1(n9935), .A2(n9934), .ZN(n9924) );
  NAND2_X1 U7830 ( .A1(n8736), .A2(n8735), .ZN(n13266) );
  NAND2_X1 U7831 ( .A1(n7055), .A2(n10377), .ZN(n13075) );
  NOR2_X1 U7832 ( .A1(n10376), .A2(n10375), .ZN(n10377) );
  NAND2_X1 U7833 ( .A1(n7311), .A2(n7313), .ZN(n7310) );
  NAND2_X1 U7834 ( .A1(n8401), .A2(n7303), .ZN(n7308) );
  NOR2_X1 U7835 ( .A1(n7304), .A2(n13896), .ZN(n7303) );
  XNOR2_X1 U7836 ( .A(n9286), .B(n8400), .ZN(n7304) );
  INV_X1 U7837 ( .A(n8409), .ZN(n7314) );
  OR2_X1 U7838 ( .A1(n8272), .A2(n8335), .ZN(n8273) );
  NOR2_X1 U7839 ( .A1(n14914), .A2(n14913), .ZN(n14912) );
  NOR2_X2 U7840 ( .A1(n14912), .A2(n7176), .ZN(n15197) );
  AOI21_X1 U7841 ( .B1(n14914), .B2(n14913), .A(n7177), .ZN(n7176) );
  INV_X1 U7842 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n7177) );
  INV_X1 U7843 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7205) );
  NAND2_X1 U7844 ( .A1(n14225), .A2(n6737), .ZN(n7440) );
  OAI21_X1 U7845 ( .B1(n9038), .B2(n9037), .A(n9036), .ZN(n9045) );
  NAND2_X1 U7846 ( .A1(n9035), .A2(n9034), .ZN(n9036) );
  NAND2_X1 U7847 ( .A1(n11429), .A2(n6669), .ZN(n6986) );
  NAND2_X1 U7848 ( .A1(n13652), .A2(n9226), .ZN(n6987) );
  OAI21_X1 U7849 ( .B1(n7642), .B2(n9061), .A(n7646), .ZN(n9067) );
  NAND2_X1 U7850 ( .A1(n7645), .A2(n7643), .ZN(n9066) );
  NAND2_X1 U7851 ( .A1(n9089), .A2(n6727), .ZN(n6990) );
  NOR2_X1 U7852 ( .A1(n9089), .A2(n6727), .ZN(n6991) );
  INV_X1 U7853 ( .A(n14295), .ZN(n6802) );
  INV_X1 U7854 ( .A(n14305), .ZN(n7412) );
  AND2_X1 U7855 ( .A1(n6999), .A2(n9125), .ZN(n6995) );
  NAND2_X1 U7856 ( .A1(n7666), .A2(n7664), .ZN(n9126) );
  AND2_X1 U7857 ( .A1(n6999), .A2(n6730), .ZN(n6996) );
  INV_X1 U7858 ( .A(n9157), .ZN(n6998) );
  OR2_X1 U7859 ( .A1(n7418), .A2(n14338), .ZN(n7416) );
  OR2_X1 U7860 ( .A1(n7418), .A2(n14339), .ZN(n7417) );
  NOR2_X1 U7861 ( .A1(n14343), .A2(n14342), .ZN(n7418) );
  NAND2_X1 U7862 ( .A1(n14343), .A2(n14342), .ZN(n7419) );
  NOR2_X1 U7863 ( .A1(n7421), .A2(n14353), .ZN(n7432) );
  NAND2_X1 U7864 ( .A1(n9183), .A2(n9182), .ZN(n7651) );
  INV_X1 U7865 ( .A(n9182), .ZN(n7649) );
  INV_X1 U7866 ( .A(n9183), .ZN(n7650) );
  NAND2_X1 U7867 ( .A1(n6705), .A2(n7432), .ZN(n7422) );
  AOI21_X1 U7868 ( .B1(n7429), .B2(n7433), .A(n7428), .ZN(n7427) );
  INV_X1 U7869 ( .A(n7426), .ZN(n7429) );
  INV_X1 U7870 ( .A(n14354), .ZN(n7428) );
  NAND2_X1 U7871 ( .A1(n7278), .A2(n13135), .ZN(n7277) );
  INV_X1 U7872 ( .A(n12968), .ZN(n7278) );
  INV_X1 U7873 ( .A(n9193), .ZN(n6977) );
  INV_X1 U7874 ( .A(P3_IR_REG_8__SCAN_IN), .ZN(n8427) );
  AOI21_X1 U7875 ( .B1(n7458), .B2(n7459), .A(n14433), .ZN(n7456) );
  AOI21_X1 U7876 ( .B1(n7210), .B2(n7212), .A(n7208), .ZN(n7207) );
  INV_X1 U7877 ( .A(n7965), .ZN(n7208) );
  NAND2_X1 U7878 ( .A1(n9790), .A2(n7354), .ZN(n9791) );
  NAND2_X1 U7879 ( .A1(n11514), .A2(n7355), .ZN(n7354) );
  OR2_X1 U7880 ( .A1(n12983), .A2(n9789), .ZN(n9790) );
  NAND2_X1 U7881 ( .A1(n11681), .A2(n7356), .ZN(n7355) );
  INV_X1 U7882 ( .A(n12684), .ZN(n8454) );
  NAND2_X1 U7883 ( .A1(n10914), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n7301) );
  NAND2_X1 U7884 ( .A1(n10980), .A2(n7023), .ZN(n10994) );
  OR2_X1 U7885 ( .A1(n10982), .A2(n10981), .ZN(n7023) );
  NAND2_X1 U7886 ( .A1(n13049), .A2(n6789), .ZN(n13051) );
  INV_X1 U7887 ( .A(n11923), .ZN(n10366) );
  OR2_X1 U7888 ( .A1(n12842), .A2(n12838), .ZN(n7391) );
  NAND2_X1 U7889 ( .A1(n7393), .A2(n7121), .ZN(n7120) );
  NAND2_X1 U7890 ( .A1(n7122), .A2(n13126), .ZN(n7121) );
  AND2_X1 U7891 ( .A1(n12842), .A2(n6723), .ZN(n7039) );
  NAND2_X1 U7892 ( .A1(n13110), .A2(n8955), .ZN(n7040) );
  INV_X1 U7893 ( .A(n13187), .ZN(n7066) );
  OR2_X1 U7894 ( .A1(n13240), .A2(n13248), .ZN(n12930) );
  INV_X1 U7895 ( .A(n7387), .ZN(n7386) );
  OAI21_X1 U7896 ( .B1(n8656), .B2(n7388), .A(n12828), .ZN(n7387) );
  INV_X1 U7897 ( .A(n12903), .ZN(n7388) );
  AND2_X1 U7898 ( .A1(n7628), .A2(n12891), .ZN(n7627) );
  NAND2_X1 U7899 ( .A1(n7629), .A2(n7631), .ZN(n7628) );
  INV_X1 U7900 ( .A(n7632), .ZN(n7629) );
  INV_X1 U7901 ( .A(n7631), .ZN(n7630) );
  NAND2_X1 U7902 ( .A1(n12189), .A2(n11834), .ZN(n7631) );
  NOR2_X1 U7903 ( .A1(P3_IR_REG_12__SCAN_IN), .A2(P3_IR_REG_21__SCAN_IN), .ZN(
        n7400) );
  NAND2_X1 U7904 ( .A1(n8852), .A2(n7281), .ZN(n7280) );
  AND2_X1 U7905 ( .A1(n8432), .A2(n8438), .ZN(n7357) );
  NOR2_X1 U7906 ( .A1(P3_IR_REG_14__SCAN_IN), .A2(P3_IR_REG_16__SCAN_IN), .ZN(
        n8430) );
  INV_X1 U7907 ( .A(n8552), .ZN(n7043) );
  NAND2_X1 U7908 ( .A1(n10468), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n8554) );
  INV_X1 U7909 ( .A(n7579), .ZN(n7578) );
  OAI22_X1 U7910 ( .A1(n7580), .A2(n6701), .B1(n13532), .B2(n13533), .ZN(n7579) );
  INV_X1 U7911 ( .A(n13553), .ZN(n6936) );
  AND2_X1 U7912 ( .A1(n7578), .A2(n6942), .ZN(n6940) );
  INV_X1 U7913 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n8074) );
  NAND2_X1 U7914 ( .A1(n7162), .A2(n14041), .ZN(n7161) );
  INV_X1 U7915 ( .A(n7163), .ZN(n7162) );
  NAND2_X1 U7916 ( .A1(n7165), .A2(n7164), .ZN(n7163) );
  AND2_X1 U7917 ( .A1(n6709), .A2(n7506), .ZN(n7085) );
  NOR2_X1 U7918 ( .A1(n13861), .A2(n7087), .ZN(n7086) );
  INV_X1 U7919 ( .A(n8134), .ZN(n7087) );
  INV_X1 U7920 ( .A(n8305), .ZN(n7339) );
  NOR2_X1 U7921 ( .A1(n8304), .A2(n6897), .ZN(n6896) );
  INV_X1 U7922 ( .A(n8303), .ZN(n6897) );
  AND2_X1 U7923 ( .A1(n11893), .A2(n7928), .ZN(n9275) );
  INV_X1 U7924 ( .A(n8295), .ZN(n7330) );
  INV_X1 U7925 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n8283) );
  INV_X1 U7926 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n7572) );
  INV_X1 U7927 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n7302) );
  AND2_X1 U7928 ( .A1(n12610), .A2(n12609), .ZN(n12612) );
  OR2_X1 U7929 ( .A1(n14690), .A2(n12645), .ZN(n12610) );
  INV_X1 U7930 ( .A(n12348), .ZN(n7530) );
  INV_X1 U7931 ( .A(n7529), .ZN(n7528) );
  OAI21_X1 U7932 ( .B1(n12168), .B2(n12345), .A(n12348), .ZN(n7529) );
  INV_X1 U7933 ( .A(n11926), .ZN(n7516) );
  NOR2_X1 U7934 ( .A1(n7014), .A2(n7587), .ZN(n7013) );
  INV_X1 U7935 ( .A(n14657), .ZN(n7014) );
  INV_X1 U7936 ( .A(n9627), .ZN(n7151) );
  INV_X1 U7937 ( .A(n14709), .ZN(n9640) );
  NAND2_X1 U7938 ( .A1(n14442), .A2(n7449), .ZN(n7448) );
  INV_X1 U7939 ( .A(n7454), .ZN(n7449) );
  AND2_X1 U7940 ( .A1(n14747), .A2(n14331), .ZN(n7451) );
  INV_X1 U7941 ( .A(n9713), .ZN(n7154) );
  XNOR2_X1 U7942 ( .A(n14845), .B(n14761), .ZN(n12509) );
  INV_X1 U7943 ( .A(n15130), .ZN(n7483) );
  INV_X1 U7944 ( .A(n6807), .ZN(n11103) );
  NAND2_X1 U7945 ( .A1(n11099), .A2(n11103), .ZN(n11101) );
  NAND2_X1 U7946 ( .A1(n11203), .A2(n14224), .ZN(n11102) );
  NAND2_X1 U7947 ( .A1(n14210), .A2(n14387), .ZN(n14412) );
  INV_X1 U7948 ( .A(n14387), .ZN(n14213) );
  INV_X1 U7949 ( .A(n14619), .ZN(n14209) );
  NOR2_X1 U7950 ( .A1(n8391), .A2(n7237), .ZN(n7236) );
  INV_X1 U7951 ( .A(n8258), .ZN(n7237) );
  INV_X1 U7952 ( .A(n8203), .ZN(n7223) );
  NAND2_X1 U7953 ( .A1(n7213), .A2(n7930), .ZN(n7212) );
  INV_X1 U7954 ( .A(n7949), .ZN(n7213) );
  NAND2_X1 U7955 ( .A1(n7908), .A2(SI_10_), .ZN(n7930) );
  NOR2_X1 U7956 ( .A1(n7221), .A2(n7218), .ZN(n7217) );
  INV_X1 U7957 ( .A(n7867), .ZN(n7218) );
  OAI21_X1 U7958 ( .B1(n7871), .B2(n7221), .A(n7905), .ZN(n7220) );
  INV_X2 U7959 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n10191) );
  OAI21_X1 U7960 ( .B1(n10433), .B2(n10441), .A(n7009), .ZN(n7008) );
  NAND2_X1 U7961 ( .A1(n10433), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n7009) );
  NAND2_X1 U7962 ( .A1(n7008), .A2(SI_3_), .ZN(n7783) );
  NAND2_X1 U7963 ( .A1(n9901), .A2(P3_ADDR_REG_2__SCAN_IN), .ZN(n7224) );
  XNOR2_X1 U7964 ( .A(n9907), .B(P3_ADDR_REG_5__SCAN_IN), .ZN(n9942) );
  AND2_X1 U7965 ( .A1(n9911), .A2(P3_ADDR_REG_6__SCAN_IN), .ZN(n6827) );
  AOI21_X1 U7966 ( .B1(P3_ADDR_REG_8__SCAN_IN), .B2(n14574), .A(n9916), .ZN(
        n9939) );
  NOR2_X1 U7967 ( .A1(n9941), .A2(n9940), .ZN(n9916) );
  NAND2_X1 U7968 ( .A1(n11820), .A2(n6965), .ZN(n11817) );
  INV_X1 U7969 ( .A(n11815), .ZN(n6965) );
  AND2_X1 U7970 ( .A1(n6766), .A2(n9812), .ZN(n7353) );
  NAND2_X1 U7971 ( .A1(n11651), .A2(n11652), .ZN(n9813) );
  NAND2_X1 U7972 ( .A1(n15696), .A2(n12850), .ZN(n9799) );
  NAND2_X1 U7973 ( .A1(n7343), .A2(n11238), .ZN(n11534) );
  NOR2_X1 U7974 ( .A1(n11537), .A2(n6853), .ZN(n7343) );
  NOR2_X1 U7975 ( .A1(n9835), .A2(n15042), .ZN(n7374) );
  INV_X1 U7976 ( .A(n12218), .ZN(n7377) );
  OR2_X1 U7977 ( .A1(n9857), .A2(n9856), .ZN(n9860) );
  OR2_X1 U7978 ( .A1(n12769), .A2(n13159), .ZN(n12767) );
  INV_X1 U7979 ( .A(n15042), .ZN(n12180) );
  NAND2_X1 U7980 ( .A1(n7368), .A2(n6736), .ZN(n7367) );
  NAND2_X1 U7981 ( .A1(n7369), .A2(n12331), .ZN(n7368) );
  INV_X1 U7982 ( .A(n7371), .ZN(n7369) );
  NAND2_X1 U7983 ( .A1(n7247), .A2(n12981), .ZN(n7246) );
  XNOR2_X1 U7984 ( .A(n7241), .B(n7356), .ZN(n7240) );
  NOR2_X1 U7985 ( .A1(n12836), .A2(n12835), .ZN(n7242) );
  INV_X1 U7986 ( .A(n8737), .ZN(n10356) );
  NAND2_X1 U7987 ( .A1(n12684), .A2(n13437), .ZN(n8480) );
  XNOR2_X1 U7988 ( .A(n10994), .B(n7022), .ZN(n10983) );
  NAND2_X1 U7989 ( .A1(n10983), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n10996) );
  OAI21_X1 U7990 ( .B1(n11323), .B2(n7295), .A(n7294), .ZN(n11842) );
  NAND2_X1 U7991 ( .A1(n11840), .A2(n7297), .ZN(n7294) );
  OR2_X1 U7992 ( .A1(n11322), .A2(n7296), .ZN(n7295) );
  INV_X1 U7993 ( .A(n7297), .ZN(n7296) );
  NAND2_X1 U7994 ( .A1(n11846), .A2(n11847), .ZN(n11848) );
  INV_X1 U7995 ( .A(n13011), .ZN(n13050) );
  AND2_X1 U7996 ( .A1(n13011), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n6823) );
  XNOR2_X1 U7997 ( .A(n13051), .B(n13015), .ZN(n15570) );
  NOR2_X1 U7998 ( .A1(n13015), .A2(n12997), .ZN(n12998) );
  NOR2_X1 U7999 ( .A1(n15583), .A2(n6820), .ZN(n13000) );
  NOR2_X1 U8000 ( .A1(n13048), .A2(n12375), .ZN(n6820) );
  OR2_X1 U8001 ( .A1(n15616), .A2(n6797), .ZN(n7293) );
  OR2_X1 U8002 ( .A1(n14984), .A2(n7287), .ZN(n7286) );
  NOR2_X1 U8003 ( .A1(n14990), .A2(n13004), .ZN(n7287) );
  INV_X1 U8004 ( .A(n13112), .ZN(n13091) );
  AND2_X1 U8005 ( .A1(n7040), .A2(n6723), .ZN(n8956) );
  NAND2_X1 U8006 ( .A1(n7040), .A2(n7039), .ZN(n10361) );
  INV_X1 U8007 ( .A(n8858), .ZN(n8857) );
  OAI21_X1 U8008 ( .B1(n8947), .B2(n7636), .A(n8952), .ZN(n7070) );
  INV_X1 U8009 ( .A(n8942), .ZN(n7636) );
  AND2_X1 U8010 ( .A1(n12950), .A2(n12955), .ZN(n13175) );
  NAND2_X1 U8011 ( .A1(n7067), .A2(n13196), .ZN(n13190) );
  INV_X1 U8012 ( .A(n13188), .ZN(n7067) );
  OAI21_X1 U8013 ( .B1(n13209), .B2(n13204), .A(n12944), .ZN(n13197) );
  OR2_X1 U8014 ( .A1(n13215), .A2(n13224), .ZN(n13216) );
  NAND2_X1 U8015 ( .A1(n13347), .A2(n12930), .ZN(n13223) );
  INV_X1 U8016 ( .A(n13219), .ZN(n13248) );
  AOI21_X1 U8017 ( .B1(n13258), .B2(n8939), .A(n7690), .ZN(n13246) );
  INV_X1 U8018 ( .A(n12917), .ZN(n7398) );
  NAND2_X1 U8019 ( .A1(n7622), .A2(n8934), .ZN(n7621) );
  NAND2_X1 U8020 ( .A1(n8933), .A2(n8932), .ZN(n12359) );
  NAND2_X1 U8021 ( .A1(n12359), .A2(n12362), .ZN(n12358) );
  NAND2_X1 U8022 ( .A1(n8657), .A2(n8656), .ZN(n15050) );
  AND2_X1 U8023 ( .A1(n12907), .A2(n12906), .ZN(n12828) );
  INV_X1 U8024 ( .A(n15645), .ZN(n8636) );
  NAND2_X1 U8025 ( .A1(n12896), .A2(n12895), .ZN(n15645) );
  AND2_X1 U8026 ( .A1(n8559), .A2(n8924), .ZN(n7638) );
  NAND2_X1 U8027 ( .A1(n11373), .A2(n12864), .ZN(n7381) );
  AOI21_X1 U8028 ( .B1(n12857), .B2(n15677), .A(n8921), .ZN(n11374) );
  AND2_X1 U8029 ( .A1(n12963), .A2(n8967), .ZN(n15700) );
  NAND2_X1 U8030 ( .A1(n12963), .A2(n8966), .ZN(n13278) );
  NAND2_X1 U8031 ( .A1(n8813), .A2(n8812), .ZN(n12708) );
  OR2_X1 U8032 ( .A1(n11545), .A2(n8811), .ZN(n8813) );
  AND2_X1 U8033 ( .A1(n13426), .A2(n10408), .ZN(n10907) );
  AND2_X1 U8034 ( .A1(n9879), .A2(n12963), .ZN(n9881) );
  AND2_X1 U8035 ( .A1(n8984), .A2(n8986), .ZN(n10623) );
  AND2_X1 U8036 ( .A1(n12689), .A2(n12688), .ZN(n12692) );
  OR2_X1 U8037 ( .A1(n12687), .A2(n12686), .ZN(n12689) );
  OR2_X1 U8038 ( .A1(n8451), .A2(n8680), .ZN(n7637) );
  NAND3_X1 U8039 ( .A1(n8443), .A2(n6707), .A3(n8444), .ZN(n8445) );
  INV_X1 U8040 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n8459) );
  INV_X1 U8041 ( .A(n7634), .ZN(n7130) );
  AND2_X1 U8042 ( .A1(n7395), .A2(n8462), .ZN(n7131) );
  INV_X1 U8043 ( .A(n8445), .ZN(n6963) );
  NAND2_X1 U8044 ( .A1(n8896), .A2(n8895), .ZN(n10343) );
  OR2_X1 U8045 ( .A1(n8893), .A2(n8892), .ZN(n8896) );
  NAND2_X1 U8046 ( .A1(n7280), .A2(n8864), .ZN(n8879) );
  OR2_X1 U8047 ( .A1(n8851), .A2(n12327), .ZN(n8864) );
  OR2_X1 U8048 ( .A1(n8910), .A2(P3_IR_REG_21__SCAN_IN), .ZN(n8970) );
  NAND2_X1 U8049 ( .A1(n7284), .A2(n8806), .ZN(n8822) );
  AND2_X1 U8050 ( .A1(n8805), .A2(n7285), .ZN(n7284) );
  XNOR2_X1 U8051 ( .A(n8804), .B(n12138), .ZN(n8803) );
  INV_X1 U8052 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n8438) );
  INV_X1 U8053 ( .A(n8770), .ZN(n8433) );
  INV_X1 U8054 ( .A(n7261), .ZN(n7260) );
  OAI21_X1 U8055 ( .B1(n8767), .B2(n7262), .A(n8783), .ZN(n7261) );
  INV_X1 U8056 ( .A(n8780), .ZN(n7262) );
  NAND2_X1 U8057 ( .A1(n8765), .A2(n8764), .ZN(n8768) );
  NAND2_X1 U8058 ( .A1(n8763), .A2(n8762), .ZN(n8765) );
  NAND2_X1 U8059 ( .A1(n8768), .A2(n8767), .ZN(n8781) );
  NAND2_X1 U8060 ( .A1(n8698), .A2(n8444), .ZN(n8770) );
  INV_X1 U8061 ( .A(n8727), .ZN(n7256) );
  AND2_X1 U8062 ( .A1(n8727), .A2(n8711), .ZN(n8712) );
  NAND2_X1 U8063 ( .A1(n8710), .A2(n8709), .ZN(n8713) );
  NAND2_X1 U8064 ( .A1(n8713), .A2(n8712), .ZN(n8728) );
  NAND2_X1 U8065 ( .A1(n8695), .A2(n8694), .ZN(n8710) );
  NAND2_X1 U8066 ( .A1(n7273), .A2(P2_DATAO_REG_13__SCAN_IN), .ZN(n7272) );
  NAND2_X1 U8067 ( .A1(n8677), .A2(n10838), .ZN(n7274) );
  INV_X1 U8068 ( .A(n7271), .ZN(n7270) );
  AND2_X1 U8069 ( .A1(n8658), .A2(n8639), .ZN(n8640) );
  INV_X1 U8070 ( .A(n8637), .ZN(n7053) );
  AND2_X1 U8071 ( .A1(n8637), .A2(n8626), .ZN(n8627) );
  NAND2_X1 U8072 ( .A1(n8628), .A2(n8627), .ZN(n8638) );
  NAND2_X1 U8073 ( .A1(n8625), .A2(n8624), .ZN(n8628) );
  OAI21_X1 U8074 ( .B1(n8571), .B2(n7060), .A(n7057), .ZN(n8610) );
  AOI21_X1 U8075 ( .B1(n7061), .B2(n7059), .A(n7058), .ZN(n7057) );
  INV_X1 U8076 ( .A(n7061), .ZN(n7060) );
  INV_X1 U8077 ( .A(n8570), .ZN(n7059) );
  NAND2_X1 U8078 ( .A1(n8610), .A2(n8609), .ZN(n8625) );
  NAND2_X1 U8079 ( .A1(n10461), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n8587) );
  AND2_X1 U8080 ( .A1(n8606), .A2(n8589), .ZN(n8590) );
  NAND2_X1 U8081 ( .A1(n8588), .A2(n8587), .ZN(n8591) );
  AND2_X1 U8082 ( .A1(n7269), .A2(n8590), .ZN(n7268) );
  NAND2_X1 U8083 ( .A1(n8574), .A2(n8587), .ZN(n7269) );
  OR2_X1 U8084 ( .A1(n8575), .A2(n8574), .ZN(n8588) );
  NAND2_X1 U8085 ( .A1(n7063), .A2(n8572), .ZN(n8575) );
  NAND2_X1 U8086 ( .A1(n8571), .A2(n8570), .ZN(n7063) );
  AND2_X1 U8087 ( .A1(n8538), .A2(n8520), .ZN(n8536) );
  AND2_X1 U8088 ( .A1(n8518), .A2(n8505), .ZN(n8516) );
  OR2_X1 U8089 ( .A1(n7860), .A2(n7859), .ZN(n7879) );
  NAND2_X1 U8090 ( .A1(n12246), .A2(n7561), .ZN(n12305) );
  NOR2_X1 U8091 ( .A1(n12249), .A2(n7562), .ZN(n7561) );
  INV_X1 U8092 ( .A(n12245), .ZN(n7562) );
  NAND2_X1 U8093 ( .A1(n6937), .A2(n6934), .ZN(n6933) );
  NAND2_X1 U8094 ( .A1(n6940), .A2(n6936), .ZN(n6934) );
  OAI21_X1 U8095 ( .B1(n7578), .B2(n13539), .A(n6938), .ZN(n6937) );
  NAND2_X1 U8096 ( .A1(n7578), .A2(n6939), .ZN(n6938) );
  NOR2_X1 U8097 ( .A1(n6941), .A2(n6936), .ZN(n6935) );
  OR2_X1 U8098 ( .A1(n7580), .A2(n6942), .ZN(n6941) );
  INV_X1 U8099 ( .A(n6933), .ZN(n6931) );
  INV_X1 U8100 ( .A(n6940), .ZN(n6932) );
  NAND2_X1 U8101 ( .A1(n6910), .A2(n11500), .ZN(n6909) );
  INV_X1 U8102 ( .A(n7586), .ZN(n6910) );
  INV_X1 U8103 ( .A(n13599), .ZN(n13454) );
  OR2_X1 U8104 ( .A1(n12469), .A2(n12470), .ZN(n13442) );
  INV_X1 U8105 ( .A(n8169), .ZN(n8167) );
  NAND2_X1 U8106 ( .A1(n13522), .A2(n13521), .ZN(n13520) );
  OR2_X1 U8107 ( .A1(n8105), .A2(n8104), .ZN(n8128) );
  INV_X1 U8108 ( .A(n11881), .ZN(n7577) );
  OR2_X1 U8109 ( .A1(n12081), .A2(n7576), .ZN(n7575) );
  INV_X1 U8110 ( .A(n12066), .ZN(n7576) );
  NAND2_X1 U8111 ( .A1(n12470), .A2(n13441), .ZN(n6894) );
  INV_X1 U8112 ( .A(n13449), .ZN(n6890) );
  OR2_X1 U8113 ( .A1(n8228), .A2(n13620), .ZN(n8247) );
  NOR2_X1 U8114 ( .A1(n7679), .A2(n7680), .ZN(n9254) );
  NOR3_X1 U8115 ( .A1(n14025), .A2(n9049), .A3(n13725), .ZN(n7679) );
  AND2_X1 U8116 ( .A1(n9247), .A2(n9229), .ZN(n9230) );
  NAND2_X1 U8117 ( .A1(n9252), .A2(n9251), .ZN(n9253) );
  INV_X1 U8118 ( .A(n9249), .ZN(n9252) );
  NAND2_X1 U8119 ( .A1(n9205), .A2(n9206), .ZN(n7663) );
  AND2_X1 U8120 ( .A1(n8343), .A2(n8342), .ZN(n9225) );
  AND2_X1 U8121 ( .A1(n8219), .A2(n8218), .ZN(n13486) );
  OR2_X1 U8122 ( .A1(n7775), .A2(n7747), .ZN(n7749) );
  OR2_X1 U8123 ( .A1(n7775), .A2(n7752), .ZN(n7754) );
  INV_X1 U8124 ( .A(n13723), .ZN(n13732) );
  NAND2_X1 U8125 ( .A1(n13947), .A2(n8254), .ZN(n8272) );
  NAND2_X1 U8126 ( .A1(n13771), .A2(n8236), .ZN(n8238) );
  NOR2_X1 U8127 ( .A1(n13841), .A2(n7161), .ZN(n13792) );
  NOR2_X1 U8128 ( .A1(n13841), .A2(n7163), .ZN(n13812) );
  AND2_X1 U8129 ( .A1(n6918), .A2(n7320), .ZN(n6919) );
  AOI21_X1 U8130 ( .B1(n7322), .B2(n13809), .A(n7321), .ZN(n7320) );
  AND2_X1 U8131 ( .A1(n13809), .A2(n8178), .ZN(n7503) );
  NAND2_X1 U8132 ( .A1(n13827), .A2(n8328), .ZN(n13803) );
  NAND2_X1 U8133 ( .A1(n13803), .A2(n13804), .ZN(n13802) );
  AND2_X1 U8134 ( .A1(n8328), .A2(n8177), .ZN(n13828) );
  OR2_X1 U8135 ( .A1(n13821), .A2(n13828), .ZN(n13819) );
  NAND2_X1 U8136 ( .A1(n7315), .A2(n7317), .ZN(n13836) );
  AOI21_X1 U8137 ( .B1(n13861), .B2(n7318), .A(n6741), .ZN(n7317) );
  INV_X1 U8138 ( .A(n8327), .ZN(n7318) );
  OR2_X1 U8139 ( .A1(n13848), .A2(n13836), .ZN(n13838) );
  NAND2_X1 U8140 ( .A1(n13872), .A2(n8327), .ZN(n13862) );
  NAND2_X1 U8141 ( .A1(n13873), .A2(n13874), .ZN(n13872) );
  NAND2_X1 U8142 ( .A1(n8068), .A2(n8067), .ZN(n13909) );
  OR2_X1 U8143 ( .A1(n13909), .A2(n13908), .ZN(n13911) );
  AND2_X1 U8144 ( .A1(n6724), .A2(n8321), .ZN(n7334) );
  NAND2_X1 U8145 ( .A1(n12388), .A2(n12389), .ZN(n8322) );
  NAND2_X1 U8146 ( .A1(n7498), .A2(n7496), .ZN(n7495) );
  NOR2_X1 U8147 ( .A1(n12268), .A2(n7497), .ZN(n7496) );
  INV_X1 U8148 ( .A(n8007), .ZN(n7497) );
  NAND2_X1 U8149 ( .A1(n7495), .A2(n7493), .ZN(n12385) );
  NOR2_X1 U8150 ( .A1(n12389), .A2(n7494), .ZN(n7493) );
  INV_X1 U8151 ( .A(n8024), .ZN(n7494) );
  OR2_X1 U8152 ( .A1(n8311), .A2(n6764), .ZN(n6944) );
  NAND2_X1 U8153 ( .A1(n7090), .A2(n12090), .ZN(n7987) );
  NOR2_X1 U8154 ( .A1(n8312), .A2(n6950), .ZN(n6949) );
  INV_X1 U8155 ( .A(n8310), .ZN(n6950) );
  AOI21_X1 U8156 ( .B1(n7096), .B2(n7094), .A(n7093), .ZN(n7090) );
  NAND2_X1 U8157 ( .A1(n11897), .A2(n8308), .ZN(n11964) );
  NAND2_X1 U8158 ( .A1(n11770), .A2(n7929), .ZN(n11891) );
  NAND2_X1 U8159 ( .A1(n8306), .A2(n7338), .ZN(n11895) );
  NAND2_X1 U8160 ( .A1(n6898), .A2(n6896), .ZN(n8306) );
  NAND2_X1 U8161 ( .A1(n11641), .A2(n7886), .ZN(n11607) );
  NAND2_X1 U8162 ( .A1(n11646), .A2(n11645), .ZN(n6898) );
  NAND2_X1 U8163 ( .A1(n8297), .A2(n8296), .ZN(n11600) );
  NAND2_X1 U8164 ( .A1(n11599), .A2(n7082), .ZN(n7081) );
  INV_X1 U8165 ( .A(n7846), .ZN(n7082) );
  NAND2_X1 U8166 ( .A1(n7505), .A2(n15476), .ZN(n7504) );
  INV_X1 U8167 ( .A(n10858), .ZN(n7075) );
  NAND2_X1 U8168 ( .A1(n8139), .A2(n8138), .ZN(n13859) );
  NAND2_X1 U8169 ( .A1(n8355), .A2(n8354), .ZN(n8361) );
  INV_X1 U8170 ( .A(n8274), .ZN(n7700) );
  AND2_X1 U8171 ( .A1(n14151), .A2(n12607), .ZN(n14096) );
  AND2_X1 U8172 ( .A1(n14087), .A2(n7545), .ZN(n7544) );
  OR2_X1 U8173 ( .A1(n14189), .A2(n12634), .ZN(n7545) );
  NOR2_X1 U8174 ( .A1(n11711), .A2(n7685), .ZN(n11736) );
  AOI21_X1 U8175 ( .B1(n7547), .B2(n7551), .A(n6748), .ZN(n7104) );
  NAND2_X1 U8176 ( .A1(n9300), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9607) );
  INV_X1 U8177 ( .A(n9597), .ZN(n9300) );
  INV_X1 U8178 ( .A(n12586), .ZN(n7546) );
  AOI21_X1 U8179 ( .B1(n7104), .B2(n7548), .A(n7102), .ZN(n7101) );
  INV_X1 U8180 ( .A(n14161), .ZN(n7102) );
  INV_X1 U8181 ( .A(n7104), .ZN(n7103) );
  AND2_X1 U8182 ( .A1(n14095), .A2(n12597), .ZN(n14171) );
  NOR2_X1 U8183 ( .A1(n6828), .A2(n14454), .ZN(n14450) );
  NOR2_X1 U8184 ( .A1(n14449), .A2(n6830), .ZN(n6829) );
  AND2_X1 U8185 ( .A1(n9639), .A2(n9638), .ZN(n14344) );
  INV_X1 U8186 ( .A(n6841), .ZN(n14380) );
  NAND4_X1 U8187 ( .A1(n9364), .A2(n9365), .A3(n9367), .A4(n9366), .ZN(n14503)
         );
  INV_X1 U8188 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9900) );
  NAND2_X1 U8189 ( .A1(n14410), .A2(n14409), .ZN(n14462) );
  NAND2_X1 U8190 ( .A1(n6814), .A2(n6813), .ZN(n12525) );
  NAND2_X1 U8191 ( .A1(n7158), .A2(n14446), .ZN(n6814) );
  NAND2_X1 U8192 ( .A1(n14647), .A2(n7589), .ZN(n7158) );
  AND2_X1 U8193 ( .A1(n9681), .A2(n9306), .ZN(n14088) );
  NAND2_X1 U8194 ( .A1(n7474), .A2(n7478), .ZN(n12523) );
  NAND2_X1 U8195 ( .A1(n12525), .A2(n15317), .ZN(n6857) );
  NOR2_X1 U8196 ( .A1(n14658), .A2(n14657), .ZN(n12521) );
  NAND2_X1 U8197 ( .A1(n14648), .A2(n14657), .ZN(n14647) );
  NAND2_X1 U8198 ( .A1(n14797), .A2(n7682), .ZN(n14648) );
  OR2_X1 U8199 ( .A1(n14801), .A2(n14191), .ZN(n7682) );
  NOR2_X2 U8200 ( .A1(n14685), .A2(n14674), .ZN(n14668) );
  OR2_X1 U8201 ( .A1(n14806), .A2(n14665), .ZN(n7445) );
  NAND2_X1 U8202 ( .A1(n14814), .A2(n7615), .ZN(n14682) );
  AND2_X1 U8203 ( .A1(n14683), .A2(n9652), .ZN(n7615) );
  OR2_X1 U8204 ( .A1(n14693), .A2(n7443), .ZN(n14680) );
  NAND2_X1 U8205 ( .A1(n9738), .A2(n7444), .ZN(n7443) );
  INV_X1 U8206 ( .A(n9737), .ZN(n7444) );
  XNOR2_X1 U8207 ( .A(n14820), .B(n14344), .ZN(n14709) );
  INV_X1 U8208 ( .A(n9615), .ZN(n7603) );
  NAND2_X1 U8209 ( .A1(n7610), .A2(n9615), .ZN(n7604) );
  NAND2_X1 U8210 ( .A1(n14728), .A2(n14727), .ZN(n14726) );
  NAND2_X1 U8211 ( .A1(n14746), .A2(n14763), .ZN(n7454) );
  INV_X1 U8212 ( .A(n14442), .ZN(n14727) );
  OR2_X1 U8213 ( .A1(n14758), .A2(n14488), .ZN(n7609) );
  NOR2_X1 U8214 ( .A1(n14747), .A2(n7606), .ZN(n7605) );
  INV_X1 U8215 ( .A(n7609), .ZN(n7606) );
  NAND2_X1 U8216 ( .A1(n7608), .A2(n7610), .ZN(n7607) );
  INV_X1 U8217 ( .A(n14756), .ZN(n7608) );
  NAND2_X1 U8218 ( .A1(n7446), .A2(n7451), .ZN(n14737) );
  NOR2_X1 U8219 ( .A1(n9588), .A2(n7157), .ZN(n7156) );
  INV_X1 U8220 ( .A(n9571), .ZN(n7157) );
  NAND2_X1 U8221 ( .A1(n15120), .A2(n15130), .ZN(n9572) );
  NAND2_X1 U8222 ( .A1(n12322), .A2(n14437), .ZN(n7484) );
  NAND2_X1 U8223 ( .A1(n7484), .A2(n7481), .ZN(n15127) );
  NOR2_X1 U8224 ( .A1(n14437), .A2(n7612), .ZN(n7611) );
  INV_X1 U8225 ( .A(n9544), .ZN(n7612) );
  AOI21_X1 U8226 ( .B1(n7139), .B2(n7141), .A(n14954), .ZN(n7138) );
  INV_X1 U8227 ( .A(n14298), .ZN(n14438) );
  AOI21_X1 U8228 ( .B1(n7469), .B2(n7471), .A(n6742), .ZN(n7467) );
  NOR2_X1 U8229 ( .A1(n9521), .A2(n9520), .ZN(n9537) );
  INV_X1 U8230 ( .A(n7592), .ZN(n7141) );
  NAND2_X1 U8231 ( .A1(n9505), .A2(n9504), .ZN(n14917) );
  NAND2_X1 U8232 ( .A1(n9495), .A2(n9494), .ZN(n14279) );
  NAND2_X1 U8233 ( .A1(n11973), .A2(n15181), .ZN(n14918) );
  NAND2_X1 U8234 ( .A1(n9475), .A2(n9474), .ZN(n11805) );
  NAND2_X1 U8235 ( .A1(n9728), .A2(n9727), .ZN(n11911) );
  AND2_X1 U8236 ( .A1(n9407), .A2(n7144), .ZN(n7142) );
  NOR2_X1 U8237 ( .A1(n7600), .A2(n7145), .ZN(n7144) );
  INV_X1 U8238 ( .A(n9435), .ZN(n7145) );
  NAND2_X1 U8239 ( .A1(n7147), .A2(n9435), .ZN(n7146) );
  OR2_X1 U8240 ( .A1(n14426), .A2(n7599), .ZN(n7147) );
  NOR2_X1 U8241 ( .A1(n14425), .A2(n7600), .ZN(n7599) );
  OAI21_X1 U8242 ( .B1(n11203), .B2(n14224), .A(n11102), .ZN(n11210) );
  NAND2_X1 U8243 ( .A1(n9339), .A2(n9338), .ZN(n14786) );
  NAND2_X1 U8244 ( .A1(n14892), .A2(n10483), .ZN(n14820) );
  INV_X1 U8245 ( .A(n14224), .ZN(n15281) );
  AOI21_X1 U8246 ( .B1(n9231), .B2(n9215), .A(n9217), .ZN(n7200) );
  NOR2_X1 U8247 ( .A1(n9217), .A2(n7196), .ZN(n7195) );
  INV_X1 U8248 ( .A(n9215), .ZN(n7196) );
  AND2_X2 U8249 ( .A1(n9558), .A2(n7135), .ZN(n9320) );
  NOR2_X1 U8250 ( .A1(n9398), .A2(n9314), .ZN(n7135) );
  INV_X1 U8251 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n9313) );
  INV_X1 U8252 ( .A(n7019), .ZN(n7018) );
  AOI21_X1 U8253 ( .B1(n7019), .B2(n7017), .A(n6790), .ZN(n7016) );
  AND2_X1 U8254 ( .A1(n6785), .A2(n8146), .ZN(n7019) );
  AND2_X1 U8255 ( .A1(n6685), .A2(n7113), .ZN(n7112) );
  INV_X1 U8256 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n7113) );
  NAND2_X1 U8257 ( .A1(n7559), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9352) );
  NAND2_X1 U8258 ( .A1(n8008), .A2(n7994), .ZN(n8010) );
  OAI21_X1 U8259 ( .B1(n7785), .B2(SI_4_), .A(n7811), .ZN(n7787) );
  OAI21_X1 U8260 ( .B1(n7008), .B2(SI_3_), .A(n7783), .ZN(n7766) );
  INV_X1 U8261 ( .A(n7764), .ZN(n7763) );
  NAND2_X1 U8262 ( .A1(n6884), .A2(n9376), .ZN(n6883) );
  NAND2_X1 U8263 ( .A1(n6879), .A2(SI_1_), .ZN(n7722) );
  XNOR2_X1 U8264 ( .A(n9942), .B(P1_ADDR_REG_5__SCAN_IN), .ZN(n9958) );
  NOR2_X2 U8265 ( .A1(n14903), .A2(n9964), .ZN(n9967) );
  NAND2_X1 U8266 ( .A1(n14906), .A2(n9971), .ZN(n9973) );
  NOR2_X1 U8267 ( .A1(n9937), .A2(n9936), .ZN(n9921) );
  OAI21_X1 U8268 ( .B1(n12721), .B2(n6955), .A(n6953), .ZN(n9873) );
  AOI21_X1 U8269 ( .B1(n11172), .B2(n11171), .A(n9804), .ZN(n11240) );
  NAND2_X1 U8270 ( .A1(n8787), .A2(n8786), .ZN(n13225) );
  NAND2_X1 U8271 ( .A1(n10347), .A2(n10346), .ZN(n13095) );
  NAND2_X1 U8272 ( .A1(n12758), .A2(n6738), .ZN(n12711) );
  INV_X1 U8273 ( .A(n12709), .ZN(n7360) );
  INV_X1 U8274 ( .A(n10675), .ZN(n13277) );
  OAI21_X1 U8275 ( .B1(n9842), .B2(n9841), .A(n9840), .ZN(n12740) );
  OAI21_X1 U8276 ( .B1(n12732), .B2(n12730), .A(n10675), .ZN(n9840) );
  NOR2_X1 U8277 ( .A1(n12740), .A2(n12741), .ZN(n12739) );
  NAND2_X1 U8278 ( .A1(n8752), .A2(n8751), .ZN(n13251) );
  NAND2_X1 U8279 ( .A1(n11240), .A2(n11239), .ZN(n11238) );
  AOI21_X1 U8280 ( .B1(n10485), .B2(n12805), .A(n8682), .ZN(n12364) );
  NAND2_X1 U8281 ( .A1(n8824), .A2(n8823), .ZN(n13181) );
  INV_X1 U8282 ( .A(n13234), .ZN(n13263) );
  INV_X1 U8283 ( .A(n12788), .ZN(n12777) );
  NAND2_X1 U8284 ( .A1(n7289), .A2(n7027), .ZN(n8499) );
  NAND2_X1 U8285 ( .A1(n8446), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8551) );
  XNOR2_X1 U8286 ( .A(n11842), .B(n11857), .ZN(n15551) );
  NAND2_X1 U8287 ( .A1(n11850), .A2(n11851), .ZN(n13049) );
  NOR2_X1 U8288 ( .A1(n15618), .A2(n15617), .ZN(n15616) );
  XNOR2_X1 U8289 ( .A(n7293), .B(n14974), .ZN(n14968) );
  NOR2_X1 U8290 ( .A1(n14968), .A2(n14969), .ZN(n14967) );
  NOR2_X1 U8291 ( .A1(n14986), .A2(n14985), .ZN(n14984) );
  XNOR2_X1 U8292 ( .A(n7286), .B(n15016), .ZN(n15007) );
  NOR2_X1 U8293 ( .A1(n15007), .A2(n15008), .ZN(n15006) );
  NOR2_X1 U8294 ( .A1(n15034), .A2(n15033), .ZN(n15035) );
  NAND2_X1 U8295 ( .A1(n13141), .A2(n12954), .ZN(n13136) );
  OR2_X1 U8296 ( .A1(n8856), .A2(n10909), .ZN(n13325) );
  AND2_X1 U8297 ( .A1(n13074), .A2(n15739), .ZN(n7054) );
  AND2_X1 U8298 ( .A1(n13106), .A2(n15734), .ZN(n7118) );
  INV_X1 U8299 ( .A(n6908), .ZN(n6905) );
  NAND2_X1 U8300 ( .A1(n6854), .A2(n6912), .ZN(n7858) );
  AND2_X1 U8301 ( .A1(n6915), .A2(n9234), .ZN(n6912) );
  NAND2_X1 U8302 ( .A1(n11501), .A2(n11500), .ZN(n11508) );
  INV_X1 U8303 ( .A(n13766), .ZN(n13948) );
  NAND2_X1 U8304 ( .A1(n8034), .A2(n8033), .ZN(n12475) );
  AND2_X1 U8305 ( .A1(n11272), .A2(n11266), .ZN(n6878) );
  NAND2_X1 U8306 ( .A1(n8149), .A2(n8148), .ZN(n13975) );
  INV_X1 U8307 ( .A(n9029), .ZN(n9256) );
  NAND4_X1 U8308 ( .A1(n7738), .A2(n7737), .A3(n7736), .A4(n7735), .ZN(n13656)
         );
  NOR2_X1 U8309 ( .A1(n13714), .A2(n6863), .ZN(n6862) );
  OR2_X1 U8310 ( .A1(n15453), .A2(n13718), .ZN(n6863) );
  NAND2_X1 U8311 ( .A1(n13715), .A2(n15450), .ZN(n6864) );
  OAI21_X1 U8312 ( .B1(n7194), .B2(n7913), .A(n7191), .ZN(n13729) );
  AOI21_X1 U8313 ( .B1(n9233), .B2(n7189), .A(n7192), .ZN(n7191) );
  NAND2_X1 U8314 ( .A1(n15470), .A2(n11044), .ZN(n13916) );
  AND2_X1 U8315 ( .A1(n13919), .A2(n11390), .ZN(n13933) );
  AND2_X1 U8316 ( .A1(n13741), .A2(n7314), .ZN(n7307) );
  INV_X1 U8317 ( .A(n9224), .ZN(n13744) );
  NAND2_X1 U8318 ( .A1(n6926), .A2(n6925), .ZN(n14030) );
  INV_X1 U8319 ( .A(n13752), .ZN(n6926) );
  NAND2_X1 U8320 ( .A1(n7794), .A2(n7793), .ZN(n11400) );
  INV_X1 U8321 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n7727) );
  AND3_X1 U8322 ( .A1(n9555), .A2(n9554), .A3(n9553), .ZN(n15132) );
  OAI22_X1 U8323 ( .A1(n11197), .A2(n11196), .B1(n11195), .B2(n11194), .ZN(
        n11198) );
  NAND2_X1 U8324 ( .A1(n9564), .A2(n9563), .ZN(n14309) );
  INV_X1 U8325 ( .A(n14323), .ZN(n14845) );
  NAND4_X1 U8326 ( .A1(n9434), .A2(n9433), .A3(n9432), .A4(n9431), .ZN(n14497)
         );
  AOI21_X1 U8327 ( .B1(n10400), .B2(n15125), .A(n10399), .ZN(n10401) );
  AOI21_X1 U8328 ( .B1(n9746), .B2(n15160), .A(n6792), .ZN(n10402) );
  OR2_X1 U8329 ( .A1(n10483), .A2(n14512), .ZN(n7509) );
  NAND2_X1 U8330 ( .A1(n14908), .A2(n14907), .ZN(n14906) );
  XNOR2_X1 U8331 ( .A(n9973), .B(n9972), .ZN(n14911) );
  NAND2_X1 U8332 ( .A1(n6819), .A2(n6818), .ZN(n7182) );
  INV_X1 U8333 ( .A(n15198), .ZN(n6818) );
  NAND2_X1 U8334 ( .A1(n6870), .A2(n6869), .ZN(n7201) );
  INV_X1 U8335 ( .A(n15215), .ZN(n6869) );
  INV_X1 U8336 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n7230) );
  INV_X1 U8337 ( .A(n14237), .ZN(n14238) );
  NAND2_X1 U8338 ( .A1(n9049), .A2(n13656), .ZN(n9041) );
  NAND2_X1 U8339 ( .A1(n11129), .A2(n6669), .ZN(n9042) );
  NAND2_X1 U8340 ( .A1(n11129), .A2(n9049), .ZN(n9039) );
  OR2_X1 U8341 ( .A1(n7437), .A2(n14252), .ZN(n7436) );
  INV_X1 U8342 ( .A(n14251), .ZN(n7437) );
  INV_X1 U8343 ( .A(n7644), .ZN(n7642) );
  NAND2_X1 U8344 ( .A1(n7641), .A2(n7647), .ZN(n7646) );
  INV_X1 U8345 ( .A(n9060), .ZN(n7647) );
  AND2_X1 U8346 ( .A1(n7644), .A2(n9068), .ZN(n7643) );
  NAND2_X1 U8347 ( .A1(n14263), .A2(n14265), .ZN(n7414) );
  NAND2_X1 U8348 ( .A1(n7656), .A2(n6740), .ZN(n6973) );
  NAND2_X1 U8349 ( .A1(n9076), .A2(n6690), .ZN(n7657) );
  NAND2_X1 U8350 ( .A1(n9082), .A2(n9083), .ZN(n6971) );
  NOR2_X1 U8351 ( .A1(n6704), .A2(n6972), .ZN(n6970) );
  NAND2_X1 U8352 ( .A1(n6704), .A2(n6972), .ZN(n6969) );
  OR2_X1 U8353 ( .A1(n7435), .A2(n14277), .ZN(n7434) );
  INV_X1 U8354 ( .A(n14276), .ZN(n7435) );
  AOI21_X1 U8355 ( .B1(n6990), .B2(n6991), .A(n6751), .ZN(n6988) );
  NOR2_X1 U8356 ( .A1(n6730), .A2(n7665), .ZN(n7664) );
  INV_X1 U8357 ( .A(n7667), .ZN(n7665) );
  OR2_X1 U8358 ( .A1(n6711), .A2(n7669), .ZN(n7667) );
  NAND2_X1 U8359 ( .A1(n6711), .A2(n7669), .ZN(n7668) );
  NOR2_X1 U8360 ( .A1(n7410), .A2(n14306), .ZN(n7407) );
  INV_X1 U8361 ( .A(n14315), .ZN(n7410) );
  NAND2_X1 U8362 ( .A1(n14315), .A2(n7409), .ZN(n7408) );
  INV_X1 U8363 ( .A(n7411), .ZN(n7409) );
  AOI21_X1 U8364 ( .B1(n7413), .B2(n14298), .A(n7412), .ZN(n7411) );
  INV_X1 U8365 ( .A(n9162), .ZN(n6992) );
  AOI21_X1 U8366 ( .B1(n7415), .B2(n7420), .A(n6754), .ZN(n14347) );
  OAI21_X1 U8367 ( .B1(n14340), .B2(n7417), .A(n7416), .ZN(n7415) );
  OAI21_X1 U8368 ( .B1(n6978), .B2(n6980), .A(n7648), .ZN(n9188) );
  NAND2_X1 U8369 ( .A1(n7650), .A2(n7649), .ZN(n7648) );
  AOI21_X1 U8370 ( .B1(n6985), .B2(n6984), .A(n6979), .ZN(n6978) );
  NOR2_X1 U8371 ( .A1(n6705), .A2(n7427), .ZN(n7424) );
  NAND2_X1 U8372 ( .A1(n7276), .A2(n7275), .ZN(n12976) );
  NAND2_X1 U8373 ( .A1(n13090), .A2(n12969), .ZN(n7275) );
  INV_X1 U8374 ( .A(n12976), .ZN(n12973) );
  NOR3_X1 U8375 ( .A1(n13086), .A2(n12842), .A3(n13111), .ZN(n12967) );
  NOR2_X1 U8376 ( .A1(n12842), .A2(n12818), .ZN(n7393) );
  NAND2_X1 U8377 ( .A1(n6976), .A2(n6975), .ZN(n9196) );
  NAND2_X1 U8378 ( .A1(n9192), .A2(n9191), .ZN(n6975) );
  CLKBUF_X1 U8379 ( .A(n14421), .Z(n6807) );
  NOR2_X1 U8380 ( .A1(n14233), .A2(n15293), .ZN(n7508) );
  NAND2_X1 U8381 ( .A1(n8047), .A2(n10834), .ZN(n8071) );
  INV_X1 U8382 ( .A(n11820), .ZN(n9815) );
  NAND2_X1 U8383 ( .A1(n7300), .A2(n7299), .ZN(n7298) );
  NOR2_X1 U8384 ( .A1(n10976), .A2(n10975), .ZN(n10977) );
  INV_X1 U8385 ( .A(n6821), .ZN(n11320) );
  OAI21_X1 U8386 ( .B1(n11162), .B2(n11161), .A(n6822), .ZN(n6821) );
  NAND2_X1 U8387 ( .A1(n11163), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n6822) );
  NAND2_X1 U8388 ( .A1(n11853), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n7297) );
  NAND2_X1 U8389 ( .A1(n15585), .A2(n13053), .ZN(n13054) );
  OR2_X1 U8390 ( .A1(n13079), .A2(n13092), .ZN(n12834) );
  NAND2_X1 U8391 ( .A1(n8901), .A2(n8900), .ZN(n8958) );
  INV_X1 U8392 ( .A(n8902), .ZN(n8901) );
  INV_X1 U8393 ( .A(n7123), .ZN(n7122) );
  OAI21_X1 U8394 ( .B1(n13126), .B2(n12954), .A(n12965), .ZN(n7123) );
  OR2_X1 U8395 ( .A1(n8950), .A2(n7065), .ZN(n8951) );
  AND2_X1 U8396 ( .A1(n13173), .A2(n8949), .ZN(n7065) );
  NAND2_X1 U8397 ( .A1(n13232), .A2(n8942), .ZN(n13215) );
  NOR2_X1 U8398 ( .A1(n7623), .A2(n7620), .ZN(n7619) );
  INV_X1 U8399 ( .A(n8932), .ZN(n7620) );
  INV_X1 U8400 ( .A(n8934), .ZN(n7623) );
  NAND2_X1 U8401 ( .A1(n7633), .A2(n12038), .ZN(n7632) );
  INV_X1 U8402 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n11333) );
  OR2_X1 U8403 ( .A1(n11947), .A2(n11797), .ZN(n12878) );
  INV_X1 U8404 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n8527) );
  OR2_X1 U8405 ( .A1(n11673), .A2(n11569), .ZN(n12868) );
  NAND2_X1 U8406 ( .A1(n7126), .A2(n15681), .ZN(n12861) );
  NAND2_X1 U8407 ( .A1(n15679), .A2(n15678), .ZN(n12853) );
  INV_X1 U8408 ( .A(n8821), .ZN(n7283) );
  NAND2_X1 U8409 ( .A1(n7259), .A2(n7257), .ZN(n8804) );
  AOI21_X1 U8410 ( .B1(n7260), .B2(n7262), .A(n7258), .ZN(n7257) );
  INV_X1 U8411 ( .A(n8793), .ZN(n7258) );
  OR2_X1 U8412 ( .A1(n8715), .A2(P3_IR_REG_14__SCAN_IN), .ZN(n8733) );
  NOR2_X1 U8413 ( .A1(n7267), .A2(n7062), .ZN(n7061) );
  INV_X1 U8414 ( .A(n8572), .ZN(n7062) );
  INV_X1 U8415 ( .A(n7268), .ZN(n7267) );
  INV_X1 U8416 ( .A(n7264), .ZN(n7058) );
  AOI21_X1 U8417 ( .B1(n7268), .B2(n7266), .A(n7265), .ZN(n7264) );
  INV_X1 U8418 ( .A(n8606), .ZN(n7265) );
  INV_X1 U8419 ( .A(n8587), .ZN(n7266) );
  OR2_X1 U8420 ( .A1(n6720), .A2(P3_IR_REG_7__SCAN_IN), .ZN(n8604) );
  NAND2_X1 U8421 ( .A1(n7580), .A2(n6942), .ZN(n6939) );
  NAND2_X1 U8422 ( .A1(n7581), .A2(n13497), .ZN(n7580) );
  INV_X1 U8423 ( .A(n13534), .ZN(n7581) );
  INV_X1 U8424 ( .A(n13539), .ZN(n6942) );
  AND2_X1 U8425 ( .A1(n8035), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8056) );
  INV_X1 U8426 ( .A(n13613), .ZN(n7582) );
  NOR2_X1 U8427 ( .A1(n8020), .A2(n8019), .ZN(n8035) );
  OAI22_X1 U8428 ( .A1(n9228), .A2(n9227), .B1(n9205), .B2(n9206), .ZN(n7662)
         );
  OR2_X1 U8429 ( .A1(n7879), .A2(n7878), .ZN(n7896) );
  OAI21_X1 U8430 ( .B1(n13675), .B2(n15400), .A(n15410), .ZN(n13676) );
  INV_X1 U8431 ( .A(n13828), .ZN(n7502) );
  NOR2_X1 U8432 ( .A1(n7319), .A2(n9279), .ZN(n7316) );
  INV_X1 U8433 ( .A(n13861), .ZN(n7319) );
  INV_X1 U8434 ( .A(n8313), .ZN(n6948) );
  INV_X1 U8435 ( .A(n7092), .ZN(n7091) );
  OAI21_X1 U8436 ( .B1(n7094), .B2(n7093), .A(n7172), .ZN(n7092) );
  OR2_X1 U8437 ( .A1(n7896), .A2(n11764), .ZN(n7921) );
  NAND2_X1 U8438 ( .A1(n7920), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n7937) );
  INV_X1 U8439 ( .A(n7921), .ZN(n7920) );
  NAND2_X1 U8440 ( .A1(n13838), .A2(n6921), .ZN(n13827) );
  OR2_X1 U8441 ( .A1(n7819), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n7832) );
  INV_X1 U8442 ( .A(P2_RD_REG_SCAN_IN), .ZN(n6876) );
  INV_X1 U8443 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n6877) );
  INV_X1 U8444 ( .A(P1_RD_REG_SCAN_IN), .ZN(n7715) );
  AOI21_X1 U8445 ( .B1(n14096), .B2(n7540), .A(n7539), .ZN(n7538) );
  INV_X1 U8446 ( .A(n14096), .ZN(n7541) );
  NOR2_X1 U8447 ( .A1(n7556), .A2(n12572), .ZN(n7555) );
  INV_X1 U8448 ( .A(n12565), .ZN(n7556) );
  NOR2_X1 U8449 ( .A1(n7533), .A2(n7111), .ZN(n7110) );
  INV_X1 U8450 ( .A(n12538), .ZN(n7111) );
  INV_X1 U8451 ( .A(n12549), .ZN(n7533) );
  INV_X1 U8452 ( .A(n7531), .ZN(n7107) );
  AOI21_X1 U8453 ( .B1(n12549), .B2(n7532), .A(n6729), .ZN(n7531) );
  INV_X1 U8454 ( .A(n15103), .ZN(n7532) );
  NAND2_X1 U8455 ( .A1(n12487), .A2(n12488), .ZN(n12503) );
  AND2_X1 U8456 ( .A1(n14398), .A2(n14397), .ZN(n14401) );
  AND2_X1 U8457 ( .A1(n14394), .A2(n7405), .ZN(n7404) );
  NAND2_X1 U8458 ( .A1(n14370), .A2(n14371), .ZN(n7405) );
  NAND2_X1 U8459 ( .A1(n14446), .A2(n14445), .ZN(n6830) );
  OR2_X1 U8460 ( .A1(n14369), .A2(n14480), .ZN(n9689) );
  NOR2_X1 U8461 ( .A1(n14446), .A2(n7590), .ZN(n7015) );
  NOR2_X1 U8462 ( .A1(n14786), .A2(n14793), .ZN(n7507) );
  NOR2_X1 U8463 ( .A1(n14711), .A2(n14812), .ZN(n7511) );
  NOR2_X1 U8464 ( .A1(n14757), .A2(n14758), .ZN(n6872) );
  AND2_X1 U8465 ( .A1(n9299), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9565) );
  INV_X1 U8466 ( .A(n9567), .ZN(n9299) );
  INV_X1 U8467 ( .A(n7470), .ZN(n7469) );
  OAI21_X1 U8468 ( .B1(n7593), .B2(n7471), .A(n14954), .ZN(n7470) );
  INV_X1 U8469 ( .A(n9734), .ZN(n7471) );
  INV_X1 U8470 ( .A(n9730), .ZN(n7461) );
  AND3_X1 U8471 ( .A1(n7508), .A2(n11341), .A3(n15303), .ZN(n11450) );
  NAND2_X1 U8472 ( .A1(n14222), .A2(n14214), .ZN(n6838) );
  INV_X1 U8473 ( .A(n7601), .ZN(n14217) );
  NAND2_X1 U8474 ( .A1(n14503), .A2(n10815), .ZN(n7601) );
  INV_X1 U8475 ( .A(n7513), .ZN(n12316) );
  INV_X1 U8476 ( .A(n7234), .ZN(n7233) );
  OAI21_X1 U8477 ( .B1(n7236), .B2(n7235), .A(n9208), .ZN(n7234) );
  INV_X1 U8478 ( .A(n8395), .ZN(n7235) );
  INV_X1 U8479 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n9312) );
  INV_X1 U8480 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n9758) );
  INV_X1 U8481 ( .A(n7021), .ZN(n7017) );
  AND2_X1 U8482 ( .A1(n8045), .A2(n8029), .ZN(n8043) );
  INV_X1 U8483 ( .A(n8009), .ZN(n7206) );
  AND2_X1 U8484 ( .A1(n8025), .A2(n8013), .ZN(n8014) );
  XNOR2_X1 U8485 ( .A(n7967), .B(n10457), .ZN(n7965) );
  INV_X1 U8486 ( .A(n7211), .ZN(n7210) );
  OAI21_X1 U8487 ( .B1(n7910), .B2(n7212), .A(n7948), .ZN(n7211) );
  OAI21_X1 U8488 ( .B1(n7889), .B2(SI_9_), .A(n7907), .ZN(n7904) );
  INV_X1 U8489 ( .A(n7811), .ZN(n7215) );
  INV_X1 U8490 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n10195) );
  NOR2_X1 U8491 ( .A1(n9915), .A2(n9914), .ZN(n9941) );
  NOR2_X1 U8492 ( .A1(n9837), .A2(n7374), .ZN(n7373) );
  INV_X1 U8493 ( .A(n9861), .ZN(n7345) );
  NAND2_X1 U8494 ( .A1(n9813), .A2(n7353), .ZN(n11818) );
  NAND2_X1 U8495 ( .A1(n8814), .A2(n10223), .ZN(n8825) );
  NAND2_X1 U8496 ( .A1(n9862), .A2(n9861), .ZN(n12747) );
  AND2_X1 U8497 ( .A1(n8580), .A2(n11333), .ZN(n8597) );
  INV_X1 U8498 ( .A(n15696), .ZN(n11025) );
  NAND2_X1 U8499 ( .A1(n9847), .A2(n13235), .ZN(n9848) );
  OR2_X1 U8500 ( .A1(n8796), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n8815) );
  NAND2_X1 U8501 ( .A1(n8788), .A2(n10192), .ZN(n8796) );
  INV_X1 U8502 ( .A(n8789), .ZN(n8788) );
  OAI21_X1 U8503 ( .B1(n12046), .B2(n9829), .A(n9828), .ZN(n12177) );
  NAND2_X1 U8504 ( .A1(n8754), .A2(n8753), .ZN(n8774) );
  INV_X1 U8505 ( .A(n8755), .ZN(n8754) );
  OR2_X1 U8506 ( .A1(n8774), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8789) );
  NAND2_X1 U8507 ( .A1(n9813), .A2(n9812), .ZN(n11698) );
  NAND2_X1 U8508 ( .A1(n8720), .A2(n8719), .ZN(n8738) );
  INV_X1 U8509 ( .A(n8721), .ZN(n8720) );
  AND2_X1 U8510 ( .A1(n12331), .A2(n7373), .ZN(n7370) );
  INV_X1 U8511 ( .A(n12982), .ZN(n7244) );
  OAI21_X1 U8512 ( .B1(n7300), .B2(n7299), .A(n7298), .ZN(n10915) );
  NOR2_X1 U8513 ( .A1(n10936), .A2(n10935), .ZN(n10939) );
  INV_X1 U8514 ( .A(n7298), .ZN(n10936) );
  XNOR2_X1 U8515 ( .A(n10977), .B(n7022), .ZN(n10978) );
  NOR2_X1 U8516 ( .A1(n10978), .A2(n8523), .ZN(n11001) );
  NOR2_X1 U8517 ( .A1(n11001), .A2(n7288), .ZN(n11162) );
  NOR2_X1 U8518 ( .A1(n10977), .A2(n7022), .ZN(n7288) );
  NAND2_X1 U8519 ( .A1(n10996), .A2(n10997), .ZN(n10998) );
  NAND2_X1 U8520 ( .A1(n11328), .A2(n11329), .ZN(n11330) );
  NAND2_X1 U8521 ( .A1(n15569), .A2(n13052), .ZN(n15586) );
  NAND2_X1 U8522 ( .A1(n15586), .A2(n15587), .ZN(n15585) );
  XNOR2_X1 U8523 ( .A(n13054), .B(n13020), .ZN(n15602) );
  NAND2_X1 U8524 ( .A1(n7394), .A2(n12970), .ZN(n12798) );
  NOR2_X1 U8525 ( .A1(n12971), .A2(n7390), .ZN(n7389) );
  INV_X1 U8526 ( .A(n7391), .ZN(n7390) );
  NAND2_X1 U8527 ( .A1(n12970), .A2(n10363), .ZN(n13086) );
  INV_X1 U8528 ( .A(n13086), .ZN(n13090) );
  INV_X1 U8529 ( .A(n12673), .ZN(n13092) );
  OAI21_X2 U8530 ( .B1(n13110), .B2(n7038), .A(n7036), .ZN(n13089) );
  AOI21_X1 U8531 ( .B1(n7039), .B2(n7037), .A(n6755), .ZN(n7036) );
  INV_X1 U8532 ( .A(n7039), .ZN(n7038) );
  INV_X1 U8533 ( .A(n8955), .ZN(n7037) );
  OR2_X1 U8534 ( .A1(n12818), .A2(n12837), .ZN(n13111) );
  OR2_X1 U8535 ( .A1(n13325), .A2(n13160), .ZN(n12954) );
  OR2_X1 U8536 ( .A1(n8839), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8858) );
  AND2_X1 U8537 ( .A1(n12843), .A2(n12844), .ZN(n13193) );
  INV_X1 U8538 ( .A(n12939), .ZN(n7399) );
  AND2_X1 U8539 ( .A1(n12939), .A2(n12940), .ZN(n13224) );
  AOI21_X1 U8540 ( .B1(n13250), .B2(n7380), .A(n7379), .ZN(n7378) );
  NAND2_X1 U8541 ( .A1(n13265), .A2(n7129), .ZN(n7128) );
  AND2_X1 U8542 ( .A1(n13264), .A2(n13250), .ZN(n7129) );
  OR2_X1 U8543 ( .A1(n13231), .A2(n12934), .ZN(n13232) );
  AND2_X1 U8544 ( .A1(n12920), .A2(n12924), .ZN(n13280) );
  OR2_X1 U8545 ( .A1(n8703), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8721) );
  NAND2_X1 U8546 ( .A1(n8685), .A2(n8684), .ZN(n8703) );
  INV_X1 U8547 ( .A(n8686), .ZN(n8685) );
  AOI21_X1 U8548 ( .B1(n7386), .B2(n7388), .A(n7385), .ZN(n7384) );
  INV_X1 U8549 ( .A(n12906), .ZN(n7385) );
  NAND2_X1 U8550 ( .A1(n8668), .A2(n12220), .ZN(n8686) );
  INV_X1 U8551 ( .A(n8669), .ZN(n8668) );
  INV_X1 U8552 ( .A(n13292), .ZN(n12373) );
  NAND2_X1 U8553 ( .A1(n12372), .A2(n15051), .ZN(n7639) );
  NOR2_X1 U8554 ( .A1(n12372), .A2(n15051), .ZN(n7640) );
  OR2_X1 U8555 ( .A1(n8648), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8669) );
  AOI21_X1 U8556 ( .B1(n7627), .B2(n7630), .A(n6716), .ZN(n7624) );
  OR2_X1 U8557 ( .A1(n8614), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8648) );
  NAND2_X1 U8558 ( .A1(n8597), .A2(n8596), .ZN(n8614) );
  NAND2_X1 U8559 ( .A1(n7626), .A2(n7631), .ZN(n12188) );
  NAND2_X1 U8560 ( .A1(n12030), .A2(n7632), .ZN(n7626) );
  INV_X1 U8561 ( .A(n12029), .ZN(n12886) );
  NOR2_X1 U8562 ( .A1(n8560), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8580) );
  NAND2_X1 U8563 ( .A1(n12884), .A2(n12883), .ZN(n12819) );
  OR2_X1 U8564 ( .A1(n8545), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8560) );
  NOR2_X1 U8565 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n8526) );
  NAND2_X1 U8566 ( .A1(n12853), .A2(n12854), .ZN(n11370) );
  AND3_X1 U8567 ( .A1(n8477), .A2(n8478), .A3(n8476), .ZN(n15695) );
  NAND2_X1 U8568 ( .A1(n8884), .A2(n8883), .ZN(n13118) );
  INV_X1 U8569 ( .A(n15730), .ZN(n15070) );
  AND2_X1 U8570 ( .A1(n7635), .A2(n6777), .ZN(n6961) );
  NAND2_X1 U8571 ( .A1(n12692), .A2(n12691), .ZN(n12802) );
  OR2_X1 U8572 ( .A1(n10349), .A2(n10348), .ZN(n10352) );
  NAND2_X1 U8573 ( .A1(n8879), .A2(n8878), .ZN(n8881) );
  NOR2_X1 U8574 ( .A1(n8445), .A2(n7634), .ZN(n8973) );
  XNOR2_X1 U8575 ( .A(n8972), .B(n8971), .ZN(n10910) );
  OAI21_X1 U8576 ( .B1(n8970), .B2(P3_IR_REG_22__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8972) );
  XNOR2_X1 U8577 ( .A(n8437), .B(P3_IR_REG_20__SCAN_IN), .ZN(n9015) );
  NAND2_X1 U8578 ( .A1(n7253), .A2(n7251), .ZN(n8763) );
  AOI21_X1 U8579 ( .B1(n7254), .B2(n7256), .A(n7252), .ZN(n7251) );
  INV_X1 U8580 ( .A(n8745), .ZN(n7252) );
  OR2_X1 U8581 ( .A1(n8733), .A2(P3_IR_REG_15__SCAN_IN), .ZN(n8748) );
  NAND2_X1 U8582 ( .A1(n7271), .A2(n7274), .ZN(n8695) );
  AND2_X1 U8583 ( .A1(n8709), .A2(n8693), .ZN(n8694) );
  NOR2_X1 U8584 ( .A1(n6697), .A2(P3_IR_REG_12__SCAN_IN), .ZN(n8698) );
  NAND2_X1 U8585 ( .A1(n7050), .A2(n7048), .ZN(n8662) );
  AOI21_X1 U8586 ( .B1(n7051), .B2(n7053), .A(n7049), .ZN(n7048) );
  NAND2_X1 U8587 ( .A1(n8628), .A2(n7051), .ZN(n7050) );
  INV_X1 U8588 ( .A(n8658), .ZN(n7049) );
  AND2_X1 U8589 ( .A1(n8675), .A2(n8660), .ZN(n8661) );
  NAND2_X1 U8590 ( .A1(n8662), .A2(n8661), .ZN(n8676) );
  NAND2_X1 U8591 ( .A1(n8555), .A2(n8554), .ZN(n8571) );
  AOI21_X1 U8592 ( .B1(n7044), .B2(n7047), .A(n7043), .ZN(n7042) );
  INV_X1 U8593 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n8534) );
  INV_X1 U8594 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n8488) );
  AND2_X1 U8595 ( .A1(n8503), .A2(n8491), .ZN(n8501) );
  AND2_X1 U8596 ( .A1(n8464), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n8486) );
  OR2_X1 U8597 ( .A1(n7979), .A2(n7978), .ZN(n7999) );
  NAND2_X1 U8598 ( .A1(n8151), .A2(n8150), .ZN(n8169) );
  INV_X1 U8599 ( .A(n8152), .ZN(n8151) );
  OR2_X1 U8600 ( .A1(n8128), .A2(n8127), .ZN(n8152) );
  NAND2_X1 U8601 ( .A1(n13491), .A2(n6701), .ZN(n13611) );
  OR2_X1 U8602 ( .A1(n7999), .A2(n12251), .ZN(n8020) );
  INV_X1 U8603 ( .A(n8332), .ZN(n9291) );
  NAND2_X1 U8604 ( .A1(n12137), .A2(n13718), .ZN(n11045) );
  NOR3_X1 U8605 ( .A1(n13661), .A2(n10712), .A3(n13665), .ZN(n13659) );
  AOI21_X1 U8606 ( .B1(n15380), .B2(n10775), .A(n10774), .ZN(n10773) );
  OR2_X1 U8607 ( .A1(n7874), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n7890) );
  OAI21_X1 U8608 ( .B1(n11232), .B2(n11230), .A(n11231), .ZN(n13673) );
  NAND2_X1 U8609 ( .A1(n15437), .A2(n13680), .ZN(n15452) );
  INV_X1 U8610 ( .A(n7195), .ZN(n7190) );
  NAND2_X1 U8611 ( .A1(n9286), .A2(n7312), .ZN(n7311) );
  NAND2_X1 U8612 ( .A1(n8272), .A2(n8335), .ZN(n8390) );
  INV_X1 U8613 ( .A(n9284), .ZN(n8335) );
  AND2_X1 U8614 ( .A1(n8264), .A2(n8248), .ZN(n13764) );
  AOI21_X1 U8615 ( .B1(n6919), .B2(n6920), .A(n6747), .ZN(n6917) );
  OAI21_X1 U8616 ( .B1(n13821), .B2(n7501), .A(n7499), .ZN(n13791) );
  OR2_X1 U8617 ( .A1(n7503), .A2(n7500), .ZN(n7499) );
  NAND2_X1 U8618 ( .A1(n7502), .A2(n8201), .ZN(n7501) );
  INV_X1 U8619 ( .A(n8201), .ZN(n7500) );
  NAND2_X1 U8620 ( .A1(n13791), .A2(n7321), .ZN(n13790) );
  INV_X1 U8621 ( .A(n7506), .ZN(n7084) );
  NAND2_X1 U8622 ( .A1(n6900), .A2(n6899), .ZN(n13894) );
  AOI21_X1 U8623 ( .B1(n6901), .B2(n6904), .A(n6746), .ZN(n6899) );
  NOR2_X1 U8624 ( .A1(n6749), .A2(n6902), .ZN(n6901) );
  OR2_X1 U8625 ( .A1(n13895), .A2(n13894), .ZN(n13898) );
  NAND2_X1 U8626 ( .A1(n7175), .A2(n7174), .ZN(n13914) );
  INV_X1 U8627 ( .A(n14053), .ZN(n7174) );
  NAND2_X1 U8628 ( .A1(n12385), .A2(n8042), .ZN(n12422) );
  AND2_X1 U8629 ( .A1(n10505), .A2(n10501), .ZN(n13617) );
  INV_X1 U8630 ( .A(n13615), .ZN(n13602) );
  OR2_X1 U8631 ( .A1(n7937), .A2(n7936), .ZN(n7956) );
  NAND2_X1 U8632 ( .A1(n7954), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n7979) );
  INV_X1 U8633 ( .A(n7956), .ZN(n7954) );
  NAND2_X1 U8634 ( .A1(n7335), .A2(n6895), .ZN(n11897) );
  INV_X1 U8635 ( .A(n7336), .ZN(n7335) );
  NAND2_X1 U8636 ( .A1(n6898), .A2(n6686), .ZN(n6895) );
  OAI21_X1 U8637 ( .B1(n7338), .B2(n7337), .A(n11892), .ZN(n7336) );
  NOR2_X1 U8638 ( .A1(n7079), .A2(n6714), .ZN(n7078) );
  INV_X1 U8639 ( .A(n7081), .ZN(n7079) );
  NAND2_X1 U8640 ( .A1(n7328), .A2(n7329), .ZN(n11577) );
  AOI21_X1 U8641 ( .B1(n11526), .B2(n7330), .A(n6713), .ZN(n7329) );
  NAND2_X1 U8642 ( .A1(n10854), .A2(n7759), .ZN(n10865) );
  NOR2_X2 U8643 ( .A1(n11129), .A2(n10855), .ZN(n10872) );
  CLKBUF_X1 U8644 ( .A(n8289), .Z(n10825) );
  NOR2_X1 U8645 ( .A1(n9029), .A2(n13718), .ZN(n11493) );
  OR3_X1 U8646 ( .A1(n13763), .A2(n13762), .A3(n8410), .ZN(n13950) );
  OR2_X1 U8647 ( .A1(n8381), .A2(P2_IR_REG_23__SCAN_IN), .ZN(n8383) );
  OR2_X1 U8648 ( .A1(n8383), .A2(P2_IR_REG_24__SCAN_IN), .ZN(n8358) );
  NAND2_X1 U8649 ( .A1(n7974), .A2(n7699), .ZN(n8274) );
  NOR2_X1 U8650 ( .A1(n7569), .A2(n7655), .ZN(n7567) );
  NAND2_X1 U8651 ( .A1(n7570), .A2(n7718), .ZN(n7569) );
  AND2_X1 U8652 ( .A1(n7694), .A2(n7572), .ZN(n7570) );
  NAND2_X1 U8653 ( .A1(n7571), .A2(n6692), .ZN(n8080) );
  INV_X1 U8654 ( .A(n8077), .ZN(n7571) );
  INV_X1 U8655 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n8464) );
  NAND2_X1 U8656 ( .A1(n15101), .A2(n15103), .ZN(n15089) );
  NAND2_X1 U8657 ( .A1(n7525), .A2(n7528), .ZN(n12410) );
  OR2_X1 U8658 ( .A1(n12169), .A2(n12345), .ZN(n7525) );
  NOR2_X1 U8659 ( .A1(n9468), .A2(n9467), .ZN(n9480) );
  OR2_X1 U8660 ( .A1(n9595), .A2(n9594), .ZN(n9597) );
  INV_X1 U8661 ( .A(n7552), .ZN(n7551) );
  OR2_X1 U8662 ( .A1(n9453), .A2(n9452), .ZN(n9468) );
  AND2_X1 U8663 ( .A1(n12628), .A2(n12626), .ZN(n14121) );
  AND2_X1 U8664 ( .A1(n14120), .A2(n12615), .ZN(n14152) );
  AND2_X1 U8665 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n9416) );
  INV_X1 U8666 ( .A(n12350), .ZN(n7523) );
  AOI21_X1 U8667 ( .B1(n7528), .B2(n12345), .A(n7527), .ZN(n7526) );
  NOR2_X1 U8668 ( .A1(n6710), .A2(n12168), .ZN(n7527) );
  OR2_X1 U8669 ( .A1(n9607), .A2(n14164), .ZN(n9619) );
  INV_X1 U8670 ( .A(n9631), .ZN(n9302) );
  CLKBUF_X1 U8671 ( .A(n12503), .Z(n12486) );
  NAND2_X1 U8672 ( .A1(n9496), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n9507) );
  AND2_X1 U8673 ( .A1(n9480), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n9496) );
  NOR2_X1 U8674 ( .A1(n14180), .A2(n7553), .ZN(n7552) );
  INV_X1 U8675 ( .A(n12571), .ZN(n7553) );
  NAND2_X1 U8676 ( .A1(n14130), .A2(n7555), .ZN(n7554) );
  OAI21_X1 U8677 ( .B1(n11712), .B2(n7518), .A(n7515), .ZN(n11929) );
  OR2_X1 U8678 ( .A1(n11713), .A2(n11926), .ZN(n7518) );
  NAND2_X1 U8679 ( .A1(n9416), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n9429) );
  NOR2_X1 U8680 ( .A1(n9429), .A2(n9428), .ZN(n9440) );
  NAND2_X1 U8681 ( .A1(n9298), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9567) );
  INV_X1 U8682 ( .A(n9551), .ZN(n9298) );
  AOI21_X1 U8683 ( .B1(n7110), .B2(n7108), .A(n7107), .ZN(n7106) );
  INV_X1 U8684 ( .A(n7110), .ZN(n7109) );
  INV_X1 U8685 ( .A(n7673), .ZN(n7108) );
  AND3_X1 U8686 ( .A1(n9543), .A2(n9542), .A3(n9541), .ZN(n14948) );
  NAND2_X1 U8687 ( .A1(n14374), .A2(n14373), .ZN(n14417) );
  NOR2_X1 U8688 ( .A1(n14639), .A2(n14393), .ZN(n14630) );
  NAND2_X1 U8689 ( .A1(n7012), .A2(n7010), .ZN(n14637) );
  NAND2_X1 U8690 ( .A1(n7011), .A2(n7588), .ZN(n7010) );
  NAND2_X1 U8691 ( .A1(n14648), .A2(n7013), .ZN(n7012) );
  INV_X1 U8692 ( .A(n7015), .ZN(n7011) );
  NAND2_X1 U8693 ( .A1(n14668), .A2(n14656), .ZN(n14649) );
  OR2_X1 U8694 ( .A1(n14793), .A2(n14666), .ZN(n9677) );
  NAND2_X1 U8695 ( .A1(n7511), .A2(n14690), .ZN(n14685) );
  OR2_X1 U8696 ( .A1(n9643), .A2(n14098), .ZN(n9655) );
  INV_X1 U8697 ( .A(n7511), .ZN(n14696) );
  NAND2_X1 U8698 ( .A1(n9640), .A2(n14727), .ZN(n7150) );
  NOR2_X1 U8699 ( .A1(n6743), .A2(n6680), .ZN(n7149) );
  NAND2_X1 U8700 ( .A1(n14729), .A2(n14820), .ZN(n14711) );
  AND2_X1 U8701 ( .A1(n7451), .A2(n14442), .ZN(n7450) );
  NAND2_X1 U8702 ( .A1(n7448), .A2(n6687), .ZN(n7447) );
  NAND2_X1 U8703 ( .A1(n6872), .A2(n14746), .ZN(n14742) );
  INV_X1 U8704 ( .A(n6872), .ZN(n14760) );
  NAND2_X1 U8705 ( .A1(n7153), .A2(n7152), .ZN(n14756) );
  NAND2_X1 U8706 ( .A1(n6762), .A2(n14326), .ZN(n7152) );
  NAND2_X1 U8707 ( .A1(n9572), .A2(n6726), .ZN(n7153) );
  AND2_X1 U8708 ( .A1(n9363), .A2(n9362), .ZN(n14162) );
  NAND2_X1 U8709 ( .A1(n9565), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9595) );
  NAND2_X1 U8710 ( .A1(n7481), .A2(n9556), .ZN(n7480) );
  NAND2_X1 U8711 ( .A1(n7513), .A2(n7512), .ZN(n15121) );
  OR2_X1 U8712 ( .A1(n9507), .A2(n9506), .ZN(n9521) );
  NAND2_X1 U8713 ( .A1(n7455), .A2(n7458), .ZN(n11968) );
  NAND2_X1 U8714 ( .A1(n11911), .A2(n7460), .ZN(n7455) );
  OR2_X1 U8715 ( .A1(n11915), .A2(n14266), .ZN(n11916) );
  NAND2_X1 U8716 ( .A1(n11624), .A2(n15320), .ZN(n11915) );
  NAND2_X1 U8717 ( .A1(n7146), .A2(n6815), .ZN(n9448) );
  AND2_X1 U8718 ( .A1(n7143), .A2(n9446), .ZN(n6815) );
  AND2_X1 U8719 ( .A1(n11450), .A2(n12127), .ZN(n11624) );
  NAND2_X1 U8720 ( .A1(n11341), .A2(n15288), .ZN(n11471) );
  NAND2_X1 U8721 ( .A1(n11101), .A2(n9397), .ZN(n11340) );
  NOR2_X2 U8722 ( .A1(n11217), .A2(n14228), .ZN(n11341) );
  NAND2_X1 U8723 ( .A1(n7601), .A2(n14222), .ZN(n14418) );
  INV_X1 U8724 ( .A(n14391), .ZN(n14393) );
  NOR2_X1 U8725 ( .A1(n14445), .A2(n7614), .ZN(n7613) );
  INV_X1 U8726 ( .A(n9664), .ZN(n7614) );
  AND2_X1 U8727 ( .A1(n14682), .A2(n9664), .ZN(n14670) );
  INV_X1 U8728 ( .A(n14309), .ZN(n15148) );
  AND2_X1 U8729 ( .A1(n14928), .A2(n15313), .ZN(n15155) );
  NAND2_X1 U8730 ( .A1(n7468), .A2(n9734), .ZN(n14955) );
  NAND2_X1 U8731 ( .A1(n14924), .A2(n7593), .ZN(n7468) );
  XNOR2_X1 U8732 ( .A(n9233), .B(n9232), .ZN(n14372) );
  NAND2_X1 U8733 ( .A1(n7232), .A2(n8395), .ZN(n9209) );
  XNOR2_X1 U8734 ( .A(n8392), .B(n8391), .ZN(n12661) );
  XNOR2_X1 U8735 ( .A(n8256), .B(n8244), .ZN(n14079) );
  INV_X1 U8736 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n9764) );
  XNOR2_X1 U8737 ( .A(n8240), .B(n8225), .ZN(n12478) );
  XNOR2_X1 U8738 ( .A(n8182), .B(SI_22_), .ZN(n9628) );
  NOR2_X2 U8739 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n9700) );
  XNOR2_X1 U8740 ( .A(n6684), .B(n8145), .ZN(n12153) );
  NAND2_X1 U8741 ( .A1(n8137), .A2(n7021), .ZN(n7020) );
  XNOR2_X1 U8742 ( .A(n8137), .B(n6859), .ZN(n12015) );
  XNOR2_X1 U8743 ( .A(n8135), .B(n11515), .ZN(n6859) );
  INV_X1 U8744 ( .A(n9320), .ZN(n9573) );
  CLKBUF_X1 U8745 ( .A(n9558), .Z(n9559) );
  OR2_X1 U8746 ( .A1(n9491), .A2(n9490), .ZN(n9547) );
  NAND2_X1 U8747 ( .A1(n7931), .A2(n7930), .ZN(n7950) );
  NAND2_X1 U8748 ( .A1(n7005), .A2(n7907), .ZN(n7911) );
  INV_X1 U8749 ( .A(n7220), .ZN(n7219) );
  AND2_X1 U8750 ( .A1(n9476), .A2(n9464), .ZN(n14594) );
  XNOR2_X1 U8751 ( .A(n7906), .B(n7904), .ZN(n10487) );
  NAND2_X1 U8752 ( .A1(n7888), .A2(n7887), .ZN(n7906) );
  NAND2_X1 U8753 ( .A1(n6854), .A2(n7867), .ZN(n7872) );
  NAND2_X1 U8754 ( .A1(n7872), .A2(n7871), .ZN(n7888) );
  NAND2_X1 U8755 ( .A1(n7848), .A2(n6913), .ZN(n6915) );
  NOR2_X1 U8756 ( .A1(n7851), .A2(n6914), .ZN(n6913) );
  INV_X1 U8757 ( .A(n7847), .ZN(n6914) );
  NOR2_X1 U8759 ( .A1(n9409), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n9412) );
  AND2_X1 U8760 ( .A1(n9412), .A2(n9411), .ZN(n9560) );
  OR2_X1 U8761 ( .A1(n9398), .A2(P1_IR_REG_3__SCAN_IN), .ZN(n9409) );
  NAND2_X1 U8762 ( .A1(n9379), .A2(n9310), .ZN(n9398) );
  INV_X1 U8763 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n9310) );
  INV_X1 U8764 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n9952) );
  AND2_X1 U8765 ( .A1(n9900), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n7226) );
  XNOR2_X1 U8766 ( .A(n9901), .B(P3_ADDR_REG_2__SCAN_IN), .ZN(n9947) );
  XNOR2_X1 U8767 ( .A(n9943), .B(P1_ADDR_REG_4__SCAN_IN), .ZN(n9945) );
  NOR2_X1 U8768 ( .A1(n9908), .A2(n9909), .ZN(n9962) );
  XNOR2_X1 U8769 ( .A(n9912), .B(n9913), .ZN(n9966) );
  XOR2_X1 U8770 ( .A(n9941), .B(n9940), .Z(n9969) );
  OAI21_X1 U8771 ( .B1(n15202), .B2(n15201), .A(n7180), .ZN(n7179) );
  OAI22_X1 U8772 ( .A1(n9981), .A2(n9923), .B1(P1_ADDR_REG_13__SCAN_IN), .B2(
        n9979), .ZN(n9934) );
  XNOR2_X1 U8773 ( .A(n12819), .B(n9870), .ZN(n11820) );
  NAND2_X1 U8774 ( .A1(n7366), .A2(n7371), .ZN(n12332) );
  NAND2_X1 U8775 ( .A1(n12218), .A2(n7373), .ZN(n7366) );
  NAND2_X1 U8776 ( .A1(n12747), .A2(n7344), .ZN(n12695) );
  NAND2_X1 U8777 ( .A1(n8838), .A2(n8837), .ZN(n13163) );
  OAI211_X1 U8778 ( .C1(SI_10_), .C2(n12806), .A(n8635), .B(n8634), .ZN(n15647) );
  OR2_X1 U8779 ( .A1(n9845), .A2(n13248), .ZN(n6958) );
  NAND2_X1 U8780 ( .A1(n6952), .A2(n6728), .ZN(n12682) );
  NAND2_X1 U8781 ( .A1(n12721), .A2(n6953), .ZN(n6952) );
  NAND2_X1 U8782 ( .A1(n6953), .A2(n6955), .ZN(n6951) );
  INV_X1 U8783 ( .A(n7351), .ZN(n7350) );
  OAI21_X1 U8784 ( .B1(n7353), .B2(n7352), .A(n11831), .ZN(n7351) );
  INV_X1 U8785 ( .A(n9817), .ZN(n7352) );
  NAND2_X1 U8786 ( .A1(n11818), .A2(n9817), .ZN(n11832) );
  NAND3_X1 U8787 ( .A1(n7342), .A2(n7341), .A3(n9800), .ZN(n11027) );
  NAND2_X1 U8788 ( .A1(n12758), .A2(n9852), .ZN(n12710) );
  AOI21_X1 U8789 ( .B1(n13151), .B2(n10356), .A(n8863), .ZN(n12726) );
  AOI21_X1 U8790 ( .B1(n7364), .B2(n7367), .A(n7362), .ZN(n7361) );
  INV_X1 U8791 ( .A(n12435), .ZN(n7362) );
  NAND2_X1 U8792 ( .A1(n11534), .A2(n9809), .ZN(n11651) );
  NAND2_X1 U8793 ( .A1(n9849), .A2(n9848), .ZN(n12760) );
  NAND2_X1 U8794 ( .A1(n7375), .A2(n7372), .ZN(n12282) );
  INV_X1 U8795 ( .A(n7374), .ZN(n7372) );
  NAND2_X1 U8796 ( .A1(n7377), .A2(n7376), .ZN(n7375) );
  OAI21_X1 U8797 ( .B1(n9859), .B2(n9858), .A(n9860), .ZN(n12769) );
  NAND2_X1 U8798 ( .A1(n11027), .A2(n7341), .ZN(n11172) );
  NOR2_X1 U8799 ( .A1(n12739), .A2(n9844), .ZN(n12781) );
  NAND2_X1 U8800 ( .A1(n12781), .A2(n12780), .ZN(n12779) );
  NAND2_X1 U8801 ( .A1(n9891), .A2(n9890), .ZN(n12790) );
  AND2_X1 U8802 ( .A1(n9879), .A2(n9878), .ZN(n12794) );
  AND2_X1 U8803 ( .A1(n8877), .A2(n8876), .ZN(n13149) );
  NAND2_X1 U8804 ( .A1(n6957), .A2(n6956), .ZN(n12786) );
  AND2_X1 U8805 ( .A1(n9875), .A2(n10907), .ZN(n12788) );
  NAND2_X1 U8806 ( .A1(n8718), .A2(n8717), .ZN(n13282) );
  NAND2_X1 U8807 ( .A1(n7240), .A2(n9003), .ZN(n7239) );
  OR2_X1 U8808 ( .A1(n7246), .A2(n15708), .ZN(n7245) );
  NAND4_X1 U8809 ( .A1(n8674), .A2(n8673), .A3(n8672), .A4(n8671), .ZN(n15042)
         );
  OR2_X1 U8810 ( .A1(n11986), .A2(n8481), .ZN(n8482) );
  OR2_X1 U8811 ( .A1(n8524), .A2(n8452), .ZN(n8458) );
  NAND2_X1 U8812 ( .A1(n8680), .A2(P3_IR_REG_2__SCAN_IN), .ZN(n7028) );
  NAND3_X1 U8813 ( .A1(n7030), .A2(n7029), .A3(P3_IR_REG_2__SCAN_IN), .ZN(
        n7025) );
  XNOR2_X1 U8814 ( .A(n8515), .B(P3_IR_REG_4__SCAN_IN), .ZN(n10982) );
  NOR2_X1 U8815 ( .A1(P3_IR_REG_2__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .ZN(
        n7349) );
  AOI22_X1 U8816 ( .A1(n11155), .A2(n11154), .B1(n11153), .B2(n11152), .ZN(
        n11316) );
  NOR2_X1 U8817 ( .A1(n11323), .A2(n11322), .ZN(n11841) );
  NOR2_X1 U8818 ( .A1(n11843), .A2(n15550), .ZN(n11845) );
  NAND2_X1 U8819 ( .A1(n15561), .A2(n11849), .ZN(n11850) );
  NOR2_X1 U8820 ( .A1(n15568), .A2(n8651), .ZN(n15567) );
  NAND2_X1 U8821 ( .A1(n7292), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n7291) );
  NAND2_X1 U8822 ( .A1(n12998), .A2(n7292), .ZN(n7290) );
  INV_X1 U8823 ( .A(n15584), .ZN(n7292) );
  AOI21_X1 U8824 ( .B1(n13015), .B2(n13014), .A(n15578), .ZN(n15595) );
  AOI21_X1 U8825 ( .B1(n13020), .B2(n13019), .A(n15608), .ZN(n15633) );
  INV_X1 U8826 ( .A(n7293), .ZN(n13002) );
  AOI21_X1 U8827 ( .B1(n13028), .B2(n13058), .A(n14977), .ZN(n15002) );
  NOR2_X1 U8828 ( .A1(n15006), .A2(n13006), .ZN(n15034) );
  INV_X1 U8829 ( .A(n7286), .ZN(n13005) );
  AND2_X1 U8830 ( .A1(n10921), .A2(n10917), .ZN(n15032) );
  INV_X1 U8831 ( .A(n13065), .ZN(n7033) );
  XNOR2_X1 U8832 ( .A(n7035), .B(n13064), .ZN(n7034) );
  NAND2_X1 U8833 ( .A1(n15024), .A2(n6799), .ZN(n7035) );
  NAND2_X1 U8834 ( .A1(n15540), .A2(n7356), .ZN(n7032) );
  NOR2_X1 U8835 ( .A1(n15035), .A2(n6868), .ZN(n13009) );
  NOR2_X1 U8836 ( .A1(n15023), .A2(n13007), .ZN(n6868) );
  XNOR2_X1 U8837 ( .A(n12798), .B(n10364), .ZN(n13074) );
  OAI21_X1 U8838 ( .B1(n8969), .B2(n15707), .A(n7117), .ZN(n13101) );
  AOI21_X1 U8839 ( .B1(n8957), .B2(n15703), .A(n6817), .ZN(n7117) );
  INV_X1 U8840 ( .A(n8968), .ZN(n6817) );
  NAND2_X1 U8841 ( .A1(n8868), .A2(n8867), .ZN(n13134) );
  AND2_X1 U8842 ( .A1(n13190), .A2(n8944), .ZN(n13174) );
  NAND2_X1 U8843 ( .A1(n8773), .A2(n8772), .ZN(n13240) );
  NAND2_X1 U8844 ( .A1(n13265), .A2(n13264), .ZN(n8744) );
  NAND2_X1 U8845 ( .A1(n12358), .A2(n8934), .ZN(n13290) );
  NAND2_X1 U8846 ( .A1(n15050), .A2(n12903), .ZN(n12369) );
  INV_X1 U8847 ( .A(n15054), .ZN(n15649) );
  NAND2_X1 U8848 ( .A1(n7397), .A2(n12894), .ZN(n15646) );
  NAND2_X1 U8849 ( .A1(n11676), .A2(n8924), .ZN(n11788) );
  AND2_X1 U8850 ( .A1(n8506), .A2(n7127), .ZN(n12021) );
  AND2_X1 U8851 ( .A1(n8507), .A2(n6721), .ZN(n7127) );
  NOR2_X1 U8852 ( .A1(n15053), .A2(n15730), .ZN(n15673) );
  AND2_X1 U8853 ( .A1(n8467), .A2(n8466), .ZN(n7396) );
  OR2_X1 U8854 ( .A1(n11362), .A2(n15708), .ZN(n15675) );
  INV_X1 U8855 ( .A(n15673), .ZN(n13297) );
  AOI22_X1 U8856 ( .A1(n12800), .A2(n12805), .B1(SI_30_), .B2(n12799), .ZN(
        n13373) );
  INV_X1 U8857 ( .A(n13118), .ZN(n13381) );
  AND2_X1 U8858 ( .A1(n13319), .A2(n13318), .ZN(n13382) );
  AOI21_X1 U8859 ( .B1(n11513), .B2(n12805), .A(n8795), .ZN(n13402) );
  NAND2_X1 U8860 ( .A1(n8702), .A2(n8701), .ZN(n13423) );
  INV_X1 U8861 ( .A(n12021), .ZN(n7126) );
  AND2_X1 U8862 ( .A1(n8988), .A2(n8987), .ZN(n13425) );
  AND2_X1 U8863 ( .A1(n10910), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13426) );
  OAI21_X1 U8864 ( .B1(n12692), .B2(n12691), .A(n12802), .ZN(n12800) );
  XNOR2_X1 U8865 ( .A(n10349), .B(n10345), .ZN(n12664) );
  NAND2_X1 U8866 ( .A1(n6706), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8460) );
  NAND2_X1 U8867 ( .A1(n8461), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8463) );
  NOR2_X1 U8868 ( .A1(n7634), .A2(n6964), .ZN(n6962) );
  NAND2_X1 U8869 ( .A1(n7279), .A2(n8864), .ZN(n8865) );
  NAND2_X1 U8870 ( .A1(n8822), .A2(n8821), .ZN(n8834) );
  XNOR2_X1 U8871 ( .A(n8436), .B(n8435), .ZN(n11693) );
  NAND2_X1 U8872 ( .A1(n8910), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8912) );
  INV_X1 U8873 ( .A(n9015), .ZN(n11514) );
  XNOR2_X1 U8874 ( .A(n8439), .B(n8438), .ZN(n13037) );
  OAI21_X1 U8875 ( .B1(n8768), .B2(n7262), .A(n7260), .ZN(n8794) );
  NAND2_X1 U8876 ( .A1(n8781), .A2(n8780), .ZN(n8784) );
  INV_X1 U8877 ( .A(SI_16_), .ZN(n10711) );
  OAI21_X1 U8878 ( .B1(n8713), .B2(n7256), .A(n7254), .ZN(n8746) );
  NAND2_X1 U8879 ( .A1(n8728), .A2(n8727), .ZN(n8731) );
  INV_X1 U8880 ( .A(SI_15_), .ZN(n10594) );
  NAND2_X1 U8881 ( .A1(n7270), .A2(n7274), .ZN(n8692) );
  NAND2_X1 U8882 ( .A1(n7272), .A2(n7274), .ZN(n8678) );
  INV_X1 U8883 ( .A(SI_12_), .ZN(n10457) );
  OAI21_X1 U8884 ( .B1(n8628), .B2(n7053), .A(n7051), .ZN(n8659) );
  NAND2_X1 U8885 ( .A1(n8638), .A2(n8637), .ZN(n8641) );
  INV_X1 U8886 ( .A(SI_11_), .ZN(n10450) );
  NAND2_X1 U8887 ( .A1(n7263), .A2(n7268), .ZN(n8607) );
  NAND2_X1 U8888 ( .A1(n8575), .A2(n8587), .ZN(n7263) );
  INV_X1 U8889 ( .A(n11325), .ZN(n11853) );
  INV_X1 U8890 ( .A(n11153), .ZN(n11163) );
  OAI21_X1 U8891 ( .B1(n8519), .B2(n7047), .A(n7044), .ZN(n8553) );
  NAND2_X1 U8892 ( .A1(n8519), .A2(n8518), .ZN(n8537) );
  NAND2_X1 U8893 ( .A1(n12246), .A2(n12245), .ZN(n12248) );
  NAND2_X1 U8894 ( .A1(n11875), .A2(n6679), .ZN(n12067) );
  NAND2_X1 U8895 ( .A1(n11875), .A2(n11874), .ZN(n11882) );
  NAND2_X1 U8896 ( .A1(n7560), .A2(n11266), .ZN(n13511) );
  NOR2_X1 U8897 ( .A1(n6933), .A2(n6935), .ZN(n6929) );
  OAI211_X1 U8898 ( .C1(n13554), .C2(n6932), .A(n6928), .B(n6931), .ZN(n13540)
         );
  OAI21_X1 U8899 ( .B1(n11436), .B2(n6907), .A(n6906), .ZN(n11664) );
  NAND2_X1 U8900 ( .A1(n11660), .A2(n11500), .ZN(n6907) );
  NAND2_X1 U8901 ( .A1(n6908), .A2(n11660), .ZN(n6906) );
  INV_X1 U8902 ( .A(n7584), .ZN(n7583) );
  OAI21_X1 U8903 ( .B1(n13521), .B2(n7585), .A(n13584), .ZN(n7584) );
  INV_X1 U8904 ( .A(n6703), .ZN(n7585) );
  NAND2_X1 U8905 ( .A1(n6888), .A2(n6892), .ZN(n13561) );
  NAND2_X1 U8906 ( .A1(n13442), .A2(n13441), .ZN(n13562) );
  NAND2_X1 U8907 ( .A1(n12469), .A2(n13441), .ZN(n6888) );
  NAND2_X1 U8908 ( .A1(n9025), .A2(n11491), .ZN(n11125) );
  AND2_X1 U8909 ( .A1(n13520), .A2(n13461), .ZN(n13581) );
  INV_X1 U8910 ( .A(n7574), .ZN(n7573) );
  OAI21_X1 U8911 ( .B1(n6679), .B2(n7575), .A(n7674), .ZN(n7574) );
  AOI21_X1 U8912 ( .B1(n6892), .B2(n6891), .A(n6890), .ZN(n6889) );
  INV_X1 U8913 ( .A(n13441), .ZN(n6891) );
  NAND2_X1 U8914 ( .A1(n11436), .A2(n11417), .ZN(n11423) );
  NAND2_X1 U8915 ( .A1(n11436), .A2(n7586), .ZN(n11501) );
  NAND2_X1 U8916 ( .A1(n13491), .A2(n13490), .ZN(n13614) );
  AND2_X1 U8917 ( .A1(n8247), .A2(n8229), .ZN(n13779) );
  AND2_X1 U8918 ( .A1(n7183), .A2(n9254), .ZN(n7002) );
  NAND2_X1 U8919 ( .A1(n7774), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n7750) );
  AND2_X1 U8920 ( .A1(n10796), .A2(n10795), .ZN(n11069) );
  AOI21_X1 U8921 ( .B1(n10788), .B2(n11070), .A(n11064), .ZN(n15395) );
  OR2_X1 U8922 ( .A1(n15409), .A2(n15408), .ZN(n15410) );
  OR2_X1 U8923 ( .A1(n13699), .A2(n13698), .ZN(n13711) );
  NAND2_X1 U8924 ( .A1(n7170), .A2(n11777), .ZN(n13939) );
  INV_X1 U8925 ( .A(n14029), .ZN(n13736) );
  NOR2_X1 U8926 ( .A1(n13760), .A2(n7490), .ZN(n7489) );
  INV_X1 U8927 ( .A(n8237), .ZN(n7490) );
  NAND2_X1 U8928 ( .A1(n8238), .A2(n8237), .ZN(n13761) );
  OR3_X1 U8929 ( .A1(n13793), .A2(n13792), .A3(n8410), .ZN(n13958) );
  OR2_X1 U8930 ( .A1(n13789), .A2(n13788), .ZN(n13959) );
  OAI21_X1 U8931 ( .B1(n13838), .B2(n6920), .A(n6919), .ZN(n13787) );
  NAND2_X1 U8932 ( .A1(n13819), .A2(n7503), .ZN(n13808) );
  AND2_X1 U8933 ( .A1(n13819), .A2(n8178), .ZN(n7691) );
  AND2_X1 U8934 ( .A1(n13840), .A2(n13839), .ZN(n13977) );
  NAND2_X1 U8935 ( .A1(n7088), .A2(n8134), .ZN(n13853) );
  NAND2_X1 U8936 ( .A1(n8113), .A2(n6709), .ZN(n7088) );
  NAND2_X1 U8937 ( .A1(n13862), .A2(n13861), .ZN(n13864) );
  NAND2_X1 U8938 ( .A1(n8113), .A2(n8112), .ZN(n13871) );
  NAND2_X1 U8939 ( .A1(n13911), .A2(n8089), .ZN(n13887) );
  NAND2_X1 U8940 ( .A1(n8322), .A2(n7334), .ZN(n7332) );
  NAND2_X1 U8941 ( .A1(n8322), .A2(n8321), .ZN(n12424) );
  NAND2_X1 U8942 ( .A1(n7495), .A2(n8024), .ZN(n12387) );
  NAND2_X1 U8943 ( .A1(n7498), .A2(n8007), .ZN(n12269) );
  NAND2_X1 U8944 ( .A1(n6944), .A2(n6946), .ZN(n12258) );
  NAND2_X1 U8945 ( .A1(n6945), .A2(n8313), .ZN(n12199) );
  NAND2_X1 U8946 ( .A1(n8311), .A2(n6949), .ZN(n6945) );
  INV_X1 U8947 ( .A(n7090), .ZN(n12054) );
  NAND2_X1 U8948 ( .A1(n8311), .A2(n8310), .ZN(n12056) );
  NAND2_X1 U8949 ( .A1(n7096), .A2(n7945), .ZN(n11957) );
  NAND2_X1 U8950 ( .A1(n8306), .A2(n8305), .ZN(n11773) );
  INV_X1 U8951 ( .A(n13933), .ZN(n13824) );
  NAND2_X1 U8952 ( .A1(n6898), .A2(n8303), .ZN(n11614) );
  NAND2_X1 U8953 ( .A1(n11575), .A2(n7846), .ZN(n11591) );
  AND2_X1 U8954 ( .A1(n7080), .A2(n7081), .ZN(n11590) );
  NAND2_X1 U8955 ( .A1(n7331), .A2(n8295), .ZN(n11525) );
  NAND2_X1 U8956 ( .A1(n11088), .A2(n11087), .ZN(n7331) );
  NAND2_X1 U8957 ( .A1(n7076), .A2(n10858), .ZN(n10853) );
  INV_X1 U8958 ( .A(n13922), .ZN(n13930) );
  INV_X1 U8959 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n6924) );
  INV_X1 U8960 ( .A(n13729), .ZN(n14025) );
  INV_X1 U8961 ( .A(n13859), .ZN(n14048) );
  NAND2_X1 U8962 ( .A1(n8018), .A2(n8017), .ZN(n12310) );
  INV_X1 U8963 ( .A(n13932), .ZN(n11459) );
  AND2_X1 U8964 ( .A1(n11277), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15470) );
  MUX2_X1 U8965 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7725), .S(
        P2_IR_REG_29__SCAN_IN), .Z(n7729) );
  XNOR2_X1 U8966 ( .A(n8362), .B(P2_IR_REG_26__SCAN_IN), .ZN(n12479) );
  NAND2_X2 U8967 ( .A1(n8285), .A2(n8381), .ZN(n12531) );
  INV_X1 U8968 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n11735) );
  INV_X1 U8969 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n11549) );
  INV_X1 U8970 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n10499) );
  INV_X1 U8971 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n10491) );
  INV_X1 U8972 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n10490) );
  INV_X1 U8973 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n10469) );
  INV_X1 U8974 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n10458) );
  INV_X1 U8975 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n10431) );
  INV_X1 U8976 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n10468) );
  INV_X1 U8977 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n10413) );
  INV_X1 U8978 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n10410) );
  INV_X1 U8979 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n10412) );
  OAI21_X1 U8980 ( .B1(n14188), .B2(n12634), .A(n7544), .ZN(n14086) );
  NAND2_X1 U8981 ( .A1(n15089), .A2(n12549), .ZN(n15093) );
  AND2_X1 U8982 ( .A1(n9528), .A2(n9527), .ZN(n15087) );
  NAND2_X1 U8983 ( .A1(n14094), .A2(n14095), .ZN(n7537) );
  NOR2_X1 U8984 ( .A1(n11198), .A2(n11199), .ZN(n11711) );
  NAND2_X1 U8985 ( .A1(n9657), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n9386) );
  AOI21_X1 U8986 ( .B1(n7544), .B2(n12634), .A(n12643), .ZN(n7543) );
  NAND2_X1 U8987 ( .A1(n6851), .A2(n12168), .ZN(n12347) );
  CLKBUF_X1 U8988 ( .A(n12169), .Z(n6851) );
  NAND2_X1 U8989 ( .A1(n12587), .A2(n12586), .ZN(n14114) );
  OAI21_X1 U8990 ( .B1(n14130), .B2(n7103), .A(n7101), .ZN(n12587) );
  NAND2_X1 U8991 ( .A1(n12486), .A2(n7673), .ZN(n12539) );
  INV_X1 U8992 ( .A(n7521), .ZN(n11741) );
  NAND2_X1 U8993 ( .A1(n7100), .A2(n7104), .ZN(n14160) );
  NAND2_X1 U8994 ( .A1(n14130), .A2(n7547), .ZN(n7100) );
  AOI21_X1 U8995 ( .B1(n7101), .B2(n7103), .A(n6761), .ZN(n7098) );
  NAND2_X1 U8996 ( .A1(n14130), .A2(n7101), .ZN(n7099) );
  NAND2_X1 U8997 ( .A1(n7554), .A2(n12571), .ZN(n14179) );
  NAND2_X1 U8998 ( .A1(n10741), .A2(n10740), .ZN(n15092) );
  AND2_X1 U8999 ( .A1(n10726), .A2(n15136), .ZN(n15111) );
  XNOR2_X1 U9000 ( .A(n12556), .B(n12557), .ZN(n14200) );
  NAND2_X1 U9001 ( .A1(n14200), .A2(n14199), .ZN(n14198) );
  INV_X1 U9002 ( .A(n15092), .ZN(n15114) );
  NAND2_X1 U9003 ( .A1(n9331), .A2(n9330), .ZN(n14481) );
  INV_X1 U9004 ( .A(n11203), .ZN(n14502) );
  CLKBUF_X1 U9005 ( .A(n14503), .Z(n6847) );
  INV_X1 U9006 ( .A(n14462), .ZN(n14772) );
  INV_X1 U9007 ( .A(n14417), .ZN(n14775) );
  INV_X1 U9008 ( .A(n12525), .ZN(n14789) );
  INV_X1 U9009 ( .A(n14786), .ZN(n14093) );
  NAND2_X1 U9010 ( .A1(n6857), .A2(n6856), .ZN(n6855) );
  AOI21_X1 U9011 ( .B1(n12522), .B2(n12523), .A(n15175), .ZN(n6858) );
  INV_X1 U9012 ( .A(n12524), .ZN(n6856) );
  NAND2_X1 U9013 ( .A1(n9666), .A2(n9665), .ZN(n14674) );
  NAND2_X1 U9014 ( .A1(n14680), .A2(n7445), .ZN(n14663) );
  AND2_X1 U9015 ( .A1(n14814), .A2(n9652), .ZN(n14684) );
  NAND2_X1 U9016 ( .A1(n14726), .A2(n9627), .ZN(n14708) );
  NAND2_X1 U9017 ( .A1(n14737), .A2(n7454), .ZN(n14723) );
  NAND2_X1 U9018 ( .A1(n7607), .A2(n7605), .ZN(n14748) );
  AND2_X1 U9019 ( .A1(n7446), .A2(n14331), .ZN(n14738) );
  AND2_X1 U9020 ( .A1(n9593), .A2(n9592), .ZN(n14323) );
  NAND2_X1 U9021 ( .A1(n7155), .A2(n9713), .ZN(n12510) );
  NAND2_X1 U9022 ( .A1(n9572), .A2(n7156), .ZN(n7155) );
  NAND2_X1 U9023 ( .A1(n9572), .A2(n9571), .ZN(n12444) );
  NAND2_X1 U9024 ( .A1(n7484), .A2(n14303), .ZN(n15129) );
  NAND2_X1 U9025 ( .A1(n15163), .A2(n9544), .ZN(n12315) );
  NAND2_X1 U9026 ( .A1(n9534), .A2(n9533), .ZN(n15164) );
  AND2_X1 U9027 ( .A1(n9519), .A2(n9518), .ZN(n15112) );
  NAND2_X1 U9028 ( .A1(n7137), .A2(n7139), .ZN(n14953) );
  OR2_X1 U9029 ( .A1(n9487), .A2(n7141), .ZN(n7137) );
  INV_X1 U9030 ( .A(n14957), .ZN(n14920) );
  OAI21_X1 U9031 ( .B1(n9487), .B2(n7597), .A(n7594), .ZN(n14916) );
  NAND2_X1 U9032 ( .A1(n9487), .A2(n9486), .ZN(n11972) );
  NAND2_X1 U9033 ( .A1(n7462), .A2(n9730), .ZN(n11803) );
  NAND2_X1 U9034 ( .A1(n7464), .A2(n7463), .ZN(n7462) );
  AND2_X1 U9035 ( .A1(n7143), .A2(n7146), .ZN(n11479) );
  NAND2_X1 U9036 ( .A1(n7598), .A2(n9423), .ZN(n11443) );
  NAND2_X1 U9037 ( .A1(n11464), .A2(n14425), .ZN(n7598) );
  NAND2_X1 U9038 ( .A1(n14407), .A2(n10411), .ZN(n9382) );
  AND2_X1 U9039 ( .A1(n15143), .A2(n10393), .ZN(n14717) );
  AOI21_X1 U9040 ( .B1(n14782), .B2(n15337), .A(n14781), .ZN(n14783) );
  NAND2_X1 U9041 ( .A1(n7199), .A2(n7188), .ZN(n7187) );
  INV_X1 U9042 ( .A(n7200), .ZN(n7188) );
  INV_X1 U9043 ( .A(n9324), .ZN(n14878) );
  NAND2_X1 U9044 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_29__SCAN_IN), 
        .ZN(n7617) );
  NAND2_X1 U9045 ( .A1(n9322), .A2(n9424), .ZN(n7616) );
  XNOR2_X1 U9046 ( .A(n9761), .B(P1_IR_REG_24__SCAN_IN), .ZN(n12328) );
  OAI21_X1 U9047 ( .B1(n9770), .B2(P1_IR_REG_23__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9761) );
  XNOR2_X1 U9048 ( .A(n8164), .B(n8163), .ZN(n12301) );
  XNOR2_X1 U9049 ( .A(n9629), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n14892) );
  OR2_X1 U9050 ( .A1(n9628), .A2(n6671), .ZN(n9629) );
  INV_X1 U9051 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n9709) );
  INV_X1 U9052 ( .A(n9352), .ZN(n9350) );
  INV_X1 U9053 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n11691) );
  INV_X1 U9054 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n11547) );
  INV_X1 U9055 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n10748) );
  INV_X1 U9056 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n10497) );
  INV_X1 U9057 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n10493) );
  INV_X1 U9058 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n10488) );
  INV_X1 U9059 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n10472) );
  INV_X1 U9060 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n10461) );
  NAND2_X1 U9061 ( .A1(n6854), .A2(n6915), .ZN(n10460) );
  INV_X1 U9062 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n10438) );
  INV_X1 U9063 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n10443) );
  INV_X1 U9064 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n10436) );
  INV_X1 U9065 ( .A(n7789), .ZN(n7786) );
  NAND2_X1 U9066 ( .A1(n7770), .A2(n7784), .ZN(n10440) );
  INV_X1 U9067 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n10462) );
  NAND2_X1 U9068 ( .A1(n6885), .A2(n7722), .ZN(n7741) );
  NOR2_X1 U9069 ( .A1(n9954), .A2(n15766), .ZN(n14900) );
  XNOR2_X1 U9070 ( .A(n9945), .B(P2_ADDR_REG_4__SCAN_IN), .ZN(n15753) );
  XNOR2_X1 U9071 ( .A(n9967), .B(P2_ADDR_REG_7__SCAN_IN), .ZN(n15760) );
  INV_X1 U9072 ( .A(n9969), .ZN(n7222) );
  AND2_X2 U9073 ( .A1(n7178), .A2(n6718), .ZN(n14914) );
  NAND2_X1 U9074 ( .A1(n7521), .A2(n7520), .ZN(n7519) );
  INV_X1 U9075 ( .A(n11740), .ZN(n7520) );
  NAND2_X1 U9076 ( .A1(n11238), .A2(n9807), .ZN(n11536) );
  NOR2_X1 U9077 ( .A1(n6788), .A2(n6832), .ZN(n6831) );
  NOR2_X1 U9078 ( .A1(n15751), .A2(n10381), .ZN(n6832) );
  NOR2_X1 U9079 ( .A1(n6691), .A2(n6834), .ZN(n6833) );
  NOR2_X1 U9080 ( .A1(n15741), .A2(n10378), .ZN(n6834) );
  NAND2_X1 U9081 ( .A1(n7116), .A2(n7114), .ZN(P3_U3454) );
  NOR2_X1 U9082 ( .A1(n6787), .A2(n7115), .ZN(n7114) );
  OR2_X1 U9083 ( .A1(n9021), .A2(n15743), .ZN(n7116) );
  NOR2_X1 U9084 ( .A1(n15741), .A2(n9009), .ZN(n7115) );
  OAI21_X1 U9085 ( .B1(n11436), .B2(n6911), .A(n6905), .ZN(n11661) );
  NAND2_X1 U9086 ( .A1(n13512), .A2(n11273), .ZN(n11275) );
  NAND2_X1 U9087 ( .A1(n6865), .A2(n6861), .ZN(n13721) );
  NAND2_X1 U9088 ( .A1(n6864), .A2(n6862), .ZN(n6861) );
  NAND2_X1 U9089 ( .A1(n13719), .A2(n13718), .ZN(n6865) );
  AND3_X1 U9090 ( .A1(n7308), .A2(n7309), .A3(n7314), .ZN(n13747) );
  AOI21_X1 U9091 ( .B1(n13744), .B2(n14002), .A(n8414), .ZN(n8415) );
  NAND2_X1 U9092 ( .A1(n15536), .A2(n6924), .ZN(n6923) );
  OAI21_X1 U9093 ( .B1(n14023), .B2(n15523), .A(n7167), .ZN(P2_U3498) );
  NOR2_X1 U9094 ( .A1(n7169), .A2(n7168), .ZN(n7167) );
  NOR2_X1 U9095 ( .A1(n15524), .A2(n14024), .ZN(n7168) );
  NOR2_X1 U9096 ( .A1(n14025), .A2(n14062), .ZN(n7169) );
  AOI21_X1 U9097 ( .B1(n13744), .B2(n8423), .A(n8422), .ZN(n8424) );
  OR2_X1 U9098 ( .A1(n15524), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n7097) );
  OR2_X1 U9099 ( .A1(n14474), .A2(n14473), .ZN(n6809) );
  INV_X1 U9100 ( .A(n10403), .ZN(n10404) );
  OAI21_X1 U9101 ( .B1(n10402), .B2(n14765), .A(n10401), .ZN(n10403) );
  NAND2_X1 U9102 ( .A1(n15355), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n7472) );
  NAND2_X1 U9103 ( .A1(n14776), .A2(n15358), .ZN(n7473) );
  INV_X1 U9104 ( .A(n7178), .ZN(n14909) );
  INV_X1 U9105 ( .A(n7182), .ZN(n15196) );
  INV_X1 U9106 ( .A(n7201), .ZN(n15213) );
  INV_X1 U9107 ( .A(n14895), .ZN(n6849) );
  XNOR2_X1 U9108 ( .A(n10340), .B(n9992), .ZN(n7227) );
  INV_X1 U9109 ( .A(n12090), .ZN(n7172) );
  AND4_X2 U9110 ( .A1(n7654), .A2(n7854), .A3(n7791), .A4(n7653), .ZN(n6677)
         );
  AND2_X1 U9112 ( .A1(n12867), .A2(n12876), .ZN(n6678) );
  INV_X1 U9113 ( .A(n14923), .ZN(n7593) );
  INV_X1 U9114 ( .A(n9286), .ZN(n7313) );
  NAND2_X1 U9115 ( .A1(n14881), .A2(n9324), .ZN(n9392) );
  INV_X1 U9116 ( .A(n9392), .ZN(n9383) );
  AND2_X1 U9117 ( .A1(n7577), .A2(n11874), .ZN(n6679) );
  XNOR2_X1 U9118 ( .A(n7637), .B(P3_IR_REG_29__SCAN_IN), .ZN(n8453) );
  AND2_X1 U9119 ( .A1(n14820), .A2(n14344), .ZN(n6680) );
  AND2_X1 U9120 ( .A1(n14210), .A2(n14387), .ZN(n6681) );
  INV_X1 U9121 ( .A(n9282), .ZN(n7321) );
  OR2_X1 U9122 ( .A1(n9174), .A2(n9175), .ZN(n6682) );
  OR2_X1 U9123 ( .A1(n12205), .A2(n13644), .ZN(n6683) );
  INV_X1 U9124 ( .A(n9739), .ZN(n7476) );
  AND2_X1 U9125 ( .A1(n7020), .A2(n6785), .ZN(n6684) );
  INV_X1 U9126 ( .A(n14493), .ZN(n12492) );
  INV_X1 U9127 ( .A(n12219), .ZN(n7376) );
  AND2_X1 U9128 ( .A1(n9700), .A2(n9315), .ZN(n6685) );
  NAND2_X1 U9129 ( .A1(n9606), .A2(n9605), .ZN(n14832) );
  INV_X1 U9130 ( .A(n14832), .ZN(n14746) );
  AND2_X1 U9131 ( .A1(n6896), .A2(n11893), .ZN(n6686) );
  OR2_X1 U9132 ( .A1(n7453), .A2(n14827), .ZN(n6687) );
  AND2_X1 U9133 ( .A1(n6957), .A2(n12717), .ZN(n6688) );
  AOI21_X1 U9134 ( .B1(n13804), .B2(n7324), .A(n7323), .ZN(n7322) );
  AND2_X1 U9135 ( .A1(n7465), .A2(n14493), .ZN(n6689) );
  AND2_X1 U9136 ( .A1(n12930), .A2(n12935), .ZN(n12934) );
  AND2_X1 U9137 ( .A1(n6987), .A2(n6986), .ZN(n6690) );
  NAND2_X1 U9138 ( .A1(n8166), .A2(n8165), .ZN(n13970) );
  INV_X1 U9139 ( .A(n13970), .ZN(n7165) );
  INV_X1 U9140 ( .A(n12925), .ZN(n7380) );
  INV_X1 U9141 ( .A(n14151), .ZN(n7539) );
  AND2_X1 U9142 ( .A1(n13079), .A2(n10379), .ZN(n6691) );
  AND4_X1 U9143 ( .A1(n8076), .A2(n8075), .A3(n8074), .A4(n8073), .ZN(n6692)
         );
  INV_X2 U9144 ( .A(n9371), .ZN(n9591) );
  NAND2_X2 U9145 ( .A1(n11490), .A2(n12137), .ZN(n8410) );
  OR2_X1 U9146 ( .A1(n15121), .A2(n14309), .ZN(n6693) );
  OR2_X1 U9147 ( .A1(n13914), .A2(n13893), .ZN(n6694) );
  AND3_X1 U9148 ( .A1(n9395), .A2(n9396), .A3(n9393), .ZN(n6695) );
  AND2_X1 U9149 ( .A1(n9177), .A2(n9176), .ZN(n6696) );
  AND2_X1 U9150 ( .A1(n7718), .A2(n7694), .ZN(n7720) );
  INV_X1 U9151 ( .A(n13656), .ZN(n7492) );
  OR2_X1 U9152 ( .A1(n8446), .A2(n8440), .ZN(n6697) );
  NAND2_X1 U9153 ( .A1(n8973), .A2(n8448), .ZN(n8976) );
  AND2_X1 U9154 ( .A1(n7537), .A2(n14096), .ZN(n6698) );
  OR3_X1 U9155 ( .A1(n8452), .A2(P3_IR_REG_1__SCAN_IN), .A3(
        P3_IR_REG_0__SCAN_IN), .ZN(n6699) );
  AND2_X1 U9156 ( .A1(n7554), .A2(n7552), .ZN(n6700) );
  AND2_X1 U9157 ( .A1(n7582), .A2(n13490), .ZN(n6701) );
  AND2_X1 U9158 ( .A1(n14668), .A2(n7507), .ZN(n6702) );
  AND2_X1 U9159 ( .A1(n13461), .A2(n13582), .ZN(n6703) );
  INV_X1 U9160 ( .A(n9174), .ZN(n7672) );
  NAND4_X1 U9161 ( .A1(n7756), .A2(n7755), .A3(n7754), .A4(n7753), .ZN(n9025)
         );
  AND2_X1 U9162 ( .A1(n9078), .A2(n9077), .ZN(n6704) );
  AND2_X1 U9163 ( .A1(n7426), .A2(n14355), .ZN(n6705) );
  INV_X1 U9164 ( .A(n11927), .ZN(n7517) );
  OR2_X1 U9165 ( .A1(n7132), .A2(n8445), .ZN(n6706) );
  AND4_X1 U9166 ( .A1(n8441), .A2(n8442), .A3(n7400), .A4(n8432), .ZN(n6707)
         );
  OR2_X1 U9167 ( .A1(n13986), .A2(n13638), .ZN(n6708) );
  AND2_X1 U9168 ( .A1(n8112), .A2(n6708), .ZN(n6709) );
  NAND2_X1 U9169 ( .A1(n12346), .A2(n7530), .ZN(n6710) );
  NAND2_X1 U9170 ( .A1(n14130), .A2(n12565), .ZN(n14140) );
  INV_X1 U9171 ( .A(n14433), .ZN(n7597) );
  AND2_X1 U9172 ( .A1(n9118), .A2(n9117), .ZN(n6711) );
  NOR2_X1 U9173 ( .A1(n13181), .A2(n13159), .ZN(n6712) );
  INV_X1 U9174 ( .A(n10995), .ZN(n7022) );
  AND2_X1 U9175 ( .A1(n11523), .A2(n11089), .ZN(n6713) );
  AND2_X1 U9176 ( .A1(n11594), .A2(n13651), .ZN(n6714) );
  INV_X1 U9177 ( .A(n8400), .ZN(n7312) );
  OR2_X1 U9178 ( .A1(n13541), .A2(n13536), .ZN(n8400) );
  NAND2_X2 U9179 ( .A1(n9394), .A2(n6695), .ZN(n14500) );
  INV_X1 U9180 ( .A(n14500), .ZN(n6811) );
  AND2_X1 U9181 ( .A1(n11526), .A2(n11087), .ZN(n6715) );
  AND2_X1 U9182 ( .A1(n15639), .A2(n12195), .ZN(n6716) );
  AND3_X1 U9183 ( .A1(n7713), .A2(n7714), .A3(n6881), .ZN(n6717) );
  OR2_X1 U9184 ( .A1(n9972), .A2(n9973), .ZN(n6718) );
  AND2_X1 U9185 ( .A1(n14053), .A2(n9160), .ZN(n6719) );
  INV_X1 U9186 ( .A(n14445), .ZN(n14669) );
  AND2_X1 U9187 ( .A1(n9349), .A2(n9348), .ZN(n14656) );
  INV_X1 U9188 ( .A(n14656), .ZN(n14793) );
  OR2_X1 U9189 ( .A1(n8446), .A2(P3_IR_REG_6__SCAN_IN), .ZN(n6720) );
  OR2_X1 U9190 ( .A1(n8465), .A2(n10929), .ZN(n6721) );
  OR2_X1 U9191 ( .A1(n13155), .A2(n13164), .ZN(n13156) );
  AND2_X1 U9192 ( .A1(n9376), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n6722) );
  NAND2_X1 U9193 ( .A1(n7977), .A2(n7976), .ZN(n12090) );
  NAND2_X1 U9194 ( .A1(n13118), .A2(n13127), .ZN(n6723) );
  OR2_X1 U9195 ( .A1(n13443), .A2(n9146), .ZN(n6724) );
  NAND2_X1 U9196 ( .A1(n9706), .A2(n9707), .ZN(n14381) );
  MUX2_X1 U9197 ( .A(n14487), .B(n14827), .S(n14335), .Z(n14341) );
  NAND2_X1 U9198 ( .A1(n12964), .A2(n12965), .ZN(n13126) );
  INV_X1 U9199 ( .A(n13126), .ZN(n13135) );
  AND2_X1 U9200 ( .A1(n6682), .A2(n6696), .ZN(n6725) );
  XNOR2_X1 U9201 ( .A(n13948), .B(n13631), .ZN(n13760) );
  INV_X1 U9202 ( .A(n11500), .ZN(n6911) );
  AND2_X1 U9203 ( .A1(n14326), .A2(n7156), .ZN(n6726) );
  AND2_X1 U9204 ( .A1(n9085), .A2(n9084), .ZN(n6727) );
  AND2_X1 U9205 ( .A1(n6951), .A2(n9874), .ZN(n6728) );
  AND2_X1 U9206 ( .A1(n12551), .A2(n12550), .ZN(n6729) );
  AND2_X1 U9207 ( .A1(n9122), .A2(n9121), .ZN(n6730) );
  OR2_X1 U9208 ( .A1(n13118), .A2(n9893), .ZN(n12839) );
  INV_X1 U9209 ( .A(n14690), .ZN(n14806) );
  AND2_X1 U9210 ( .A1(n9654), .A2(n9653), .ZN(n14690) );
  AND2_X1 U9211 ( .A1(n12934), .A2(n7378), .ZN(n6731) );
  XOR2_X1 U9212 ( .A(n14775), .B(n14478), .Z(n6732) );
  OR2_X1 U9213 ( .A1(n13385), .A2(n13149), .ZN(n6733) );
  INV_X1 U9214 ( .A(n7548), .ZN(n7547) );
  NAND2_X1 U9215 ( .A1(n12580), .A2(n7549), .ZN(n7548) );
  AND2_X1 U9216 ( .A1(n8210), .A2(n8209), .ZN(n14041) );
  INV_X1 U9217 ( .A(n14041), .ZN(n13797) );
  INV_X1 U9218 ( .A(n11893), .ZN(n7337) );
  AND2_X1 U9219 ( .A1(n13520), .A2(n6703), .ZN(n6734) );
  AND2_X1 U9220 ( .A1(n8636), .A2(n12894), .ZN(n6735) );
  NAND2_X1 U9221 ( .A1(n9838), .A2(n12438), .ZN(n6736) );
  INV_X1 U9222 ( .A(n14352), .ZN(n7421) );
  INV_X1 U9223 ( .A(n7166), .ZN(n13822) );
  NOR2_X1 U9224 ( .A1(n13841), .A2(n13970), .ZN(n7166) );
  NAND2_X1 U9225 ( .A1(n14224), .A2(n14502), .ZN(n6737) );
  AND2_X1 U9226 ( .A1(n7360), .A2(n9852), .ZN(n6738) );
  INV_X1 U9227 ( .A(n6947), .ZN(n6946) );
  OAI21_X1 U9228 ( .B1(n8315), .B2(n6750), .A(n6683), .ZN(n6947) );
  OR2_X1 U9229 ( .A1(n9047), .A2(n9046), .ZN(n6739) );
  AND2_X1 U9230 ( .A1(n14303), .A2(n14304), .ZN(n14437) );
  INV_X1 U9231 ( .A(n14437), .ZN(n9556) );
  OR2_X1 U9232 ( .A1(n6690), .A2(n9076), .ZN(n6740) );
  AND2_X1 U9233 ( .A1(n13859), .A2(n13579), .ZN(n6741) );
  INV_X1 U9234 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n7027) );
  AND2_X1 U9235 ( .A1(n15112), .A2(n14491), .ZN(n6742) );
  AND2_X1 U9236 ( .A1(n9640), .A2(n7151), .ZN(n6743) );
  OR2_X1 U9237 ( .A1(n14693), .A2(n9737), .ZN(n6744) );
  INV_X1 U9238 ( .A(n9247), .ZN(n9288) );
  NOR2_X1 U9239 ( .A1(n14917), .A2(n15108), .ZN(n6745) );
  NOR2_X1 U9240 ( .A1(n14053), .A2(n9160), .ZN(n6746) );
  NOR2_X1 U9241 ( .A1(n14041), .A2(n13633), .ZN(n6747) );
  NOR2_X1 U9242 ( .A1(n12582), .A2(n12581), .ZN(n6748) );
  INV_X1 U9243 ( .A(n7588), .ZN(n7587) );
  NAND2_X1 U9244 ( .A1(n14093), .A2(n14192), .ZN(n7588) );
  AND2_X1 U9245 ( .A1(n14332), .A2(n14331), .ZN(n14755) );
  INV_X1 U9246 ( .A(n14755), .ZN(n7610) );
  OR2_X1 U9247 ( .A1(n6719), .A2(n7333), .ZN(n6749) );
  INV_X1 U9248 ( .A(n7590), .ZN(n7589) );
  NOR2_X1 U9249 ( .A1(n14656), .A2(n14666), .ZN(n7590) );
  OR2_X1 U9250 ( .A1(n6949), .A2(n6948), .ZN(n6750) );
  AND2_X1 U9251 ( .A1(n9092), .A2(n9091), .ZN(n6751) );
  INV_X1 U9252 ( .A(n9423), .ZN(n7600) );
  AND2_X1 U9253 ( .A1(n11019), .A2(n11020), .ZN(n6752) );
  INV_X1 U9254 ( .A(n14306), .ZN(n7413) );
  NAND2_X1 U9255 ( .A1(n8433), .A2(n7357), .ZN(n6753) );
  NOR2_X1 U9256 ( .A1(n7418), .A2(n7419), .ZN(n6754) );
  NOR2_X1 U9257 ( .A1(n10362), .A2(n13112), .ZN(n6755) );
  NOR2_X1 U9258 ( .A1(n9836), .A2(n12373), .ZN(n6756) );
  NOR2_X1 U9259 ( .A1(n14093), .A2(n14481), .ZN(n6757) );
  NAND2_X1 U9260 ( .A1(n8433), .A2(n8432), .ZN(n6758) );
  AND2_X1 U9261 ( .A1(n12723), .A2(n12722), .ZN(n6759) );
  INV_X1 U9262 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n10441) );
  NAND2_X1 U9263 ( .A1(n13893), .A2(n13639), .ZN(n6760) );
  INV_X1 U9264 ( .A(n7964), .ZN(n7093) );
  OR2_X1 U9265 ( .A1(n14113), .A2(n7546), .ZN(n6761) );
  INV_X1 U9266 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n8680) );
  OR2_X1 U9267 ( .A1(n9604), .A2(n7154), .ZN(n6762) );
  NOR2_X1 U9268 ( .A1(n10736), .A2(n10735), .ZN(n6763) );
  NAND2_X1 U9269 ( .A1(P3_ADDR_REG_0__SCAN_IN), .A2(n9952), .ZN(n9951) );
  INV_X1 U9270 ( .A(n9951), .ZN(n6874) );
  OR2_X1 U9271 ( .A1(n8315), .A2(n6948), .ZN(n6764) );
  AND2_X1 U9272 ( .A1(n13295), .A2(n7621), .ZN(n6765) );
  NOR2_X1 U9273 ( .A1(n11697), .A2(n9815), .ZN(n6766) );
  AND2_X1 U9274 ( .A1(n14405), .A2(n14404), .ZN(n6767) );
  NOR2_X1 U9275 ( .A1(n13755), .A2(n14022), .ZN(n6768) );
  OR2_X1 U9276 ( .A1(n8446), .A2(n8445), .ZN(n6769) );
  AND2_X1 U9277 ( .A1(n7526), .A2(n7523), .ZN(n6770) );
  NOR2_X1 U9278 ( .A1(n14087), .A2(n12634), .ZN(n6771) );
  AND2_X1 U9279 ( .A1(n14369), .A2(n14368), .ZN(n6772) );
  AND2_X1 U9280 ( .A1(n13118), .A2(n9893), .ZN(n12837) );
  AND2_X1 U9281 ( .A1(n7800), .A2(n13653), .ZN(n6773) );
  OR2_X1 U9282 ( .A1(n14370), .A2(n14371), .ZN(n6774) );
  OR2_X1 U9283 ( .A1(n14265), .A2(n14263), .ZN(n6775) );
  OR2_X1 U9284 ( .A1(n14278), .A2(n14276), .ZN(n6776) );
  INV_X1 U9285 ( .A(n14369), .ZN(n14780) );
  NAND2_X1 U9286 ( .A1(n9679), .A2(n9678), .ZN(n14369) );
  AND2_X1 U9287 ( .A1(n8459), .A2(n8462), .ZN(n6777) );
  OR2_X1 U9288 ( .A1(n14251), .A2(n14253), .ZN(n6778) );
  AND2_X1 U9289 ( .A1(n7964), .A2(n7944), .ZN(n6779) );
  OR2_X1 U9290 ( .A1(n7086), .A2(n7084), .ZN(n6780) );
  AND2_X1 U9291 ( .A1(n7423), .A2(n7422), .ZN(n6781) );
  NAND2_X1 U9292 ( .A1(n13828), .A2(n13826), .ZN(n6922) );
  AND2_X1 U9293 ( .A1(n7357), .A2(n8434), .ZN(n6782) );
  AND2_X1 U9294 ( .A1(n7408), .A2(n14322), .ZN(n6783) );
  INV_X1 U9295 ( .A(n6893), .ZN(n6892) );
  NAND2_X1 U9296 ( .A1(n13563), .A2(n6894), .ZN(n6893) );
  OR2_X1 U9297 ( .A1(n7672), .A2(n7671), .ZN(n6784) );
  INV_X1 U9298 ( .A(n7482), .ZN(n7481) );
  NAND2_X1 U9299 ( .A1(n7483), .A2(n14303), .ZN(n7482) );
  NAND2_X1 U9300 ( .A1(n9550), .A2(n9549), .ZN(n12552) );
  INV_X1 U9301 ( .A(n12552), .ZN(n7512) );
  INV_X1 U9302 ( .A(n15557), .ZN(n11857) );
  INV_X1 U9303 ( .A(n12362), .ZN(n7622) );
  NAND2_X1 U9304 ( .A1(n8899), .A2(n8898), .ZN(n10362) );
  INV_X1 U9305 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n7491) );
  NAND2_X1 U9306 ( .A1(n8136), .A2(n11515), .ZN(n6785) );
  NAND2_X1 U9307 ( .A1(n8744), .A2(n12925), .ZN(n13249) );
  NAND2_X1 U9308 ( .A1(n12539), .A2(n12538), .ZN(n15101) );
  INV_X1 U9309 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n10212) );
  INV_X1 U9310 ( .A(n13965), .ZN(n7164) );
  AND4_X1 U9311 ( .A1(n8655), .A2(n8654), .A3(n8653), .A4(n8652), .ZN(n12372)
         );
  INV_X1 U9312 ( .A(n12933), .ZN(n7379) );
  NAND2_X1 U9313 ( .A1(n7128), .A2(n7378), .ZN(n13241) );
  INV_X1 U9314 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n7915) );
  OR2_X1 U9315 ( .A1(n12596), .A2(n12595), .ZN(n14095) );
  INV_X1 U9316 ( .A(n14095), .ZN(n7540) );
  AND2_X1 U9317 ( .A1(n9614), .A2(n9613), .ZN(n14336) );
  NOR2_X1 U9318 ( .A1(n15567), .A2(n12998), .ZN(n6786) );
  INV_X1 U9319 ( .A(n7175), .ZN(n13913) );
  AND2_X1 U9320 ( .A1(n10362), .A2(n10379), .ZN(n6787) );
  AND2_X1 U9321 ( .A1(n13079), .A2(n10382), .ZN(n6788) );
  OR2_X1 U9322 ( .A1(n13050), .A2(n8617), .ZN(n6789) );
  INV_X1 U9323 ( .A(n8323), .ZN(n7333) );
  NAND2_X1 U9324 ( .A1(n10354), .A2(n10353), .ZN(n13079) );
  AND2_X1 U9325 ( .A1(n8147), .A2(SI_21_), .ZN(n6790) );
  AND2_X1 U9326 ( .A1(n7607), .A2(n7609), .ZN(n6791) );
  AND2_X1 U9327 ( .A1(n14480), .A2(n14762), .ZN(n6792) );
  AND2_X1 U9328 ( .A1(n7332), .A2(n8323), .ZN(n6793) );
  INV_X1 U9329 ( .A(n15751), .ZN(n15749) );
  INV_X1 U9330 ( .A(n14487), .ZN(n7453) );
  AOI21_X1 U9331 ( .B1(n7460), .B2(n14431), .A(n6689), .ZN(n7458) );
  AND2_X1 U9332 ( .A1(n12067), .A2(n12066), .ZN(n6794) );
  AND2_X1 U9333 ( .A1(n8396), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n6795) );
  NAND2_X1 U9334 ( .A1(n11945), .A2(n8926), .ZN(n12030) );
  INV_X1 U9335 ( .A(n13048), .ZN(n15590) );
  AOI21_X1 U9336 ( .B1(n12218), .B2(n7370), .A(n7367), .ZN(n12434) );
  INV_X1 U9337 ( .A(n7519), .ZN(n11928) );
  AND2_X1 U9338 ( .A1(n11050), .A2(n11049), .ZN(n13591) );
  INV_X1 U9339 ( .A(n13591), .ZN(n13627) );
  OR2_X1 U9340 ( .A1(n9839), .A2(n13291), .ZN(n6796) );
  AND2_X1 U9341 ( .A1(n15625), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n6797) );
  INV_X1 U9342 ( .A(n14431), .ZN(n7463) );
  INV_X1 U9343 ( .A(n7460), .ZN(n7459) );
  INV_X1 U9344 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n7231) );
  OAI21_X1 U9345 ( .B1(n12046), .B2(n9830), .A(n9833), .ZN(n12176) );
  INV_X1 U9346 ( .A(n12176), .ZN(n6967) );
  OR2_X1 U9347 ( .A1(n7200), .A2(n7913), .ZN(n6798) );
  OAI21_X1 U9348 ( .B1(n7198), .B2(n6798), .A(n9218), .ZN(n7192) );
  INV_X1 U9349 ( .A(n12189), .ZN(n7633) );
  INV_X1 U9350 ( .A(n11662), .ZN(n7159) );
  NAND2_X1 U9351 ( .A1(n9479), .A2(n9478), .ZN(n14275) );
  INV_X1 U9352 ( .A(n14275), .ZN(n7465) );
  AND2_X2 U9353 ( .A1(n11098), .A2(n11097), .ZN(n15358) );
  OR2_X1 U9354 ( .A1(n9027), .A2(n8334), .ZN(n13906) );
  NAND2_X1 U9355 ( .A1(n9795), .A2(n9794), .ZN(n9801) );
  INV_X1 U9356 ( .A(n7199), .ZN(n7198) );
  NAND2_X1 U9357 ( .A1(n9217), .A2(n9215), .ZN(n7199) );
  OR2_X1 U9358 ( .A1(n15023), .A2(n13063), .ZN(n6799) );
  INV_X1 U9359 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n7717) );
  INV_X1 U9360 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n7716) );
  INV_X1 U9361 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n9901) );
  INV_X1 U9362 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n6968) );
  INV_X1 U9363 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n7402) );
  OR2_X1 U9364 ( .A1(n6805), .A2(n14297), .ZN(n7406) );
  OAI21_X1 U9365 ( .B1(n14225), .B2(n14227), .A(n14421), .ZN(n7438) );
  NAND2_X1 U9366 ( .A1(n6800), .A2(n6774), .ZN(n6846) );
  OR2_X2 U9367 ( .A1(n14366), .A2(n14367), .ZN(n6800) );
  NOR2_X1 U9368 ( .A1(n14358), .A2(n14359), .ZN(n6801) );
  AOI21_X1 U9369 ( .B1(n14357), .B2(n14356), .A(n6801), .ZN(n14362) );
  NAND2_X1 U9370 ( .A1(n6803), .A2(n6802), .ZN(n6806) );
  NAND2_X1 U9371 ( .A1(n14241), .A2(n14240), .ZN(n14244) );
  OAI21_X1 U9372 ( .B1(n7425), .B2(n7424), .A(n6781), .ZN(n14358) );
  OAI21_X1 U9373 ( .B1(n6846), .B2(n6845), .A(n7404), .ZN(n14406) );
  NAND2_X1 U9374 ( .A1(n14334), .A2(n14333), .ZN(n14340) );
  INV_X1 U9375 ( .A(n14296), .ZN(n6803) );
  OAI21_X1 U9376 ( .B1(n14327), .B2(n14326), .A(n14325), .ZN(n14328) );
  NAND2_X1 U9377 ( .A1(n14215), .A2(n14337), .ZN(n6837) );
  OAI211_X1 U9378 ( .C1(n12322), .C2(n7482), .A(n9736), .B(n7480), .ZN(n12449)
         );
  AOI22_X1 U9379 ( .A1(n12509), .A2(n12511), .B1(n14323), .B2(n14761), .ZN(
        n14754) );
  NOR2_X1 U9380 ( .A1(n14695), .A2(n14694), .ZN(n14693) );
  OAI21_X1 U9381 ( .B1(n7457), .B2(n11911), .A(n7456), .ZN(n9733) );
  NAND2_X1 U9382 ( .A1(n7466), .A2(n7467), .ZN(n12226) );
  NAND2_X1 U9383 ( .A1(n9715), .A2(n6807), .ZN(n11105) );
  NAND2_X1 U9384 ( .A1(n11207), .A2(n14422), .ZN(n11206) );
  AOI21_X1 U9385 ( .B1(n14634), .B2(n9740), .A(n6772), .ZN(n9741) );
  NAND2_X1 U9386 ( .A1(n11620), .A2(n14429), .ZN(n9728) );
  OAI22_X1 U9387 ( .A1(n12648), .A2(n10815), .B1(n11208), .B2(n10816), .ZN(
        n10817) );
  AOI21_X1 U9388 ( .B1(n7450), .B2(n7452), .A(n7447), .ZN(n14710) );
  AOI21_X2 U9389 ( .B1(n7519), .B2(n7517), .A(n11929), .ZN(n12123) );
  NAND2_X1 U9390 ( .A1(n6804), .A2(n15114), .ZN(n14092) );
  NAND2_X1 U9391 ( .A1(n7105), .A2(n14086), .ZN(n6804) );
  NAND2_X1 U9392 ( .A1(n6806), .A2(n7407), .ZN(n6805) );
  INV_X1 U9393 ( .A(n6812), .ZN(n11181) );
  NAND4_X1 U9394 ( .A1(n9374), .A2(n9375), .A3(n9372), .A4(n9373), .ZN(n6812)
         );
  OAI21_X2 U9395 ( .B1(n14505), .B2(n10730), .A(n11180), .ZN(n14219) );
  OAI21_X1 U9396 ( .B1(n14362), .B2(n14361), .A(n14360), .ZN(n14363) );
  NAND2_X1 U9397 ( .A1(n6812), .A2(n10730), .ZN(n11180) );
  AOI21_X1 U9398 ( .B1(n14296), .B2(n14295), .A(n14294), .ZN(n14297) );
  NAND2_X1 U9399 ( .A1(n9706), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9702) );
  INV_X2 U9400 ( .A(n14337), .ZN(n14229) );
  OAI21_X1 U9401 ( .B1(n14476), .B2(n14475), .A(n6809), .ZN(P1_U3242) );
  NAND2_X1 U9402 ( .A1(n6810), .A2(n14223), .ZN(n14226) );
  NAND2_X1 U9403 ( .A1(n14220), .A2(n14221), .ZN(n6810) );
  AOI21_X1 U9404 ( .B1(n14219), .B2(n14218), .A(n14217), .ZN(n14220) );
  OR2_X1 U9405 ( .A1(n9371), .A2(n7491), .ZN(n7510) );
  MUX2_X1 U9406 ( .A(n14224), .B(n14502), .S(n14337), .Z(n14225) );
  XNOR2_X1 U9407 ( .A(n6811), .B(n6672), .ZN(n14421) );
  NAND2_X1 U9408 ( .A1(n15207), .A2(n15208), .ZN(n15204) );
  INV_X1 U9409 ( .A(n15197), .ZN(n6819) );
  NAND2_X1 U9410 ( .A1(n9735), .A2(n14299), .ZN(n12322) );
  INV_X1 U9411 ( .A(n6838), .ZN(n14216) );
  AOI22_X1 U9412 ( .A1(n14710), .A2(n14709), .B1(n14718), .B2(n14344), .ZN(
        n14695) );
  NAND2_X1 U9413 ( .A1(n14647), .A2(n7015), .ZN(n6813) );
  NAND2_X1 U9414 ( .A1(n6816), .A2(n7566), .ZN(n13544) );
  NAND2_X1 U9415 ( .A1(n7565), .A2(n7681), .ZN(n6816) );
  INV_X4 U9416 ( .A(n8524), .ZN(n11984) );
  NAND2_X1 U9417 ( .A1(n13125), .A2(n13126), .ZN(n13124) );
  NAND2_X1 U9418 ( .A1(n6931), .A2(n6932), .ZN(n6930) );
  NAND2_X1 U9419 ( .A1(n8026), .A2(n8025), .ZN(n8044) );
  OAI21_X1 U9420 ( .B1(n15040), .B2(n7640), .A(n7639), .ZN(n12370) );
  NOR2_X1 U9421 ( .A1(n7118), .A2(n13101), .ZN(n9021) );
  NOR2_X1 U9422 ( .A1(n13231), .A2(n12934), .ZN(n7069) );
  INV_X1 U9423 ( .A(n15217), .ZN(n6826) );
  NAND2_X1 U9424 ( .A1(n9985), .A2(P2_ADDR_REG_16__SCAN_IN), .ZN(n6825) );
  NAND2_X1 U9425 ( .A1(n11261), .A2(n11262), .ZN(n7560) );
  NAND2_X2 U9426 ( .A1(n12467), .A2(n12466), .ZN(n12469) );
  AOI21_X1 U9427 ( .B1(n13455), .B2(n13454), .A(n7676), .ZN(n13519) );
  NAND2_X1 U9428 ( .A1(n12034), .A2(n12889), .ZN(n12187) );
  NAND2_X1 U9429 ( .A1(n13165), .A2(n13164), .ZN(n13167) );
  NAND2_X1 U9430 ( .A1(n7383), .A2(n7384), .ZN(n12363) );
  OAI21_X1 U9431 ( .B1(n13296), .B2(n7398), .A(n12916), .ZN(n13281) );
  AOI21_X1 U9432 ( .B1(n13141), .B2(n7122), .A(n7120), .ZN(n7119) );
  NOR2_X1 U9433 ( .A1(n11164), .A2(n8563), .ZN(n11323) );
  NOR2_X1 U9434 ( .A1(n15552), .A2(n15551), .ZN(n15550) );
  NAND2_X1 U9435 ( .A1(n10959), .A2(n7301), .ZN(n7300) );
  NAND2_X1 U9436 ( .A1(n11303), .A2(n10913), .ZN(n10960) );
  INV_X1 U9437 ( .A(n11301), .ZN(n6867) );
  NAND2_X1 U9438 ( .A1(n14236), .A2(n14237), .ZN(n14235) );
  NAND2_X1 U9439 ( .A1(n6836), .A2(n14232), .ZN(n14236) );
  INV_X1 U9440 ( .A(n14453), .ZN(n14470) );
  NAND2_X1 U9441 ( .A1(n14406), .A2(n6767), .ZN(n14453) );
  NAND2_X1 U9442 ( .A1(n9320), .A2(n7557), .ZN(n7559) );
  NAND2_X1 U9443 ( .A1(n9701), .A2(n6685), .ZN(n9706) );
  NAND2_X1 U9444 ( .A1(n14363), .A2(n7401), .ZN(n14366) );
  MUX2_X2 U9445 ( .A(n14213), .B(n14381), .S(n14382), .Z(n14337) );
  OAI21_X1 U9446 ( .B1(n6838), .B2(n14337), .A(n6837), .ZN(n14221) );
  NAND2_X1 U9447 ( .A1(n8015), .A2(n8014), .ZN(n8026) );
  NAND2_X1 U9448 ( .A1(n7868), .A2(n7217), .ZN(n7006) );
  NAND2_X1 U9449 ( .A1(n6824), .A2(n7439), .ZN(n6836) );
  NAND2_X1 U9450 ( .A1(n14226), .A2(n7440), .ZN(n6824) );
  NAND2_X2 U9451 ( .A1(n15206), .A2(n15204), .ZN(n15210) );
  NOR2_X2 U9452 ( .A1(n14964), .A2(n14965), .ZN(n14963) );
  AND2_X2 U9453 ( .A1(n6826), .A2(n6825), .ZN(n14964) );
  NAND2_X1 U9454 ( .A1(n6850), .A2(n6849), .ZN(n6873) );
  NAND2_X1 U9455 ( .A1(n7074), .A2(n7717), .ZN(n7073) );
  NAND2_X1 U9456 ( .A1(n7007), .A2(n8008), .ZN(n8015) );
  NAND4_X1 U9457 ( .A1(n6732), .A2(n6829), .A3(n14447), .A4(n14448), .ZN(n6828) );
  NAND2_X1 U9458 ( .A1(n7006), .A2(n7219), .ZN(n7005) );
  NAND2_X1 U9459 ( .A1(n7852), .A2(n7851), .ZN(n7868) );
  NAND2_X1 U9460 ( .A1(n13611), .A2(n13497), .ZN(n13535) );
  NAND2_X1 U9461 ( .A1(n7322), .A2(n6922), .ZN(n6918) );
  INV_X2 U9462 ( .A(n13537), .ZN(n13498) );
  NAND2_X4 U9463 ( .A1(n11052), .A2(n9029), .ZN(n13537) );
  AOI21_X1 U9464 ( .B1(n13738), .B2(n15491), .A(n8412), .ZN(n8420) );
  NAND3_X1 U9465 ( .A1(n13512), .A2(n11274), .A3(n11273), .ZN(n11412) );
  NAND2_X1 U9466 ( .A1(n11792), .A2(n8925), .ZN(n11946) );
  OAI21_X1 U9467 ( .B1(n10380), .B2(n15749), .A(n6831), .ZN(P3_U3488) );
  OAI21_X1 U9468 ( .B1(n10380), .B2(n15743), .A(n6833), .ZN(P3_U3456) );
  NAND2_X1 U9469 ( .A1(n7625), .A2(n7624), .ZN(n15638) );
  NOR2_X1 U9470 ( .A1(n13089), .A2(n13090), .ZN(n13088) );
  NAND2_X1 U9471 ( .A1(n8952), .A2(n7069), .ZN(n7068) );
  MUX2_X2 U9472 ( .A(n13940), .B(n14023), .S(n15539), .Z(n13941) );
  OR2_X1 U9473 ( .A1(n11085), .A2(n11400), .ZN(n11518) );
  OR2_X2 U9474 ( .A1(n13932), .A2(n11053), .ZN(n10855) );
  AND2_X2 U9475 ( .A1(n13776), .A2(n13766), .ZN(n13763) );
  NOR2_X2 U9476 ( .A1(n6835), .A2(n13841), .ZN(n13776) );
  XOR2_X1 U9477 ( .A(n13731), .B(n13729), .Z(n7170) );
  NAND2_X1 U9478 ( .A1(n7406), .A2(n6783), .ZN(n14327) );
  NAND2_X1 U9479 ( .A1(n14287), .A2(n14286), .ZN(n14288) );
  OAI21_X1 U9480 ( .B1(n14470), .B2(n14469), .A(n7687), .ZN(n6848) );
  NOR2_X2 U9481 ( .A1(n6840), .A2(n9309), .ZN(n9558) );
  NAND4_X1 U9482 ( .A1(n9308), .A2(n9307), .A3(n10298), .A4(n10191), .ZN(n6840) );
  INV_X2 U9483 ( .A(n14503), .ZN(n11208) );
  NAND2_X1 U9484 ( .A1(n6842), .A2(n7436), .ZN(n14256) );
  NAND3_X1 U9485 ( .A1(n14249), .A2(n14248), .A3(n6778), .ZN(n6842) );
  NAND2_X1 U9486 ( .A1(n6843), .A2(n7414), .ZN(n14269) );
  NAND3_X1 U9487 ( .A1(n14261), .A2(n14260), .A3(n6775), .ZN(n6843) );
  NAND2_X1 U9488 ( .A1(n6844), .A2(n7434), .ZN(n14282) );
  NAND3_X1 U9489 ( .A1(n14274), .A2(n14273), .A3(n6776), .ZN(n6844) );
  NAND2_X2 U9490 ( .A1(n9391), .A2(n9390), .ZN(n14228) );
  NOR2_X1 U9491 ( .A1(n6768), .A2(n7689), .ZN(n6925) );
  NAND3_X1 U9492 ( .A1(n7824), .A2(n7504), .A3(n7077), .ZN(n7080) );
  OAI21_X1 U9493 ( .B1(n14030), .B2(n15536), .A(n6923), .ZN(n8387) );
  NAND2_X1 U9494 ( .A1(n8390), .A2(n8273), .ZN(n13755) );
  NOR2_X1 U9495 ( .A1(n6848), .A2(n14471), .ZN(n14476) );
  XNOR2_X1 U9496 ( .A(n11400), .B(n13654), .ZN(n11087) );
  NAND2_X1 U9497 ( .A1(n6873), .A2(n14894), .ZN(n6860) );
  INV_X1 U9498 ( .A(n14896), .ZN(n6850) );
  AND2_X2 U9499 ( .A1(n9703), .A2(n9770), .ZN(n9742) );
  NAND2_X2 U9500 ( .A1(n12598), .A2(n14171), .ZN(n14094) );
  OR2_X4 U9501 ( .A1(n14132), .A2(n14133), .ZN(n14130) );
  NAND2_X1 U9502 ( .A1(n14187), .A2(n6771), .ZN(n7105) );
  OAI21_X1 U9503 ( .B1(n14347), .B2(n14346), .A(n14345), .ZN(n14348) );
  NAND2_X1 U9504 ( .A1(n6963), .A2(n6962), .ZN(n8461) );
  NAND2_X1 U9505 ( .A1(n7070), .A2(n7068), .ZN(n13155) );
  NAND2_X1 U9506 ( .A1(n7618), .A2(n6765), .ZN(n13289) );
  INV_X1 U9507 ( .A(n12370), .ZN(n8931) );
  NAND2_X1 U9508 ( .A1(n12779), .A2(n6958), .ZN(n12702) );
  NAND2_X1 U9509 ( .A1(n7363), .A2(n7361), .ZN(n12732) );
  NAND2_X1 U9510 ( .A1(n12711), .A2(n9855), .ZN(n9857) );
  NAND2_X1 U9511 ( .A1(n7346), .A2(n7345), .ZN(n7344) );
  INV_X1 U9512 ( .A(n9807), .ZN(n6853) );
  NAND2_X1 U9513 ( .A1(n12177), .A2(n12372), .ZN(n6966) );
  OAI21_X1 U9514 ( .B1(n7784), .B2(n7787), .A(n7214), .ZN(n7816) );
  NAND2_X1 U9515 ( .A1(n6881), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n6880) );
  NOR2_X1 U9516 ( .A1(n9962), .A2(n9961), .ZN(n9910) );
  NOR2_X2 U9517 ( .A1(n6858), .A2(n6855), .ZN(n14788) );
  AOI21_X2 U9518 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(n9986), .A(n14963), .ZN(
        n14896) );
  NAND2_X1 U9519 ( .A1(n14362), .A2(n14361), .ZN(n7401) );
  INV_X1 U9520 ( .A(n14351), .ZN(n7425) );
  XNOR2_X1 U9521 ( .A(n6860), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(SUB_1596_U62)
         );
  NAND2_X1 U9522 ( .A1(n15556), .A2(n15553), .ZN(n11859) );
  NAND2_X1 U9523 ( .A1(n11855), .A2(n11856), .ZN(n15556) );
  OAI211_X1 U9524 ( .C1(n7034), .C2(n15541), .A(n7033), .B(n7032), .ZN(n7031)
         );
  INV_X1 U9525 ( .A(n7031), .ZN(n13066) );
  NAND2_X1 U9526 ( .A1(n15439), .A2(n15438), .ZN(n15437) );
  NAND2_X1 U9527 ( .A1(n15760), .A2(n15761), .ZN(n15759) );
  NAND2_X1 U9528 ( .A1(n6866), .A2(P2_ADDR_REG_11__SCAN_IN), .ZN(n7181) );
  NAND2_X1 U9529 ( .A1(n15197), .A2(n15198), .ZN(n6866) );
  INV_X1 U9530 ( .A(n15214), .ZN(n6870) );
  INV_X1 U9531 ( .A(n9958), .ZN(n6871) );
  NOR2_X1 U9532 ( .A1(n10939), .A2(n10938), .ZN(n10976) );
  XNOR2_X1 U9533 ( .A(n11320), .B(n11321), .ZN(n11164) );
  NAND2_X1 U9534 ( .A1(n7473), .A2(n7472), .ZN(P1_U3557) );
  OAI211_X1 U9535 ( .C1(n10390), .C2(n15155), .A(n9754), .B(n10402), .ZN(
        n14776) );
  NOR2_X1 U9536 ( .A1(n9946), .A2(P1_ADDR_REG_3__SCAN_IN), .ZN(n9904) );
  XNOR2_X2 U9537 ( .A(n9902), .B(n10195), .ZN(n9946) );
  INV_X1 U9538 ( .A(n9949), .ZN(n6875) );
  NAND2_X1 U9539 ( .A1(n15214), .A2(n15215), .ZN(n7203) );
  NAND2_X1 U9540 ( .A1(n7203), .A2(P2_ADDR_REG_15__SCAN_IN), .ZN(n7202) );
  XNOR2_X1 U9541 ( .A(n9953), .B(n9950), .ZN(n15767) );
  XNOR2_X1 U9542 ( .A(n9949), .B(n6874), .ZN(n9953) );
  OR2_X1 U9543 ( .A1(n9948), .A2(n9947), .ZN(n7225) );
  NAND2_X1 U9544 ( .A1(n7229), .A2(n14894), .ZN(n7228) );
  XNOR2_X1 U9545 ( .A(n7228), .B(n7227), .ZN(SUB_1596_U4) );
  NAND3_X1 U9546 ( .A1(n6877), .A2(n6876), .A3(P2_ADDR_REG_19__SCAN_IN), .ZN(
        n7004) );
  INV_X1 U9547 ( .A(n10433), .ZN(n6881) );
  NAND2_X1 U9548 ( .A1(n6880), .A2(n7071), .ZN(n6879) );
  NAND3_X1 U9549 ( .A1(n6880), .A2(n7071), .A3(n6886), .ZN(n6885) );
  AND2_X1 U9550 ( .A1(n6883), .A2(n6882), .ZN(n7739) );
  AOI21_X1 U9551 ( .B1(n10433), .B2(n8464), .A(n10454), .ZN(n6882) );
  INV_X1 U9552 ( .A(n10433), .ZN(n6884) );
  INV_X1 U9553 ( .A(SI_1_), .ZN(n6886) );
  NAND2_X1 U9554 ( .A1(n6887), .A2(n6889), .ZN(n13600) );
  NAND2_X1 U9555 ( .A1(n12388), .A2(n6901), .ZN(n6900) );
  NAND2_X1 U9556 ( .A1(n11507), .A2(n6909), .ZN(n6908) );
  NAND2_X1 U9557 ( .A1(n7848), .A2(n7847), .ZN(n7852) );
  NAND2_X1 U9558 ( .A1(n13838), .A2(n6919), .ZN(n6916) );
  NAND2_X1 U9559 ( .A1(n6917), .A2(n6916), .ZN(n13773) );
  INV_X1 U9560 ( .A(n7322), .ZN(n6920) );
  INV_X1 U9561 ( .A(n6922), .ZN(n6921) );
  NAND2_X1 U9562 ( .A1(n13554), .A2(n6929), .ZN(n6927) );
  NAND2_X1 U9563 ( .A1(n13554), .A2(n6935), .ZN(n6928) );
  OAI211_X1 U9564 ( .C1(n13554), .C2(n6930), .A(n13591), .B(n6927), .ZN(n7565)
         );
  NAND2_X1 U9565 ( .A1(n13554), .A2(n13553), .ZN(n13491) );
  NAND2_X1 U9566 ( .A1(n12721), .A2(n9869), .ZN(n6957) );
  INV_X1 U9567 ( .A(n7395), .ZN(n6964) );
  NAND3_X1 U9568 ( .A1(n6707), .A2(n8533), .A3(n7395), .ZN(n6959) );
  NAND3_X1 U9569 ( .A1(n8443), .A2(n6961), .A3(n8444), .ZN(n6960) );
  AND2_X2 U9570 ( .A1(n6967), .A2(n6966), .ZN(n12218) );
  NAND2_X2 U9571 ( .A1(n8453), .A2(n12684), .ZN(n8524) );
  INV_X1 U9572 ( .A(n9079), .ZN(n6972) );
  INV_X1 U9573 ( .A(n9179), .ZN(n6979) );
  NAND4_X1 U9574 ( .A1(n6983), .A2(n6982), .A3(n7651), .A4(n6981), .ZN(n6980)
         );
  NAND2_X1 U9575 ( .A1(n6696), .A2(n9179), .ZN(n6981) );
  NAND2_X1 U9576 ( .A1(n9169), .A2(n6725), .ZN(n6982) );
  NAND2_X1 U9577 ( .A1(n7670), .A2(n6725), .ZN(n6983) );
  NAND2_X1 U9578 ( .A1(n9169), .A2(n6682), .ZN(n6984) );
  NAND2_X1 U9579 ( .A1(n7670), .A2(n6682), .ZN(n6985) );
  OAI21_X1 U9580 ( .B1(n9090), .B2(n6991), .A(n6990), .ZN(n9097) );
  NAND2_X1 U9581 ( .A1(n6989), .A2(n6988), .ZN(n9096) );
  NAND2_X1 U9582 ( .A1(n9090), .A2(n6990), .ZN(n6989) );
  NAND2_X1 U9583 ( .A1(n9126), .A2(n6995), .ZN(n6993) );
  NAND2_X1 U9584 ( .A1(n9127), .A2(n6996), .ZN(n6994) );
  NAND3_X1 U9585 ( .A1(n6994), .A2(n6993), .A3(n6998), .ZN(n9163) );
  NAND4_X1 U9586 ( .A1(n6994), .A2(n6993), .A3(n6998), .A4(n6992), .ZN(n6997)
         );
  NAND2_X1 U9587 ( .A1(n6997), .A2(n9161), .ZN(n9165) );
  INV_X1 U9588 ( .A(n9138), .ZN(n6999) );
  NAND2_X2 U9589 ( .A1(n8282), .A2(n7000), .ZN(n7714) );
  NAND3_X1 U9590 ( .A1(n9253), .A2(n7663), .A3(n9230), .ZN(n7003) );
  NAND2_X1 U9591 ( .A1(n7004), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n7072) );
  NAND2_X1 U9592 ( .A1(n7994), .A2(n7206), .ZN(n7007) );
  NAND2_X1 U9593 ( .A1(n7993), .A2(SI_14_), .ZN(n7994) );
  NAND3_X1 U9594 ( .A1(n7027), .A2(P3_IR_REG_31__SCAN_IN), .A3(
        P3_IR_REG_1__SCAN_IN), .ZN(n7024) );
  NAND3_X1 U9595 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(n7027), .A3(
        P3_IR_REG_31__SCAN_IN), .ZN(n7026) );
  NAND2_X1 U9596 ( .A1(n8519), .A2(n7044), .ZN(n7041) );
  NAND2_X1 U9597 ( .A1(n7041), .A2(n7042), .ZN(n8555) );
  NOR2_X1 U9598 ( .A1(n13075), .A2(n7054), .ZN(n10380) );
  NAND2_X1 U9599 ( .A1(n7056), .A2(n15703), .ZN(n7055) );
  XNOR2_X1 U9600 ( .A(n10365), .B(n10364), .ZN(n7056) );
  OAI22_X1 U9601 ( .A1(n7064), .A2(n13188), .B1(n8945), .B2(n8944), .ZN(n8950)
         );
  INV_X1 U9602 ( .A(n13193), .ZN(n13196) );
  NOR2_X1 U9603 ( .A1(n13193), .A2(n7066), .ZN(n13173) );
  NAND3_X1 U9604 ( .A1(n7716), .A2(n7715), .A3(P3_ADDR_REG_19__SCAN_IN), .ZN(
        n7074) );
  NAND2_X1 U9605 ( .A1(n10852), .A2(n7075), .ZN(n10854) );
  XNOR2_X1 U9606 ( .A(n11129), .B(n13656), .ZN(n10858) );
  INV_X1 U9607 ( .A(n10852), .ZN(n7076) );
  NAND2_X1 U9608 ( .A1(n7080), .A2(n7078), .ZN(n11639) );
  NAND3_X1 U9609 ( .A1(n7824), .A2(n9272), .A3(n7504), .ZN(n11575) );
  NAND2_X1 U9610 ( .A1(n8113), .A2(n7085), .ZN(n7083) );
  NAND2_X1 U9611 ( .A1(n7083), .A2(n6780), .ZN(n13849) );
  NAND2_X1 U9612 ( .A1(n11891), .A2(n6779), .ZN(n7089) );
  NAND2_X1 U9613 ( .A1(n11891), .A2(n7944), .ZN(n7096) );
  NAND2_X1 U9614 ( .A1(n7089), .A2(n7091), .ZN(n7986) );
  NAND2_X2 U9615 ( .A1(n7099), .A2(n7098), .ZN(n14111) );
  OAI21_X1 U9616 ( .B1(n14130), .B2(n7551), .A(n7547), .ZN(n14105) );
  NAND2_X1 U9617 ( .A1(n9701), .A2(n7112), .ZN(n9770) );
  NAND2_X1 U9618 ( .A1(n9701), .A2(n9700), .ZN(n9704) );
  INV_X1 U9619 ( .A(n7119), .ZN(n7392) );
  NAND2_X1 U9620 ( .A1(n12021), .A2(n7124), .ZN(n12864) );
  INV_X1 U9621 ( .A(n15681), .ZN(n7124) );
  XNOR2_X1 U9622 ( .A(n12021), .B(n7125), .ZN(n9805) );
  OAI22_X1 U9623 ( .A1(n13424), .A2(n7126), .B1(n15741), .B2(n8494), .ZN(
        n11377) );
  OAI22_X1 U9624 ( .A1(n13367), .A2(n7126), .B1(n15751), .B2(n11379), .ZN(
        n11380) );
  NAND2_X1 U9625 ( .A1(n7131), .A2(n7130), .ZN(n7132) );
  OAI21_X2 U9626 ( .B1(n12363), .B2(n7133), .A(n12911), .ZN(n13296) );
  INV_X1 U9627 ( .A(n9755), .ZN(n7134) );
  NAND2_X1 U9628 ( .A1(n7136), .A2(n7138), .ZN(n9530) );
  NAND2_X1 U9629 ( .A1(n9487), .A2(n7139), .ZN(n7136) );
  NAND2_X1 U9630 ( .A1(n9408), .A2(n7142), .ZN(n7143) );
  INV_X1 U9631 ( .A(n14728), .ZN(n7148) );
  OAI21_X1 U9632 ( .B1(n7148), .B2(n7150), .A(n7149), .ZN(n14705) );
  XNOR2_X2 U9633 ( .A(n7403), .B(P1_IR_REG_30__SCAN_IN), .ZN(n9324) );
  NOR2_X2 U9634 ( .A1(n11636), .A2(n11755), .ZN(n11776) );
  INV_X1 U9635 ( .A(n11635), .ZN(n7160) );
  AND2_X2 U9636 ( .A1(n11583), .A2(n15482), .ZN(n11593) );
  NAND2_X1 U9637 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n8283), .ZN(n7710) );
  NAND2_X1 U9638 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n7744) );
  OAI22_X1 U9639 ( .A1(n7708), .A2(P2_IR_REG_31__SCAN_IN), .B1(n7707), .B2(
        n14065), .ZN(n7712) );
  NAND2_X1 U9640 ( .A1(n7819), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7792) );
  NAND2_X1 U9641 ( .A1(n7972), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7973) );
  NAND2_X1 U9642 ( .A1(n8077), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7951) );
  NAND2_X1 U9643 ( .A1(n8080), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8078) );
  OAI21_X1 U9644 ( .B1(n8277), .B2(P2_IR_REG_19__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8279) );
  NAND2_X1 U9645 ( .A1(n7726), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7725) );
  NAND2_X1 U9646 ( .A1(n7995), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7996) );
  NAND2_X1 U9647 ( .A1(n8282), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8281) );
  NAND2_X1 U9648 ( .A1(n8052), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8030) );
  OAI21_X1 U9649 ( .B1(n8052), .B2(n8051), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n8053) );
  NAND2_X1 U9650 ( .A1(n8031), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8032) );
  NAND2_X1 U9651 ( .A1(n8381), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8382) );
  NAND2_X1 U9652 ( .A1(n8345), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8407) );
  NAND2_X1 U9653 ( .A1(n7932), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7917) );
  OAI21_X1 U9654 ( .B1(n7932), .B2(P2_IR_REG_10__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n7933) );
  NOR2_X2 U9655 ( .A1(n12263), .A2(n12310), .ZN(n12392) );
  NOR2_X2 U9656 ( .A1(n6694), .A2(n13986), .ZN(n13882) );
  NOR2_X2 U9657 ( .A1(n12427), .A2(n13443), .ZN(n7175) );
  NAND2_X1 U9658 ( .A1(n15202), .A2(n15201), .ZN(n15200) );
  INV_X1 U9659 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7180) );
  AND2_X2 U9660 ( .A1(n7182), .A2(n7181), .ZN(n15202) );
  NAND3_X1 U9661 ( .A1(n7193), .A2(n7194), .A3(n7187), .ZN(n14875) );
  NAND2_X1 U9662 ( .A1(n9233), .A2(n7195), .ZN(n7193) );
  NOR2_X1 U9663 ( .A1(n7913), .A2(n7190), .ZN(n7189) );
  AND2_X2 U9664 ( .A1(n7202), .A2(n7201), .ZN(n15219) );
  OAI21_X1 U9665 ( .B1(n7911), .B2(n7212), .A(n7210), .ZN(n7966) );
  NAND2_X1 U9666 ( .A1(n7209), .A2(n7207), .ZN(n7970) );
  NAND2_X1 U9667 ( .A1(n7911), .A2(n7210), .ZN(n7209) );
  AOI21_X1 U9668 ( .B1(n7788), .B2(n7216), .A(n7215), .ZN(n7214) );
  INV_X1 U9669 ( .A(n7783), .ZN(n7216) );
  NAND2_X1 U9670 ( .A1(n7789), .A2(n7788), .ZN(n7812) );
  NAND2_X1 U9671 ( .A1(n7784), .A2(n7783), .ZN(n7789) );
  OAI21_X2 U9672 ( .B1(n7769), .B2(n7768), .A(n7767), .ZN(n7784) );
  AND2_X2 U9673 ( .A1(n7225), .A2(n7224), .ZN(n9902) );
  NOR2_X2 U9674 ( .A1(n9904), .A2(n9903), .ZN(n9905) );
  NAND2_X1 U9675 ( .A1(n8259), .A2(n7236), .ZN(n7232) );
  NAND2_X1 U9676 ( .A1(n8259), .A2(n8258), .ZN(n8392) );
  NOR2_X1 U9677 ( .A1(n6722), .A2(n8486), .ZN(n10455) );
  XNOR2_X1 U9678 ( .A(n7238), .B(n8486), .ZN(n10444) );
  INV_X1 U9679 ( .A(n8487), .ZN(n7238) );
  NAND3_X1 U9680 ( .A1(n7245), .A2(n7243), .A3(n7239), .ZN(n12984) );
  NAND3_X1 U9681 ( .A1(n12816), .A2(n12817), .A3(n7242), .ZN(n7241) );
  NAND2_X1 U9682 ( .A1(n7246), .A2(n7244), .ZN(n7243) );
  NAND2_X1 U9683 ( .A1(n7248), .A2(n12817), .ZN(n7247) );
  NAND2_X1 U9684 ( .A1(n7250), .A2(n7249), .ZN(n7248) );
  INV_X1 U9685 ( .A(n12977), .ZN(n7249) );
  NAND2_X1 U9686 ( .A1(n12978), .A2(n12979), .ZN(n7250) );
  NAND2_X1 U9687 ( .A1(n8713), .A2(n7254), .ZN(n7253) );
  NAND2_X1 U9688 ( .A1(n8768), .A2(n7260), .ZN(n7259) );
  INV_X1 U9689 ( .A(n8677), .ZN(n7273) );
  NAND3_X1 U9690 ( .A1(n12967), .A2(n12966), .A3(n7277), .ZN(n7276) );
  INV_X1 U9691 ( .A(n7280), .ZN(n7279) );
  NAND2_X1 U9692 ( .A1(n8864), .A2(n8852), .ZN(n8853) );
  INV_X1 U9693 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7281) );
  NAND2_X1 U9694 ( .A1(n8806), .A2(n8805), .ZN(n8809) );
  INV_X1 U9695 ( .A(n8808), .ZN(n7285) );
  NAND2_X1 U9696 ( .A1(n8881), .A2(n8880), .ZN(n8893) );
  NAND2_X1 U9697 ( .A1(n8850), .A2(n8849), .ZN(n8851) );
  NAND2_X1 U9698 ( .A1(n8072), .A2(n8071), .ZN(n8117) );
  INV_X1 U9699 ( .A(n9246), .ZN(n9248) );
  NOR2_X1 U9700 ( .A1(n7327), .A2(n8855), .ZN(n7326) );
  NOR2_X2 U9701 ( .A1(n11518), .A2(n11523), .ZN(n11583) );
  NOR2_X1 U9702 ( .A1(n10915), .A2(n12018), .ZN(n10935) );
  NAND2_X1 U9703 ( .A1(n7970), .A2(n7969), .ZN(n7992) );
  NAND2_X1 U9704 ( .A1(n8117), .A2(n8116), .ZN(n8124) );
  NOR2_X1 U9705 ( .A1(n11845), .A2(n11844), .ZN(n12996) );
  NAND2_X1 U9706 ( .A1(n10352), .A2(n10351), .ZN(n12687) );
  NAND2_X1 U9707 ( .A1(n8847), .A2(n8846), .ZN(n8850) );
  NAND2_X1 U9708 ( .A1(n8803), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n8806) );
  NAND2_X1 U9709 ( .A1(n12808), .A2(n12807), .ZN(n12812) );
  NAND2_X1 U9710 ( .A1(n8046), .A2(n8045), .ZN(n8070) );
  NAND4_X1 U9711 ( .A1(n7695), .A2(n7915), .A3(n7302), .A4(n7891), .ZN(n7655)
         );
  NAND3_X1 U9712 ( .A1(n7308), .A2(n7309), .A3(n7307), .ZN(n8412) );
  NAND2_X1 U9713 ( .A1(n7306), .A2(n7305), .ZN(n7309) );
  INV_X1 U9714 ( .A(n8401), .ZN(n7305) );
  AND2_X1 U9715 ( .A1(n7310), .A2(n13906), .ZN(n7306) );
  NAND2_X1 U9716 ( .A1(n13873), .A2(n7316), .ZN(n7315) );
  NOR2_X1 U9717 ( .A1(n7692), .A2(n7325), .ZN(n7745) );
  NOR2_X1 U9718 ( .A1(n7913), .A2(n10466), .ZN(n7325) );
  NAND2_X1 U9719 ( .A1(n11088), .A2(n6715), .ZN(n7328) );
  NOR2_X1 U9720 ( .A1(n11774), .A2(n7339), .ZN(n7338) );
  NAND3_X1 U9721 ( .A1(n7568), .A2(n7652), .A3(n6677), .ZN(n7972) );
  AND4_X2 U9722 ( .A1(n7568), .A2(n7652), .A3(n6677), .A4(n7340), .ZN(n7974)
         );
  NOR2_X1 U9723 ( .A1(n9797), .A2(n9801), .ZN(n11028) );
  INV_X1 U9724 ( .A(n9801), .ZN(n7341) );
  INV_X1 U9725 ( .A(n9797), .ZN(n7342) );
  INV_X1 U9726 ( .A(n9862), .ZN(n7346) );
  NAND3_X1 U9727 ( .A1(n12747), .A2(n13178), .A3(n7344), .ZN(n12694) );
  AND3_X2 U9728 ( .A1(n7348), .A2(n7347), .A3(n8426), .ZN(n8533) );
  NAND3_X1 U9729 ( .A1(n7349), .A2(n8426), .A3(n7030), .ZN(n8514) );
  INV_X2 U9730 ( .A(n9791), .ZN(n9870) );
  NAND2_X1 U9731 ( .A1(n8433), .A2(n6782), .ZN(n8910) );
  NAND2_X1 U9732 ( .A1(n12218), .A2(n7364), .ZN(n7363) );
  NAND3_X1 U9733 ( .A1(n7382), .A2(n12863), .A3(n7381), .ZN(n11559) );
  NAND3_X1 U9734 ( .A1(n12864), .A2(n12854), .A3(n12853), .ZN(n7382) );
  NAND2_X1 U9735 ( .A1(n11369), .A2(n12864), .ZN(n11560) );
  NAND2_X1 U9736 ( .A1(n11370), .A2(n12821), .ZN(n11369) );
  INV_X1 U9737 ( .A(n11373), .ZN(n12821) );
  NAND2_X1 U9738 ( .A1(n8657), .A2(n7386), .ZN(n7383) );
  NAND2_X1 U9739 ( .A1(n7392), .A2(n7391), .ZN(n13085) );
  NAND2_X1 U9740 ( .A1(n7392), .A2(n7389), .ZN(n7394) );
  NAND2_X1 U9741 ( .A1(n14340), .A2(n14339), .ZN(n7420) );
  INV_X1 U9742 ( .A(n7438), .ZN(n7439) );
  NAND2_X1 U9743 ( .A1(n14754), .A2(n14755), .ZN(n7452) );
  CLKBUF_X1 U9744 ( .A(n7452), .Z(n7446) );
  NOR2_X1 U9745 ( .A1(n14432), .A2(n7461), .ZN(n7460) );
  NAND2_X1 U9746 ( .A1(n14924), .A2(n7469), .ZN(n7466) );
  NAND2_X1 U9747 ( .A1(n14658), .A2(n9739), .ZN(n7474) );
  NAND2_X4 U9748 ( .A1(n9745), .A2(n14883), .ZN(n10483) );
  NAND2_X2 U9749 ( .A1(n9335), .A2(n9334), .ZN(n9745) );
  NAND2_X2 U9750 ( .A1(n10483), .A2(n8855), .ZN(n9370) );
  NAND2_X1 U9751 ( .A1(n13909), .A2(n8089), .ZN(n7487) );
  INV_X1 U9752 ( .A(n8089), .ZN(n7488) );
  NAND2_X1 U9753 ( .A1(n7824), .A2(n7504), .ZN(n11573) );
  NAND2_X1 U9754 ( .A1(n11082), .A2(n6773), .ZN(n7505) );
  NAND2_X1 U9755 ( .A1(n11082), .A2(n7800), .ZN(n11517) );
  NAND3_X1 U9756 ( .A1(n14780), .A2(n7507), .A3(n14668), .ZN(n14639) );
  NAND2_X1 U9757 ( .A1(n7508), .A2(n11341), .ZN(n11472) );
  NOR2_X2 U9758 ( .A1(n11916), .A2(n14275), .ZN(n11973) );
  NOR2_X2 U9759 ( .A1(n6693), .A2(n14851), .ZN(n12514) );
  NOR2_X2 U9760 ( .A1(n14956), .A2(n15164), .ZN(n7513) );
  AND2_X1 U9761 ( .A1(n6763), .A2(n7514), .ZN(n10737) );
  NAND2_X1 U9762 ( .A1(n10732), .A2(n10731), .ZN(n7514) );
  NAND3_X1 U9763 ( .A1(n7524), .A2(n6770), .A3(n7522), .ZN(n12411) );
  NAND2_X1 U9764 ( .A1(n12169), .A2(n7528), .ZN(n7522) );
  OR2_X2 U9765 ( .A1(n12169), .A2(n6710), .ZN(n7524) );
  NAND3_X1 U9766 ( .A1(n7524), .A2(n7526), .A3(n7522), .ZN(n12349) );
  NAND2_X1 U9767 ( .A1(n14094), .A2(n7538), .ZN(n7534) );
  NAND2_X1 U9768 ( .A1(n7534), .A2(n7535), .ZN(n14119) );
  NAND2_X1 U9769 ( .A1(n7542), .A2(n7543), .ZN(n12652) );
  NAND2_X1 U9770 ( .A1(n14188), .A2(n7544), .ZN(n7542) );
  NAND2_X1 U9771 ( .A1(n9320), .A2(n9318), .ZN(n9575) );
  INV_X1 U9772 ( .A(n7559), .ZN(n9701) );
  NAND2_X2 U9773 ( .A1(n7563), .A2(n13718), .ZN(n11052) );
  OAI21_X1 U9774 ( .B1(n13540), .B2(n13627), .A(n14032), .ZN(n7566) );
  NAND3_X1 U9775 ( .A1(n6677), .A2(n7720), .A3(n7568), .ZN(n8077) );
  INV_X1 U9776 ( .A(n7655), .ZN(n7568) );
  OAI21_X1 U9777 ( .B1(n11875), .B2(n7575), .A(n7573), .ZN(n12086) );
  OAI21_X1 U9778 ( .B1(n13519), .B2(n7585), .A(n7583), .ZN(n13545) );
  AND2_X1 U9779 ( .A1(n11425), .A2(n11417), .ZN(n7586) );
  NAND2_X1 U9780 ( .A1(n9320), .A2(n9319), .ZN(n7591) );
  NAND2_X1 U9781 ( .A1(n9408), .A2(n9407), .ZN(n11464) );
  OAI21_X1 U9782 ( .B1(n14217), .B2(n14337), .A(n7602), .ZN(n14223) );
  NAND2_X1 U9783 ( .A1(n14222), .A2(n14337), .ZN(n7602) );
  NAND2_X1 U9784 ( .A1(n15163), .A2(n7611), .ZN(n12313) );
  OAI211_X1 U9785 ( .C1(n9323), .C2(n7617), .A(n14872), .B(n7616), .ZN(n14881)
         );
  NAND2_X2 U9786 ( .A1(n13124), .A2(n6733), .ZN(n13110) );
  NAND2_X1 U9787 ( .A1(n8933), .A2(n7619), .ZN(n7618) );
  NAND2_X1 U9788 ( .A1(n12030), .A2(n7627), .ZN(n7625) );
  NAND2_X1 U9789 ( .A1(n8533), .A2(n8534), .ZN(n8446) );
  NAND2_X1 U9790 ( .A1(n9061), .A2(n7646), .ZN(n7645) );
  INV_X1 U9791 ( .A(n9059), .ZN(n7641) );
  NAND2_X1 U9792 ( .A1(n9059), .A2(n9060), .ZN(n7644) );
  AND3_X2 U9793 ( .A1(n7696), .A2(n7694), .A3(n7718), .ZN(n7652) );
  NOR2_X2 U9794 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n7654) );
  INV_X1 U9795 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n7653) );
  NAND3_X1 U9796 ( .A1(n9072), .A2(n9071), .A3(n7657), .ZN(n7656) );
  NAND2_X1 U9797 ( .A1(n7660), .A2(n7658), .ZN(n9090) );
  NAND2_X1 U9798 ( .A1(n7661), .A2(n7659), .ZN(n7658) );
  INV_X1 U9799 ( .A(n9083), .ZN(n7659) );
  INV_X1 U9800 ( .A(n9082), .ZN(n7661) );
  NAND2_X1 U9801 ( .A1(n9120), .A2(n7668), .ZN(n7666) );
  NAND2_X1 U9802 ( .A1(n7666), .A2(n7667), .ZN(n9127) );
  OAI21_X1 U9803 ( .B1(n9171), .B2(n9170), .A(n6784), .ZN(n7670) );
  INV_X1 U9804 ( .A(n9175), .ZN(n7671) );
  OR2_X1 U9805 ( .A1(n9332), .A2(n9424), .ZN(n9333) );
  NAND2_X1 U9806 ( .A1(n11664), .A2(n11663), .ZN(n11759) );
  OAI21_X1 U9807 ( .B1(n7762), .B2(n7763), .A(n7761), .ZN(n7770) );
  CLKBUF_X1 U9808 ( .A(n9745), .Z(n12662) );
  OR2_X1 U9809 ( .A1(n8811), .A2(n10444), .ZN(n8477) );
  NAND2_X4 U9810 ( .A1(n8465), .A2(n6884), .ZN(n8811) );
  INV_X1 U9811 ( .A(n14236), .ZN(n14239) );
  NAND2_X1 U9812 ( .A1(n9792), .A2(n9791), .ZN(n9795) );
  CLKBUF_X1 U9813 ( .A(n13519), .Z(n13522) );
  XNOR2_X1 U9814 ( .A(n8399), .B(n7313), .ZN(n13738) );
  CLKBUF_X1 U9815 ( .A(n12123), .Z(n11935) );
  NAND2_X2 U9816 ( .A1(n9866), .A2(n12748), .ZN(n12721) );
  NAND2_X1 U9817 ( .A1(n8929), .A2(n8928), .ZN(n15040) );
  XNOR2_X1 U9818 ( .A(n13109), .B(n13111), .ZN(n13312) );
  AND2_X1 U9819 ( .A1(n10565), .A2(n6676), .ZN(n15261) );
  NAND2_X1 U9820 ( .A1(n8931), .A2(n8930), .ZN(n8933) );
  NAND2_X1 U9821 ( .A1(n9793), .A2(n9870), .ZN(n9794) );
  OAI222_X1 U9822 ( .A1(n13440), .A2(n12668), .B1(P3_U3151), .B2(n12667), .C1(
        n12666), .C2(n12665), .ZN(P3_U3267) );
  INV_X1 U9823 ( .A(n8453), .ZN(n13437) );
  NAND2_X1 U9824 ( .A1(n9116), .A2(n9115), .ZN(n9120) );
  NAND2_X1 U9825 ( .A1(n9294), .A2(n9260), .ZN(n9261) );
  NAND4_X4 U9826 ( .A1(n8485), .A2(n8484), .A3(n8483), .A4(n8482), .ZN(n15698)
         );
  NAND4_X2 U9827 ( .A1(n8474), .A2(n8473), .A3(n8472), .A4(n8471), .ZN(n15682)
         );
  NAND2_X1 U9828 ( .A1(n7734), .A2(n14074), .ZN(n7777) );
  AND2_X1 U9829 ( .A1(n11385), .A2(n13916), .ZN(n13926) );
  INV_X1 U9830 ( .A(n14062), .ZN(n8423) );
  AND2_X2 U9831 ( .A1(n11384), .A2(n8419), .ZN(n15524) );
  OR2_X1 U9832 ( .A1(n11362), .A2(n9877), .ZN(n12797) );
  INV_X1 U9833 ( .A(n12797), .ZN(n9897) );
  OR2_X1 U9834 ( .A1(n15743), .A2(n15730), .ZN(n13424) );
  AND2_X1 U9835 ( .A1(n12504), .A2(n12502), .ZN(n7673) );
  AND2_X1 U9836 ( .A1(n12110), .A2(n12107), .ZN(n7674) );
  NAND2_X1 U9837 ( .A1(n13191), .A2(n13190), .ZN(n7675) );
  AND2_X1 U9838 ( .A1(n13453), .A2(n13452), .ZN(n7676) );
  NOR2_X1 U9839 ( .A1(n9496), .A2(n9481), .ZN(n7677) );
  AND2_X1 U9840 ( .A1(n7989), .A2(n10486), .ZN(n7678) );
  AND3_X1 U9841 ( .A1(n14025), .A2(n9049), .A3(n13725), .ZN(n7680) );
  AND2_X1 U9842 ( .A1(n13541), .A2(n13597), .ZN(n7681) );
  AND3_X1 U9843 ( .A1(n9318), .A2(n9758), .A3(n9764), .ZN(n7683) );
  AND2_X1 U9844 ( .A1(n12158), .A2(n12157), .ZN(n7684) );
  INV_X1 U9845 ( .A(n12137), .ZN(n8333) );
  AND2_X1 U9846 ( .A1(n11710), .A2(n11709), .ZN(n7685) );
  AND2_X2 U9847 ( .A1(n8385), .A2(n11043), .ZN(n15539) );
  INV_X1 U9848 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n8596) );
  INV_X1 U9849 ( .A(n15685), .ZN(n15703) );
  INV_X1 U9850 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n10222) );
  INV_X1 U9851 ( .A(n12934), .ZN(n13242) );
  NOR2_X1 U9852 ( .A1(n7712), .A2(n7711), .ZN(n7686) );
  INV_X1 U9853 ( .A(n8559), .ZN(n12820) );
  AND3_X1 U9854 ( .A1(n14468), .A2(n14467), .A3(n14466), .ZN(n7687) );
  INV_X1 U9855 ( .A(n15047), .ZN(n8656) );
  OR2_X1 U9856 ( .A1(n10390), .A2(n14750), .ZN(n7688) );
  NOR3_X1 U9857 ( .A1(n8411), .A2(n8352), .A3(n8410), .ZN(n7689) );
  NOR2_X1 U9858 ( .A1(n8938), .A2(n13259), .ZN(n7690) );
  NAND2_X1 U9859 ( .A1(n8845), .A2(n8844), .ZN(n13146) );
  INV_X1 U9860 ( .A(n13809), .ZN(n13804) );
  AND2_X1 U9861 ( .A1(n7821), .A2(n13663), .ZN(n7692) );
  OR2_X1 U9862 ( .A1(n9055), .A2(n9054), .ZN(n7693) );
  INV_X1 U9863 ( .A(n14277), .ZN(n14278) );
  OAI21_X1 U9864 ( .B1(n9141), .B2(n9140), .A(n9139), .ZN(n9138) );
  AOI21_X1 U9865 ( .B1(n9171), .B2(n9170), .A(n9168), .ZN(n9169) );
  INV_X1 U9866 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n7696) );
  INV_X1 U9867 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n9311) );
  INV_X1 U9868 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n7695) );
  OAI21_X1 U9869 ( .B1(n11313), .B2(n10912), .A(n10913), .ZN(n11301) );
  INV_X1 U9870 ( .A(n8871), .ZN(n8870) );
  INV_X1 U9871 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n8447) );
  INV_X1 U9872 ( .A(n12535), .ZN(n12536) );
  INV_X1 U9873 ( .A(n13127), .ZN(n9893) );
  INV_X1 U9874 ( .A(n9831), .ZN(n9826) );
  OR2_X1 U9875 ( .A1(n8958), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n10355) );
  INV_X1 U9876 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n12220) );
  INV_X1 U9877 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n8448) );
  INV_X1 U9878 ( .A(n13536), .ZN(n8388) );
  OR2_X1 U9879 ( .A1(n7777), .A2(n10712), .ZN(n7753) );
  OR3_X1 U9880 ( .A1(n14465), .A2(n14477), .A3(n14464), .ZN(n14466) );
  INV_X1 U9881 ( .A(n14402), .ZN(n14403) );
  INV_X1 U9882 ( .A(n9668), .ZN(n9303) );
  INV_X1 U9883 ( .A(n9619), .ZN(n9301) );
  INV_X1 U9884 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n9467) );
  OR2_X1 U9885 ( .A1(n9655), .A2(n14155), .ZN(n9668) );
  INV_X1 U9886 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n9315) );
  NOR2_X1 U9887 ( .A1(n9827), .A2(n9826), .ZN(n9828) );
  OR2_X1 U9888 ( .A1(n8885), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8902) );
  INV_X1 U9889 ( .A(n10355), .ZN(n13070) );
  AND2_X1 U9890 ( .A1(n12951), .A2(n13139), .ZN(n12960) );
  AND2_X1 U9891 ( .A1(n12990), .A2(n7356), .ZN(n9004) );
  OR2_X1 U9892 ( .A1(n8804), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8805) );
  NOR2_X1 U9893 ( .A1(P3_IR_REG_17__SCAN_IN), .A2(P3_IR_REG_15__SCAN_IN), .ZN(
        n8431) );
  AND2_X1 U9894 ( .A1(n8624), .A2(n8608), .ZN(n8609) );
  NAND2_X1 U9895 ( .A1(n10413), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n8538) );
  INV_X1 U9896 ( .A(n11276), .ZN(n11274) );
  NAND2_X1 U9897 ( .A1(n8056), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8105) );
  NAND2_X1 U9898 ( .A1(n13541), .A2(n8388), .ZN(n8389) );
  NAND2_X1 U9899 ( .A1(n8167), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n8192) );
  INV_X1 U9900 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n7703) );
  NAND2_X1 U9901 ( .A1(n9302), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n9643) );
  INV_X1 U9902 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n9428) );
  NAND2_X1 U9903 ( .A1(n14401), .A2(n14403), .ZN(n14404) );
  NAND2_X1 U9904 ( .A1(n9303), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n9670) );
  NAND2_X1 U9905 ( .A1(n9301), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n9631) );
  AND2_X1 U9906 ( .A1(n14812), .A2(n14174), .ZN(n9737) );
  NAND2_X1 U9907 ( .A1(n8240), .A2(n12290), .ZN(n8241) );
  NAND2_X1 U9908 ( .A1(n7869), .A2(SI_8_), .ZN(n7887) );
  NOR2_X1 U9909 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n9966), .ZN(n9914) );
  NOR2_X1 U9910 ( .A1(n9978), .A2(n9977), .ZN(n9922) );
  NAND2_X1 U9911 ( .A1(n8857), .A2(n12753), .ZN(n8871) );
  AND2_X1 U9912 ( .A1(n11993), .A2(n11992), .ZN(n13069) );
  INV_X1 U9913 ( .A(n15573), .ZN(n13015) );
  AND2_X1 U9914 ( .A1(n10920), .A2(n10918), .ZN(n10921) );
  INV_X1 U9915 ( .A(n13159), .ZN(n13195) );
  NAND2_X1 U9916 ( .A1(n13279), .A2(n12924), .ZN(n13265) );
  INV_X1 U9917 ( .A(n13425), .ZN(n11360) );
  OR2_X1 U9918 ( .A1(n13069), .A2(n13068), .ZN(n13368) );
  INV_X1 U9919 ( .A(n10362), .ZN(n13104) );
  INV_X1 U9920 ( .A(n15700), .ZN(n13276) );
  AND3_X1 U9921 ( .A1(n8431), .A2(n8430), .A3(n8697), .ZN(n8444) );
  AND2_X1 U9922 ( .A1(n8554), .A2(n8539), .ZN(n8552) );
  INV_X1 U9923 ( .A(n13510), .ZN(n11272) );
  INV_X1 U9924 ( .A(n8262), .ZN(n8264) );
  OR2_X1 U9925 ( .A1(n8192), .A2(n13572), .ZN(n8213) );
  INV_X1 U9926 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n11764) );
  XNOR2_X1 U9927 ( .A(n13473), .B(n13471), .ZN(n13590) );
  INV_X1 U9928 ( .A(n11424), .ZN(n11425) );
  INV_X1 U9929 ( .A(n13605), .ZN(n13621) );
  OR2_X1 U9930 ( .A1(n13750), .A2(n8338), .ZN(n8270) );
  INV_X1 U9931 ( .A(n8403), .ZN(n9220) );
  INV_X1 U9932 ( .A(n9272), .ZN(n11576) );
  NAND2_X1 U9933 ( .A1(n10865), .A2(n10864), .ZN(n10867) );
  OR2_X1 U9934 ( .A1(n10505), .A2(n11048), .ZN(n13615) );
  INV_X1 U9935 ( .A(n13906), .ZN(n13896) );
  INV_X1 U9936 ( .A(n8358), .ZN(n8355) );
  AND2_X1 U9937 ( .A1(n6763), .A2(n12646), .ZN(n10813) );
  NOR2_X1 U9938 ( .A1(n10819), .A2(n10818), .ZN(n11018) );
  OR2_X1 U9939 ( .A1(n14641), .A2(n9692), .ZN(n9688) );
  INV_X1 U9940 ( .A(n14717), .ZN(n15141) );
  INV_X1 U9941 ( .A(n11210), .ZN(n14422) );
  INV_X1 U9942 ( .A(n15334), .ZN(n15310) );
  OR2_X1 U9943 ( .A1(n10388), .A2(n14209), .ZN(n14928) );
  AND2_X1 U9944 ( .A1(n8071), .A2(n8049), .ZN(n8069) );
  AND2_X1 U9945 ( .A1(n7760), .A2(n7766), .ZN(n7761) );
  AND2_X1 U9946 ( .A1(n14555), .A2(n9942), .ZN(n9908) );
  INV_X1 U9947 ( .A(n9895), .ZN(n9896) );
  INV_X1 U9948 ( .A(n6852), .ZN(n10909) );
  INV_X1 U9949 ( .A(n11693), .ZN(n12990) );
  INV_X1 U9950 ( .A(n12726), .ZN(n13160) );
  INV_X1 U9951 ( .A(n15541), .ZN(n15628) );
  INV_X1 U9952 ( .A(n15675), .ZN(n15710) );
  INV_X1 U9953 ( .A(n13367), .ZN(n10382) );
  OR2_X1 U9954 ( .A1(n9017), .A2(n13425), .ZN(n9020) );
  INV_X1 U9955 ( .A(n13424), .ZN(n10379) );
  NAND2_X1 U9956 ( .A1(n11693), .A2(n11681), .ZN(n15730) );
  OR2_X1 U9957 ( .A1(n15680), .A2(n15734), .ZN(n15739) );
  AND2_X1 U9958 ( .A1(n11693), .A2(n15689), .ZN(n15734) );
  INV_X1 U9959 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n8568) );
  OR2_X1 U9960 ( .A1(n11055), .A2(n11123), .ZN(n11456) );
  AND2_X1 U9961 ( .A1(n8270), .A2(n8269), .ZN(n13536) );
  NOR2_X1 U9962 ( .A1(n11068), .A2(n11067), .ZN(n11232) );
  AND2_X1 U9963 ( .A1(n10523), .A2(n14081), .ZN(n15450) );
  AND2_X1 U9964 ( .A1(n15359), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15453) );
  INV_X1 U9965 ( .A(n9279), .ZN(n13874) );
  INV_X1 U9966 ( .A(n9275), .ZN(n11774) );
  AND2_X1 U9967 ( .A1(n13919), .A2(n11387), .ZN(n13924) );
  NOR2_X1 U9968 ( .A1(n8413), .A2(n15539), .ZN(n8414) );
  INV_X1 U9969 ( .A(n15465), .ZN(n11043) );
  INV_X1 U9970 ( .A(n15516), .ZN(n15508) );
  AND2_X1 U9971 ( .A1(n10406), .A2(n10500), .ZN(n11277) );
  NAND2_X1 U9972 ( .A1(n9537), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9551) );
  AND2_X1 U9973 ( .A1(n10741), .A2(n11095), .ZN(n14195) );
  OR2_X1 U9974 ( .A1(n10721), .A2(P1_U3086), .ZN(n14472) );
  AND2_X1 U9975 ( .A1(n9347), .A2(n9346), .ZN(n14666) );
  INV_X1 U9976 ( .A(n9657), .ZN(n9692) );
  AND2_X1 U9977 ( .A1(n10618), .A2(n10617), .ZN(n10889) );
  INV_X1 U9978 ( .A(n15266), .ZN(n15232) );
  INV_X1 U9979 ( .A(n15248), .ZN(n15258) );
  INV_X1 U9980 ( .A(n12509), .ZN(n14441) );
  INV_X1 U9981 ( .A(n14750), .ZN(n15126) );
  AND2_X1 U9982 ( .A1(n10394), .A2(n14619), .ZN(n15125) );
  AND2_X1 U9983 ( .A1(n11096), .A2(n11095), .ZN(n11098) );
  INV_X1 U9984 ( .A(n15160), .ZN(n15175) );
  INV_X1 U9985 ( .A(n15155), .ZN(n15337) );
  AND3_X1 U9986 ( .A1(n9785), .A2(n10720), .A3(n9784), .ZN(n11097) );
  NAND2_X1 U9987 ( .A1(n9766), .A2(n9767), .ZN(n10474) );
  AND2_X1 U9988 ( .A1(n10920), .A2(n10919), .ZN(n15623) );
  AOI21_X1 U9989 ( .B1(n10362), .B2(n9897), .A(n9896), .ZN(n9898) );
  INV_X1 U9990 ( .A(n12790), .ZN(n12440) );
  INV_X1 U9991 ( .A(n12372), .ZN(n15640) );
  INV_X1 U9992 ( .A(n15540), .ZN(n15626) );
  INV_X1 U9993 ( .A(n15032), .ZN(n15636) );
  AND2_X1 U9994 ( .A1(n13129), .A2(n13128), .ZN(n13319) );
  INV_X1 U9995 ( .A(n15693), .ZN(n13303) );
  NAND2_X1 U9996 ( .A1(n15751), .A2(n15070), .ZN(n13367) );
  AND3_X2 U9997 ( .A1(n11359), .A2(n9020), .A3(n9019), .ZN(n15751) );
  INV_X1 U9998 ( .A(n12812), .ZN(n13370) );
  INV_X2 U9999 ( .A(n15743), .ZN(n15741) );
  AND2_X1 U10000 ( .A1(n9008), .A2(n9007), .ZN(n15743) );
  INV_X1 U10001 ( .A(SI_17_), .ZN(n10834) );
  INV_X1 U10002 ( .A(SI_13_), .ZN(n10486) );
  INV_X1 U10003 ( .A(n10982), .ZN(n10937) );
  INV_X1 U10004 ( .A(n13624), .ZN(n13597) );
  NAND2_X1 U10005 ( .A1(n11280), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13607) );
  INV_X1 U10006 ( .A(n13486), .ZN(n13633) );
  INV_X1 U10007 ( .A(n13924), .ZN(n13902) );
  NAND2_X1 U10008 ( .A1(n13541), .A2(n14002), .ZN(n8386) );
  INV_X1 U10009 ( .A(n15539), .ZN(n15536) );
  INV_X1 U10010 ( .A(n15524), .ZN(n15523) );
  OR2_X1 U10011 ( .A1(n15467), .A2(n15463), .ZN(n15464) );
  INV_X1 U10012 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n11689) );
  NAND2_X1 U10013 ( .A1(n11200), .A2(P1_STATE_REG_SCAN_IN), .ZN(n15119) );
  INV_X1 U10014 ( .A(n14368), .ZN(n14480) );
  INV_X1 U10015 ( .A(n14324), .ZN(n14761) );
  INV_X1 U10016 ( .A(n15087), .ZN(n14491) );
  OR2_X1 U10017 ( .A1(n10407), .A2(n10734), .ZN(n14501) );
  OR2_X1 U10018 ( .A1(n10698), .A2(n14520), .ZN(n15266) );
  INV_X1 U10019 ( .A(n15125), .ZN(n14958) );
  OR2_X1 U10020 ( .A1(n10720), .A2(n10738), .ZN(n15136) );
  INV_X1 U10021 ( .A(n15143), .ZN(n14765) );
  INV_X1 U10022 ( .A(n15358), .ZN(n15355) );
  NAND2_X1 U10023 ( .A1(n15339), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n9787) );
  INV_X1 U10024 ( .A(n15341), .ZN(n15339) );
  AND2_X2 U10025 ( .A1(n9786), .A2(n11097), .ZN(n15341) );
  AND2_X1 U10026 ( .A1(n10482), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10478) );
  INV_X1 U10027 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n11733) );
  INV_X1 U10028 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10838) );
  NAND2_X1 U10029 ( .A1(n15753), .A2(n15754), .ZN(n15752) );
  XNOR2_X1 U10030 ( .A(n10339), .B(n10338), .ZN(n10340) );
  AND2_X1 U10031 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10503), .ZN(P2_U3947) );
  INV_X1 U10032 ( .A(n14501), .ZN(P1_U4016) );
  NAND2_X1 U10033 ( .A1(n7688), .A2(n10404), .ZN(P1_U3356) );
  NAND2_X1 U10034 ( .A1(n9788), .A2(n9787), .ZN(P1_U3525) );
  NOR2_X4 U10035 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n7718) );
  NOR2_X1 U10036 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), 
        .ZN(n8076) );
  NOR2_X1 U10037 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), 
        .ZN(n7698) );
  NOR2_X1 U10038 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), 
        .ZN(n7697) );
  NAND4_X1 U10039 ( .A1(n8076), .A2(n7698), .A3(n7697), .A4(n8074), .ZN(n7704)
         );
  INV_X1 U10040 ( .A(n7704), .ZN(n7699) );
  NAND2_X2 U10041 ( .A1(n7700), .A2(n7703), .ZN(n8282) );
  AND2_X1 U10042 ( .A1(P2_IR_REG_28__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), 
        .ZN(n7707) );
  NOR2_X1 U10043 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), 
        .ZN(n7702) );
  NOR2_X1 U10044 ( .A1(P2_IR_REG_26__SCAN_IN), .A2(P2_IR_REG_25__SCAN_IN), 
        .ZN(n7701) );
  AND2_X1 U10045 ( .A1(n7702), .A2(n7701), .ZN(n7709) );
  NOR2_X1 U10046 ( .A1(P2_IR_REG_28__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), 
        .ZN(n7708) );
  NAND4_X1 U10047 ( .A1(n7709), .A2(n7708), .A3(n7703), .A4(n8283), .ZN(n7705)
         );
  NOR2_X1 U10048 ( .A1(n7705), .A2(n7704), .ZN(n7706) );
  NAND2_X1 U10049 ( .A1(n7974), .A2(n7706), .ZN(n7726) );
  INV_X1 U10050 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n14065) );
  INV_X1 U10051 ( .A(n7709), .ZN(n8344) );
  NOR2_X1 U10052 ( .A1(n8344), .A2(n7710), .ZN(n7711) );
  INV_X1 U10053 ( .A(n10433), .ZN(n8855) );
  NOR2_X1 U10054 ( .A1(n7718), .A2(n14065), .ZN(n7719) );
  MUX2_X1 U10055 ( .A(n14065), .B(n7719), .S(P2_IR_REG_2__SCAN_IN), .Z(n7721)
         );
  NOR2_X1 U10056 ( .A1(n7721), .A2(n7720), .ZN(n10524) );
  AOI22_X1 U10057 ( .A1(n6717), .A2(P1_DATAO_REG_2__SCAN_IN), .B1(n10524), 
        .B2(n7821), .ZN(n7724) );
  INV_X1 U10058 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n9376) );
  INV_X1 U10059 ( .A(SI_0_), .ZN(n10454) );
  NAND2_X1 U10060 ( .A1(n7743), .A2(n7722), .ZN(n7769) );
  NAND2_X1 U10061 ( .A1(n7769), .A2(SI_2_), .ZN(n7760) );
  OAI21_X1 U10062 ( .B1(n7769), .B2(SI_2_), .A(n7760), .ZN(n7762) );
  MUX2_X1 U10063 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(P1_DATAO_REG_2__SCAN_IN), 
        .S(n10433), .Z(n7764) );
  XNOR2_X1 U10064 ( .A(n7762), .B(n7764), .ZN(n10411) );
  NAND2_X1 U10065 ( .A1(n10411), .A2(n7818), .ZN(n7723) );
  INV_X1 U10066 ( .A(n7726), .ZN(n7728) );
  NAND2_X1 U10067 ( .A1(n7728), .A2(n7727), .ZN(n7730) );
  INV_X1 U10068 ( .A(n7734), .ZN(n14069) );
  NAND2_X1 U10069 ( .A1(n7774), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n7738) );
  INV_X1 U10070 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n7732) );
  NAND2_X1 U10071 ( .A1(n8253), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n7736) );
  INV_X1 U10072 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n10525) );
  OR2_X1 U10073 ( .A1(n7777), .A2(n10525), .ZN(n7735) );
  NAND2_X1 U10074 ( .A1(n6717), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n7746) );
  INV_X1 U10075 ( .A(n7739), .ZN(n7740) );
  NAND2_X1 U10076 ( .A1(n7741), .A2(n7740), .ZN(n7742) );
  NAND2_X1 U10077 ( .A1(n7743), .A2(n7742), .ZN(n10466) );
  XNOR2_X1 U10078 ( .A(n7744), .B(P2_IR_REG_1__SCAN_IN), .ZN(n13663) );
  NAND2_X1 U10079 ( .A1(n8253), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n7751) );
  INV_X1 U10080 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n7747) );
  INV_X1 U10081 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n13935) );
  OR2_X1 U10082 ( .A1(n7777), .A2(n13935), .ZN(n7748) );
  XNOR2_X1 U10083 ( .A(n11459), .B(n13658), .ZN(n8289) );
  NAND2_X1 U10084 ( .A1(n8253), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n7756) );
  NAND2_X1 U10085 ( .A1(n7774), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n7755) );
  INV_X1 U10086 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n7752) );
  INV_X1 U10087 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n10712) );
  NAND2_X1 U10088 ( .A1(n10433), .A2(SI_0_), .ZN(n7757) );
  XNOR2_X1 U10089 ( .A(n7757), .B(n8464), .ZN(n14084) );
  INV_X1 U10090 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n13665) );
  MUX2_X1 U10091 ( .A(n14084), .B(n13665), .S(n7821), .Z(n11491) );
  INV_X1 U10092 ( .A(n11491), .ZN(n11053) );
  NAND2_X1 U10093 ( .A1(n9025), .A2(n11053), .ZN(n10824) );
  NAND2_X1 U10094 ( .A1(n8289), .A2(n10824), .ZN(n10823) );
  INV_X1 U10095 ( .A(n13658), .ZN(n11122) );
  NAND2_X1 U10096 ( .A1(n11122), .A2(n11459), .ZN(n7758) );
  NAND2_X1 U10097 ( .A1(n10823), .A2(n7758), .ZN(n10852) );
  OR2_X1 U10098 ( .A1(n11129), .A2(n13656), .ZN(n7759) );
  INV_X1 U10099 ( .A(SI_2_), .ZN(n10424) );
  NOR2_X1 U10100 ( .A1(n7763), .A2(n10424), .ZN(n7768) );
  NOR2_X1 U10101 ( .A1(n7764), .A2(SI_2_), .ZN(n7765) );
  NOR2_X1 U10102 ( .A1(n7766), .A2(n7765), .ZN(n7767) );
  OR2_X1 U10103 ( .A1(n10440), .A2(n7913), .ZN(n7773) );
  OR2_X1 U10104 ( .A1(n7720), .A2(n14065), .ZN(n7771) );
  XNOR2_X1 U10105 ( .A(n7771), .B(P2_IR_REG_3__SCAN_IN), .ZN(n10526) );
  AOI22_X1 U10106 ( .A1(n6717), .A2(P1_DATAO_REG_3__SCAN_IN), .B1(n10526), 
        .B2(n7821), .ZN(n7772) );
  NAND2_X1 U10107 ( .A1(n9219), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n7781) );
  OR2_X1 U10108 ( .A1(n8338), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n7780) );
  INV_X1 U10109 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n7776) );
  OR2_X1 U10110 ( .A1(n8403), .A2(n7776), .ZN(n7779) );
  INV_X1 U10111 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n11396) );
  OR2_X1 U10112 ( .A1(n9223), .A2(n11396), .ZN(n7778) );
  INV_X1 U10113 ( .A(n13655), .ZN(n11090) );
  XNOR2_X1 U10114 ( .A(n13515), .B(n11090), .ZN(n10864) );
  OR2_X1 U10115 ( .A1(n13515), .A2(n13655), .ZN(n7782) );
  NAND2_X1 U10116 ( .A1(n10867), .A2(n7782), .ZN(n11084) );
  MUX2_X1 U10117 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(P1_DATAO_REG_4__SCAN_IN), 
        .S(n10433), .Z(n7785) );
  NAND2_X1 U10118 ( .A1(n7785), .A2(SI_4_), .ZN(n7811) );
  NAND2_X1 U10119 ( .A1(n7786), .A2(n7787), .ZN(n7790) );
  INV_X1 U10120 ( .A(n7787), .ZN(n7788) );
  NAND2_X1 U10121 ( .A1(n7790), .A2(n7812), .ZN(n10435) );
  OR2_X1 U10122 ( .A1(n10435), .A2(n7913), .ZN(n7794) );
  NAND2_X1 U10123 ( .A1(n7720), .A2(n7791), .ZN(n7819) );
  XNOR2_X1 U10124 ( .A(n7792), .B(P2_IR_REG_4__SCAN_IN), .ZN(n10527) );
  AOI22_X1 U10125 ( .A1(n6717), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n10527), 
        .B2(n7821), .ZN(n7793) );
  NAND2_X1 U10126 ( .A1(n9219), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n7799) );
  NAND2_X1 U10127 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n7803) );
  OAI21_X1 U10128 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(P2_REG3_REG_3__SCAN_IN), 
        .A(n7803), .ZN(n11402) );
  OR2_X1 U10129 ( .A1(n8338), .A2(n11402), .ZN(n7798) );
  INV_X1 U10130 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n7795) );
  OR2_X1 U10131 ( .A1(n8403), .A2(n7795), .ZN(n7797) );
  INV_X1 U10132 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n11407) );
  OR2_X1 U10133 ( .A1(n9223), .A2(n11407), .ZN(n7796) );
  NAND4_X1 U10134 ( .A1(n7799), .A2(n7798), .A3(n7797), .A4(n7796), .ZN(n13654) );
  INV_X1 U10135 ( .A(n11087), .ZN(n11083) );
  NAND2_X1 U10136 ( .A1(n11084), .A2(n11083), .ZN(n11082) );
  OR2_X1 U10137 ( .A1(n11400), .A2(n13654), .ZN(n7800) );
  NAND2_X1 U10138 ( .A1(n9219), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n7810) );
  INV_X1 U10139 ( .A(n7803), .ZN(n7801) );
  NAND2_X1 U10140 ( .A1(n7801), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7839) );
  INV_X1 U10141 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n7802) );
  NAND2_X1 U10142 ( .A1(n7803), .A2(n7802), .ZN(n7804) );
  NAND2_X1 U10143 ( .A1(n7839), .A2(n7804), .ZN(n11521) );
  OR2_X1 U10144 ( .A1(n8338), .A2(n11521), .ZN(n7809) );
  INV_X1 U10145 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n7805) );
  OR2_X1 U10146 ( .A1(n8403), .A2(n7805), .ZN(n7808) );
  INV_X1 U10147 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n7806) );
  OR2_X1 U10148 ( .A1(n9223), .A2(n7806), .ZN(n7807) );
  NAND4_X1 U10149 ( .A1(n7810), .A2(n7809), .A3(n7808), .A4(n7807), .ZN(n13653) );
  INV_X1 U10150 ( .A(n13653), .ZN(n11089) );
  MUX2_X1 U10151 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n10433), .Z(n7813) );
  NAND2_X1 U10152 ( .A1(n7813), .A2(SI_5_), .ZN(n7825) );
  OAI21_X1 U10153 ( .B1(n7813), .B2(SI_5_), .A(n7825), .ZN(n7814) );
  INV_X1 U10154 ( .A(n7814), .ZN(n7815) );
  NAND2_X1 U10155 ( .A1(n7816), .A2(n7815), .ZN(n7826) );
  OR2_X1 U10156 ( .A1(n7816), .A2(n7815), .ZN(n7817) );
  AND2_X1 U10157 ( .A1(n7826), .A2(n7817), .ZN(n10442) );
  NAND2_X1 U10158 ( .A1(n10442), .A2(n9234), .ZN(n7823) );
  NAND2_X1 U10159 ( .A1(n7832), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7820) );
  XNOR2_X1 U10160 ( .A(n7820), .B(P2_IR_REG_5__SCAN_IN), .ZN(n10766) );
  AOI22_X1 U10161 ( .A1(n6717), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n10766), 
        .B2(n7821), .ZN(n7822) );
  NAND2_X1 U10162 ( .A1(n7823), .A2(n7822), .ZN(n11523) );
  INV_X1 U10163 ( .A(n11523), .ZN(n15476) );
  NAND2_X1 U10164 ( .A1(n11517), .A2(n11089), .ZN(n7824) );
  NAND2_X1 U10165 ( .A1(n7826), .A2(n7825), .ZN(n7830) );
  MUX2_X1 U10166 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n10432), .Z(n7827) );
  OAI21_X1 U10167 ( .B1(SI_6_), .B2(n7827), .A(n7847), .ZN(n7828) );
  INV_X1 U10168 ( .A(n7828), .ZN(n7829) );
  OR2_X1 U10169 ( .A1(n7830), .A2(n7829), .ZN(n7831) );
  NAND2_X1 U10170 ( .A1(n7848), .A2(n7831), .ZN(n10437) );
  OR2_X1 U10171 ( .A1(n10437), .A2(n7913), .ZN(n7836) );
  INV_X1 U10172 ( .A(n7832), .ZN(n7833) );
  NAND2_X1 U10173 ( .A1(n7833), .A2(n7653), .ZN(n7853) );
  NAND2_X1 U10174 ( .A1(n7853), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7834) );
  XNOR2_X1 U10175 ( .A(n7834), .B(P2_IR_REG_6__SCAN_IN), .ZN(n10542) );
  AOI22_X1 U10176 ( .A1(n6717), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n10542), 
        .B2(n7821), .ZN(n7835) );
  NAND2_X1 U10177 ( .A1(n9219), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n7845) );
  INV_X1 U10178 ( .A(n7839), .ZN(n7837) );
  NAND2_X1 U10179 ( .A1(n7837), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n7860) );
  INV_X1 U10180 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n7838) );
  NAND2_X1 U10181 ( .A1(n7839), .A2(n7838), .ZN(n7840) );
  NAND2_X1 U10182 ( .A1(n7860), .A2(n7840), .ZN(n11585) );
  OR2_X1 U10183 ( .A1(n8338), .A2(n11585), .ZN(n7844) );
  INV_X1 U10184 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n7841) );
  OR2_X1 U10185 ( .A1(n8403), .A2(n7841), .ZN(n7843) );
  INV_X1 U10186 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n11582) );
  OR2_X1 U10187 ( .A1(n9223), .A2(n11582), .ZN(n7842) );
  NAND4_X1 U10188 ( .A1(n7845), .A2(n7844), .A3(n7843), .A4(n7842), .ZN(n13652) );
  INV_X1 U10189 ( .A(n13652), .ZN(n9075) );
  XNOR2_X1 U10190 ( .A(n11429), .B(n9075), .ZN(n9272) );
  NAND2_X1 U10191 ( .A1(n11429), .A2(n13652), .ZN(n7846) );
  MUX2_X1 U10192 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n6671), .Z(n7849) );
  NAND2_X1 U10193 ( .A1(n7849), .A2(SI_7_), .ZN(n7867) );
  OAI21_X1 U10194 ( .B1(n7849), .B2(SI_7_), .A(n7867), .ZN(n7850) );
  INV_X1 U10195 ( .A(n7850), .ZN(n7851) );
  INV_X1 U10196 ( .A(n7853), .ZN(n7855) );
  NAND2_X1 U10197 ( .A1(n7855), .A2(n7854), .ZN(n7874) );
  NAND2_X1 U10198 ( .A1(n7874), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7856) );
  XNOR2_X1 U10199 ( .A(n7856), .B(P2_IR_REG_7__SCAN_IN), .ZN(n10749) );
  AOI22_X1 U10200 ( .A1(n6717), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n10749), 
        .B2(n7821), .ZN(n7857) );
  NAND2_X1 U10201 ( .A1(n7858), .A2(n7857), .ZN(n11594) );
  NAND2_X1 U10202 ( .A1(n9219), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7866) );
  INV_X1 U10203 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n7859) );
  NAND2_X1 U10204 ( .A1(n7860), .A2(n7859), .ZN(n7861) );
  NAND2_X1 U10205 ( .A1(n7879), .A2(n7861), .ZN(n11595) );
  OR2_X1 U10206 ( .A1(n8338), .A2(n11595), .ZN(n7865) );
  INV_X1 U10207 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n7862) );
  OR2_X1 U10208 ( .A1(n8403), .A2(n7862), .ZN(n7864) );
  OR2_X1 U10209 ( .A1(n9223), .A2(n10755), .ZN(n7863) );
  NAND4_X1 U10210 ( .A1(n7866), .A2(n7865), .A3(n7864), .A4(n7863), .ZN(n13651) );
  INV_X1 U10211 ( .A(n13651), .ZN(n8299) );
  XNOR2_X1 U10212 ( .A(n11594), .B(n8299), .ZN(n11599) );
  MUX2_X1 U10213 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n6671), .Z(n7869) );
  OAI21_X1 U10214 ( .B1(SI_8_), .B2(n7869), .A(n7887), .ZN(n7870) );
  INV_X1 U10215 ( .A(n7870), .ZN(n7871) );
  OR2_X1 U10216 ( .A1(n7872), .A2(n7871), .ZN(n7873) );
  NAND2_X1 U10217 ( .A1(n7888), .A2(n7873), .ZN(n10471) );
  OR2_X1 U10218 ( .A1(n10471), .A2(n7913), .ZN(n7877) );
  NAND2_X1 U10219 ( .A1(n7890), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7875) );
  XNOR2_X1 U10220 ( .A(n7875), .B(P2_IR_REG_8__SCAN_IN), .ZN(n10784) );
  AOI22_X1 U10221 ( .A1(n6717), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n10784), 
        .B2(n7821), .ZN(n7876) );
  NAND2_X1 U10222 ( .A1(n7877), .A2(n7876), .ZN(n11662) );
  NAND2_X1 U10223 ( .A1(n9219), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n7885) );
  INV_X1 U10224 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n7878) );
  NAND2_X1 U10225 ( .A1(n7879), .A2(n7878), .ZN(n7880) );
  NAND2_X1 U10226 ( .A1(n7896), .A2(n7880), .ZN(n11642) );
  OR2_X1 U10227 ( .A1(n8338), .A2(n11642), .ZN(n7884) );
  INV_X1 U10228 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n7881) );
  OR2_X1 U10229 ( .A1(n8403), .A2(n7881), .ZN(n7883) );
  INV_X1 U10230 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n10757) );
  OR2_X1 U10231 ( .A1(n9223), .A2(n10757), .ZN(n7882) );
  NAND4_X1 U10232 ( .A1(n7885), .A2(n7884), .A3(n7883), .A4(n7882), .ZN(n13650) );
  INV_X1 U10233 ( .A(n13650), .ZN(n8302) );
  XNOR2_X1 U10234 ( .A(n11662), .B(n8302), .ZN(n11638) );
  NAND2_X1 U10235 ( .A1(n11639), .A2(n11638), .ZN(n11641) );
  NAND2_X1 U10236 ( .A1(n11662), .A2(n13650), .ZN(n7886) );
  MUX2_X1 U10237 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n6671), .Z(n7889) );
  NAND2_X1 U10238 ( .A1(n7889), .A2(SI_9_), .ZN(n7907) );
  NAND2_X1 U10239 ( .A1(n10487), .A2(n9234), .ZN(n7895) );
  INV_X1 U10240 ( .A(n7890), .ZN(n7892) );
  INV_X1 U10241 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n7891) );
  NAND2_X1 U10242 ( .A1(n7892), .A2(n7891), .ZN(n7914) );
  NAND2_X1 U10243 ( .A1(n7914), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7893) );
  XNOR2_X1 U10244 ( .A(n7893), .B(P2_IR_REG_9__SCAN_IN), .ZN(n10794) );
  AOI22_X1 U10245 ( .A1(n8396), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n10794), 
        .B2(n7821), .ZN(n7894) );
  NAND2_X1 U10246 ( .A1(n7895), .A2(n7894), .ZN(n11755) );
  NAND2_X1 U10247 ( .A1(n9219), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n7902) );
  NAND2_X1 U10248 ( .A1(n7896), .A2(n11764), .ZN(n7897) );
  NAND2_X1 U10249 ( .A1(n7921), .A2(n7897), .ZN(n11610) );
  OR2_X1 U10250 ( .A1(n8338), .A2(n11610), .ZN(n7901) );
  INV_X1 U10251 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n7898) );
  OR2_X1 U10252 ( .A1(n8403), .A2(n7898), .ZN(n7900) );
  INV_X1 U10253 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n10788) );
  OR2_X1 U10254 ( .A1(n9223), .A2(n10788), .ZN(n7899) );
  NAND4_X1 U10255 ( .A1(n7902), .A2(n7901), .A3(n7900), .A4(n7899), .ZN(n13649) );
  XNOR2_X1 U10256 ( .A(n11755), .B(n13649), .ZN(n9273) );
  INV_X1 U10257 ( .A(n9273), .ZN(n11613) );
  NAND2_X1 U10258 ( .A1(n11607), .A2(n11613), .ZN(n11606) );
  NAND2_X1 U10259 ( .A1(n11755), .A2(n13649), .ZN(n7903) );
  NAND2_X1 U10260 ( .A1(n11606), .A2(n7903), .ZN(n11771) );
  INV_X1 U10261 ( .A(n7904), .ZN(n7905) );
  MUX2_X1 U10262 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n6671), .Z(n7908) );
  OAI21_X1 U10263 ( .B1(SI_10_), .B2(n7908), .A(n7930), .ZN(n7909) );
  INV_X1 U10264 ( .A(n7909), .ZN(n7910) );
  OR2_X1 U10265 ( .A1(n7911), .A2(n7910), .ZN(n7912) );
  NAND2_X1 U10266 ( .A1(n7931), .A2(n7912), .ZN(n10492) );
  OR2_X1 U10267 ( .A1(n10492), .A2(n7913), .ZN(n7919) );
  INV_X1 U10268 ( .A(n7914), .ZN(n7916) );
  NAND2_X1 U10269 ( .A1(n7916), .A2(n7915), .ZN(n7932) );
  XNOR2_X1 U10270 ( .A(n7917), .B(P2_IR_REG_10__SCAN_IN), .ZN(n11072) );
  AOI22_X1 U10271 ( .A1(n11072), .A2(n7821), .B1(n6717), .B2(
        P1_DATAO_REG_10__SCAN_IN), .ZN(n7918) );
  NAND2_X1 U10272 ( .A1(n9219), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n7927) );
  INV_X1 U10273 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n11884) );
  NAND2_X1 U10274 ( .A1(n7921), .A2(n11884), .ZN(n7922) );
  NAND2_X1 U10275 ( .A1(n7937), .A2(n7922), .ZN(n11780) );
  OR2_X1 U10276 ( .A1(n8338), .A2(n11780), .ZN(n7926) );
  INV_X1 U10277 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n7923) );
  OR2_X1 U10278 ( .A1(n8403), .A2(n7923), .ZN(n7925) );
  INV_X1 U10279 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n11065) );
  OR2_X1 U10280 ( .A1(n9223), .A2(n11065), .ZN(n7924) );
  NAND4_X1 U10281 ( .A1(n7927), .A2(n7926), .A3(n7925), .A4(n7924), .ZN(n13648) );
  INV_X1 U10282 ( .A(n13648), .ZN(n9094) );
  NAND2_X1 U10283 ( .A1(n15507), .A2(n9094), .ZN(n11893) );
  OR2_X1 U10284 ( .A1(n15507), .A2(n9094), .ZN(n7928) );
  NAND2_X1 U10285 ( .A1(n11771), .A2(n11774), .ZN(n11770) );
  NAND2_X1 U10286 ( .A1(n15507), .A2(n13648), .ZN(n7929) );
  MUX2_X1 U10287 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(P1_DATAO_REG_11__SCAN_IN), 
        .S(n6671), .Z(n7946) );
  XNOR2_X1 U10288 ( .A(n7950), .B(n7949), .ZN(n10496) );
  NAND2_X1 U10289 ( .A1(n10496), .A2(n9234), .ZN(n7935) );
  XNOR2_X1 U10290 ( .A(n7933), .B(P2_IR_REG_11__SCAN_IN), .ZN(n11229) );
  AOI22_X1 U10291 ( .A1(n11229), .A2(n7821), .B1(P1_DATAO_REG_11__SCAN_IN), 
        .B2(n8396), .ZN(n7934) );
  NAND2_X1 U10292 ( .A1(n9219), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n7943) );
  INV_X1 U10293 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n7936) );
  NAND2_X1 U10294 ( .A1(n7937), .A2(n7936), .ZN(n7938) );
  NAND2_X1 U10295 ( .A1(n7956), .A2(n7938), .ZN(n11903) );
  OR2_X1 U10296 ( .A1(n8338), .A2(n11903), .ZN(n7942) );
  INV_X1 U10297 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n7939) );
  OR2_X1 U10298 ( .A1(n8403), .A2(n7939), .ZN(n7941) );
  INV_X1 U10299 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n11066) );
  OR2_X1 U10300 ( .A1(n9223), .A2(n11066), .ZN(n7940) );
  NAND4_X1 U10301 ( .A1(n7943), .A2(n7942), .A3(n7941), .A4(n7940), .ZN(n13647) );
  OR2_X1 U10302 ( .A1(n12068), .A2(n13647), .ZN(n7944) );
  NAND2_X1 U10303 ( .A1(n12068), .A2(n13647), .ZN(n7945) );
  INV_X1 U10304 ( .A(n7946), .ZN(n7947) );
  NAND2_X1 U10305 ( .A1(n7947), .A2(n10450), .ZN(n7948) );
  MUX2_X1 U10306 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(P1_DATAO_REG_12__SCAN_IN), 
        .S(n6671), .Z(n7967) );
  XNOR2_X1 U10307 ( .A(n7966), .B(n7965), .ZN(n10745) );
  NAND2_X1 U10308 ( .A1(n10745), .A2(n9234), .ZN(n7953) );
  XNOR2_X1 U10309 ( .A(n7951), .B(P2_IR_REG_12__SCAN_IN), .ZN(n13674) );
  AOI22_X1 U10310 ( .A1(n8396), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n13674), 
        .B2(n7821), .ZN(n7952) );
  INV_X1 U10311 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7955) );
  NAND2_X1 U10312 ( .A1(n7956), .A2(n7955), .ZN(n7957) );
  NAND2_X1 U10313 ( .A1(n7979), .A2(n7957), .ZN(n12113) );
  OR2_X1 U10314 ( .A1(n8338), .A2(n12113), .ZN(n7962) );
  INV_X1 U10315 ( .A(n9219), .ZN(n8402) );
  INV_X1 U10316 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n13687) );
  OR2_X1 U10317 ( .A1(n8402), .A2(n13687), .ZN(n7961) );
  INV_X1 U10318 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n7958) );
  OR2_X1 U10319 ( .A1(n8403), .A2(n7958), .ZN(n7960) );
  INV_X1 U10320 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n11960) );
  OR2_X1 U10321 ( .A1(n9223), .A2(n11960), .ZN(n7959) );
  NAND4_X1 U10322 ( .A1(n7962), .A2(n7961), .A3(n7960), .A4(n7959), .ZN(n13646) );
  AND2_X1 U10323 ( .A1(n14019), .A2(n13646), .ZN(n7963) );
  OR2_X1 U10324 ( .A1(n14019), .A2(n13646), .ZN(n7964) );
  INV_X1 U10325 ( .A(n7967), .ZN(n7968) );
  NAND2_X1 U10326 ( .A1(n7968), .A2(n10457), .ZN(n7969) );
  MUX2_X1 U10327 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(P1_DATAO_REG_13__SCAN_IN), 
        .S(n6671), .Z(n7990) );
  XNOR2_X1 U10328 ( .A(n7990), .B(n10486), .ZN(n7971) );
  XNOR2_X1 U10329 ( .A(n7992), .B(n7971), .ZN(n10836) );
  NAND2_X1 U10330 ( .A1(n10836), .A2(n9234), .ZN(n7977) );
  MUX2_X1 U10331 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7973), .S(
        P2_IR_REG_13__SCAN_IN), .Z(n7975) );
  INV_X1 U10332 ( .A(n7974), .ZN(n7995) );
  AND2_X1 U10333 ( .A1(n7975), .A2(n7995), .ZN(n13689) );
  AOI22_X1 U10334 ( .A1(n8396), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n13689), 
        .B2(n7821), .ZN(n7976) );
  INV_X1 U10335 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n7978) );
  NAND2_X1 U10336 ( .A1(n7979), .A2(n7978), .ZN(n7980) );
  AND2_X1 U10337 ( .A1(n7999), .A2(n7980), .ZN(n12089) );
  NAND2_X1 U10338 ( .A1(n8253), .A2(n12089), .ZN(n7985) );
  INV_X1 U10339 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n13690) );
  OR2_X1 U10340 ( .A1(n8402), .A2(n13690), .ZN(n7984) );
  INV_X1 U10341 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n7981) );
  OR2_X1 U10342 ( .A1(n8403), .A2(n7981), .ZN(n7983) );
  INV_X1 U10343 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n13675) );
  OR2_X1 U10344 ( .A1(n9223), .A2(n13675), .ZN(n7982) );
  NAND4_X1 U10345 ( .A1(n7985), .A2(n7984), .A3(n7983), .A4(n7982), .ZN(n13645) );
  NAND2_X1 U10346 ( .A1(n7986), .A2(n13645), .ZN(n7988) );
  NAND2_X1 U10347 ( .A1(n7988), .A2(n7987), .ZN(n12210) );
  INV_X1 U10348 ( .A(n7990), .ZN(n7989) );
  NAND2_X1 U10349 ( .A1(n7990), .A2(SI_13_), .ZN(n7991) );
  MUX2_X1 U10350 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(P1_DATAO_REG_14__SCAN_IN), 
        .S(n6671), .Z(n8009) );
  XNOR2_X1 U10351 ( .A(n8010), .B(n8009), .ZN(n11350) );
  NAND2_X1 U10352 ( .A1(n11350), .A2(n9234), .ZN(n7998) );
  XNOR2_X1 U10353 ( .A(n7996), .B(P2_IR_REG_14__SCAN_IN), .ZN(n15417) );
  AOI22_X1 U10354 ( .A1(n8396), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n15417), 
        .B2(n7821), .ZN(n7997) );
  INV_X1 U10355 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n12251) );
  NAND2_X1 U10356 ( .A1(n7999), .A2(n12251), .ZN(n8000) );
  NAND2_X1 U10357 ( .A1(n8020), .A2(n8000), .ZN(n12250) );
  INV_X1 U10358 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n8001) );
  OR2_X1 U10359 ( .A1(n8403), .A2(n8001), .ZN(n8003) );
  INV_X1 U10360 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n13692) );
  OR2_X1 U10361 ( .A1(n8402), .A2(n13692), .ZN(n8002) );
  AND2_X1 U10362 ( .A1(n8003), .A2(n8002), .ZN(n8005) );
  INV_X1 U10363 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n12206) );
  OR2_X1 U10364 ( .A1(n9223), .A2(n12206), .ZN(n8004) );
  OAI211_X1 U10365 ( .C1(n12250), .C2(n8338), .A(n8005), .B(n8004), .ZN(n13644) );
  XNOR2_X1 U10366 ( .A(n12277), .B(n13644), .ZN(n12209) );
  INV_X1 U10367 ( .A(n12209), .ZN(n8006) );
  NAND2_X1 U10368 ( .A1(n12277), .A2(n13644), .ZN(n8007) );
  MUX2_X1 U10369 ( .A(n11547), .B(n11549), .S(n6671), .Z(n8011) );
  NAND2_X1 U10370 ( .A1(n8011), .A2(n10594), .ZN(n8025) );
  INV_X1 U10371 ( .A(n8011), .ZN(n8012) );
  NAND2_X1 U10372 ( .A1(n8012), .A2(SI_15_), .ZN(n8013) );
  OR2_X1 U10373 ( .A1(n8015), .A2(n8014), .ZN(n8016) );
  NAND2_X1 U10374 ( .A1(n8026), .A2(n8016), .ZN(n11546) );
  NAND2_X1 U10375 ( .A1(n11546), .A2(n9234), .ZN(n8018) );
  NAND2_X1 U10376 ( .A1(n7974), .A2(n8074), .ZN(n8052) );
  XNOR2_X1 U10377 ( .A(n8030), .B(P2_IR_REG_15__SCAN_IN), .ZN(n15426) );
  AOI22_X1 U10378 ( .A1(n8396), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n15426), 
        .B2(n7821), .ZN(n8017) );
  INV_X1 U10379 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n12265) );
  INV_X1 U10380 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n8019) );
  INV_X1 U10381 ( .A(n8035), .ZN(n8037) );
  NAND2_X1 U10382 ( .A1(n8020), .A2(n8019), .ZN(n8021) );
  NAND2_X1 U10383 ( .A1(n8037), .A2(n8021), .ZN(n12308) );
  OR2_X1 U10384 ( .A1(n12308), .A2(n8338), .ZN(n8023) );
  AOI22_X1 U10385 ( .A1(n9220), .A2(P2_REG0_REG_15__SCAN_IN), .B1(n9219), .B2(
        P2_REG1_REG_15__SCAN_IN), .ZN(n8022) );
  OAI211_X1 U10386 ( .C1(n9223), .C2(n12265), .A(n8023), .B(n8022), .ZN(n13643) );
  INV_X1 U10387 ( .A(n13643), .ZN(n8317) );
  XNOR2_X1 U10388 ( .A(n12310), .B(n8317), .ZN(n12257) );
  INV_X1 U10389 ( .A(n12257), .ZN(n12268) );
  OR2_X1 U10390 ( .A1(n12310), .A2(n13643), .ZN(n8024) );
  MUX2_X1 U10391 ( .A(n11691), .B(n11689), .S(n6671), .Z(n8027) );
  NAND2_X1 U10392 ( .A1(n8027), .A2(n10711), .ZN(n8045) );
  INV_X1 U10393 ( .A(n8027), .ZN(n8028) );
  NAND2_X1 U10394 ( .A1(n8028), .A2(SI_16_), .ZN(n8029) );
  XNOR2_X1 U10395 ( .A(n8044), .B(n8043), .ZN(n11688) );
  NAND2_X1 U10396 ( .A1(n11688), .A2(n9234), .ZN(n8034) );
  INV_X1 U10397 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n8073) );
  NAND2_X1 U10398 ( .A1(n8030), .A2(n8073), .ZN(n8031) );
  XNOR2_X1 U10399 ( .A(n8032), .B(P2_IR_REG_16__SCAN_IN), .ZN(n15436) );
  AOI22_X1 U10400 ( .A1(n8396), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n15436), 
        .B2(n7821), .ZN(n8033) );
  INV_X1 U10401 ( .A(n8056), .ZN(n8058) );
  INV_X1 U10402 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n8036) );
  NAND2_X1 U10403 ( .A1(n8037), .A2(n8036), .ZN(n8038) );
  NAND2_X1 U10404 ( .A1(n8058), .A2(n8038), .ZN(n12473) );
  AOI22_X1 U10405 ( .A1(n9220), .A2(P2_REG0_REG_16__SCAN_IN), .B1(n9219), .B2(
        P2_REG1_REG_16__SCAN_IN), .ZN(n8040) );
  INV_X1 U10406 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n12393) );
  OR2_X1 U10407 ( .A1(n9223), .A2(n12393), .ZN(n8039) );
  OAI211_X1 U10408 ( .C1(n12473), .C2(n8338), .A(n8040), .B(n8039), .ZN(n13642) );
  NAND2_X1 U10409 ( .A1(n12475), .A2(n13642), .ZN(n8042) );
  OR2_X1 U10410 ( .A1(n12475), .A2(n13642), .ZN(n8041) );
  NAND2_X1 U10411 ( .A1(n8042), .A2(n8041), .ZN(n12389) );
  NAND2_X1 U10412 ( .A1(n8044), .A2(n8043), .ZN(n8046) );
  MUX2_X1 U10413 ( .A(n11733), .B(n11735), .S(n6671), .Z(n8047) );
  INV_X1 U10414 ( .A(n8047), .ZN(n8048) );
  NAND2_X1 U10415 ( .A1(n8048), .A2(SI_17_), .ZN(n8049) );
  XNOR2_X1 U10416 ( .A(n8070), .B(n8069), .ZN(n11732) );
  NAND2_X1 U10417 ( .A1(n11732), .A2(n9234), .ZN(n8055) );
  INV_X1 U10418 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n8050) );
  NAND2_X1 U10419 ( .A1(n8073), .A2(n8050), .ZN(n8051) );
  XNOR2_X1 U10420 ( .A(n8053), .B(P2_IR_REG_17__SCAN_IN), .ZN(n15454) );
  AOI22_X1 U10421 ( .A1(n8396), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n15454), 
        .B2(n7821), .ZN(n8054) );
  INV_X1 U10422 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8057) );
  NAND2_X1 U10423 ( .A1(n8058), .A2(n8057), .ZN(n8059) );
  NAND2_X1 U10424 ( .A1(n8105), .A2(n8059), .ZN(n12428) );
  OR2_X1 U10425 ( .A1(n12428), .A2(n8338), .ZN(n8065) );
  INV_X1 U10426 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8062) );
  NAND2_X1 U10427 ( .A1(n9220), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n8061) );
  INV_X1 U10428 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n14007) );
  OR2_X1 U10429 ( .A1(n8402), .A2(n14007), .ZN(n8060) );
  OAI211_X1 U10430 ( .C1(n8062), .C2(n9223), .A(n8061), .B(n8060), .ZN(n8063)
         );
  INV_X1 U10431 ( .A(n8063), .ZN(n8064) );
  NAND2_X1 U10432 ( .A1(n8065), .A2(n8064), .ZN(n13641) );
  XNOR2_X1 U10433 ( .A(n13443), .B(n13641), .ZN(n12423) );
  INV_X1 U10434 ( .A(n12423), .ZN(n8066) );
  NAND2_X1 U10435 ( .A1(n12422), .A2(n8066), .ZN(n8068) );
  NAND2_X1 U10436 ( .A1(n13443), .A2(n13641), .ZN(n8067) );
  NAND2_X1 U10437 ( .A1(n8070), .A2(n8069), .ZN(n8072) );
  INV_X1 U10438 ( .A(SI_18_), .ZN(n10879) );
  XNOR2_X1 U10439 ( .A(n8117), .B(n10879), .ZN(n8090) );
  MUX2_X1 U10440 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(P1_DATAO_REG_18__SCAN_IN), 
        .S(n6671), .Z(n8118) );
  XNOR2_X1 U10441 ( .A(n8090), .B(n8118), .ZN(n11979) );
  NAND2_X1 U10442 ( .A1(n11979), .A2(n9234), .ZN(n8083) );
  NOR2_X1 U10443 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), 
        .ZN(n8075) );
  MUX2_X1 U10444 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8078), .S(
        P2_IR_REG_18__SCAN_IN), .Z(n8079) );
  INV_X1 U10445 ( .A(n8079), .ZN(n8081) );
  NOR2_X1 U10446 ( .A1(n8081), .A2(n8097), .ZN(n13710) );
  AOI22_X1 U10447 ( .A1(n8396), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n13710), 
        .B2(n7821), .ZN(n8082) );
  XNOR2_X1 U10448 ( .A(n8105), .B(P2_REG3_REG_18__SCAN_IN), .ZN(n13601) );
  NAND2_X1 U10449 ( .A1(n13601), .A2(n8253), .ZN(n8088) );
  INV_X1 U10450 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n13918) );
  NAND2_X1 U10451 ( .A1(n9220), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n8085) );
  INV_X1 U10452 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n13699) );
  OR2_X1 U10453 ( .A1(n8402), .A2(n13699), .ZN(n8084) );
  OAI211_X1 U10454 ( .C1(n13918), .C2(n9223), .A(n8085), .B(n8084), .ZN(n8086)
         );
  INV_X1 U10455 ( .A(n8086), .ZN(n8087) );
  NAND2_X1 U10456 ( .A1(n8088), .A2(n8087), .ZN(n13640) );
  INV_X1 U10457 ( .A(n13640), .ZN(n9160) );
  XNOR2_X1 U10458 ( .A(n14053), .B(n9160), .ZN(n13904) );
  INV_X1 U10459 ( .A(n13904), .ZN(n13908) );
  OR2_X1 U10460 ( .A1(n14053), .A2(n13640), .ZN(n8089) );
  INV_X1 U10461 ( .A(n8090), .ZN(n8092) );
  NOR2_X1 U10462 ( .A1(n8117), .A2(n10879), .ZN(n8091) );
  AOI21_X1 U10463 ( .B1(n8092), .B2(n8118), .A(n8091), .ZN(n8096) );
  MUX2_X1 U10464 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n6671), .Z(n8093) );
  NAND2_X1 U10465 ( .A1(n8093), .A2(SI_19_), .ZN(n8121) );
  INV_X1 U10466 ( .A(n8093), .ZN(n8094) );
  INV_X1 U10467 ( .A(SI_19_), .ZN(n11119) );
  NAND2_X1 U10468 ( .A1(n8094), .A2(n11119), .ZN(n8119) );
  AND2_X1 U10469 ( .A1(n8121), .A2(n8119), .ZN(n8095) );
  XNOR2_X1 U10470 ( .A(n8096), .B(n8095), .ZN(n12025) );
  NAND2_X1 U10471 ( .A1(n12025), .A2(n9234), .ZN(n8101) );
  INV_X1 U10472 ( .A(n8097), .ZN(n8277) );
  NAND2_X1 U10473 ( .A1(n8277), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8099) );
  INV_X1 U10474 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n8098) );
  XNOR2_X2 U10475 ( .A(n8099), .B(n8098), .ZN(n13718) );
  INV_X1 U10476 ( .A(n13718), .ZN(n9289) );
  AOI22_X1 U10477 ( .A1(n8396), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n9289), 
        .B2(n7821), .ZN(n8100) );
  INV_X1 U10478 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n8103) );
  INV_X1 U10479 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n8102) );
  OAI21_X1 U10480 ( .B1(n8105), .B2(n8103), .A(n8102), .ZN(n8106) );
  NAND2_X1 U10481 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(P2_REG3_REG_19__SCAN_IN), 
        .ZN(n8104) );
  NAND2_X1 U10482 ( .A1(n8106), .A2(n8128), .ZN(n13888) );
  OR2_X1 U10483 ( .A1(n13888), .A2(n8338), .ZN(n8111) );
  INV_X1 U10484 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n13889) );
  NAND2_X1 U10485 ( .A1(n9220), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n8108) );
  NAND2_X1 U10486 ( .A1(n9219), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n8107) );
  OAI211_X1 U10487 ( .C1(n9223), .C2(n13889), .A(n8108), .B(n8107), .ZN(n8109)
         );
  INV_X1 U10488 ( .A(n8109), .ZN(n8110) );
  NAND2_X1 U10489 ( .A1(n8111), .A2(n8110), .ZN(n13639) );
  OR2_X1 U10490 ( .A1(n13893), .A2(n13639), .ZN(n8112) );
  INV_X1 U10491 ( .A(n8118), .ZN(n8114) );
  OAI21_X1 U10492 ( .B1(n10879), .B2(n8114), .A(n8121), .ZN(n8115) );
  INV_X1 U10493 ( .A(n8115), .ZN(n8116) );
  NOR2_X1 U10494 ( .A1(n8118), .A2(SI_18_), .ZN(n8122) );
  INV_X1 U10495 ( .A(n8119), .ZN(n8120) );
  AOI21_X1 U10496 ( .B1(n8122), .B2(n8121), .A(n8120), .ZN(n8123) );
  INV_X1 U10497 ( .A(SI_20_), .ZN(n11515) );
  MUX2_X1 U10498 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(P1_DATAO_REG_20__SCAN_IN), 
        .S(n6671), .Z(n8135) );
  NAND2_X1 U10499 ( .A1(n12015), .A2(n9234), .ZN(n8126) );
  NAND2_X1 U10500 ( .A1(n8396), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8125) );
  INV_X1 U10501 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n8127) );
  NAND2_X1 U10502 ( .A1(n8128), .A2(n8127), .ZN(n8129) );
  NAND2_X1 U10503 ( .A1(n8152), .A2(n8129), .ZN(n13877) );
  INV_X1 U10504 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n13878) );
  NAND2_X1 U10505 ( .A1(n9220), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n8131) );
  NAND2_X1 U10506 ( .A1(n9219), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n8130) );
  OAI211_X1 U10507 ( .C1(n13878), .C2(n9223), .A(n8131), .B(n8130), .ZN(n8132)
         );
  INV_X1 U10508 ( .A(n8132), .ZN(n8133) );
  OAI21_X1 U10509 ( .B1(n13877), .B2(n8338), .A(n8133), .ZN(n13638) );
  NAND2_X1 U10510 ( .A1(n13986), .A2(n13638), .ZN(n8134) );
  INV_X1 U10511 ( .A(n8135), .ZN(n8136) );
  MUX2_X1 U10512 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n6671), .Z(n8147) );
  XNOR2_X1 U10513 ( .A(n8147), .B(SI_21_), .ZN(n8145) );
  NAND2_X1 U10514 ( .A1(n12153), .A2(n9234), .ZN(n8139) );
  NAND2_X1 U10515 ( .A1(n8396), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n8138) );
  XNOR2_X1 U10516 ( .A(n8152), .B(P2_REG3_REG_21__SCAN_IN), .ZN(n13855) );
  NAND2_X1 U10517 ( .A1(n13855), .A2(n8253), .ZN(n8144) );
  INV_X1 U10518 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n13857) );
  NAND2_X1 U10519 ( .A1(n9220), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n8141) );
  NAND2_X1 U10520 ( .A1(n9219), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n8140) );
  OAI211_X1 U10521 ( .C1(n13857), .C2(n9223), .A(n8141), .B(n8140), .ZN(n8142)
         );
  INV_X1 U10522 ( .A(n8142), .ZN(n8143) );
  NAND2_X1 U10523 ( .A1(n8144), .A2(n8143), .ZN(n13637) );
  XNOR2_X1 U10524 ( .A(n13859), .B(n13637), .ZN(n13861) );
  INV_X1 U10525 ( .A(n8145), .ZN(n8146) );
  MUX2_X1 U10526 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .S(n6671), .Z(n8183) );
  XNOR2_X1 U10527 ( .A(n9628), .B(n8183), .ZN(n12530) );
  NAND2_X1 U10528 ( .A1(n12530), .A2(n9234), .ZN(n8149) );
  NAND2_X1 U10529 ( .A1(n8396), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n8148) );
  AND2_X1 U10530 ( .A1(P2_REG3_REG_22__SCAN_IN), .A2(P2_REG3_REG_21__SCAN_IN), 
        .ZN(n8150) );
  INV_X1 U10531 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n13548) );
  INV_X1 U10532 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n13593) );
  OAI21_X1 U10533 ( .B1(n8152), .B2(n13548), .A(n13593), .ZN(n8153) );
  AND2_X1 U10534 ( .A1(n8169), .A2(n8153), .ZN(n13843) );
  NAND2_X1 U10535 ( .A1(n13843), .A2(n8253), .ZN(n8158) );
  INV_X1 U10536 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n13846) );
  NAND2_X1 U10537 ( .A1(n9220), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n8155) );
  NAND2_X1 U10538 ( .A1(n9219), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n8154) );
  OAI211_X1 U10539 ( .C1(n13846), .C2(n9223), .A(n8155), .B(n8154), .ZN(n8156)
         );
  INV_X1 U10540 ( .A(n8156), .ZN(n8157) );
  NAND2_X1 U10541 ( .A1(n8158), .A2(n8157), .ZN(n13636) );
  INV_X1 U10542 ( .A(n13636), .ZN(n13505) );
  XNOR2_X1 U10543 ( .A(n13975), .B(n13505), .ZN(n13848) );
  NAND2_X1 U10544 ( .A1(n13849), .A2(n13848), .ZN(n13847) );
  NAND2_X1 U10545 ( .A1(n13975), .A2(n13636), .ZN(n8159) );
  INV_X1 U10546 ( .A(n9628), .ZN(n8160) );
  NAND2_X1 U10547 ( .A1(n8160), .A2(n8183), .ZN(n8162) );
  NAND2_X1 U10548 ( .A1(n8182), .A2(SI_22_), .ZN(n8161) );
  NAND2_X1 U10549 ( .A1(n8162), .A2(n8161), .ZN(n8164) );
  MUX2_X1 U10550 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n6671), .Z(n8185) );
  XNOR2_X1 U10551 ( .A(n8185), .B(SI_23_), .ZN(n8163) );
  NAND2_X1 U10552 ( .A1(n12301), .A2(n9234), .ZN(n8166) );
  NAND2_X1 U10553 ( .A1(n8396), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n8165) );
  INV_X1 U10554 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8168) );
  NAND2_X1 U10555 ( .A1(n8169), .A2(n8168), .ZN(n8170) );
  NAND2_X1 U10556 ( .A1(n8192), .A2(n8170), .ZN(n13832) );
  OR2_X1 U10557 ( .A1(n13832), .A2(n8338), .ZN(n8175) );
  INV_X1 U10558 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n13823) );
  NAND2_X1 U10559 ( .A1(n9220), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n8172) );
  NAND2_X1 U10560 ( .A1(n9219), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n8171) );
  OAI211_X1 U10561 ( .C1(n9223), .C2(n13823), .A(n8172), .B(n8171), .ZN(n8173)
         );
  INV_X1 U10562 ( .A(n8173), .ZN(n8174) );
  NAND2_X1 U10563 ( .A1(n8175), .A2(n8174), .ZN(n13635) );
  INV_X1 U10564 ( .A(n13635), .ZN(n8176) );
  NAND2_X1 U10565 ( .A1(n13970), .A2(n8176), .ZN(n8328) );
  OR2_X1 U10566 ( .A1(n13970), .A2(n8176), .ZN(n8177) );
  OR2_X1 U10567 ( .A1(n13970), .A2(n13635), .ZN(n8178) );
  INV_X1 U10568 ( .A(n8185), .ZN(n8179) );
  INV_X1 U10569 ( .A(SI_23_), .ZN(n11829) );
  NAND2_X1 U10570 ( .A1(n8179), .A2(n11829), .ZN(n8186) );
  OAI21_X1 U10571 ( .B1(SI_22_), .B2(n8183), .A(n8186), .ZN(n8180) );
  INV_X1 U10572 ( .A(n8180), .ZN(n8181) );
  INV_X1 U10573 ( .A(n8183), .ZN(n8184) );
  INV_X1 U10574 ( .A(SI_22_), .ZN(n10097) );
  NOR2_X1 U10575 ( .A1(n8184), .A2(n10097), .ZN(n8187) );
  AOI22_X1 U10576 ( .A1(n8187), .A2(n8186), .B1(n8185), .B2(SI_23_), .ZN(n8188) );
  MUX2_X1 U10577 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n6671), .Z(n8203) );
  XNOR2_X1 U10578 ( .A(n8202), .B(n8203), .ZN(n12325) );
  NAND2_X1 U10579 ( .A1(n12325), .A2(n9234), .ZN(n8191) );
  NAND2_X1 U10580 ( .A1(n8396), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n8190) );
  INV_X1 U10581 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n13572) );
  NAND2_X1 U10582 ( .A1(n8192), .A2(n13572), .ZN(n8193) );
  AND2_X1 U10583 ( .A1(n8213), .A2(n8193), .ZN(n13813) );
  NAND2_X1 U10584 ( .A1(n13813), .A2(n8253), .ZN(n8199) );
  INV_X1 U10585 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n8196) );
  NAND2_X1 U10586 ( .A1(n9220), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n8195) );
  NAND2_X1 U10587 ( .A1(n9219), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n8194) );
  OAI211_X1 U10588 ( .C1(n8196), .C2(n9223), .A(n8195), .B(n8194), .ZN(n8197)
         );
  INV_X1 U10589 ( .A(n8197), .ZN(n8198) );
  NAND2_X1 U10590 ( .A1(n8199), .A2(n8198), .ZN(n13634) );
  INV_X1 U10591 ( .A(n13634), .ZN(n13555) );
  NAND2_X1 U10592 ( .A1(n13965), .A2(n13555), .ZN(n13785) );
  OR2_X1 U10593 ( .A1(n13965), .A2(n13555), .ZN(n8200) );
  NAND2_X1 U10594 ( .A1(n13785), .A2(n8200), .ZN(n13809) );
  NAND2_X1 U10595 ( .A1(n13965), .A2(n13634), .ZN(n8201) );
  NAND2_X1 U10596 ( .A1(n8204), .A2(SI_24_), .ZN(n8205) );
  INV_X1 U10597 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n12381) );
  INV_X1 U10598 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n12384) );
  MUX2_X1 U10599 ( .A(n12381), .B(n12384), .S(n6671), .Z(n8206) );
  INV_X1 U10600 ( .A(SI_25_), .ZN(n12216) );
  NAND2_X1 U10601 ( .A1(n8206), .A2(n12216), .ZN(n8223) );
  INV_X1 U10602 ( .A(n8206), .ZN(n8207) );
  NAND2_X1 U10603 ( .A1(n8207), .A2(SI_25_), .ZN(n8208) );
  NAND2_X1 U10604 ( .A1(n8223), .A2(n8208), .ZN(n8221) );
  XNOR2_X1 U10605 ( .A(n8222), .B(n8221), .ZN(n12379) );
  NAND2_X1 U10606 ( .A1(n12379), .A2(n9234), .ZN(n8210) );
  NAND2_X1 U10607 ( .A1(n8396), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n8209) );
  INV_X1 U10608 ( .A(n8213), .ZN(n8211) );
  NAND2_X1 U10609 ( .A1(n8211), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n8228) );
  INV_X1 U10610 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8212) );
  NAND2_X1 U10611 ( .A1(n8213), .A2(n8212), .ZN(n8214) );
  NAND2_X1 U10612 ( .A1(n8228), .A2(n8214), .ZN(n13795) );
  OR2_X1 U10613 ( .A1(n13795), .A2(n8338), .ZN(n8219) );
  INV_X1 U10614 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n13794) );
  NAND2_X1 U10615 ( .A1(n9220), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n8216) );
  NAND2_X1 U10616 ( .A1(n9219), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n8215) );
  OAI211_X1 U10617 ( .C1(n13794), .C2(n9223), .A(n8216), .B(n8215), .ZN(n8217)
         );
  INV_X1 U10618 ( .A(n8217), .ZN(n8218) );
  XNOR2_X1 U10619 ( .A(n13797), .B(n13633), .ZN(n9282) );
  NAND2_X1 U10620 ( .A1(n14041), .A2(n13486), .ZN(n8220) );
  NAND2_X1 U10621 ( .A1(n13790), .A2(n8220), .ZN(n13771) );
  INV_X1 U10622 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n14890) );
  INV_X1 U10623 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n8894) );
  MUX2_X1 U10624 ( .A(n14890), .B(n8894), .S(n6671), .Z(n8239) );
  XNOR2_X1 U10625 ( .A(n8239), .B(SI_26_), .ZN(n8225) );
  NAND2_X1 U10626 ( .A1(n12478), .A2(n9234), .ZN(n8227) );
  NAND2_X1 U10627 ( .A1(n8396), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n8226) );
  INV_X1 U10628 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n13620) );
  NAND2_X1 U10629 ( .A1(n8228), .A2(n13620), .ZN(n8229) );
  NAND2_X1 U10630 ( .A1(n13779), .A2(n8253), .ZN(n8235) );
  INV_X1 U10631 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8232) );
  NAND2_X1 U10632 ( .A1(n9220), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n8231) );
  NAND2_X1 U10633 ( .A1(n9219), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n8230) );
  OAI211_X1 U10634 ( .C1(n9223), .C2(n8232), .A(n8231), .B(n8230), .ZN(n8233)
         );
  INV_X1 U10635 ( .A(n8233), .ZN(n8234) );
  NAND2_X1 U10636 ( .A1(n8235), .A2(n8234), .ZN(n13632) );
  NAND2_X1 U10637 ( .A1(n13778), .A2(n13632), .ZN(n8236) );
  OR2_X1 U10638 ( .A1(n13778), .A2(n13632), .ZN(n8237) );
  INV_X1 U10639 ( .A(SI_26_), .ZN(n12290) );
  MUX2_X1 U10640 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(P1_DATAO_REG_27__SCAN_IN), 
        .S(n6671), .Z(n8257) );
  INV_X1 U10641 ( .A(n8257), .ZN(n8243) );
  XNOR2_X1 U10642 ( .A(n8243), .B(SI_27_), .ZN(n8244) );
  INV_X1 U10643 ( .A(n8247), .ZN(n8245) );
  INV_X1 U10644 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n8246) );
  NAND2_X1 U10645 ( .A1(n8247), .A2(n8246), .ZN(n8248) );
  INV_X1 U10646 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n8251) );
  NAND2_X1 U10647 ( .A1(n9220), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n8250) );
  NAND2_X1 U10648 ( .A1(n9219), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n8249) );
  OAI211_X1 U10649 ( .C1(n8251), .C2(n9223), .A(n8250), .B(n8249), .ZN(n8252)
         );
  INV_X1 U10650 ( .A(n13616), .ZN(n13631) );
  OR2_X1 U10651 ( .A1(n13766), .A2(n13616), .ZN(n8254) );
  NOR2_X1 U10652 ( .A1(n8257), .A2(SI_27_), .ZN(n8255) );
  NAND2_X1 U10653 ( .A1(n8257), .A2(SI_27_), .ZN(n8258) );
  MUX2_X1 U10654 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(P1_DATAO_REG_28__SCAN_IN), 
        .S(n6671), .Z(n8393) );
  XNOR2_X1 U10655 ( .A(n8393), .B(SI_28_), .ZN(n8391) );
  NAND2_X1 U10656 ( .A1(n12661), .A2(n9234), .ZN(n8261) );
  NAND2_X1 U10657 ( .A1(n8396), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n8260) );
  NAND2_X1 U10658 ( .A1(n8262), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n13740) );
  INV_X1 U10659 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8263) );
  NAND2_X1 U10660 ( .A1(n8264), .A2(n8263), .ZN(n8265) );
  NAND2_X1 U10661 ( .A1(n13740), .A2(n8265), .ZN(n13750) );
  INV_X1 U10662 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n13748) );
  NAND2_X1 U10663 ( .A1(n9219), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n8267) );
  NAND2_X1 U10664 ( .A1(n9220), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n8266) );
  OAI211_X1 U10665 ( .C1(n13748), .C2(n9223), .A(n8267), .B(n8266), .ZN(n8268)
         );
  INV_X1 U10666 ( .A(n8268), .ZN(n8269) );
  NAND2_X1 U10667 ( .A1(n13541), .A2(n13536), .ZN(n8271) );
  NAND2_X1 U10668 ( .A1(n8274), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8275) );
  NAND2_X2 U10669 ( .A1(n8276), .A2(n8282), .ZN(n8332) );
  INV_X1 U10670 ( .A(n8332), .ZN(n8280) );
  INV_X1 U10671 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n8278) );
  XNOR2_X1 U10672 ( .A(n8279), .B(n8278), .ZN(n8286) );
  AND2_X1 U10673 ( .A1(n9289), .A2(n12137), .ZN(n8287) );
  NAND2_X1 U10674 ( .A1(n12531), .A2(n8287), .ZN(n15511) );
  NAND2_X1 U10675 ( .A1(n11052), .A2(n15511), .ZN(n15491) );
  INV_X1 U10676 ( .A(n15491), .ZN(n14022) );
  INV_X1 U10677 ( .A(n13639), .ZN(n13578) );
  NAND2_X1 U10678 ( .A1(n13893), .A2(n13578), .ZN(n8324) );
  OR2_X1 U10679 ( .A1(n13893), .A2(n13578), .ZN(n8288) );
  NAND2_X1 U10680 ( .A1(n8324), .A2(n8288), .ZN(n13895) );
  INV_X1 U10681 ( .A(n9025), .ZN(n8290) );
  NAND2_X1 U10682 ( .A1(n8290), .A2(n11053), .ZN(n9031) );
  OAI22_X1 U10683 ( .A1(n10825), .A2(n9031), .B1(n11459), .B2(n13658), .ZN(
        n10859) );
  NAND2_X1 U10684 ( .A1(n10859), .A2(n10858), .ZN(n8292) );
  NAND2_X1 U10685 ( .A1(n11129), .A2(n7492), .ZN(n8291) );
  NAND2_X1 U10686 ( .A1(n8292), .A2(n8291), .ZN(n10869) );
  INV_X1 U10687 ( .A(n10864), .ZN(n10868) );
  NAND2_X1 U10688 ( .A1(n10869), .A2(n10868), .ZN(n8294) );
  NAND2_X1 U10689 ( .A1(n13515), .A2(n11090), .ZN(n8293) );
  NAND2_X1 U10690 ( .A1(n8294), .A2(n8293), .ZN(n11088) );
  INV_X1 U10691 ( .A(n13654), .ZN(n10870) );
  NAND2_X1 U10692 ( .A1(n11400), .A2(n10870), .ZN(n8295) );
  XNOR2_X1 U10693 ( .A(n11523), .B(n13653), .ZN(n11526) );
  NAND2_X1 U10694 ( .A1(n11577), .A2(n11576), .ZN(n8297) );
  NAND2_X1 U10695 ( .A1(n11429), .A2(n9075), .ZN(n8296) );
  INV_X1 U10696 ( .A(n11599), .ZN(n8298) );
  NAND2_X1 U10697 ( .A1(n11600), .A2(n8298), .ZN(n8301) );
  NAND2_X1 U10698 ( .A1(n11594), .A2(n8299), .ZN(n8300) );
  INV_X1 U10699 ( .A(n11638), .ZN(n11645) );
  NAND2_X1 U10700 ( .A1(n11662), .A2(n8302), .ZN(n8303) );
  INV_X1 U10701 ( .A(n13649), .ZN(n9088) );
  AND2_X1 U10702 ( .A1(n11755), .A2(n9088), .ZN(n8304) );
  OR2_X1 U10703 ( .A1(n11755), .A2(n9088), .ZN(n8305) );
  XNOR2_X1 U10704 ( .A(n12068), .B(n13647), .ZN(n11892) );
  INV_X1 U10705 ( .A(n13647), .ZN(n8307) );
  NAND2_X1 U10706 ( .A1(n12068), .A2(n8307), .ZN(n8308) );
  INV_X1 U10707 ( .A(n13646), .ZN(n9269) );
  OR2_X1 U10708 ( .A1(n14019), .A2(n9269), .ZN(n8309) );
  NAND2_X1 U10709 ( .A1(n11964), .A2(n8309), .ZN(n8311) );
  NAND2_X1 U10710 ( .A1(n14019), .A2(n9269), .ZN(n8310) );
  INV_X1 U10711 ( .A(n13645), .ZN(n9268) );
  AND2_X1 U10712 ( .A1(n12090), .A2(n9268), .ZN(n8312) );
  OR2_X1 U10713 ( .A1(n12090), .A2(n9268), .ZN(n8313) );
  INV_X1 U10714 ( .A(n13644), .ZN(n8314) );
  NOR2_X1 U10715 ( .A1(n12277), .A2(n8314), .ZN(n8315) );
  INV_X1 U10716 ( .A(n12277), .ZN(n12205) );
  AND2_X1 U10717 ( .A1(n12310), .A2(n8317), .ZN(n8316) );
  OR2_X1 U10718 ( .A1(n12310), .A2(n8317), .ZN(n8318) );
  NAND2_X1 U10719 ( .A1(n8319), .A2(n8318), .ZN(n12388) );
  INV_X1 U10720 ( .A(n13642), .ZN(n8320) );
  OR2_X1 U10721 ( .A1(n12475), .A2(n8320), .ZN(n8321) );
  INV_X1 U10722 ( .A(n13641), .ZN(n9146) );
  NAND2_X1 U10723 ( .A1(n13443), .A2(n9146), .ZN(n8323) );
  NAND2_X1 U10724 ( .A1(n13898), .A2(n8324), .ZN(n13873) );
  INV_X1 U10725 ( .A(n13638), .ZN(n8325) );
  NAND2_X1 U10726 ( .A1(n13986), .A2(n8325), .ZN(n8327) );
  OR2_X1 U10727 ( .A1(n13986), .A2(n8325), .ZN(n8326) );
  NAND2_X1 U10728 ( .A1(n8327), .A2(n8326), .ZN(n9279) );
  INV_X1 U10729 ( .A(n13637), .ZN(n13579) );
  OR2_X1 U10730 ( .A1(n13975), .A2(n13505), .ZN(n13826) );
  INV_X1 U10731 ( .A(n13632), .ZN(n13556) );
  OR2_X1 U10732 ( .A1(n13778), .A2(n13556), .ZN(n9267) );
  NAND2_X1 U10733 ( .A1(n13773), .A2(n9267), .ZN(n8329) );
  NAND2_X1 U10734 ( .A1(n13778), .A2(n13556), .ZN(n9266) );
  NAND2_X1 U10735 ( .A1(n8329), .A2(n9266), .ZN(n13756) );
  NAND2_X1 U10736 ( .A1(n13756), .A2(n13760), .ZN(n8331) );
  OR2_X1 U10737 ( .A1(n13766), .A2(n13631), .ZN(n8330) );
  NAND2_X1 U10738 ( .A1(n8331), .A2(n8330), .ZN(n8336) );
  NOR2_X1 U10739 ( .A1(n12531), .A2(n13718), .ZN(n9027) );
  AND2_X1 U10740 ( .A1(n9291), .A2(n8333), .ZN(n8334) );
  NAND2_X1 U10741 ( .A1(n8336), .A2(n8335), .ZN(n8337) );
  NAND3_X1 U10742 ( .A1(n8401), .A2(n13906), .A3(n8337), .ZN(n8351) );
  OR2_X1 U10743 ( .A1(n13740), .A2(n8338), .ZN(n8343) );
  INV_X1 U10744 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n13739) );
  NAND2_X1 U10745 ( .A1(n9219), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n8340) );
  NAND2_X1 U10746 ( .A1(n9220), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n8339) );
  OAI211_X1 U10747 ( .C1(n13739), .C2(n9223), .A(n8340), .B(n8339), .ZN(n8341)
         );
  INV_X1 U10748 ( .A(n8341), .ZN(n8342) );
  OR2_X1 U10749 ( .A1(n8381), .A2(n8344), .ZN(n8345) );
  INV_X1 U10750 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n8346) );
  NAND2_X1 U10751 ( .A1(n8407), .A2(n8346), .ZN(n8347) );
  NAND2_X1 U10752 ( .A1(n8347), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8348) );
  XNOR2_X1 U10753 ( .A(n8348), .B(P2_IR_REG_28__SCAN_IN), .ZN(n10505) );
  NOR2_X1 U10754 ( .A1(n12531), .A2(n8332), .ZN(n10501) );
  INV_X1 U10755 ( .A(n10501), .ZN(n11048) );
  INV_X1 U10756 ( .A(n13617), .ZN(n13577) );
  OR2_X1 U10757 ( .A1(n13616), .A2(n13577), .ZN(n8349) );
  OAI21_X1 U10758 ( .B1(n9225), .B2(n13615), .A(n8349), .ZN(n13542) );
  INV_X1 U10759 ( .A(n13542), .ZN(n8350) );
  NAND2_X1 U10760 ( .A1(n8351), .A2(n8350), .ZN(n13752) );
  INV_X1 U10761 ( .A(n13778), .ZN(n14037) );
  INV_X1 U10762 ( .A(n12475), .ZN(n14063) );
  INV_X1 U10763 ( .A(n15507), .ZN(n11890) );
  INV_X1 U10764 ( .A(n13515), .ZN(n11144) );
  NAND2_X1 U10765 ( .A1(n10872), .A2(n11144), .ZN(n11085) );
  INV_X1 U10766 ( .A(n11429), .ZN(n15482) );
  INV_X1 U10767 ( .A(n11594), .ZN(n15488) );
  NAND2_X1 U10768 ( .A1(n11890), .A2(n11776), .ZN(n11901) );
  OR2_X2 U10769 ( .A1(n12068), .A2(n11901), .ZN(n11958) );
  NAND2_X1 U10770 ( .A1(n14063), .A2(n12392), .ZN(n12427) );
  NAND2_X1 U10771 ( .A1(n13882), .A2(n14048), .ZN(n13854) );
  OR2_X2 U10772 ( .A1(n13975), .A2(n13854), .ZN(n13841) );
  AND2_X2 U10773 ( .A1(n14032), .A2(n13763), .ZN(n8411) );
  NOR2_X1 U10774 ( .A1(n14032), .A2(n13763), .ZN(n8352) );
  NAND2_X1 U10775 ( .A1(n8358), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8353) );
  MUX2_X1 U10776 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8353), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n8356) );
  INV_X1 U10777 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n8354) );
  NAND2_X1 U10778 ( .A1(n8356), .A2(n8361), .ZN(n12382) );
  NAND2_X1 U10779 ( .A1(n8383), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8357) );
  MUX2_X1 U10780 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8357), .S(
        P2_IR_REG_24__SCAN_IN), .Z(n8359) );
  NAND2_X1 U10781 ( .A1(n8359), .A2(n8358), .ZN(n12326) );
  XNOR2_X1 U10782 ( .A(n12326), .B(P2_B_REG_SCAN_IN), .ZN(n8360) );
  NAND2_X1 U10783 ( .A1(n12382), .A2(n8360), .ZN(n8363) );
  NAND2_X1 U10784 ( .A1(n8361), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8362) );
  NAND2_X1 U10785 ( .A1(n8363), .A2(n12479), .ZN(n8377) );
  NOR4_X1 U10786 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n8372) );
  OR4_X1 U10787 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n8369) );
  NOR4_X1 U10788 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n8367) );
  NOR4_X1 U10789 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n8366) );
  NOR4_X1 U10790 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n8365) );
  NOR4_X1 U10791 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n8364) );
  NAND4_X1 U10792 ( .A1(n8367), .A2(n8366), .A3(n8365), .A4(n8364), .ZN(n8368)
         );
  NOR4_X1 U10793 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        n8369), .A4(n8368), .ZN(n8371) );
  NOR4_X1 U10794 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n8370) );
  AND3_X1 U10795 ( .A1(n8372), .A2(n8371), .A3(n8370), .ZN(n8373) );
  NOR2_X1 U10796 ( .A1(n8377), .A2(n8373), .ZN(n11037) );
  INV_X1 U10797 ( .A(n11037), .ZN(n8375) );
  INV_X1 U10798 ( .A(n12382), .ZN(n8374) );
  OAI22_X1 U10799 ( .A1(n8377), .A2(P2_D_REG_1__SCAN_IN), .B1(n12479), .B2(
        n8374), .ZN(n15469) );
  NOR2_X1 U10800 ( .A1(n15511), .A2(n9291), .ZN(n11044) );
  INV_X1 U10801 ( .A(n11044), .ZN(n11038) );
  NAND3_X1 U10802 ( .A1(n8375), .A2(n15469), .A3(n11038), .ZN(n8418) );
  NAND2_X1 U10803 ( .A1(n10501), .A2(n11045), .ZN(n11040) );
  INV_X1 U10804 ( .A(n11040), .ZN(n8376) );
  NOR2_X1 U10805 ( .A1(n8418), .A2(n8376), .ZN(n8385) );
  INV_X1 U10806 ( .A(n8377), .ZN(n15463) );
  INV_X1 U10807 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n15466) );
  INV_X1 U10808 ( .A(n12326), .ZN(n8378) );
  NOR2_X1 U10809 ( .A1(n12479), .A2(n8378), .ZN(n8379) );
  AOI21_X1 U10810 ( .B1(n15463), .B2(n15466), .A(n8379), .ZN(n11036) );
  NOR2_X1 U10811 ( .A1(n12382), .A2(n12326), .ZN(n8380) );
  NAND2_X1 U10812 ( .A1(n8380), .A2(n12479), .ZN(n10406) );
  MUX2_X1 U10813 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8382), .S(
        P2_IR_REG_23__SCAN_IN), .Z(n8384) );
  NAND2_X1 U10814 ( .A1(n8384), .A2(n8383), .ZN(n10500) );
  NAND2_X1 U10815 ( .A1(n11036), .A2(n15470), .ZN(n15465) );
  NAND2_X1 U10816 ( .A1(n11490), .A2(n11045), .ZN(n15516) );
  NAND2_X1 U10817 ( .A1(n15539), .A2(n15508), .ZN(n14016) );
  NAND2_X1 U10818 ( .A1(n8387), .A2(n8386), .ZN(P2_U3527) );
  NAND2_X1 U10819 ( .A1(n8390), .A2(n8389), .ZN(n8399) );
  INV_X1 U10820 ( .A(n8393), .ZN(n8394) );
  INV_X1 U10821 ( .A(SI_28_), .ZN(n12668) );
  NAND2_X1 U10822 ( .A1(n8394), .A2(n12668), .ZN(n8395) );
  MUX2_X1 U10823 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(P1_DATAO_REG_29__SCAN_IN), 
        .S(n6671), .Z(n9210) );
  INV_X1 U10824 ( .A(SI_29_), .ZN(n13439) );
  XNOR2_X1 U10825 ( .A(n9210), .B(n13439), .ZN(n9208) );
  NAND2_X1 U10826 ( .A1(n14071), .A2(n9234), .ZN(n8398) );
  NAND2_X1 U10827 ( .A1(n8396), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n8397) );
  INV_X1 U10828 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n13944) );
  OR2_X1 U10829 ( .A1(n8402), .A2(n13944), .ZN(n8406) );
  INV_X1 U10830 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n13733) );
  OR2_X1 U10831 ( .A1(n9223), .A2(n13733), .ZN(n8405) );
  INV_X1 U10832 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n14027) );
  OR2_X1 U10833 ( .A1(n8403), .A2(n14027), .ZN(n8404) );
  AND3_X1 U10834 ( .A1(n8406), .A2(n8405), .A3(n8404), .ZN(n9240) );
  XNOR2_X1 U10835 ( .A(n8407), .B(P2_IR_REG_27__SCAN_IN), .ZN(n14081) );
  NAND2_X1 U10836 ( .A1(n14081), .A2(P2_B_REG_SCAN_IN), .ZN(n8408) );
  NAND2_X1 U10837 ( .A1(n13602), .A2(n8408), .ZN(n13727) );
  OAI22_X1 U10838 ( .A1(n13536), .A2(n13577), .B1(n9240), .B2(n13727), .ZN(
        n8409) );
  NAND2_X1 U10839 ( .A1(n9224), .A2(n8411), .ZN(n13723) );
  OAI211_X1 U10840 ( .C1(n9224), .C2(n8411), .A(n11777), .B(n13723), .ZN(
        n13741) );
  OR2_X1 U10841 ( .A1(n8420), .A2(n15536), .ZN(n8416) );
  INV_X1 U10842 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n8413) );
  NAND2_X1 U10843 ( .A1(n8416), .A2(n8415), .ZN(P2_U3528) );
  NAND2_X1 U10844 ( .A1(n15470), .A2(n11040), .ZN(n8417) );
  NOR2_X1 U10845 ( .A1(n8417), .A2(n11036), .ZN(n11384) );
  INV_X1 U10846 ( .A(n8418), .ZN(n8419) );
  OR2_X1 U10847 ( .A1(n8420), .A2(n15523), .ZN(n8425) );
  NAND2_X1 U10848 ( .A1(n15524), .A2(n15508), .ZN(n14062) );
  INV_X1 U10849 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n8421) );
  NOR2_X1 U10850 ( .A1(n15524), .A2(n8421), .ZN(n8422) );
  NAND2_X1 U10851 ( .A1(n8425), .A2(n8424), .ZN(P2_U3496) );
  INV_X1 U10852 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n9009) );
  NOR2_X1 U10853 ( .A1(P3_IR_REG_6__SCAN_IN), .A2(P3_IR_REG_10__SCAN_IN), .ZN(
        n8429) );
  NAND4_X1 U10854 ( .A1(n8429), .A2(n8428), .A3(n8427), .A4(n8568), .ZN(n8440)
         );
  INV_X1 U10855 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n8432) );
  INV_X1 U10856 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n8434) );
  NAND2_X1 U10857 ( .A1(n8970), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8436) );
  INV_X1 U10858 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n8435) );
  NAND2_X1 U10859 ( .A1(n6753), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8437) );
  NAND2_X1 U10860 ( .A1(n6758), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8439) );
  NAND2_X1 U10861 ( .A1(n11514), .A2(n7356), .ZN(n15708) );
  INV_X1 U10862 ( .A(n15708), .ZN(n15689) );
  INV_X1 U10863 ( .A(n8440), .ZN(n8443) );
  NOR2_X1 U10864 ( .A1(P3_IR_REG_22__SCAN_IN), .A2(P3_IR_REG_19__SCAN_IN), 
        .ZN(n8442) );
  NOR2_X1 U10865 ( .A1(P3_IR_REG_20__SCAN_IN), .A2(P3_IR_REG_23__SCAN_IN), 
        .ZN(n8441) );
  INV_X1 U10866 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n8449) );
  NAND2_X1 U10867 ( .A1(n8451), .A2(n8449), .ZN(n13431) );
  INV_X1 U10868 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n8452) );
  NAND2_X2 U10869 ( .A1(n8453), .A2(n8454), .ZN(n8737) );
  INV_X1 U10870 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n11364) );
  OR2_X1 U10871 ( .A1(n8737), .A2(n11364), .ZN(n8457) );
  NAND2_X1 U10872 ( .A1(n8798), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n8456) );
  NAND2_X2 U10873 ( .A1(n8454), .A2(n13437), .ZN(n11986) );
  INV_X1 U10874 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n10911) );
  OR2_X1 U10875 ( .A1(n11986), .A2(n10911), .ZN(n8455) );
  XNOR2_X2 U10876 ( .A(n8460), .B(n8459), .ZN(n12667) );
  INV_X1 U10877 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n8462) );
  NAND2_X1 U10878 ( .A1(n8465), .A2(n6671), .ZN(n8623) );
  OR2_X1 U10879 ( .A1(n8623), .A2(n10454), .ZN(n8468) );
  OR2_X1 U10880 ( .A1(n8811), .A2(n10455), .ZN(n8467) );
  OR2_X1 U10881 ( .A1(n8465), .A2(n7030), .ZN(n8466) );
  INV_X1 U10882 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n8469) );
  OR2_X1 U10883 ( .A1(n11986), .A2(n8469), .ZN(n8474) );
  INV_X1 U10884 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n11305) );
  OR2_X1 U10885 ( .A1(n8737), .A2(n11305), .ZN(n8473) );
  INV_X1 U10886 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n8470) );
  OR2_X1 U10887 ( .A1(n8480), .A2(n8470), .ZN(n8472) );
  NAND2_X1 U10888 ( .A1(n11984), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n8471) );
  OR2_X1 U10889 ( .A1(n8623), .A2(n6886), .ZN(n8478) );
  XNOR2_X1 U10890 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n8487) );
  NAND2_X1 U10891 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), 
        .ZN(n8475) );
  XNOR2_X2 U10892 ( .A(n8475), .B(n7029), .ZN(n11313) );
  OR2_X1 U10893 ( .A1(n8465), .A2(n11313), .ZN(n8476) );
  NAND2_X1 U10894 ( .A1(n9799), .A2(n12845), .ZN(n15679) );
  NAND2_X1 U10895 ( .A1(n11984), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n8485) );
  INV_X1 U10896 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n11173) );
  OR2_X1 U10897 ( .A1(n8737), .A2(n11173), .ZN(n8484) );
  INV_X1 U10898 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n8479) );
  OR2_X1 U10899 ( .A1(n8480), .A2(n8479), .ZN(n8483) );
  INV_X1 U10900 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n8481) );
  NAND2_X1 U10901 ( .A1(n8487), .A2(n8486), .ZN(n8490) );
  NAND2_X1 U10902 ( .A1(n8488), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8489) );
  NAND2_X1 U10903 ( .A1(n8490), .A2(n8489), .ZN(n8502) );
  NAND2_X1 U10904 ( .A1(n10412), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n8503) );
  NAND2_X1 U10905 ( .A1(n10462), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n8491) );
  XNOR2_X1 U10906 ( .A(n8502), .B(n8501), .ZN(n10422) );
  OR2_X1 U10907 ( .A1(n8811), .A2(n10422), .ZN(n8493) );
  OR2_X1 U10908 ( .A1(n8623), .A2(SI_2_), .ZN(n8492) );
  OAI211_X1 U10909 ( .C1(n10967), .C2(n8465), .A(n8493), .B(n8492), .ZN(n15687) );
  NAND2_X1 U10910 ( .A1(n15698), .A2(n15687), .ZN(n12859) );
  INV_X1 U10911 ( .A(n12857), .ZN(n15678) );
  NAND2_X1 U10912 ( .A1(n11984), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n8498) );
  OR2_X1 U10913 ( .A1(n8737), .A2(P3_REG3_REG_3__SCAN_IN), .ZN(n8497) );
  INV_X1 U10914 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n8494) );
  OR2_X1 U10915 ( .A1(n11989), .A2(n8494), .ZN(n8496) );
  INV_X1 U10916 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n12018) );
  OR2_X1 U10917 ( .A1(n11986), .A2(n12018), .ZN(n8495) );
  NAND2_X1 U10918 ( .A1(n8499), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8500) );
  XNOR2_X1 U10919 ( .A(n8500), .B(P3_IR_REG_3__SCAN_IN), .ZN(n10929) );
  NAND2_X1 U10920 ( .A1(n8502), .A2(n8501), .ZN(n8504) );
  NAND2_X1 U10921 ( .A1(n8504), .A2(n8503), .ZN(n8517) );
  NAND2_X1 U10922 ( .A1(n10441), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n8505) );
  XNOR2_X1 U10923 ( .A(n8517), .B(n8516), .ZN(n10445) );
  OR2_X1 U10924 ( .A1(n8811), .A2(n10445), .ZN(n8507) );
  OR2_X1 U10925 ( .A1(n12806), .A2(SI_3_), .ZN(n8506) );
  NAND2_X1 U10926 ( .A1(n8960), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n8513) );
  INV_X1 U10927 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n10981) );
  OR2_X1 U10928 ( .A1(n8524), .A2(n10981), .ZN(n8512) );
  AND2_X1 U10929 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n8508) );
  NOR2_X1 U10930 ( .A1(n8526), .A2(n8508), .ZN(n15676) );
  OR2_X1 U10931 ( .A1(n8737), .A2(n15676), .ZN(n8511) );
  INV_X1 U10932 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n8509) );
  OR2_X1 U10933 ( .A1(n11989), .A2(n8509), .ZN(n8510) );
  NAND4_X1 U10934 ( .A1(n8513), .A2(n8512), .A3(n8511), .A4(n8510), .ZN(n11673) );
  NAND2_X1 U10935 ( .A1(n8514), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8515) );
  NAND2_X1 U10936 ( .A1(n8517), .A2(n8516), .ZN(n8519) );
  NAND2_X1 U10937 ( .A1(n10436), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n8520) );
  XNOR2_X1 U10938 ( .A(n8537), .B(n8536), .ZN(n10414) );
  OR2_X1 U10939 ( .A1(n8811), .A2(n10414), .ZN(n8522) );
  OR2_X1 U10940 ( .A1(n12806), .A2(SI_4_), .ZN(n8521) );
  OAI211_X1 U10941 ( .C1(n10982), .C2(n6852), .A(n8522), .B(n8521), .ZN(n11569) );
  NAND2_X1 U10942 ( .A1(n11673), .A2(n11569), .ZN(n12869) );
  NAND2_X1 U10943 ( .A1(n12868), .A2(n12869), .ZN(n11563) );
  INV_X1 U10944 ( .A(n11563), .ZN(n12863) );
  NAND2_X1 U10945 ( .A1(n11559), .A2(n12868), .ZN(n11672) );
  NAND2_X1 U10946 ( .A1(n8798), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n8532) );
  INV_X1 U10947 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n8523) );
  OR2_X1 U10948 ( .A1(n11986), .A2(n8523), .ZN(n8531) );
  INV_X1 U10949 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n8525) );
  OR2_X1 U10950 ( .A1(n8524), .A2(n8525), .ZN(n8530) );
  NAND2_X1 U10951 ( .A1(n8526), .A2(n8527), .ZN(n8545) );
  OR2_X1 U10952 ( .A1(n8527), .A2(n8526), .ZN(n8528) );
  AND2_X1 U10953 ( .A1(n8545), .A2(n8528), .ZN(n11683) );
  OR2_X1 U10954 ( .A1(n8737), .A2(n11683), .ZN(n8529) );
  NAND4_X1 U10955 ( .A1(n8532), .A2(n8531), .A3(n8530), .A4(n8529), .ZN(n12995) );
  OR2_X1 U10956 ( .A1(n8533), .A2(n8680), .ZN(n8535) );
  XNOR2_X1 U10957 ( .A(n8535), .B(n8534), .ZN(n10995) );
  NAND2_X1 U10958 ( .A1(n10443), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n8539) );
  XNOR2_X1 U10959 ( .A(n8553), .B(n8552), .ZN(n10425) );
  OR2_X1 U10960 ( .A1(n8811), .A2(n10425), .ZN(n8541) );
  OR2_X1 U10961 ( .A1(n12806), .A2(SI_5_), .ZN(n8540) );
  OAI211_X1 U10962 ( .C1(n7022), .C2(n6852), .A(n8541), .B(n8540), .ZN(n11682)
         );
  OR2_X1 U10963 ( .A1(n12995), .A2(n11682), .ZN(n12867) );
  NAND2_X1 U10964 ( .A1(n12995), .A2(n11682), .ZN(n12876) );
  NAND2_X1 U10965 ( .A1(n11672), .A2(n6678), .ZN(n8542) );
  NAND2_X1 U10966 ( .A1(n8542), .A2(n12867), .ZN(n11786) );
  NAND2_X1 U10967 ( .A1(n8798), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n8550) );
  INV_X1 U10968 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n8543) );
  OR2_X1 U10969 ( .A1(n11986), .A2(n8543), .ZN(n8549) );
  INV_X1 U10970 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n8544) );
  OR2_X1 U10971 ( .A1(n8524), .A2(n8544), .ZN(n8548) );
  NAND2_X1 U10972 ( .A1(n8545), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8546) );
  AND2_X1 U10973 ( .A1(n8560), .A2(n8546), .ZN(n15666) );
  OR2_X1 U10974 ( .A1(n8737), .A2(n15666), .ZN(n8547) );
  NAND4_X1 U10975 ( .A1(n8550), .A2(n8549), .A3(n8548), .A4(n8547), .ZN(n11947) );
  XNOR2_X1 U10976 ( .A(n8551), .B(P3_IR_REG_6__SCAN_IN), .ZN(n11153) );
  INV_X1 U10977 ( .A(SI_6_), .ZN(n10452) );
  OR2_X1 U10978 ( .A1(n12806), .A2(n10452), .ZN(n8558) );
  XNOR2_X1 U10979 ( .A(n10431), .B(P2_DATAO_REG_6__SCAN_IN), .ZN(n8556) );
  XNOR2_X1 U10980 ( .A(n8571), .B(n8556), .ZN(n10453) );
  OR2_X1 U10981 ( .A1(n8811), .A2(n10453), .ZN(n8557) );
  OAI211_X1 U10982 ( .C1(n6852), .C2(n11163), .A(n8558), .B(n8557), .ZN(n15664) );
  INV_X1 U10983 ( .A(n15664), .ZN(n11797) );
  NAND2_X1 U10984 ( .A1(n11947), .A2(n11797), .ZN(n12877) );
  NAND2_X1 U10985 ( .A1(n12878), .A2(n12877), .ZN(n8559) );
  NAND2_X1 U10986 ( .A1(n11786), .A2(n12820), .ZN(n11785) );
  NAND2_X1 U10987 ( .A1(n11785), .A2(n12878), .ZN(n11943) );
  NAND2_X1 U10988 ( .A1(n8798), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n8567) );
  AND2_X1 U10989 ( .A1(n8560), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8561) );
  NOR2_X1 U10990 ( .A1(n8580), .A2(n8561), .ZN(n15659) );
  OR2_X1 U10991 ( .A1(n8737), .A2(n15659), .ZN(n8566) );
  INV_X1 U10992 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n8562) );
  OR2_X1 U10993 ( .A1(n8524), .A2(n8562), .ZN(n8565) );
  INV_X1 U10994 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n8563) );
  OR2_X1 U10995 ( .A1(n11986), .A2(n8563), .ZN(n8564) );
  NAND4_X1 U10996 ( .A1(n8567), .A2(n8566), .A3(n8565), .A4(n8564), .ZN(n12031) );
  NAND2_X1 U10997 ( .A1(n6720), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8569) );
  XNOR2_X1 U10998 ( .A(n8569), .B(n8568), .ZN(n11327) );
  INV_X1 U10999 ( .A(n11327), .ZN(n11321) );
  NAND2_X1 U11000 ( .A1(n10438), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n8570) );
  NAND2_X1 U11001 ( .A1(n10431), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n8572) );
  NAND2_X1 U11002 ( .A1(n10458), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n8573) );
  NAND2_X1 U11003 ( .A1(n8587), .A2(n8573), .ZN(n8574) );
  NAND2_X1 U11004 ( .A1(n8575), .A2(n8574), .ZN(n8576) );
  AND2_X1 U11005 ( .A1(n8588), .A2(n8576), .ZN(n10417) );
  OR2_X1 U11006 ( .A1(n8811), .A2(n10417), .ZN(n8578) );
  OR2_X1 U11007 ( .A1(n8623), .A2(SI_7_), .ZN(n8577) );
  OAI211_X1 U11008 ( .C1(n11321), .C2(n6852), .A(n8578), .B(n8577), .ZN(n11953) );
  OR2_X1 U11009 ( .A1(n12031), .A2(n11953), .ZN(n12884) );
  NAND2_X1 U11010 ( .A1(n12031), .A2(n11953), .ZN(n12883) );
  INV_X1 U11011 ( .A(n12819), .ZN(n12880) );
  NAND2_X1 U11012 ( .A1(n11943), .A2(n12880), .ZN(n11942) );
  NAND2_X1 U11013 ( .A1(n11942), .A2(n12884), .ZN(n12032) );
  NAND2_X1 U11014 ( .A1(n8798), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n8585) );
  INV_X1 U11015 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n12041) );
  OR2_X1 U11016 ( .A1(n11986), .A2(n12041), .ZN(n8584) );
  INV_X1 U11017 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n8579) );
  OR2_X1 U11018 ( .A1(n8524), .A2(n8579), .ZN(n8583) );
  NOR2_X1 U11019 ( .A1(n8580), .A2(n11333), .ZN(n8581) );
  OR2_X1 U11020 ( .A1(n8597), .A2(n8581), .ZN(n12039) );
  INV_X1 U11021 ( .A(n12039), .ZN(n11839) );
  OR2_X1 U11022 ( .A1(n8737), .A2(n11839), .ZN(n8582) );
  NAND4_X1 U11023 ( .A1(n8585), .A2(n8584), .A3(n8583), .A4(n8582), .ZN(n12189) );
  NAND2_X1 U11024 ( .A1(n8604), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8586) );
  XNOR2_X1 U11025 ( .A(n8586), .B(P3_IR_REG_8__SCAN_IN), .ZN(n11325) );
  NAND2_X1 U11026 ( .A1(n10469), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n8589) );
  OR2_X1 U11027 ( .A1(n8591), .A2(n8590), .ZN(n8592) );
  NAND2_X1 U11028 ( .A1(n8607), .A2(n8592), .ZN(n10420) );
  OR2_X1 U11029 ( .A1(n8811), .A2(n10420), .ZN(n8594) );
  INV_X1 U11030 ( .A(SI_8_), .ZN(n10421) );
  OR2_X1 U11031 ( .A1(n12806), .A2(n10421), .ZN(n8593) );
  OAI211_X1 U11032 ( .C1(n6852), .C2(n11853), .A(n8594), .B(n8593), .ZN(n11834) );
  INV_X1 U11033 ( .A(n11834), .ZN(n12038) );
  OR2_X1 U11034 ( .A1(n12189), .A2(n12038), .ZN(n12889) );
  NAND2_X1 U11035 ( .A1(n12189), .A2(n12038), .ZN(n12888) );
  NAND2_X1 U11036 ( .A1(n12889), .A2(n12888), .ZN(n12029) );
  NAND2_X1 U11037 ( .A1(n12032), .A2(n12886), .ZN(n12034) );
  NAND2_X1 U11038 ( .A1(n8960), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n8603) );
  INV_X1 U11039 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n8595) );
  OR2_X1 U11040 ( .A1(n8524), .A2(n8595), .ZN(n8602) );
  OR2_X1 U11041 ( .A1(n8597), .A2(n8596), .ZN(n8598) );
  AND2_X1 U11042 ( .A1(n8614), .A2(n8598), .ZN(n12193) );
  OR2_X1 U11043 ( .A1(n8737), .A2(n12193), .ZN(n8601) );
  INV_X1 U11044 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n8599) );
  OR2_X1 U11045 ( .A1(n11989), .A2(n8599), .ZN(n8600) );
  NAND4_X1 U11046 ( .A1(n8603), .A2(n8602), .A3(n8601), .A4(n8600), .ZN(n15639) );
  NOR2_X1 U11047 ( .A1(n8604), .A2(P3_IR_REG_8__SCAN_IN), .ZN(n8631) );
  OR2_X1 U11048 ( .A1(n8631), .A2(n8680), .ZN(n8605) );
  INV_X1 U11049 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n8630) );
  XNOR2_X1 U11050 ( .A(n8605), .B(n8630), .ZN(n15557) );
  OR2_X1 U11051 ( .A1(n12806), .A2(SI_9_), .ZN(n8613) );
  NAND2_X1 U11052 ( .A1(n10488), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n8624) );
  NAND2_X1 U11053 ( .A1(n10490), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n8608) );
  OR2_X1 U11054 ( .A1(n8610), .A2(n8609), .ZN(n8611) );
  AND2_X1 U11055 ( .A1(n8625), .A2(n8611), .ZN(n10428) );
  OR2_X1 U11056 ( .A1(n8811), .A2(n10428), .ZN(n8612) );
  OAI211_X1 U11057 ( .C1(n11857), .C2(n6852), .A(n8613), .B(n8612), .ZN(n15731) );
  NAND2_X1 U11058 ( .A1(n15639), .A2(n15731), .ZN(n12893) );
  OR2_X1 U11059 ( .A1(n15639), .A2(n15731), .ZN(n12894) );
  NAND2_X1 U11060 ( .A1(n8798), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n8622) );
  NAND2_X1 U11061 ( .A1(n8614), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8615) );
  NAND2_X1 U11062 ( .A1(n8648), .A2(n8615), .ZN(n15642) );
  INV_X1 U11063 ( .A(n15642), .ZN(n8616) );
  OR2_X1 U11064 ( .A1(n8737), .A2(n8616), .ZN(n8621) );
  INV_X1 U11065 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n8617) );
  OR2_X1 U11066 ( .A1(n8524), .A2(n8617), .ZN(n8620) );
  INV_X1 U11067 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n8618) );
  OR2_X1 U11068 ( .A1(n11986), .A2(n8618), .ZN(n8619) );
  NAND4_X1 U11069 ( .A1(n8622), .A2(n8621), .A3(n8620), .A4(n8619), .ZN(n15043) );
  NAND2_X1 U11070 ( .A1(n10493), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n8637) );
  NAND2_X1 U11071 ( .A1(n10491), .A2(P2_DATAO_REG_10__SCAN_IN), .ZN(n8626) );
  OR2_X1 U11072 ( .A1(n8628), .A2(n8627), .ZN(n8629) );
  NAND2_X1 U11073 ( .A1(n8638), .A2(n8629), .ZN(n10448) );
  NAND2_X1 U11074 ( .A1(n10448), .A2(n12805), .ZN(n8635) );
  NAND2_X1 U11075 ( .A1(n8631), .A2(n8630), .ZN(n8643) );
  NAND2_X1 U11076 ( .A1(n8643), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8633) );
  INV_X1 U11077 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n8632) );
  XNOR2_X1 U11078 ( .A(n8633), .B(n8632), .ZN(n13011) );
  OR2_X1 U11079 ( .A1(n6852), .A2(n13050), .ZN(n8634) );
  OR2_X1 U11080 ( .A1(n15043), .A2(n15647), .ZN(n12896) );
  NAND2_X1 U11081 ( .A1(n15043), .A2(n15647), .ZN(n12895) );
  INV_X1 U11082 ( .A(n15048), .ZN(n8657) );
  NAND2_X1 U11083 ( .A1(n10497), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n8658) );
  NAND2_X1 U11084 ( .A1(n10499), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n8639) );
  OR2_X1 U11085 ( .A1(n8641), .A2(n8640), .ZN(n8642) );
  NAND2_X1 U11086 ( .A1(n8659), .A2(n8642), .ZN(n10451) );
  NAND2_X1 U11087 ( .A1(n10451), .A2(n12805), .ZN(n8647) );
  OAI21_X1 U11088 ( .B1(n8643), .B2(P3_IR_REG_10__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8645) );
  INV_X1 U11089 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n8644) );
  XNOR2_X1 U11090 ( .A(n8645), .B(n8644), .ZN(n15573) );
  AOI22_X1 U11091 ( .A1(n12799), .A2(n10450), .B1(n10909), .B2(n15573), .ZN(
        n8646) );
  NAND2_X1 U11092 ( .A1(n8647), .A2(n8646), .ZN(n15051) );
  INV_X1 U11093 ( .A(n15051), .ZN(n12184) );
  NAND2_X1 U11094 ( .A1(n8798), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n8655) );
  NAND2_X1 U11095 ( .A1(n8648), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8649) );
  AND2_X1 U11096 ( .A1(n8669), .A2(n8649), .ZN(n15046) );
  OR2_X1 U11097 ( .A1(n8737), .A2(n15046), .ZN(n8654) );
  INV_X1 U11098 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n8650) );
  OR2_X1 U11099 ( .A1(n8524), .A2(n8650), .ZN(n8653) );
  INV_X1 U11100 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n8651) );
  OR2_X1 U11101 ( .A1(n11986), .A2(n8651), .ZN(n8652) );
  OR2_X1 U11102 ( .A1(n12184), .A2(n12372), .ZN(n12902) );
  NAND2_X1 U11103 ( .A1(n12184), .A2(n12372), .ZN(n12903) );
  NAND2_X1 U11104 ( .A1(n12902), .A2(n12903), .ZN(n15047) );
  NAND2_X1 U11105 ( .A1(n10748), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n8675) );
  INV_X1 U11106 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n10746) );
  NAND2_X1 U11107 ( .A1(n10746), .A2(P2_DATAO_REG_12__SCAN_IN), .ZN(n8660) );
  OR2_X1 U11108 ( .A1(n8662), .A2(n8661), .ZN(n8663) );
  NAND2_X1 U11109 ( .A1(n8676), .A2(n8663), .ZN(n10456) );
  OR2_X1 U11110 ( .A1(n10456), .A2(n8811), .ZN(n8666) );
  NAND2_X1 U11111 ( .A1(n6697), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8664) );
  XNOR2_X1 U11112 ( .A(n8664), .B(P3_IR_REG_12__SCAN_IN), .ZN(n13048) );
  AOI22_X1 U11113 ( .A1(n12799), .A2(SI_12_), .B1(n10909), .B2(n13048), .ZN(
        n8665) );
  NAND2_X1 U11114 ( .A1(n8666), .A2(n8665), .ZN(n15069) );
  NAND2_X1 U11115 ( .A1(n8798), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n8674) );
  INV_X1 U11116 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n12375) );
  OR2_X1 U11117 ( .A1(n11986), .A2(n12375), .ZN(n8673) );
  INV_X1 U11118 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n8667) );
  OR2_X1 U11119 ( .A1(n8524), .A2(n8667), .ZN(n8672) );
  NAND2_X1 U11120 ( .A1(n8669), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n8670) );
  AND2_X1 U11121 ( .A1(n8686), .A2(n8670), .ZN(n12374) );
  OR2_X1 U11122 ( .A1(n8737), .A2(n12374), .ZN(n8671) );
  OR2_X1 U11123 ( .A1(n15069), .A2(n12180), .ZN(n12907) );
  NAND2_X1 U11124 ( .A1(n15069), .A2(n12180), .ZN(n12906) );
  INV_X1 U11125 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n10837) );
  NAND2_X1 U11126 ( .A1(n8678), .A2(n10837), .ZN(n8679) );
  NAND2_X1 U11127 ( .A1(n8692), .A2(n8679), .ZN(n10485) );
  OR2_X1 U11128 ( .A1(n8698), .A2(n8680), .ZN(n8681) );
  XNOR2_X1 U11129 ( .A(n8681), .B(n8697), .ZN(n15605) );
  INV_X1 U11130 ( .A(n15605), .ZN(n13020) );
  OAI22_X1 U11131 ( .A1(n12806), .A2(SI_13_), .B1(n13020), .B2(n6852), .ZN(
        n8682) );
  NAND2_X1 U11132 ( .A1(n8798), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n8691) );
  INV_X1 U11133 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n8683) );
  OR2_X1 U11134 ( .A1(n11986), .A2(n8683), .ZN(n8690) );
  OR2_X1 U11135 ( .A1(n8524), .A2(n15064), .ZN(n8689) );
  INV_X1 U11136 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n8684) );
  NAND2_X1 U11137 ( .A1(n8686), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n8687) );
  AND2_X1 U11138 ( .A1(n8703), .A2(n8687), .ZN(n12365) );
  OR2_X1 U11139 ( .A1(n8737), .A2(n12365), .ZN(n8688) );
  NAND4_X1 U11140 ( .A1(n8691), .A2(n8690), .A3(n8689), .A4(n8688), .ZN(n13292) );
  NAND2_X1 U11141 ( .A1(n12364), .A2(n12373), .ZN(n12912) );
  OR2_X1 U11142 ( .A1(n12364), .A2(n12373), .ZN(n12911) );
  INV_X1 U11143 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n11353) );
  NAND2_X1 U11144 ( .A1(n11353), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n8709) );
  INV_X1 U11145 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n11351) );
  NAND2_X1 U11146 ( .A1(n11351), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n8693) );
  OR2_X1 U11147 ( .A1(n8695), .A2(n8694), .ZN(n8696) );
  NAND2_X1 U11148 ( .A1(n8710), .A2(n8696), .ZN(n10494) );
  NAND2_X1 U11149 ( .A1(n10494), .A2(n12805), .ZN(n8702) );
  INV_X1 U11150 ( .A(SI_14_), .ZN(n10495) );
  NAND2_X1 U11151 ( .A1(n8698), .A2(n8697), .ZN(n8715) );
  NAND2_X1 U11152 ( .A1(n8715), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8700) );
  INV_X1 U11153 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n8699) );
  XNOR2_X1 U11154 ( .A(n8700), .B(n8699), .ZN(n15625) );
  AOI22_X1 U11155 ( .A1(n12799), .A2(n10495), .B1(n10909), .B2(n15625), .ZN(
        n8701) );
  NAND2_X1 U11156 ( .A1(n8960), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n8708) );
  INV_X1 U11157 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n13365) );
  OR2_X1 U11158 ( .A1(n8524), .A2(n13365), .ZN(n8707) );
  NAND2_X1 U11159 ( .A1(n8703), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8704) );
  AND2_X1 U11160 ( .A1(n8721), .A2(n8704), .ZN(n13298) );
  OR2_X1 U11161 ( .A1(n8737), .A2(n13298), .ZN(n8706) );
  INV_X1 U11162 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n13421) );
  OR2_X1 U11163 ( .A1(n11989), .A2(n13421), .ZN(n8705) );
  NAND4_X1 U11164 ( .A1(n8708), .A2(n8707), .A3(n8706), .A4(n8705), .ZN(n12438) );
  NAND2_X1 U11165 ( .A1(n13423), .A2(n12438), .ZN(n12917) );
  OR2_X1 U11166 ( .A1(n13423), .A2(n12438), .ZN(n12916) );
  NAND2_X1 U11167 ( .A1(n11547), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n8727) );
  NAND2_X1 U11168 ( .A1(n11549), .A2(P2_DATAO_REG_15__SCAN_IN), .ZN(n8711) );
  OR2_X1 U11169 ( .A1(n8713), .A2(n8712), .ZN(n8714) );
  NAND2_X1 U11170 ( .A1(n8728), .A2(n8714), .ZN(n10593) );
  OR2_X1 U11171 ( .A1(n10593), .A2(n8811), .ZN(n8718) );
  NAND2_X1 U11172 ( .A1(n8733), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8716) );
  XNOR2_X1 U11173 ( .A(n8716), .B(P3_IR_REG_15__SCAN_IN), .ZN(n13058) );
  AOI22_X1 U11174 ( .A1(n12799), .A2(SI_15_), .B1(n10909), .B2(n13058), .ZN(
        n8717) );
  NAND2_X1 U11175 ( .A1(n8798), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n8726) );
  INV_X1 U11176 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n13361) );
  OR2_X1 U11177 ( .A1(n8524), .A2(n13361), .ZN(n8725) );
  INV_X1 U11178 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n14969) );
  OR2_X1 U11179 ( .A1(n11986), .A2(n14969), .ZN(n8724) );
  INV_X1 U11180 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n8719) );
  NAND2_X1 U11181 ( .A1(n8721), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8722) );
  AND2_X1 U11182 ( .A1(n8738), .A2(n8722), .ZN(n13283) );
  OR2_X1 U11183 ( .A1(n8737), .A2(n13283), .ZN(n8723) );
  NAND4_X1 U11184 ( .A1(n8726), .A2(n8725), .A3(n8724), .A4(n8723), .ZN(n13291) );
  INV_X1 U11185 ( .A(n13291), .ZN(n13262) );
  OR2_X1 U11186 ( .A1(n13282), .A2(n13262), .ZN(n12920) );
  NAND2_X1 U11187 ( .A1(n13282), .A2(n13262), .ZN(n12924) );
  NAND2_X1 U11188 ( .A1(n13281), .A2(n13280), .ZN(n13279) );
  NAND2_X1 U11189 ( .A1(n11691), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n8745) );
  NAND2_X1 U11190 ( .A1(n11689), .A2(P2_DATAO_REG_16__SCAN_IN), .ZN(n8729) );
  AND2_X1 U11191 ( .A1(n8745), .A2(n8729), .ZN(n8730) );
  OR2_X1 U11192 ( .A1(n8731), .A2(n8730), .ZN(n8732) );
  NAND2_X1 U11193 ( .A1(n8746), .A2(n8732), .ZN(n10710) );
  OR2_X1 U11194 ( .A1(n10710), .A2(n8811), .ZN(n8736) );
  NAND2_X1 U11195 ( .A1(n8748), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8734) );
  XNOR2_X1 U11196 ( .A(n8734), .B(P3_IR_REG_16__SCAN_IN), .ZN(n14990) );
  AOI22_X1 U11197 ( .A1(n12799), .A2(SI_16_), .B1(n10909), .B2(n14990), .ZN(
        n8735) );
  NAND2_X1 U11198 ( .A1(n8738), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n8739) );
  NAND2_X1 U11199 ( .A1(n8755), .A2(n8739), .ZN(n13267) );
  NAND2_X1 U11200 ( .A1(n10356), .A2(n13267), .ZN(n8743) );
  INV_X1 U11201 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n13004) );
  OR2_X1 U11202 ( .A1(n11986), .A2(n13004), .ZN(n8742) );
  INV_X1 U11203 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n13357) );
  OR2_X1 U11204 ( .A1(n8524), .A2(n13357), .ZN(n8741) );
  INV_X1 U11205 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n13413) );
  OR2_X1 U11206 ( .A1(n11989), .A2(n13413), .ZN(n8740) );
  NAND4_X1 U11207 ( .A1(n8743), .A2(n8742), .A3(n8741), .A4(n8740), .ZN(n10675) );
  OR2_X1 U11208 ( .A1(n13266), .A2(n13277), .ZN(n12921) );
  NAND2_X1 U11209 ( .A1(n13266), .A2(n13277), .ZN(n12925) );
  NAND2_X1 U11210 ( .A1(n12921), .A2(n12925), .ZN(n13259) );
  INV_X1 U11211 ( .A(n13259), .ZN(n13264) );
  NAND2_X1 U11212 ( .A1(n11733), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n8764) );
  NAND2_X1 U11213 ( .A1(n11735), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n8747) );
  NAND2_X1 U11214 ( .A1(n8764), .A2(n8747), .ZN(n8761) );
  XNOR2_X1 U11215 ( .A(n8763), .B(n8761), .ZN(n10833) );
  NAND2_X1 U11216 ( .A1(n10833), .A2(n12805), .ZN(n8752) );
  OAI21_X1 U11217 ( .B1(n8748), .B2(P3_IR_REG_16__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8749) );
  MUX2_X1 U11218 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8749), .S(
        P3_IR_REG_17__SCAN_IN), .Z(n8750) );
  NAND2_X1 U11219 ( .A1(n8750), .A2(n8770), .ZN(n15016) );
  AOI22_X1 U11220 ( .A1(n12799), .A2(SI_17_), .B1(n10909), .B2(n13060), .ZN(
        n8751) );
  INV_X1 U11221 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n8753) );
  NAND2_X1 U11222 ( .A1(n8755), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n8756) );
  NAND2_X1 U11223 ( .A1(n8774), .A2(n8756), .ZN(n13252) );
  NAND2_X1 U11224 ( .A1(n10356), .A2(n13252), .ZN(n8760) );
  INV_X1 U11225 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n13353) );
  OR2_X1 U11226 ( .A1(n8524), .A2(n13353), .ZN(n8759) );
  INV_X1 U11227 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n13409) );
  OR2_X1 U11228 ( .A1(n11989), .A2(n13409), .ZN(n8758) );
  INV_X1 U11229 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n15008) );
  OR2_X1 U11230 ( .A1(n11986), .A2(n15008), .ZN(n8757) );
  NAND4_X1 U11231 ( .A1(n8760), .A2(n8759), .A3(n8758), .A4(n8757), .ZN(n13234) );
  OR2_X1 U11232 ( .A1(n13251), .A2(n13263), .ZN(n12931) );
  NAND2_X1 U11233 ( .A1(n13251), .A2(n13263), .ZN(n12933) );
  NAND2_X1 U11234 ( .A1(n12931), .A2(n12933), .ZN(n13245) );
  INV_X1 U11235 ( .A(n13245), .ZN(n13250) );
  INV_X1 U11236 ( .A(n8761), .ZN(n8762) );
  INV_X1 U11237 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n11983) );
  NAND2_X1 U11238 ( .A1(n11983), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n8780) );
  INV_X1 U11239 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n11980) );
  NAND2_X1 U11240 ( .A1(n11980), .A2(P2_DATAO_REG_18__SCAN_IN), .ZN(n8766) );
  AND2_X1 U11241 ( .A1(n8780), .A2(n8766), .ZN(n8767) );
  OR2_X1 U11242 ( .A1(n8768), .A2(n8767), .ZN(n8769) );
  NAND2_X1 U11243 ( .A1(n8781), .A2(n8769), .ZN(n10878) );
  OR2_X1 U11244 ( .A1(n10878), .A2(n8811), .ZN(n8773) );
  NAND2_X1 U11245 ( .A1(n8770), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8771) );
  XNOR2_X1 U11246 ( .A(n8771), .B(P3_IR_REG_18__SCAN_IN), .ZN(n15023) );
  AOI22_X1 U11247 ( .A1(n12799), .A2(SI_18_), .B1(n10909), .B2(n15023), .ZN(
        n8772) );
  NAND2_X1 U11248 ( .A1(n8774), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8775) );
  NAND2_X1 U11249 ( .A1(n8789), .A2(n8775), .ZN(n13237) );
  NAND2_X1 U11250 ( .A1(n13237), .A2(n10356), .ZN(n8779) );
  NAND2_X1 U11251 ( .A1(n8960), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n8778) );
  INV_X1 U11252 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n13063) );
  OR2_X1 U11253 ( .A1(n8524), .A2(n13063), .ZN(n8777) );
  NAND2_X1 U11254 ( .A1(n8798), .A2(P3_REG0_REG_18__SCAN_IN), .ZN(n8776) );
  NAND4_X1 U11255 ( .A1(n8779), .A2(n8778), .A3(n8777), .A4(n8776), .ZN(n13219) );
  NAND2_X1 U11256 ( .A1(n13240), .A2(n13248), .ZN(n12935) );
  INV_X1 U11257 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n12026) );
  NAND2_X1 U11258 ( .A1(n12026), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n8793) );
  INV_X1 U11259 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n12028) );
  NAND2_X1 U11260 ( .A1(n12028), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n8782) );
  AND2_X1 U11261 ( .A1(n8793), .A2(n8782), .ZN(n8783) );
  OR2_X1 U11262 ( .A1(n8784), .A2(n8783), .ZN(n8785) );
  NAND2_X1 U11263 ( .A1(n8794), .A2(n8785), .ZN(n11120) );
  OR2_X1 U11264 ( .A1(n11120), .A2(n8811), .ZN(n8787) );
  AOI22_X1 U11265 ( .A1(n12799), .A2(SI_19_), .B1(n7356), .B2(n10909), .ZN(
        n8786) );
  INV_X1 U11266 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n13008) );
  INV_X1 U11267 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n10192) );
  NAND2_X1 U11268 ( .A1(n8789), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8790) );
  NAND2_X1 U11269 ( .A1(n8796), .A2(n8790), .ZN(n13226) );
  NAND2_X1 U11270 ( .A1(n13226), .A2(n10356), .ZN(n8792) );
  AOI22_X1 U11271 ( .A1(n8798), .A2(P3_REG0_REG_19__SCAN_IN), .B1(n11984), 
        .B2(P3_REG1_REG_19__SCAN_IN), .ZN(n8791) );
  OAI211_X1 U11272 ( .C1(n11986), .C2(n13008), .A(n8792), .B(n8791), .ZN(
        n13235) );
  INV_X1 U11273 ( .A(n13235), .ZN(n13207) );
  NAND2_X1 U11274 ( .A1(n13225), .A2(n13207), .ZN(n12940) );
  INV_X1 U11275 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n12138) );
  XNOR2_X1 U11276 ( .A(n8803), .B(P2_DATAO_REG_20__SCAN_IN), .ZN(n11513) );
  NOR2_X1 U11277 ( .A1(n12806), .A2(n11515), .ZN(n8795) );
  INV_X1 U11278 ( .A(P3_REG2_REG_20__SCAN_IN), .ZN(n8801) );
  NAND2_X1 U11279 ( .A1(n8796), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n8797) );
  NAND2_X1 U11280 ( .A1(n8815), .A2(n8797), .ZN(n13210) );
  NAND2_X1 U11281 ( .A1(n13210), .A2(n10356), .ZN(n8800) );
  AOI22_X1 U11282 ( .A1(n8798), .A2(P3_REG0_REG_20__SCAN_IN), .B1(n11984), 
        .B2(P3_REG1_REG_20__SCAN_IN), .ZN(n8799) );
  OAI211_X1 U11283 ( .C1(n11986), .C2(n8801), .A(n8800), .B(n8799), .ZN(n13220) );
  NAND2_X1 U11284 ( .A1(n13402), .A2(n6674), .ZN(n12944) );
  OR2_X1 U11285 ( .A1(n13402), .A2(n6674), .ZN(n12945) );
  NAND2_X1 U11286 ( .A1(n12944), .A2(n12945), .ZN(n13204) );
  INV_X1 U11287 ( .A(n13204), .ZN(n8802) );
  INV_X1 U11288 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n12154) );
  NAND2_X1 U11289 ( .A1(n12154), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n8821) );
  INV_X1 U11290 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n12660) );
  NAND2_X1 U11291 ( .A1(n12660), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n8807) );
  NAND2_X1 U11292 ( .A1(n8821), .A2(n8807), .ZN(n8808) );
  NAND2_X1 U11293 ( .A1(n8809), .A2(n8808), .ZN(n8810) );
  NAND2_X1 U11294 ( .A1(n8822), .A2(n8810), .ZN(n11545) );
  INV_X1 U11295 ( .A(SI_21_), .ZN(n11544) );
  OR2_X1 U11296 ( .A1(n12806), .A2(n11544), .ZN(n8812) );
  INV_X1 U11297 ( .A(n8815), .ZN(n8814) );
  INV_X1 U11298 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n10223) );
  NAND2_X1 U11299 ( .A1(n8815), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n8816) );
  NAND2_X1 U11300 ( .A1(n8825), .A2(n8816), .ZN(n13198) );
  INV_X1 U11301 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n13396) );
  NAND2_X1 U11302 ( .A1(n11984), .A2(P3_REG1_REG_21__SCAN_IN), .ZN(n8818) );
  NAND2_X1 U11303 ( .A1(n8960), .A2(P3_REG2_REG_21__SCAN_IN), .ZN(n8817) );
  OAI211_X1 U11304 ( .C1(n11989), .C2(n13396), .A(n8818), .B(n8817), .ZN(n8819) );
  AOI21_X2 U11305 ( .B1(n13198), .B2(n10356), .A(n8819), .ZN(n13208) );
  NAND2_X1 U11306 ( .A1(n12708), .A2(n13208), .ZN(n12844) );
  NAND2_X1 U11307 ( .A1(n13197), .A2(n12844), .ZN(n8820) );
  OR2_X1 U11308 ( .A1(n12708), .A2(n13208), .ZN(n12843) );
  NAND2_X1 U11309 ( .A1(n8820), .A2(n12843), .ZN(n13180) );
  INV_X1 U11310 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n12533) );
  XNOR2_X1 U11311 ( .A(n12533), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n8833) );
  XNOR2_X1 U11312 ( .A(n8834), .B(n8833), .ZN(n11695) );
  NAND2_X1 U11313 ( .A1(n11695), .A2(n12805), .ZN(n8824) );
  OR2_X1 U11314 ( .A1(n12806), .A2(n10097), .ZN(n8823) );
  OR2_X2 U11315 ( .A1(n8825), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8839) );
  NAND2_X1 U11316 ( .A1(n8825), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8826) );
  NAND2_X1 U11317 ( .A1(n8839), .A2(n8826), .ZN(n13182) );
  NAND2_X1 U11318 ( .A1(n13182), .A2(n10356), .ZN(n8831) );
  INV_X1 U11319 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n13392) );
  NAND2_X1 U11320 ( .A1(n8960), .A2(P3_REG2_REG_22__SCAN_IN), .ZN(n8828) );
  NAND2_X1 U11321 ( .A1(n11984), .A2(P3_REG1_REG_22__SCAN_IN), .ZN(n8827) );
  OAI211_X1 U11322 ( .C1(n13392), .C2(n11989), .A(n8828), .B(n8827), .ZN(n8829) );
  INV_X1 U11323 ( .A(n8829), .ZN(n8830) );
  NAND2_X1 U11324 ( .A1(n13181), .A2(n13195), .ZN(n12955) );
  NAND2_X1 U11325 ( .A1(n13180), .A2(n12955), .ZN(n8832) );
  NAND2_X1 U11326 ( .A1(n8832), .A2(n12950), .ZN(n13165) );
  NAND2_X1 U11327 ( .A1(n12533), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n8835) );
  XNOR2_X1 U11328 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .ZN(n8846) );
  XNOR2_X1 U11329 ( .A(n8847), .B(n8846), .ZN(n11827) );
  NAND2_X1 U11330 ( .A1(n11827), .A2(n12805), .ZN(n8838) );
  OR2_X1 U11331 ( .A1(n12806), .A2(n11829), .ZN(n8837) );
  NAND2_X1 U11332 ( .A1(n8839), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8840) );
  NAND2_X1 U11333 ( .A1(n8858), .A2(n8840), .ZN(n13168) );
  NAND2_X1 U11334 ( .A1(n13168), .A2(n10356), .ZN(n8845) );
  INV_X1 U11335 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n13388) );
  NAND2_X1 U11336 ( .A1(n8960), .A2(P3_REG2_REG_23__SCAN_IN), .ZN(n8842) );
  NAND2_X1 U11337 ( .A1(n11984), .A2(P3_REG1_REG_23__SCAN_IN), .ZN(n8841) );
  OAI211_X1 U11338 ( .C1(n13388), .C2(n11989), .A(n8842), .B(n8841), .ZN(n8843) );
  INV_X1 U11339 ( .A(n8843), .ZN(n8844) );
  XNOR2_X1 U11340 ( .A(n13163), .B(n13146), .ZN(n13164) );
  INV_X1 U11341 ( .A(SI_24_), .ZN(n12064) );
  INV_X1 U11342 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n8848) );
  NAND2_X1 U11343 ( .A1(n8848), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n8849) );
  INV_X1 U11344 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n12327) );
  NAND2_X1 U11345 ( .A1(n8851), .A2(n12327), .ZN(n8852) );
  NAND2_X1 U11346 ( .A1(n8853), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n8854) );
  NAND2_X1 U11347 ( .A1(n8865), .A2(n8854), .ZN(n12063) );
  MUX2_X1 U11348 ( .A(n12064), .B(n12063), .S(n8855), .Z(n8856) );
  INV_X1 U11349 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n12753) );
  NAND2_X1 U11350 ( .A1(n8858), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n8859) );
  NAND2_X1 U11351 ( .A1(n8871), .A2(n8859), .ZN(n13151) );
  INV_X1 U11352 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n8862) );
  NAND2_X1 U11353 ( .A1(n8960), .A2(P3_REG2_REG_24__SCAN_IN), .ZN(n8861) );
  NAND2_X1 U11354 ( .A1(n11984), .A2(P3_REG1_REG_24__SCAN_IN), .ZN(n8860) );
  OAI211_X1 U11355 ( .C1(n8862), .C2(n11989), .A(n8861), .B(n8860), .ZN(n8863)
         );
  XNOR2_X1 U11356 ( .A(n13325), .B(n13160), .ZN(n13144) );
  INV_X1 U11357 ( .A(n13144), .ZN(n12951) );
  INV_X1 U11358 ( .A(n13146), .ZN(n13178) );
  OR2_X1 U11359 ( .A1(n13163), .A2(n13178), .ZN(n13139) );
  NAND2_X1 U11360 ( .A1(n13167), .A2(n12960), .ZN(n13141) );
  XNOR2_X1 U11361 ( .A(n12384), .B(P2_DATAO_REG_25__SCAN_IN), .ZN(n8866) );
  XNOR2_X1 U11362 ( .A(n8879), .B(n8866), .ZN(n12214) );
  NAND2_X1 U11363 ( .A1(n12214), .A2(n12805), .ZN(n8868) );
  OR2_X1 U11364 ( .A1(n12806), .A2(n12216), .ZN(n8867) );
  INV_X1 U11365 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n8869) );
  NAND2_X1 U11366 ( .A1(n8871), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n8872) );
  NAND2_X1 U11367 ( .A1(n8885), .A2(n8872), .ZN(n13130) );
  NAND2_X1 U11368 ( .A1(n13130), .A2(n10356), .ZN(n8877) );
  INV_X1 U11369 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n13383) );
  NAND2_X1 U11370 ( .A1(n8960), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n8874) );
  NAND2_X1 U11371 ( .A1(n11984), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n8873) );
  OAI211_X1 U11372 ( .C1(n13383), .C2(n11989), .A(n8874), .B(n8873), .ZN(n8875) );
  INV_X1 U11373 ( .A(n8875), .ZN(n8876) );
  OR2_X1 U11374 ( .A1(n13134), .A2(n13149), .ZN(n12964) );
  NAND2_X1 U11375 ( .A1(n13134), .A2(n13149), .ZN(n12965) );
  NAND2_X1 U11376 ( .A1(n12384), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n8878) );
  NAND2_X1 U11377 ( .A1(n12381), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n8880) );
  XNOR2_X1 U11378 ( .A(n8894), .B(P2_DATAO_REG_26__SCAN_IN), .ZN(n8882) );
  XNOR2_X1 U11379 ( .A(n8893), .B(n8882), .ZN(n12288) );
  NAND2_X1 U11380 ( .A1(n12288), .A2(n12805), .ZN(n8884) );
  OR2_X1 U11381 ( .A1(n12806), .A2(n12290), .ZN(n8883) );
  NAND2_X1 U11382 ( .A1(n8885), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8886) );
  NAND2_X1 U11383 ( .A1(n8902), .A2(n8886), .ZN(n13117) );
  NAND2_X1 U11384 ( .A1(n13117), .A2(n10356), .ZN(n8891) );
  INV_X1 U11385 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n13379) );
  NAND2_X1 U11386 ( .A1(n11984), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n8888) );
  NAND2_X1 U11387 ( .A1(n8960), .A2(P3_REG2_REG_26__SCAN_IN), .ZN(n8887) );
  OAI211_X1 U11388 ( .C1(n11989), .C2(n13379), .A(n8888), .B(n8887), .ZN(n8889) );
  INV_X1 U11389 ( .A(n8889), .ZN(n8890) );
  AND2_X1 U11390 ( .A1(n14890), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n8892) );
  NAND2_X1 U11391 ( .A1(n8894), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n8895) );
  XNOR2_X1 U11392 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(P2_DATAO_REG_27__SCAN_IN), 
        .ZN(n8897) );
  XNOR2_X1 U11393 ( .A(n10343), .B(n8897), .ZN(n12340) );
  NAND2_X1 U11394 ( .A1(n12340), .A2(n12805), .ZN(n8899) );
  INV_X1 U11395 ( .A(SI_27_), .ZN(n12341) );
  OR2_X1 U11396 ( .A1(n8623), .A2(n12341), .ZN(n8898) );
  INV_X1 U11397 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n8900) );
  NAND2_X1 U11398 ( .A1(n8902), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n8903) );
  NAND2_X1 U11399 ( .A1(n8958), .A2(n8903), .ZN(n13102) );
  NAND2_X1 U11400 ( .A1(n13102), .A2(n10356), .ZN(n8908) );
  NAND2_X1 U11401 ( .A1(n11984), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n8905) );
  NAND2_X1 U11402 ( .A1(n8960), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n8904) );
  OAI211_X1 U11403 ( .C1(n11989), .C2(n9009), .A(n8905), .B(n8904), .ZN(n8906)
         );
  INV_X1 U11404 ( .A(n8906), .ZN(n8907) );
  NAND2_X2 U11405 ( .A1(n8908), .A2(n8907), .ZN(n13112) );
  NAND2_X1 U11406 ( .A1(n10362), .A2(n13091), .ZN(n13083) );
  OAI21_X2 U11407 ( .B1(n10362), .B2(n13091), .A(n13083), .ZN(n12842) );
  INV_X1 U11408 ( .A(n8969), .ZN(n13106) );
  OAI21_X1 U11409 ( .B1(n11693), .B2(n9015), .A(n7356), .ZN(n8913) );
  INV_X1 U11410 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n8911) );
  NAND2_X1 U11411 ( .A1(n8913), .A2(n11681), .ZN(n8915) );
  OAI21_X1 U11412 ( .B1(n9015), .B2(n12848), .A(n11693), .ZN(n8914) );
  NAND2_X1 U11413 ( .A1(n8915), .A2(n8914), .ZN(n9883) );
  NAND2_X1 U11414 ( .A1(n9883), .A2(n15730), .ZN(n10898) );
  NAND2_X1 U11415 ( .A1(n11514), .A2(n13037), .ZN(n12982) );
  OR2_X1 U11416 ( .A1(n10898), .A2(n12982), .ZN(n8917) );
  AND2_X1 U11417 ( .A1(n9015), .A2(n13037), .ZN(n8916) );
  NAND2_X1 U11418 ( .A1(n12990), .A2(n8916), .ZN(n9018) );
  NAND2_X1 U11419 ( .A1(n8917), .A2(n9018), .ZN(n15680) );
  INV_X1 U11420 ( .A(n15680), .ZN(n15707) );
  INV_X1 U11421 ( .A(n13134), .ZN(n13385) );
  INV_X1 U11422 ( .A(n15695), .ZN(n9796) );
  NOR2_X1 U11423 ( .A1(n15682), .A2(n9796), .ZN(n9793) );
  INV_X1 U11424 ( .A(n9793), .ZN(n8919) );
  INV_X1 U11425 ( .A(n11368), .ZN(n10902) );
  NAND2_X1 U11426 ( .A1(n15699), .A2(n10902), .ZN(n15701) );
  NAND2_X1 U11427 ( .A1(n15702), .A2(n15701), .ZN(n8918) );
  NAND2_X1 U11428 ( .A1(n8919), .A2(n8918), .ZN(n15677) );
  INV_X1 U11429 ( .A(n15687), .ZN(n8920) );
  NOR2_X1 U11430 ( .A1(n15698), .A2(n8920), .ZN(n8921) );
  NAND2_X1 U11431 ( .A1(n11374), .A2(n11373), .ZN(n11372) );
  NAND2_X1 U11432 ( .A1(n15681), .A2(n12021), .ZN(n8922) );
  NAND2_X1 U11433 ( .A1(n11372), .A2(n8922), .ZN(n11564) );
  NAND2_X1 U11434 ( .A1(n11564), .A2(n11563), .ZN(n11562) );
  INV_X1 U11435 ( .A(n11569), .ZN(n15672) );
  NAND2_X1 U11436 ( .A1(n11673), .A2(n15672), .ZN(n8923) );
  NAND2_X1 U11437 ( .A1(n11562), .A2(n8923), .ZN(n11674) );
  OR2_X2 U11438 ( .A1(n11674), .A2(n6678), .ZN(n11676) );
  INV_X1 U11439 ( .A(n12995), .ZN(n11790) );
  NAND2_X1 U11440 ( .A1(n11790), .A2(n11682), .ZN(n8924) );
  NAND2_X1 U11441 ( .A1(n11947), .A2(n15664), .ZN(n8925) );
  NAND2_X1 U11442 ( .A1(n11946), .A2(n12819), .ZN(n11945) );
  INV_X1 U11443 ( .A(n11953), .ZN(n15657) );
  NAND2_X1 U11444 ( .A1(n12031), .A2(n15657), .ZN(n8926) );
  NAND2_X1 U11445 ( .A1(n12894), .A2(n12893), .ZN(n12891) );
  INV_X1 U11446 ( .A(n15731), .ZN(n12195) );
  NAND2_X1 U11447 ( .A1(n15638), .A2(n15645), .ZN(n8929) );
  INV_X1 U11448 ( .A(n15647), .ZN(n8927) );
  NAND2_X1 U11449 ( .A1(n15043), .A2(n8927), .ZN(n8928) );
  INV_X1 U11450 ( .A(n12828), .ZN(n8930) );
  NAND2_X1 U11451 ( .A1(n15069), .A2(n15042), .ZN(n8932) );
  NAND2_X1 U11452 ( .A1(n12911), .A2(n12912), .ZN(n12362) );
  NAND2_X1 U11453 ( .A1(n12364), .A2(n13292), .ZN(n8934) );
  NAND2_X1 U11454 ( .A1(n12916), .A2(n12917), .ZN(n13295) );
  INV_X1 U11455 ( .A(n12438), .ZN(n13275) );
  OR2_X1 U11456 ( .A1(n13423), .A2(n13275), .ZN(n8935) );
  NAND2_X1 U11457 ( .A1(n13289), .A2(n8935), .ZN(n13273) );
  OR2_X1 U11458 ( .A1(n13282), .A2(n13291), .ZN(n8936) );
  NAND2_X1 U11459 ( .A1(n13273), .A2(n8936), .ZN(n13258) );
  NAND2_X1 U11460 ( .A1(n13282), .A2(n13291), .ZN(n13257) );
  NAND2_X1 U11461 ( .A1(n13266), .A2(n10675), .ZN(n8937) );
  AND2_X1 U11462 ( .A1(n13257), .A2(n8937), .ZN(n8939) );
  INV_X1 U11463 ( .A(n8937), .ZN(n8938) );
  NAND2_X1 U11464 ( .A1(n13246), .A2(n13245), .ZN(n8941) );
  NAND2_X1 U11465 ( .A1(n13251), .A2(n13234), .ZN(n8940) );
  NAND2_X1 U11466 ( .A1(n8941), .A2(n8940), .ZN(n13231) );
  OR2_X1 U11467 ( .A1(n13240), .A2(n13219), .ZN(n8942) );
  NAND2_X1 U11468 ( .A1(n13181), .A2(n13159), .ZN(n8949) );
  INV_X1 U11469 ( .A(n8949), .ZN(n8945) );
  INV_X1 U11470 ( .A(n13208), .ZN(n12771) );
  OR2_X1 U11471 ( .A1(n12708), .A2(n12771), .ZN(n8944) );
  OR2_X1 U11472 ( .A1(n13402), .A2(n6673), .ZN(n8948) );
  INV_X1 U11473 ( .A(n8948), .ZN(n8943) );
  OR2_X1 U11474 ( .A1(n8943), .A2(n13204), .ZN(n13188) );
  OR2_X1 U11475 ( .A1(n13224), .A2(n8950), .ZN(n8946) );
  OR2_X1 U11476 ( .A1(n8946), .A2(n6712), .ZN(n8947) );
  NAND2_X1 U11477 ( .A1(n13225), .A2(n13235), .ZN(n13203) );
  AND2_X1 U11478 ( .A1(n13203), .A2(n8948), .ZN(n13187) );
  OR2_X1 U11479 ( .A1(n6712), .A2(n8951), .ZN(n8952) );
  NAND2_X1 U11480 ( .A1(n13163), .A2(n13146), .ZN(n8953) );
  NAND2_X1 U11481 ( .A1(n13145), .A2(n13144), .ZN(n13143) );
  OR2_X1 U11482 ( .A1(n13325), .A2(n12726), .ZN(n8954) );
  NAND2_X1 U11483 ( .A1(n13143), .A2(n8954), .ZN(n13125) );
  NAND2_X1 U11484 ( .A1(n13381), .A2(n9893), .ZN(n8955) );
  OAI21_X1 U11485 ( .B1(n8956), .B2(n12842), .A(n10361), .ZN(n8957) );
  NOR2_X1 U11486 ( .A1(n11681), .A2(n11514), .ZN(n12985) );
  NOR2_X2 U11487 ( .A1(n9004), .A2(n12985), .ZN(n15685) );
  NAND2_X1 U11488 ( .A1(n8958), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n8959) );
  NAND2_X1 U11489 ( .A1(n10355), .A2(n8959), .ZN(n13096) );
  NAND2_X1 U11490 ( .A1(n13096), .A2(n10356), .ZN(n8965) );
  INV_X1 U11491 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n13375) );
  NAND2_X1 U11492 ( .A1(n8960), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n8962) );
  NAND2_X1 U11493 ( .A1(n11984), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n8961) );
  OAI211_X1 U11494 ( .C1(n13375), .C2(n11989), .A(n8962), .B(n8961), .ZN(n8963) );
  INV_X1 U11495 ( .A(n8963), .ZN(n8964) );
  NAND2_X2 U11496 ( .A1(n8965), .A2(n8964), .ZN(n11923) );
  INV_X1 U11497 ( .A(n12667), .ZN(n12987) );
  INV_X1 U11498 ( .A(n13029), .ZN(n13039) );
  NAND2_X1 U11499 ( .A1(n12987), .A2(n13039), .ZN(n10916) );
  AND2_X1 U11500 ( .A1(n6852), .A2(n10916), .ZN(n8967) );
  INV_X1 U11501 ( .A(n8967), .ZN(n8966) );
  AOI22_X1 U11502 ( .A1(n11923), .A2(n15697), .B1(n15700), .B2(n13127), .ZN(
        n8968) );
  INV_X1 U11503 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n8971) );
  INV_X1 U11504 ( .A(n8973), .ZN(n8974) );
  NAND2_X1 U11505 ( .A1(n8974), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8975) );
  MUX2_X1 U11506 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8975), .S(
        P3_IR_REG_25__SCAN_IN), .Z(n8977) );
  NAND2_X1 U11507 ( .A1(n8977), .A2(n8976), .ZN(n12217) );
  INV_X1 U11508 ( .A(n12217), .ZN(n8981) );
  NAND2_X1 U11509 ( .A1(n8976), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8978) );
  XNOR2_X1 U11510 ( .A(n8978), .B(P3_IR_REG_26__SCAN_IN), .ZN(n8986) );
  NAND2_X1 U11511 ( .A1(n6769), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8979) );
  XNOR2_X1 U11512 ( .A(n8979), .B(n8447), .ZN(n12065) );
  INV_X1 U11513 ( .A(n12065), .ZN(n8980) );
  NAND3_X1 U11514 ( .A1(n8981), .A2(n8986), .A3(n8980), .ZN(n10408) );
  INV_X1 U11515 ( .A(n10907), .ZN(n8982) );
  NOR2_X1 U11516 ( .A1(n8982), .A2(n12982), .ZN(n9879) );
  XNOR2_X1 U11517 ( .A(n12065), .B(P3_B_REG_SCAN_IN), .ZN(n8983) );
  NAND2_X1 U11518 ( .A1(n12217), .A2(n8983), .ZN(n8984) );
  INV_X1 U11519 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n8985) );
  NAND2_X1 U11520 ( .A1(n10623), .A2(n8985), .ZN(n8988) );
  INV_X1 U11521 ( .A(n8986), .ZN(n12291) );
  NAND2_X1 U11522 ( .A1(n12291), .A2(n12217), .ZN(n8987) );
  INV_X1 U11523 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n8989) );
  NAND2_X1 U11524 ( .A1(n10623), .A2(n8989), .ZN(n8991) );
  NAND2_X1 U11525 ( .A1(n12291), .A2(n12065), .ZN(n8990) );
  NAND2_X1 U11526 ( .A1(n8991), .A2(n8990), .ZN(n9789) );
  INV_X1 U11527 ( .A(n9789), .ZN(n13427) );
  AND2_X1 U11528 ( .A1(n13425), .A2(n13427), .ZN(n9013) );
  NOR2_X1 U11529 ( .A1(P3_D_REG_17__SCAN_IN), .A2(P3_D_REG_22__SCAN_IN), .ZN(
        n8995) );
  NOR4_X1 U11530 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        P3_D_REG_25__SCAN_IN), .A4(P3_D_REG_20__SCAN_IN), .ZN(n8994) );
  NOR4_X1 U11531 ( .A1(P3_D_REG_29__SCAN_IN), .A2(P3_D_REG_10__SCAN_IN), .A3(
        P3_D_REG_31__SCAN_IN), .A4(P3_D_REG_14__SCAN_IN), .ZN(n8993) );
  NOR4_X1 U11532 ( .A1(P3_D_REG_19__SCAN_IN), .A2(P3_D_REG_18__SCAN_IN), .A3(
        P3_D_REG_27__SCAN_IN), .A4(P3_D_REG_24__SCAN_IN), .ZN(n8992) );
  NAND4_X1 U11533 ( .A1(n8995), .A2(n8994), .A3(n8993), .A4(n8992), .ZN(n9001)
         );
  NOR4_X1 U11534 ( .A1(P3_D_REG_9__SCAN_IN), .A2(P3_D_REG_16__SCAN_IN), .A3(
        P3_D_REG_15__SCAN_IN), .A4(P3_D_REG_30__SCAN_IN), .ZN(n8999) );
  NOR4_X1 U11535 ( .A1(P3_D_REG_11__SCAN_IN), .A2(P3_D_REG_21__SCAN_IN), .A3(
        P3_D_REG_12__SCAN_IN), .A4(P3_D_REG_26__SCAN_IN), .ZN(n8998) );
  NOR4_X1 U11536 ( .A1(P3_D_REG_3__SCAN_IN), .A2(P3_D_REG_5__SCAN_IN), .A3(
        P3_D_REG_4__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n8997) );
  NOR4_X1 U11537 ( .A1(P3_D_REG_13__SCAN_IN), .A2(P3_D_REG_28__SCAN_IN), .A3(
        P3_D_REG_23__SCAN_IN), .A4(P3_D_REG_6__SCAN_IN), .ZN(n8996) );
  NAND4_X1 U11538 ( .A1(n8999), .A2(n8998), .A3(n8997), .A4(n8996), .ZN(n9000)
         );
  OAI21_X1 U11539 ( .B1(n9001), .B2(n9000), .A(n10623), .ZN(n9010) );
  NAND2_X1 U11540 ( .A1(n9013), .A2(n9010), .ZN(n9882) );
  INV_X1 U11541 ( .A(n9882), .ZN(n9002) );
  NAND2_X1 U11542 ( .A1(n9881), .A2(n9002), .ZN(n9008) );
  NAND2_X1 U11543 ( .A1(n11681), .A2(n9015), .ZN(n12983) );
  INV_X1 U11544 ( .A(n12983), .ZN(n9003) );
  NAND2_X1 U11545 ( .A1(n9004), .A2(n9003), .ZN(n9887) );
  AND2_X1 U11546 ( .A1(n9789), .A2(n11360), .ZN(n9012) );
  NAND2_X1 U11547 ( .A1(n9012), .A2(n9010), .ZN(n9880) );
  INV_X1 U11548 ( .A(n9880), .ZN(n9888) );
  NAND2_X1 U11549 ( .A1(n9883), .A2(n9888), .ZN(n9005) );
  OAI21_X1 U11550 ( .B1(n9887), .B2(n9882), .A(n9005), .ZN(n9006) );
  NAND2_X1 U11551 ( .A1(n9006), .A2(n10907), .ZN(n9007) );
  INV_X1 U11552 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n9022) );
  INV_X1 U11553 ( .A(n9010), .ZN(n9011) );
  NOR3_X1 U11554 ( .A1(n9013), .A2(n9012), .A3(n9011), .ZN(n9014) );
  AND2_X1 U11555 ( .A1(n10907), .A2(n9014), .ZN(n11359) );
  OAI22_X1 U11556 ( .A1(n15730), .A2(n9015), .B1(n7356), .B2(n11693), .ZN(
        n9016) );
  AOI21_X1 U11557 ( .B1(n9016), .B2(n12982), .A(n12963), .ZN(n9017) );
  NAND2_X1 U11558 ( .A1(n12975), .A2(n9018), .ZN(n11356) );
  NAND2_X1 U11559 ( .A1(n12963), .A2(n12982), .ZN(n9884) );
  NAND2_X1 U11560 ( .A1(n11356), .A2(n9884), .ZN(n11357) );
  NAND2_X1 U11561 ( .A1(n11357), .A2(n13425), .ZN(n9019) );
  MUX2_X1 U11562 ( .A(n9022), .B(n9021), .S(n15751), .Z(n9024) );
  NAND2_X1 U11563 ( .A1(n10362), .A2(n10382), .ZN(n9023) );
  NAND2_X1 U11564 ( .A1(n9024), .A2(n9023), .ZN(P3_U3486) );
  NAND2_X1 U11565 ( .A1(n9291), .A2(n11045), .ZN(n9026) );
  AOI21_X1 U11566 ( .B1(n9027), .B2(n12137), .A(n9026), .ZN(n9028) );
  INV_X1 U11567 ( .A(n9028), .ZN(n9237) );
  NAND2_X1 U11568 ( .A1(n11125), .A2(n6669), .ZN(n9030) );
  OAI21_X1 U11569 ( .B1(n11125), .B2(n9237), .A(n9030), .ZN(n9033) );
  NAND2_X1 U11570 ( .A1(n9031), .A2(n9029), .ZN(n9032) );
  NAND2_X1 U11571 ( .A1(n9033), .A2(n9032), .ZN(n9038) );
  NAND2_X1 U11572 ( .A1(n9049), .A2(n13932), .ZN(n9035) );
  NAND2_X1 U11573 ( .A1(n9239), .A2(n13658), .ZN(n9034) );
  NAND2_X1 U11574 ( .A1(n9038), .A2(n9037), .ZN(n9044) );
  NAND2_X1 U11575 ( .A1(n9239), .A2(n13656), .ZN(n9040) );
  NAND2_X1 U11576 ( .A1(n9040), .A2(n9039), .ZN(n9047) );
  NAND2_X1 U11577 ( .A1(n9047), .A2(n9046), .ZN(n9043) );
  NAND3_X1 U11578 ( .A1(n9045), .A2(n9044), .A3(n9043), .ZN(n9048) );
  NAND2_X1 U11579 ( .A1(n9048), .A2(n6739), .ZN(n9055) );
  INV_X1 U11580 ( .A(n9049), .ZN(n9129) );
  NAND2_X1 U11581 ( .A1(n13515), .A2(n9129), .ZN(n9051) );
  NAND2_X1 U11582 ( .A1(n13655), .A2(n9226), .ZN(n9050) );
  NAND2_X1 U11583 ( .A1(n9051), .A2(n9050), .ZN(n9054) );
  AOI22_X1 U11584 ( .A1(n13515), .A2(n9226), .B1(n9239), .B2(n13655), .ZN(
        n9052) );
  AOI21_X1 U11585 ( .B1(n9055), .B2(n9054), .A(n9052), .ZN(n9053) );
  INV_X1 U11586 ( .A(n9053), .ZN(n9056) );
  NAND2_X1 U11587 ( .A1(n9056), .A2(n7693), .ZN(n9061) );
  NAND2_X1 U11588 ( .A1(n11400), .A2(n9226), .ZN(n9058) );
  NAND2_X1 U11589 ( .A1(n9129), .A2(n13654), .ZN(n9057) );
  NAND2_X1 U11590 ( .A1(n9058), .A2(n9057), .ZN(n9060) );
  AOI22_X1 U11591 ( .A1(n11400), .A2(n9239), .B1(n9226), .B2(n13654), .ZN(
        n9059) );
  NAND2_X1 U11592 ( .A1(n11523), .A2(n6669), .ZN(n9063) );
  NAND2_X1 U11593 ( .A1(n13653), .A2(n9226), .ZN(n9062) );
  NAND2_X1 U11594 ( .A1(n9063), .A2(n9062), .ZN(n9068) );
  NAND2_X1 U11595 ( .A1(n11523), .A2(n9226), .ZN(n9064) );
  OAI21_X1 U11596 ( .B1(n11089), .B2(n9226), .A(n9064), .ZN(n9065) );
  NAND2_X1 U11597 ( .A1(n9066), .A2(n9065), .ZN(n9072) );
  INV_X1 U11598 ( .A(n9067), .ZN(n9070) );
  INV_X1 U11599 ( .A(n9068), .ZN(n9069) );
  NAND2_X1 U11600 ( .A1(n9070), .A2(n9069), .ZN(n9071) );
  NAND2_X1 U11601 ( .A1(n11429), .A2(n9226), .ZN(n9074) );
  NAND2_X1 U11602 ( .A1(n9129), .A2(n13652), .ZN(n9073) );
  NAND2_X1 U11603 ( .A1(n9074), .A2(n9073), .ZN(n9076) );
  NAND2_X1 U11604 ( .A1(n11594), .A2(n9129), .ZN(n9078) );
  NAND2_X1 U11605 ( .A1(n13651), .A2(n9226), .ZN(n9077) );
  AOI22_X1 U11606 ( .A1(n11594), .A2(n9226), .B1(n13651), .B2(n9239), .ZN(
        n9079) );
  NAND2_X1 U11607 ( .A1(n11662), .A2(n9226), .ZN(n9081) );
  NAND2_X1 U11608 ( .A1(n9129), .A2(n13650), .ZN(n9080) );
  NAND2_X1 U11609 ( .A1(n9081), .A2(n9080), .ZN(n9083) );
  AOI22_X1 U11610 ( .A1(n11662), .A2(n6669), .B1(n9241), .B2(n13650), .ZN(
        n9082) );
  NAND2_X1 U11611 ( .A1(n11755), .A2(n9129), .ZN(n9085) );
  NAND2_X1 U11612 ( .A1(n13649), .A2(n9226), .ZN(n9084) );
  NAND2_X1 U11613 ( .A1(n11755), .A2(n9226), .ZN(n9087) );
  OAI21_X1 U11614 ( .B1(n9088), .B2(n9226), .A(n9087), .ZN(n9089) );
  NAND2_X1 U11615 ( .A1(n15507), .A2(n9226), .ZN(n9092) );
  NAND2_X1 U11616 ( .A1(n9129), .A2(n13648), .ZN(n9091) );
  NAND2_X1 U11617 ( .A1(n15507), .A2(n9129), .ZN(n9093) );
  OAI21_X1 U11618 ( .B1(n9094), .B2(n9239), .A(n9093), .ZN(n9095) );
  NAND2_X1 U11619 ( .A1(n9096), .A2(n9095), .ZN(n9100) );
  INV_X1 U11620 ( .A(n9097), .ZN(n9098) );
  NAND2_X1 U11621 ( .A1(n9098), .A2(n6751), .ZN(n9099) );
  NAND2_X1 U11622 ( .A1(n9100), .A2(n9099), .ZN(n9105) );
  NAND2_X1 U11623 ( .A1(n12068), .A2(n9129), .ZN(n9102) );
  NAND2_X1 U11624 ( .A1(n13647), .A2(n9226), .ZN(n9101) );
  NAND2_X1 U11625 ( .A1(n9102), .A2(n9101), .ZN(n9104) );
  AOI22_X1 U11626 ( .A1(n12068), .A2(n9226), .B1(n13647), .B2(n6669), .ZN(
        n9103) );
  AOI21_X1 U11627 ( .B1(n9105), .B2(n9104), .A(n9103), .ZN(n9107) );
  NOR2_X1 U11628 ( .A1(n9105), .A2(n9104), .ZN(n9106) );
  NAND2_X1 U11629 ( .A1(n14019), .A2(n9226), .ZN(n9109) );
  NAND2_X1 U11630 ( .A1(n9239), .A2(n13646), .ZN(n9108) );
  NAND2_X1 U11631 ( .A1(n9109), .A2(n9108), .ZN(n9110) );
  NAND2_X1 U11632 ( .A1(n9111), .A2(n9110), .ZN(n9114) );
  NAND2_X1 U11633 ( .A1(n14019), .A2(n9129), .ZN(n9112) );
  OAI21_X1 U11634 ( .B1(n9269), .B2(n9239), .A(n9112), .ZN(n9113) );
  NAND2_X1 U11635 ( .A1(n9114), .A2(n9113), .ZN(n9115) );
  NAND2_X1 U11636 ( .A1(n12090), .A2(n9129), .ZN(n9118) );
  NAND2_X1 U11637 ( .A1(n13645), .A2(n9241), .ZN(n9117) );
  AOI22_X1 U11638 ( .A1(n12090), .A2(n9226), .B1(n13645), .B2(n9239), .ZN(
        n9119) );
  NAND2_X1 U11639 ( .A1(n12277), .A2(n9241), .ZN(n9122) );
  NAND2_X1 U11640 ( .A1(n9129), .A2(n13644), .ZN(n9121) );
  NAND2_X1 U11641 ( .A1(n12277), .A2(n9129), .ZN(n9124) );
  NAND2_X1 U11642 ( .A1(n13644), .A2(n9241), .ZN(n9123) );
  NAND2_X1 U11643 ( .A1(n9124), .A2(n9123), .ZN(n9125) );
  AND2_X1 U11644 ( .A1(n13643), .A2(n9239), .ZN(n9128) );
  AOI21_X1 U11645 ( .B1(n12310), .B2(n9241), .A(n9128), .ZN(n9141) );
  NAND2_X1 U11646 ( .A1(n12310), .A2(n9129), .ZN(n9131) );
  NAND2_X1 U11647 ( .A1(n13643), .A2(n9241), .ZN(n9130) );
  NAND2_X1 U11648 ( .A1(n9131), .A2(n9130), .ZN(n9140) );
  AND2_X1 U11649 ( .A1(n13641), .A2(n9241), .ZN(n9132) );
  AOI21_X1 U11650 ( .B1(n13443), .B2(n9129), .A(n9132), .ZN(n9149) );
  NAND2_X1 U11651 ( .A1(n13443), .A2(n9241), .ZN(n9134) );
  NAND2_X1 U11652 ( .A1(n13641), .A2(n6669), .ZN(n9133) );
  NAND2_X1 U11653 ( .A1(n9134), .A2(n9133), .ZN(n9147) );
  AND2_X1 U11654 ( .A1(n13642), .A2(n9241), .ZN(n9135) );
  AOI21_X1 U11655 ( .B1(n12475), .B2(n9129), .A(n9135), .ZN(n9143) );
  NAND2_X1 U11656 ( .A1(n12475), .A2(n9226), .ZN(n9137) );
  NAND2_X1 U11657 ( .A1(n13642), .A2(n9239), .ZN(n9136) );
  NAND2_X1 U11658 ( .A1(n9137), .A2(n9136), .ZN(n9142) );
  AOI22_X1 U11659 ( .A1(n9149), .A2(n9147), .B1(n9143), .B2(n9142), .ZN(n9139)
         );
  INV_X1 U11660 ( .A(n9139), .ZN(n9156) );
  NAND2_X1 U11661 ( .A1(n9141), .A2(n9140), .ZN(n9155) );
  INV_X1 U11662 ( .A(n9142), .ZN(n9145) );
  INV_X1 U11663 ( .A(n9143), .ZN(n9144) );
  NAND2_X1 U11664 ( .A1(n9145), .A2(n9144), .ZN(n9148) );
  INV_X1 U11665 ( .A(n13443), .ZN(n14058) );
  NAND3_X1 U11666 ( .A1(n9148), .A2(n9146), .A3(n14058), .ZN(n9153) );
  INV_X1 U11667 ( .A(n9147), .ZN(n9152) );
  INV_X1 U11668 ( .A(n9148), .ZN(n9151) );
  INV_X1 U11669 ( .A(n9149), .ZN(n9150) );
  AOI22_X1 U11670 ( .A1(n9153), .A2(n9152), .B1(n9151), .B2(n9150), .ZN(n9154)
         );
  OAI21_X1 U11671 ( .B1(n9156), .B2(n9155), .A(n9154), .ZN(n9157) );
  AND2_X1 U11672 ( .A1(n13640), .A2(n9239), .ZN(n9158) );
  AOI21_X1 U11673 ( .B1(n14053), .B2(n9241), .A(n9158), .ZN(n9162) );
  NAND2_X1 U11674 ( .A1(n14053), .A2(n9239), .ZN(n9159) );
  OAI21_X1 U11675 ( .B1(n9160), .B2(n9129), .A(n9159), .ZN(n9161) );
  NAND2_X1 U11676 ( .A1(n9163), .A2(n9162), .ZN(n9164) );
  NAND2_X1 U11677 ( .A1(n9165), .A2(n9164), .ZN(n9171) );
  NAND2_X1 U11678 ( .A1(n13893), .A2(n6669), .ZN(n9167) );
  NAND2_X1 U11679 ( .A1(n13639), .A2(n9241), .ZN(n9166) );
  NAND2_X1 U11680 ( .A1(n9167), .A2(n9166), .ZN(n9170) );
  AOI22_X1 U11681 ( .A1(n13893), .A2(n9226), .B1(n13639), .B2(n9239), .ZN(
        n9168) );
  NAND2_X1 U11682 ( .A1(n13986), .A2(n9241), .ZN(n9173) );
  NAND2_X1 U11683 ( .A1(n13638), .A2(n6669), .ZN(n9172) );
  NAND2_X1 U11684 ( .A1(n9173), .A2(n9172), .ZN(n9175) );
  AOI22_X1 U11685 ( .A1(n13986), .A2(n9129), .B1(n9241), .B2(n13638), .ZN(
        n9174) );
  NAND2_X1 U11686 ( .A1(n13859), .A2(n6669), .ZN(n9177) );
  NAND2_X1 U11687 ( .A1(n13637), .A2(n9241), .ZN(n9176) );
  NAND2_X1 U11688 ( .A1(n13859), .A2(n9241), .ZN(n9178) );
  OAI21_X1 U11689 ( .B1(n13579), .B2(n9049), .A(n9178), .ZN(n9179) );
  NAND2_X1 U11690 ( .A1(n13975), .A2(n9241), .ZN(n9181) );
  NAND2_X1 U11691 ( .A1(n13636), .A2(n9239), .ZN(n9180) );
  NAND2_X1 U11692 ( .A1(n9181), .A2(n9180), .ZN(n9183) );
  AOI22_X1 U11693 ( .A1(n13975), .A2(n6669), .B1(n9241), .B2(n13636), .ZN(
        n9182) );
  NAND2_X1 U11694 ( .A1(n13970), .A2(n6669), .ZN(n9185) );
  NAND2_X1 U11695 ( .A1(n13635), .A2(n9241), .ZN(n9184) );
  NAND2_X1 U11696 ( .A1(n9185), .A2(n9184), .ZN(n9187) );
  AOI22_X1 U11697 ( .A1(n13970), .A2(n9226), .B1(n13635), .B2(n9086), .ZN(
        n9186) );
  AOI21_X1 U11698 ( .B1(n9188), .B2(n9187), .A(n9186), .ZN(n9190) );
  NOR2_X1 U11699 ( .A1(n9188), .A2(n9187), .ZN(n9189) );
  AOI22_X1 U11700 ( .A1(n13965), .A2(n9226), .B1(n13634), .B2(n6669), .ZN(
        n9191) );
  AOI22_X1 U11701 ( .A1(n13965), .A2(n6669), .B1(n9241), .B2(n13634), .ZN(
        n9193) );
  INV_X1 U11702 ( .A(n9196), .ZN(n9198) );
  OAI22_X1 U11703 ( .A1(n14041), .A2(n9241), .B1(n13486), .B2(n6669), .ZN(
        n9195) );
  INV_X1 U11704 ( .A(n9195), .ZN(n9197) );
  AOI22_X1 U11705 ( .A1(n13797), .A2(n9241), .B1(n13633), .B2(n6669), .ZN(
        n9194) );
  AOI22_X1 U11706 ( .A1(n13778), .A2(n9226), .B1(n13632), .B2(n6669), .ZN(
        n9199) );
  NOR2_X1 U11707 ( .A1(n9200), .A2(n9199), .ZN(n9204) );
  AOI22_X1 U11708 ( .A1(n13778), .A2(n6669), .B1(n9241), .B2(n13632), .ZN(
        n9203) );
  INV_X1 U11709 ( .A(n9199), .ZN(n9202) );
  INV_X1 U11710 ( .A(n9200), .ZN(n9201) );
  OAI22_X1 U11711 ( .A1(n9204), .A2(n9203), .B1(n9202), .B2(n9201), .ZN(n9207)
         );
  OAI22_X1 U11712 ( .A1(n13766), .A2(n9049), .B1(n13616), .B2(n6669), .ZN(
        n9206) );
  AOI22_X1 U11713 ( .A1(n13541), .A2(n9226), .B1(n8388), .B2(n6669), .ZN(n9228) );
  OAI22_X1 U11714 ( .A1(n14032), .A2(n9241), .B1(n13536), .B2(n6669), .ZN(
        n9227) );
  AOI22_X1 U11715 ( .A1(n13948), .A2(n9226), .B1(n13631), .B2(n9239), .ZN(
        n9205) );
  INV_X1 U11716 ( .A(n9210), .ZN(n9211) );
  NAND2_X1 U11717 ( .A1(n9211), .A2(n13439), .ZN(n9212) );
  MUX2_X1 U11718 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n6671), .Z(n9214) );
  XNOR2_X1 U11719 ( .A(n9214), .B(SI_30_), .ZN(n9231) );
  NAND2_X1 U11720 ( .A1(n9214), .A2(SI_30_), .ZN(n9215) );
  MUX2_X1 U11721 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n6671), .Z(n9216) );
  XNOR2_X1 U11722 ( .A(n9216), .B(SI_31_), .ZN(n9217) );
  NAND2_X1 U11723 ( .A1(n8396), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n9218) );
  INV_X1 U11724 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n13724) );
  NAND2_X1 U11725 ( .A1(n9219), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n9222) );
  NAND2_X1 U11726 ( .A1(n9220), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n9221) );
  OAI211_X1 U11727 ( .C1(n9223), .C2(n13724), .A(n9222), .B(n9221), .ZN(n13725) );
  XNOR2_X1 U11728 ( .A(n13729), .B(n13725), .ZN(n9247) );
  OAI22_X1 U11729 ( .A1(n9224), .A2(n9049), .B1(n9225), .B2(n6669), .ZN(n9242)
         );
  INV_X1 U11730 ( .A(n9225), .ZN(n13630) );
  AOI22_X1 U11731 ( .A1(n13744), .A2(n9226), .B1(n13630), .B2(n6669), .ZN(
        n9243) );
  AOI22_X1 U11732 ( .A1(n9242), .A2(n9243), .B1(n9228), .B2(n9227), .ZN(n9229)
         );
  INV_X1 U11733 ( .A(n9231), .ZN(n9232) );
  NAND2_X1 U11734 ( .A1(n14372), .A2(n9234), .ZN(n9236) );
  NAND2_X1 U11735 ( .A1(n8396), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n9235) );
  AOI21_X1 U11736 ( .B1(n9239), .B2(n13725), .A(n9237), .ZN(n9238) );
  OAI22_X1 U11737 ( .A1(n14029), .A2(n9239), .B1(n9240), .B2(n9238), .ZN(n9250) );
  INV_X1 U11738 ( .A(n9240), .ZN(n13629) );
  AOI22_X1 U11739 ( .A1(n13736), .A2(n6669), .B1(n9241), .B2(n13629), .ZN(
        n9249) );
  INV_X1 U11740 ( .A(n9242), .ZN(n9245) );
  INV_X1 U11741 ( .A(n9243), .ZN(n9244) );
  AOI22_X1 U11742 ( .A1(n9250), .A2(n9249), .B1(n9245), .B2(n9244), .ZN(n9246)
         );
  INV_X1 U11743 ( .A(n9250), .ZN(n9251) );
  INV_X1 U11744 ( .A(n9294), .ZN(n9258) );
  OAI21_X1 U11745 ( .B1(n8332), .B2(n9289), .A(n11045), .ZN(n9255) );
  AOI21_X1 U11746 ( .B1(n9256), .B2(n12531), .A(n9255), .ZN(n9257) );
  NAND2_X1 U11747 ( .A1(n9258), .A2(n9257), .ZN(n9263) );
  INV_X1 U11748 ( .A(n10500), .ZN(n10405) );
  NAND2_X1 U11749 ( .A1(n10405), .A2(P2_STATE_REG_SCAN_IN), .ZN(n12298) );
  INV_X1 U11750 ( .A(n12298), .ZN(n9262) );
  MUX2_X1 U11751 ( .A(n7564), .B(n9291), .S(n8333), .Z(n9259) );
  NAND2_X1 U11752 ( .A1(n9259), .A2(n9289), .ZN(n9260) );
  NAND3_X1 U11753 ( .A1(n9263), .A2(n9262), .A3(n9261), .ZN(n9297) );
  INV_X1 U11754 ( .A(n11045), .ZN(n9264) );
  NAND4_X1 U11755 ( .A1(n15470), .A2(n9264), .A3(n13617), .A4(n14081), .ZN(
        n9265) );
  OAI211_X1 U11756 ( .C1(n7564), .C2(n12298), .A(n9265), .B(P2_B_REG_SCAN_IN), 
        .ZN(n9296) );
  XOR2_X1 U11757 ( .A(n13629), .B(n13736), .Z(n9287) );
  NAND2_X1 U11758 ( .A1(n9267), .A2(n9266), .ZN(n13772) );
  XNOR2_X1 U11759 ( .A(n12090), .B(n9268), .ZN(n12055) );
  XNOR2_X1 U11760 ( .A(n14019), .B(n9269), .ZN(n11963) );
  NAND2_X1 U11761 ( .A1(n9031), .A2(n11125), .ZN(n15474) );
  NOR4_X1 U11762 ( .A1(n10864), .A2(n10825), .A3(n12137), .A4(n15474), .ZN(
        n9270) );
  NAND4_X1 U11763 ( .A1(n11526), .A2(n9270), .A3(n10858), .A4(n11087), .ZN(
        n9271) );
  NOR4_X1 U11764 ( .A1(n11638), .A2(n11599), .A3(n9272), .A4(n9271), .ZN(n9274) );
  NAND4_X1 U11765 ( .A1(n9275), .A2(n9274), .A3(n11892), .A4(n9273), .ZN(n9276) );
  NOR4_X1 U11766 ( .A1(n12257), .A2(n12055), .A3(n11963), .A4(n9276), .ZN(
        n9277) );
  NAND4_X1 U11767 ( .A1(n12389), .A2(n12423), .A3(n9277), .A4(n12209), .ZN(
        n9278) );
  NOR4_X1 U11768 ( .A1(n9279), .A2(n13904), .A3(n9278), .A4(n13895), .ZN(n9280) );
  NAND3_X1 U11769 ( .A1(n13828), .A2(n9280), .A3(n13861), .ZN(n9281) );
  NOR4_X1 U11770 ( .A1(n13772), .A2(n9281), .A3(n13848), .A4(n13809), .ZN(
        n9283) );
  NAND4_X1 U11771 ( .A1(n9284), .A2(n9283), .A3(n13760), .A4(n9282), .ZN(n9285) );
  XNOR2_X1 U11772 ( .A(n9290), .B(n9289), .ZN(n9292) );
  NOR3_X1 U11773 ( .A1(n9292), .A2(n9291), .A3(n12298), .ZN(n9293) );
  OAI21_X1 U11774 ( .B1(n9294), .B2(n8333), .A(n9293), .ZN(n9295) );
  NAND3_X1 U11775 ( .A1(n9297), .A2(n9296), .A3(n9295), .ZN(P2_U3328) );
  NAND2_X1 U11776 ( .A1(n9440), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n9453) );
  INV_X1 U11777 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n9452) );
  INV_X1 U11778 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n9506) );
  INV_X1 U11779 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n9520) );
  INV_X1 U11780 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n9594) );
  INV_X1 U11781 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n14164) );
  INV_X1 U11782 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n14098) );
  INV_X1 U11783 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n14155) );
  INV_X1 U11784 ( .A(n9670), .ZN(n9304) );
  NAND2_X1 U11785 ( .A1(n9304), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n9341) );
  INV_X1 U11786 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n9305) );
  NAND2_X1 U11787 ( .A1(n9341), .A2(n9305), .ZN(n9306) );
  NOR2_X1 U11788 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n9308) );
  INV_X2 U11789 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n10298) );
  NAND4_X1 U11790 ( .A1(n9545), .A2(n9489), .A3(n9436), .A4(n9515), .ZN(n9309)
         );
  NOR2_X2 U11791 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n9379) );
  NAND4_X1 U11792 ( .A1(n9313), .A2(n9312), .A3(n9411), .A4(n9311), .ZN(n9314)
         );
  NOR2_X1 U11793 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), 
        .ZN(n9317) );
  NOR2_X1 U11794 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), 
        .ZN(n9316) );
  NAND4_X1 U11795 ( .A1(n9700), .A2(n9317), .A3(n9316), .A4(n9315), .ZN(n9755)
         );
  INV_X1 U11796 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n9318) );
  INV_X1 U11797 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n9321) );
  INV_X1 U11798 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n9322) );
  AND2_X4 U11799 ( .A1(n9324), .A2(n9325), .ZN(n9657) );
  NAND2_X1 U11800 ( .A1(n14088), .A2(n9657), .ZN(n9331) );
  INV_X1 U11801 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n9328) );
  INV_X2 U11802 ( .A(n9392), .ZN(n14375) );
  NAND2_X1 U11803 ( .A1(n14375), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n9327) );
  AND2_X2 U11804 ( .A1(n14878), .A2(n14881), .ZN(n9418) );
  NAND2_X1 U11805 ( .A1(n9633), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n9326) );
  OAI211_X1 U11806 ( .C1(n9328), .C2(n14380), .A(n9327), .B(n9326), .ZN(n9329)
         );
  INV_X1 U11807 ( .A(n9329), .ZN(n9330) );
  INV_X1 U11808 ( .A(n14481), .ZN(n14192) );
  MUX2_X2 U11809 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9333), .S(
        P1_IR_REG_28__SCAN_IN), .Z(n9335) );
  INV_X1 U11810 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n9336) );
  NAND2_X1 U11811 ( .A1(n14079), .A2(n14407), .ZN(n9339) );
  INV_X1 U11812 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n14886) );
  OR2_X1 U11813 ( .A1(n14408), .A2(n14886), .ZN(n9338) );
  INV_X1 U11814 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n14193) );
  NAND2_X1 U11815 ( .A1(n9670), .A2(n14193), .ZN(n9340) );
  NAND2_X1 U11816 ( .A1(n9341), .A2(n9340), .ZN(n14652) );
  OR2_X1 U11817 ( .A1(n14652), .A2(n9692), .ZN(n9347) );
  INV_X1 U11818 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n9344) );
  NAND2_X1 U11819 ( .A1(n14376), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n9343) );
  NAND2_X1 U11820 ( .A1(n14375), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n9342) );
  OAI211_X1 U11821 ( .C1(n14380), .C2(n9344), .A(n9343), .B(n9342), .ZN(n9345)
         );
  INV_X1 U11822 ( .A(n9345), .ZN(n9346) );
  NAND2_X1 U11823 ( .A1(n12478), .A2(n14407), .ZN(n9349) );
  OR2_X1 U11824 ( .A1(n14408), .A2(n14890), .ZN(n9348) );
  NAND2_X1 U11825 ( .A1(n12025), .A2(n14407), .ZN(n9355) );
  NAND2_X1 U11826 ( .A1(n9350), .A2(P1_IR_REG_19__SCAN_IN), .ZN(n9353) );
  INV_X1 U11827 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n9351) );
  NAND2_X1 U11828 ( .A1(n9352), .A2(n9351), .ZN(n9708) );
  AOI22_X1 U11829 ( .A1(n9591), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n14209), 
        .B2(n9590), .ZN(n9354) );
  INV_X1 U11830 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n9356) );
  NAND2_X1 U11831 ( .A1(n9597), .A2(n9356), .ZN(n9357) );
  NAND2_X1 U11832 ( .A1(n9607), .A2(n9357), .ZN(n14764) );
  OR2_X1 U11833 ( .A1(n14764), .A2(n9692), .ZN(n9363) );
  INV_X1 U11834 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9360) );
  NAND2_X1 U11835 ( .A1(n14375), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n9359) );
  NAND2_X1 U11836 ( .A1(n9633), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n9358) );
  OAI211_X1 U11837 ( .C1(n14380), .C2(n9360), .A(n9359), .B(n9358), .ZN(n9361)
         );
  INV_X1 U11838 ( .A(n9361), .ZN(n9362) );
  OR2_X1 U11839 ( .A1(n14758), .A2(n14162), .ZN(n14332) );
  NAND2_X1 U11840 ( .A1(n14758), .A2(n14162), .ZN(n14331) );
  NAND2_X1 U11841 ( .A1(n9383), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n9367) );
  NAND2_X1 U11842 ( .A1(n9657), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n9366) );
  NAND2_X1 U11843 ( .A1(n9418), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n9365) );
  NAND2_X1 U11844 ( .A1(n9582), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n9364) );
  INV_X1 U11845 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n9369) );
  NAND2_X1 U11846 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n9368) );
  XNOR2_X1 U11847 ( .A(n9369), .B(n9368), .ZN(n14512) );
  INV_X2 U11848 ( .A(n11189), .ZN(n10815) );
  NAND2_X1 U11849 ( .A1(n9657), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n9375) );
  NAND2_X1 U11850 ( .A1(n9383), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n9374) );
  NAND2_X1 U11851 ( .A1(n9418), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n9373) );
  NAND2_X1 U11852 ( .A1(n9582), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n9372) );
  NOR2_X1 U11853 ( .A1(n6671), .A2(n10454), .ZN(n9377) );
  XNOR2_X1 U11854 ( .A(n9377), .B(n9376), .ZN(n14893) );
  MUX2_X1 U11855 ( .A(P1_IR_REG_0__SCAN_IN), .B(n14893), .S(n10483), .Z(n10730) );
  NAND2_X1 U11856 ( .A1(n14418), .A2(n11180), .ZN(n11179) );
  NAND2_X1 U11857 ( .A1(n11208), .A2(n10815), .ZN(n9378) );
  NAND2_X1 U11858 ( .A1(n11179), .A2(n9378), .ZN(n11211) );
  INV_X1 U11859 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9424) );
  OR2_X1 U11860 ( .A1(n9379), .A2(n9424), .ZN(n9380) );
  XNOR2_X1 U11861 ( .A(n9380), .B(P1_IR_REG_2__SCAN_IN), .ZN(n14530) );
  AOI22_X1 U11862 ( .A1(n9591), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(n9590), .B2(
        n14530), .ZN(n9381) );
  NAND2_X1 U11863 ( .A1(n9383), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n9387) );
  NAND2_X1 U11864 ( .A1(n9418), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n9385) );
  NAND2_X1 U11865 ( .A1(n9582), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n9384) );
  NAND2_X1 U11866 ( .A1(n11211), .A2(n11210), .ZN(n11209) );
  NOR2_X1 U11867 ( .A1(n14224), .A2(n14502), .ZN(n14227) );
  INV_X1 U11868 ( .A(n14227), .ZN(n9388) );
  NAND2_X1 U11869 ( .A1(n11209), .A2(n9388), .ZN(n11099) );
  OR2_X1 U11870 ( .A1(n10440), .A2(n9370), .ZN(n9391) );
  NAND2_X1 U11871 ( .A1(n9398), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9389) );
  XNOR2_X1 U11872 ( .A(n9389), .B(P1_IR_REG_3__SCAN_IN), .ZN(n14546) );
  AOI22_X1 U11873 ( .A1(n9591), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(n9590), .B2(
        n14546), .ZN(n9390) );
  NAND2_X1 U11874 ( .A1(n9383), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n9396) );
  INV_X1 U11875 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n14539) );
  NAND2_X1 U11876 ( .A1(n9657), .A2(n14539), .ZN(n9395) );
  NAND2_X1 U11877 ( .A1(n14376), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n9394) );
  NAND2_X1 U11878 ( .A1(n9582), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n9393) );
  OR2_X1 U11879 ( .A1(n14500), .A2(n14228), .ZN(n9397) );
  OR2_X1 U11880 ( .A1(n10435), .A2(n9370), .ZN(n9401) );
  NAND2_X1 U11881 ( .A1(n9409), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9399) );
  XNOR2_X1 U11882 ( .A(n9399), .B(P1_IR_REG_4__SCAN_IN), .ZN(n15231) );
  AOI22_X1 U11883 ( .A1(n9591), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n9590), .B2(
        n15231), .ZN(n9400) );
  NAND2_X1 U11884 ( .A1(n9401), .A2(n9400), .ZN(n14233) );
  INV_X1 U11885 ( .A(n14233), .ZN(n15288) );
  NAND2_X1 U11886 ( .A1(n6841), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n9406) );
  NAND2_X1 U11887 ( .A1(n14375), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n9405) );
  NOR2_X1 U11888 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n9402) );
  NOR2_X1 U11889 ( .A1(n9416), .A2(n9402), .ZN(n11716) );
  NAND2_X1 U11890 ( .A1(n9657), .A2(n11716), .ZN(n9404) );
  NAND2_X1 U11891 ( .A1(n14376), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n9403) );
  NAND4_X1 U11892 ( .A1(n9406), .A2(n9405), .A3(n9404), .A4(n9403), .ZN(n14499) );
  INV_X1 U11893 ( .A(n14499), .ZN(n9718) );
  OAI21_X1 U11894 ( .B1(n11340), .B2(n15288), .A(n9718), .ZN(n9408) );
  NAND2_X1 U11895 ( .A1(n11340), .A2(n15288), .ZN(n9407) );
  NAND2_X1 U11896 ( .A1(n10442), .A2(n14407), .ZN(n9415) );
  NOR2_X1 U11897 ( .A1(n9412), .A2(n9424), .ZN(n9410) );
  MUX2_X1 U11898 ( .A(n9424), .B(n9410), .S(P1_IR_REG_5__SCAN_IN), .Z(n9413)
         );
  OR2_X1 U11899 ( .A1(n9413), .A2(n9560), .ZN(n14562) );
  INV_X1 U11900 ( .A(n14562), .ZN(n14557) );
  AOI22_X1 U11901 ( .A1(n9591), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n9590), .B2(
        n14557), .ZN(n9414) );
  NAND2_X1 U11902 ( .A1(n9415), .A2(n9414), .ZN(n15293) );
  NAND2_X1 U11903 ( .A1(n14375), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n9422) );
  NAND2_X1 U11904 ( .A1(n6841), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n9421) );
  OAI21_X1 U11905 ( .B1(n9416), .B2(P1_REG3_REG_5__SCAN_IN), .A(n9429), .ZN(
        n11744) );
  INV_X1 U11906 ( .A(n11744), .ZN(n9417) );
  NAND2_X1 U11907 ( .A1(n9657), .A2(n9417), .ZN(n9420) );
  NAND2_X1 U11908 ( .A1(n14376), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n9419) );
  XNOR2_X1 U11909 ( .A(n15293), .B(n11445), .ZN(n14425) );
  OR2_X1 U11910 ( .A1(n15293), .A2(n14498), .ZN(n9423) );
  OR2_X1 U11911 ( .A1(n10437), .A2(n9370), .ZN(n9427) );
  OR2_X1 U11912 ( .A1(n9560), .A2(n9424), .ZN(n9425) );
  XNOR2_X1 U11913 ( .A(n9425), .B(P1_IR_REG_6__SCAN_IN), .ZN(n10584) );
  AOI22_X1 U11914 ( .A1(n9591), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n9590), .B2(
        n10584), .ZN(n9426) );
  NAND2_X1 U11915 ( .A1(n9427), .A2(n9426), .ZN(n14250) );
  NAND2_X1 U11916 ( .A1(n6841), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n9434) );
  NAND2_X1 U11917 ( .A1(n14375), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n9433) );
  AND2_X1 U11918 ( .A1(n9429), .A2(n9428), .ZN(n9430) );
  NOR2_X1 U11919 ( .A1(n9440), .A2(n9430), .ZN(n11939) );
  NAND2_X1 U11920 ( .A1(n9657), .A2(n11939), .ZN(n9432) );
  NAND2_X1 U11921 ( .A1(n9633), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n9431) );
  XNOR2_X1 U11922 ( .A(n14250), .B(n14497), .ZN(n14426) );
  INV_X1 U11923 ( .A(n14250), .ZN(n15303) );
  INV_X1 U11924 ( .A(n14497), .ZN(n11933) );
  NAND2_X1 U11925 ( .A1(n15303), .A2(n11933), .ZN(n9435) );
  OR2_X1 U11926 ( .A1(n10460), .A2(n9370), .ZN(n9439) );
  NAND2_X1 U11927 ( .A1(n9560), .A2(n9436), .ZN(n9491) );
  NAND2_X1 U11928 ( .A1(n9491), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9437) );
  XNOR2_X1 U11929 ( .A(n9437), .B(n10312), .ZN(n10596) );
  AOI22_X1 U11930 ( .A1(n9591), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n9590), .B2(
        n10596), .ZN(n9438) );
  NAND2_X1 U11931 ( .A1(n9439), .A2(n9438), .ZN(n15309) );
  NAND2_X1 U11932 ( .A1(n6841), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n9445) );
  NAND2_X1 U11933 ( .A1(n14375), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n9444) );
  OR2_X1 U11934 ( .A1(n9440), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n9441) );
  AND2_X1 U11935 ( .A1(n9453), .A2(n9441), .ZN(n11486) );
  NAND2_X1 U11936 ( .A1(n9657), .A2(n11486), .ZN(n9443) );
  NAND2_X1 U11937 ( .A1(n14376), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n9442) );
  NAND4_X1 U11938 ( .A1(n9445), .A2(n9444), .A3(n9443), .A4(n9442), .ZN(n14496) );
  XNOR2_X1 U11939 ( .A(n15309), .B(n14496), .ZN(n14427) );
  INV_X1 U11940 ( .A(n14427), .ZN(n9446) );
  OR2_X1 U11941 ( .A1(n15309), .A2(n14496), .ZN(n9447) );
  NAND2_X1 U11942 ( .A1(n9448), .A2(n9447), .ZN(n11619) );
  OR2_X1 U11943 ( .A1(n10471), .A2(n9370), .ZN(n9451) );
  OR2_X1 U11944 ( .A1(n9491), .A2(n10312), .ZN(n9449) );
  NAND2_X1 U11945 ( .A1(n9449), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9461) );
  XNOR2_X1 U11946 ( .A(n9461), .B(P1_IR_REG_8__SCAN_IN), .ZN(n14576) );
  AOI22_X1 U11947 ( .A1(n9591), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n9590), .B2(
        n14576), .ZN(n9450) );
  NAND2_X1 U11948 ( .A1(n9451), .A2(n9450), .ZN(n14262) );
  NAND2_X1 U11949 ( .A1(n6841), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n9458) );
  NAND2_X1 U11950 ( .A1(n14375), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n9457) );
  NAND2_X1 U11951 ( .A1(n9453), .A2(n9452), .ZN(n9454) );
  AND2_X1 U11952 ( .A1(n9468), .A2(n9454), .ZN(n12173) );
  NAND2_X1 U11953 ( .A1(n9657), .A2(n12173), .ZN(n9456) );
  NAND2_X1 U11954 ( .A1(n14376), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n9455) );
  NAND4_X1 U11955 ( .A1(n9458), .A2(n9457), .A3(n9456), .A4(n9455), .ZN(n14495) );
  XNOR2_X1 U11956 ( .A(n14262), .B(n14495), .ZN(n14429) );
  INV_X1 U11957 ( .A(n14429), .ZN(n11618) );
  NAND2_X1 U11958 ( .A1(n11619), .A2(n11618), .ZN(n9460) );
  OR2_X1 U11959 ( .A1(n14262), .A2(n14495), .ZN(n9459) );
  NAND2_X1 U11960 ( .A1(n9460), .A2(n9459), .ZN(n11910) );
  NAND2_X1 U11961 ( .A1(n10487), .A2(n14407), .ZN(n9466) );
  INV_X1 U11962 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n10052) );
  NAND2_X1 U11963 ( .A1(n9461), .A2(n10052), .ZN(n9462) );
  NAND2_X1 U11964 ( .A1(n9462), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9463) );
  NAND2_X1 U11965 ( .A1(n9463), .A2(n10191), .ZN(n9476) );
  OR2_X1 U11966 ( .A1(n9463), .A2(n10191), .ZN(n9464) );
  AOI22_X1 U11967 ( .A1(n9590), .A2(n14594), .B1(n9591), .B2(
        P2_DATAO_REG_9__SCAN_IN), .ZN(n9465) );
  NAND2_X1 U11968 ( .A1(n9466), .A2(n9465), .ZN(n14266) );
  NAND2_X1 U11969 ( .A1(n14375), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n9473) );
  NAND2_X1 U11970 ( .A1(n6841), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n9472) );
  AND2_X1 U11971 ( .A1(n9468), .A2(n9467), .ZN(n9469) );
  NOR2_X1 U11972 ( .A1(n9480), .A2(n9469), .ZN(n12351) );
  NAND2_X1 U11973 ( .A1(n9657), .A2(n12351), .ZN(n9471) );
  NAND2_X1 U11974 ( .A1(n14376), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n9470) );
  NAND4_X1 U11975 ( .A1(n9473), .A2(n9472), .A3(n9471), .A4(n9470), .ZN(n14494) );
  INV_X1 U11976 ( .A(n14494), .ZN(n9729) );
  XNOR2_X1 U11977 ( .A(n14266), .B(n9729), .ZN(n14431) );
  NAND2_X1 U11978 ( .A1(n11910), .A2(n14431), .ZN(n9475) );
  OR2_X1 U11979 ( .A1(n14266), .A2(n14494), .ZN(n9474) );
  OR2_X1 U11980 ( .A1(n10492), .A2(n9370), .ZN(n9479) );
  NAND2_X1 U11981 ( .A1(n9476), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9477) );
  XNOR2_X1 U11982 ( .A(n9477), .B(P1_IR_REG_10__SCAN_IN), .ZN(n10605) );
  AOI22_X1 U11983 ( .A1(n10605), .A2(n9590), .B1(n9591), .B2(
        P2_DATAO_REG_10__SCAN_IN), .ZN(n9478) );
  NAND2_X1 U11984 ( .A1(n6841), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n9485) );
  NAND2_X1 U11985 ( .A1(n14375), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n9484) );
  NOR2_X1 U11986 ( .A1(n9480), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n9481) );
  NAND2_X1 U11987 ( .A1(n9657), .A2(n7677), .ZN(n9483) );
  NAND2_X1 U11988 ( .A1(n14376), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n9482) );
  NAND4_X1 U11989 ( .A1(n9485), .A2(n9484), .A3(n9483), .A4(n9482), .ZN(n14493) );
  XNOR2_X1 U11990 ( .A(n14275), .B(n12492), .ZN(n14432) );
  OR2_X1 U11991 ( .A1(n14275), .A2(n14493), .ZN(n9486) );
  NAND2_X1 U11992 ( .A1(n10496), .A2(n14407), .ZN(n9495) );
  INV_X1 U11993 ( .A(n10312), .ZN(n9488) );
  NAND4_X1 U11994 ( .A1(n9489), .A2(n10191), .A3(n10052), .A4(n9488), .ZN(
        n9490) );
  NAND2_X1 U11995 ( .A1(n9547), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9492) );
  XNOR2_X1 U11996 ( .A(n9492), .B(n10298), .ZN(n10890) );
  OAI22_X1 U11997 ( .A1(n14408), .A2(n10497), .B1(n10890), .B2(n10483), .ZN(
        n9493) );
  INV_X1 U11998 ( .A(n9493), .ZN(n9494) );
  NAND2_X1 U11999 ( .A1(n14375), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n9501) );
  OR2_X1 U12000 ( .A1(n9496), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n9497) );
  AND2_X1 U12001 ( .A1(n9507), .A2(n9497), .ZN(n12494) );
  NAND2_X1 U12002 ( .A1(n9657), .A2(n12494), .ZN(n9500) );
  NAND2_X1 U12003 ( .A1(n14376), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n9499) );
  NAND2_X1 U12004 ( .A1(n6841), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n9498) );
  NAND4_X1 U12005 ( .A1(n9501), .A2(n9500), .A3(n9499), .A4(n9498), .ZN(n14492) );
  INV_X1 U12006 ( .A(n14492), .ZN(n9731) );
  XNOR2_X1 U12007 ( .A(n14279), .B(n9731), .ZN(n14433) );
  OR2_X1 U12008 ( .A1(n14279), .A2(n14492), .ZN(n9502) );
  NAND2_X1 U12009 ( .A1(n10745), .A2(n14407), .ZN(n9505) );
  NAND2_X1 U12010 ( .A1(n9503), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9513) );
  XNOR2_X1 U12011 ( .A(n9513), .B(P1_IR_REG_12__SCAN_IN), .ZN(n10891) );
  AOI22_X1 U12012 ( .A1(n9591), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n10891), 
        .B2(n9590), .ZN(n9504) );
  NAND2_X1 U12013 ( .A1(n6841), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n9512) );
  NAND2_X1 U12014 ( .A1(n14375), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n9511) );
  NAND2_X1 U12015 ( .A1(n9507), .A2(n9506), .ZN(n9508) );
  AND2_X1 U12016 ( .A1(n9521), .A2(n9508), .ZN(n14930) );
  NAND2_X1 U12017 ( .A1(n9657), .A2(n14930), .ZN(n9510) );
  NAND2_X1 U12018 ( .A1(n9633), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n9509) );
  NAND4_X1 U12019 ( .A1(n9512), .A2(n9511), .A3(n9510), .A4(n9509), .ZN(n15108) );
  INV_X1 U12020 ( .A(n15108), .ZN(n14946) );
  XNOR2_X1 U12021 ( .A(n14917), .B(n14946), .ZN(n14923) );
  NAND2_X1 U12022 ( .A1(n10836), .A2(n14407), .ZN(n9519) );
  NAND2_X1 U12023 ( .A1(n9513), .A2(n9545), .ZN(n9514) );
  NAND2_X1 U12024 ( .A1(n9514), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9516) );
  NAND2_X1 U12025 ( .A1(n9516), .A2(n10050), .ZN(n9531) );
  OAI21_X1 U12026 ( .B1(n9516), .B2(n10050), .A(n9531), .ZN(n11255) );
  OAI22_X1 U12027 ( .A1(n11255), .A2(n10483), .B1(n14408), .B2(n10838), .ZN(
        n9517) );
  INV_X1 U12028 ( .A(n9517), .ZN(n9518) );
  INV_X1 U12029 ( .A(n15112), .ZN(n15172) );
  AND2_X1 U12030 ( .A1(n9521), .A2(n9520), .ZN(n9522) );
  OR2_X1 U12031 ( .A1(n9537), .A2(n9522), .ZN(n15118) );
  NAND2_X1 U12032 ( .A1(n14375), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n9523) );
  OAI21_X1 U12033 ( .B1(n15118), .B2(n9692), .A(n9523), .ZN(n9524) );
  INV_X1 U12034 ( .A(n9524), .ZN(n9528) );
  NAND2_X1 U12035 ( .A1(n9633), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n9526) );
  NAND2_X1 U12036 ( .A1(n6841), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n9525) );
  AND2_X1 U12037 ( .A1(n9526), .A2(n9525), .ZN(n9527) );
  XNOR2_X1 U12038 ( .A(n15172), .B(n14491), .ZN(n14954) );
  INV_X1 U12039 ( .A(n14954), .ZN(n14952) );
  NAND2_X1 U12040 ( .A1(n15112), .A2(n15087), .ZN(n9529) );
  NAND2_X1 U12041 ( .A1(n9530), .A2(n9529), .ZN(n12232) );
  NAND2_X1 U12042 ( .A1(n11350), .A2(n14407), .ZN(n9534) );
  NAND2_X1 U12043 ( .A1(n9531), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9532) );
  XNOR2_X1 U12044 ( .A(n9532), .B(P1_IR_REG_14__SCAN_IN), .ZN(n11718) );
  AOI22_X1 U12045 ( .A1(n11718), .A2(n9590), .B1(n9591), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n9533) );
  NAND2_X1 U12046 ( .A1(n6841), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n9536) );
  NAND2_X1 U12047 ( .A1(n14375), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n9535) );
  AND2_X1 U12048 ( .A1(n9536), .A2(n9535), .ZN(n9543) );
  INV_X1 U12049 ( .A(n9537), .ZN(n9539) );
  INV_X1 U12050 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n9538) );
  NAND2_X1 U12051 ( .A1(n9539), .A2(n9538), .ZN(n9540) );
  NAND2_X1 U12052 ( .A1(n9551), .A2(n9540), .ZN(n15100) );
  OR2_X1 U12053 ( .A1(n15100), .A2(n9692), .ZN(n9542) );
  NAND2_X1 U12054 ( .A1(n9633), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n9541) );
  OR2_X1 U12055 ( .A1(n15164), .A2(n14948), .ZN(n14299) );
  NAND2_X1 U12056 ( .A1(n15164), .A2(n14948), .ZN(n14300) );
  NAND2_X1 U12057 ( .A1(n14299), .A2(n14300), .ZN(n14298) );
  INV_X1 U12058 ( .A(n14948), .ZN(n15106) );
  NAND2_X1 U12059 ( .A1(n15164), .A2(n15106), .ZN(n9544) );
  NAND2_X1 U12060 ( .A1(n11546), .A2(n14407), .ZN(n9550) );
  INV_X1 U12061 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n10277) );
  NAND4_X1 U12062 ( .A1(n10298), .A2(n10050), .A3(n9545), .A4(n10277), .ZN(
        n9546) );
  OAI21_X1 U12063 ( .B1(n9547), .B2(n9546), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n9548) );
  XNOR2_X1 U12064 ( .A(n9548), .B(P1_IR_REG_15__SCAN_IN), .ZN(n12004) );
  AOI22_X1 U12065 ( .A1(n9591), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n12004), 
        .B2(n9590), .ZN(n9549) );
  INV_X1 U12066 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n14202) );
  NAND2_X1 U12067 ( .A1(n9551), .A2(n14202), .ZN(n9552) );
  NAND2_X1 U12068 ( .A1(n9567), .A2(n9552), .ZN(n14201) );
  OR2_X1 U12069 ( .A1(n14201), .A2(n9692), .ZN(n9555) );
  AOI22_X1 U12070 ( .A1(n6841), .A2(P1_REG1_REG_15__SCAN_IN), .B1(n14375), 
        .B2(P1_REG2_REG_15__SCAN_IN), .ZN(n9554) );
  NAND2_X1 U12071 ( .A1(n9633), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n9553) );
  NAND2_X1 U12072 ( .A1(n12552), .A2(n15132), .ZN(n14304) );
  INV_X1 U12073 ( .A(n15132), .ZN(n14490) );
  OR2_X1 U12074 ( .A1(n12552), .A2(n14490), .ZN(n9557) );
  NAND2_X1 U12075 ( .A1(n11688), .A2(n14407), .ZN(n9564) );
  NAND2_X1 U12076 ( .A1(n9560), .A2(n9559), .ZN(n9561) );
  NAND2_X1 U12077 ( .A1(n9561), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9562) );
  XNOR2_X1 U12078 ( .A(n9562), .B(P1_IR_REG_16__SCAN_IN), .ZN(n12008) );
  AOI22_X1 U12079 ( .A1(n9591), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n9590), 
        .B2(n12008), .ZN(n9563) );
  INV_X1 U12080 ( .A(n9565), .ZN(n9580) );
  INV_X1 U12081 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n9566) );
  NAND2_X1 U12082 ( .A1(n9567), .A2(n9566), .ZN(n9568) );
  NAND2_X1 U12083 ( .A1(n9580), .A2(n9568), .ZN(n15137) );
  AOI22_X1 U12084 ( .A1(n6841), .A2(P1_REG1_REG_16__SCAN_IN), .B1(n14375), 
        .B2(P1_REG2_REG_16__SCAN_IN), .ZN(n9570) );
  NAND2_X1 U12085 ( .A1(n9633), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n9569) );
  OAI211_X1 U12086 ( .C1(n15137), .C2(n9692), .A(n9570), .B(n9569), .ZN(n14489) );
  INV_X1 U12087 ( .A(n14489), .ZN(n14307) );
  XNOR2_X1 U12088 ( .A(n14309), .B(n14307), .ZN(n15130) );
  OR2_X1 U12089 ( .A1(n14309), .A2(n14489), .ZN(n9571) );
  NAND2_X1 U12090 ( .A1(n11732), .A2(n14407), .ZN(n9578) );
  NAND2_X1 U12091 ( .A1(n9573), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9574) );
  MUX2_X1 U12092 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9574), .S(
        P1_IR_REG_17__SCAN_IN), .Z(n9576) );
  AND2_X1 U12093 ( .A1(n9576), .A2(n9575), .ZN(n14605) );
  AOI22_X1 U12094 ( .A1(n9591), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n9590), 
        .B2(n14605), .ZN(n9577) );
  INV_X1 U12095 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n9579) );
  NAND2_X1 U12096 ( .A1(n9580), .A2(n9579), .ZN(n9581) );
  NAND2_X1 U12097 ( .A1(n9595), .A2(n9581), .ZN(n14147) );
  OR2_X1 U12098 ( .A1(n14147), .A2(n9692), .ZN(n9587) );
  INV_X1 U12099 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n12446) );
  NAND2_X1 U12100 ( .A1(n6841), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n9584) );
  NAND2_X1 U12101 ( .A1(n9633), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n9583) );
  OAI211_X1 U12102 ( .C1(n9392), .C2(n12446), .A(n9584), .B(n9583), .ZN(n9585)
         );
  INV_X1 U12103 ( .A(n9585), .ZN(n9586) );
  NAND2_X1 U12104 ( .A1(n9587), .A2(n9586), .ZN(n15135) );
  OR2_X1 U12105 ( .A1(n14851), .A2(n15135), .ZN(n9714) );
  INV_X1 U12106 ( .A(n9714), .ZN(n9588) );
  NAND2_X1 U12107 ( .A1(n14851), .A2(n15135), .ZN(n9713) );
  NAND2_X1 U12108 ( .A1(n11979), .A2(n14407), .ZN(n9593) );
  NAND2_X1 U12109 ( .A1(n9575), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9589) );
  XNOR2_X1 U12110 ( .A(n9589), .B(P1_IR_REG_18__SCAN_IN), .ZN(n14611) );
  AOI22_X1 U12111 ( .A1(n9591), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n9590), 
        .B2(n14611), .ZN(n9592) );
  NAND2_X1 U12112 ( .A1(n9595), .A2(n9594), .ZN(n9596) );
  AND2_X1 U12113 ( .A1(n9597), .A2(n9596), .ZN(n14181) );
  NAND2_X1 U12114 ( .A1(n14181), .A2(n9657), .ZN(n9603) );
  INV_X1 U12115 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9600) );
  NAND2_X1 U12116 ( .A1(n14375), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9599) );
  NAND2_X1 U12117 ( .A1(n9633), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n9598) );
  OAI211_X1 U12118 ( .C1(n9600), .C2(n14380), .A(n9599), .B(n9598), .ZN(n9601)
         );
  INV_X1 U12119 ( .A(n9601), .ZN(n9602) );
  AND2_X1 U12120 ( .A1(n9603), .A2(n9602), .ZN(n14324) );
  NAND2_X1 U12121 ( .A1(n14845), .A2(n14761), .ZN(n14329) );
  INV_X1 U12122 ( .A(n14329), .ZN(n9604) );
  OR2_X1 U12123 ( .A1(n14845), .A2(n14761), .ZN(n14326) );
  INV_X1 U12124 ( .A(n14162), .ZN(n14488) );
  NAND2_X1 U12125 ( .A1(n12015), .A2(n14407), .ZN(n9606) );
  INV_X1 U12126 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n12016) );
  OR2_X1 U12127 ( .A1(n14408), .A2(n12016), .ZN(n9605) );
  NAND2_X1 U12128 ( .A1(n9607), .A2(n14164), .ZN(n9608) );
  AND2_X1 U12129 ( .A1(n9619), .A2(n9608), .ZN(n14744) );
  NAND2_X1 U12130 ( .A1(n14744), .A2(n9657), .ZN(n9614) );
  INV_X1 U12131 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n9611) );
  NAND2_X1 U12132 ( .A1(n14375), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n9610) );
  NAND2_X1 U12133 ( .A1(n9633), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n9609) );
  OAI211_X1 U12134 ( .C1(n14380), .C2(n9611), .A(n9610), .B(n9609), .ZN(n9612)
         );
  INV_X1 U12135 ( .A(n9612), .ZN(n9613) );
  INV_X1 U12136 ( .A(n14336), .ZN(n14763) );
  XNOR2_X1 U12137 ( .A(n14832), .B(n14763), .ZN(n14747) );
  OR2_X1 U12138 ( .A1(n14746), .A2(n14336), .ZN(n9615) );
  NAND2_X1 U12139 ( .A1(n12153), .A2(n14407), .ZN(n9617) );
  OR2_X1 U12140 ( .A1(n14408), .A2(n12154), .ZN(n9616) );
  INV_X1 U12141 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n9618) );
  NAND2_X1 U12142 ( .A1(n9619), .A2(n9618), .ZN(n9620) );
  NAND2_X1 U12143 ( .A1(n9631), .A2(n9620), .ZN(n14730) );
  OR2_X1 U12144 ( .A1(n14730), .A2(n9692), .ZN(n9626) );
  INV_X1 U12145 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n9623) );
  NAND2_X1 U12146 ( .A1(n14375), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n9622) );
  NAND2_X1 U12147 ( .A1(n9633), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n9621) );
  OAI211_X1 U12148 ( .C1(n9623), .C2(n14380), .A(n9622), .B(n9621), .ZN(n9624)
         );
  INV_X1 U12149 ( .A(n9624), .ZN(n9625) );
  NAND2_X1 U12150 ( .A1(n9626), .A2(n9625), .ZN(n14487) );
  XNOR2_X1 U12151 ( .A(n14827), .B(n14487), .ZN(n14442) );
  OR2_X1 U12152 ( .A1(n14827), .A2(n14487), .ZN(n9627) );
  INV_X1 U12153 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9630) );
  NAND2_X1 U12154 ( .A1(n9631), .A2(n9630), .ZN(n9632) );
  NAND2_X1 U12155 ( .A1(n9643), .A2(n9632), .ZN(n14713) );
  OR2_X1 U12156 ( .A1(n14713), .A2(n9692), .ZN(n9639) );
  INV_X1 U12157 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n9636) );
  NAND2_X1 U12158 ( .A1(n9633), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n9635) );
  NAND2_X1 U12159 ( .A1(n14375), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n9634) );
  OAI211_X1 U12160 ( .C1(n14380), .C2(n9636), .A(n9635), .B(n9634), .ZN(n9637)
         );
  INV_X1 U12161 ( .A(n9637), .ZN(n9638) );
  INV_X1 U12162 ( .A(n14705), .ZN(n9651) );
  NAND2_X1 U12163 ( .A1(n12301), .A2(n14407), .ZN(n9642) );
  INV_X1 U12164 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n12303) );
  OR2_X1 U12165 ( .A1(n14408), .A2(n12303), .ZN(n9641) );
  NAND2_X1 U12166 ( .A1(n9643), .A2(n14098), .ZN(n9644) );
  NAND2_X1 U12167 ( .A1(n9655), .A2(n9644), .ZN(n14699) );
  OR2_X1 U12168 ( .A1(n14699), .A2(n9692), .ZN(n9650) );
  INV_X1 U12169 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n9647) );
  NAND2_X1 U12170 ( .A1(n14375), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n9646) );
  NAND2_X1 U12171 ( .A1(n14376), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n9645) );
  OAI211_X1 U12172 ( .C1(n9647), .C2(n14380), .A(n9646), .B(n9645), .ZN(n9648)
         );
  INV_X1 U12173 ( .A(n9648), .ZN(n9649) );
  NAND2_X1 U12174 ( .A1(n9650), .A2(n9649), .ZN(n14485) );
  INV_X1 U12175 ( .A(n14485), .ZN(n14174) );
  XNOR2_X1 U12176 ( .A(n14812), .B(n14174), .ZN(n14694) );
  INV_X1 U12177 ( .A(n14694), .ZN(n14704) );
  NAND2_X1 U12178 ( .A1(n14812), .A2(n14485), .ZN(n9652) );
  NAND2_X1 U12179 ( .A1(n12325), .A2(n14407), .ZN(n9654) );
  OR2_X1 U12180 ( .A1(n14408), .A2(n7281), .ZN(n9653) );
  NAND2_X1 U12181 ( .A1(n9655), .A2(n14155), .ZN(n9656) );
  AND2_X1 U12182 ( .A1(n9668), .A2(n9656), .ZN(n14687) );
  NAND2_X1 U12183 ( .A1(n14687), .A2(n9657), .ZN(n9663) );
  INV_X1 U12184 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n9660) );
  NAND2_X1 U12185 ( .A1(n14376), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n9659) );
  NAND2_X1 U12186 ( .A1(n14375), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n9658) );
  OAI211_X1 U12187 ( .C1(n14380), .C2(n9660), .A(n9659), .B(n9658), .ZN(n9661)
         );
  INV_X1 U12188 ( .A(n9661), .ZN(n9662) );
  XNOR2_X1 U12189 ( .A(n14806), .B(n14665), .ZN(n14683) );
  NAND2_X1 U12190 ( .A1(n14690), .A2(n14665), .ZN(n9664) );
  NAND2_X1 U12191 ( .A1(n12379), .A2(n14407), .ZN(n9666) );
  OR2_X1 U12192 ( .A1(n14408), .A2(n12381), .ZN(n9665) );
  INV_X1 U12193 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n9667) );
  NAND2_X1 U12194 ( .A1(n9668), .A2(n9667), .ZN(n9669) );
  NAND2_X1 U12195 ( .A1(n9670), .A2(n9669), .ZN(n14672) );
  OR2_X1 U12196 ( .A1(n14672), .A2(n9692), .ZN(n9676) );
  INV_X1 U12197 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n9673) );
  NAND2_X1 U12198 ( .A1(n14375), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n9672) );
  NAND2_X1 U12199 ( .A1(n14376), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n9671) );
  OAI211_X1 U12200 ( .C1(n9673), .C2(n14380), .A(n9672), .B(n9671), .ZN(n9674)
         );
  INV_X1 U12201 ( .A(n9674), .ZN(n9675) );
  NAND2_X1 U12202 ( .A1(n9676), .A2(n9675), .ZN(n14483) );
  XNOR2_X1 U12203 ( .A(n14674), .B(n14483), .ZN(n14445) );
  INV_X1 U12204 ( .A(n14674), .ZN(n14801) );
  INV_X1 U12205 ( .A(n14483), .ZN(n14191) );
  NAND2_X1 U12206 ( .A1(n14793), .A2(n14666), .ZN(n9739) );
  NAND2_X1 U12207 ( .A1(n12661), .A2(n14407), .ZN(n9679) );
  INV_X1 U12208 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n12663) );
  OR2_X1 U12209 ( .A1(n14408), .A2(n12663), .ZN(n9678) );
  INV_X1 U12210 ( .A(n9681), .ZN(n9680) );
  NAND2_X1 U12211 ( .A1(n9680), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n10398) );
  INV_X1 U12212 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n12654) );
  NAND2_X1 U12213 ( .A1(n9681), .A2(n12654), .ZN(n9682) );
  NAND2_X1 U12214 ( .A1(n10398), .A2(n9682), .ZN(n14641) );
  INV_X1 U12215 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n9685) );
  NAND2_X1 U12216 ( .A1(n14376), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n9684) );
  NAND2_X1 U12217 ( .A1(n14375), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n9683) );
  OAI211_X1 U12218 ( .C1(n14380), .C2(n9685), .A(n9684), .B(n9683), .ZN(n9686)
         );
  INV_X1 U12219 ( .A(n9686), .ZN(n9687) );
  NAND2_X1 U12220 ( .A1(n14369), .A2(n14480), .ZN(n9690) );
  NAND2_X1 U12221 ( .A1(n9690), .A2(n9689), .ZN(n14448) );
  INV_X1 U12222 ( .A(n14448), .ZN(n14636) );
  NAND2_X1 U12223 ( .A1(n14637), .A2(n14636), .ZN(n14635) );
  NAND2_X1 U12224 ( .A1(n14635), .A2(n9690), .ZN(n9699) );
  INV_X1 U12225 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n14880) );
  NOR2_X1 U12226 ( .A1(n14408), .A2(n14880), .ZN(n9691) );
  OR2_X1 U12227 ( .A1(n10398), .A2(n9692), .ZN(n9698) );
  INV_X1 U12228 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n9695) );
  NAND2_X1 U12229 ( .A1(n14376), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n9694) );
  NAND2_X1 U12230 ( .A1(n14375), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n9693) );
  OAI211_X1 U12231 ( .C1(n14380), .C2(n9695), .A(n9694), .B(n9693), .ZN(n9696)
         );
  INV_X1 U12232 ( .A(n9696), .ZN(n9697) );
  XNOR2_X1 U12233 ( .A(n9699), .B(n14449), .ZN(n10390) );
  INV_X1 U12234 ( .A(n14212), .ZN(n9711) );
  NAND2_X1 U12235 ( .A1(n9704), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9705) );
  NAND2_X1 U12236 ( .A1(n9708), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9710) );
  NAND2_X1 U12237 ( .A1(n9711), .A2(n14218), .ZN(n9712) );
  INV_X2 U12238 ( .A(n14218), .ZN(n10727) );
  NAND2_X1 U12239 ( .A1(n9712), .A2(n12646), .ZN(n10388) );
  OR2_X1 U12240 ( .A1(n14412), .A2(n14619), .ZN(n15313) );
  NAND2_X1 U12241 ( .A1(n9714), .A2(n9713), .ZN(n14439) );
  NAND2_X1 U12242 ( .A1(n14309), .A2(n14307), .ZN(n12450) );
  AND2_X1 U12243 ( .A1(n14439), .A2(n12450), .ZN(n9736) );
  NAND2_X1 U12244 ( .A1(n11181), .A2(n10730), .ZN(n14214) );
  NOR2_X1 U12245 ( .A1(n14216), .A2(n14217), .ZN(n11207) );
  NAND2_X1 U12246 ( .A1(n11206), .A2(n11102), .ZN(n9715) );
  NAND2_X1 U12247 ( .A1(n14228), .A2(n6811), .ZN(n9716) );
  NAND2_X1 U12248 ( .A1(n11105), .A2(n9716), .ZN(n11343) );
  OR2_X1 U12249 ( .A1(n14233), .A2(n9718), .ZN(n9717) );
  NAND2_X1 U12250 ( .A1(n11343), .A2(n9717), .ZN(n9720) );
  NAND2_X1 U12251 ( .A1(n14233), .A2(n9718), .ZN(n9719) );
  NAND2_X1 U12252 ( .A1(n9720), .A2(n9719), .ZN(n11466) );
  INV_X1 U12253 ( .A(n14425), .ZN(n11465) );
  NAND2_X1 U12254 ( .A1(n11466), .A2(n11465), .ZN(n9722) );
  NAND2_X1 U12255 ( .A1(n15293), .A2(n11445), .ZN(n9721) );
  NAND2_X1 U12256 ( .A1(n9722), .A2(n9721), .ZN(n11444) );
  NAND2_X1 U12257 ( .A1(n11444), .A2(n14426), .ZN(n9724) );
  NAND2_X1 U12258 ( .A1(n14250), .A2(n11933), .ZN(n9723) );
  INV_X1 U12259 ( .A(n14496), .ZN(n12124) );
  AND2_X1 U12260 ( .A1(n15309), .A2(n12124), .ZN(n9725) );
  OR2_X1 U12261 ( .A1(n15309), .A2(n12124), .ZN(n9726) );
  INV_X1 U12262 ( .A(n14495), .ZN(n12354) );
  OR2_X1 U12263 ( .A1(n14262), .A2(n12354), .ZN(n9727) );
  NAND2_X1 U12264 ( .A1(n14266), .A2(n9729), .ZN(n9730) );
  OR2_X1 U12265 ( .A1(n14279), .A2(n9731), .ZN(n9732) );
  NAND2_X1 U12266 ( .A1(n9733), .A2(n9732), .ZN(n14924) );
  OR2_X1 U12267 ( .A1(n14917), .A2(n14946), .ZN(n9734) );
  NAND2_X1 U12268 ( .A1(n12226), .A2(n14438), .ZN(n9735) );
  INV_X1 U12269 ( .A(n15135), .ZN(n14310) );
  OR2_X1 U12270 ( .A1(n14851), .A2(n14310), .ZN(n14313) );
  NAND2_X1 U12271 ( .A1(n12449), .A2(n14313), .ZN(n12511) );
  INV_X1 U12272 ( .A(n14827), .ZN(n14734) );
  INV_X1 U12273 ( .A(n14820), .ZN(n14718) );
  INV_X1 U12274 ( .A(n14683), .ZN(n9738) );
  NAND2_X1 U12275 ( .A1(n14780), .A2(n14480), .ZN(n9740) );
  XNOR2_X1 U12276 ( .A(n9741), .B(n14449), .ZN(n9746) );
  NAND2_X1 U12277 ( .A1(n9742), .A2(n14209), .ZN(n9744) );
  NAND2_X1 U12278 ( .A1(n9753), .A2(n14213), .ZN(n9743) );
  NAND2_X1 U12279 ( .A1(n9744), .A2(n9743), .ZN(n15160) );
  NAND2_X1 U12280 ( .A1(n9742), .A2(n9753), .ZN(n14413) );
  INV_X1 U12281 ( .A(n14413), .ZN(n9748) );
  INV_X1 U12282 ( .A(n12662), .ZN(n14520) );
  NAND2_X1 U12283 ( .A1(n9748), .A2(n14520), .ZN(n15131) );
  INV_X1 U12284 ( .A(n15131), .ZN(n14762) );
  NOR2_X1 U12285 ( .A1(n9742), .A2(n9753), .ZN(n10703) );
  AND2_X1 U12286 ( .A1(n14387), .A2(n14619), .ZN(n9773) );
  INV_X1 U12287 ( .A(n9773), .ZN(n9747) );
  NAND2_X1 U12288 ( .A1(n10703), .A2(n9747), .ZN(n15334) );
  INV_X1 U12289 ( .A(P1_B_REG_SCAN_IN), .ZN(n9749) );
  NAND2_X1 U12290 ( .A1(n9748), .A2(n12662), .ZN(n14947) );
  INV_X1 U12291 ( .A(n14947), .ZN(n15134) );
  OAI21_X1 U12292 ( .B1(n6676), .B2(n9749), .A(n15134), .ZN(n14626) );
  INV_X1 U12293 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9752) );
  NAND2_X1 U12294 ( .A1(n14375), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n9751) );
  NAND2_X1 U12295 ( .A1(n14376), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n9750) );
  OAI211_X1 U12296 ( .C1(n14380), .C2(n9752), .A(n9751), .B(n9750), .ZN(n14478) );
  INV_X1 U12297 ( .A(n14478), .ZN(n14383) );
  NOR2_X1 U12298 ( .A1(n14626), .A2(n14383), .ZN(n10395) );
  INV_X1 U12299 ( .A(n14279), .ZN(n15181) );
  INV_X1 U12300 ( .A(n14262), .ZN(n15320) );
  INV_X1 U12301 ( .A(n10730), .ZN(n11294) );
  NAND2_X1 U12302 ( .A1(n10815), .A2(n11294), .ZN(n11216) );
  OR2_X1 U12303 ( .A1(n14224), .A2(n11216), .ZN(n11217) );
  INV_X1 U12304 ( .A(n15309), .ZN(n12127) );
  NAND2_X1 U12305 ( .A1(n15112), .A2(n14957), .ZN(n14956) );
  NAND2_X1 U12306 ( .A1(n14323), .A2(n12514), .ZN(n14757) );
  INV_X1 U12307 ( .A(n15122), .ZN(n14741) );
  AOI211_X1 U12308 ( .C1(n14393), .C2(n14639), .A(n14741), .B(n14630), .ZN(
        n10400) );
  AOI211_X1 U12309 ( .C1(n15310), .C2(n14393), .A(n10395), .B(n10400), .ZN(
        n9754) );
  NOR2_X1 U12310 ( .A1(n9575), .A2(n9755), .ZN(n9759) );
  INV_X1 U12311 ( .A(n9759), .ZN(n9756) );
  NAND2_X1 U12312 ( .A1(n9756), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9757) );
  MUX2_X1 U12313 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9757), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n9760) );
  NAND2_X1 U12314 ( .A1(n9759), .A2(n9758), .ZN(n9763) );
  NAND2_X1 U12315 ( .A1(n9760), .A2(n9763), .ZN(n12380) );
  NAND2_X1 U12316 ( .A1(n12380), .A2(P1_B_REG_SCAN_IN), .ZN(n9762) );
  MUX2_X1 U12317 ( .A(n9762), .B(P1_B_REG_SCAN_IN), .S(n12328), .Z(n9766) );
  NAND2_X1 U12318 ( .A1(n9763), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9765) );
  XNOR2_X1 U12319 ( .A(n9765), .B(n9764), .ZN(n14888) );
  INV_X1 U12320 ( .A(n14888), .ZN(n9767) );
  OR2_X1 U12321 ( .A1(n10474), .A2(P1_D_REG_0__SCAN_IN), .ZN(n9768) );
  OR2_X1 U12322 ( .A1(n12328), .A2(n9767), .ZN(n10477) );
  AND2_X1 U12323 ( .A1(n9768), .A2(n10477), .ZN(n11096) );
  NOR2_X1 U12324 ( .A1(n14888), .A2(n12380), .ZN(n9769) );
  NAND2_X2 U12325 ( .A1(n12328), .A2(n9769), .ZN(n10734) );
  NAND2_X1 U12326 ( .A1(n9770), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9772) );
  INV_X1 U12327 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n9771) );
  XNOR2_X1 U12328 ( .A(n9772), .B(n9771), .ZN(n10482) );
  OAI211_X1 U12329 ( .C1(n9773), .C2(n14413), .A(n10734), .B(n10482), .ZN(
        n10721) );
  NOR2_X1 U12330 ( .A1(n11096), .A2(n14472), .ZN(n9786) );
  AND2_X1 U12331 ( .A1(n12380), .A2(n14888), .ZN(n10475) );
  INV_X1 U12332 ( .A(n10475), .ZN(n9774) );
  OAI21_X1 U12333 ( .B1(n10474), .B2(P1_D_REG_1__SCAN_IN), .A(n9774), .ZN(
        n9785) );
  NAND2_X1 U12334 ( .A1(n15122), .A2(n14209), .ZN(n10720) );
  NOR4_X1 U12335 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n9783) );
  NOR4_X1 U12336 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n9782) );
  OR4_X1 U12337 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n9780) );
  NOR4_X1 U12338 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n9778) );
  NOR4_X1 U12339 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n9777) );
  NOR4_X1 U12340 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n9776) );
  NOR4_X1 U12341 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n9775) );
  NAND4_X1 U12342 ( .A1(n9778), .A2(n9777), .A3(n9776), .A4(n9775), .ZN(n9779)
         );
  NOR4_X1 U12343 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n9780), .A4(n9779), .ZN(n9781) );
  AND3_X1 U12344 ( .A1(n9783), .A2(n9782), .A3(n9781), .ZN(n10383) );
  OR2_X1 U12345 ( .A1(n10474), .A2(n10383), .ZN(n9784) );
  NAND2_X1 U12346 ( .A1(n14776), .A2(n15341), .ZN(n9788) );
  XNOR2_X1 U12347 ( .A(n10362), .B(n9870), .ZN(n12676) );
  NOR2_X1 U12348 ( .A1(n12676), .A2(n13112), .ZN(n12671) );
  AOI21_X1 U12349 ( .B1(n12676), .B2(n13112), .A(n12671), .ZN(n9874) );
  INV_X4 U12350 ( .A(n9870), .ZN(n12669) );
  XNOR2_X1 U12351 ( .A(n13240), .B(n12669), .ZN(n9845) );
  INV_X1 U12352 ( .A(n12845), .ZN(n9792) );
  AND3_X1 U12353 ( .A1(n15682), .A2(n9870), .A3(n9796), .ZN(n9797) );
  NAND2_X1 U12354 ( .A1(n15701), .A2(n9870), .ZN(n9798) );
  NAND2_X1 U12355 ( .A1(n9799), .A2(n9798), .ZN(n9800) );
  XNOR2_X1 U12356 ( .A(n9870), .B(n15687), .ZN(n9802) );
  XNOR2_X1 U12357 ( .A(n9802), .B(n15698), .ZN(n11171) );
  INV_X1 U12358 ( .A(n9802), .ZN(n9803) );
  NOR2_X1 U12359 ( .A1(n9803), .A2(n15698), .ZN(n9804) );
  XNOR2_X1 U12360 ( .A(n9805), .B(n15681), .ZN(n11239) );
  INV_X1 U12361 ( .A(n9805), .ZN(n9806) );
  NAND2_X1 U12362 ( .A1(n9806), .A2(n15681), .ZN(n9807) );
  XNOR2_X1 U12363 ( .A(n11569), .B(n7125), .ZN(n9808) );
  XNOR2_X1 U12364 ( .A(n9808), .B(n11673), .ZN(n11537) );
  OR2_X1 U12365 ( .A1(n11673), .A2(n9808), .ZN(n9809) );
  XNOR2_X1 U12366 ( .A(n9870), .B(n11682), .ZN(n9810) );
  XNOR2_X1 U12367 ( .A(n9810), .B(n12995), .ZN(n11652) );
  INV_X1 U12368 ( .A(n9810), .ZN(n9811) );
  OR2_X1 U12369 ( .A1(n12995), .A2(n9811), .ZN(n9812) );
  XNOR2_X1 U12370 ( .A(n9870), .B(n15664), .ZN(n9814) );
  XNOR2_X1 U12371 ( .A(n9814), .B(n11947), .ZN(n11697) );
  NAND2_X1 U12372 ( .A1(n9814), .A2(n11947), .ZN(n11815) );
  NAND2_X1 U12373 ( .A1(n9815), .A2(n12031), .ZN(n9816) );
  AND2_X1 U12374 ( .A1(n11817), .A2(n9816), .ZN(n9817) );
  XNOR2_X1 U12375 ( .A(n11834), .B(n12669), .ZN(n9818) );
  XNOR2_X1 U12376 ( .A(n9818), .B(n12189), .ZN(n11831) );
  INV_X1 U12377 ( .A(n9818), .ZN(n9819) );
  NAND2_X1 U12378 ( .A1(n9819), .A2(n12189), .ZN(n9820) );
  XNOR2_X1 U12379 ( .A(n15731), .B(n12669), .ZN(n9822) );
  XNOR2_X1 U12380 ( .A(n9822), .B(n15639), .ZN(n12047) );
  XNOR2_X1 U12381 ( .A(n15647), .B(n12669), .ZN(n9821) );
  AND2_X1 U12382 ( .A1(n9821), .A2(n15043), .ZN(n9825) );
  OR2_X1 U12383 ( .A1(n12047), .A2(n9825), .ZN(n9829) );
  XNOR2_X1 U12384 ( .A(n15051), .B(n12669), .ZN(n9832) );
  INV_X1 U12385 ( .A(n9832), .ZN(n9827) );
  XNOR2_X1 U12386 ( .A(n9821), .B(n15043), .ZN(n12095) );
  INV_X1 U12387 ( .A(n12095), .ZN(n9824) );
  INV_X1 U12388 ( .A(n15639), .ZN(n12103) );
  INV_X1 U12389 ( .A(n9822), .ZN(n9823) );
  NAND2_X1 U12390 ( .A1(n12103), .A2(n9823), .ZN(n12094) );
  AND2_X1 U12391 ( .A1(n9824), .A2(n12094), .ZN(n12097) );
  OR2_X1 U12392 ( .A1(n9825), .A2(n12097), .ZN(n9831) );
  OR2_X1 U12393 ( .A1(n9829), .A2(n9832), .ZN(n9830) );
  OR2_X1 U12394 ( .A1(n9832), .A2(n9831), .ZN(n9833) );
  XNOR2_X1 U12395 ( .A(n15069), .B(n12669), .ZN(n9834) );
  XOR2_X1 U12396 ( .A(n15042), .B(n9834), .Z(n12219) );
  INV_X1 U12397 ( .A(n9834), .ZN(n9835) );
  XOR2_X1 U12398 ( .A(n12669), .B(n12364), .Z(n12280) );
  NOR2_X1 U12399 ( .A1(n12280), .A2(n13292), .ZN(n9837) );
  INV_X1 U12400 ( .A(n12280), .ZN(n9836) );
  XNOR2_X1 U12401 ( .A(n13423), .B(n12669), .ZN(n9838) );
  XOR2_X1 U12402 ( .A(n12438), .B(n9838), .Z(n12331) );
  XNOR2_X1 U12403 ( .A(n13282), .B(n9870), .ZN(n9839) );
  NAND2_X1 U12404 ( .A1(n9839), .A2(n13291), .ZN(n12435) );
  INV_X1 U12405 ( .A(n12732), .ZN(n9842) );
  XOR2_X1 U12406 ( .A(n12669), .B(n13266), .Z(n12730) );
  INV_X1 U12407 ( .A(n12730), .ZN(n9841) );
  XNOR2_X1 U12408 ( .A(n13251), .B(n12669), .ZN(n9843) );
  XOR2_X1 U12409 ( .A(n13234), .B(n9843), .Z(n12741) );
  AND2_X1 U12410 ( .A1(n9843), .A2(n13263), .ZN(n9844) );
  XNOR2_X1 U12411 ( .A(n9845), .B(n13219), .ZN(n12780) );
  XNOR2_X1 U12412 ( .A(n13225), .B(n12669), .ZN(n9846) );
  XNOR2_X1 U12413 ( .A(n9846), .B(n13235), .ZN(n12701) );
  INV_X1 U12414 ( .A(n9846), .ZN(n9847) );
  XNOR2_X1 U12415 ( .A(n13402), .B(n12669), .ZN(n9850) );
  XNOR2_X1 U12416 ( .A(n9850), .B(n6674), .ZN(n12761) );
  INV_X1 U12417 ( .A(n9850), .ZN(n9851) );
  NAND2_X1 U12418 ( .A1(n9851), .A2(n6673), .ZN(n9852) );
  XNOR2_X1 U12419 ( .A(n12708), .B(n12669), .ZN(n9853) );
  XNOR2_X1 U12420 ( .A(n9853), .B(n13208), .ZN(n12709) );
  INV_X1 U12421 ( .A(n9853), .ZN(n9854) );
  NAND2_X1 U12422 ( .A1(n9854), .A2(n12771), .ZN(n9855) );
  INV_X1 U12423 ( .A(n9857), .ZN(n9859) );
  XOR2_X1 U12424 ( .A(n12669), .B(n13181), .Z(n9856) );
  INV_X1 U12425 ( .A(n9856), .ZN(n9858) );
  NAND2_X1 U12426 ( .A1(n12767), .A2(n9860), .ZN(n9862) );
  XNOR2_X1 U12427 ( .A(n13163), .B(n12669), .ZN(n9861) );
  NAND2_X1 U12428 ( .A1(n12694), .A2(n12747), .ZN(n9866) );
  XNOR2_X1 U12429 ( .A(n13325), .B(n9870), .ZN(n9863) );
  NAND2_X1 U12430 ( .A1(n9863), .A2(n12726), .ZN(n12720) );
  INV_X1 U12431 ( .A(n9863), .ZN(n9864) );
  NAND2_X1 U12432 ( .A1(n9864), .A2(n13160), .ZN(n9865) );
  XNOR2_X1 U12433 ( .A(n13134), .B(n12669), .ZN(n9867) );
  NAND2_X1 U12434 ( .A1(n9867), .A2(n13149), .ZN(n12718) );
  AND2_X1 U12435 ( .A1(n12720), .A2(n12718), .ZN(n9869) );
  INV_X1 U12436 ( .A(n9867), .ZN(n9868) );
  INV_X1 U12437 ( .A(n13149), .ZN(n11632) );
  NAND2_X1 U12438 ( .A1(n9868), .A2(n11632), .ZN(n12717) );
  XNOR2_X1 U12439 ( .A(n13118), .B(n9870), .ZN(n9871) );
  NOR2_X1 U12440 ( .A1(n9871), .A2(n13127), .ZN(n9872) );
  AOI21_X1 U12441 ( .B1(n9871), .B2(n13127), .A(n9872), .ZN(n12787) );
  OAI21_X1 U12442 ( .B1(n9874), .B2(n9873), .A(n12682), .ZN(n9876) );
  OAI22_X1 U12443 ( .A1(n10898), .A2(n9882), .B1(n9887), .B2(n9880), .ZN(n9875) );
  NAND2_X1 U12444 ( .A1(n9876), .A2(n12788), .ZN(n9899) );
  NAND2_X1 U12445 ( .A1(n10907), .A2(n15070), .ZN(n11362) );
  AND2_X1 U12446 ( .A1(n9882), .A2(n15708), .ZN(n9877) );
  NOR2_X1 U12447 ( .A1(n13278), .A2(n9880), .ZN(n9878) );
  AND2_X1 U12448 ( .A1(n9879), .A2(n15700), .ZN(n12988) );
  NAND2_X1 U12449 ( .A1(n12988), .A2(n9888), .ZN(n12792) );
  NAND2_X1 U12450 ( .A1(n9881), .A2(n9880), .ZN(n9891) );
  NAND2_X1 U12451 ( .A1(n9883), .A2(n9882), .ZN(n9886) );
  AND3_X1 U12452 ( .A1(n9884), .A2(n10408), .A3(n10910), .ZN(n9885) );
  OAI211_X1 U12453 ( .C1(n9888), .C2(n9887), .A(n9886), .B(n9885), .ZN(n9889)
         );
  NAND2_X1 U12454 ( .A1(n9889), .A2(P3_STATE_REG_SCAN_IN), .ZN(n9890) );
  AOI22_X1 U12455 ( .A1(n13102), .A2(n12790), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n9892) );
  OAI21_X1 U12456 ( .B1(n9893), .B2(n12792), .A(n9892), .ZN(n9894) );
  AOI21_X1 U12457 ( .B1(n12794), .B2(n11923), .A(n9894), .ZN(n9895) );
  NAND2_X1 U12458 ( .A1(n9899), .A2(n9898), .ZN(P3_U3154) );
  INV_X1 U12459 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n15015) );
  INV_X1 U12460 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n9925) );
  INV_X1 U12461 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n11250) );
  XNOR2_X1 U12462 ( .A(P3_ADDR_REG_14__SCAN_IN), .B(n11250), .ZN(n9935) );
  INV_X1 U12463 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n15256) );
  INV_X1 U12464 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n10613) );
  INV_X1 U12465 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n9918) );
  INV_X1 U12466 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n14574) );
  INV_X1 U12467 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n9911) );
  NOR2_X1 U12468 ( .A1(n9902), .A2(n10195), .ZN(n9903) );
  NOR2_X1 U12469 ( .A1(n9905), .A2(n10222), .ZN(n9906) );
  INV_X1 U12470 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n15239) );
  NOR2_X1 U12471 ( .A1(n9907), .A2(n10212), .ZN(n9909) );
  INV_X1 U12472 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n14555) );
  INV_X1 U12473 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n10226) );
  XNOR2_X1 U12474 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(n10226), .ZN(n9961) );
  INV_X1 U12475 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n9913) );
  NOR2_X1 U12476 ( .A1(n9912), .A2(n9913), .ZN(n9915) );
  INV_X1 U12477 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n10040) );
  XNOR2_X1 U12478 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n10040), .ZN(n9940) );
  XNOR2_X1 U12479 ( .A(n9918), .B(P3_ADDR_REG_9__SCAN_IN), .ZN(n9938) );
  NOR2_X1 U12480 ( .A1(n9939), .A2(n9938), .ZN(n9917) );
  AOI21_X1 U12481 ( .B1(P3_ADDR_REG_9__SCAN_IN), .B2(n9918), .A(n9917), .ZN(
        n9919) );
  AND2_X1 U12482 ( .A1(n9919), .A2(P1_ADDR_REG_10__SCAN_IN), .ZN(n9975) );
  NOR2_X1 U12483 ( .A1(n9919), .A2(P1_ADDR_REG_10__SCAN_IN), .ZN(n9974) );
  NOR2_X1 U12484 ( .A1(P3_ADDR_REG_10__SCAN_IN), .A2(n9974), .ZN(n9920) );
  XNOR2_X1 U12485 ( .A(n10613), .B(P3_ADDR_REG_11__SCAN_IN), .ZN(n9936) );
  AOI21_X2 U12486 ( .B1(P3_ADDR_REG_11__SCAN_IN), .B2(n10613), .A(n9921), .ZN(
        n9978) );
  XNOR2_X1 U12487 ( .A(n15256), .B(P3_ADDR_REG_12__SCAN_IN), .ZN(n9977) );
  INV_X1 U12488 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n9979) );
  AND2_X1 U12489 ( .A1(n9979), .A2(P1_ADDR_REG_13__SCAN_IN), .ZN(n9923) );
  INV_X1 U12490 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n9931) );
  NAND2_X1 U12491 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(n9931), .ZN(n9926) );
  NOR2_X1 U12492 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(n9931), .ZN(n9930) );
  NAND2_X1 U12493 ( .A1(n9927), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n9929) );
  XOR2_X1 U12494 ( .A(P1_ADDR_REG_16__SCAN_IN), .B(n9927), .Z(n9984) );
  INV_X1 U12495 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n14994) );
  NAND2_X1 U12496 ( .A1(n9984), .A2(n14994), .ZN(n9928) );
  NAND2_X1 U12497 ( .A1(n9929), .A2(n9928), .ZN(n9987) );
  XNOR2_X1 U12498 ( .A(P1_ADDR_REG_17__SCAN_IN), .B(n9987), .ZN(n9988) );
  XOR2_X1 U12499 ( .A(n15015), .B(n9988), .Z(n14965) );
  AOI21_X1 U12500 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(n9931), .A(n9930), .ZN(
        n9933) );
  XOR2_X1 U12501 ( .A(n9933), .B(n9932), .Z(n15215) );
  XNOR2_X1 U12502 ( .A(n9935), .B(n9934), .ZN(n15211) );
  XOR2_X1 U12503 ( .A(n9937), .B(n9936), .Z(n15198) );
  XOR2_X1 U12504 ( .A(n9939), .B(n9938), .Z(n9972) );
  INV_X1 U12505 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n9944) );
  NAND2_X1 U12506 ( .A1(n9945), .A2(n9944), .ZN(n9957) );
  XOR2_X1 U12507 ( .A(n9946), .B(P1_ADDR_REG_3__SCAN_IN), .Z(n15764) );
  XOR2_X1 U12508 ( .A(n9948), .B(n9947), .Z(n14901) );
  INV_X1 U12509 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n9950) );
  NOR2_X1 U12510 ( .A1(n9953), .A2(n9950), .ZN(n9954) );
  OAI21_X1 U12511 ( .B1(P3_ADDR_REG_0__SCAN_IN), .B2(n9952), .A(n9951), .ZN(
        n15758) );
  NAND2_X1 U12512 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(n15758), .ZN(n15768) );
  NOR2_X1 U12513 ( .A1(n15768), .A2(n15767), .ZN(n15766) );
  NOR2_X1 U12514 ( .A1(n14901), .A2(n14900), .ZN(n9955) );
  NAND2_X1 U12515 ( .A1(n14901), .A2(n14900), .ZN(n14899) );
  OAI21_X1 U12516 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(n9955), .A(n14899), .ZN(
        n15763) );
  NAND2_X1 U12517 ( .A1(n15764), .A2(n15763), .ZN(n9956) );
  NOR2_X1 U12518 ( .A1(n15764), .A2(n15763), .ZN(n15762) );
  AOI21_X1 U12519 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(n9956), .A(n15762), .ZN(
        n15754) );
  NAND2_X1 U12520 ( .A1(n9958), .A2(n9959), .ZN(n9960) );
  INV_X1 U12521 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n15756) );
  NOR2_X1 U12522 ( .A1(n9963), .A2(n7231), .ZN(n9964) );
  XOR2_X1 U12523 ( .A(n9962), .B(n9961), .Z(n14905) );
  INV_X1 U12524 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n9965) );
  NAND2_X1 U12525 ( .A1(n9967), .A2(n9965), .ZN(n9968) );
  XOR2_X1 U12526 ( .A(n9966), .B(P1_ADDR_REG_7__SCAN_IN), .Z(n15761) );
  NAND2_X1 U12527 ( .A1(n9969), .A2(n9970), .ZN(n9971) );
  INV_X1 U12528 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n14907) );
  INV_X1 U12529 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n14910) );
  INV_X1 U12530 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n11863) );
  NOR2_X1 U12531 ( .A1(n9975), .A2(n9974), .ZN(n9976) );
  XNOR2_X1 U12532 ( .A(n11863), .B(n9976), .ZN(n14913) );
  XOR2_X1 U12533 ( .A(n9978), .B(n9977), .Z(n15201) );
  XNOR2_X1 U12534 ( .A(P1_ADDR_REG_13__SCAN_IN), .B(n9979), .ZN(n9980) );
  XNOR2_X1 U12535 ( .A(n9981), .B(n9980), .ZN(n9982) );
  INV_X1 U12536 ( .A(n15205), .ZN(n15206) );
  INV_X1 U12537 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n15208) );
  NAND2_X1 U12538 ( .A1(n9983), .A2(n9982), .ZN(n15207) );
  XOR2_X1 U12539 ( .A(P3_ADDR_REG_16__SCAN_IN), .B(n9984), .Z(n15218) );
  NAND2_X1 U12540 ( .A1(n15219), .A2(n15218), .ZN(n9985) );
  NAND2_X1 U12541 ( .A1(n14965), .A2(n14964), .ZN(n9986) );
  NOR2_X1 U12542 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n9987), .ZN(n9990) );
  NOR2_X1 U12543 ( .A1(n15015), .A2(n9988), .ZN(n9989) );
  NOR2_X1 U12544 ( .A1(n9990), .A2(n9989), .ZN(n9994) );
  XOR2_X1 U12545 ( .A(P3_ADDR_REG_18__SCAN_IN), .B(P1_ADDR_REG_18__SCAN_IN), 
        .Z(n9993) );
  XOR2_X1 U12546 ( .A(n9994), .B(n9993), .Z(n14895) );
  XNOR2_X1 U12547 ( .A(P3_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n9991) );
  XNOR2_X1 U12548 ( .A(n9991), .B(n7717), .ZN(n9992) );
  INV_X1 U12549 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n15271) );
  NOR2_X1 U12550 ( .A1(n9994), .A2(n9993), .ZN(n9995) );
  AOI21_X1 U12551 ( .B1(P3_ADDR_REG_18__SCAN_IN), .B2(n15271), .A(n9995), .ZN(
        n10339) );
  OAI22_X1 U12552 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(keyinput_g121), .B1(
        keyinput_g67), .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n9996) );
  AOI221_X1 U12553 ( .B1(P1_IR_REG_14__SCAN_IN), .B2(keyinput_g121), .C1(
        P3_DATAO_REG_29__SCAN_IN), .C2(keyinput_g67), .A(n9996), .ZN(n10003)
         );
  OAI22_X1 U12554 ( .A1(P3_DATAO_REG_15__SCAN_IN), .A2(keyinput_g81), .B1(
        keyinput_g79), .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n9997) );
  AOI221_X1 U12555 ( .B1(P3_DATAO_REG_15__SCAN_IN), .B2(keyinput_g81), .C1(
        P3_DATAO_REG_17__SCAN_IN), .C2(keyinput_g79), .A(n9997), .ZN(n10002)
         );
  OAI22_X1 U12556 ( .A1(n10312), .A2(keyinput_g114), .B1(keyinput_g106), .B2(
        P3_ADDR_REG_9__SCAN_IN), .ZN(n9998) );
  AOI221_X1 U12557 ( .B1(n10312), .B2(keyinput_g114), .C1(
        P3_ADDR_REG_9__SCAN_IN), .C2(keyinput_g106), .A(n9998), .ZN(n10001) );
  OAI22_X1 U12558 ( .A1(SI_10_), .A2(keyinput_g22), .B1(
        P3_DATAO_REG_5__SCAN_IN), .B2(keyinput_g91), .ZN(n9999) );
  AOI221_X1 U12559 ( .B1(SI_10_), .B2(keyinput_g22), .C1(keyinput_g91), .C2(
        P3_DATAO_REG_5__SCAN_IN), .A(n9999), .ZN(n10000) );
  NAND4_X1 U12560 ( .A1(n10003), .A2(n10002), .A3(n10001), .A4(n10000), .ZN(
        n10117) );
  OAI22_X1 U12561 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(keyinput_g40), .B1(
        keyinput_g118), .B2(P1_IR_REG_11__SCAN_IN), .ZN(n10004) );
  AOI221_X1 U12562 ( .B1(P3_REG3_REG_3__SCAN_IN), .B2(keyinput_g40), .C1(
        P1_IR_REG_11__SCAN_IN), .C2(keyinput_g118), .A(n10004), .ZN(n10029) );
  INV_X1 U12563 ( .A(P3_B_REG_SCAN_IN), .ZN(n10373) );
  OAI22_X1 U12564 ( .A1(SI_19_), .A2(keyinput_g13), .B1(P3_ADDR_REG_4__SCAN_IN), .B2(keyinput_g101), .ZN(n10005) );
  AOI221_X1 U12565 ( .B1(SI_19_), .B2(keyinput_g13), .C1(keyinput_g101), .C2(
        P3_ADDR_REG_4__SCAN_IN), .A(n10005), .ZN(n10008) );
  OAI22_X1 U12566 ( .A1(P3_REG3_REG_6__SCAN_IN), .A2(keyinput_g61), .B1(
        keyinput_g123), .B2(P1_IR_REG_16__SCAN_IN), .ZN(n10006) );
  AOI221_X1 U12567 ( .B1(P3_REG3_REG_6__SCAN_IN), .B2(keyinput_g61), .C1(
        P1_IR_REG_16__SCAN_IN), .C2(keyinput_g123), .A(n10006), .ZN(n10007) );
  OAI211_X1 U12568 ( .C1(n10373), .C2(keyinput_g64), .A(n10008), .B(n10007), 
        .ZN(n10009) );
  AOI21_X1 U12569 ( .B1(n10373), .B2(keyinput_g64), .A(n10009), .ZN(n10028) );
  AOI22_X1 U12570 ( .A1(P3_DATAO_REG_20__SCAN_IN), .A2(keyinput_g76), .B1(
        P3_REG3_REG_12__SCAN_IN), .B2(keyinput_g46), .ZN(n10010) );
  OAI221_X1 U12571 ( .B1(P3_DATAO_REG_20__SCAN_IN), .B2(keyinput_g76), .C1(
        P3_REG3_REG_12__SCAN_IN), .C2(keyinput_g46), .A(n10010), .ZN(n10017)
         );
  AOI22_X1 U12572 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(keyinput_g116), .B1(
        P3_REG3_REG_14__SCAN_IN), .B2(keyinput_g37), .ZN(n10011) );
  OAI221_X1 U12573 ( .B1(P1_IR_REG_9__SCAN_IN), .B2(keyinput_g116), .C1(
        P3_REG3_REG_14__SCAN_IN), .C2(keyinput_g37), .A(n10011), .ZN(n10016)
         );
  AOI22_X1 U12574 ( .A1(P3_REG3_REG_1__SCAN_IN), .A2(keyinput_g44), .B1(
        P3_REG3_REG_11__SCAN_IN), .B2(keyinput_g58), .ZN(n10012) );
  OAI221_X1 U12575 ( .B1(P3_REG3_REG_1__SCAN_IN), .B2(keyinput_g44), .C1(
        P3_REG3_REG_11__SCAN_IN), .C2(keyinput_g58), .A(n10012), .ZN(n10015)
         );
  AOI22_X1 U12576 ( .A1(P3_DATAO_REG_21__SCAN_IN), .A2(keyinput_g75), .B1(
        SI_7_), .B2(keyinput_g25), .ZN(n10013) );
  OAI221_X1 U12577 ( .B1(P3_DATAO_REG_21__SCAN_IN), .B2(keyinput_g75), .C1(
        SI_7_), .C2(keyinput_g25), .A(n10013), .ZN(n10014) );
  NOR4_X1 U12578 ( .A1(n10017), .A2(n10016), .A3(n10015), .A4(n10014), .ZN(
        n10027) );
  AOI22_X1 U12579 ( .A1(P3_ADDR_REG_3__SCAN_IN), .A2(keyinput_g100), .B1(SI_4_), .B2(keyinput_g28), .ZN(n10018) );
  OAI221_X1 U12580 ( .B1(P3_ADDR_REG_3__SCAN_IN), .B2(keyinput_g100), .C1(
        SI_4_), .C2(keyinput_g28), .A(n10018), .ZN(n10025) );
  AOI22_X1 U12581 ( .A1(P3_DATAO_REG_31__SCAN_IN), .A2(keyinput_g65), .B1(
        SI_16_), .B2(keyinput_g16), .ZN(n10019) );
  OAI221_X1 U12582 ( .B1(P3_DATAO_REG_31__SCAN_IN), .B2(keyinput_g65), .C1(
        SI_16_), .C2(keyinput_g16), .A(n10019), .ZN(n10024) );
  AOI22_X1 U12583 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(keyinput_g111), .B1(
        P1_IR_REG_17__SCAN_IN), .B2(keyinput_g124), .ZN(n10020) );
  OAI221_X1 U12584 ( .B1(P1_IR_REG_4__SCAN_IN), .B2(keyinput_g111), .C1(
        P1_IR_REG_17__SCAN_IN), .C2(keyinput_g124), .A(n10020), .ZN(n10023) );
  AOI22_X1 U12585 ( .A1(P3_ADDR_REG_7__SCAN_IN), .A2(keyinput_g104), .B1(
        SI_12_), .B2(keyinput_g20), .ZN(n10021) );
  OAI221_X1 U12586 ( .B1(P3_ADDR_REG_7__SCAN_IN), .B2(keyinput_g104), .C1(
        SI_12_), .C2(keyinput_g20), .A(n10021), .ZN(n10022) );
  NOR4_X1 U12587 ( .A1(n10025), .A2(n10024), .A3(n10023), .A4(n10022), .ZN(
        n10026) );
  NAND4_X1 U12588 ( .A1(n10029), .A2(n10028), .A3(n10027), .A4(n10026), .ZN(
        n10116) );
  AOI22_X1 U12589 ( .A1(P3_DATAO_REG_4__SCAN_IN), .A2(keyinput_g92), .B1(
        P3_RD_REG_SCAN_IN), .B2(keyinput_g33), .ZN(n10030) );
  OAI221_X1 U12590 ( .B1(P3_DATAO_REG_4__SCAN_IN), .B2(keyinput_g92), .C1(
        P3_RD_REG_SCAN_IN), .C2(keyinput_g33), .A(n10030), .ZN(n10038) );
  AOI22_X1 U12591 ( .A1(P3_DATAO_REG_10__SCAN_IN), .A2(keyinput_g86), .B1(
        SI_29_), .B2(keyinput_g3), .ZN(n10031) );
  OAI221_X1 U12592 ( .B1(P3_DATAO_REG_10__SCAN_IN), .B2(keyinput_g86), .C1(
        SI_29_), .C2(keyinput_g3), .A(n10031), .ZN(n10037) );
  AOI22_X1 U12593 ( .A1(P3_DATAO_REG_26__SCAN_IN), .A2(keyinput_g70), .B1(
        P3_DATAO_REG_3__SCAN_IN), .B2(keyinput_g93), .ZN(n10032) );
  OAI221_X1 U12594 ( .B1(P3_DATAO_REG_26__SCAN_IN), .B2(keyinput_g70), .C1(
        P3_DATAO_REG_3__SCAN_IN), .C2(keyinput_g93), .A(n10032), .ZN(n10036)
         );
  XNOR2_X1 U12595 ( .A(P1_IR_REG_12__SCAN_IN), .B(keyinput_g119), .ZN(n10034)
         );
  XNOR2_X1 U12596 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput_g110), .ZN(n10033)
         );
  NAND2_X1 U12597 ( .A1(n10034), .A2(n10033), .ZN(n10035) );
  NOR4_X1 U12598 ( .A1(n10038), .A2(n10037), .A3(n10036), .A4(n10035), .ZN(
        n10072) );
  INV_X1 U12599 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n15549) );
  AOI22_X1 U12600 ( .A1(n15549), .A2(keyinput_g97), .B1(n10040), .B2(
        keyinput_g105), .ZN(n10039) );
  OAI221_X1 U12601 ( .B1(n15549), .B2(keyinput_g97), .C1(n10040), .C2(
        keyinput_g105), .A(n10039), .ZN(n10048) );
  INV_X1 U12602 ( .A(P3_DATAO_REG_6__SCAN_IN), .ZN(n10666) );
  XNOR2_X1 U12603 ( .A(n10666), .B(keyinput_g90), .ZN(n10047) );
  INV_X1 U12604 ( .A(P3_DATAO_REG_12__SCAN_IN), .ZN(n10662) );
  XNOR2_X1 U12605 ( .A(n10662), .B(keyinput_g84), .ZN(n10046) );
  XNOR2_X1 U12606 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput_g112), .ZN(n10044)
         );
  XNOR2_X1 U12607 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput_g108), .ZN(n10043)
         );
  XNOR2_X1 U12608 ( .A(SI_1_), .B(keyinput_g31), .ZN(n10042) );
  XNOR2_X1 U12609 ( .A(SI_8_), .B(keyinput_g24), .ZN(n10041) );
  NAND4_X1 U12610 ( .A1(n10044), .A2(n10043), .A3(n10042), .A4(n10041), .ZN(
        n10045) );
  NOR4_X1 U12611 ( .A1(n10048), .A2(n10047), .A3(n10046), .A4(n10045), .ZN(
        n10071) );
  INV_X1 U12612 ( .A(P3_DATAO_REG_27__SCAN_IN), .ZN(n11802) );
  AOI22_X1 U12613 ( .A1(n10050), .A2(keyinput_g120), .B1(keyinput_g69), .B2(
        n11802), .ZN(n10049) );
  OAI221_X1 U12614 ( .B1(n10050), .B2(keyinput_g120), .C1(n11802), .C2(
        keyinput_g69), .A(n10049), .ZN(n10055) );
  AOI22_X1 U12615 ( .A1(n10052), .A2(keyinput_g115), .B1(n10223), .B2(
        keyinput_g45), .ZN(n10051) );
  OAI221_X1 U12616 ( .B1(n10052), .B2(keyinput_g115), .C1(n10223), .C2(
        keyinput_g45), .A(n10051), .ZN(n10054) );
  XOR2_X1 U12617 ( .A(SI_5_), .B(keyinput_g27), .Z(n10053) );
  OR3_X1 U12618 ( .A1(n10055), .A2(n10054), .A3(n10053), .ZN(n10059) );
  INV_X1 U12619 ( .A(P3_DATAO_REG_13__SCAN_IN), .ZN(n10672) );
  AOI22_X1 U12620 ( .A1(n12668), .A2(keyinput_g4), .B1(keyinput_g83), .B2(
        n10672), .ZN(n10056) );
  OAI221_X1 U12621 ( .B1(n12668), .B2(keyinput_g4), .C1(n10672), .C2(
        keyinput_g83), .A(n10056), .ZN(n10058) );
  INV_X1 U12622 ( .A(P3_DATAO_REG_16__SCAN_IN), .ZN(n10677) );
  XNOR2_X1 U12623 ( .A(n10677), .B(keyinput_g80), .ZN(n10057) );
  NOR3_X1 U12624 ( .A1(n10059), .A2(n10058), .A3(n10057), .ZN(n10070) );
  AOI22_X1 U12625 ( .A1(n11333), .A2(keyinput_g43), .B1(keyinput_g54), .B2(
        n11364), .ZN(n10060) );
  OAI221_X1 U12626 ( .B1(n11333), .B2(keyinput_g43), .C1(n11364), .C2(
        keyinput_g54), .A(n10060), .ZN(n10063) );
  XOR2_X1 U12627 ( .A(P1_IR_REG_0__SCAN_IN), .B(keyinput_g107), .Z(n10062) );
  INV_X1 U12628 ( .A(P3_DATAO_REG_9__SCAN_IN), .ZN(n10660) );
  XNOR2_X1 U12629 ( .A(n10660), .B(keyinput_g87), .ZN(n10061) );
  OR3_X1 U12630 ( .A1(n10063), .A2(n10062), .A3(n10061), .ZN(n10068) );
  INV_X1 U12631 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n10940) );
  INV_X1 U12632 ( .A(P3_ADDR_REG_1__SCAN_IN), .ZN(n10289) );
  AOI22_X1 U12633 ( .A1(n10940), .A2(keyinput_g52), .B1(keyinput_g98), .B2(
        n10289), .ZN(n10064) );
  OAI221_X1 U12634 ( .B1(n10940), .B2(keyinput_g52), .C1(n10289), .C2(
        keyinput_g98), .A(n10064), .ZN(n10067) );
  INV_X1 U12635 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n11862) );
  INV_X1 U12636 ( .A(P3_DATAO_REG_19__SCAN_IN), .ZN(n10709) );
  AOI22_X1 U12637 ( .A1(n11862), .A2(keyinput_g39), .B1(keyinput_g77), .B2(
        n10709), .ZN(n10065) );
  OAI221_X1 U12638 ( .B1(n11862), .B2(keyinput_g39), .C1(n10709), .C2(
        keyinput_g77), .A(n10065), .ZN(n10066) );
  NOR3_X1 U12639 ( .A1(n10068), .A2(n10067), .A3(n10066), .ZN(n10069) );
  NAND4_X1 U12640 ( .A1(n10072), .A2(n10071), .A3(n10070), .A4(n10069), .ZN(
        n10115) );
  AOI22_X1 U12641 ( .A1(n11173), .A2(keyinput_g59), .B1(keyinput_g6), .B2(
        n12290), .ZN(n10073) );
  OAI221_X1 U12642 ( .B1(n11173), .B2(keyinput_g59), .C1(n12290), .C2(
        keyinput_g6), .A(n10073), .ZN(n10076) );
  XOR2_X1 U12643 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput_g127), .Z(n10075) );
  INV_X1 U12644 ( .A(P3_DATAO_REG_28__SCAN_IN), .ZN(n11925) );
  XNOR2_X1 U12645 ( .A(n11925), .B(keyinput_g68), .ZN(n10074) );
  OR3_X1 U12646 ( .A1(n10076), .A2(n10075), .A3(n10074), .ZN(n10081) );
  INV_X1 U12647 ( .A(P3_DATAO_REG_24__SCAN_IN), .ZN(n11533) );
  AOI22_X1 U12648 ( .A1(P3_U3151), .A2(keyinput_g34), .B1(keyinput_g72), .B2(
        n11533), .ZN(n10077) );
  OAI221_X1 U12649 ( .B1(P3_U3151), .B2(keyinput_g34), .C1(n11533), .C2(
        keyinput_g72), .A(n10077), .ZN(n10080) );
  INV_X1 U12650 ( .A(P3_DATAO_REG_14__SCAN_IN), .ZN(n10664) );
  AOI22_X1 U12651 ( .A1(n10450), .A2(keyinput_g21), .B1(keyinput_g82), .B2(
        n10664), .ZN(n10078) );
  OAI221_X1 U12652 ( .B1(n10450), .B2(keyinput_g21), .C1(n10664), .C2(
        keyinput_g82), .A(n10078), .ZN(n10079) );
  NOR3_X1 U12653 ( .A1(n10081), .A2(n10080), .A3(n10079), .ZN(n10113) );
  INV_X1 U12654 ( .A(P3_DATAO_REG_23__SCAN_IN), .ZN(n11355) );
  AOI22_X1 U12655 ( .A1(n12216), .A2(keyinput_g7), .B1(keyinput_g73), .B2(
        n11355), .ZN(n10082) );
  OAI221_X1 U12656 ( .B1(n12216), .B2(keyinput_g7), .C1(n11355), .C2(
        keyinput_g73), .A(n10082), .ZN(n10090) );
  AOI22_X1 U12657 ( .A1(n10192), .A2(keyinput_g41), .B1(keyinput_g8), .B2(
        n12064), .ZN(n10083) );
  OAI221_X1 U12658 ( .B1(n10192), .B2(keyinput_g41), .C1(n12064), .C2(
        keyinput_g8), .A(n10083), .ZN(n10089) );
  INV_X1 U12659 ( .A(P3_REG3_REG_26__SCAN_IN), .ZN(n10203) );
  AOI22_X1 U12660 ( .A1(n10203), .A2(keyinput_g62), .B1(keyinput_g51), .B2(
        n12753), .ZN(n10084) );
  OAI221_X1 U12661 ( .B1(n10203), .B2(keyinput_g62), .C1(n12753), .C2(
        keyinput_g51), .A(n10084), .ZN(n10088) );
  INV_X1 U12662 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n11159) );
  XOR2_X1 U12663 ( .A(n11159), .B(keyinput_g35), .Z(n10086) );
  XNOR2_X1 U12664 ( .A(P1_IR_REG_2__SCAN_IN), .B(keyinput_g109), .ZN(n10085)
         );
  NAND2_X1 U12665 ( .A1(n10086), .A2(n10085), .ZN(n10087) );
  NOR4_X1 U12666 ( .A1(n10090), .A2(n10089), .A3(n10088), .A4(n10087), .ZN(
        n10112) );
  AOI22_X1 U12667 ( .A1(n12341), .A2(keyinput_g5), .B1(keyinput_g17), .B2(
        n10594), .ZN(n10091) );
  OAI221_X1 U12668 ( .B1(n12341), .B2(keyinput_g5), .C1(n10594), .C2(
        keyinput_g17), .A(n10091), .ZN(n10094) );
  INV_X1 U12669 ( .A(P3_DATAO_REG_1__SCAN_IN), .ZN(n10691) );
  XNOR2_X1 U12670 ( .A(n10691), .B(keyinput_g95), .ZN(n10093) );
  XOR2_X1 U12671 ( .A(P1_IR_REG_18__SCAN_IN), .B(keyinput_g125), .Z(n10092) );
  OR3_X1 U12672 ( .A1(n10094), .A2(n10093), .A3(n10092), .ZN(n10100) );
  INV_X1 U12673 ( .A(P3_DATAO_REG_30__SCAN_IN), .ZN(n10262) );
  AOI22_X1 U12674 ( .A1(n10262), .A2(keyinput_g66), .B1(n8869), .B2(
        keyinput_g47), .ZN(n10095) );
  OAI221_X1 U12675 ( .B1(n10262), .B2(keyinput_g66), .C1(n8869), .C2(
        keyinput_g47), .A(n10095), .ZN(n10099) );
  INV_X1 U12676 ( .A(P3_DATAO_REG_8__SCAN_IN), .ZN(n10670) );
  AOI22_X1 U12677 ( .A1(n10670), .A2(keyinput_g88), .B1(n10097), .B2(
        keyinput_g10), .ZN(n10096) );
  OAI221_X1 U12678 ( .B1(n10670), .B2(keyinput_g88), .C1(n10097), .C2(
        keyinput_g10), .A(n10096), .ZN(n10098) );
  NOR3_X1 U12679 ( .A1(n10100), .A2(n10099), .A3(n10098), .ZN(n10111) );
  INV_X1 U12680 ( .A(P3_DATAO_REG_18__SCAN_IN), .ZN(n10693) );
  AOI22_X1 U12681 ( .A1(n10693), .A2(keyinput_g78), .B1(n10212), .B2(
        keyinput_g102), .ZN(n10101) );
  OAI221_X1 U12682 ( .B1(n10693), .B2(keyinput_g78), .C1(n10212), .C2(
        keyinput_g102), .A(n10101), .ZN(n10109) );
  INV_X1 U12683 ( .A(P3_DATAO_REG_7__SCAN_IN), .ZN(n10668) );
  AOI22_X1 U12684 ( .A1(n10486), .A2(keyinput_g19), .B1(keyinput_g89), .B2(
        n10668), .ZN(n10102) );
  OAI221_X1 U12685 ( .B1(n10486), .B2(keyinput_g19), .C1(n10668), .C2(
        keyinput_g89), .A(n10102), .ZN(n10108) );
  INV_X1 U12686 ( .A(SI_31_), .ZN(n13429) );
  AOI22_X1 U12687 ( .A1(n10495), .A2(keyinput_g18), .B1(keyinput_g1), .B2(
        n13429), .ZN(n10103) );
  OAI221_X1 U12688 ( .B1(n10495), .B2(keyinput_g18), .C1(n13429), .C2(
        keyinput_g1), .A(n10103), .ZN(n10107) );
  XNOR2_X1 U12689 ( .A(SI_6_), .B(keyinput_g26), .ZN(n10105) );
  XNOR2_X1 U12690 ( .A(SI_9_), .B(keyinput_g23), .ZN(n10104) );
  NAND2_X1 U12691 ( .A1(n10105), .A2(n10104), .ZN(n10106) );
  NOR4_X1 U12692 ( .A1(n10109), .A2(n10108), .A3(n10107), .A4(n10106), .ZN(
        n10110) );
  NAND4_X1 U12693 ( .A1(n10113), .A2(n10112), .A3(n10111), .A4(n10110), .ZN(
        n10114) );
  NOR4_X1 U12694 ( .A1(n10117), .A2(n10116), .A3(n10115), .A4(n10114), .ZN(
        n10337) );
  OAI22_X1 U12695 ( .A1(P3_REG3_REG_20__SCAN_IN), .A2(keyinput_g55), .B1(
        SI_20_), .B2(keyinput_g12), .ZN(n10118) );
  AOI221_X1 U12696 ( .B1(P3_REG3_REG_20__SCAN_IN), .B2(keyinput_g55), .C1(
        keyinput_g12), .C2(SI_20_), .A(n10118), .ZN(n10125) );
  OAI22_X1 U12697 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(keyinput_g126), .B1(
        P3_DATAO_REG_25__SCAN_IN), .B2(keyinput_g71), .ZN(n10119) );
  AOI221_X1 U12698 ( .B1(P1_IR_REG_19__SCAN_IN), .B2(keyinput_g126), .C1(
        keyinput_g71), .C2(P3_DATAO_REG_25__SCAN_IN), .A(n10119), .ZN(n10124)
         );
  OAI22_X1 U12699 ( .A1(P3_REG3_REG_23__SCAN_IN), .A2(keyinput_g38), .B1(
        P1_IR_REG_6__SCAN_IN), .B2(keyinput_g113), .ZN(n10120) );
  AOI221_X1 U12700 ( .B1(P3_REG3_REG_23__SCAN_IN), .B2(keyinput_g38), .C1(
        keyinput_g113), .C2(P1_IR_REG_6__SCAN_IN), .A(n10120), .ZN(n10123) );
  OAI22_X1 U12701 ( .A1(P3_REG3_REG_5__SCAN_IN), .A2(keyinput_g49), .B1(
        P3_ADDR_REG_6__SCAN_IN), .B2(keyinput_g103), .ZN(n10121) );
  AOI221_X1 U12702 ( .B1(P3_REG3_REG_5__SCAN_IN), .B2(keyinput_g49), .C1(
        keyinput_g103), .C2(P3_ADDR_REG_6__SCAN_IN), .A(n10121), .ZN(n10122)
         );
  NAND4_X1 U12703 ( .A1(n10125), .A2(n10124), .A3(n10123), .A4(n10122), .ZN(
        n10153) );
  OAI22_X1 U12704 ( .A1(SI_21_), .A2(keyinput_g11), .B1(SI_18_), .B2(
        keyinput_g14), .ZN(n10126) );
  AOI221_X1 U12705 ( .B1(SI_21_), .B2(keyinput_g11), .C1(keyinput_g14), .C2(
        SI_18_), .A(n10126), .ZN(n10133) );
  OAI22_X1 U12706 ( .A1(P3_REG3_REG_9__SCAN_IN), .A2(keyinput_g53), .B1(
        keyinput_g0), .B2(P3_WR_REG_SCAN_IN), .ZN(n10127) );
  AOI221_X1 U12707 ( .B1(P3_REG3_REG_9__SCAN_IN), .B2(keyinput_g53), .C1(
        P3_WR_REG_SCAN_IN), .C2(keyinput_g0), .A(n10127), .ZN(n10132) );
  OAI22_X1 U12708 ( .A1(SI_2_), .A2(keyinput_g30), .B1(P3_DATAO_REG_2__SCAN_IN), .B2(keyinput_g94), .ZN(n10128) );
  AOI221_X1 U12709 ( .B1(SI_2_), .B2(keyinput_g30), .C1(keyinput_g94), .C2(
        P3_DATAO_REG_2__SCAN_IN), .A(n10128), .ZN(n10131) );
  OAI22_X1 U12710 ( .A1(P3_REG3_REG_17__SCAN_IN), .A2(keyinput_g50), .B1(
        P1_IR_REG_10__SCAN_IN), .B2(keyinput_g117), .ZN(n10129) );
  AOI221_X1 U12711 ( .B1(P3_REG3_REG_17__SCAN_IN), .B2(keyinput_g50), .C1(
        keyinput_g117), .C2(P1_IR_REG_10__SCAN_IN), .A(n10129), .ZN(n10130) );
  NAND4_X1 U12712 ( .A1(n10133), .A2(n10132), .A3(n10131), .A4(n10130), .ZN(
        n10152) );
  OAI22_X1 U12713 ( .A1(SI_3_), .A2(keyinput_g29), .B1(keyinput_g32), .B2(
        SI_0_), .ZN(n10134) );
  AOI221_X1 U12714 ( .B1(SI_3_), .B2(keyinput_g29), .C1(SI_0_), .C2(
        keyinput_g32), .A(n10134), .ZN(n10141) );
  OAI22_X1 U12715 ( .A1(P3_REG3_REG_22__SCAN_IN), .A2(keyinput_g57), .B1(
        P3_REG3_REG_18__SCAN_IN), .B2(keyinput_g60), .ZN(n10135) );
  AOI221_X1 U12716 ( .B1(P3_REG3_REG_22__SCAN_IN), .B2(keyinput_g57), .C1(
        keyinput_g60), .C2(P3_REG3_REG_18__SCAN_IN), .A(n10135), .ZN(n10140)
         );
  OAI22_X1 U12717 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(keyinput_g122), .B1(
        keyinput_g99), .B2(P3_ADDR_REG_2__SCAN_IN), .ZN(n10136) );
  AOI221_X1 U12718 ( .B1(P1_IR_REG_15__SCAN_IN), .B2(keyinput_g122), .C1(
        P3_ADDR_REG_2__SCAN_IN), .C2(keyinput_g99), .A(n10136), .ZN(n10139) );
  OAI22_X1 U12719 ( .A1(P3_REG3_REG_13__SCAN_IN), .A2(keyinput_g56), .B1(
        SI_17_), .B2(keyinput_g15), .ZN(n10137) );
  AOI221_X1 U12720 ( .B1(P3_REG3_REG_13__SCAN_IN), .B2(keyinput_g56), .C1(
        keyinput_g15), .C2(SI_17_), .A(n10137), .ZN(n10138) );
  NAND4_X1 U12721 ( .A1(n10141), .A2(n10140), .A3(n10139), .A4(n10138), .ZN(
        n10151) );
  OAI22_X1 U12722 ( .A1(P3_REG3_REG_15__SCAN_IN), .A2(keyinput_g63), .B1(
        keyinput_g2), .B2(SI_30_), .ZN(n10142) );
  AOI221_X1 U12723 ( .B1(P3_REG3_REG_15__SCAN_IN), .B2(keyinput_g63), .C1(
        SI_30_), .C2(keyinput_g2), .A(n10142), .ZN(n10149) );
  OAI22_X1 U12724 ( .A1(P3_REG3_REG_27__SCAN_IN), .A2(keyinput_g36), .B1(
        P3_DATAO_REG_0__SCAN_IN), .B2(keyinput_g96), .ZN(n10143) );
  AOI221_X1 U12725 ( .B1(P3_REG3_REG_27__SCAN_IN), .B2(keyinput_g36), .C1(
        keyinput_g96), .C2(P3_DATAO_REG_0__SCAN_IN), .A(n10143), .ZN(n10148)
         );
  OAI22_X1 U12726 ( .A1(P3_DATAO_REG_11__SCAN_IN), .A2(keyinput_g85), .B1(
        keyinput_g74), .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n10144) );
  AOI221_X1 U12727 ( .B1(P3_DATAO_REG_11__SCAN_IN), .B2(keyinput_g85), .C1(
        P3_DATAO_REG_22__SCAN_IN), .C2(keyinput_g74), .A(n10144), .ZN(n10147)
         );
  OAI22_X1 U12728 ( .A1(P3_REG3_REG_16__SCAN_IN), .A2(keyinput_g48), .B1(
        keyinput_g9), .B2(SI_23_), .ZN(n10145) );
  AOI221_X1 U12729 ( .B1(P3_REG3_REG_16__SCAN_IN), .B2(keyinput_g48), .C1(
        SI_23_), .C2(keyinput_g9), .A(n10145), .ZN(n10146) );
  NAND4_X1 U12730 ( .A1(n10149), .A2(n10148), .A3(n10147), .A4(n10146), .ZN(
        n10150) );
  NOR4_X1 U12731 ( .A1(n10153), .A2(n10152), .A3(n10151), .A4(n10150), .ZN(
        n10336) );
  AOI22_X1 U12732 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(keyinput_f120), .B1(SI_25_), .B2(keyinput_f7), .ZN(n10154) );
  OAI221_X1 U12733 ( .B1(P1_IR_REG_13__SCAN_IN), .B2(keyinput_f120), .C1(
        SI_25_), .C2(keyinput_f7), .A(n10154), .ZN(n10161) );
  AOI22_X1 U12734 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(keyinput_f109), .B1(
        P3_REG3_REG_16__SCAN_IN), .B2(keyinput_f48), .ZN(n10155) );
  OAI221_X1 U12735 ( .B1(P1_IR_REG_2__SCAN_IN), .B2(keyinput_f109), .C1(
        P3_REG3_REG_16__SCAN_IN), .C2(keyinput_f48), .A(n10155), .ZN(n10160)
         );
  AOI22_X1 U12736 ( .A1(keyinput_f86), .A2(P3_DATAO_REG_10__SCAN_IN), .B1(
        P3_ADDR_REG_8__SCAN_IN), .B2(keyinput_f105), .ZN(n10156) );
  OAI221_X1 U12737 ( .B1(keyinput_f86), .B2(P3_DATAO_REG_10__SCAN_IN), .C1(
        P3_ADDR_REG_8__SCAN_IN), .C2(keyinput_f105), .A(n10156), .ZN(n10159)
         );
  AOI22_X1 U12738 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(keyinput_f108), .B1(SI_14_), 
        .B2(keyinput_f18), .ZN(n10157) );
  OAI221_X1 U12739 ( .B1(P1_IR_REG_1__SCAN_IN), .B2(keyinput_f108), .C1(SI_14_), .C2(keyinput_f18), .A(n10157), .ZN(n10158) );
  NOR4_X1 U12740 ( .A1(n10161), .A2(n10160), .A3(n10159), .A4(n10158), .ZN(
        n10330) );
  AOI22_X1 U12741 ( .A1(SI_22_), .A2(keyinput_f10), .B1(
        P3_REG3_REG_15__SCAN_IN), .B2(keyinput_f63), .ZN(n10162) );
  OAI221_X1 U12742 ( .B1(SI_22_), .B2(keyinput_f10), .C1(
        P3_REG3_REG_15__SCAN_IN), .C2(keyinput_f63), .A(n10162), .ZN(n10187)
         );
  OAI22_X1 U12743 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(keyinput_f112), .B1(
        keyinput_f96), .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n10163) );
  AOI221_X1 U12744 ( .B1(P1_IR_REG_5__SCAN_IN), .B2(keyinput_f112), .C1(
        P3_DATAO_REG_0__SCAN_IN), .C2(keyinput_f96), .A(n10163), .ZN(n10167)
         );
  AOI22_X1 U12745 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(keyinput_f119), .B1(
        P3_STATE_REG_SCAN_IN), .B2(keyinput_f34), .ZN(n10164) );
  OAI221_X1 U12746 ( .B1(P1_IR_REG_12__SCAN_IN), .B2(keyinput_f119), .C1(
        P3_STATE_REG_SCAN_IN), .C2(keyinput_f34), .A(n10164), .ZN(n10165) );
  AOI21_X1 U12747 ( .B1(keyinput_f77), .B2(n10709), .A(n10165), .ZN(n10166) );
  OAI211_X1 U12748 ( .C1(keyinput_f77), .C2(n10709), .A(n10167), .B(n10166), 
        .ZN(n10186) );
  OAI22_X1 U12749 ( .A1(P3_REG3_REG_1__SCAN_IN), .A2(keyinput_f44), .B1(
        keyinput_f91), .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n10168) );
  AOI221_X1 U12750 ( .B1(P3_REG3_REG_1__SCAN_IN), .B2(keyinput_f44), .C1(
        P3_DATAO_REG_5__SCAN_IN), .C2(keyinput_f91), .A(n10168), .ZN(n10175)
         );
  OAI22_X1 U12751 ( .A1(SI_29_), .A2(keyinput_f3), .B1(keyinput_f20), .B2(
        SI_12_), .ZN(n10169) );
  AOI221_X1 U12752 ( .B1(SI_29_), .B2(keyinput_f3), .C1(SI_12_), .C2(
        keyinput_f20), .A(n10169), .ZN(n10174) );
  OAI22_X1 U12753 ( .A1(SI_3_), .A2(keyinput_f29), .B1(keyinput_f87), .B2(
        P3_DATAO_REG_9__SCAN_IN), .ZN(n10170) );
  AOI221_X1 U12754 ( .B1(SI_3_), .B2(keyinput_f29), .C1(
        P3_DATAO_REG_9__SCAN_IN), .C2(keyinput_f87), .A(n10170), .ZN(n10173)
         );
  OAI22_X1 U12755 ( .A1(SI_2_), .A2(keyinput_f30), .B1(
        P3_DATAO_REG_28__SCAN_IN), .B2(keyinput_f68), .ZN(n10171) );
  AOI221_X1 U12756 ( .B1(SI_2_), .B2(keyinput_f30), .C1(keyinput_f68), .C2(
        P3_DATAO_REG_28__SCAN_IN), .A(n10171), .ZN(n10172) );
  NAND4_X1 U12757 ( .A1(n10175), .A2(n10174), .A3(n10173), .A4(n10172), .ZN(
        n10185) );
  OAI22_X1 U12758 ( .A1(P3_REG3_REG_20__SCAN_IN), .A2(keyinput_f55), .B1(
        SI_31_), .B2(keyinput_f1), .ZN(n10176) );
  AOI221_X1 U12759 ( .B1(P3_REG3_REG_20__SCAN_IN), .B2(keyinput_f55), .C1(
        keyinput_f1), .C2(SI_31_), .A(n10176), .ZN(n10183) );
  OAI22_X1 U12760 ( .A1(SI_13_), .A2(keyinput_f19), .B1(P1_IR_REG_17__SCAN_IN), 
        .B2(keyinput_f124), .ZN(n10177) );
  AOI221_X1 U12761 ( .B1(SI_13_), .B2(keyinput_f19), .C1(keyinput_f124), .C2(
        P1_IR_REG_17__SCAN_IN), .A(n10177), .ZN(n10182) );
  OAI22_X1 U12762 ( .A1(P3_REG3_REG_0__SCAN_IN), .A2(keyinput_f54), .B1(
        keyinput_f117), .B2(P1_IR_REG_10__SCAN_IN), .ZN(n10178) );
  AOI221_X1 U12763 ( .B1(P3_REG3_REG_0__SCAN_IN), .B2(keyinput_f54), .C1(
        P1_IR_REG_10__SCAN_IN), .C2(keyinput_f117), .A(n10178), .ZN(n10181) );
  OAI22_X1 U12764 ( .A1(keyinput_f33), .A2(P3_RD_REG_SCAN_IN), .B1(
        keyinput_f76), .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n10179) );
  AOI221_X1 U12765 ( .B1(keyinput_f33), .B2(P3_RD_REG_SCAN_IN), .C1(
        P3_DATAO_REG_20__SCAN_IN), .C2(keyinput_f76), .A(n10179), .ZN(n10180)
         );
  NAND4_X1 U12766 ( .A1(n10183), .A2(n10182), .A3(n10181), .A4(n10180), .ZN(
        n10184) );
  NOR4_X1 U12767 ( .A1(n10187), .A2(n10186), .A3(n10185), .A4(n10184), .ZN(
        n10329) );
  INV_X1 U12768 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n10189) );
  OAI22_X1 U12769 ( .A1(n12341), .A2(keyinput_f5), .B1(n10189), .B2(
        keyinput_f99), .ZN(n10188) );
  AOI221_X1 U12770 ( .B1(n12341), .B2(keyinput_f5), .C1(keyinput_f99), .C2(
        n10189), .A(n10188), .ZN(n10200) );
  OAI22_X1 U12771 ( .A1(n10192), .A2(keyinput_f41), .B1(n10191), .B2(
        keyinput_f116), .ZN(n10190) );
  AOI221_X1 U12772 ( .B1(n10192), .B2(keyinput_f41), .C1(keyinput_f116), .C2(
        n10191), .A(n10190), .ZN(n10199) );
  OAI22_X1 U12773 ( .A1(n11544), .A2(keyinput_f11), .B1(n10693), .B2(
        keyinput_f78), .ZN(n10193) );
  AOI221_X1 U12774 ( .B1(n11544), .B2(keyinput_f11), .C1(keyinput_f78), .C2(
        n10693), .A(n10193), .ZN(n10198) );
  INV_X1 U12775 ( .A(P3_REG3_REG_23__SCAN_IN), .ZN(n10196) );
  OAI22_X1 U12776 ( .A1(n10196), .A2(keyinput_f38), .B1(n10195), .B2(
        keyinput_f100), .ZN(n10194) );
  AOI221_X1 U12777 ( .B1(n10196), .B2(keyinput_f38), .C1(keyinput_f100), .C2(
        n10195), .A(n10194), .ZN(n10197) );
  NAND4_X1 U12778 ( .A1(n10200), .A2(n10199), .A3(n10198), .A4(n10197), .ZN(
        n10236) );
  INV_X1 U12779 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n11995) );
  OAI22_X1 U12780 ( .A1(n12753), .A2(keyinput_f51), .B1(n11995), .B2(
        keyinput_f65), .ZN(n10201) );
  AOI221_X1 U12781 ( .B1(n12753), .B2(keyinput_f51), .C1(keyinput_f65), .C2(
        n11995), .A(n10201), .ZN(n10210) );
  OAI22_X1 U12782 ( .A1(n10203), .A2(keyinput_f62), .B1(n10711), .B2(
        keyinput_f16), .ZN(n10202) );
  AOI221_X1 U12783 ( .B1(n10203), .B2(keyinput_f62), .C1(keyinput_f16), .C2(
        n10711), .A(n10202), .ZN(n10209) );
  XNOR2_X1 U12784 ( .A(SI_1_), .B(keyinput_f31), .ZN(n10207) );
  XNOR2_X1 U12785 ( .A(P1_IR_REG_19__SCAN_IN), .B(keyinput_f126), .ZN(n10206)
         );
  XNOR2_X1 U12786 ( .A(P3_REG3_REG_6__SCAN_IN), .B(keyinput_f61), .ZN(n10205)
         );
  XNOR2_X1 U12787 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput_f127), .ZN(n10204)
         );
  AND4_X1 U12788 ( .A1(n10207), .A2(n10206), .A3(n10205), .A4(n10204), .ZN(
        n10208) );
  NAND3_X1 U12789 ( .A1(n10210), .A2(n10209), .A3(n10208), .ZN(n10235) );
  OAI22_X1 U12790 ( .A1(n10212), .A2(keyinput_f102), .B1(n10670), .B2(
        keyinput_f88), .ZN(n10211) );
  AOI221_X1 U12791 ( .B1(n10212), .B2(keyinput_f102), .C1(keyinput_f88), .C2(
        n10670), .A(n10211), .ZN(n10220) );
  OAI22_X1 U12792 ( .A1(n12220), .A2(keyinput_f46), .B1(n8596), .B2(
        keyinput_f53), .ZN(n10213) );
  AOI221_X1 U12793 ( .B1(n12220), .B2(keyinput_f46), .C1(keyinput_f53), .C2(
        n8596), .A(n10213), .ZN(n10219) );
  OAI22_X1 U12794 ( .A1(n11862), .A2(keyinput_f39), .B1(n12064), .B2(
        keyinput_f8), .ZN(n10214) );
  AOI221_X1 U12795 ( .B1(n11862), .B2(keyinput_f39), .C1(keyinput_f8), .C2(
        n12064), .A(n10214), .ZN(n10218) );
  XOR2_X1 U12796 ( .A(SI_4_), .B(keyinput_f28), .Z(n10216) );
  XNOR2_X1 U12797 ( .A(keyinput_f35), .B(n11159), .ZN(n10215) );
  NOR2_X1 U12798 ( .A1(n10216), .A2(n10215), .ZN(n10217) );
  NAND4_X1 U12799 ( .A1(n10220), .A2(n10219), .A3(n10218), .A4(n10217), .ZN(
        n10234) );
  OAI22_X1 U12800 ( .A1(n10223), .A2(keyinput_f45), .B1(n10222), .B2(
        keyinput_f101), .ZN(n10221) );
  AOI221_X1 U12801 ( .B1(n10223), .B2(keyinput_f45), .C1(keyinput_f101), .C2(
        n10222), .A(n10221), .ZN(n10232) );
  OAI22_X1 U12802 ( .A1(n10879), .A2(keyinput_f14), .B1(n10450), .B2(
        keyinput_f21), .ZN(n10224) );
  AOI221_X1 U12803 ( .B1(n10879), .B2(keyinput_f14), .C1(keyinput_f21), .C2(
        n10450), .A(n10224), .ZN(n10231) );
  OAI22_X1 U12804 ( .A1(n10940), .A2(keyinput_f52), .B1(n12290), .B2(
        keyinput_f6), .ZN(n10225) );
  AOI221_X1 U12805 ( .B1(n10940), .B2(keyinput_f52), .C1(keyinput_f6), .C2(
        n12290), .A(n10225), .ZN(n10230) );
  XOR2_X1 U12806 ( .A(P1_IR_REG_18__SCAN_IN), .B(keyinput_f125), .Z(n10228) );
  XNOR2_X1 U12807 ( .A(keyinput_f103), .B(n10226), .ZN(n10227) );
  NOR2_X1 U12808 ( .A1(n10228), .A2(n10227), .ZN(n10229) );
  NAND4_X1 U12809 ( .A1(n10232), .A2(n10231), .A3(n10230), .A4(n10229), .ZN(
        n10233) );
  NOR4_X1 U12810 ( .A1(n10236), .A2(n10235), .A3(n10234), .A4(n10233), .ZN(
        n10328) );
  AOI22_X1 U12811 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(keyinput_f113), .B1(
        P3_B_REG_SCAN_IN), .B2(keyinput_f64), .ZN(n10237) );
  OAI221_X1 U12812 ( .B1(P1_IR_REG_6__SCAN_IN), .B2(keyinput_f113), .C1(
        P3_B_REG_SCAN_IN), .C2(keyinput_f64), .A(n10237), .ZN(n10244) );
  AOI22_X1 U12813 ( .A1(keyinput_f85), .A2(P3_DATAO_REG_11__SCAN_IN), .B1(
        keyinput_f72), .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n10238) );
  OAI221_X1 U12814 ( .B1(keyinput_f85), .B2(P3_DATAO_REG_11__SCAN_IN), .C1(
        keyinput_f72), .C2(P3_DATAO_REG_24__SCAN_IN), .A(n10238), .ZN(n10243)
         );
  AOI22_X1 U12815 ( .A1(keyinput_f93), .A2(P3_DATAO_REG_3__SCAN_IN), .B1(
        keyinput_f94), .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n10239) );
  OAI221_X1 U12816 ( .B1(keyinput_f93), .B2(P3_DATAO_REG_3__SCAN_IN), .C1(
        keyinput_f94), .C2(P3_DATAO_REG_2__SCAN_IN), .A(n10239), .ZN(n10242)
         );
  AOI22_X1 U12817 ( .A1(keyinput_f67), .A2(P3_DATAO_REG_29__SCAN_IN), .B1(
        P1_IR_REG_16__SCAN_IN), .B2(keyinput_f123), .ZN(n10240) );
  OAI221_X1 U12818 ( .B1(keyinput_f67), .B2(P3_DATAO_REG_29__SCAN_IN), .C1(
        P1_IR_REG_16__SCAN_IN), .C2(keyinput_f123), .A(n10240), .ZN(n10241) );
  NOR4_X1 U12819 ( .A1(n10244), .A2(n10243), .A3(n10242), .A4(n10241), .ZN(
        n10275) );
  AOI22_X1 U12820 ( .A1(P3_ADDR_REG_7__SCAN_IN), .A2(keyinput_f104), .B1(SI_7_), .B2(keyinput_f25), .ZN(n10245) );
  OAI221_X1 U12821 ( .B1(P3_ADDR_REG_7__SCAN_IN), .B2(keyinput_f104), .C1(
        SI_7_), .C2(keyinput_f25), .A(n10245), .ZN(n10252) );
  AOI22_X1 U12822 ( .A1(keyinput_f89), .A2(P3_DATAO_REG_7__SCAN_IN), .B1(
        P3_REG3_REG_8__SCAN_IN), .B2(keyinput_f43), .ZN(n10246) );
  OAI221_X1 U12823 ( .B1(keyinput_f89), .B2(P3_DATAO_REG_7__SCAN_IN), .C1(
        P3_REG3_REG_8__SCAN_IN), .C2(keyinput_f43), .A(n10246), .ZN(n10251) );
  AOI22_X1 U12824 ( .A1(keyinput_f81), .A2(P3_DATAO_REG_15__SCAN_IN), .B1(
        SI_20_), .B2(keyinput_f12), .ZN(n10247) );
  OAI221_X1 U12825 ( .B1(keyinput_f81), .B2(P3_DATAO_REG_15__SCAN_IN), .C1(
        SI_20_), .C2(keyinput_f12), .A(n10247), .ZN(n10250) );
  AOI22_X1 U12826 ( .A1(keyinput_f84), .A2(P3_DATAO_REG_12__SCAN_IN), .B1(
        keyinput_f74), .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n10248) );
  OAI221_X1 U12827 ( .B1(keyinput_f84), .B2(P3_DATAO_REG_12__SCAN_IN), .C1(
        keyinput_f74), .C2(P3_DATAO_REG_22__SCAN_IN), .A(n10248), .ZN(n10249)
         );
  NOR4_X1 U12828 ( .A1(n10252), .A2(n10251), .A3(n10250), .A4(n10249), .ZN(
        n10274) );
  AOI22_X1 U12829 ( .A1(keyinput_f79), .A2(P3_DATAO_REG_17__SCAN_IN), .B1(
        SI_28_), .B2(keyinput_f4), .ZN(n10253) );
  OAI221_X1 U12830 ( .B1(keyinput_f79), .B2(P3_DATAO_REG_17__SCAN_IN), .C1(
        SI_28_), .C2(keyinput_f4), .A(n10253), .ZN(n10260) );
  AOI22_X1 U12831 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(keyinput_f115), .B1(
        P3_REG3_REG_17__SCAN_IN), .B2(keyinput_f50), .ZN(n10254) );
  OAI221_X1 U12832 ( .B1(P1_IR_REG_8__SCAN_IN), .B2(keyinput_f115), .C1(
        P3_REG3_REG_17__SCAN_IN), .C2(keyinput_f50), .A(n10254), .ZN(n10259)
         );
  AOI22_X1 U12833 ( .A1(keyinput_f70), .A2(P3_DATAO_REG_26__SCAN_IN), .B1(
        keyinput_f73), .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n10255) );
  OAI221_X1 U12834 ( .B1(keyinput_f70), .B2(P3_DATAO_REG_26__SCAN_IN), .C1(
        keyinput_f73), .C2(P3_DATAO_REG_23__SCAN_IN), .A(n10255), .ZN(n10258)
         );
  AOI22_X1 U12835 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(keyinput_f110), .B1(
        P3_REG3_REG_27__SCAN_IN), .B2(keyinput_f36), .ZN(n10256) );
  OAI221_X1 U12836 ( .B1(P1_IR_REG_3__SCAN_IN), .B2(keyinput_f110), .C1(
        P3_REG3_REG_27__SCAN_IN), .C2(keyinput_f36), .A(n10256), .ZN(n10257)
         );
  NOR4_X1 U12837 ( .A1(n10260), .A2(n10259), .A3(n10258), .A4(n10257), .ZN(
        n10273) );
  AOI22_X1 U12838 ( .A1(n10666), .A2(keyinput_f90), .B1(keyinput_f66), .B2(
        n10262), .ZN(n10261) );
  OAI221_X1 U12839 ( .B1(n10666), .B2(keyinput_f90), .C1(n10262), .C2(
        keyinput_f66), .A(n10261), .ZN(n10271) );
  AOI22_X1 U12840 ( .A1(keyinput_f82), .A2(P3_DATAO_REG_14__SCAN_IN), .B1(
        keyinput_f69), .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n10263) );
  OAI221_X1 U12841 ( .B1(keyinput_f82), .B2(P3_DATAO_REG_14__SCAN_IN), .C1(
        keyinput_f69), .C2(P3_DATAO_REG_27__SCAN_IN), .A(n10263), .ZN(n10270)
         );
  INV_X1 U12842 ( .A(SI_10_), .ZN(n10449) );
  INV_X1 U12843 ( .A(P3_REG3_REG_18__SCAN_IN), .ZN(n10265) );
  AOI22_X1 U12844 ( .A1(n10449), .A2(keyinput_f22), .B1(n10265), .B2(
        keyinput_f60), .ZN(n10264) );
  OAI221_X1 U12845 ( .B1(n10449), .B2(keyinput_f22), .C1(n10265), .C2(
        keyinput_f60), .A(n10264), .ZN(n10269) );
  XOR2_X1 U12846 ( .A(P3_ADDR_REG_9__SCAN_IN), .B(keyinput_f106), .Z(n10267)
         );
  XNOR2_X1 U12847 ( .A(SI_9_), .B(keyinput_f23), .ZN(n10266) );
  NAND2_X1 U12848 ( .A1(n10267), .A2(n10266), .ZN(n10268) );
  NOR4_X1 U12849 ( .A1(n10271), .A2(n10270), .A3(n10269), .A4(n10268), .ZN(
        n10272) );
  NAND4_X1 U12850 ( .A1(n10275), .A2(n10274), .A3(n10273), .A4(n10272), .ZN(
        n10326) );
  AOI22_X1 U12851 ( .A1(n10277), .A2(keyinput_f121), .B1(n10454), .B2(
        keyinput_f32), .ZN(n10276) );
  OAI221_X1 U12852 ( .B1(n10277), .B2(keyinput_f121), .C1(n10454), .C2(
        keyinput_f32), .A(n10276), .ZN(n10325) );
  INV_X1 U12853 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n12179) );
  INV_X1 U12854 ( .A(P3_DATAO_REG_21__SCAN_IN), .ZN(n11012) );
  OAI22_X1 U12855 ( .A1(n12179), .A2(keyinput_f58), .B1(n11012), .B2(
        keyinput_f75), .ZN(n10278) );
  AOI221_X1 U12856 ( .B1(n12179), .B2(keyinput_f58), .C1(keyinput_f75), .C2(
        n11012), .A(n10278), .ZN(n10285) );
  XOR2_X1 U12857 ( .A(n10677), .B(keyinput_f80), .Z(n10284) );
  XNOR2_X1 U12858 ( .A(keyinput_f0), .B(P3_WR_REG_SCAN_IN), .ZN(n10283) );
  XOR2_X1 U12859 ( .A(SI_5_), .B(keyinput_f27), .Z(n10281) );
  INV_X1 U12860 ( .A(P3_REG3_REG_22__SCAN_IN), .ZN(n10279) );
  XNOR2_X1 U12861 ( .A(keyinput_f57), .B(n10279), .ZN(n10280) );
  NOR2_X1 U12862 ( .A1(n10281), .A2(n10280), .ZN(n10282) );
  NAND4_X1 U12863 ( .A1(n10285), .A2(n10284), .A3(n10283), .A4(n10282), .ZN(
        n10324) );
  INV_X1 U12864 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n10287) );
  INV_X1 U12865 ( .A(P3_DATAO_REG_25__SCAN_IN), .ZN(n11634) );
  AOI22_X1 U12866 ( .A1(n10287), .A2(keyinput_f122), .B1(keyinput_f71), .B2(
        n11634), .ZN(n10286) );
  OAI221_X1 U12867 ( .B1(n10287), .B2(keyinput_f122), .C1(n11634), .C2(
        keyinput_f71), .A(n10286), .ZN(n10296) );
  AOI22_X1 U12868 ( .A1(n10289), .A2(keyinput_f98), .B1(n8869), .B2(
        keyinput_f47), .ZN(n10288) );
  OAI221_X1 U12869 ( .B1(n10289), .B2(keyinput_f98), .C1(n8869), .C2(
        keyinput_f47), .A(n10288), .ZN(n10295) );
  AOI22_X1 U12870 ( .A1(n8527), .A2(keyinput_f49), .B1(keyinput_f17), .B2(
        n10594), .ZN(n10290) );
  OAI221_X1 U12871 ( .B1(n8527), .B2(keyinput_f49), .C1(n10594), .C2(
        keyinput_f17), .A(n10290), .ZN(n10294) );
  XNOR2_X1 U12872 ( .A(P1_IR_REG_0__SCAN_IN), .B(keyinput_f107), .ZN(n10292)
         );
  XNOR2_X1 U12873 ( .A(SI_23_), .B(keyinput_f9), .ZN(n10291) );
  NAND2_X1 U12874 ( .A1(n10292), .A2(n10291), .ZN(n10293) );
  NOR4_X1 U12875 ( .A1(n10296), .A2(n10295), .A3(n10294), .A4(n10293), .ZN(
        n10322) );
  INV_X1 U12876 ( .A(P3_DATAO_REG_4__SCAN_IN), .ZN(n10658) );
  AOI22_X1 U12877 ( .A1(n10298), .A2(keyinput_f118), .B1(keyinput_f92), .B2(
        n10658), .ZN(n10297) );
  OAI221_X1 U12878 ( .B1(n10298), .B2(keyinput_f118), .C1(n10658), .C2(
        keyinput_f92), .A(n10297), .ZN(n10300) );
  XNOR2_X1 U12879 ( .A(n10691), .B(keyinput_f95), .ZN(n10299) );
  NOR2_X1 U12880 ( .A1(n10300), .A2(n10299), .ZN(n10308) );
  INV_X1 U12881 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n12020) );
  AOI22_X1 U12882 ( .A1(n10672), .A2(keyinput_f83), .B1(n12020), .B2(
        keyinput_f40), .ZN(n10301) );
  OAI221_X1 U12883 ( .B1(n10672), .B2(keyinput_f83), .C1(n12020), .C2(
        keyinput_f40), .A(n10301), .ZN(n10302) );
  INV_X1 U12884 ( .A(n10302), .ZN(n10307) );
  INV_X1 U12885 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n12333) );
  AOI22_X1 U12886 ( .A1(n12333), .A2(keyinput_f37), .B1(keyinput_f97), .B2(
        n15549), .ZN(n10303) );
  OAI221_X1 U12887 ( .B1(n12333), .B2(keyinput_f37), .C1(n15549), .C2(
        keyinput_f97), .A(n10303), .ZN(n10304) );
  INV_X1 U12888 ( .A(n10304), .ZN(n10306) );
  XNOR2_X1 U12889 ( .A(SI_6_), .B(keyinput_f26), .ZN(n10305) );
  AND4_X1 U12890 ( .A1(n10308), .A2(n10307), .A3(n10306), .A4(n10305), .ZN(
        n10321) );
  INV_X1 U12891 ( .A(SI_30_), .ZN(n10310) );
  AOI22_X1 U12892 ( .A1(n8684), .A2(keyinput_f56), .B1(keyinput_f2), .B2(
        n10310), .ZN(n10309) );
  OAI221_X1 U12893 ( .B1(n8684), .B2(keyinput_f56), .C1(n10310), .C2(
        keyinput_f2), .A(n10309), .ZN(n10319) );
  AOI22_X1 U12894 ( .A1(n11173), .A2(keyinput_f59), .B1(keyinput_f15), .B2(
        n10834), .ZN(n10311) );
  OAI221_X1 U12895 ( .B1(n11173), .B2(keyinput_f59), .C1(n10834), .C2(
        keyinput_f15), .A(n10311), .ZN(n10318) );
  XNOR2_X1 U12896 ( .A(SI_19_), .B(keyinput_f13), .ZN(n10316) );
  XNOR2_X1 U12897 ( .A(SI_8_), .B(keyinput_f24), .ZN(n10315) );
  XNOR2_X1 U12898 ( .A(n10312), .B(keyinput_f114), .ZN(n10314) );
  XNOR2_X1 U12899 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput_f111), .ZN(n10313)
         );
  NAND4_X1 U12900 ( .A1(n10316), .A2(n10315), .A3(n10314), .A4(n10313), .ZN(
        n10317) );
  NOR3_X1 U12901 ( .A1(n10319), .A2(n10318), .A3(n10317), .ZN(n10320) );
  NAND3_X1 U12902 ( .A1(n10322), .A2(n10321), .A3(n10320), .ZN(n10323) );
  NOR4_X1 U12903 ( .A1(n10326), .A2(n10325), .A3(n10324), .A4(n10323), .ZN(
        n10327) );
  NAND4_X1 U12904 ( .A1(n10330), .A2(n10329), .A3(n10328), .A4(n10327), .ZN(
        n10332) );
  AOI21_X1 U12905 ( .B1(keyinput_f42), .B2(n10332), .A(P3_REG3_REG_28__SCAN_IN), .ZN(n10334) );
  INV_X1 U12906 ( .A(keyinput_f42), .ZN(n10331) );
  AOI21_X1 U12907 ( .B1(n10332), .B2(n10331), .A(keyinput_g42), .ZN(n10333) );
  AOI22_X1 U12908 ( .A1(keyinput_g42), .A2(n10334), .B1(
        P3_REG3_REG_28__SCAN_IN), .B2(n10333), .ZN(n10335) );
  AOI21_X1 U12909 ( .B1(n10337), .B2(n10336), .A(n10335), .ZN(n10338) );
  INV_X1 U12910 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n10378) );
  INV_X1 U12911 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n10341) );
  AND2_X1 U12912 ( .A1(n10341), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n10342) );
  NAND2_X1 U12913 ( .A1(n14886), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n10344) );
  INV_X1 U12914 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n10350) );
  XNOR2_X1 U12915 ( .A(n10350), .B(P2_DATAO_REG_28__SCAN_IN), .ZN(n10345) );
  NAND2_X1 U12916 ( .A1(n12664), .A2(n12805), .ZN(n10347) );
  OR2_X1 U12917 ( .A1(n12806), .A2(n12668), .ZN(n10346) );
  NAND2_X1 U12918 ( .A1(n13095), .A2(n10366), .ZN(n10363) );
  NAND2_X1 U12919 ( .A1(n10363), .A2(n13083), .ZN(n12971) );
  AND2_X1 U12920 ( .A1(n12663), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n10348) );
  NAND2_X1 U12921 ( .A1(n10350), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n10351) );
  XNOR2_X1 U12922 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .ZN(n12685) );
  XNOR2_X1 U12923 ( .A(n12687), .B(n12685), .ZN(n13436) );
  NAND2_X1 U12924 ( .A1(n13436), .A2(n12805), .ZN(n10354) );
  OR2_X1 U12925 ( .A1(n12806), .A2(n13439), .ZN(n10353) );
  NAND2_X1 U12926 ( .A1(n13070), .A2(n10356), .ZN(n11993) );
  NAND2_X1 U12927 ( .A1(n11984), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n10358) );
  INV_X1 U12928 ( .A(P3_REG2_REG_29__SCAN_IN), .ZN(n13077) );
  OR2_X1 U12929 ( .A1(n11986), .A2(n13077), .ZN(n10357) );
  OAI211_X1 U12930 ( .C1(n10378), .C2(n11989), .A(n10358), .B(n10357), .ZN(
        n10359) );
  INV_X1 U12931 ( .A(n10359), .ZN(n10360) );
  NAND2_X1 U12932 ( .A1(n11993), .A2(n10360), .ZN(n12673) );
  NAND2_X1 U12933 ( .A1(n13079), .A2(n13092), .ZN(n12810) );
  NAND2_X1 U12934 ( .A1(n12834), .A2(n12810), .ZN(n10364) );
  AOI21_X1 U12935 ( .B1(n13095), .B2(n11923), .A(n13088), .ZN(n10365) );
  NOR2_X1 U12936 ( .A1(n13276), .A2(n10366), .ZN(n10376) );
  INV_X1 U12937 ( .A(P3_REG0_REG_30__SCAN_IN), .ZN(n10370) );
  NAND2_X1 U12938 ( .A1(n11984), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n10369) );
  INV_X1 U12939 ( .A(P3_REG2_REG_30__SCAN_IN), .ZN(n10367) );
  OR2_X1 U12940 ( .A1(n11986), .A2(n10367), .ZN(n10368) );
  OAI211_X1 U12941 ( .C1(n10370), .C2(n11989), .A(n10369), .B(n10368), .ZN(
        n10371) );
  INV_X1 U12942 ( .A(n10371), .ZN(n10372) );
  AND2_X1 U12943 ( .A1(n11993), .A2(n10372), .ZN(n12809) );
  NOR2_X1 U12944 ( .A1(n12667), .A2(n10373), .ZN(n10374) );
  OR2_X1 U12945 ( .A1(n13278), .A2(n10374), .ZN(n13068) );
  NOR2_X1 U12946 ( .A1(n12809), .A2(n13068), .ZN(n10375) );
  INV_X1 U12947 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n10381) );
  INV_X1 U12948 ( .A(n10474), .ZN(n10385) );
  NAND2_X1 U12949 ( .A1(n10383), .A2(P1_D_REG_1__SCAN_IN), .ZN(n10384) );
  AOI21_X1 U12950 ( .B1(n10385), .B2(n10384), .A(n10475), .ZN(n10719) );
  INV_X1 U12951 ( .A(n14472), .ZN(n11095) );
  AND2_X1 U12952 ( .A1(n10719), .A2(n11095), .ZN(n10387) );
  INV_X1 U12953 ( .A(n11096), .ZN(n10386) );
  NAND2_X1 U12954 ( .A1(n10387), .A2(n10386), .ZN(n10391) );
  NAND2_X1 U12955 ( .A1(n10734), .A2(n10478), .ZN(n10738) );
  NAND2_X2 U12956 ( .A1(n10391), .A2(n15136), .ZN(n15143) );
  INV_X1 U12957 ( .A(n10388), .ZN(n10389) );
  NAND2_X1 U12958 ( .A1(n15143), .A2(n10389), .ZN(n14750) );
  INV_X1 U12959 ( .A(n10391), .ZN(n10394) );
  NAND2_X1 U12960 ( .A1(n14381), .A2(n14213), .ZN(n14459) );
  INV_X1 U12961 ( .A(n14459), .ZN(n10392) );
  NAND2_X1 U12962 ( .A1(n14210), .A2(n10392), .ZN(n14950) );
  INV_X1 U12963 ( .A(n14950), .ZN(n10393) );
  NAND2_X1 U12964 ( .A1(n14393), .A2(n14717), .ZN(n10397) );
  INV_X1 U12965 ( .A(n15143), .ZN(n14931) );
  AOI22_X1 U12966 ( .A1(n14931), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n10395), 
        .B2(n10394), .ZN(n10396) );
  OAI211_X1 U12967 ( .C1(n15136), .C2(n10398), .A(n10397), .B(n10396), .ZN(
        n10399) );
  NOR2_X1 U12968 ( .A1(n10406), .A2(n10405), .ZN(n10503) );
  INV_X1 U12969 ( .A(n10478), .ZN(n10407) );
  INV_X1 U12970 ( .A(n10408), .ZN(n10409) );
  AND2_X4 U12971 ( .A1(n13426), .A2(n10409), .ZN(P3_U3897) );
  NOR2_X1 U12972 ( .A1(n6671), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14080) );
  INV_X1 U12973 ( .A(n14080), .ZN(n14072) );
  NAND2_X1 U12974 ( .A1(n6671), .A2(P2_U3088), .ZN(n14083) );
  INV_X1 U12975 ( .A(n10526), .ZN(n15360) );
  OAI222_X1 U12976 ( .A1(n14072), .A2(n10410), .B1(n14083), .B2(n10440), .C1(
        n15360), .C2(P2_U3088), .ZN(P2_U3324) );
  INV_X1 U12977 ( .A(n10411), .ZN(n10463) );
  INV_X1 U12978 ( .A(n10524), .ZN(n10689) );
  OAI222_X1 U12979 ( .A1(n14072), .A2(n10412), .B1(n14083), .B2(n10463), .C1(
        n10689), .C2(P2_U3088), .ZN(P2_U3325) );
  INV_X1 U12980 ( .A(n10527), .ZN(n15373) );
  OAI222_X1 U12981 ( .A1(n14072), .A2(n10413), .B1(n14083), .B2(n10435), .C1(
        n15373), .C2(P2_U3088), .ZN(P2_U3323) );
  INV_X1 U12982 ( .A(SI_4_), .ZN(n10416) );
  NOR2_X1 U12983 ( .A1(n6671), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13433) );
  INV_X2 U12984 ( .A(n13433), .ZN(n12666) );
  INV_X1 U12985 ( .A(n10414), .ZN(n10415) );
  OAI222_X1 U12986 ( .A1(P3_U3151), .A2(n10937), .B1(n13440), .B2(n10416), 
        .C1(n12666), .C2(n10415), .ZN(P3_U3291) );
  INV_X1 U12987 ( .A(SI_7_), .ZN(n10419) );
  INV_X1 U12988 ( .A(n10417), .ZN(n10418) );
  OAI222_X1 U12989 ( .A1(P3_U3151), .A2(n11327), .B1(n13440), .B2(n10419), 
        .C1(n12666), .C2(n10418), .ZN(P3_U3288) );
  OAI222_X1 U12990 ( .A1(P3_U3151), .A2(n11853), .B1(n13440), .B2(n10421), 
        .C1(n12666), .C2(n10420), .ZN(P3_U3287) );
  INV_X1 U12991 ( .A(n10967), .ZN(n10914) );
  INV_X1 U12992 ( .A(n10422), .ZN(n10423) );
  OAI222_X1 U12993 ( .A1(P3_U3151), .A2(n10914), .B1(n13440), .B2(n10424), 
        .C1(n12666), .C2(n10423), .ZN(P3_U3293) );
  INV_X1 U12994 ( .A(SI_5_), .ZN(n10427) );
  INV_X1 U12995 ( .A(n10425), .ZN(n10426) );
  OAI222_X1 U12996 ( .A1(P3_U3151), .A2(n10995), .B1(n13440), .B2(n10427), 
        .C1(n12666), .C2(n10426), .ZN(P3_U3290) );
  INV_X1 U12997 ( .A(SI_9_), .ZN(n10430) );
  INV_X1 U12998 ( .A(n10428), .ZN(n10429) );
  OAI222_X1 U12999 ( .A1(P3_U3151), .A2(n15557), .B1(n13440), .B2(n10430), 
        .C1(n12666), .C2(n10429), .ZN(P3_U3286) );
  INV_X1 U13000 ( .A(n10542), .ZN(n10533) );
  OAI222_X1 U13001 ( .A1(n14072), .A2(n10431), .B1(n14083), .B2(n10437), .C1(
        n10533), .C2(P2_U3088), .ZN(P2_U3321) );
  NAND2_X1 U13002 ( .A1(n6671), .A2(P1_U3086), .ZN(n14891) );
  CLKBUF_X1 U13003 ( .A(n14891), .Z(n14869) );
  NOR2_X1 U13004 ( .A1(n6671), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14874) );
  INV_X2 U13005 ( .A(n14874), .ZN(n14885) );
  INV_X1 U13006 ( .A(n15231), .ZN(n10434) );
  OAI222_X1 U13007 ( .A1(n14869), .A2(n10436), .B1(n14885), .B2(n10435), .C1(
        n10434), .C2(P1_U3086), .ZN(P1_U3351) );
  INV_X1 U13008 ( .A(n10584), .ZN(n10851) );
  OAI222_X1 U13009 ( .A1(n14869), .A2(n10438), .B1(n14885), .B2(n10437), .C1(
        n10851), .C2(P1_U3086), .ZN(P1_U3349) );
  INV_X1 U13010 ( .A(n14546), .ZN(n10439) );
  OAI222_X1 U13011 ( .A1(n14869), .A2(n10441), .B1(n14885), .B2(n10440), .C1(
        n10439), .C2(P1_U3086), .ZN(P1_U3352) );
  INV_X1 U13012 ( .A(n10442), .ZN(n10467) );
  OAI222_X1 U13013 ( .A1(n14869), .A2(n10443), .B1(n14885), .B2(n10467), .C1(
        n14562), .C2(P1_U3086), .ZN(P1_U3350) );
  OAI222_X1 U13014 ( .A1(n12666), .A2(n10444), .B1(n13440), .B2(n6886), .C1(
        P3_U3151), .C2(n11313), .ZN(P3_U3294) );
  INV_X1 U13015 ( .A(SI_3_), .ZN(n10447) );
  INV_X1 U13016 ( .A(n10445), .ZN(n10446) );
  OAI222_X1 U13017 ( .A1(P3_U3151), .A2(n7299), .B1(n13440), .B2(n10447), .C1(
        n12666), .C2(n10446), .ZN(P3_U3292) );
  OAI222_X1 U13018 ( .A1(P3_U3151), .A2(n13011), .B1(n13440), .B2(n10449), 
        .C1(n12666), .C2(n10448), .ZN(P3_U3285) );
  OAI222_X1 U13019 ( .A1(n15573), .A2(P3_U3151), .B1(n12666), .B2(n10451), 
        .C1(n13440), .C2(n10450), .ZN(P3_U3284) );
  OAI222_X1 U13020 ( .A1(P3_U3151), .A2(n11163), .B1(n12666), .B2(n10453), 
        .C1(n10452), .C2(n13440), .ZN(P3_U3289) );
  OAI222_X1 U13021 ( .A1(P3_U3151), .A2(n7030), .B1(n12666), .B2(n10455), .C1(
        n10454), .C2(n13440), .ZN(P3_U3295) );
  OAI222_X1 U13022 ( .A1(n13440), .A2(n10457), .B1(n12666), .B2(n10456), .C1(
        n15590), .C2(P3_U3151), .ZN(P3_U3283) );
  INV_X1 U13023 ( .A(n10749), .ZN(n10756) );
  OAI222_X1 U13024 ( .A1(n14072), .A2(n10458), .B1(n14083), .B2(n10460), .C1(
        n10756), .C2(P2_U3088), .ZN(P2_U3320) );
  INV_X1 U13025 ( .A(n10596), .ZN(n10459) );
  OAI222_X1 U13026 ( .A1(n14891), .A2(n10461), .B1(n14885), .B2(n10460), .C1(
        n10459), .C2(P1_U3086), .ZN(P1_U3348) );
  INV_X1 U13027 ( .A(n14530), .ZN(n10464) );
  OAI222_X1 U13028 ( .A1(P1_U3086), .A2(n10464), .B1(n14885), .B2(n10463), 
        .C1(n10462), .C2(n14869), .ZN(P1_U3353) );
  OAI222_X1 U13029 ( .A1(P1_U3086), .A2(n14512), .B1(n14885), .B2(n10466), 
        .C1(n7491), .C2(n14869), .ZN(P1_U3354) );
  CLKBUF_X1 U13030 ( .A(n14083), .Z(n14075) );
  AOI22_X1 U13031 ( .A1(n14080), .A2(P1_DATAO_REG_1__SCAN_IN), .B1(n13663), 
        .B2(P2_STATE_REG_SCAN_IN), .ZN(n10465) );
  OAI21_X1 U13032 ( .B1(n10466), .B2(n14075), .A(n10465), .ZN(P2_U3326) );
  INV_X1 U13033 ( .A(n10766), .ZN(n10780) );
  OAI222_X1 U13034 ( .A1(n14072), .A2(n10468), .B1(n14075), .B2(n10467), .C1(
        n10780), .C2(P2_U3088), .ZN(P2_U3322) );
  INV_X1 U13035 ( .A(n10784), .ZN(n10782) );
  OAI222_X1 U13036 ( .A1(n14072), .A2(n10469), .B1(n14075), .B2(n10471), .C1(
        n10782), .C2(P2_U3088), .ZN(P2_U3319) );
  INV_X1 U13037 ( .A(n14576), .ZN(n10470) );
  OAI222_X1 U13038 ( .A1(n14869), .A2(n10472), .B1(n14885), .B2(n10471), .C1(
        n10470), .C2(P1_U3086), .ZN(P1_U3347) );
  INV_X1 U13039 ( .A(n10738), .ZN(n10473) );
  NAND2_X1 U13040 ( .A1(n10474), .A2(n10473), .ZN(n15272) );
  INV_X1 U13041 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n10476) );
  AOI22_X1 U13042 ( .A1(n15272), .A2(n10476), .B1(n10475), .B2(n10478), .ZN(
        P1_U3446) );
  INV_X1 U13043 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n10480) );
  INV_X1 U13044 ( .A(n10477), .ZN(n10479) );
  AOI22_X1 U13045 ( .A1(n15272), .A2(n10480), .B1(n10479), .B2(n10478), .ZN(
        P1_U3445) );
  NAND2_X1 U13046 ( .A1(n9025), .A2(P2_U3947), .ZN(n10481) );
  OAI21_X1 U13047 ( .B1(n9376), .B2(P2_U3947), .A(n10481), .ZN(P2_U3531) );
  INV_X1 U13048 ( .A(n10482), .ZN(n10484) );
  NAND2_X1 U13049 ( .A1(n10484), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14475) );
  NAND2_X1 U13050 ( .A1(n10738), .A2(n14475), .ZN(n10564) );
  OAI21_X1 U13051 ( .B1(n10484), .B2(n14413), .A(n10483), .ZN(n10562) );
  NAND2_X1 U13052 ( .A1(n10564), .A2(n10562), .ZN(n15270) );
  INV_X1 U13053 ( .A(n15270), .ZN(n14593) );
  NOR2_X1 U13054 ( .A1(n14593), .A2(P1_U4016), .ZN(P1_U3085) );
  OAI222_X1 U13055 ( .A1(P3_U3151), .A2(n15605), .B1(n13440), .B2(n10486), 
        .C1(n12666), .C2(n10485), .ZN(P3_U3282) );
  INV_X1 U13056 ( .A(n10487), .ZN(n10489) );
  INV_X1 U13057 ( .A(n14594), .ZN(n14590) );
  OAI222_X1 U13058 ( .A1(n14869), .A2(n10488), .B1(n14885), .B2(n10489), .C1(
        P1_U3086), .C2(n14590), .ZN(P1_U3346) );
  INV_X1 U13059 ( .A(n10794), .ZN(n11070) );
  OAI222_X1 U13060 ( .A1(n14072), .A2(n10490), .B1(n14075), .B2(n10489), .C1(
        P2_U3088), .C2(n11070), .ZN(P2_U3318) );
  INV_X1 U13061 ( .A(n11072), .ZN(n15387) );
  OAI222_X1 U13062 ( .A1(n14072), .A2(n10491), .B1(n14075), .B2(n10492), .C1(
        n15387), .C2(P2_U3088), .ZN(P2_U3317) );
  INV_X1 U13063 ( .A(n10605), .ZN(n10812) );
  OAI222_X1 U13064 ( .A1(n14869), .A2(n10493), .B1(n14885), .B2(n10492), .C1(
        n10812), .C2(P1_U3086), .ZN(P1_U3345) );
  OAI222_X1 U13065 ( .A1(P3_U3151), .A2(n15625), .B1(n13440), .B2(n10495), 
        .C1(n12666), .C2(n10494), .ZN(P3_U3281) );
  INV_X1 U13066 ( .A(n10496), .ZN(n10498) );
  OAI222_X1 U13067 ( .A1(n14869), .A2(n10497), .B1(n14885), .B2(n10498), .C1(
        P1_U3086), .C2(n10890), .ZN(P1_U3344) );
  INV_X1 U13068 ( .A(n11229), .ZN(n11223) );
  OAI222_X1 U13069 ( .A1(n14072), .A2(n10499), .B1(n14075), .B2(n10498), .C1(
        P2_U3088), .C2(n11223), .ZN(P2_U3316) );
  AOI21_X1 U13070 ( .B1(n10501), .B2(n10500), .A(n7821), .ZN(n10502) );
  OR2_X1 U13071 ( .A1(n10503), .A2(n10502), .ZN(n10507) );
  INV_X1 U13072 ( .A(n10505), .ZN(n10504) );
  AND2_X1 U13073 ( .A1(n10507), .A2(n10504), .ZN(n15359) );
  INV_X1 U13074 ( .A(n15453), .ZN(n15401) );
  NOR2_X2 U13075 ( .A1(n10507), .A2(P2_U3088), .ZN(n15448) );
  NAND2_X1 U13076 ( .A1(P2_U3088), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n11427) );
  INV_X1 U13077 ( .A(n11427), .ZN(n10522) );
  NAND2_X1 U13078 ( .A1(n10505), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14077) );
  INV_X1 U13079 ( .A(n14077), .ZN(n10506) );
  AND2_X1 U13080 ( .A1(n10507), .A2(n10506), .ZN(n10523) );
  INV_X1 U13081 ( .A(n14081), .ZN(n10508) );
  NAND2_X1 U13082 ( .A1(n10523), .A2(n10508), .ZN(n15375) );
  INV_X1 U13083 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10509) );
  MUX2_X1 U13084 ( .A(n10509), .B(P2_REG1_REG_2__SCAN_IN), .S(n10524), .Z(
        n10679) );
  INV_X1 U13085 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10510) );
  MUX2_X1 U13086 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n10510), .S(n13663), .Z(
        n10512) );
  AND2_X1 U13087 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n10511) );
  NAND2_X1 U13088 ( .A1(n10512), .A2(n10511), .ZN(n13667) );
  NAND2_X1 U13089 ( .A1(n13663), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n10513) );
  AND2_X1 U13090 ( .A1(n13667), .A2(n10513), .ZN(n10680) );
  NOR2_X1 U13091 ( .A1(n10679), .A2(n10680), .ZN(n10678) );
  AOI21_X1 U13092 ( .B1(P2_REG1_REG_2__SCAN_IN), .B2(n10524), .A(n10678), .ZN(
        n15367) );
  INV_X1 U13093 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10514) );
  MUX2_X1 U13094 ( .A(n10514), .B(P2_REG1_REG_3__SCAN_IN), .S(n10526), .Z(
        n15366) );
  NOR2_X1 U13095 ( .A1(n15367), .A2(n15366), .ZN(n15365) );
  AOI21_X1 U13096 ( .B1(n10526), .B2(P2_REG1_REG_3__SCAN_IN), .A(n15365), .ZN(
        n15378) );
  INV_X1 U13097 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10515) );
  MUX2_X1 U13098 ( .A(n10515), .B(P2_REG1_REG_4__SCAN_IN), .S(n10527), .Z(
        n15377) );
  NOR2_X1 U13099 ( .A1(n15378), .A2(n15377), .ZN(n15376) );
  NOR2_X1 U13100 ( .A1(n15373), .A2(n10515), .ZN(n10765) );
  INV_X1 U13101 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10516) );
  MUX2_X1 U13102 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n10516), .S(n10766), .Z(
        n10517) );
  OAI21_X1 U13103 ( .B1(n15376), .B2(n10765), .A(n10517), .ZN(n10769) );
  NAND2_X1 U13104 ( .A1(n10766), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n10519) );
  INV_X1 U13105 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n15528) );
  MUX2_X1 U13106 ( .A(n15528), .B(P2_REG1_REG_6__SCAN_IN), .S(n10542), .Z(
        n10518) );
  AOI21_X1 U13107 ( .B1(n10769), .B2(n10519), .A(n10518), .ZN(n10537) );
  AND3_X1 U13108 ( .A1(n10769), .A2(n10519), .A3(n10518), .ZN(n10520) );
  NOR3_X1 U13109 ( .A1(n15375), .A2(n10537), .A3(n10520), .ZN(n10521) );
  AOI211_X1 U13110 ( .C1(n15448), .C2(P2_ADDR_REG_6__SCAN_IN), .A(n10522), .B(
        n10521), .ZN(n10532) );
  MUX2_X1 U13111 ( .A(n13935), .B(P2_REG2_REG_1__SCAN_IN), .S(n13663), .Z(
        n13661) );
  AOI21_X1 U13112 ( .B1(n13663), .B2(P2_REG2_REG_1__SCAN_IN), .A(n13659), .ZN(
        n10684) );
  MUX2_X1 U13113 ( .A(n10525), .B(P2_REG2_REG_2__SCAN_IN), .S(n10524), .Z(
        n10683) );
  OR2_X1 U13114 ( .A1(n10684), .A2(n10683), .ZN(n10686) );
  OAI21_X1 U13115 ( .B1(n10525), .B2(n10689), .A(n10686), .ZN(n15364) );
  MUX2_X1 U13116 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n11396), .S(n10526), .Z(
        n15363) );
  NAND2_X1 U13117 ( .A1(n15364), .A2(n15363), .ZN(n15362) );
  OAI21_X1 U13118 ( .B1(n11396), .B2(n15360), .A(n15362), .ZN(n15382) );
  MUX2_X1 U13119 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n11407), .S(n10527), .Z(
        n15381) );
  NAND2_X1 U13120 ( .A1(n15382), .A2(n15381), .ZN(n15380) );
  NAND2_X1 U13121 ( .A1(n10527), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n10775) );
  MUX2_X1 U13122 ( .A(n7806), .B(P2_REG2_REG_5__SCAN_IN), .S(n10766), .Z(
        n10774) );
  NOR2_X1 U13123 ( .A1(n10780), .A2(n7806), .ZN(n10529) );
  MUX2_X1 U13124 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n11582), .S(n10542), .Z(
        n10528) );
  OAI21_X1 U13125 ( .B1(n10773), .B2(n10529), .A(n10528), .ZN(n10545) );
  OR3_X1 U13126 ( .A1(n10773), .A2(n10529), .A3(n10528), .ZN(n10530) );
  NAND3_X1 U13127 ( .A1(n15450), .A2(n10545), .A3(n10530), .ZN(n10531) );
  OAI211_X1 U13128 ( .C1(n15401), .C2(n10533), .A(n10532), .B(n10531), .ZN(
        P2_U3220) );
  NAND2_X1 U13129 ( .A1(P2_U3088), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n11509) );
  INV_X1 U13130 ( .A(n11509), .ZN(n10541) );
  NOR2_X1 U13131 ( .A1(n10533), .A2(n15528), .ZN(n10536) );
  INV_X1 U13132 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n10534) );
  MUX2_X1 U13133 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n10534), .S(n10749), .Z(
        n10535) );
  OAI21_X1 U13134 ( .B1(n10537), .B2(n10536), .A(n10535), .ZN(n10752) );
  INV_X1 U13135 ( .A(n10752), .ZN(n10539) );
  NOR3_X1 U13136 ( .A1(n10537), .A2(n10536), .A3(n10535), .ZN(n10538) );
  NOR3_X1 U13137 ( .A1(n10539), .A2(n10538), .A3(n15375), .ZN(n10540) );
  AOI211_X1 U13138 ( .C1(n15448), .C2(P2_ADDR_REG_7__SCAN_IN), .A(n10541), .B(
        n10540), .ZN(n10549) );
  NAND2_X1 U13139 ( .A1(n10542), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n10544) );
  INV_X1 U13140 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n10755) );
  MUX2_X1 U13141 ( .A(n10755), .B(P2_REG2_REG_7__SCAN_IN), .S(n10749), .Z(
        n10543) );
  AOI21_X1 U13142 ( .B1(n10545), .B2(n10544), .A(n10543), .ZN(n10760) );
  INV_X1 U13143 ( .A(n10760), .ZN(n10547) );
  NAND3_X1 U13144 ( .A1(n10545), .A2(n10544), .A3(n10543), .ZN(n10546) );
  NAND3_X1 U13145 ( .A1(n15450), .A2(n10547), .A3(n10546), .ZN(n10548) );
  OAI211_X1 U13146 ( .C1(n15401), .C2(n10756), .A(n10549), .B(n10548), .ZN(
        P2_U3221) );
  INV_X1 U13147 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n15345) );
  MUX2_X1 U13148 ( .A(n15345), .B(P1_REG1_REG_5__SCAN_IN), .S(n14562), .Z(
        n14560) );
  INV_X1 U13149 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10550) );
  MUX2_X1 U13150 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n10550), .S(n14530), .Z(
        n10553) );
  INV_X1 U13151 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10551) );
  MUX2_X1 U13152 ( .A(n10551), .B(P1_REG1_REG_1__SCAN_IN), .S(n14512), .Z(
        n14510) );
  AND2_X1 U13153 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n14511) );
  NAND2_X1 U13154 ( .A1(n14510), .A2(n14511), .ZN(n14527) );
  OR2_X1 U13155 ( .A1(n14512), .A2(n10551), .ZN(n14526) );
  NAND2_X1 U13156 ( .A1(n14527), .A2(n14526), .ZN(n10552) );
  NAND2_X1 U13157 ( .A1(n10553), .A2(n10552), .ZN(n14544) );
  NAND2_X1 U13158 ( .A1(n14530), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n14542) );
  NAND2_X1 U13159 ( .A1(n14544), .A2(n14542), .ZN(n10556) );
  INV_X1 U13160 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n10554) );
  MUX2_X1 U13161 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n10554), .S(n14546), .Z(
        n10555) );
  NAND2_X1 U13162 ( .A1(n10556), .A2(n10555), .ZN(n15223) );
  NAND2_X1 U13163 ( .A1(n14546), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n15222) );
  NAND2_X1 U13164 ( .A1(n15223), .A2(n15222), .ZN(n10559) );
  INV_X1 U13165 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n10557) );
  MUX2_X1 U13166 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n10557), .S(n15231), .Z(
        n10558) );
  NAND2_X1 U13167 ( .A1(n10559), .A2(n10558), .ZN(n15225) );
  NAND2_X1 U13168 ( .A1(n15231), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n10560) );
  AND2_X1 U13169 ( .A1(n15225), .A2(n10560), .ZN(n14559) );
  NAND2_X1 U13170 ( .A1(n14560), .A2(n14559), .ZN(n14558) );
  NAND2_X1 U13171 ( .A1(n14562), .A2(n15345), .ZN(n10561) );
  NAND2_X1 U13172 ( .A1(n14558), .A2(n10561), .ZN(n10847) );
  INV_X1 U13173 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n15347) );
  MUX2_X1 U13174 ( .A(n15347), .B(P1_REG1_REG_6__SCAN_IN), .S(n10584), .Z(
        n10846) );
  OR2_X1 U13175 ( .A1(n10847), .A2(n10846), .ZN(n10844) );
  NAND2_X1 U13176 ( .A1(n10584), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n10567) );
  INV_X1 U13177 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n15349) );
  MUX2_X1 U13178 ( .A(n15349), .B(P1_REG1_REG_7__SCAN_IN), .S(n10596), .Z(
        n10566) );
  AOI21_X1 U13179 ( .B1(n10844), .B2(n10567), .A(n10566), .ZN(n10595) );
  INV_X1 U13180 ( .A(n10562), .ZN(n10563) );
  NAND2_X1 U13181 ( .A1(n10564), .A2(n10563), .ZN(n10698) );
  INV_X1 U13182 ( .A(n10698), .ZN(n10565) );
  NAND3_X1 U13183 ( .A1(n10844), .A2(n10567), .A3(n10566), .ZN(n10568) );
  NAND2_X1 U13184 ( .A1(n15261), .A2(n10568), .ZN(n10592) );
  INV_X1 U13185 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n10569) );
  NAND2_X1 U13186 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n12130) );
  OAI21_X1 U13187 ( .B1(n15270), .B2(n10569), .A(n12130), .ZN(n10570) );
  AOI21_X1 U13188 ( .B1(n10596), .B2(n15232), .A(n10570), .ZN(n10591) );
  OR3_X1 U13189 ( .A1(n10698), .A2(n6676), .A3(n12662), .ZN(n15248) );
  INV_X1 U13190 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n11470) );
  MUX2_X1 U13191 ( .A(n11470), .B(P1_REG2_REG_5__SCAN_IN), .S(n14562), .Z(
        n10581) );
  INV_X1 U13192 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n14531) );
  MUX2_X1 U13193 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n14531), .S(n14530), .Z(
        n10574) );
  INV_X1 U13194 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n10571) );
  MUX2_X1 U13195 ( .A(n10571), .B(P1_REG2_REG_1__SCAN_IN), .S(n14512), .Z(
        n10572) );
  AND2_X1 U13196 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n14519) );
  NAND2_X1 U13197 ( .A1(n10572), .A2(n14519), .ZN(n14533) );
  OR2_X1 U13198 ( .A1(n14512), .A2(n10571), .ZN(n14532) );
  NAND2_X1 U13199 ( .A1(n14533), .A2(n14532), .ZN(n10573) );
  NAND2_X1 U13200 ( .A1(n10574), .A2(n10573), .ZN(n14549) );
  NAND2_X1 U13201 ( .A1(n14530), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n14547) );
  NAND2_X1 U13202 ( .A1(n14549), .A2(n14547), .ZN(n10576) );
  INV_X1 U13203 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n11140) );
  MUX2_X1 U13204 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n11140), .S(n14546), .Z(
        n10575) );
  NAND2_X1 U13205 ( .A1(n10576), .A2(n10575), .ZN(n15228) );
  NAND2_X1 U13206 ( .A1(n14546), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n15227) );
  NAND2_X1 U13207 ( .A1(n15228), .A2(n15227), .ZN(n10579) );
  INV_X1 U13208 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n10577) );
  MUX2_X1 U13209 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n10577), .S(n15231), .Z(
        n10578) );
  NAND2_X1 U13210 ( .A1(n10579), .A2(n10578), .ZN(n15230) );
  NAND2_X1 U13211 ( .A1(n15231), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n14563) );
  NAND2_X1 U13212 ( .A1(n15230), .A2(n14563), .ZN(n10580) );
  NAND2_X1 U13213 ( .A1(n10581), .A2(n10580), .ZN(n14566) );
  NAND2_X1 U13214 ( .A1(n14557), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n10582) );
  NAND2_X1 U13215 ( .A1(n14566), .A2(n10582), .ZN(n10842) );
  INV_X1 U13216 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n10583) );
  MUX2_X1 U13217 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n10583), .S(n10584), .Z(
        n10841) );
  NAND2_X1 U13218 ( .A1(n10842), .A2(n10841), .ZN(n10840) );
  NAND2_X1 U13219 ( .A1(n10584), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n10588) );
  NAND2_X1 U13220 ( .A1(n10840), .A2(n10588), .ZN(n10586) );
  INV_X1 U13221 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n11484) );
  MUX2_X1 U13222 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n11484), .S(n10596), .Z(
        n10585) );
  NAND2_X1 U13223 ( .A1(n10586), .A2(n10585), .ZN(n14579) );
  MUX2_X1 U13224 ( .A(n11484), .B(P1_REG2_REG_7__SCAN_IN), .S(n10596), .Z(
        n10587) );
  NAND3_X1 U13225 ( .A1(n10840), .A2(n10588), .A3(n10587), .ZN(n10589) );
  NAND3_X1 U13226 ( .A1(n15258), .A2(n14579), .A3(n10589), .ZN(n10590) );
  OAI211_X1 U13227 ( .C1(n10595), .C2(n10592), .A(n10591), .B(n10590), .ZN(
        P1_U3250) );
  INV_X1 U13228 ( .A(n13058), .ZN(n14974) );
  OAI222_X1 U13229 ( .A1(P3_U3151), .A2(n14974), .B1(n13440), .B2(n10594), 
        .C1(n12666), .C2(n10593), .ZN(P3_U3280) );
  AOI21_X1 U13230 ( .B1(n10596), .B2(P1_REG1_REG_7__SCAN_IN), .A(n10595), .ZN(
        n14571) );
  INV_X1 U13231 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n15351) );
  MUX2_X1 U13232 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n15351), .S(n14576), .Z(
        n14570) );
  AND2_X1 U13233 ( .A1(n14571), .A2(n14570), .ZN(n14587) );
  NOR2_X1 U13234 ( .A1(n14576), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n14585) );
  INV_X1 U13235 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n15353) );
  MUX2_X1 U13236 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n15353), .S(n14594), .Z(
        n14586) );
  OAI21_X1 U13237 ( .B1(n14587), .B2(n14585), .A(n14586), .ZN(n14584) );
  OAI21_X1 U13238 ( .B1(n14594), .B2(P1_REG1_REG_9__SCAN_IN), .A(n14584), .ZN(
        n10803) );
  INV_X1 U13239 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n15356) );
  MUX2_X1 U13240 ( .A(n15356), .B(P1_REG1_REG_10__SCAN_IN), .S(n10605), .Z(
        n10802) );
  NOR2_X1 U13241 ( .A1(n10803), .A2(n10802), .ZN(n10801) );
  AOI21_X1 U13242 ( .B1(n10605), .B2(P1_REG1_REG_10__SCAN_IN), .A(n10801), 
        .ZN(n10618) );
  INV_X1 U13243 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n15185) );
  INV_X1 U13244 ( .A(n15261), .ZN(n15243) );
  NOR3_X1 U13245 ( .A1(n10618), .A2(n15185), .A3(n15243), .ZN(n10608) );
  NAND2_X1 U13246 ( .A1(n10596), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n14578) );
  NAND2_X1 U13247 ( .A1(n14579), .A2(n14578), .ZN(n10599) );
  INV_X1 U13248 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n10597) );
  MUX2_X1 U13249 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n10597), .S(n14576), .Z(
        n10598) );
  NAND2_X1 U13250 ( .A1(n10599), .A2(n10598), .ZN(n14597) );
  NAND2_X1 U13251 ( .A1(n14576), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n14596) );
  NAND2_X1 U13252 ( .A1(n14597), .A2(n14596), .ZN(n10602) );
  INV_X1 U13253 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n10600) );
  MUX2_X1 U13254 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n10600), .S(n14594), .Z(
        n10601) );
  NAND2_X1 U13255 ( .A1(n10602), .A2(n10601), .ZN(n14599) );
  NAND2_X1 U13256 ( .A1(n14594), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n10603) );
  NAND2_X1 U13257 ( .A1(n14599), .A2(n10603), .ZN(n10807) );
  INV_X1 U13258 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n10604) );
  MUX2_X1 U13259 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n10604), .S(n10605), .Z(
        n10806) );
  NAND2_X1 U13260 ( .A1(n10807), .A2(n10806), .ZN(n10805) );
  NAND2_X1 U13261 ( .A1(n10605), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n10606) );
  NAND2_X1 U13262 ( .A1(n10805), .A2(n10606), .ZN(n10612) );
  NOR3_X1 U13263 ( .A1(n10612), .A2(P1_REG2_REG_11__SCAN_IN), .A3(n15248), 
        .ZN(n10607) );
  NOR3_X1 U13264 ( .A1(n10608), .A2(n15232), .A3(n10607), .ZN(n10622) );
  AOI21_X1 U13265 ( .B1(n10890), .B2(P1_REG2_REG_11__SCAN_IN), .A(n10612), 
        .ZN(n10609) );
  NOR2_X1 U13266 ( .A1(n10609), .A2(n15248), .ZN(n10615) );
  INV_X1 U13267 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n10610) );
  MUX2_X1 U13268 ( .A(n10610), .B(P1_REG2_REG_11__SCAN_IN), .S(n10890), .Z(
        n10611) );
  NAND2_X1 U13269 ( .A1(n10612), .A2(n10611), .ZN(n10881) );
  NAND2_X1 U13270 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n12490)
         );
  OAI21_X1 U13271 ( .B1(n15270), .B2(n10613), .A(n12490), .ZN(n10614) );
  AOI21_X1 U13272 ( .B1(n10615), .B2(n10881), .A(n10614), .ZN(n10621) );
  INV_X1 U13273 ( .A(n10890), .ZN(n10616) );
  NOR3_X1 U13274 ( .A1(n10618), .A2(P1_REG1_REG_11__SCAN_IN), .A3(n10616), 
        .ZN(n10619) );
  MUX2_X1 U13275 ( .A(n15185), .B(P1_REG1_REG_11__SCAN_IN), .S(n10890), .Z(
        n10617) );
  OAI21_X1 U13276 ( .B1(n10619), .B2(n10889), .A(n15261), .ZN(n10620) );
  OAI211_X1 U13277 ( .C1(n10622), .C2(n10890), .A(n10621), .B(n10620), .ZN(
        P1_U3254) );
  INV_X1 U13278 ( .A(n13426), .ZN(n10624) );
  NOR2_X1 U13279 ( .A1(n10624), .A2(n10623), .ZN(n10626) );
  CLKBUF_X1 U13280 ( .A(n10626), .Z(n10656) );
  INV_X1 U13281 ( .A(P3_D_REG_8__SCAN_IN), .ZN(n10625) );
  NOR2_X1 U13282 ( .A1(n10656), .A2(n10625), .ZN(P3_U3257) );
  INV_X1 U13283 ( .A(P3_D_REG_5__SCAN_IN), .ZN(n10627) );
  NOR2_X1 U13284 ( .A1(n10656), .A2(n10627), .ZN(P3_U3260) );
  INV_X1 U13285 ( .A(P3_D_REG_11__SCAN_IN), .ZN(n10628) );
  NOR2_X1 U13286 ( .A1(n10656), .A2(n10628), .ZN(P3_U3254) );
  INV_X1 U13287 ( .A(P3_D_REG_6__SCAN_IN), .ZN(n10629) );
  NOR2_X1 U13288 ( .A1(n10656), .A2(n10629), .ZN(P3_U3259) );
  INV_X1 U13289 ( .A(P3_D_REG_2__SCAN_IN), .ZN(n10630) );
  NOR2_X1 U13290 ( .A1(n10656), .A2(n10630), .ZN(P3_U3263) );
  INV_X1 U13291 ( .A(P3_D_REG_23__SCAN_IN), .ZN(n10631) );
  NOR2_X1 U13292 ( .A1(n10626), .A2(n10631), .ZN(P3_U3242) );
  INV_X1 U13293 ( .A(P3_D_REG_7__SCAN_IN), .ZN(n10632) );
  NOR2_X1 U13294 ( .A1(n10626), .A2(n10632), .ZN(P3_U3258) );
  INV_X1 U13295 ( .A(P3_D_REG_21__SCAN_IN), .ZN(n10633) );
  NOR2_X1 U13296 ( .A1(n10626), .A2(n10633), .ZN(P3_U3244) );
  INV_X1 U13297 ( .A(P3_D_REG_20__SCAN_IN), .ZN(n10634) );
  NOR2_X1 U13298 ( .A1(n10626), .A2(n10634), .ZN(P3_U3245) );
  INV_X1 U13299 ( .A(P3_D_REG_19__SCAN_IN), .ZN(n10635) );
  NOR2_X1 U13300 ( .A1(n10656), .A2(n10635), .ZN(P3_U3246) );
  INV_X1 U13301 ( .A(P3_D_REG_3__SCAN_IN), .ZN(n10636) );
  NOR2_X1 U13302 ( .A1(n10626), .A2(n10636), .ZN(P3_U3262) );
  INV_X1 U13303 ( .A(P3_D_REG_17__SCAN_IN), .ZN(n10637) );
  NOR2_X1 U13304 ( .A1(n10656), .A2(n10637), .ZN(P3_U3248) );
  INV_X1 U13305 ( .A(P3_D_REG_16__SCAN_IN), .ZN(n10638) );
  NOR2_X1 U13306 ( .A1(n10656), .A2(n10638), .ZN(P3_U3249) );
  INV_X1 U13307 ( .A(P3_D_REG_15__SCAN_IN), .ZN(n10639) );
  NOR2_X1 U13308 ( .A1(n10656), .A2(n10639), .ZN(P3_U3250) );
  INV_X1 U13309 ( .A(P3_D_REG_31__SCAN_IN), .ZN(n10640) );
  NOR2_X1 U13310 ( .A1(n10626), .A2(n10640), .ZN(P3_U3234) );
  INV_X1 U13311 ( .A(P3_D_REG_30__SCAN_IN), .ZN(n10641) );
  NOR2_X1 U13312 ( .A1(n10626), .A2(n10641), .ZN(P3_U3235) );
  INV_X1 U13313 ( .A(P3_D_REG_29__SCAN_IN), .ZN(n10642) );
  NOR2_X1 U13314 ( .A1(n10626), .A2(n10642), .ZN(P3_U3236) );
  INV_X1 U13315 ( .A(P3_D_REG_28__SCAN_IN), .ZN(n10643) );
  NOR2_X1 U13316 ( .A1(n10626), .A2(n10643), .ZN(P3_U3237) );
  INV_X1 U13317 ( .A(P3_D_REG_27__SCAN_IN), .ZN(n10644) );
  NOR2_X1 U13318 ( .A1(n10626), .A2(n10644), .ZN(P3_U3238) );
  INV_X1 U13319 ( .A(P3_D_REG_26__SCAN_IN), .ZN(n10645) );
  NOR2_X1 U13320 ( .A1(n10626), .A2(n10645), .ZN(P3_U3239) );
  INV_X1 U13321 ( .A(P3_D_REG_25__SCAN_IN), .ZN(n10646) );
  NOR2_X1 U13322 ( .A1(n10656), .A2(n10646), .ZN(P3_U3240) );
  INV_X1 U13323 ( .A(P3_D_REG_24__SCAN_IN), .ZN(n10647) );
  NOR2_X1 U13324 ( .A1(n10656), .A2(n10647), .ZN(P3_U3241) );
  INV_X1 U13325 ( .A(P3_D_REG_9__SCAN_IN), .ZN(n10648) );
  NOR2_X1 U13326 ( .A1(n10656), .A2(n10648), .ZN(P3_U3256) );
  INV_X1 U13327 ( .A(P3_D_REG_12__SCAN_IN), .ZN(n10649) );
  NOR2_X1 U13328 ( .A1(n10656), .A2(n10649), .ZN(P3_U3253) );
  INV_X1 U13329 ( .A(P3_D_REG_4__SCAN_IN), .ZN(n10650) );
  NOR2_X1 U13330 ( .A1(n10656), .A2(n10650), .ZN(P3_U3261) );
  INV_X1 U13331 ( .A(P3_D_REG_13__SCAN_IN), .ZN(n10651) );
  NOR2_X1 U13332 ( .A1(n10656), .A2(n10651), .ZN(P3_U3252) );
  INV_X1 U13333 ( .A(P3_D_REG_10__SCAN_IN), .ZN(n10652) );
  NOR2_X1 U13334 ( .A1(n10656), .A2(n10652), .ZN(P3_U3255) );
  INV_X1 U13335 ( .A(P3_D_REG_18__SCAN_IN), .ZN(n10653) );
  NOR2_X1 U13336 ( .A1(n10656), .A2(n10653), .ZN(P3_U3247) );
  INV_X1 U13337 ( .A(P3_D_REG_22__SCAN_IN), .ZN(n10654) );
  NOR2_X1 U13338 ( .A1(n10656), .A2(n10654), .ZN(P3_U3243) );
  INV_X1 U13339 ( .A(P3_D_REG_14__SCAN_IN), .ZN(n10655) );
  NOR2_X1 U13340 ( .A1(n10656), .A2(n10655), .ZN(P3_U3251) );
  NAND2_X1 U13341 ( .A1(P3_U3897), .A2(n11673), .ZN(n10657) );
  OAI21_X1 U13342 ( .B1(P3_U3897), .B2(n10658), .A(n10657), .ZN(P3_U3495) );
  NAND2_X1 U13343 ( .A1(P3_U3897), .A2(n15639), .ZN(n10659) );
  OAI21_X1 U13344 ( .B1(P3_U3897), .B2(n10660), .A(n10659), .ZN(P3_U3500) );
  NAND2_X1 U13345 ( .A1(P3_U3897), .A2(n15042), .ZN(n10661) );
  OAI21_X1 U13346 ( .B1(P3_U3897), .B2(n10662), .A(n10661), .ZN(P3_U3503) );
  NAND2_X1 U13347 ( .A1(P3_U3897), .A2(n12438), .ZN(n10663) );
  OAI21_X1 U13348 ( .B1(P3_U3897), .B2(n10664), .A(n10663), .ZN(P3_U3505) );
  NAND2_X1 U13349 ( .A1(P3_U3897), .A2(n11947), .ZN(n10665) );
  OAI21_X1 U13350 ( .B1(P3_U3897), .B2(n10666), .A(n10665), .ZN(P3_U3497) );
  NAND2_X1 U13351 ( .A1(P3_U3897), .A2(n12031), .ZN(n10667) );
  OAI21_X1 U13352 ( .B1(P3_U3897), .B2(n10668), .A(n10667), .ZN(P3_U3498) );
  NAND2_X1 U13353 ( .A1(P3_U3897), .A2(n12189), .ZN(n10669) );
  OAI21_X1 U13354 ( .B1(P3_U3897), .B2(n10670), .A(n10669), .ZN(P3_U3499) );
  NAND2_X1 U13355 ( .A1(P3_U3897), .A2(n13292), .ZN(n10671) );
  OAI21_X1 U13356 ( .B1(P3_U3897), .B2(n10672), .A(n10671), .ZN(P3_U3504) );
  INV_X1 U13357 ( .A(P3_DATAO_REG_15__SCAN_IN), .ZN(n10674) );
  NAND2_X1 U13358 ( .A1(P3_U3897), .A2(n13291), .ZN(n10673) );
  OAI21_X1 U13359 ( .B1(P3_U3897), .B2(n10674), .A(n10673), .ZN(P3_U3506) );
  NAND2_X1 U13360 ( .A1(P3_U3897), .A2(n10675), .ZN(n10676) );
  OAI21_X1 U13361 ( .B1(P3_U3897), .B2(n10677), .A(n10676), .ZN(P3_U3507) );
  INV_X1 U13362 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n11550) );
  NOR2_X1 U13363 ( .A1(n11550), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10682) );
  AOI211_X1 U13364 ( .C1(n10680), .C2(n10679), .A(n10678), .B(n15375), .ZN(
        n10681) );
  AOI211_X1 U13365 ( .C1(n15448), .C2(P2_ADDR_REG_2__SCAN_IN), .A(n10682), .B(
        n10681), .ZN(n10688) );
  NAND2_X1 U13366 ( .A1(n10684), .A2(n10683), .ZN(n10685) );
  NAND3_X1 U13367 ( .A1(n15450), .A2(n10686), .A3(n10685), .ZN(n10687) );
  OAI211_X1 U13368 ( .C1(n15401), .C2(n10689), .A(n10688), .B(n10687), .ZN(
        P2_U3216) );
  NAND2_X1 U13369 ( .A1(P3_U3897), .A2(n15682), .ZN(n10690) );
  OAI21_X1 U13370 ( .B1(P3_U3897), .B2(n10691), .A(n10690), .ZN(P3_U3492) );
  NAND2_X1 U13371 ( .A1(n13219), .A2(P3_U3897), .ZN(n10692) );
  OAI21_X1 U13372 ( .B1(P3_U3897), .B2(n10693), .A(n10692), .ZN(P3_U3509) );
  INV_X1 U13373 ( .A(n6676), .ZN(n10695) );
  NOR2_X1 U13374 ( .A1(n6676), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n10694) );
  NOR2_X1 U13375 ( .A1(n12662), .A2(n10694), .ZN(n14523) );
  OAI21_X1 U13376 ( .B1(n10695), .B2(P1_REG1_REG_0__SCAN_IN), .A(n14523), .ZN(
        n10696) );
  MUX2_X1 U13377 ( .A(n10696), .B(n14523), .S(P1_IR_REG_0__SCAN_IN), .Z(n10697) );
  INV_X1 U13378 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n11289) );
  OAI22_X1 U13379 ( .A1(n10698), .A2(n10697), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n11289), .ZN(n10701) );
  INV_X1 U13380 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n10699) );
  NOR3_X1 U13381 ( .A1(n15243), .A2(P1_REG1_REG_0__SCAN_IN), .A3(n10699), .ZN(
        n10700) );
  AOI211_X1 U13382 ( .C1(n14593), .C2(P1_ADDR_REG_0__SCAN_IN), .A(n10701), .B(
        n10700), .ZN(n10702) );
  INV_X1 U13383 ( .A(n10702), .ZN(P1_U3243) );
  INV_X1 U13384 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n10707) );
  INV_X1 U13385 ( .A(n10703), .ZN(n10705) );
  INV_X1 U13386 ( .A(n11181), .ZN(n14505) );
  INV_X1 U13387 ( .A(n14219), .ZN(n14419) );
  OAI21_X1 U13388 ( .B1(n15337), .B2(n15160), .A(n14419), .ZN(n10704) );
  NAND2_X1 U13389 ( .A1(n6847), .A2(n15134), .ZN(n11290) );
  OAI211_X1 U13390 ( .C1(n10705), .C2(n11294), .A(n10704), .B(n11290), .ZN(
        n14854) );
  NAND2_X1 U13391 ( .A1(n15341), .A2(n14854), .ZN(n10706) );
  OAI21_X1 U13392 ( .B1(n15341), .B2(n10707), .A(n10706), .ZN(P1_U3459) );
  NAND2_X1 U13393 ( .A1(n13235), .A2(P3_U3897), .ZN(n10708) );
  OAI21_X1 U13394 ( .B1(P3_U3897), .B2(n10709), .A(n10708), .ZN(P3_U3510) );
  INV_X1 U13395 ( .A(n14990), .ZN(n13047) );
  OAI222_X1 U13396 ( .A1(P3_U3151), .A2(n13047), .B1(n13440), .B2(n10711), 
        .C1(n12666), .C2(n10710), .ZN(P3_U3279) );
  NAND2_X1 U13397 ( .A1(n15450), .A2(n10712), .ZN(n10713) );
  OAI211_X1 U13398 ( .C1(P2_REG1_REG_0__SCAN_IN), .C2(n15375), .A(n15401), .B(
        n10713), .ZN(n10714) );
  INV_X1 U13399 ( .A(n10714), .ZN(n10716) );
  INV_X1 U13400 ( .A(n15375), .ZN(n15456) );
  AOI22_X1 U13401 ( .A1(n15456), .A2(P2_REG1_REG_0__SCAN_IN), .B1(n15450), 
        .B2(P2_REG2_REG_0__SCAN_IN), .ZN(n10715) );
  MUX2_X1 U13402 ( .A(n10716), .B(n10715), .S(n13665), .Z(n10718) );
  AOI22_X1 U13403 ( .A1(n15448), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3088), .ZN(n10717) );
  NAND2_X1 U13404 ( .A1(n10718), .A2(n10717), .ZN(P2_U3214) );
  NAND2_X1 U13405 ( .A1(n10719), .A2(n11096), .ZN(n10724) );
  NAND2_X1 U13406 ( .A1(n10724), .A2(n10720), .ZN(n10723) );
  INV_X1 U13407 ( .A(n10721), .ZN(n10722) );
  NAND2_X1 U13408 ( .A1(n10723), .A2(n10722), .ZN(n11200) );
  OR2_X1 U13409 ( .A1(n11200), .A2(P1_U3086), .ZN(n11021) );
  INV_X1 U13410 ( .A(n11021), .ZN(n10744) );
  INV_X1 U13411 ( .A(n10724), .ZN(n10741) );
  AND2_X1 U13412 ( .A1(n14195), .A2(n15134), .ZN(n15107) );
  NOR2_X1 U13413 ( .A1(n10738), .A2(n14950), .ZN(n10725) );
  NAND2_X1 U13414 ( .A1(n10741), .A2(n10725), .ZN(n10726) );
  NAND2_X4 U13415 ( .A1(n10734), .A2(n10727), .ZN(n12648) );
  NAND2_X1 U13416 ( .A1(n10728), .A2(n6808), .ZN(n10732) );
  INV_X1 U13417 ( .A(n10734), .ZN(n10729) );
  AOI22_X1 U13418 ( .A1(n11192), .A2(n10730), .B1(n10729), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n10731) );
  INV_X1 U13419 ( .A(n11192), .ZN(n10816) );
  NOR2_X1 U13420 ( .A1(n11181), .A2(n10816), .ZN(n10736) );
  INV_X1 U13421 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n10733) );
  OAI22_X1 U13422 ( .A1(n12648), .A2(n11294), .B1(n10734), .B2(n10733), .ZN(
        n10735) );
  NOR2_X1 U13423 ( .A1(n10814), .A2(n10737), .ZN(n14518) );
  NAND2_X1 U13424 ( .A1(n15334), .A2(n14413), .ZN(n10739) );
  NOR2_X1 U13425 ( .A1(n10739), .A2(n10738), .ZN(n10740) );
  OAI22_X1 U13426 ( .A1(n15111), .A2(n11294), .B1(n14518), .B2(n15092), .ZN(
        n10742) );
  AOI21_X1 U13427 ( .B1(n15107), .B2(n6847), .A(n10742), .ZN(n10743) );
  OAI21_X1 U13428 ( .B1(n10744), .B2(n11289), .A(n10743), .ZN(P1_U3232) );
  INV_X1 U13429 ( .A(n13674), .ZN(n13688) );
  INV_X1 U13430 ( .A(n10745), .ZN(n10747) );
  OAI222_X1 U13431 ( .A1(P2_U3088), .A2(n13688), .B1(n14075), .B2(n10747), 
        .C1(n10746), .C2(n14072), .ZN(P2_U3315) );
  INV_X1 U13432 ( .A(n10891), .ZN(n15252) );
  OAI222_X1 U13433 ( .A1(n14869), .A2(n10748), .B1(n14885), .B2(n10747), .C1(
        n15252), .C2(P1_U3086), .ZN(P1_U3343) );
  NAND2_X1 U13434 ( .A1(n10749), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n10751) );
  INV_X1 U13435 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n15531) );
  MUX2_X1 U13436 ( .A(n15531), .B(P2_REG1_REG_8__SCAN_IN), .S(n10784), .Z(
        n10750) );
  AOI21_X1 U13437 ( .B1(n10752), .B2(n10751), .A(n10750), .ZN(n10783) );
  NAND3_X1 U13438 ( .A1(n10752), .A2(n10751), .A3(n10750), .ZN(n10753) );
  NAND2_X1 U13439 ( .A1(n10753), .A2(n15456), .ZN(n10764) );
  INV_X1 U13440 ( .A(n15448), .ZN(n13722) );
  NAND2_X1 U13441 ( .A1(P2_U3088), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n11666) );
  OAI21_X1 U13442 ( .B1(n13722), .B2(n14907), .A(n11666), .ZN(n10754) );
  AOI21_X1 U13443 ( .B1(n10784), .B2(n15453), .A(n10754), .ZN(n10763) );
  NOR2_X1 U13444 ( .A1(n10756), .A2(n10755), .ZN(n10759) );
  MUX2_X1 U13445 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n10757), .S(n10784), .Z(
        n10758) );
  OAI21_X1 U13446 ( .B1(n10760), .B2(n10759), .A(n10758), .ZN(n10781) );
  OR3_X1 U13447 ( .A1(n10760), .A2(n10759), .A3(n10758), .ZN(n10761) );
  NAND3_X1 U13448 ( .A1(n15450), .A2(n10781), .A3(n10761), .ZN(n10762) );
  OAI211_X1 U13449 ( .C1(n10783), .C2(n10764), .A(n10763), .B(n10762), .ZN(
        P2_U3222) );
  INV_X1 U13450 ( .A(n10765), .ZN(n10768) );
  MUX2_X1 U13451 ( .A(n10516), .B(P2_REG1_REG_5__SCAN_IN), .S(n10766), .Z(
        n10767) );
  NAND2_X1 U13452 ( .A1(n10768), .A2(n10767), .ZN(n10770) );
  OAI211_X1 U13453 ( .C1(n15376), .C2(n10770), .A(n15456), .B(n10769), .ZN(
        n10771) );
  NAND2_X1 U13454 ( .A1(P2_U3088), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n11439) );
  OAI211_X1 U13455 ( .C1(n15756), .C2(n13722), .A(n10771), .B(n11439), .ZN(
        n10772) );
  INV_X1 U13456 ( .A(n10772), .ZN(n10779) );
  INV_X1 U13457 ( .A(n10773), .ZN(n10777) );
  NAND3_X1 U13458 ( .A1(n15380), .A2(n10775), .A3(n10774), .ZN(n10776) );
  NAND3_X1 U13459 ( .A1(n15450), .A2(n10777), .A3(n10776), .ZN(n10778) );
  OAI211_X1 U13460 ( .C1(n15401), .C2(n10780), .A(n10779), .B(n10778), .ZN(
        P2_U3219) );
  INV_X1 U13461 ( .A(n15450), .ZN(n15407) );
  NOR2_X1 U13462 ( .A1(n15407), .A2(n10788), .ZN(n10786) );
  OAI21_X1 U13463 ( .B1(n10757), .B2(n10782), .A(n10781), .ZN(n10789) );
  AOI21_X1 U13464 ( .B1(n10784), .B2(P2_REG1_REG_8__SCAN_IN), .A(n10783), .ZN(
        n10796) );
  INV_X1 U13465 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n15533) );
  NOR3_X1 U13466 ( .A1(n10796), .A2(n15533), .A3(n15375), .ZN(n10785) );
  AOI211_X1 U13467 ( .C1(n10786), .C2(n10789), .A(n15453), .B(n10785), .ZN(
        n10800) );
  AND2_X1 U13468 ( .A1(P2_U3088), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n10793) );
  MUX2_X1 U13469 ( .A(n10788), .B(P2_REG2_REG_9__SCAN_IN), .S(n10794), .Z(
        n10787) );
  NOR2_X1 U13470 ( .A1(n10789), .A2(n10787), .ZN(n11064) );
  INV_X1 U13471 ( .A(n11064), .ZN(n10791) );
  NAND3_X1 U13472 ( .A1(n10789), .A2(n11070), .A3(n10788), .ZN(n10790) );
  AOI21_X1 U13473 ( .B1(n10791), .B2(n10790), .A(n15407), .ZN(n10792) );
  AOI211_X1 U13474 ( .C1(n15448), .C2(P2_ADDR_REG_9__SCAN_IN), .A(n10793), .B(
        n10792), .ZN(n10799) );
  NOR3_X1 U13475 ( .A1(n10796), .A2(n10794), .A3(P2_REG1_REG_9__SCAN_IN), .ZN(
        n10797) );
  MUX2_X1 U13476 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n15533), .S(n10794), .Z(
        n10795) );
  OAI21_X1 U13477 ( .B1(n10797), .B2(n11069), .A(n15456), .ZN(n10798) );
  OAI211_X1 U13478 ( .C1(n10800), .C2(n11070), .A(n10799), .B(n10798), .ZN(
        P2_U3223) );
  AOI211_X1 U13479 ( .C1(n10803), .C2(n10802), .A(n15243), .B(n10801), .ZN(
        n10804) );
  INV_X1 U13480 ( .A(n10804), .ZN(n10811) );
  NAND2_X1 U13481 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3086), .ZN(n12416)
         );
  OAI211_X1 U13482 ( .C1(n10807), .C2(n10806), .A(n15258), .B(n10805), .ZN(
        n10808) );
  NAND2_X1 U13483 ( .A1(n12416), .A2(n10808), .ZN(n10809) );
  AOI21_X1 U13484 ( .B1(n14593), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n10809), 
        .ZN(n10810) );
  OAI211_X1 U13485 ( .C1(n15266), .C2(n10812), .A(n10811), .B(n10810), .ZN(
        P1_U3253) );
  NOR2_X1 U13486 ( .A1(n10814), .A2(n10813), .ZN(n10819) );
  XNOR2_X1 U13487 ( .A(n10817), .B(n12646), .ZN(n11017) );
  OAI22_X1 U13488 ( .A1(n11014), .A2(n11208), .B1(n10815), .B2(n12645), .ZN(
        n11016) );
  XNOR2_X1 U13489 ( .A(n11017), .B(n11016), .ZN(n10818) );
  AOI21_X1 U13490 ( .B1(n10819), .B2(n10818), .A(n11018), .ZN(n10822) );
  INV_X1 U13491 ( .A(n15111), .ZN(n15097) );
  AOI22_X1 U13492 ( .A1(n11189), .A2(n15097), .B1(n15107), .B2(n14502), .ZN(
        n10821) );
  NAND2_X1 U13493 ( .A1(n14195), .A2(n14762), .ZN(n15086) );
  INV_X1 U13494 ( .A(n15086), .ZN(n15109) );
  AOI22_X1 U13495 ( .A1(n15109), .A2(n6808), .B1(P1_REG3_REG_1__SCAN_IN), .B2(
        n11021), .ZN(n10820) );
  OAI211_X1 U13496 ( .C1(n10822), .C2(n15092), .A(n10821), .B(n10820), .ZN(
        P1_U3222) );
  OAI21_X1 U13497 ( .B1(n10825), .B2(n10824), .A(n10823), .ZN(n13927) );
  INV_X1 U13498 ( .A(n13927), .ZN(n10830) );
  XNOR2_X1 U13499 ( .A(n10825), .B(n9031), .ZN(n10827) );
  AOI22_X1 U13500 ( .A1(n13602), .A2(n13656), .B1(n13617), .B2(n9025), .ZN(
        n11458) );
  OAI21_X1 U13501 ( .B1(n10830), .B2(n11052), .A(n11458), .ZN(n10826) );
  AOI21_X1 U13502 ( .B1(n10827), .B2(n13906), .A(n10826), .ZN(n13934) );
  AOI21_X1 U13503 ( .B1(n11053), .B2(n13932), .A(n13912), .ZN(n10828) );
  AND2_X1 U13504 ( .A1(n10855), .A2(n10828), .ZN(n13929) );
  INV_X1 U13505 ( .A(n13929), .ZN(n10829) );
  OAI211_X1 U13506 ( .C1(n10830), .C2(n15511), .A(n13934), .B(n10829), .ZN(
        n11149) );
  OAI22_X1 U13507 ( .A1(n14016), .A2(n11459), .B1(n15539), .B2(n10510), .ZN(
        n10831) );
  AOI21_X1 U13508 ( .B1(n15539), .B2(n11149), .A(n10831), .ZN(n10832) );
  INV_X1 U13509 ( .A(n10832), .ZN(P2_U3500) );
  INV_X1 U13510 ( .A(n10833), .ZN(n10835) );
  OAI222_X1 U13511 ( .A1(n15016), .A2(P3_U3151), .B1(n12666), .B2(n10835), 
        .C1(n10834), .C2(n13440), .ZN(P3_U3278) );
  INV_X1 U13512 ( .A(n10836), .ZN(n10839) );
  INV_X1 U13513 ( .A(n13689), .ZN(n15400) );
  OAI222_X1 U13514 ( .A1(n14072), .A2(n10837), .B1(n14075), .B2(n10839), .C1(
        n15400), .C2(P2_U3088), .ZN(P2_U3314) );
  OAI222_X1 U13515 ( .A1(P1_U3086), .A2(n11255), .B1(n14885), .B2(n10839), 
        .C1(n10838), .C2(n14869), .ZN(P1_U3342) );
  NAND2_X1 U13516 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3086), .ZN(n11936) );
  OAI211_X1 U13517 ( .C1(n10842), .C2(n10841), .A(n15258), .B(n10840), .ZN(
        n10843) );
  NAND2_X1 U13518 ( .A1(n11936), .A2(n10843), .ZN(n10849) );
  INV_X1 U13519 ( .A(n10844), .ZN(n10845) );
  AOI211_X1 U13520 ( .C1(n10847), .C2(n10846), .A(n10845), .B(n15243), .ZN(
        n10848) );
  AOI211_X1 U13521 ( .C1(n14593), .C2(P1_ADDR_REG_6__SCAN_IN), .A(n10849), .B(
        n10848), .ZN(n10850) );
  OAI21_X1 U13522 ( .B1(n10851), .B2(n15266), .A(n10850), .ZN(P1_U3249) );
  NAND2_X1 U13523 ( .A1(n10854), .A2(n10853), .ZN(n11555) );
  NAND2_X1 U13524 ( .A1(n11129), .A2(n10855), .ZN(n10856) );
  NAND2_X1 U13525 ( .A1(n10856), .A2(n11777), .ZN(n10857) );
  NOR2_X1 U13526 ( .A1(n10872), .A2(n10857), .ZN(n11554) );
  XNOR2_X1 U13527 ( .A(n10859), .B(n10858), .ZN(n10861) );
  NAND2_X1 U13528 ( .A1(n13617), .A2(n13658), .ZN(n10860) );
  OAI21_X1 U13529 ( .B1(n13615), .B2(n11090), .A(n10860), .ZN(n11046) );
  AOI21_X1 U13530 ( .B1(n10861), .B2(n13906), .A(n11046), .ZN(n11558) );
  INV_X1 U13531 ( .A(n11558), .ZN(n10862) );
  AOI211_X1 U13532 ( .C1(n15491), .C2(n11555), .A(n11554), .B(n10862), .ZN(
        n11132) );
  INV_X1 U13533 ( .A(n14016), .ZN(n14002) );
  AOI22_X1 U13534 ( .A1(n14002), .A2(n11129), .B1(n15536), .B2(
        P2_REG1_REG_2__SCAN_IN), .ZN(n10863) );
  OAI21_X1 U13535 ( .B1(n11132), .B2(n15536), .A(n10863), .ZN(P2_U3501) );
  OR2_X1 U13536 ( .A1(n10865), .A2(n10864), .ZN(n10866) );
  NAND2_X1 U13537 ( .A1(n10867), .A2(n10866), .ZN(n11394) );
  INV_X1 U13538 ( .A(n11394), .ZN(n10873) );
  XNOR2_X1 U13539 ( .A(n10869), .B(n10868), .ZN(n10871) );
  OAI22_X1 U13540 ( .A1(n13577), .A2(n7492), .B1(n10870), .B2(n13615), .ZN(
        n13514) );
  AOI21_X1 U13541 ( .B1(n10871), .B2(n13906), .A(n13514), .ZN(n11395) );
  OAI211_X1 U13542 ( .C1(n10872), .C2(n11144), .A(n11777), .B(n11085), .ZN(
        n11388) );
  OAI211_X1 U13543 ( .C1(n10873), .C2(n14022), .A(n11395), .B(n11388), .ZN(
        n11146) );
  INV_X1 U13544 ( .A(n11146), .ZN(n10875) );
  AOI22_X1 U13545 ( .A1(n14002), .A2(n13515), .B1(n15536), .B2(
        P2_REG1_REG_3__SCAN_IN), .ZN(n10874) );
  OAI21_X1 U13546 ( .B1(n10875), .B2(n15536), .A(n10874), .ZN(P2_U3502) );
  NOR2_X1 U13547 ( .A1(n12790), .A2(P3_U3151), .ZN(n11174) );
  AND2_X1 U13548 ( .A1(n15699), .A2(n11368), .ZN(n12846) );
  INV_X1 U13549 ( .A(n12846), .ZN(n12849) );
  NAND2_X1 U13550 ( .A1(n11025), .A2(n12849), .ZN(n12823) );
  INV_X1 U13551 ( .A(n12794), .ZN(n12774) );
  INV_X1 U13552 ( .A(n15682), .ZN(n10901) );
  OAI22_X1 U13553 ( .A1(n12774), .A2(n10901), .B1(n11368), .B2(n12797), .ZN(
        n10876) );
  AOI21_X1 U13554 ( .B1(n12788), .B2(n12823), .A(n10876), .ZN(n10877) );
  OAI21_X1 U13555 ( .B1(n11174), .B2(n11364), .A(n10877), .ZN(P3_U3172) );
  INV_X1 U13556 ( .A(n15023), .ZN(n13046) );
  OAI222_X1 U13557 ( .A1(P3_U3151), .A2(n13046), .B1(n13440), .B2(n10879), 
        .C1(n12666), .C2(n10878), .ZN(P3_U3277) );
  NOR2_X1 U13558 ( .A1(n15266), .A2(n11255), .ZN(n10888) );
  NAND2_X1 U13559 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n15116)
         );
  NOR2_X1 U13560 ( .A1(n10891), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n10882) );
  INV_X1 U13561 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n10880) );
  AOI22_X1 U13562 ( .A1(n10891), .A2(n10880), .B1(P1_REG2_REG_12__SCAN_IN), 
        .B2(n15252), .ZN(n15247) );
  OAI21_X1 U13563 ( .B1(n10890), .B2(n10610), .A(n10881), .ZN(n15246) );
  NOR2_X1 U13564 ( .A1(n15247), .A2(n15246), .ZN(n15245) );
  NOR2_X1 U13565 ( .A1(n10882), .A2(n15245), .ZN(n10885) );
  INV_X1 U13566 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n10883) );
  MUX2_X1 U13567 ( .A(n10883), .B(P1_REG2_REG_13__SCAN_IN), .S(n11255), .Z(
        n10884) );
  NAND2_X1 U13568 ( .A1(n10884), .A2(n10885), .ZN(n11254) );
  OAI211_X1 U13569 ( .C1(n10885), .C2(n10884), .A(n11254), .B(n15258), .ZN(
        n10886) );
  NAND2_X1 U13570 ( .A1(n15116), .A2(n10886), .ZN(n10887) );
  AOI211_X1 U13571 ( .C1(n14593), .C2(P1_ADDR_REG_13__SCAN_IN), .A(n10888), 
        .B(n10887), .ZN(n10897) );
  AOI21_X1 U13572 ( .B1(n15185), .B2(n10890), .A(n10889), .ZN(n15242) );
  INV_X1 U13573 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n14944) );
  AOI22_X1 U13574 ( .A1(n10891), .A2(n14944), .B1(P1_REG1_REG_12__SCAN_IN), 
        .B2(n15252), .ZN(n15241) );
  NOR2_X1 U13575 ( .A1(n15242), .A2(n15241), .ZN(n15240) );
  NOR2_X1 U13576 ( .A1(n10891), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n10892) );
  NOR2_X1 U13577 ( .A1(n15240), .A2(n10892), .ZN(n10895) );
  INV_X1 U13578 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n10893) );
  MUX2_X1 U13579 ( .A(n10893), .B(P1_REG1_REG_13__SCAN_IN), .S(n11255), .Z(
        n10894) );
  NAND2_X1 U13580 ( .A1(n10895), .A2(n10894), .ZN(n11247) );
  OAI211_X1 U13581 ( .C1(n10895), .C2(n10894), .A(n15261), .B(n11247), .ZN(
        n10896) );
  NAND2_X1 U13582 ( .A1(n10897), .A2(n10896), .ZN(P1_U3256) );
  INV_X1 U13583 ( .A(n10898), .ZN(n10899) );
  OAI21_X1 U13584 ( .B1(n10899), .B2(n15703), .A(n12823), .ZN(n10900) );
  OAI21_X1 U13585 ( .B1(n10901), .B2(n13278), .A(n10900), .ZN(n11366) );
  AOI21_X1 U13586 ( .B1(n15070), .B2(n10902), .A(n11366), .ZN(n11035) );
  NAND2_X1 U13587 ( .A1(n15743), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n10903) );
  OAI21_X1 U13588 ( .B1(n11035), .B2(n15743), .A(n10903), .ZN(P3_U3390) );
  MUX2_X1 U13589 ( .A(P3_REG2_REG_3__SCAN_IN), .B(P3_REG1_REG_3__SCAN_IN), .S(
        n13027), .Z(n10932) );
  XOR2_X1 U13590 ( .A(n10929), .B(n10932), .Z(n10933) );
  MUX2_X1 U13591 ( .A(P3_REG2_REG_1__SCAN_IN), .B(P3_REG1_REG_1__SCAN_IN), .S(
        n13029), .Z(n10904) );
  XNOR2_X1 U13592 ( .A(n10904), .B(n11313), .ZN(n11296) );
  MUX2_X1 U13593 ( .A(n10911), .B(n8452), .S(n13029), .Z(n15543) );
  NAND2_X1 U13594 ( .A1(n15543), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n15542) );
  OAI22_X1 U13595 ( .A1(n11296), .A2(n15542), .B1(n10904), .B2(n11313), .ZN(
        n10952) );
  MUX2_X1 U13596 ( .A(P3_REG2_REG_2__SCAN_IN), .B(P3_REG1_REG_2__SCAN_IN), .S(
        n13029), .Z(n10905) );
  XNOR2_X1 U13597 ( .A(n10905), .B(n10967), .ZN(n10953) );
  INV_X1 U13598 ( .A(n10905), .ZN(n10906) );
  AOI22_X1 U13599 ( .A1(n10952), .A2(n10953), .B1(n10967), .B2(n10906), .ZN(
        n10934) );
  XOR2_X1 U13600 ( .A(n10934), .B(n10933), .Z(n10931) );
  NAND2_X1 U13601 ( .A1(P3_U3897), .A2(n12667), .ZN(n15611) );
  OR2_X1 U13602 ( .A1(n10910), .A2(P3_U3151), .ZN(n12992) );
  INV_X1 U13603 ( .A(n12992), .ZN(n10908) );
  OR2_X1 U13604 ( .A1(n10908), .A2(n10907), .ZN(n10920) );
  AOI21_X1 U13605 ( .B1(n12963), .B2(n10910), .A(n10909), .ZN(n10918) );
  MUX2_X1 U13606 ( .A(n10921), .B(P3_U3897), .S(n12987), .Z(n15540) );
  XNOR2_X1 U13607 ( .A(n10967), .B(P3_REG2_REG_2__SCAN_IN), .ZN(n10961) );
  NOR2_X1 U13608 ( .A1(n10911), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n10912) );
  NAND2_X1 U13609 ( .A1(n7289), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n10913) );
  NAND2_X1 U13610 ( .A1(n10961), .A2(n10960), .ZN(n10959) );
  AOI21_X1 U13611 ( .B1(n12018), .B2(n10915), .A(n10935), .ZN(n10927) );
  INV_X1 U13612 ( .A(n10916), .ZN(n10917) );
  INV_X1 U13613 ( .A(n10918), .ZN(n10919) );
  NOR2_X1 U13614 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12020), .ZN(n11241) );
  NAND2_X1 U13615 ( .A1(n10921), .A2(n13027), .ZN(n15541) );
  INV_X1 U13616 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n10923) );
  MUX2_X1 U13617 ( .A(n10923), .B(P3_REG1_REG_2__SCAN_IN), .S(n10967), .Z(
        n10956) );
  AND2_X1 U13618 ( .A1(P3_REG1_REG_0__SCAN_IN), .A2(n7030), .ZN(n10922) );
  OAI21_X1 U13619 ( .B1(n11313), .B2(n10922), .A(n6699), .ZN(n11298) );
  INV_X1 U13620 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n11297) );
  OR2_X1 U13621 ( .A1(n11298), .A2(n11297), .ZN(n11300) );
  NAND2_X1 U13622 ( .A1(n11300), .A2(n6699), .ZN(n10955) );
  NAND2_X1 U13623 ( .A1(n10956), .A2(n10955), .ZN(n10954) );
  OAI21_X1 U13624 ( .B1(n10967), .B2(n10923), .A(n10954), .ZN(n10941) );
  XNOR2_X1 U13625 ( .A(n10941), .B(n10929), .ZN(n10942) );
  XOR2_X1 U13626 ( .A(P3_REG1_REG_3__SCAN_IN), .B(n10942), .Z(n10924) );
  NOR2_X1 U13627 ( .A1(n15541), .A2(n10924), .ZN(n10925) );
  AOI211_X1 U13628 ( .C1(n15623), .C2(P3_ADDR_REG_3__SCAN_IN), .A(n11241), .B(
        n10925), .ZN(n10926) );
  OAI21_X1 U13629 ( .B1(n10927), .B2(n15636), .A(n10926), .ZN(n10928) );
  AOI21_X1 U13630 ( .B1(n10929), .B2(n15540), .A(n10928), .ZN(n10930) );
  OAI21_X1 U13631 ( .B1(n10931), .B2(n15611), .A(n10930), .ZN(P3_U3185) );
  MUX2_X1 U13632 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n13027), .Z(n10970) );
  XNOR2_X1 U13633 ( .A(n10970), .B(n10982), .ZN(n10972) );
  OAI22_X1 U13634 ( .A1(n10934), .A2(n10933), .B1(n10932), .B2(n7299), .ZN(
        n10973) );
  XOR2_X1 U13635 ( .A(n10973), .B(n10972), .Z(n10951) );
  NAND2_X1 U13636 ( .A1(n10937), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n10974) );
  OAI21_X1 U13637 ( .B1(n10937), .B2(P3_REG2_REG_4__SCAN_IN), .A(n10974), .ZN(
        n10938) );
  AOI21_X1 U13638 ( .B1(n10939), .B2(n10938), .A(n10976), .ZN(n10948) );
  NOR2_X1 U13639 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10940), .ZN(n11538) );
  MUX2_X1 U13640 ( .A(P3_REG1_REG_4__SCAN_IN), .B(n10981), .S(n10982), .Z(
        n10944) );
  AOI22_X1 U13641 ( .A1(n10942), .A2(P3_REG1_REG_3__SCAN_IN), .B1(n7299), .B2(
        n10941), .ZN(n10943) );
  NOR2_X1 U13642 ( .A1(n10943), .A2(n10944), .ZN(n10979) );
  AOI21_X1 U13643 ( .B1(n10944), .B2(n10943), .A(n10979), .ZN(n10945) );
  NOR2_X1 U13644 ( .A1(n15541), .A2(n10945), .ZN(n10946) );
  AOI211_X1 U13645 ( .C1(n15623), .C2(P3_ADDR_REG_4__SCAN_IN), .A(n11538), .B(
        n10946), .ZN(n10947) );
  OAI21_X1 U13646 ( .B1(n10948), .B2(n15636), .A(n10947), .ZN(n10949) );
  AOI21_X1 U13647 ( .B1(n10982), .B2(n15540), .A(n10949), .ZN(n10950) );
  OAI21_X1 U13648 ( .B1(n10951), .B2(n15611), .A(n10950), .ZN(P3_U3186) );
  XOR2_X1 U13649 ( .A(n10952), .B(n10953), .Z(n10969) );
  OAI21_X1 U13650 ( .B1(n10956), .B2(n10955), .A(n10954), .ZN(n10957) );
  NAND2_X1 U13651 ( .A1(n15628), .A2(n10957), .ZN(n10965) );
  NOR2_X1 U13652 ( .A1(n11173), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10958) );
  AOI21_X1 U13653 ( .B1(n15623), .B2(P3_ADDR_REG_2__SCAN_IN), .A(n10958), .ZN(
        n10964) );
  OAI21_X1 U13654 ( .B1(n10961), .B2(n10960), .A(n10959), .ZN(n10962) );
  NAND2_X1 U13655 ( .A1(n15032), .A2(n10962), .ZN(n10963) );
  NAND3_X1 U13656 ( .A1(n10965), .A2(n10964), .A3(n10963), .ZN(n10966) );
  AOI21_X1 U13657 ( .B1(n10967), .B2(n15540), .A(n10966), .ZN(n10968) );
  OAI21_X1 U13658 ( .B1(n10969), .B2(n15611), .A(n10968), .ZN(P3_U3184) );
  MUX2_X1 U13659 ( .A(P3_REG2_REG_5__SCAN_IN), .B(P3_REG1_REG_5__SCAN_IN), .S(
        n13027), .Z(n10991) );
  XNOR2_X1 U13660 ( .A(n10991), .B(n10995), .ZN(n10992) );
  INV_X1 U13661 ( .A(n10970), .ZN(n10971) );
  AOI22_X1 U13662 ( .A1(n10973), .A2(n10972), .B1(n10982), .B2(n10971), .ZN(
        n10993) );
  XOR2_X1 U13663 ( .A(n10992), .B(n10993), .Z(n10990) );
  INV_X1 U13664 ( .A(n10974), .ZN(n10975) );
  AOI21_X1 U13665 ( .B1(n10978), .B2(n8523), .A(n11001), .ZN(n10987) );
  NOR2_X1 U13666 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n8527), .ZN(n11653) );
  AOI21_X1 U13667 ( .B1(n15623), .B2(P3_ADDR_REG_5__SCAN_IN), .A(n11653), .ZN(
        n10986) );
  INV_X1 U13668 ( .A(n10979), .ZN(n10980) );
  OAI21_X1 U13669 ( .B1(P3_REG1_REG_5__SCAN_IN), .B2(n10983), .A(n10996), .ZN(
        n10984) );
  NAND2_X1 U13670 ( .A1(n15628), .A2(n10984), .ZN(n10985) );
  OAI211_X1 U13671 ( .C1(n15636), .C2(n10987), .A(n10986), .B(n10985), .ZN(
        n10988) );
  AOI21_X1 U13672 ( .B1(n7022), .B2(n15540), .A(n10988), .ZN(n10989) );
  OAI21_X1 U13673 ( .B1(n10990), .B2(n15611), .A(n10989), .ZN(P3_U3187) );
  MUX2_X1 U13674 ( .A(P3_REG2_REG_6__SCAN_IN), .B(P3_REG1_REG_6__SCAN_IN), .S(
        n13027), .Z(n11151) );
  XNOR2_X1 U13675 ( .A(n11151), .B(n11153), .ZN(n11154) );
  OAI22_X1 U13676 ( .A1(n10993), .A2(n10992), .B1(n10991), .B2(n10995), .ZN(
        n11155) );
  XOR2_X1 U13677 ( .A(n11154), .B(n11155), .Z(n11010) );
  AOI22_X1 U13678 ( .A1(n11153), .A2(n8544), .B1(P3_REG1_REG_6__SCAN_IN), .B2(
        n11163), .ZN(n10999) );
  NAND2_X1 U13679 ( .A1(n10995), .A2(n10994), .ZN(n10997) );
  NAND2_X1 U13680 ( .A1(n10999), .A2(n10998), .ZN(n11156) );
  OAI21_X1 U13681 ( .B1(n10999), .B2(n10998), .A(n11156), .ZN(n11000) );
  INV_X1 U13682 ( .A(n11000), .ZN(n11007) );
  NAND2_X1 U13683 ( .A1(P3_REG2_REG_6__SCAN_IN), .A2(n11163), .ZN(n11002) );
  OAI21_X1 U13684 ( .B1(P3_REG2_REG_6__SCAN_IN), .B2(n11163), .A(n11002), .ZN(
        n11161) );
  XNOR2_X1 U13685 ( .A(n11162), .B(n11161), .ZN(n11003) );
  NAND2_X1 U13686 ( .A1(n15032), .A2(n11003), .ZN(n11006) );
  INV_X1 U13687 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n11004) );
  NOR2_X1 U13688 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11004), .ZN(n11700) );
  AOI21_X1 U13689 ( .B1(n15623), .B2(P3_ADDR_REG_6__SCAN_IN), .A(n11700), .ZN(
        n11005) );
  OAI211_X1 U13690 ( .C1(n15541), .C2(n11007), .A(n11006), .B(n11005), .ZN(
        n11008) );
  AOI21_X1 U13691 ( .B1(n11153), .B2(n15540), .A(n11008), .ZN(n11009) );
  OAI21_X1 U13692 ( .B1(n11010), .B2(n15611), .A(n11009), .ZN(P3_U3188) );
  NAND2_X1 U13693 ( .A1(n12771), .A2(P3_U3897), .ZN(n11011) );
  OAI21_X1 U13694 ( .B1(P3_U3897), .B2(n11012), .A(n11011), .ZN(P3_U3512) );
  OAI22_X1 U13695 ( .A1(n15281), .A2(n12648), .B1(n11203), .B2(n12645), .ZN(
        n11013) );
  XNOR2_X1 U13696 ( .A(n11013), .B(n12646), .ZN(n11195) );
  NAND2_X1 U13697 ( .A1(n14224), .A2(n11192), .ZN(n11015) );
  OAI21_X1 U13698 ( .B1(n12644), .B2(n11203), .A(n11015), .ZN(n11194) );
  XNOR2_X1 U13699 ( .A(n11195), .B(n11194), .ZN(n11196) );
  INV_X1 U13700 ( .A(n11016), .ZN(n11020) );
  INV_X1 U13701 ( .A(n11017), .ZN(n11019) );
  XOR2_X1 U13702 ( .A(n11196), .B(n11197), .Z(n11024) );
  AOI22_X1 U13703 ( .A1(n15109), .A2(n6847), .B1(n15097), .B2(n14224), .ZN(
        n11023) );
  AOI22_X1 U13704 ( .A1(n15107), .A2(n14500), .B1(n11021), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n11022) );
  OAI211_X1 U13705 ( .C1(n11024), .C2(n15092), .A(n11023), .B(n11022), .ZN(
        P1_U3237) );
  NAND3_X1 U13706 ( .A1(n15702), .A2(n11025), .A3(n12669), .ZN(n11026) );
  OAI211_X1 U13707 ( .C1(n11028), .C2(n15701), .A(n11027), .B(n11026), .ZN(
        n11029) );
  NAND2_X1 U13708 ( .A1(n11029), .A2(n12788), .ZN(n11033) );
  INV_X1 U13709 ( .A(n12792), .ZN(n12770) );
  INV_X1 U13710 ( .A(n15698), .ZN(n11030) );
  OAI22_X1 U13711 ( .A1(n12774), .A2(n11030), .B1(n15695), .B2(n12797), .ZN(
        n11031) );
  AOI21_X1 U13712 ( .B1(n12770), .B2(n15699), .A(n11031), .ZN(n11032) );
  OAI211_X1 U13713 ( .C1(n11174), .C2(n11305), .A(n11033), .B(n11032), .ZN(
        P3_U3162) );
  NAND2_X1 U13714 ( .A1(n15749), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n11034) );
  OAI21_X1 U13715 ( .B1(n11035), .B2(n15749), .A(n11034), .ZN(P3_U3459) );
  INV_X1 U13716 ( .A(n11036), .ZN(n11039) );
  OR2_X1 U13717 ( .A1(n15469), .A2(n11037), .ZN(n11042) );
  OAI21_X1 U13718 ( .B1(n11039), .B2(n11042), .A(n11038), .ZN(n11041) );
  NAND2_X1 U13719 ( .A1(n11041), .A2(n11040), .ZN(n11279) );
  INV_X1 U13720 ( .A(n15470), .ZN(n15467) );
  NOR2_X1 U13721 ( .A1(n11279), .A2(n15467), .ZN(n11121) );
  INV_X1 U13722 ( .A(n11042), .ZN(n11383) );
  NAND2_X1 U13723 ( .A1(n11043), .A2(n11383), .ZN(n11047) );
  NAND2_X1 U13724 ( .A1(n11490), .A2(n8333), .ZN(n11389) );
  OAI21_X2 U13725 ( .B1(n11047), .B2(n11389), .A(n13916), .ZN(n13624) );
  AOI22_X1 U13726 ( .A1(n11129), .A2(n13624), .B1(n13605), .B2(n11046), .ZN(
        n11063) );
  INV_X1 U13727 ( .A(n11047), .ZN(n11050) );
  AND2_X1 U13728 ( .A1(n11048), .A2(n15516), .ZN(n11049) );
  XNOR2_X1 U13729 ( .A(n13537), .B(n13932), .ZN(n11056) );
  NAND2_X1 U13730 ( .A1(n13658), .A2(n8410), .ZN(n11057) );
  XNOR2_X1 U13731 ( .A(n11056), .B(n11057), .ZN(n11457) );
  AND2_X1 U13732 ( .A1(n13537), .A2(n11491), .ZN(n11055) );
  NAND2_X1 U13733 ( .A1(n11053), .A2(n11777), .ZN(n11054) );
  NAND2_X1 U13734 ( .A1(n9031), .A2(n11054), .ZN(n11123) );
  NAND2_X1 U13735 ( .A1(n11457), .A2(n11456), .ZN(n11060) );
  INV_X1 U13736 ( .A(n11056), .ZN(n11058) );
  NAND2_X1 U13737 ( .A1(n11058), .A2(n11057), .ZN(n11059) );
  NAND2_X1 U13738 ( .A1(n11060), .A2(n11059), .ZN(n11262) );
  XNOR2_X1 U13739 ( .A(n11129), .B(n13537), .ZN(n11265) );
  NAND2_X1 U13740 ( .A1(n13656), .A2(n8410), .ZN(n11263) );
  XNOR2_X1 U13741 ( .A(n11265), .B(n11263), .ZN(n11261) );
  XNOR2_X1 U13742 ( .A(n11262), .B(n11261), .ZN(n11061) );
  NAND2_X1 U13743 ( .A1(n13591), .A2(n11061), .ZN(n11062) );
  OAI211_X1 U13744 ( .C1(n11121), .C2(n11550), .A(n11063), .B(n11062), .ZN(
        P2_U3209) );
  MUX2_X1 U13745 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n11065), .S(n11072), .Z(
        n15394) );
  NAND2_X1 U13746 ( .A1(n15395), .A2(n15394), .ZN(n15393) );
  OAI21_X1 U13747 ( .B1(n11065), .B2(n15387), .A(n15393), .ZN(n11068) );
  MUX2_X1 U13748 ( .A(n11066), .B(P2_REG2_REG_11__SCAN_IN), .S(n11229), .Z(
        n11067) );
  AOI21_X1 U13749 ( .B1(n11068), .B2(n11067), .A(n11232), .ZN(n11081) );
  AOI21_X1 U13750 ( .B1(n15533), .B2(n11070), .A(n11069), .ZN(n15392) );
  INV_X1 U13751 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n11071) );
  MUX2_X1 U13752 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n11071), .S(n11072), .Z(
        n15391) );
  NAND2_X1 U13753 ( .A1(n15392), .A2(n15391), .ZN(n15390) );
  NAND2_X1 U13754 ( .A1(n11072), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n11074) );
  INV_X1 U13755 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n15537) );
  MUX2_X1 U13756 ( .A(n15537), .B(P2_REG1_REG_11__SCAN_IN), .S(n11229), .Z(
        n11073) );
  AOI21_X1 U13757 ( .B1(n15390), .B2(n11074), .A(n11073), .ZN(n11225) );
  INV_X1 U13758 ( .A(n11225), .ZN(n11076) );
  NAND3_X1 U13759 ( .A1(n15390), .A2(n11074), .A3(n11073), .ZN(n11075) );
  NAND3_X1 U13760 ( .A1(n11076), .A2(n15456), .A3(n11075), .ZN(n11080) );
  INV_X1 U13761 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n11077) );
  NAND2_X1 U13762 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_U3088), .ZN(n12071)
         );
  OAI21_X1 U13763 ( .B1(n13722), .B2(n11077), .A(n12071), .ZN(n11078) );
  AOI21_X1 U13764 ( .B1(n11229), .B2(n15453), .A(n11078), .ZN(n11079) );
  OAI211_X1 U13765 ( .C1(n11081), .C2(n15407), .A(n11080), .B(n11079), .ZN(
        P2_U3225) );
  OAI21_X1 U13766 ( .B1(n11084), .B2(n11083), .A(n11082), .ZN(n11405) );
  AOI21_X1 U13767 ( .B1(n11085), .B2(n11400), .A(n13912), .ZN(n11086) );
  NAND2_X1 U13768 ( .A1(n11086), .A2(n11518), .ZN(n11399) );
  INV_X1 U13769 ( .A(n11399), .ZN(n11093) );
  XNOR2_X1 U13770 ( .A(n11088), .B(n11087), .ZN(n11091) );
  OAI22_X1 U13771 ( .A1(n13577), .A2(n11090), .B1(n11089), .B2(n13615), .ZN(
        n11281) );
  AOI21_X1 U13772 ( .B1(n11091), .B2(n13906), .A(n11281), .ZN(n11406) );
  INV_X1 U13773 ( .A(n11406), .ZN(n11092) );
  AOI211_X1 U13774 ( .C1(n15491), .C2(n11405), .A(n11093), .B(n11092), .ZN(
        n11135) );
  AOI22_X1 U13775 ( .A1(n14002), .A2(n11400), .B1(n15536), .B2(
        P2_REG1_REG_4__SCAN_IN), .ZN(n11094) );
  OAI21_X1 U13776 ( .B1(n11135), .B2(n15536), .A(n11094), .ZN(P2_U3503) );
  OR2_X1 U13777 ( .A1(n11099), .A2(n11103), .ZN(n11100) );
  NAND2_X1 U13778 ( .A1(n11101), .A2(n11100), .ZN(n11107) );
  INV_X1 U13779 ( .A(n11107), .ZN(n11143) );
  NAND3_X1 U13780 ( .A1(n11206), .A2(n11103), .A3(n11102), .ZN(n11104) );
  NAND2_X1 U13781 ( .A1(n11105), .A2(n11104), .ZN(n11106) );
  NAND2_X1 U13782 ( .A1(n11106), .A2(n15160), .ZN(n11110) );
  INV_X1 U13783 ( .A(n14928), .ZN(n15317) );
  NAND2_X1 U13784 ( .A1(n11107), .A2(n15317), .ZN(n11109) );
  AOI22_X1 U13785 ( .A1(n15134), .A2(n14499), .B1(n14762), .B2(n14502), .ZN(
        n11108) );
  AND3_X1 U13786 ( .A1(n11110), .A2(n11109), .A3(n11108), .ZN(n11139) );
  INV_X1 U13787 ( .A(n11217), .ZN(n11112) );
  INV_X1 U13788 ( .A(n11341), .ZN(n11111) );
  OAI211_X1 U13789 ( .C1(n6672), .C2(n11112), .A(n11111), .B(n15122), .ZN(
        n11137) );
  INV_X1 U13790 ( .A(n11137), .ZN(n11113) );
  AOI21_X1 U13791 ( .B1(n15310), .B2(n14228), .A(n11113), .ZN(n11114) );
  OAI211_X1 U13792 ( .C1(n11143), .C2(n15313), .A(n11139), .B(n11114), .ZN(
        n11116) );
  NAND2_X1 U13793 ( .A1(n11116), .A2(n15358), .ZN(n11115) );
  OAI21_X1 U13794 ( .B1(n15358), .B2(n10554), .A(n11115), .ZN(P1_U3531) );
  INV_X1 U13795 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n11118) );
  NAND2_X1 U13796 ( .A1(n11116), .A2(n15341), .ZN(n11117) );
  OAI21_X1 U13797 ( .B1(n15341), .B2(n11118), .A(n11117), .ZN(P1_U3468) );
  OAI222_X1 U13798 ( .A1(n12666), .A2(n11120), .B1(n13440), .B2(n11119), .C1(
        P3_U3151), .C2(n13037), .ZN(P3_U3276) );
  INV_X1 U13799 ( .A(n11121), .ZN(n11461) );
  NAND2_X1 U13800 ( .A1(n11461), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n11128) );
  NOR2_X1 U13801 ( .A1(n13615), .A2(n11122), .ZN(n11494) );
  INV_X1 U13802 ( .A(n11123), .ZN(n11124) );
  OAI21_X1 U13803 ( .B1(n11777), .B2(n11125), .A(n11124), .ZN(n11126) );
  AOI22_X1 U13804 ( .A1(n13605), .A2(n11494), .B1(n13591), .B2(n11126), .ZN(
        n11127) );
  OAI211_X1 U13805 ( .C1(n13597), .C2(n11491), .A(n11128), .B(n11127), .ZN(
        P2_U3204) );
  INV_X1 U13806 ( .A(n11129), .ZN(n11551) );
  OAI22_X1 U13807 ( .A1(n14062), .A2(n11551), .B1(n15524), .B2(n7732), .ZN(
        n11130) );
  INV_X1 U13808 ( .A(n11130), .ZN(n11131) );
  OAI21_X1 U13809 ( .B1(n11132), .B2(n15523), .A(n11131), .ZN(P2_U3436) );
  NOR2_X1 U13810 ( .A1(n15524), .A2(n7795), .ZN(n11133) );
  AOI21_X1 U13811 ( .B1(n8423), .B2(n11400), .A(n11133), .ZN(n11134) );
  OAI21_X1 U13812 ( .B1(n11135), .B2(n15523), .A(n11134), .ZN(P2_U3442) );
  NAND2_X1 U13813 ( .A1(n14218), .A2(n14209), .ZN(n14414) );
  INV_X1 U13814 ( .A(n14414), .ZN(n11136) );
  NAND2_X1 U13815 ( .A1(n15143), .A2(n11136), .ZN(n14921) );
  OAI22_X1 U13816 ( .A1(n14958), .A2(n11137), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(n15136), .ZN(n11138) );
  AOI21_X1 U13817 ( .B1(n14717), .B2(n14228), .A(n11138), .ZN(n11142) );
  MUX2_X1 U13818 ( .A(n11140), .B(n11139), .S(n15143), .Z(n11141) );
  OAI211_X1 U13819 ( .C1(n11143), .C2(n14921), .A(n11142), .B(n11141), .ZN(
        P1_U3290) );
  OAI22_X1 U13820 ( .A1(n14062), .A2(n11144), .B1(n15524), .B2(n7776), .ZN(
        n11145) );
  AOI21_X1 U13821 ( .B1(n15524), .B2(n11146), .A(n11145), .ZN(n11147) );
  INV_X1 U13822 ( .A(n11147), .ZN(P2_U3439) );
  OAI22_X1 U13823 ( .A1(n14062), .A2(n11459), .B1(n15524), .B2(n7747), .ZN(
        n11148) );
  AOI21_X1 U13824 ( .B1(n15524), .B2(n11149), .A(n11148), .ZN(n11150) );
  INV_X1 U13825 ( .A(n11150), .ZN(P2_U3433) );
  MUX2_X1 U13826 ( .A(P3_REG2_REG_7__SCAN_IN), .B(P3_REG1_REG_7__SCAN_IN), .S(
        n13027), .Z(n11314) );
  XNOR2_X1 U13827 ( .A(n11314), .B(n11327), .ZN(n11315) );
  INV_X1 U13828 ( .A(n11151), .ZN(n11152) );
  XOR2_X1 U13829 ( .A(n11315), .B(n11316), .Z(n11170) );
  NAND2_X1 U13830 ( .A1(P3_REG1_REG_6__SCAN_IN), .A2(n11163), .ZN(n11157) );
  NAND2_X1 U13831 ( .A1(n11157), .A2(n11156), .ZN(n11326) );
  XOR2_X1 U13832 ( .A(n11326), .B(n11327), .Z(n11158) );
  NAND2_X1 U13833 ( .A1(P3_REG1_REG_7__SCAN_IN), .A2(n11158), .ZN(n11328) );
  OAI21_X1 U13834 ( .B1(P3_REG1_REG_7__SCAN_IN), .B2(n11158), .A(n11328), .ZN(
        n11168) );
  NOR2_X1 U13835 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11159), .ZN(n11822) );
  AOI21_X1 U13836 ( .B1(n15623), .B2(P3_ADDR_REG_7__SCAN_IN), .A(n11822), .ZN(
        n11160) );
  OAI21_X1 U13837 ( .B1(n15626), .B2(n11327), .A(n11160), .ZN(n11167) );
  AOI21_X1 U13838 ( .B1(n11164), .B2(n8563), .A(n11323), .ZN(n11165) );
  NOR2_X1 U13839 ( .A1(n11165), .A2(n15636), .ZN(n11166) );
  AOI211_X1 U13840 ( .C1(n15628), .C2(n11168), .A(n11167), .B(n11166), .ZN(
        n11169) );
  OAI21_X1 U13841 ( .B1(n11170), .B2(n15611), .A(n11169), .ZN(P3_U3189) );
  XOR2_X1 U13842 ( .A(n11172), .B(n11171), .Z(n11178) );
  OAI22_X1 U13843 ( .A1(n12774), .A2(n7124), .B1(n12797), .B2(n15687), .ZN(
        n11176) );
  NOR2_X1 U13844 ( .A1(n11174), .A2(n11173), .ZN(n11175) );
  AOI211_X1 U13845 ( .C1(n12770), .C2(n15682), .A(n11176), .B(n11175), .ZN(
        n11177) );
  OAI21_X1 U13846 ( .B1(n11178), .B2(n12777), .A(n11177), .ZN(P3_U3177) );
  OAI21_X1 U13847 ( .B1(n14418), .B2(n11180), .A(n11179), .ZN(n15278) );
  OAI22_X1 U13848 ( .A1(n11203), .A2(n14947), .B1(n11181), .B2(n15131), .ZN(
        n11186) );
  OAI21_X1 U13849 ( .B1(n10815), .B2(n11294), .A(n11216), .ZN(n11187) );
  XNOR2_X1 U13850 ( .A(n11187), .B(n11208), .ZN(n11183) );
  INV_X1 U13851 ( .A(n14418), .ZN(n11182) );
  MUX2_X1 U13852 ( .A(n11183), .B(n11182), .S(n6808), .Z(n11184) );
  NOR2_X1 U13853 ( .A1(n11184), .A2(n15175), .ZN(n11185) );
  AOI211_X1 U13854 ( .C1(n15317), .C2(n15278), .A(n11186), .B(n11185), .ZN(
        n15275) );
  NOR2_X1 U13855 ( .A1(n11187), .A2(n14741), .ZN(n15273) );
  INV_X1 U13856 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n14506) );
  OAI22_X1 U13857 ( .A1(n15143), .A2(n10571), .B1(n14506), .B2(n15136), .ZN(
        n11188) );
  AOI21_X1 U13858 ( .B1(n15125), .B2(n15273), .A(n11188), .ZN(n11191) );
  INV_X1 U13859 ( .A(n14921), .ZN(n11220) );
  AOI22_X1 U13860 ( .A1(n11220), .A2(n15278), .B1(n14717), .B2(n11189), .ZN(
        n11190) );
  OAI211_X1 U13861 ( .C1(n15275), .C2(n14765), .A(n11191), .B(n11190), .ZN(
        P1_U3292) );
  INV_X4 U13862 ( .A(n11192), .ZN(n12645) );
  AOI22_X1 U13863 ( .A1(n14228), .A2(n12635), .B1(n12621), .B2(n14500), .ZN(
        n11193) );
  XNOR2_X1 U13864 ( .A(n11193), .B(n12646), .ZN(n11708) );
  AOI22_X1 U13865 ( .A1(n10728), .A2(n14500), .B1(n12621), .B2(n14228), .ZN(
        n11707) );
  XNOR2_X1 U13866 ( .A(n11708), .B(n11707), .ZN(n11199) );
  AOI211_X1 U13867 ( .C1(n11199), .C2(n11198), .A(n15092), .B(n11711), .ZN(
        n11205) );
  AOI22_X1 U13868 ( .A1(n14228), .A2(n15097), .B1(n15107), .B2(n14499), .ZN(
        n11202) );
  MUX2_X1 U13869 ( .A(n15119), .B(P1_STATE_REG_SCAN_IN), .S(
        P1_REG3_REG_3__SCAN_IN), .Z(n11201) );
  OAI211_X1 U13870 ( .C1(n11203), .C2(n15086), .A(n11202), .B(n11201), .ZN(
        n11204) );
  OR2_X1 U13871 ( .A1(n11205), .A2(n11204), .ZN(P1_U3218) );
  OAI21_X1 U13872 ( .B1(n14422), .B2(n11207), .A(n11206), .ZN(n11215) );
  OAI22_X1 U13873 ( .A1(n6811), .A2(n14947), .B1(n11208), .B2(n15131), .ZN(
        n11214) );
  OAI21_X1 U13874 ( .B1(n11211), .B2(n11210), .A(n11209), .ZN(n15285) );
  INV_X1 U13875 ( .A(n15285), .ZN(n11212) );
  NOR2_X1 U13876 ( .A1(n11212), .A2(n14928), .ZN(n11213) );
  AOI211_X1 U13877 ( .C1(n15160), .C2(n11215), .A(n11214), .B(n11213), .ZN(
        n15282) );
  INV_X1 U13878 ( .A(n11216), .ZN(n11218) );
  OAI211_X1 U13879 ( .C1(n15281), .C2(n11218), .A(n15122), .B(n11217), .ZN(
        n15280) );
  INV_X1 U13880 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n14524) );
  OAI22_X1 U13881 ( .A1(n14958), .A2(n15280), .B1(n14524), .B2(n15136), .ZN(
        n11219) );
  AOI21_X1 U13882 ( .B1(n14931), .B2(P1_REG2_REG_2__SCAN_IN), .A(n11219), .ZN(
        n11222) );
  AOI22_X1 U13883 ( .A1(n11220), .A2(n15285), .B1(n14717), .B2(n14224), .ZN(
        n11221) );
  OAI211_X1 U13884 ( .C1(n15282), .C2(n14765), .A(n11222), .B(n11221), .ZN(
        P1_U3291) );
  XNOR2_X1 U13885 ( .A(n13674), .B(P2_REG1_REG_12__SCAN_IN), .ZN(n11227) );
  NOR2_X1 U13886 ( .A1(n11223), .A2(n15537), .ZN(n11224) );
  OR2_X1 U13887 ( .A1(n11225), .A2(n11224), .ZN(n11226) );
  NOR3_X1 U13888 ( .A1(n11225), .A2(n11224), .A3(n11227), .ZN(n13686) );
  AOI21_X1 U13889 ( .B1(n11227), .B2(n11226), .A(n13686), .ZN(n11237) );
  NAND2_X1 U13890 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3088), .ZN(n12114)
         );
  OAI21_X1 U13891 ( .B1(n13722), .B2(n7180), .A(n12114), .ZN(n11228) );
  AOI21_X1 U13892 ( .B1(n13674), .B2(n15453), .A(n11228), .ZN(n11236) );
  NOR2_X1 U13893 ( .A1(n11229), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n11230) );
  MUX2_X1 U13894 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n11960), .S(n13674), .Z(
        n11231) );
  INV_X1 U13895 ( .A(n13673), .ZN(n11234) );
  NOR3_X1 U13896 ( .A1(n11232), .A2(n11231), .A3(n11230), .ZN(n11233) );
  OAI21_X1 U13897 ( .B1(n11234), .B2(n11233), .A(n15450), .ZN(n11235) );
  OAI211_X1 U13898 ( .C1(n11237), .C2(n15375), .A(n11236), .B(n11235), .ZN(
        P2_U3226) );
  OAI211_X1 U13899 ( .C1(n11240), .C2(n11239), .A(n11238), .B(n12788), .ZN(
        n11246) );
  INV_X1 U13900 ( .A(n11673), .ZN(n11243) );
  AOI21_X1 U13901 ( .B1(n9897), .B2(n12021), .A(n11241), .ZN(n11242) );
  OAI21_X1 U13902 ( .B1(n11243), .B2(n12774), .A(n11242), .ZN(n11244) );
  AOI21_X1 U13903 ( .B1(n12770), .B2(n15698), .A(n11244), .ZN(n11245) );
  OAI211_X1 U13904 ( .C1(P3_REG3_REG_3__SCAN_IN), .C2(n12440), .A(n11246), .B(
        n11245), .ZN(P3_U3158) );
  INV_X1 U13905 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n15170) );
  INV_X1 U13906 ( .A(n11718), .ZN(n11723) );
  AOI22_X1 U13907 ( .A1(n11718), .A2(n15170), .B1(P1_REG1_REG_14__SCAN_IN), 
        .B2(n11723), .ZN(n11249) );
  OAI21_X1 U13908 ( .B1(n11255), .B2(n10893), .A(n11247), .ZN(n11248) );
  NOR2_X1 U13909 ( .A1(n11249), .A2(n11248), .ZN(n11722) );
  AOI21_X1 U13910 ( .B1(n11249), .B2(n11248), .A(n11722), .ZN(n11260) );
  NAND2_X1 U13911 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n15098)
         );
  OAI21_X1 U13912 ( .B1(n15270), .B2(n11250), .A(n15098), .ZN(n11251) );
  AOI21_X1 U13913 ( .B1(n11718), .B2(n15232), .A(n11251), .ZN(n11259) );
  INV_X1 U13914 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n11252) );
  MUX2_X1 U13915 ( .A(n11252), .B(P1_REG2_REG_14__SCAN_IN), .S(n11718), .Z(
        n11253) );
  INV_X1 U13916 ( .A(n11253), .ZN(n11257) );
  OAI21_X1 U13917 ( .B1(n11255), .B2(n10883), .A(n11254), .ZN(n11256) );
  NAND2_X1 U13918 ( .A1(n11257), .A2(n11256), .ZN(n11719) );
  OAI211_X1 U13919 ( .C1(n11257), .C2(n11256), .A(n15258), .B(n11719), .ZN(
        n11258) );
  OAI211_X1 U13920 ( .C1(n11260), .C2(n15243), .A(n11259), .B(n11258), .ZN(
        P1_U3257) );
  XNOR2_X1 U13921 ( .A(n11400), .B(n13498), .ZN(n11411) );
  NAND2_X1 U13922 ( .A1(n13654), .A2(n13912), .ZN(n11410) );
  XNOR2_X1 U13923 ( .A(n11411), .B(n11410), .ZN(n11276) );
  INV_X1 U13924 ( .A(n11263), .ZN(n11264) );
  OR2_X1 U13925 ( .A1(n11265), .A2(n11264), .ZN(n11266) );
  XNOR2_X1 U13926 ( .A(n13515), .B(n13537), .ZN(n11267) );
  AND2_X1 U13927 ( .A1(n13655), .A2(n8410), .ZN(n11268) );
  NAND2_X1 U13928 ( .A1(n11267), .A2(n11268), .ZN(n11273) );
  INV_X1 U13929 ( .A(n11267), .ZN(n11270) );
  INV_X1 U13930 ( .A(n11268), .ZN(n11269) );
  NAND2_X1 U13931 ( .A1(n11270), .A2(n11269), .ZN(n11271) );
  NAND2_X1 U13932 ( .A1(n11273), .A2(n11271), .ZN(n13510) );
  INV_X1 U13933 ( .A(n11412), .ZN(n11435) );
  AOI21_X1 U13934 ( .B1(n11276), .B2(n11275), .A(n11435), .ZN(n11287) );
  INV_X1 U13935 ( .A(n11402), .ZN(n11285) );
  INV_X1 U13936 ( .A(n11277), .ZN(n11278) );
  OR2_X1 U13937 ( .A1(n11279), .A2(n11278), .ZN(n11280) );
  INV_X1 U13938 ( .A(n13607), .ZN(n13623) );
  INV_X1 U13939 ( .A(n11400), .ZN(n11283) );
  AOI22_X1 U13940 ( .A1(n13605), .A2(n11281), .B1(P2_REG3_REG_4__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11282) );
  OAI21_X1 U13941 ( .B1(n13597), .B2(n11283), .A(n11282), .ZN(n11284) );
  AOI21_X1 U13942 ( .B1(n11285), .B2(n13623), .A(n11284), .ZN(n11286) );
  OAI21_X1 U13943 ( .B1(n11287), .B2(n13627), .A(n11286), .ZN(P2_U3202) );
  NAND2_X1 U13944 ( .A1(n15143), .A2(n14619), .ZN(n11628) );
  INV_X1 U13945 ( .A(n11628), .ZN(n11288) );
  AOI21_X1 U13946 ( .B1(n15122), .B2(n11288), .A(n14717), .ZN(n11295) );
  OAI22_X1 U13947 ( .A1(n14931), .A2(n11290), .B1(n11289), .B2(n15136), .ZN(
        n11292) );
  NAND2_X1 U13948 ( .A1(n15143), .A2(n15160), .ZN(n14959) );
  AOI21_X1 U13949 ( .B1(n14750), .B2(n14959), .A(n14219), .ZN(n11291) );
  AOI211_X1 U13950 ( .C1(n14765), .C2(P1_REG2_REG_0__SCAN_IN), .A(n11292), .B(
        n11291), .ZN(n11293) );
  OAI21_X1 U13951 ( .B1(n11295), .B2(n11294), .A(n11293), .ZN(P1_U3293) );
  INV_X1 U13952 ( .A(n15611), .ZN(n15630) );
  XNOR2_X1 U13953 ( .A(n15542), .B(n11296), .ZN(n11311) );
  NAND2_X1 U13954 ( .A1(n11298), .A2(n11297), .ZN(n11299) );
  AND2_X1 U13955 ( .A1(n11300), .A2(n11299), .ZN(n11309) );
  NAND2_X1 U13956 ( .A1(n11301), .A2(n8469), .ZN(n11302) );
  NAND2_X1 U13957 ( .A1(n11303), .A2(n11302), .ZN(n11304) );
  NAND2_X1 U13958 ( .A1(n15032), .A2(n11304), .ZN(n11308) );
  NOR2_X1 U13959 ( .A1(n11305), .A2(P3_STATE_REG_SCAN_IN), .ZN(n11306) );
  AOI21_X1 U13960 ( .B1(n15623), .B2(P3_ADDR_REG_1__SCAN_IN), .A(n11306), .ZN(
        n11307) );
  OAI211_X1 U13961 ( .C1(n11309), .C2(n15541), .A(n11308), .B(n11307), .ZN(
        n11310) );
  AOI21_X1 U13962 ( .B1(n15630), .B2(n11311), .A(n11310), .ZN(n11312) );
  OAI21_X1 U13963 ( .B1(n11313), .B2(n15626), .A(n11312), .ZN(P3_U3183) );
  OAI22_X1 U13964 ( .A1(n11316), .A2(n11315), .B1(n11314), .B2(n11327), .ZN(
        n11318) );
  MUX2_X1 U13965 ( .A(P3_REG2_REG_8__SCAN_IN), .B(P3_REG1_REG_8__SCAN_IN), .S(
        n13027), .Z(n11854) );
  XNOR2_X1 U13966 ( .A(n11854), .B(n11325), .ZN(n11317) );
  NAND2_X1 U13967 ( .A1(n11318), .A2(n11317), .ZN(n11855) );
  OAI21_X1 U13968 ( .B1(n11318), .B2(n11317), .A(n11855), .ZN(n11319) );
  NAND2_X1 U13969 ( .A1(n11319), .A2(n15630), .ZN(n11339) );
  NOR2_X1 U13970 ( .A1(n11321), .A2(n11320), .ZN(n11322) );
  NAND2_X1 U13971 ( .A1(P3_REG2_REG_8__SCAN_IN), .A2(n11853), .ZN(n11324) );
  OAI21_X1 U13972 ( .B1(P3_REG2_REG_8__SCAN_IN), .B2(n11853), .A(n11324), .ZN(
        n11840) );
  XNOR2_X1 U13973 ( .A(n11841), .B(n11840), .ZN(n11337) );
  AOI22_X1 U13974 ( .A1(P3_REG1_REG_8__SCAN_IN), .A2(n11853), .B1(n11325), 
        .B2(n8579), .ZN(n11331) );
  NAND2_X1 U13975 ( .A1(n11327), .A2(n11326), .ZN(n11329) );
  OAI21_X1 U13976 ( .B1(n11331), .B2(n11330), .A(n11846), .ZN(n11332) );
  NAND2_X1 U13977 ( .A1(n11332), .A2(n15628), .ZN(n11335) );
  NOR2_X1 U13978 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11333), .ZN(n11833) );
  AOI21_X1 U13979 ( .B1(n15623), .B2(P3_ADDR_REG_8__SCAN_IN), .A(n11833), .ZN(
        n11334) );
  OAI211_X1 U13980 ( .C1(n15626), .C2(n11853), .A(n11335), .B(n11334), .ZN(
        n11336) );
  AOI21_X1 U13981 ( .B1(n15032), .B2(n11337), .A(n11336), .ZN(n11338) );
  NAND2_X1 U13982 ( .A1(n11339), .A2(n11338), .ZN(P3_U3190) );
  XNOR2_X1 U13983 ( .A(n14233), .B(n14499), .ZN(n14420) );
  XOR2_X1 U13984 ( .A(n11340), .B(n14420), .Z(n15291) );
  OAI211_X1 U13985 ( .C1(n11341), .C2(n15288), .A(n11471), .B(n15122), .ZN(
        n15287) );
  INV_X1 U13986 ( .A(n15136), .ZN(n14929) );
  AOI22_X1 U13987 ( .A1(n14717), .A2(n14233), .B1(n11716), .B2(n14929), .ZN(
        n11342) );
  OAI21_X1 U13988 ( .B1(n14958), .B2(n15287), .A(n11342), .ZN(n11348) );
  XNOR2_X1 U13989 ( .A(n11343), .B(n14420), .ZN(n11344) );
  NAND2_X1 U13990 ( .A1(n11344), .A2(n15160), .ZN(n11346) );
  AOI22_X1 U13991 ( .A1(n15134), .A2(n14498), .B1(n14762), .B2(n14500), .ZN(
        n11345) );
  NAND2_X1 U13992 ( .A1(n11346), .A2(n11345), .ZN(n15289) );
  MUX2_X1 U13993 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n15289), .S(n15143), .Z(
        n11347) );
  AOI211_X1 U13994 ( .C1(n15126), .C2(n15291), .A(n11348), .B(n11347), .ZN(
        n11349) );
  INV_X1 U13995 ( .A(n11349), .ZN(P1_U3289) );
  INV_X1 U13996 ( .A(n11350), .ZN(n11352) );
  INV_X1 U13997 ( .A(n15417), .ZN(n13691) );
  OAI222_X1 U13998 ( .A1(n14072), .A2(n11351), .B1(n14083), .B2(n11352), .C1(
        n13691), .C2(P2_U3088), .ZN(P2_U3313) );
  OAI222_X1 U13999 ( .A1(n14869), .A2(n11353), .B1(n14885), .B2(n11352), .C1(
        n11723), .C2(P1_U3086), .ZN(P1_U3341) );
  NAND2_X1 U14000 ( .A1(n13146), .A2(P3_U3897), .ZN(n11354) );
  OAI21_X1 U14001 ( .B1(P3_U3897), .B2(n11355), .A(n11354), .ZN(P3_U3514) );
  INV_X1 U14002 ( .A(n11356), .ZN(n11361) );
  NAND2_X1 U14003 ( .A1(n11357), .A2(n11360), .ZN(n11358) );
  OAI211_X1 U14004 ( .C1(n11361), .C2(n11360), .A(n11359), .B(n11358), .ZN(
        n11363) );
  OR2_X1 U14005 ( .A1(n11363), .A2(n15689), .ZN(n15053) );
  OAI22_X1 U14006 ( .A1(n15693), .A2(n10911), .B1(n11364), .B2(n15675), .ZN(
        n11365) );
  AOI21_X1 U14007 ( .B1(n15693), .B2(n11366), .A(n11365), .ZN(n11367) );
  OAI21_X1 U14008 ( .B1(n11368), .B2(n13297), .A(n11367), .ZN(P3_U3233) );
  OAI21_X1 U14009 ( .B1(n11370), .B2(n12821), .A(n11369), .ZN(n11371) );
  INV_X1 U14010 ( .A(n11371), .ZN(n12024) );
  INV_X1 U14011 ( .A(n15739), .ZN(n15065) );
  OAI211_X1 U14012 ( .C1(n11374), .C2(n11373), .A(n11372), .B(n15703), .ZN(
        n11376) );
  AOI22_X1 U14013 ( .A1(n15700), .A2(n15698), .B1(n11673), .B2(n15697), .ZN(
        n11375) );
  AND2_X1 U14014 ( .A1(n11376), .A2(n11375), .ZN(n12019) );
  OAI21_X1 U14015 ( .B1(n12024), .B2(n15065), .A(n12019), .ZN(n11381) );
  AOI21_X1 U14016 ( .B1(n11381), .B2(n15741), .A(n11377), .ZN(n11378) );
  INV_X1 U14017 ( .A(n11378), .ZN(P3_U3399) );
  INV_X1 U14018 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n11379) );
  AOI21_X1 U14019 ( .B1(n11381), .B2(n15751), .A(n11380), .ZN(n11382) );
  INV_X1 U14020 ( .A(n11382), .ZN(P3_U3462) );
  NAND2_X1 U14021 ( .A1(n11384), .A2(n11383), .ZN(n11385) );
  INV_X1 U14022 ( .A(n11493), .ZN(n11386) );
  NAND2_X1 U14023 ( .A1(n11052), .A2(n11386), .ZN(n11387) );
  INV_X2 U14024 ( .A(n13926), .ZN(n13919) );
  NAND2_X1 U14025 ( .A1(n13919), .A2(n13718), .ZN(n13922) );
  NOR2_X1 U14026 ( .A1(n13922), .A2(n11388), .ZN(n11393) );
  INV_X1 U14027 ( .A(n11389), .ZN(n11390) );
  NAND2_X1 U14028 ( .A1(n13933), .A2(n13515), .ZN(n11391) );
  OAI21_X1 U14029 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(n13916), .A(n11391), .ZN(
        n11392) );
  AOI211_X1 U14030 ( .C1(n13924), .C2(n11394), .A(n11393), .B(n11392), .ZN(
        n11398) );
  MUX2_X1 U14031 ( .A(n11396), .B(n11395), .S(n13919), .Z(n11397) );
  NAND2_X1 U14032 ( .A1(n11398), .A2(n11397), .ZN(P2_U3262) );
  NOR2_X1 U14033 ( .A1(n13922), .A2(n11399), .ZN(n11404) );
  NAND2_X1 U14034 ( .A1(n13933), .A2(n11400), .ZN(n11401) );
  OAI21_X1 U14035 ( .B1(n13916), .B2(n11402), .A(n11401), .ZN(n11403) );
  AOI211_X1 U14036 ( .C1(n13924), .C2(n11405), .A(n11404), .B(n11403), .ZN(
        n11409) );
  MUX2_X1 U14037 ( .A(n11407), .B(n11406), .S(n13919), .Z(n11408) );
  NAND2_X1 U14038 ( .A1(n11409), .A2(n11408), .ZN(P2_U3261) );
  NAND2_X1 U14039 ( .A1(n11411), .A2(n11410), .ZN(n11432) );
  NAND2_X1 U14040 ( .A1(n11412), .A2(n11432), .ZN(n11413) );
  XNOR2_X1 U14041 ( .A(n11523), .B(n13485), .ZN(n11414) );
  NAND2_X1 U14042 ( .A1(n13653), .A2(n13912), .ZN(n11415) );
  XNOR2_X1 U14043 ( .A(n11414), .B(n11415), .ZN(n11433) );
  NAND2_X1 U14044 ( .A1(n11413), .A2(n11433), .ZN(n11436) );
  INV_X1 U14045 ( .A(n11414), .ZN(n11416) );
  NAND2_X1 U14046 ( .A1(n11416), .A2(n11415), .ZN(n11417) );
  XNOR2_X1 U14047 ( .A(n11429), .B(n13537), .ZN(n11418) );
  AND2_X1 U14048 ( .A1(n13652), .A2(n8410), .ZN(n11419) );
  NAND2_X1 U14049 ( .A1(n11418), .A2(n11419), .ZN(n11500) );
  INV_X1 U14050 ( .A(n11418), .ZN(n11421) );
  INV_X1 U14051 ( .A(n11419), .ZN(n11420) );
  NAND2_X1 U14052 ( .A1(n11421), .A2(n11420), .ZN(n11422) );
  NAND2_X1 U14053 ( .A1(n11500), .A2(n11422), .ZN(n11424) );
  AOI21_X1 U14054 ( .B1(n11423), .B2(n11424), .A(n13627), .ZN(n11426) );
  NAND2_X1 U14055 ( .A1(n11426), .A2(n11501), .ZN(n11431) );
  AOI22_X1 U14056 ( .A1(n13602), .A2(n13651), .B1(n13617), .B2(n13653), .ZN(
        n11579) );
  OAI21_X1 U14057 ( .B1(n13621), .B2(n11579), .A(n11427), .ZN(n11428) );
  AOI21_X1 U14058 ( .B1(n11429), .B2(n13624), .A(n11428), .ZN(n11430) );
  OAI211_X1 U14059 ( .C1(n13607), .C2(n11585), .A(n11431), .B(n11430), .ZN(
        P2_U3211) );
  INV_X1 U14060 ( .A(n11432), .ZN(n11434) );
  NOR3_X1 U14061 ( .A1(n11435), .A2(n11434), .A3(n11433), .ZN(n11438) );
  INV_X1 U14062 ( .A(n11436), .ZN(n11437) );
  OAI21_X1 U14063 ( .B1(n11438), .B2(n11437), .A(n13591), .ZN(n11442) );
  AOI22_X1 U14064 ( .A1(n13602), .A2(n13652), .B1(n13617), .B2(n13654), .ZN(
        n11527) );
  OAI21_X1 U14065 ( .B1(n13621), .B2(n11527), .A(n11439), .ZN(n11440) );
  AOI21_X1 U14066 ( .B1(n11523), .B2(n13624), .A(n11440), .ZN(n11441) );
  OAI211_X1 U14067 ( .C1(n13607), .C2(n11521), .A(n11442), .B(n11441), .ZN(
        P2_U3199) );
  XNOR2_X1 U14068 ( .A(n11443), .B(n14426), .ZN(n15301) );
  XNOR2_X1 U14069 ( .A(n11444), .B(n14426), .ZN(n11447) );
  OAI22_X1 U14070 ( .A1(n12124), .A2(n14947), .B1(n11445), .B2(n15131), .ZN(
        n11446) );
  AOI21_X1 U14071 ( .B1(n11447), .B2(n15160), .A(n11446), .ZN(n11448) );
  OAI21_X1 U14072 ( .B1(n15301), .B2(n14928), .A(n11448), .ZN(n15304) );
  NAND2_X1 U14073 ( .A1(n15304), .A2(n15143), .ZN(n11455) );
  INV_X1 U14074 ( .A(n11939), .ZN(n11449) );
  OAI22_X1 U14075 ( .A1(n15143), .A2(n10583), .B1(n11449), .B2(n15136), .ZN(
        n11453) );
  INV_X1 U14076 ( .A(n11472), .ZN(n11451) );
  INV_X1 U14077 ( .A(n11450), .ZN(n11485) );
  OAI211_X1 U14078 ( .C1(n15303), .C2(n11451), .A(n11485), .B(n15122), .ZN(
        n15302) );
  NOR2_X1 U14079 ( .A1(n15302), .A2(n11628), .ZN(n11452) );
  AOI211_X1 U14080 ( .C1(n14717), .C2(n14250), .A(n11453), .B(n11452), .ZN(
        n11454) );
  OAI211_X1 U14081 ( .C1(n15301), .C2(n14921), .A(n11455), .B(n11454), .ZN(
        P1_U3287) );
  XOR2_X1 U14082 ( .A(n11457), .B(n11456), .Z(n11463) );
  OAI22_X1 U14083 ( .A1(n11459), .A2(n13597), .B1(n13621), .B2(n11458), .ZN(
        n11460) );
  AOI21_X1 U14084 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(n11461), .A(n11460), .ZN(
        n11462) );
  OAI21_X1 U14085 ( .B1(n11463), .B2(n13627), .A(n11462), .ZN(P2_U3194) );
  XNOR2_X1 U14086 ( .A(n11464), .B(n14425), .ZN(n15299) );
  INV_X1 U14087 ( .A(n15299), .ZN(n11478) );
  XNOR2_X1 U14088 ( .A(n11466), .B(n11465), .ZN(n11469) );
  NAND2_X1 U14089 ( .A1(n15134), .A2(n14497), .ZN(n11468) );
  NAND2_X1 U14090 ( .A1(n14762), .A2(n14499), .ZN(n11467) );
  NAND2_X1 U14091 ( .A1(n11468), .A2(n11467), .ZN(n11745) );
  AOI21_X1 U14092 ( .B1(n11469), .B2(n15160), .A(n11745), .ZN(n15297) );
  MUX2_X1 U14093 ( .A(n11470), .B(n15297), .S(n15143), .Z(n11477) );
  AOI21_X1 U14094 ( .B1(n11471), .B2(n15293), .A(n14741), .ZN(n11473) );
  NAND2_X1 U14095 ( .A1(n11473), .A2(n11472), .ZN(n15295) );
  INV_X1 U14096 ( .A(n15295), .ZN(n11475) );
  INV_X1 U14097 ( .A(n15293), .ZN(n11747) );
  OAI22_X1 U14098 ( .A1(n15141), .A2(n11747), .B1(n11744), .B2(n15136), .ZN(
        n11474) );
  AOI21_X1 U14099 ( .B1(n15125), .B2(n11475), .A(n11474), .ZN(n11476) );
  OAI211_X1 U14100 ( .C1(n14750), .C2(n11478), .A(n11477), .B(n11476), .ZN(
        P1_U3288) );
  XNOR2_X1 U14101 ( .A(n11479), .B(n14427), .ZN(n15314) );
  XNOR2_X1 U14102 ( .A(n11480), .B(n14427), .ZN(n11483) );
  NAND2_X1 U14103 ( .A1(n15134), .A2(n14495), .ZN(n11482) );
  NAND2_X1 U14104 ( .A1(n14762), .A2(n14497), .ZN(n11481) );
  NAND2_X1 U14105 ( .A1(n11482), .A2(n11481), .ZN(n12128) );
  AOI21_X1 U14106 ( .B1(n11483), .B2(n15160), .A(n12128), .ZN(n15312) );
  MUX2_X1 U14107 ( .A(n11484), .B(n15312), .S(n15143), .Z(n11489) );
  AOI211_X1 U14108 ( .C1(n15309), .C2(n11485), .A(n14741), .B(n11624), .ZN(
        n15308) );
  INV_X1 U14109 ( .A(n11486), .ZN(n12131) );
  OAI22_X1 U14110 ( .A1(n15141), .A2(n12127), .B1(n12131), .B2(n15136), .ZN(
        n11487) );
  AOI21_X1 U14111 ( .B1(n15308), .B2(n15125), .A(n11487), .ZN(n11488) );
  OAI211_X1 U14112 ( .C1(n14750), .C2(n15314), .A(n11489), .B(n11488), .ZN(
        P1_U3286) );
  INV_X1 U14113 ( .A(n11490), .ZN(n11492) );
  NOR2_X1 U14114 ( .A1(n11492), .A2(n11491), .ZN(n15473) );
  AND2_X1 U14115 ( .A1(n13919), .A2(n11493), .ZN(n13928) );
  AOI22_X1 U14116 ( .A1(n13930), .A2(n15473), .B1(n13928), .B2(n15474), .ZN(
        n11499) );
  INV_X1 U14117 ( .A(n15473), .ZN(n11496) );
  NAND2_X1 U14118 ( .A1(n13896), .A2(n11052), .ZN(n11495) );
  AOI21_X1 U14119 ( .B1(n15474), .B2(n11495), .A(n11494), .ZN(n15471) );
  OAI21_X1 U14120 ( .B1(n12137), .B2(n11496), .A(n15471), .ZN(n11497) );
  INV_X1 U14121 ( .A(n13916), .ZN(n13931) );
  AOI22_X1 U14122 ( .A1(n13919), .A2(n11497), .B1(P2_REG3_REG_0__SCAN_IN), 
        .B2(n13931), .ZN(n11498) );
  OAI211_X1 U14123 ( .C1(n10712), .C2(n13919), .A(n11499), .B(n11498), .ZN(
        P2_U3265) );
  XNOR2_X1 U14124 ( .A(n11594), .B(n13485), .ZN(n11502) );
  AND2_X1 U14125 ( .A1(n13651), .A2(n13912), .ZN(n11503) );
  NAND2_X1 U14126 ( .A1(n11502), .A2(n11503), .ZN(n11660) );
  INV_X1 U14127 ( .A(n11502), .ZN(n11505) );
  INV_X1 U14128 ( .A(n11503), .ZN(n11504) );
  NAND2_X1 U14129 ( .A1(n11505), .A2(n11504), .ZN(n11506) );
  AND2_X1 U14130 ( .A1(n11660), .A2(n11506), .ZN(n11507) );
  OAI211_X1 U14131 ( .C1(n11508), .C2(n11507), .A(n11661), .B(n13591), .ZN(
        n11512) );
  AOI22_X1 U14132 ( .A1(n13602), .A2(n13650), .B1(n13617), .B2(n13652), .ZN(
        n11601) );
  OAI21_X1 U14133 ( .B1(n13621), .B2(n11601), .A(n11509), .ZN(n11510) );
  AOI21_X1 U14134 ( .B1(n11594), .B2(n13624), .A(n11510), .ZN(n11511) );
  OAI211_X1 U14135 ( .C1(n13607), .C2(n11595), .A(n11512), .B(n11511), .ZN(
        P2_U3185) );
  INV_X1 U14136 ( .A(n11513), .ZN(n11516) );
  OAI222_X1 U14137 ( .A1(n12666), .A2(n11516), .B1(n13440), .B2(n11515), .C1(
        P3_U3151), .C2(n11514), .ZN(P3_U3275) );
  XOR2_X1 U14138 ( .A(n11526), .B(n11517), .Z(n15479) );
  INV_X1 U14139 ( .A(n11518), .ZN(n11520) );
  INV_X1 U14140 ( .A(n11583), .ZN(n11519) );
  OAI211_X1 U14141 ( .C1(n15476), .C2(n11520), .A(n11519), .B(n11777), .ZN(
        n15475) );
  INV_X1 U14142 ( .A(n11521), .ZN(n11522) );
  AOI22_X1 U14143 ( .A1(n13933), .A2(n11523), .B1(n13931), .B2(n11522), .ZN(
        n11524) );
  OAI21_X1 U14144 ( .B1(n13922), .B2(n15475), .A(n11524), .ZN(n11530) );
  XOR2_X1 U14145 ( .A(n11526), .B(n11525), .Z(n11528) );
  OAI21_X1 U14146 ( .B1(n11528), .B2(n13896), .A(n11527), .ZN(n15477) );
  MUX2_X1 U14147 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n15477), .S(n13919), .Z(
        n11529) );
  AOI211_X1 U14148 ( .C1(n13924), .C2(n15479), .A(n11530), .B(n11529), .ZN(
        n11531) );
  INV_X1 U14149 ( .A(n11531), .ZN(P2_U3260) );
  NAND2_X1 U14150 ( .A1(n13160), .A2(P3_U3897), .ZN(n11532) );
  OAI21_X1 U14151 ( .B1(P3_U3897), .B2(n11533), .A(n11532), .ZN(P3_U3515) );
  INV_X1 U14152 ( .A(n11534), .ZN(n11535) );
  AOI21_X1 U14153 ( .B1(n11537), .B2(n11536), .A(n11535), .ZN(n11543) );
  AOI21_X1 U14154 ( .B1(n9897), .B2(n15672), .A(n11538), .ZN(n11539) );
  OAI21_X1 U14155 ( .B1(n11790), .B2(n12774), .A(n11539), .ZN(n11541) );
  NOR2_X1 U14156 ( .A1(n12440), .A2(n15676), .ZN(n11540) );
  AOI211_X1 U14157 ( .C1(n12770), .C2(n15681), .A(n11541), .B(n11540), .ZN(
        n11542) );
  OAI21_X1 U14158 ( .B1(n11543), .B2(n12777), .A(n11542), .ZN(P3_U3170) );
  OAI222_X1 U14159 ( .A1(n12666), .A2(n11545), .B1(n13440), .B2(n11544), .C1(
        P3_U3151), .C2(n11681), .ZN(P3_U3274) );
  INV_X1 U14160 ( .A(n11546), .ZN(n11548) );
  INV_X1 U14161 ( .A(n12004), .ZN(n11726) );
  OAI222_X1 U14162 ( .A1(n14869), .A2(n11547), .B1(n14885), .B2(n11548), .C1(
        P1_U3086), .C2(n11726), .ZN(P1_U3340) );
  INV_X1 U14163 ( .A(n15426), .ZN(n13694) );
  OAI222_X1 U14164 ( .A1(n14072), .A2(n11549), .B1(n14083), .B2(n11548), .C1(
        P2_U3088), .C2(n13694), .ZN(P2_U3312) );
  OAI22_X1 U14165 ( .A1(n13919), .A2(n10525), .B1(n11550), .B2(n13916), .ZN(
        n11553) );
  NOR2_X1 U14166 ( .A1(n13824), .A2(n11551), .ZN(n11552) );
  AOI211_X1 U14167 ( .C1(n11554), .C2(n13930), .A(n11553), .B(n11552), .ZN(
        n11557) );
  NAND2_X1 U14168 ( .A1(n13924), .A2(n11555), .ZN(n11556) );
  OAI211_X1 U14169 ( .C1(n13926), .C2(n11558), .A(n11557), .B(n11556), .ZN(
        P2_U3263) );
  OAI21_X1 U14170 ( .B1(n11560), .B2(n12863), .A(n11559), .ZN(n11561) );
  INV_X1 U14171 ( .A(n11561), .ZN(n15669) );
  OAI211_X1 U14172 ( .C1(n11564), .C2(n11563), .A(n11562), .B(n15703), .ZN(
        n11566) );
  AOI22_X1 U14173 ( .A1(n15700), .A2(n15681), .B1(n12995), .B2(n15697), .ZN(
        n11565) );
  AND2_X1 U14174 ( .A1(n11566), .A2(n11565), .ZN(n15667) );
  OAI21_X1 U14175 ( .B1(n15669), .B2(n15065), .A(n15667), .ZN(n11571) );
  OAI22_X1 U14176 ( .A1(n11569), .A2(n13424), .B1(n15741), .B2(n8509), .ZN(
        n11567) );
  AOI21_X1 U14177 ( .B1(n11571), .B2(n15741), .A(n11567), .ZN(n11568) );
  INV_X1 U14178 ( .A(n11568), .ZN(P3_U3402) );
  OAI22_X1 U14179 ( .A1(n13367), .A2(n11569), .B1(n15751), .B2(n10981), .ZN(
        n11570) );
  AOI21_X1 U14180 ( .B1(n11571), .B2(n15751), .A(n11570), .ZN(n11572) );
  INV_X1 U14181 ( .A(n11572), .ZN(P3_U3463) );
  NAND2_X1 U14182 ( .A1(n11573), .A2(n11576), .ZN(n11574) );
  NAND2_X1 U14183 ( .A1(n11575), .A2(n11574), .ZN(n15480) );
  XNOR2_X1 U14184 ( .A(n11577), .B(n11576), .ZN(n11578) );
  NAND2_X1 U14185 ( .A1(n11578), .A2(n13906), .ZN(n11580) );
  NAND2_X1 U14186 ( .A1(n11580), .A2(n11579), .ZN(n15483) );
  INV_X1 U14187 ( .A(n15483), .ZN(n11581) );
  MUX2_X1 U14188 ( .A(n11582), .B(n11581), .S(n13919), .Z(n11589) );
  OAI21_X1 U14189 ( .B1(n11583), .B2(n15482), .A(n11777), .ZN(n11584) );
  OR2_X1 U14190 ( .A1(n11584), .A2(n11593), .ZN(n15481) );
  INV_X1 U14191 ( .A(n15481), .ZN(n11587) );
  OAI22_X1 U14192 ( .A1(n13824), .A2(n15482), .B1(n13916), .B2(n11585), .ZN(
        n11586) );
  AOI21_X1 U14193 ( .B1(n13930), .B2(n11587), .A(n11586), .ZN(n11588) );
  OAI211_X1 U14194 ( .C1(n13902), .C2(n15480), .A(n11589), .B(n11588), .ZN(
        P2_U3259) );
  OAI21_X1 U14195 ( .B1(n11591), .B2(n11599), .A(n11590), .ZN(n11592) );
  INV_X1 U14196 ( .A(n11592), .ZN(n15492) );
  OAI211_X1 U14197 ( .C1(n11593), .C2(n15488), .A(n11777), .B(n11635), .ZN(
        n15487) );
  NAND2_X1 U14198 ( .A1(n13933), .A2(n11594), .ZN(n11598) );
  INV_X1 U14199 ( .A(n11595), .ZN(n11596) );
  NAND2_X1 U14200 ( .A1(n13931), .A2(n11596), .ZN(n11597) );
  OAI211_X1 U14201 ( .C1(n15487), .C2(n13922), .A(n11598), .B(n11597), .ZN(
        n11604) );
  XNOR2_X1 U14202 ( .A(n11600), .B(n11599), .ZN(n11602) );
  OAI21_X1 U14203 ( .B1(n11602), .B2(n13896), .A(n11601), .ZN(n15489) );
  MUX2_X1 U14204 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n15489), .S(n13919), .Z(
        n11603) );
  AOI211_X1 U14205 ( .C1(n13924), .C2(n15492), .A(n11604), .B(n11603), .ZN(
        n11605) );
  INV_X1 U14206 ( .A(n11605), .ZN(P2_U3258) );
  OAI21_X1 U14207 ( .B1(n11607), .B2(n11613), .A(n11606), .ZN(n15499) );
  NAND2_X1 U14208 ( .A1(n11755), .A2(n11636), .ZN(n11608) );
  NAND2_X1 U14209 ( .A1(n11608), .A2(n11777), .ZN(n11609) );
  NOR2_X1 U14210 ( .A1(n11776), .A2(n11609), .ZN(n15502) );
  INV_X1 U14211 ( .A(n11755), .ZN(n15500) );
  INV_X1 U14212 ( .A(n11610), .ZN(n11767) );
  AOI22_X1 U14213 ( .A1(n13926), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n11767), 
        .B2(n13931), .ZN(n11611) );
  OAI21_X1 U14214 ( .B1(n13824), .B2(n15500), .A(n11611), .ZN(n11612) );
  AOI21_X1 U14215 ( .B1(n15502), .B2(n13930), .A(n11612), .ZN(n11617) );
  XNOR2_X1 U14216 ( .A(n11614), .B(n11613), .ZN(n11615) );
  AOI22_X1 U14217 ( .A1(n13602), .A2(n13648), .B1(n13617), .B2(n13650), .ZN(
        n11765) );
  OAI21_X1 U14218 ( .B1(n11615), .B2(n13896), .A(n11765), .ZN(n15501) );
  NAND2_X1 U14219 ( .A1(n15501), .A2(n13919), .ZN(n11616) );
  OAI211_X1 U14220 ( .C1(n15499), .C2(n13902), .A(n11617), .B(n11616), .ZN(
        P2_U3256) );
  XNOR2_X1 U14221 ( .A(n11619), .B(n11618), .ZN(n15323) );
  INV_X1 U14222 ( .A(n15323), .ZN(n11631) );
  XNOR2_X1 U14223 ( .A(n11620), .B(n14429), .ZN(n11623) );
  NAND2_X1 U14224 ( .A1(n15134), .A2(n14494), .ZN(n11622) );
  NAND2_X1 U14225 ( .A1(n14762), .A2(n14496), .ZN(n11621) );
  AND2_X1 U14226 ( .A1(n11622), .A2(n11621), .ZN(n12171) );
  OAI21_X1 U14227 ( .B1(n11623), .B2(n15175), .A(n12171), .ZN(n15321) );
  OAI211_X1 U14228 ( .C1(n15320), .C2(n11624), .A(n15122), .B(n11915), .ZN(
        n15319) );
  INV_X1 U14229 ( .A(n12173), .ZN(n11625) );
  OAI22_X1 U14230 ( .A1(n15143), .A2(n10597), .B1(n11625), .B2(n15136), .ZN(
        n11626) );
  AOI21_X1 U14231 ( .B1(n14717), .B2(n14262), .A(n11626), .ZN(n11627) );
  OAI21_X1 U14232 ( .B1(n15319), .B2(n11628), .A(n11627), .ZN(n11629) );
  AOI21_X1 U14233 ( .B1(n15321), .B2(n15143), .A(n11629), .ZN(n11630) );
  OAI21_X1 U14234 ( .B1(n14750), .B2(n11631), .A(n11630), .ZN(P1_U3285) );
  NAND2_X1 U14235 ( .A1(n11632), .A2(P3_U3897), .ZN(n11633) );
  OAI21_X1 U14236 ( .B1(P3_U3897), .B2(n11634), .A(n11633), .ZN(P3_U3516) );
  AOI21_X1 U14237 ( .B1(n11635), .B2(n11662), .A(n13912), .ZN(n11637) );
  NAND2_X1 U14238 ( .A1(n11637), .A2(n11636), .ZN(n15493) );
  OR2_X1 U14239 ( .A1(n11639), .A2(n11638), .ZN(n11640) );
  AND2_X1 U14240 ( .A1(n11641), .A2(n11640), .ZN(n15496) );
  NAND2_X1 U14241 ( .A1(n15496), .A2(n13924), .ZN(n11644) );
  INV_X1 U14242 ( .A(n11642), .ZN(n11669) );
  AOI22_X1 U14243 ( .A1(n13933), .A2(n11662), .B1(n11669), .B2(n13931), .ZN(
        n11643) );
  OAI211_X1 U14244 ( .C1(n13922), .C2(n15493), .A(n11644), .B(n11643), .ZN(
        n11650) );
  XNOR2_X1 U14245 ( .A(n11646), .B(n11645), .ZN(n11647) );
  NAND2_X1 U14246 ( .A1(n11647), .A2(n13906), .ZN(n11648) );
  AOI22_X1 U14247 ( .A1(n13602), .A2(n13649), .B1(n13617), .B2(n13651), .ZN(
        n11667) );
  NAND2_X1 U14248 ( .A1(n11648), .A2(n11667), .ZN(n15495) );
  MUX2_X1 U14249 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n15495), .S(n13919), .Z(
        n11649) );
  OR2_X1 U14250 ( .A1(n11650), .A2(n11649), .ZN(P2_U3257) );
  XOR2_X1 U14251 ( .A(n11652), .B(n11651), .Z(n11659) );
  NAND2_X1 U14252 ( .A1(n12794), .A2(n11947), .ZN(n11655) );
  INV_X1 U14253 ( .A(n11653), .ZN(n11654) );
  OAI211_X1 U14254 ( .C1(n12797), .C2(n11682), .A(n11655), .B(n11654), .ZN(
        n11657) );
  NOR2_X1 U14255 ( .A1(n12440), .A2(n11683), .ZN(n11656) );
  AOI211_X1 U14256 ( .C1(n12770), .C2(n11673), .A(n11657), .B(n11656), .ZN(
        n11658) );
  OAI21_X1 U14257 ( .B1(n11659), .B2(n12777), .A(n11658), .ZN(P3_U3167) );
  XNOR2_X1 U14258 ( .A(n11662), .B(n13485), .ZN(n11752) );
  NAND2_X1 U14259 ( .A1(n13650), .A2(n8410), .ZN(n11753) );
  XNOR2_X1 U14260 ( .A(n11752), .B(n11753), .ZN(n11663) );
  OAI21_X1 U14261 ( .B1(n11664), .B2(n11663), .A(n11759), .ZN(n11665) );
  NAND2_X1 U14262 ( .A1(n11665), .A2(n13591), .ZN(n11671) );
  OAI21_X1 U14263 ( .B1(n13621), .B2(n11667), .A(n11666), .ZN(n11668) );
  AOI21_X1 U14264 ( .B1(n11669), .B2(n13623), .A(n11668), .ZN(n11670) );
  OAI211_X1 U14265 ( .C1(n7159), .C2(n13597), .A(n11671), .B(n11670), .ZN(
        P2_U3193) );
  XNOR2_X1 U14266 ( .A(n11672), .B(n6678), .ZN(n15722) );
  NAND2_X1 U14267 ( .A1(n15722), .A2(n15680), .ZN(n11680) );
  AOI22_X1 U14268 ( .A1(n15700), .A2(n11673), .B1(n11947), .B2(n15697), .ZN(
        n11679) );
  NAND2_X1 U14269 ( .A1(n11674), .A2(n6678), .ZN(n11675) );
  NAND2_X1 U14270 ( .A1(n11676), .A2(n11675), .ZN(n11677) );
  NAND2_X1 U14271 ( .A1(n11677), .A2(n15703), .ZN(n11678) );
  AND3_X1 U14272 ( .A1(n11680), .A2(n11679), .A3(n11678), .ZN(n15724) );
  OR2_X1 U14273 ( .A1(n11681), .A2(n15708), .ZN(n15690) );
  INV_X1 U14274 ( .A(n15690), .ZN(n12017) );
  AND2_X1 U14275 ( .A1(n15693), .A2(n12017), .ZN(n15711) );
  INV_X1 U14276 ( .A(n15053), .ZN(n15648) );
  NOR2_X1 U14277 ( .A1(n11682), .A2(n15730), .ZN(n15721) );
  INV_X1 U14278 ( .A(n11683), .ZN(n11684) );
  AOI22_X1 U14279 ( .A1(n15648), .A2(n15721), .B1(n15710), .B2(n11684), .ZN(
        n11685) );
  OAI21_X1 U14280 ( .B1(n8523), .B2(n15693), .A(n11685), .ZN(n11686) );
  AOI21_X1 U14281 ( .B1(n15722), .B2(n15711), .A(n11686), .ZN(n11687) );
  OAI21_X1 U14282 ( .B1(n15724), .B2(n13303), .A(n11687), .ZN(P3_U3228) );
  INV_X1 U14283 ( .A(n15436), .ZN(n13696) );
  INV_X1 U14284 ( .A(n11688), .ZN(n11690) );
  OAI222_X1 U14285 ( .A1(P2_U3088), .A2(n13696), .B1(n14083), .B2(n11690), 
        .C1(n11689), .C2(n14072), .ZN(P2_U3311) );
  INV_X1 U14286 ( .A(n12008), .ZN(n12145) );
  OAI222_X1 U14287 ( .A1(n14891), .A2(n11691), .B1(n14885), .B2(n11690), .C1(
        n12145), .C2(P1_U3086), .ZN(P1_U3339) );
  NOR2_X1 U14288 ( .A1(n13440), .A2(SI_22_), .ZN(n11692) );
  AOI21_X1 U14289 ( .B1(n11693), .B2(P3_STATE_REG_SCAN_IN), .A(n11692), .ZN(
        n11694) );
  OAI21_X1 U14290 ( .B1(n11695), .B2(n12666), .A(n11694), .ZN(n11696) );
  INV_X1 U14291 ( .A(n11696), .ZN(P3_U3273) );
  AOI21_X1 U14292 ( .B1(n11698), .B2(n11697), .A(n12777), .ZN(n11699) );
  OR2_X1 U14293 ( .A1(n11698), .A2(n11697), .ZN(n11816) );
  NAND2_X1 U14294 ( .A1(n11699), .A2(n11816), .ZN(n11704) );
  INV_X1 U14295 ( .A(n12031), .ZN(n11789) );
  AOI21_X1 U14296 ( .B1(n9897), .B2(n15664), .A(n11700), .ZN(n11701) );
  OAI21_X1 U14297 ( .B1(n11789), .B2(n12774), .A(n11701), .ZN(n11702) );
  AOI21_X1 U14298 ( .B1(n12770), .B2(n12995), .A(n11702), .ZN(n11703) );
  OAI211_X1 U14299 ( .C1(n15666), .C2(n12440), .A(n11704), .B(n11703), .ZN(
        P3_U3179) );
  INV_X1 U14300 ( .A(n15119), .ZN(n14205) );
  AOI22_X1 U14301 ( .A1(n15109), .A2(n14500), .B1(n15107), .B2(n14498), .ZN(
        n11705) );
  NAND2_X1 U14302 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n15237) );
  OAI211_X1 U14303 ( .C1(n15288), .C2(n15111), .A(n11705), .B(n15237), .ZN(
        n11715) );
  AOI22_X1 U14304 ( .A1(n14233), .A2(n12635), .B1(n12621), .B2(n14499), .ZN(
        n11706) );
  XNOR2_X1 U14305 ( .A(n11706), .B(n12646), .ZN(n11713) );
  INV_X1 U14306 ( .A(n11707), .ZN(n11710) );
  INV_X1 U14307 ( .A(n11708), .ZN(n11709) );
  AOI22_X1 U14308 ( .A1(n10728), .A2(n14499), .B1(n14233), .B2(n12621), .ZN(
        n11737) );
  AOI211_X1 U14309 ( .C1(n11713), .C2(n11712), .A(n15092), .B(n11741), .ZN(
        n11714) );
  AOI211_X1 U14310 ( .C1(n14205), .C2(n11716), .A(n11715), .B(n11714), .ZN(
        n11717) );
  INV_X1 U14311 ( .A(n11717), .ZN(P1_U3230) );
  NAND2_X1 U14312 ( .A1(n11718), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n11720) );
  NAND2_X1 U14313 ( .A1(n11720), .A2(n11719), .ZN(n11996) );
  XNOR2_X1 U14314 ( .A(n12004), .B(n11996), .ZN(n11721) );
  NOR2_X1 U14315 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n11721), .ZN(n11997) );
  AOI21_X1 U14316 ( .B1(P1_REG2_REG_15__SCAN_IN), .B2(n11721), .A(n11997), 
        .ZN(n11731) );
  AOI21_X1 U14317 ( .B1(n11723), .B2(n15170), .A(n11722), .ZN(n12003) );
  XNOR2_X1 U14318 ( .A(n12004), .B(n12003), .ZN(n11724) );
  NOR2_X1 U14319 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n11724), .ZN(n12005) );
  AOI21_X1 U14320 ( .B1(P1_REG1_REG_15__SCAN_IN), .B2(n11724), .A(n12005), 
        .ZN(n11725) );
  OR2_X1 U14321 ( .A1(n11725), .A2(n15243), .ZN(n11730) );
  NOR2_X1 U14322 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n14202), .ZN(n11728) );
  NOR2_X1 U14323 ( .A1(n15266), .A2(n11726), .ZN(n11727) );
  AOI211_X1 U14324 ( .C1(n14593), .C2(P1_ADDR_REG_15__SCAN_IN), .A(n11728), 
        .B(n11727), .ZN(n11729) );
  OAI211_X1 U14325 ( .C1(n11731), .C2(n15248), .A(n11730), .B(n11729), .ZN(
        P1_U3258) );
  INV_X1 U14326 ( .A(n11732), .ZN(n11734) );
  INV_X1 U14327 ( .A(n14605), .ZN(n12152) );
  OAI222_X1 U14328 ( .A1(n14891), .A2(n11733), .B1(n14885), .B2(n11734), .C1(
        n12152), .C2(P1_U3086), .ZN(P1_U3338) );
  INV_X1 U14329 ( .A(n15454), .ZN(n13697) );
  OAI222_X1 U14330 ( .A1(n14072), .A2(n11735), .B1(n14083), .B2(n11734), .C1(
        n13697), .C2(P2_U3088), .ZN(P2_U3310) );
  INV_X1 U14331 ( .A(n11736), .ZN(n11739) );
  INV_X1 U14332 ( .A(n11737), .ZN(n11738) );
  AOI22_X1 U14333 ( .A1(n15293), .A2(n12635), .B1(n12621), .B2(n14498), .ZN(
        n11742) );
  XNOR2_X1 U14334 ( .A(n11742), .B(n12646), .ZN(n11926) );
  AOI22_X1 U14335 ( .A1(n15293), .A2(n12621), .B1(n10728), .B2(n14498), .ZN(
        n11927) );
  XNOR2_X1 U14336 ( .A(n11926), .B(n7517), .ZN(n11743) );
  XNOR2_X1 U14337 ( .A(n11928), .B(n11743), .ZN(n11750) );
  NOR2_X1 U14338 ( .A1(n15119), .A2(n11744), .ZN(n11749) );
  NAND2_X1 U14339 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n14554) );
  NAND2_X1 U14340 ( .A1(n14195), .A2(n11745), .ZN(n11746) );
  OAI211_X1 U14341 ( .C1(n15111), .C2(n11747), .A(n14554), .B(n11746), .ZN(
        n11748) );
  AOI211_X1 U14342 ( .C1(n11750), .C2(n15114), .A(n11749), .B(n11748), .ZN(
        n11751) );
  INV_X1 U14343 ( .A(n11751), .ZN(P1_U3227) );
  INV_X1 U14344 ( .A(n11759), .ZN(n11757) );
  INV_X1 U14345 ( .A(n11752), .ZN(n11754) );
  NAND2_X1 U14346 ( .A1(n11754), .A2(n11753), .ZN(n11758) );
  INV_X1 U14347 ( .A(n11758), .ZN(n11756) );
  XNOR2_X1 U14348 ( .A(n11755), .B(n13485), .ZN(n11871) );
  NAND2_X1 U14349 ( .A1(n13649), .A2(n13912), .ZN(n11872) );
  XNOR2_X1 U14350 ( .A(n11871), .B(n11872), .ZN(n11760) );
  NOR3_X1 U14351 ( .A1(n11757), .A2(n11756), .A3(n11760), .ZN(n11763) );
  NAND2_X1 U14352 ( .A1(n11759), .A2(n11758), .ZN(n11761) );
  INV_X1 U14353 ( .A(n11875), .ZN(n11762) );
  OAI21_X1 U14354 ( .B1(n11763), .B2(n11762), .A(n13591), .ZN(n11769) );
  OAI22_X1 U14355 ( .A1(n13621), .A2(n11765), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11764), .ZN(n11766) );
  AOI21_X1 U14356 ( .B1(n11767), .B2(n13623), .A(n11766), .ZN(n11768) );
  OAI211_X1 U14357 ( .C1(n15500), .C2(n13597), .A(n11769), .B(n11768), .ZN(
        P2_U3203) );
  OAI21_X1 U14358 ( .B1(n11771), .B2(n11774), .A(n11770), .ZN(n15510) );
  INV_X1 U14359 ( .A(n11895), .ZN(n11772) );
  AOI21_X1 U14360 ( .B1(n11774), .B2(n11773), .A(n11772), .ZN(n11775) );
  AOI22_X1 U14361 ( .A1(n13602), .A2(n13647), .B1(n13617), .B2(n13649), .ZN(
        n11885) );
  OAI21_X1 U14362 ( .B1(n11775), .B2(n13896), .A(n11885), .ZN(n15505) );
  INV_X1 U14363 ( .A(n11776), .ZN(n11779) );
  INV_X1 U14364 ( .A(n11901), .ZN(n11778) );
  AOI211_X1 U14365 ( .C1(n15507), .C2(n11779), .A(n8410), .B(n11778), .ZN(
        n15506) );
  NAND2_X1 U14366 ( .A1(n15506), .A2(n13930), .ZN(n11782) );
  INV_X1 U14367 ( .A(n11780), .ZN(n11887) );
  AOI22_X1 U14368 ( .A1(n13926), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n11887), 
        .B2(n13931), .ZN(n11781) );
  OAI211_X1 U14369 ( .C1(n11890), .C2(n13824), .A(n11782), .B(n11781), .ZN(
        n11783) );
  AOI21_X1 U14370 ( .B1(n15505), .B2(n13919), .A(n11783), .ZN(n11784) );
  OAI21_X1 U14371 ( .B1(n13902), .B2(n15510), .A(n11784), .ZN(P2_U3255) );
  OAI21_X1 U14372 ( .B1(n11786), .B2(n12820), .A(n11785), .ZN(n11787) );
  INV_X1 U14373 ( .A(n11787), .ZN(n15661) );
  AOI21_X1 U14374 ( .B1(n11788), .B2(n12820), .A(n15685), .ZN(n11793) );
  OAI22_X1 U14375 ( .A1(n11790), .A2(n13276), .B1(n11789), .B2(n13278), .ZN(
        n11791) );
  AOI21_X1 U14376 ( .B1(n11793), .B2(n11792), .A(n11791), .ZN(n15660) );
  OAI21_X1 U14377 ( .B1(n15065), .B2(n15661), .A(n15660), .ZN(n11799) );
  INV_X1 U14378 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n11794) );
  OAI22_X1 U14379 ( .A1(n11797), .A2(n13424), .B1(n15741), .B2(n11794), .ZN(
        n11795) );
  AOI21_X1 U14380 ( .B1(n11799), .B2(n15741), .A(n11795), .ZN(n11796) );
  INV_X1 U14381 ( .A(n11796), .ZN(P3_U3408) );
  OAI22_X1 U14382 ( .A1(n13367), .A2(n11797), .B1(n15751), .B2(n8544), .ZN(
        n11798) );
  AOI21_X1 U14383 ( .B1(n11799), .B2(n15751), .A(n11798), .ZN(n11800) );
  INV_X1 U14384 ( .A(n11800), .ZN(P3_U3465) );
  NAND2_X1 U14385 ( .A1(n13112), .A2(P3_U3897), .ZN(n11801) );
  OAI21_X1 U14386 ( .B1(P3_U3897), .B2(n11802), .A(n11801), .ZN(P3_U3518) );
  XNOR2_X1 U14387 ( .A(n11803), .B(n14432), .ZN(n11804) );
  NAND2_X1 U14388 ( .A1(n14762), .A2(n14494), .ZN(n12418) );
  OAI21_X1 U14389 ( .B1(n11804), .B2(n15175), .A(n12418), .ZN(n15335) );
  INV_X1 U14390 ( .A(n15335), .ZN(n11814) );
  XNOR2_X1 U14391 ( .A(n11805), .B(n14432), .ZN(n15338) );
  NAND2_X1 U14392 ( .A1(n14275), .A2(n11916), .ZN(n11806) );
  NAND2_X1 U14393 ( .A1(n11806), .A2(n15122), .ZN(n11807) );
  OR2_X1 U14394 ( .A1(n11973), .A2(n11807), .ZN(n11809) );
  NAND2_X1 U14395 ( .A1(n15134), .A2(n14492), .ZN(n11808) );
  AND2_X1 U14396 ( .A1(n11809), .A2(n11808), .ZN(n15333) );
  AOI22_X1 U14397 ( .A1(n14765), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n7677), 
        .B2(n14929), .ZN(n11811) );
  NAND2_X1 U14398 ( .A1(n14275), .A2(n14717), .ZN(n11810) );
  OAI211_X1 U14399 ( .C1(n15333), .C2(n14958), .A(n11811), .B(n11810), .ZN(
        n11812) );
  AOI21_X1 U14400 ( .B1(n15338), .B2(n15126), .A(n11812), .ZN(n11813) );
  OAI21_X1 U14401 ( .B1(n11814), .B2(n14765), .A(n11813), .ZN(P1_U3283) );
  NAND2_X1 U14402 ( .A1(n11816), .A2(n11815), .ZN(n11821) );
  AND2_X1 U14403 ( .A1(n11818), .A2(n11817), .ZN(n11819) );
  OAI211_X1 U14404 ( .C1(n11821), .C2(n11820), .A(n11819), .B(n12788), .ZN(
        n11826) );
  AOI21_X1 U14405 ( .B1(n9897), .B2(n15657), .A(n11822), .ZN(n11823) );
  OAI21_X1 U14406 ( .B1(n7633), .B2(n12774), .A(n11823), .ZN(n11824) );
  AOI21_X1 U14407 ( .B1(n12770), .B2(n11947), .A(n11824), .ZN(n11825) );
  OAI211_X1 U14408 ( .C1(n15659), .C2(n12440), .A(n11826), .B(n11825), .ZN(
        P3_U3153) );
  NAND2_X1 U14409 ( .A1(n11827), .A2(n13433), .ZN(n11828) );
  OAI211_X1 U14410 ( .C1(n11829), .C2(n13440), .A(n11828), .B(n12992), .ZN(
        P3_U3272) );
  OAI211_X1 U14411 ( .C1(n11832), .C2(n11831), .A(n11830), .B(n12788), .ZN(
        n11838) );
  AOI21_X1 U14412 ( .B1(n9897), .B2(n11834), .A(n11833), .ZN(n11835) );
  OAI21_X1 U14413 ( .B1(n12103), .B2(n12774), .A(n11835), .ZN(n11836) );
  AOI21_X1 U14414 ( .B1(n12770), .B2(n12031), .A(n11836), .ZN(n11837) );
  OAI211_X1 U14415 ( .C1(n11839), .C2(n12440), .A(n11838), .B(n11837), .ZN(
        P3_U3161) );
  NOR2_X1 U14416 ( .A1(n11857), .A2(n11842), .ZN(n11843) );
  INV_X1 U14417 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n15552) );
  AOI22_X1 U14418 ( .A1(n13050), .A2(P3_REG2_REG_10__SCAN_IN), .B1(n8618), 
        .B2(n13011), .ZN(n11844) );
  AOI21_X1 U14419 ( .B1(n11845), .B2(n11844), .A(n12996), .ZN(n11870) );
  AOI22_X1 U14420 ( .A1(n13050), .A2(n8617), .B1(P3_REG1_REG_10__SCAN_IN), 
        .B2(n13011), .ZN(n11851) );
  NAND2_X1 U14421 ( .A1(P3_REG1_REG_8__SCAN_IN), .A2(n11853), .ZN(n11847) );
  NAND2_X1 U14422 ( .A1(n15557), .A2(n11848), .ZN(n11849) );
  NAND2_X1 U14423 ( .A1(P3_REG1_REG_9__SCAN_IN), .A2(n15562), .ZN(n15561) );
  OAI21_X1 U14424 ( .B1(n11851), .B2(n11850), .A(n13049), .ZN(n11868) );
  MUX2_X1 U14425 ( .A(n15552), .B(n8595), .S(n13027), .Z(n11858) );
  INV_X1 U14426 ( .A(n11858), .ZN(n11852) );
  NAND2_X1 U14427 ( .A1(n11852), .A2(n15557), .ZN(n15553) );
  OR2_X1 U14428 ( .A1(n11854), .A2(n11853), .ZN(n11856) );
  NAND2_X1 U14429 ( .A1(n11858), .A2(n11857), .ZN(n15554) );
  NAND2_X1 U14430 ( .A1(n11859), .A2(n15554), .ZN(n11861) );
  MUX2_X1 U14431 ( .A(P3_REG2_REG_10__SCAN_IN), .B(P3_REG1_REG_10__SCAN_IN), 
        .S(n13027), .Z(n13012) );
  XNOR2_X1 U14432 ( .A(n13012), .B(n13050), .ZN(n11860) );
  NAND2_X1 U14433 ( .A1(n11861), .A2(n11860), .ZN(n13010) );
  OAI21_X1 U14434 ( .B1(n11861), .B2(n11860), .A(n13010), .ZN(n11865) );
  NOR2_X1 U14435 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11862), .ZN(n12101) );
  INV_X1 U14436 ( .A(n15623), .ZN(n15548) );
  NOR2_X1 U14437 ( .A1(n15548), .A2(n11863), .ZN(n11864) );
  AOI211_X1 U14438 ( .C1(n15630), .C2(n11865), .A(n12101), .B(n11864), .ZN(
        n11866) );
  OAI21_X1 U14439 ( .B1(n13011), .B2(n15626), .A(n11866), .ZN(n11867) );
  AOI21_X1 U14440 ( .B1(n11868), .B2(n15628), .A(n11867), .ZN(n11869) );
  OAI21_X1 U14441 ( .B1(n11870), .B2(n15636), .A(n11869), .ZN(P3_U3192) );
  INV_X1 U14442 ( .A(n11871), .ZN(n11873) );
  NAND2_X1 U14443 ( .A1(n11873), .A2(n11872), .ZN(n11874) );
  XNOR2_X1 U14444 ( .A(n15507), .B(n13537), .ZN(n11876) );
  AND2_X1 U14445 ( .A1(n13648), .A2(n13912), .ZN(n11877) );
  NAND2_X1 U14446 ( .A1(n11876), .A2(n11877), .ZN(n12066) );
  INV_X1 U14447 ( .A(n11876), .ZN(n11879) );
  INV_X1 U14448 ( .A(n11877), .ZN(n11878) );
  NAND2_X1 U14449 ( .A1(n11879), .A2(n11878), .ZN(n11880) );
  NAND2_X1 U14450 ( .A1(n12066), .A2(n11880), .ZN(n11881) );
  AOI21_X1 U14451 ( .B1(n11882), .B2(n11881), .A(n13627), .ZN(n11883) );
  NAND2_X1 U14452 ( .A1(n11883), .A2(n12067), .ZN(n11889) );
  OAI22_X1 U14453 ( .A1(n13621), .A2(n11885), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11884), .ZN(n11886) );
  AOI21_X1 U14454 ( .B1(n11887), .B2(n13623), .A(n11886), .ZN(n11888) );
  OAI211_X1 U14455 ( .C1(n11890), .C2(n13597), .A(n11889), .B(n11888), .ZN(
        P2_U3189) );
  XNOR2_X1 U14456 ( .A(n11891), .B(n11892), .ZN(n15520) );
  INV_X1 U14457 ( .A(n11052), .ZN(n15514) );
  INV_X1 U14458 ( .A(n11892), .ZN(n11894) );
  NAND3_X1 U14459 ( .A1(n11895), .A2(n11894), .A3(n11893), .ZN(n11896) );
  NAND2_X1 U14460 ( .A1(n11897), .A2(n11896), .ZN(n11898) );
  NAND2_X1 U14461 ( .A1(n11898), .A2(n13906), .ZN(n11899) );
  AOI22_X1 U14462 ( .A1(n13602), .A2(n13646), .B1(n13617), .B2(n13648), .ZN(
        n12072) );
  NAND2_X1 U14463 ( .A1(n11899), .A2(n12072), .ZN(n11900) );
  AOI21_X1 U14464 ( .B1(n15520), .B2(n15514), .A(n11900), .ZN(n15522) );
  AOI21_X1 U14465 ( .B1(n12068), .B2(n11901), .A(n13912), .ZN(n11902) );
  NAND2_X1 U14466 ( .A1(n11902), .A2(n11958), .ZN(n15515) );
  INV_X1 U14467 ( .A(n11903), .ZN(n12074) );
  AOI22_X1 U14468 ( .A1(n13926), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n12074), 
        .B2(n13931), .ZN(n11905) );
  NAND2_X1 U14469 ( .A1(n12068), .A2(n13933), .ZN(n11904) );
  OAI211_X1 U14470 ( .C1(n15515), .C2(n13922), .A(n11905), .B(n11904), .ZN(
        n11906) );
  AOI21_X1 U14471 ( .B1(n15520), .B2(n13928), .A(n11906), .ZN(n11907) );
  OAI21_X1 U14472 ( .B1(n15522), .B2(n13926), .A(n11907), .ZN(P2_U3254) );
  INV_X1 U14473 ( .A(P3_DATAO_REG_29__SCAN_IN), .ZN(n11909) );
  NAND2_X1 U14474 ( .A1(n12673), .A2(P3_U3897), .ZN(n11908) );
  OAI21_X1 U14475 ( .B1(P3_U3897), .B2(n11909), .A(n11908), .ZN(P3_U3520) );
  XOR2_X1 U14476 ( .A(n11910), .B(n14431), .Z(n15325) );
  XNOR2_X1 U14477 ( .A(n11911), .B(n14431), .ZN(n11913) );
  OAI22_X1 U14478 ( .A1(n12354), .A2(n15131), .B1(n12492), .B2(n14947), .ZN(
        n11912) );
  AOI21_X1 U14479 ( .B1(n11913), .B2(n15160), .A(n11912), .ZN(n11914) );
  OAI21_X1 U14480 ( .B1(n15325), .B2(n14928), .A(n11914), .ZN(n15328) );
  NAND2_X1 U14481 ( .A1(n15328), .A2(n15143), .ZN(n11922) );
  INV_X1 U14482 ( .A(n14266), .ZN(n15327) );
  INV_X1 U14483 ( .A(n11915), .ZN(n11917) );
  OAI211_X1 U14484 ( .C1(n15327), .C2(n11917), .A(n15122), .B(n11916), .ZN(
        n15326) );
  INV_X1 U14485 ( .A(n15326), .ZN(n11920) );
  AOI22_X1 U14486 ( .A1(n14931), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n12351), 
        .B2(n14929), .ZN(n11918) );
  OAI21_X1 U14487 ( .B1(n15327), .B2(n15141), .A(n11918), .ZN(n11919) );
  AOI21_X1 U14488 ( .B1(n11920), .B2(n15125), .A(n11919), .ZN(n11921) );
  OAI211_X1 U14489 ( .C1(n15325), .C2(n14921), .A(n11922), .B(n11921), .ZN(
        P1_U3284) );
  NAND2_X1 U14490 ( .A1(n11923), .A2(P3_U3897), .ZN(n11924) );
  OAI21_X1 U14491 ( .B1(P3_U3897), .B2(n11925), .A(n11924), .ZN(P3_U3519) );
  NAND2_X1 U14492 ( .A1(n14250), .A2(n12635), .ZN(n11931) );
  NAND2_X1 U14493 ( .A1(n12621), .A2(n14497), .ZN(n11930) );
  NAND2_X1 U14494 ( .A1(n11931), .A2(n11930), .ZN(n11932) );
  XNOR2_X1 U14495 ( .A(n11932), .B(n12618), .ZN(n12120) );
  NOR2_X1 U14496 ( .A1(n12644), .A2(n11933), .ZN(n11934) );
  AOI21_X1 U14497 ( .B1(n14250), .B2(n12621), .A(n11934), .ZN(n12121) );
  XNOR2_X1 U14498 ( .A(n12120), .B(n12121), .ZN(n12122) );
  XNOR2_X1 U14499 ( .A(n11935), .B(n12122), .ZN(n11941) );
  AOI22_X1 U14500 ( .A1(n15109), .A2(n14498), .B1(n15107), .B2(n14496), .ZN(
        n11937) );
  OAI211_X1 U14501 ( .C1(n15303), .C2(n15111), .A(n11937), .B(n11936), .ZN(
        n11938) );
  AOI21_X1 U14502 ( .B1(n11939), .B2(n14205), .A(n11938), .ZN(n11940) );
  OAI21_X1 U14503 ( .B1(n11941), .B2(n15092), .A(n11940), .ZN(P1_U3239) );
  OAI21_X1 U14504 ( .B1(n11943), .B2(n12880), .A(n11942), .ZN(n11944) );
  INV_X1 U14505 ( .A(n11944), .ZN(n15654) );
  OAI211_X1 U14506 ( .C1(n11946), .C2(n12819), .A(n11945), .B(n15703), .ZN(
        n11949) );
  AOI22_X1 U14507 ( .A1(n15700), .A2(n11947), .B1(n12189), .B2(n15697), .ZN(
        n11948) );
  AND2_X1 U14508 ( .A1(n11949), .A2(n11948), .ZN(n15653) );
  OAI21_X1 U14509 ( .B1(n15654), .B2(n15065), .A(n15653), .ZN(n11955) );
  OAI22_X1 U14510 ( .A1(n13367), .A2(n11953), .B1(n15751), .B2(n8562), .ZN(
        n11950) );
  AOI21_X1 U14511 ( .B1(n11955), .B2(n15751), .A(n11950), .ZN(n11951) );
  INV_X1 U14512 ( .A(n11951), .ZN(P3_U3466) );
  INV_X1 U14513 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n11952) );
  OAI22_X1 U14514 ( .A1(n11953), .A2(n13424), .B1(n15741), .B2(n11952), .ZN(
        n11954) );
  AOI21_X1 U14515 ( .B1(n11955), .B2(n15741), .A(n11954), .ZN(n11956) );
  INV_X1 U14516 ( .A(n11956), .ZN(P3_U3411) );
  XNOR2_X1 U14517 ( .A(n11957), .B(n11963), .ZN(n14021) );
  AOI211_X1 U14518 ( .C1(n14019), .C2(n11958), .A(n8410), .B(n7173), .ZN(
        n14018) );
  INV_X1 U14519 ( .A(n14019), .ZN(n11959) );
  NOR2_X1 U14520 ( .A1(n11959), .A2(n13824), .ZN(n11962) );
  OAI22_X1 U14521 ( .A1(n13919), .A2(n11960), .B1(n12113), .B2(n13916), .ZN(
        n11961) );
  AOI211_X1 U14522 ( .C1(n14018), .C2(n13930), .A(n11962), .B(n11961), .ZN(
        n11967) );
  XNOR2_X1 U14523 ( .A(n11964), .B(n11963), .ZN(n11965) );
  AOI22_X1 U14524 ( .A1(n13602), .A2(n13645), .B1(n13617), .B2(n13647), .ZN(
        n12115) );
  OAI21_X1 U14525 ( .B1(n11965), .B2(n13896), .A(n12115), .ZN(n14017) );
  NAND2_X1 U14526 ( .A1(n14017), .A2(n13919), .ZN(n11966) );
  OAI211_X1 U14527 ( .C1(n14021), .C2(n13902), .A(n11967), .B(n11966), .ZN(
        P2_U3253) );
  XNOR2_X1 U14528 ( .A(n11968), .B(n14433), .ZN(n11969) );
  NAND2_X1 U14529 ( .A1(n11969), .A2(n15160), .ZN(n11971) );
  AOI22_X1 U14530 ( .A1(n15134), .A2(n15108), .B1(n14762), .B2(n14493), .ZN(
        n11970) );
  NAND2_X1 U14531 ( .A1(n11971), .A2(n11970), .ZN(n15184) );
  INV_X1 U14532 ( .A(n15184), .ZN(n11978) );
  XNOR2_X1 U14533 ( .A(n11972), .B(n14433), .ZN(n15179) );
  OAI211_X1 U14534 ( .C1(n15181), .C2(n11973), .A(n15122), .B(n14918), .ZN(
        n15180) );
  AOI22_X1 U14535 ( .A1(n14765), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n12494), 
        .B2(n14929), .ZN(n11975) );
  NAND2_X1 U14536 ( .A1(n14279), .A2(n14717), .ZN(n11974) );
  OAI211_X1 U14537 ( .C1(n15180), .C2(n14958), .A(n11975), .B(n11974), .ZN(
        n11976) );
  AOI21_X1 U14538 ( .B1(n15179), .B2(n15126), .A(n11976), .ZN(n11977) );
  OAI21_X1 U14539 ( .B1(n11978), .B2(n14765), .A(n11977), .ZN(P1_U3282) );
  INV_X1 U14540 ( .A(n13710), .ZN(n11981) );
  INV_X1 U14541 ( .A(n11979), .ZN(n11982) );
  OAI222_X1 U14542 ( .A1(P2_U3088), .A2(n11981), .B1(n14083), .B2(n11982), 
        .C1(n11980), .C2(n14072), .ZN(P2_U3309) );
  INV_X1 U14543 ( .A(n14611), .ZN(n15265) );
  OAI222_X1 U14544 ( .A1(n14891), .A2(n11983), .B1(n14885), .B2(n11982), .C1(
        n15265), .C2(P1_U3086), .ZN(P1_U3337) );
  INV_X1 U14545 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n11990) );
  NAND2_X1 U14546 ( .A1(n11984), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n11988) );
  INV_X1 U14547 ( .A(P3_REG2_REG_31__SCAN_IN), .ZN(n11985) );
  OR2_X1 U14548 ( .A1(n11986), .A2(n11985), .ZN(n11987) );
  OAI211_X1 U14549 ( .C1(n11990), .C2(n11989), .A(n11988), .B(n11987), .ZN(
        n11991) );
  INV_X1 U14550 ( .A(n11991), .ZN(n11992) );
  INV_X1 U14551 ( .A(n13069), .ZN(n12811) );
  NAND2_X1 U14552 ( .A1(n12811), .A2(P3_U3897), .ZN(n11994) );
  OAI21_X1 U14553 ( .B1(P3_U3897), .B2(n11995), .A(n11994), .ZN(P3_U3522) );
  NOR2_X1 U14554 ( .A1(n12004), .A2(n11996), .ZN(n11998) );
  NOR2_X1 U14555 ( .A1(n11998), .A2(n11997), .ZN(n12002) );
  INV_X1 U14556 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n12000) );
  NAND2_X1 U14557 ( .A1(n12008), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n12140) );
  INV_X1 U14558 ( .A(n12140), .ZN(n11999) );
  AOI21_X1 U14559 ( .B1(n12000), .B2(n12145), .A(n11999), .ZN(n12001) );
  NAND2_X1 U14560 ( .A1(n12001), .A2(n12002), .ZN(n12139) );
  OAI211_X1 U14561 ( .C1(n12002), .C2(n12001), .A(n15258), .B(n12139), .ZN(
        n12014) );
  NAND2_X1 U14562 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n14134)
         );
  NOR2_X1 U14563 ( .A1(n12004), .A2(n12003), .ZN(n12006) );
  NOR2_X1 U14564 ( .A1(n12006), .A2(n12005), .ZN(n12010) );
  NOR2_X1 U14565 ( .A1(n12008), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n12007) );
  AOI21_X1 U14566 ( .B1(n12008), .B2(P1_REG1_REG_16__SCAN_IN), .A(n12007), 
        .ZN(n12009) );
  NAND2_X1 U14567 ( .A1(n12009), .A2(n12010), .ZN(n12144) );
  OAI211_X1 U14568 ( .C1(n12010), .C2(n12009), .A(n15261), .B(n12144), .ZN(
        n12011) );
  NAND2_X1 U14569 ( .A1(n14134), .A2(n12011), .ZN(n12012) );
  AOI21_X1 U14570 ( .B1(n14593), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n12012), 
        .ZN(n12013) );
  OAI211_X1 U14571 ( .C1(n15266), .C2(n12145), .A(n12014), .B(n12013), .ZN(
        P1_U3259) );
  INV_X1 U14572 ( .A(n12015), .ZN(n12136) );
  OAI222_X1 U14573 ( .A1(n14891), .A2(n12016), .B1(n14885), .B2(n12136), .C1(
        n14387), .C2(P1_U3086), .ZN(P1_U3335) );
  OR2_X1 U14574 ( .A1(n15680), .A2(n12017), .ZN(n15652) );
  NAND2_X1 U14575 ( .A1(n15693), .A2(n15652), .ZN(n15054) );
  MUX2_X1 U14576 ( .A(n12019), .B(n12018), .S(n15714), .Z(n12023) );
  AOI22_X1 U14577 ( .A1(n15673), .A2(n12021), .B1(n15710), .B2(n12020), .ZN(
        n12022) );
  OAI211_X1 U14578 ( .C1(n12024), .C2(n15054), .A(n12023), .B(n12022), .ZN(
        P3_U3230) );
  INV_X1 U14579 ( .A(n12025), .ZN(n12027) );
  OAI222_X1 U14580 ( .A1(n14891), .A2(n12026), .B1(n14885), .B2(n12027), .C1(
        P1_U3086), .C2(n14619), .ZN(P1_U3336) );
  OAI222_X1 U14581 ( .A1(n14072), .A2(n12028), .B1(n14083), .B2(n12027), .C1(
        n13718), .C2(P2_U3088), .ZN(P2_U3308) );
  XNOR2_X1 U14582 ( .A(n12030), .B(n12029), .ZN(n12037) );
  AOI22_X1 U14583 ( .A1(n15700), .A2(n12031), .B1(n15639), .B2(n15697), .ZN(
        n12036) );
  OR2_X1 U14584 ( .A1(n12032), .A2(n12886), .ZN(n12033) );
  NAND2_X1 U14585 ( .A1(n12034), .A2(n12033), .ZN(n15728) );
  NAND2_X1 U14586 ( .A1(n15728), .A2(n15680), .ZN(n12035) );
  OAI211_X1 U14587 ( .C1(n12037), .C2(n15685), .A(n12036), .B(n12035), .ZN(
        n15726) );
  INV_X1 U14588 ( .A(n15726), .ZN(n12044) );
  NOR2_X1 U14589 ( .A1(n12038), .A2(n15730), .ZN(n15727) );
  AOI22_X1 U14590 ( .A1(n15648), .A2(n15727), .B1(n15710), .B2(n12039), .ZN(
        n12040) );
  OAI21_X1 U14591 ( .B1(n12041), .B2(n15693), .A(n12040), .ZN(n12042) );
  AOI21_X1 U14592 ( .B1(n15728), .B2(n15711), .A(n12042), .ZN(n12043) );
  OAI21_X1 U14593 ( .B1(n12044), .B2(n13303), .A(n12043), .ZN(P3_U3225) );
  OR2_X1 U14594 ( .A1(n12046), .A2(n12047), .ZN(n12098) );
  INV_X1 U14595 ( .A(n12098), .ZN(n12045) );
  AOI21_X1 U14596 ( .B1(n12047), .B2(n12046), .A(n12045), .ZN(n12053) );
  INV_X1 U14597 ( .A(n12193), .ZN(n12051) );
  NOR2_X1 U14598 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n8596), .ZN(n15560) );
  AOI21_X1 U14599 ( .B1(n12794), .B2(n15043), .A(n15560), .ZN(n12049) );
  NAND2_X1 U14600 ( .A1(n9897), .A2(n12195), .ZN(n12048) );
  OAI211_X1 U14601 ( .C1(n12792), .C2(n7633), .A(n12049), .B(n12048), .ZN(
        n12050) );
  AOI21_X1 U14602 ( .B1(n12051), .B2(n12790), .A(n12050), .ZN(n12052) );
  OAI21_X1 U14603 ( .B1(n12053), .B2(n12777), .A(n12052), .ZN(P3_U3171) );
  XNOR2_X1 U14604 ( .A(n12054), .B(n12055), .ZN(n15084) );
  INV_X1 U14605 ( .A(n15084), .ZN(n12062) );
  XNOR2_X1 U14606 ( .A(n12056), .B(n12055), .ZN(n12057) );
  AOI22_X1 U14607 ( .A1(n13602), .A2(n13644), .B1(n13617), .B2(n13646), .ZN(
        n12087) );
  OAI21_X1 U14608 ( .B1(n12057), .B2(n13896), .A(n12087), .ZN(n15082) );
  OAI211_X1 U14609 ( .C1(n7172), .C2(n7173), .A(n11777), .B(n12204), .ZN(
        n15081) );
  AOI22_X1 U14610 ( .A1(n13926), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n12089), 
        .B2(n13931), .ZN(n12059) );
  NAND2_X1 U14611 ( .A1(n12090), .A2(n13933), .ZN(n12058) );
  OAI211_X1 U14612 ( .C1(n15081), .C2(n13922), .A(n12059), .B(n12058), .ZN(
        n12060) );
  AOI21_X1 U14613 ( .B1(n15082), .B2(n13919), .A(n12060), .ZN(n12061) );
  OAI21_X1 U14614 ( .B1(n12062), .B2(n13902), .A(n12061), .ZN(P2_U3252) );
  OAI222_X1 U14615 ( .A1(P3_U3151), .A2(n12065), .B1(n13440), .B2(n12064), 
        .C1(n12666), .C2(n12063), .ZN(P3_U3271) );
  INV_X1 U14616 ( .A(n12068), .ZN(n15517) );
  XNOR2_X1 U14617 ( .A(n12068), .B(n13485), .ZN(n12078) );
  AND2_X1 U14618 ( .A1(n13647), .A2(n13912), .ZN(n12077) );
  INV_X1 U14619 ( .A(n12077), .ZN(n12079) );
  XNOR2_X1 U14620 ( .A(n12078), .B(n12079), .ZN(n12069) );
  NAND2_X1 U14621 ( .A1(n6794), .A2(n12069), .ZN(n12108) );
  OAI21_X1 U14622 ( .B1(n6794), .B2(n12069), .A(n12108), .ZN(n12070) );
  NAND2_X1 U14623 ( .A1(n12070), .A2(n13591), .ZN(n12076) );
  OAI21_X1 U14624 ( .B1(n13621), .B2(n12072), .A(n12071), .ZN(n12073) );
  AOI21_X1 U14625 ( .B1(n12074), .B2(n13623), .A(n12073), .ZN(n12075) );
  OAI211_X1 U14626 ( .C1(n15517), .C2(n13597), .A(n12076), .B(n12075), .ZN(
        P2_U3208) );
  AND2_X1 U14627 ( .A1(n12078), .A2(n12077), .ZN(n12081) );
  XNOR2_X1 U14628 ( .A(n14019), .B(n13498), .ZN(n12082) );
  NAND2_X1 U14629 ( .A1(n13646), .A2(n13912), .ZN(n12083) );
  NAND2_X1 U14630 ( .A1(n12082), .A2(n12083), .ZN(n12110) );
  INV_X1 U14631 ( .A(n12078), .ZN(n12080) );
  NAND2_X1 U14632 ( .A1(n12080), .A2(n12079), .ZN(n12107) );
  INV_X1 U14633 ( .A(n12082), .ZN(n12085) );
  INV_X1 U14634 ( .A(n12083), .ZN(n12084) );
  NAND2_X1 U14635 ( .A1(n12085), .A2(n12084), .ZN(n12109) );
  XNOR2_X1 U14636 ( .A(n12090), .B(n13537), .ZN(n12244) );
  NAND2_X1 U14637 ( .A1(n13645), .A2(n8410), .ZN(n12242) );
  XNOR2_X1 U14638 ( .A(n12244), .B(n12242), .ZN(n12240) );
  XNOR2_X1 U14639 ( .A(n12241), .B(n12240), .ZN(n12093) );
  AND2_X1 U14640 ( .A1(P2_U3088), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n15403) );
  NOR2_X1 U14641 ( .A1(n13621), .A2(n12087), .ZN(n12088) );
  AOI211_X1 U14642 ( .C1(n13623), .C2(n12089), .A(n15403), .B(n12088), .ZN(
        n12092) );
  NAND2_X1 U14643 ( .A1(n12090), .A2(n13624), .ZN(n12091) );
  OAI211_X1 U14644 ( .C1(n12093), .C2(n13627), .A(n12092), .B(n12091), .ZN(
        P2_U3206) );
  NAND2_X1 U14645 ( .A1(n12098), .A2(n12094), .ZN(n12096) );
  AOI21_X1 U14646 ( .B1(n12096), .B2(n12095), .A(n12777), .ZN(n12100) );
  NAND2_X1 U14647 ( .A1(n12098), .A2(n12097), .ZN(n12099) );
  NAND2_X1 U14648 ( .A1(n12100), .A2(n12099), .ZN(n12106) );
  AOI21_X1 U14649 ( .B1(n12794), .B2(n15640), .A(n12101), .ZN(n12102) );
  OAI21_X1 U14650 ( .B1(n12792), .B2(n12103), .A(n12102), .ZN(n12104) );
  AOI21_X1 U14651 ( .B1(n15642), .B2(n12790), .A(n12104), .ZN(n12105) );
  OAI211_X1 U14652 ( .C1(n12797), .C2(n15647), .A(n12106), .B(n12105), .ZN(
        P3_U3157) );
  NAND2_X1 U14653 ( .A1(n12108), .A2(n12107), .ZN(n12112) );
  NAND2_X1 U14654 ( .A1(n12110), .A2(n12109), .ZN(n12111) );
  XNOR2_X1 U14655 ( .A(n12112), .B(n12111), .ZN(n12119) );
  NOR2_X1 U14656 ( .A1(n13607), .A2(n12113), .ZN(n12117) );
  OAI21_X1 U14657 ( .B1(n13621), .B2(n12115), .A(n12114), .ZN(n12116) );
  AOI211_X1 U14658 ( .C1(n14019), .C2(n13624), .A(n12117), .B(n12116), .ZN(
        n12118) );
  OAI21_X1 U14659 ( .B1(n12119), .B2(n13627), .A(n12118), .ZN(P2_U3196) );
  OAI22_X2 U14660 ( .A1(n12123), .A2(n12122), .B1(n12121), .B2(n12120), .ZN(
        n12160) );
  NOR2_X1 U14661 ( .A1(n12644), .A2(n12124), .ZN(n12125) );
  AOI21_X1 U14662 ( .B1(n15309), .B2(n12621), .A(n12125), .ZN(n12156) );
  AOI22_X1 U14663 ( .A1(n15309), .A2(n12635), .B1(n12621), .B2(n14496), .ZN(
        n12126) );
  XNOR2_X1 U14664 ( .A(n12126), .B(n12646), .ZN(n12155) );
  XOR2_X1 U14665 ( .A(n12156), .B(n12155), .Z(n12159) );
  XOR2_X1 U14666 ( .A(n12160), .B(n12159), .Z(n12134) );
  NOR2_X1 U14667 ( .A1(n12127), .A2(n15111), .ZN(n12133) );
  NAND2_X1 U14668 ( .A1(n14195), .A2(n12128), .ZN(n12129) );
  OAI211_X1 U14669 ( .C1(n15119), .C2(n12131), .A(n12130), .B(n12129), .ZN(
        n12132) );
  AOI211_X1 U14670 ( .C1(n12134), .C2(n15114), .A(n12133), .B(n12132), .ZN(
        n12135) );
  INV_X1 U14671 ( .A(n12135), .ZN(P1_U3213) );
  OAI222_X1 U14672 ( .A1(n14072), .A2(n12138), .B1(P2_U3088), .B2(n12137), 
        .C1(n14075), .C2(n12136), .ZN(P2_U3307) );
  NAND2_X1 U14673 ( .A1(n12140), .A2(n12139), .ZN(n12143) );
  NAND2_X1 U14674 ( .A1(n14605), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n14610) );
  INV_X1 U14675 ( .A(n14610), .ZN(n12141) );
  AOI21_X1 U14676 ( .B1(n12446), .B2(n12152), .A(n12141), .ZN(n12142) );
  NAND2_X1 U14677 ( .A1(n12142), .A2(n12143), .ZN(n14609) );
  OAI211_X1 U14678 ( .C1(n12143), .C2(n12142), .A(n15258), .B(n14609), .ZN(
        n12151) );
  NAND2_X1 U14679 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n14144)
         );
  XNOR2_X1 U14680 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n12152), .ZN(n12147) );
  INV_X1 U14681 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n15152) );
  OAI21_X1 U14682 ( .B1(n15152), .B2(n12145), .A(n12144), .ZN(n12146) );
  NAND2_X1 U14683 ( .A1(n12147), .A2(n12146), .ZN(n14603) );
  OAI211_X1 U14684 ( .C1(n12147), .C2(n12146), .A(n14603), .B(n15261), .ZN(
        n12148) );
  NAND2_X1 U14685 ( .A1(n14144), .A2(n12148), .ZN(n12149) );
  AOI21_X1 U14686 ( .B1(n14593), .B2(P1_ADDR_REG_17__SCAN_IN), .A(n12149), 
        .ZN(n12150) );
  OAI211_X1 U14687 ( .C1(n15266), .C2(n12152), .A(n12151), .B(n12150), .ZN(
        P1_U3260) );
  INV_X1 U14688 ( .A(n12153), .ZN(n12659) );
  OAI222_X1 U14689 ( .A1(n14891), .A2(n12154), .B1(n14885), .B2(n12659), .C1(
        P1_U3086), .C2(n14381), .ZN(P1_U3334) );
  INV_X1 U14690 ( .A(n12155), .ZN(n12158) );
  INV_X1 U14691 ( .A(n12156), .ZN(n12157) );
  AOI21_X2 U14692 ( .B1(n12160), .B2(n12159), .A(n7684), .ZN(n12169) );
  NAND2_X1 U14693 ( .A1(n14262), .A2(n12635), .ZN(n12162) );
  NAND2_X1 U14694 ( .A1(n12621), .A2(n14495), .ZN(n12161) );
  NAND2_X1 U14695 ( .A1(n12162), .A2(n12161), .ZN(n12163) );
  XNOR2_X1 U14696 ( .A(n12163), .B(n12646), .ZN(n12167) );
  NAND2_X1 U14697 ( .A1(n14262), .A2(n12621), .ZN(n12165) );
  NAND2_X1 U14698 ( .A1(n10728), .A2(n14495), .ZN(n12164) );
  NAND2_X1 U14699 ( .A1(n12165), .A2(n12164), .ZN(n12166) );
  NOR2_X1 U14700 ( .A1(n12167), .A2(n12166), .ZN(n12345) );
  AOI21_X1 U14701 ( .B1(n12167), .B2(n12166), .A(n12345), .ZN(n12168) );
  OAI21_X1 U14702 ( .B1(n6851), .B2(n12168), .A(n12347), .ZN(n12170) );
  NAND2_X1 U14703 ( .A1(n12170), .A2(n15114), .ZN(n12175) );
  INV_X1 U14704 ( .A(n14195), .ZN(n14203) );
  NAND2_X1 U14705 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n14573) );
  OAI21_X1 U14706 ( .B1(n14203), .B2(n12171), .A(n14573), .ZN(n12172) );
  AOI21_X1 U14707 ( .B1(n12173), .B2(n14205), .A(n12172), .ZN(n12174) );
  OAI211_X1 U14708 ( .C1(n15320), .C2(n15111), .A(n12175), .B(n12174), .ZN(
        P1_U3221) );
  NAND2_X1 U14709 ( .A1(n6967), .A2(n12177), .ZN(n12178) );
  XNOR2_X1 U14710 ( .A(n12178), .B(n12372), .ZN(n12186) );
  NOR2_X1 U14711 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12179), .ZN(n15571) );
  NOR2_X1 U14712 ( .A1(n12774), .A2(n12180), .ZN(n12181) );
  AOI211_X1 U14713 ( .C1(n12770), .C2(n15043), .A(n15571), .B(n12181), .ZN(
        n12182) );
  OAI21_X1 U14714 ( .B1(n15046), .B2(n12440), .A(n12182), .ZN(n12183) );
  AOI21_X1 U14715 ( .B1(n12184), .B2(n9897), .A(n12183), .ZN(n12185) );
  OAI21_X1 U14716 ( .B1(n12186), .B2(n12777), .A(n12185), .ZN(P3_U3176) );
  XOR2_X1 U14717 ( .A(n12891), .B(n12187), .Z(n15735) );
  INV_X1 U14718 ( .A(n15735), .ZN(n12198) );
  INV_X1 U14719 ( .A(n15711), .ZN(n13121) );
  XNOR2_X1 U14720 ( .A(n12188), .B(n12891), .ZN(n12192) );
  NAND2_X1 U14721 ( .A1(n15735), .A2(n15680), .ZN(n12191) );
  AOI22_X1 U14722 ( .A1(n15700), .A2(n12189), .B1(n15043), .B2(n15697), .ZN(
        n12190) );
  OAI211_X1 U14723 ( .C1(n15685), .C2(n12192), .A(n12191), .B(n12190), .ZN(
        n15732) );
  NAND2_X1 U14724 ( .A1(n15732), .A2(n15693), .ZN(n12197) );
  OAI22_X1 U14725 ( .A1(n15693), .A2(n15552), .B1(n12193), .B2(n15675), .ZN(
        n12194) );
  AOI21_X1 U14726 ( .B1(n15673), .B2(n12195), .A(n12194), .ZN(n12196) );
  OAI211_X1 U14727 ( .C1(n12198), .C2(n13121), .A(n12197), .B(n12196), .ZN(
        P3_U3224) );
  XNOR2_X1 U14728 ( .A(n12199), .B(n12209), .ZN(n12202) );
  NAND2_X1 U14729 ( .A1(n13643), .A2(n13602), .ZN(n12201) );
  NAND2_X1 U14730 ( .A1(n13617), .A2(n13645), .ZN(n12200) );
  AND2_X1 U14731 ( .A1(n12201), .A2(n12200), .ZN(n12252) );
  OAI21_X1 U14732 ( .B1(n12202), .B2(n13896), .A(n12252), .ZN(n12274) );
  INV_X1 U14733 ( .A(n12274), .ZN(n12213) );
  INV_X1 U14734 ( .A(n12263), .ZN(n12203) );
  AOI211_X1 U14735 ( .C1(n12277), .C2(n12204), .A(n8410), .B(n12203), .ZN(
        n12273) );
  NOR2_X1 U14736 ( .A1(n12205), .A2(n13824), .ZN(n12208) );
  OAI22_X1 U14737 ( .A1(n13919), .A2(n12206), .B1(n12250), .B2(n13916), .ZN(
        n12207) );
  AOI211_X1 U14738 ( .C1(n12273), .C2(n13930), .A(n12208), .B(n12207), .ZN(
        n12212) );
  XNOR2_X1 U14739 ( .A(n12210), .B(n12209), .ZN(n12275) );
  NAND2_X1 U14740 ( .A1(n12275), .A2(n13924), .ZN(n12211) );
  OAI211_X1 U14741 ( .C1(n13926), .C2(n12213), .A(n12212), .B(n12211), .ZN(
        P2_U3251) );
  INV_X1 U14742 ( .A(n12214), .ZN(n12215) );
  OAI222_X1 U14743 ( .A1(P3_U3151), .A2(n12217), .B1(n13440), .B2(n12216), 
        .C1(n12666), .C2(n12215), .ZN(P3_U3270) );
  XOR2_X1 U14744 ( .A(n12219), .B(n12218), .Z(n12225) );
  NOR2_X1 U14745 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12220), .ZN(n15588) );
  NOR2_X1 U14746 ( .A1(n12774), .A2(n12373), .ZN(n12221) );
  AOI211_X1 U14747 ( .C1(n12770), .C2(n15640), .A(n15588), .B(n12221), .ZN(
        n12222) );
  OAI21_X1 U14748 ( .B1(n12374), .B2(n12440), .A(n12222), .ZN(n12223) );
  AOI21_X1 U14749 ( .B1(n9897), .B2(n15069), .A(n12223), .ZN(n12224) );
  OAI21_X1 U14750 ( .B1(n12225), .B2(n12777), .A(n12224), .ZN(P3_U3164) );
  XNOR2_X1 U14751 ( .A(n12226), .B(n14298), .ZN(n12228) );
  OAI22_X1 U14752 ( .A1(n15132), .A2(n14947), .B1(n15087), .B2(n15131), .ZN(
        n12227) );
  AOI21_X1 U14753 ( .B1(n12228), .B2(n15160), .A(n12227), .ZN(n15169) );
  OAI22_X1 U14754 ( .A1(n15143), .A2(n11252), .B1(n15100), .B2(n15136), .ZN(
        n12231) );
  AOI21_X1 U14755 ( .B1(n15164), .B2(n14956), .A(n14741), .ZN(n12229) );
  NAND2_X1 U14756 ( .A1(n12229), .A2(n12316), .ZN(n15166) );
  NOR2_X1 U14757 ( .A1(n15166), .A2(n14958), .ZN(n12230) );
  AOI211_X1 U14758 ( .C1(n14717), .C2(n15164), .A(n12231), .B(n12230), .ZN(
        n12234) );
  NAND2_X1 U14759 ( .A1(n12232), .A2(n14438), .ZN(n15162) );
  NAND3_X1 U14760 ( .A1(n15163), .A2(n15162), .A3(n15126), .ZN(n12233) );
  OAI211_X1 U14761 ( .C1(n15169), .C2(n14765), .A(n12234), .B(n12233), .ZN(
        P1_U3279) );
  XNOR2_X1 U14762 ( .A(n12277), .B(n13498), .ZN(n12235) );
  NAND2_X1 U14763 ( .A1(n13644), .A2(n13912), .ZN(n12236) );
  NAND2_X1 U14764 ( .A1(n12235), .A2(n12236), .ZN(n12304) );
  INV_X1 U14765 ( .A(n12235), .ZN(n12238) );
  INV_X1 U14766 ( .A(n12236), .ZN(n12237) );
  NAND2_X1 U14767 ( .A1(n12238), .A2(n12237), .ZN(n12239) );
  NAND2_X1 U14768 ( .A1(n12304), .A2(n12239), .ZN(n12249) );
  INV_X1 U14769 ( .A(n12242), .ZN(n12243) );
  NAND2_X1 U14770 ( .A1(n12244), .A2(n12243), .ZN(n12245) );
  INV_X1 U14771 ( .A(n12305), .ZN(n12247) );
  AOI21_X1 U14772 ( .B1(n12249), .B2(n12248), .A(n12247), .ZN(n12256) );
  NOR2_X1 U14773 ( .A1(n13607), .A2(n12250), .ZN(n12254) );
  OAI22_X1 U14774 ( .A1(n13621), .A2(n12252), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12251), .ZN(n12253) );
  AOI211_X1 U14775 ( .C1(n12277), .C2(n13624), .A(n12254), .B(n12253), .ZN(
        n12255) );
  OAI21_X1 U14776 ( .B1(n12256), .B2(n13627), .A(n12255), .ZN(P2_U3187) );
  XNOR2_X1 U14777 ( .A(n12258), .B(n12257), .ZN(n12262) );
  NAND2_X1 U14778 ( .A1(n13642), .A2(n13602), .ZN(n12260) );
  NAND2_X1 U14779 ( .A1(n13617), .A2(n13644), .ZN(n12259) );
  NAND2_X1 U14780 ( .A1(n12260), .A2(n12259), .ZN(n12306) );
  INV_X1 U14781 ( .A(n12306), .ZN(n12261) );
  OAI21_X1 U14782 ( .B1(n12262), .B2(n13896), .A(n12261), .ZN(n12292) );
  INV_X1 U14783 ( .A(n12292), .ZN(n12272) );
  AOI211_X1 U14784 ( .C1(n12310), .C2(n12263), .A(n8410), .B(n12392), .ZN(
        n12293) );
  INV_X1 U14785 ( .A(n12310), .ZN(n12264) );
  NOR2_X1 U14786 ( .A1(n12264), .A2(n13824), .ZN(n12267) );
  OAI22_X1 U14787 ( .A1(n13919), .A2(n12265), .B1(n12308), .B2(n13916), .ZN(
        n12266) );
  AOI211_X1 U14788 ( .C1(n12293), .C2(n13930), .A(n12267), .B(n12266), .ZN(
        n12271) );
  XNOR2_X1 U14789 ( .A(n12269), .B(n12268), .ZN(n12294) );
  NAND2_X1 U14790 ( .A1(n12294), .A2(n13924), .ZN(n12270) );
  OAI211_X1 U14791 ( .C1(n13926), .C2(n12272), .A(n12271), .B(n12270), .ZN(
        P2_U3250) );
  AOI211_X1 U14792 ( .C1(n15491), .C2(n12275), .A(n12274), .B(n12273), .ZN(
        n12279) );
  AOI22_X1 U14793 ( .A1(n12277), .A2(n14002), .B1(P2_REG1_REG_14__SCAN_IN), 
        .B2(n15536), .ZN(n12276) );
  OAI21_X1 U14794 ( .B1(n12279), .B2(n15536), .A(n12276), .ZN(P2_U3513) );
  AOI22_X1 U14795 ( .A1(n12277), .A2(n8423), .B1(P2_REG0_REG_14__SCAN_IN), 
        .B2(n15523), .ZN(n12278) );
  OAI21_X1 U14796 ( .B1(n12279), .B2(n15523), .A(n12278), .ZN(P2_U3472) );
  XNOR2_X1 U14797 ( .A(n12280), .B(n13292), .ZN(n12281) );
  XNOR2_X1 U14798 ( .A(n12282), .B(n12281), .ZN(n12287) );
  NOR2_X1 U14799 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n8684), .ZN(n15603) );
  NOR2_X1 U14800 ( .A1(n12774), .A2(n13275), .ZN(n12283) );
  AOI211_X1 U14801 ( .C1(n12770), .C2(n15042), .A(n15603), .B(n12283), .ZN(
        n12284) );
  OAI21_X1 U14802 ( .B1(n12365), .B2(n12440), .A(n12284), .ZN(n12285) );
  AOI21_X1 U14803 ( .B1(n12364), .B2(n9897), .A(n12285), .ZN(n12286) );
  OAI21_X1 U14804 ( .B1(n12287), .B2(n12777), .A(n12286), .ZN(P3_U3174) );
  INV_X1 U14805 ( .A(n12288), .ZN(n12289) );
  OAI222_X1 U14806 ( .A1(P3_U3151), .A2(n12291), .B1(n13440), .B2(n12290), 
        .C1(n12666), .C2(n12289), .ZN(P3_U3269) );
  AOI211_X1 U14807 ( .C1(n15491), .C2(n12294), .A(n12293), .B(n12292), .ZN(
        n12297) );
  AOI22_X1 U14808 ( .A1(n12310), .A2(n8423), .B1(P2_REG0_REG_15__SCAN_IN), 
        .B2(n15523), .ZN(n12295) );
  OAI21_X1 U14809 ( .B1(n12297), .B2(n15523), .A(n12295), .ZN(P2_U3475) );
  AOI22_X1 U14810 ( .A1(n12310), .A2(n14002), .B1(P2_REG1_REG_15__SCAN_IN), 
        .B2(n15536), .ZN(n12296) );
  OAI21_X1 U14811 ( .B1(n12297), .B2(n15536), .A(n12296), .ZN(P2_U3514) );
  INV_X1 U14812 ( .A(n12301), .ZN(n12300) );
  NAND2_X1 U14813 ( .A1(n14080), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n12299) );
  OAI211_X1 U14814 ( .C1(n12300), .C2(n14083), .A(n12299), .B(n12298), .ZN(
        P2_U3304) );
  NAND2_X1 U14815 ( .A1(n12301), .A2(n14874), .ZN(n12302) );
  OAI211_X1 U14816 ( .C1(n12303), .C2(n14869), .A(n12302), .B(n14475), .ZN(
        P1_U3332) );
  XNOR2_X1 U14817 ( .A(n12310), .B(n13485), .ZN(n12463) );
  AND2_X1 U14818 ( .A1(n13643), .A2(n13912), .ZN(n12461) );
  XNOR2_X1 U14819 ( .A(n12462), .B(n12461), .ZN(n12312) );
  AND2_X1 U14820 ( .A1(P2_U3088), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n15425) );
  AOI21_X1 U14821 ( .B1(n13605), .B2(n12306), .A(n15425), .ZN(n12307) );
  OAI21_X1 U14822 ( .B1(n12308), .B2(n13607), .A(n12307), .ZN(n12309) );
  AOI21_X1 U14823 ( .B1(n12310), .B2(n13624), .A(n12309), .ZN(n12311) );
  OAI21_X1 U14824 ( .B1(n12312), .B2(n13627), .A(n12311), .ZN(P2_U3213) );
  INV_X1 U14825 ( .A(n12313), .ZN(n12314) );
  AOI21_X1 U14826 ( .B1(n14437), .B2(n12315), .A(n12314), .ZN(n15156) );
  NAND2_X1 U14827 ( .A1(n12552), .A2(n12316), .ZN(n12317) );
  NAND3_X1 U14828 ( .A1(n15121), .A2(n15122), .A3(n12317), .ZN(n15154) );
  INV_X1 U14829 ( .A(n15154), .ZN(n12321) );
  AOI22_X1 U14830 ( .A1(n14489), .A2(n15134), .B1(n15106), .B2(n14762), .ZN(
        n15153) );
  OAI22_X1 U14831 ( .A1(n14931), .A2(n15153), .B1(n14201), .B2(n15136), .ZN(
        n12318) );
  AOI21_X1 U14832 ( .B1(P1_REG2_REG_15__SCAN_IN), .B2(n14765), .A(n12318), 
        .ZN(n12319) );
  OAI21_X1 U14833 ( .B1(n7512), .B2(n15141), .A(n12319), .ZN(n12320) );
  AOI21_X1 U14834 ( .B1(n12321), .B2(n15125), .A(n12320), .ZN(n12324) );
  XOR2_X1 U14835 ( .A(n14437), .B(n12322), .Z(n15159) );
  INV_X1 U14836 ( .A(n14959), .ZN(n14721) );
  NAND2_X1 U14837 ( .A1(n15159), .A2(n14721), .ZN(n12323) );
  OAI211_X1 U14838 ( .C1(n15156), .C2(n14750), .A(n12324), .B(n12323), .ZN(
        P1_U3278) );
  INV_X1 U14839 ( .A(n12325), .ZN(n12330) );
  OAI222_X1 U14840 ( .A1(n14072), .A2(n12327), .B1(n14075), .B2(n12330), .C1(
        n12326), .C2(P2_U3088), .ZN(P2_U3303) );
  INV_X1 U14841 ( .A(n12328), .ZN(n12329) );
  OAI222_X1 U14842 ( .A1(n14891), .A2(n7281), .B1(n14885), .B2(n12330), .C1(
        P1_U3086), .C2(n12329), .ZN(P1_U3331) );
  XNOR2_X1 U14843 ( .A(n12332), .B(n12331), .ZN(n12339) );
  INV_X1 U14844 ( .A(n13423), .ZN(n12337) );
  NOR2_X1 U14845 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12333), .ZN(n15622) );
  NOR2_X1 U14846 ( .A1(n12774), .A2(n13262), .ZN(n12334) );
  AOI211_X1 U14847 ( .C1(n12770), .C2(n13292), .A(n15622), .B(n12334), .ZN(
        n12335) );
  OAI21_X1 U14848 ( .B1(n13298), .B2(n12440), .A(n12335), .ZN(n12336) );
  AOI21_X1 U14849 ( .B1(n12337), .B2(n9897), .A(n12336), .ZN(n12338) );
  OAI21_X1 U14850 ( .B1(n12339), .B2(n12777), .A(n12338), .ZN(P3_U3155) );
  INV_X1 U14851 ( .A(n12340), .ZN(n12342) );
  OAI222_X1 U14852 ( .A1(P3_U3151), .A2(n13027), .B1(n12666), .B2(n12342), 
        .C1(n12341), .C2(n13440), .ZN(P3_U3268) );
  AOI22_X1 U14853 ( .A1(n14266), .A2(n12635), .B1(n12621), .B2(n14494), .ZN(
        n12344) );
  XOR2_X1 U14854 ( .A(n12646), .B(n12344), .Z(n12350) );
  AOI22_X1 U14855 ( .A1(n14266), .A2(n12621), .B1(n10728), .B2(n14494), .ZN(
        n12348) );
  INV_X1 U14856 ( .A(n12345), .ZN(n12346) );
  INV_X1 U14857 ( .A(n12411), .ZN(n12409) );
  AOI21_X1 U14858 ( .B1(n12350), .B2(n12349), .A(n12409), .ZN(n12357) );
  AND2_X1 U14859 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n14592) );
  AOI21_X1 U14860 ( .B1(n15107), .B2(n14493), .A(n14592), .ZN(n12353) );
  NAND2_X1 U14861 ( .A1(n14205), .A2(n12351), .ZN(n12352) );
  OAI211_X1 U14862 ( .C1(n12354), .C2(n15086), .A(n12353), .B(n12352), .ZN(
        n12355) );
  AOI21_X1 U14863 ( .B1(n14266), .B2(n15097), .A(n12355), .ZN(n12356) );
  OAI21_X1 U14864 ( .B1(n12357), .B2(n15092), .A(n12356), .ZN(P1_U3231) );
  OAI211_X1 U14865 ( .C1(n12359), .C2(n12362), .A(n12358), .B(n15703), .ZN(
        n12361) );
  AOI22_X1 U14866 ( .A1(n15700), .A2(n15042), .B1(n12438), .B2(n15697), .ZN(
        n12360) );
  AND2_X1 U14867 ( .A1(n12361), .A2(n12360), .ZN(n15060) );
  XNOR2_X1 U14868 ( .A(n12363), .B(n7622), .ZN(n15063) );
  NAND2_X1 U14869 ( .A1(n12364), .A2(n15070), .ZN(n15059) );
  NOR2_X1 U14870 ( .A1(n15059), .A2(n15053), .ZN(n12367) );
  OAI22_X1 U14871 ( .A1(n15693), .A2(n8683), .B1(n12365), .B2(n15675), .ZN(
        n12366) );
  AOI211_X1 U14872 ( .C1(n15063), .C2(n15649), .A(n12367), .B(n12366), .ZN(
        n12368) );
  OAI21_X1 U14873 ( .B1(n15060), .B2(n13303), .A(n12368), .ZN(P3_U3220) );
  XOR2_X1 U14874 ( .A(n12369), .B(n12828), .Z(n15066) );
  XNOR2_X1 U14875 ( .A(n12370), .B(n12828), .ZN(n12371) );
  OAI222_X1 U14876 ( .A1(n13278), .A2(n12373), .B1(n13276), .B2(n12372), .C1(
        n15685), .C2(n12371), .ZN(n15067) );
  NAND2_X1 U14877 ( .A1(n15067), .A2(n15693), .ZN(n12378) );
  OAI22_X1 U14878 ( .A1(n15693), .A2(n12375), .B1(n12374), .B2(n15675), .ZN(
        n12376) );
  AOI21_X1 U14879 ( .B1(n15673), .B2(n15069), .A(n12376), .ZN(n12377) );
  OAI211_X1 U14880 ( .C1(n15054), .C2(n15066), .A(n12378), .B(n12377), .ZN(
        P3_U3221) );
  INV_X1 U14881 ( .A(n12379), .ZN(n12383) );
  OAI222_X1 U14882 ( .A1(n14891), .A2(n12381), .B1(n14885), .B2(n12383), .C1(
        P1_U3086), .C2(n12380), .ZN(P1_U3330) );
  OAI222_X1 U14883 ( .A1(n14072), .A2(n12384), .B1(n14075), .B2(n12383), .C1(
        n12382), .C2(P2_U3088), .ZN(P2_U3302) );
  INV_X1 U14884 ( .A(n12385), .ZN(n12386) );
  AOI21_X1 U14885 ( .B1(n12389), .B2(n12387), .A(n12386), .ZN(n14013) );
  XOR2_X1 U14886 ( .A(n12389), .B(n12388), .Z(n12390) );
  NAND2_X1 U14887 ( .A1(n12390), .A2(n13906), .ZN(n14011) );
  AND2_X1 U14888 ( .A1(n13643), .A2(n13617), .ZN(n12391) );
  AOI21_X1 U14889 ( .B1(n13641), .B2(n13602), .A(n12391), .ZN(n14010) );
  AOI21_X1 U14890 ( .B1(n14011), .B2(n14010), .A(n13926), .ZN(n12397) );
  OAI211_X1 U14891 ( .C1(n14063), .C2(n12392), .A(n11777), .B(n12427), .ZN(
        n14009) );
  OAI22_X1 U14892 ( .A1(n13919), .A2(n12393), .B1(n12473), .B2(n13916), .ZN(
        n12394) );
  AOI21_X1 U14893 ( .B1(n12475), .B2(n13933), .A(n12394), .ZN(n12395) );
  OAI21_X1 U14894 ( .B1(n14009), .B2(n13922), .A(n12395), .ZN(n12396) );
  AOI211_X1 U14895 ( .C1(n14013), .C2(n13924), .A(n12397), .B(n12396), .ZN(
        n12398) );
  INV_X1 U14896 ( .A(n12398), .ZN(P2_U3249) );
  INV_X1 U14897 ( .A(n12410), .ZN(n12408) );
  NAND2_X1 U14898 ( .A1(n14275), .A2(n12635), .ZN(n12400) );
  NAND2_X1 U14899 ( .A1(n12621), .A2(n14493), .ZN(n12399) );
  NAND2_X1 U14900 ( .A1(n12400), .A2(n12399), .ZN(n12401) );
  XNOR2_X1 U14901 ( .A(n12401), .B(n12618), .ZN(n12403) );
  NOR2_X1 U14902 ( .A1(n12644), .A2(n12492), .ZN(n12402) );
  AOI21_X1 U14903 ( .B1(n14275), .B2(n12621), .A(n12402), .ZN(n12404) );
  NAND2_X1 U14904 ( .A1(n12403), .A2(n12404), .ZN(n12484) );
  INV_X1 U14905 ( .A(n12403), .ZN(n12406) );
  INV_X1 U14906 ( .A(n12404), .ZN(n12405) );
  NAND2_X1 U14907 ( .A1(n12406), .A2(n12405), .ZN(n12407) );
  AND2_X1 U14908 ( .A1(n12484), .A2(n12407), .ZN(n12412) );
  NOR3_X1 U14909 ( .A1(n12409), .A2(n12408), .A3(n12412), .ZN(n12415) );
  NAND2_X1 U14910 ( .A1(n12411), .A2(n12410), .ZN(n12413) );
  NAND2_X1 U14911 ( .A1(n12413), .A2(n12412), .ZN(n12485) );
  INV_X1 U14912 ( .A(n12485), .ZN(n12414) );
  OAI21_X1 U14913 ( .B1(n12415), .B2(n12414), .A(n15114), .ZN(n12421) );
  NAND2_X1 U14914 ( .A1(n15107), .A2(n14492), .ZN(n12417) );
  OAI211_X1 U14915 ( .C1(n14203), .C2(n12418), .A(n12417), .B(n12416), .ZN(
        n12419) );
  AOI21_X1 U14916 ( .B1(n7677), .B2(n14205), .A(n12419), .ZN(n12420) );
  OAI211_X1 U14917 ( .C1(n7465), .C2(n15111), .A(n12421), .B(n12420), .ZN(
        P1_U3217) );
  XNOR2_X1 U14918 ( .A(n12422), .B(n12423), .ZN(n14006) );
  INV_X1 U14919 ( .A(n14006), .ZN(n12433) );
  XNOR2_X1 U14920 ( .A(n12424), .B(n12423), .ZN(n12426) );
  AND2_X1 U14921 ( .A1(n13642), .A2(n13617), .ZN(n12425) );
  AOI21_X1 U14922 ( .B1(n13640), .B2(n13602), .A(n12425), .ZN(n13565) );
  OAI21_X1 U14923 ( .B1(n12426), .B2(n13896), .A(n13565), .ZN(n14005) );
  AOI211_X1 U14924 ( .C1(n13443), .C2(n12427), .A(n8410), .B(n7175), .ZN(
        n14004) );
  NAND2_X1 U14925 ( .A1(n14004), .A2(n13930), .ZN(n12430) );
  INV_X1 U14926 ( .A(n12428), .ZN(n13567) );
  AOI22_X1 U14927 ( .A1(n13926), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n13567), 
        .B2(n13931), .ZN(n12429) );
  OAI211_X1 U14928 ( .C1(n14058), .C2(n13824), .A(n12430), .B(n12429), .ZN(
        n12431) );
  AOI21_X1 U14929 ( .B1(n13919), .B2(n14005), .A(n12431), .ZN(n12432) );
  OAI21_X1 U14930 ( .B1(n12433), .B2(n13902), .A(n12432), .ZN(P2_U3248) );
  NAND2_X1 U14931 ( .A1(n6796), .A2(n12435), .ZN(n12436) );
  XNOR2_X1 U14932 ( .A(n12434), .B(n12436), .ZN(n12443) );
  AND2_X1 U14933 ( .A1(P3_U3151), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n14972) );
  NOR2_X1 U14934 ( .A1(n12774), .A2(n13277), .ZN(n12437) );
  AOI211_X1 U14935 ( .C1(n12770), .C2(n12438), .A(n14972), .B(n12437), .ZN(
        n12439) );
  OAI21_X1 U14936 ( .B1(n13283), .B2(n12440), .A(n12439), .ZN(n12441) );
  AOI21_X1 U14937 ( .B1(n9897), .B2(n13282), .A(n12441), .ZN(n12442) );
  OAI21_X1 U14938 ( .B1(n12443), .B2(n12777), .A(n12442), .ZN(P3_U3181) );
  XNOR2_X1 U14939 ( .A(n12444), .B(n14439), .ZN(n14853) );
  AOI211_X1 U14940 ( .C1(n14851), .C2(n6693), .A(n14741), .B(n12514), .ZN(
        n14849) );
  INV_X1 U14941 ( .A(n14851), .ZN(n12445) );
  NOR2_X1 U14942 ( .A1(n12445), .A2(n15141), .ZN(n12448) );
  OAI22_X1 U14943 ( .A1(n15143), .A2(n12446), .B1(n14147), .B2(n15136), .ZN(
        n12447) );
  AOI211_X1 U14944 ( .C1(n14849), .C2(n15125), .A(n12448), .B(n12447), .ZN(
        n12455) );
  NAND2_X1 U14945 ( .A1(n12449), .A2(n15160), .ZN(n12453) );
  AOI21_X1 U14946 ( .B1(n15127), .B2(n12450), .A(n14439), .ZN(n12452) );
  AOI22_X1 U14947 ( .A1(n14761), .A2(n15134), .B1(n14762), .B2(n14489), .ZN(
        n12451) );
  OAI21_X1 U14948 ( .B1(n12453), .B2(n12452), .A(n12451), .ZN(n14850) );
  NAND2_X1 U14949 ( .A1(n14850), .A2(n15143), .ZN(n12454) );
  OAI211_X1 U14950 ( .C1(n14853), .C2(n14750), .A(n12455), .B(n12454), .ZN(
        P1_U3276) );
  XNOR2_X1 U14951 ( .A(n12475), .B(n13498), .ZN(n12456) );
  NAND2_X1 U14952 ( .A1(n13642), .A2(n13912), .ZN(n12457) );
  NAND2_X1 U14953 ( .A1(n12456), .A2(n12457), .ZN(n13441) );
  INV_X1 U14954 ( .A(n12456), .ZN(n12459) );
  INV_X1 U14955 ( .A(n12457), .ZN(n12458) );
  NAND2_X1 U14956 ( .A1(n12459), .A2(n12458), .ZN(n12460) );
  NAND2_X1 U14957 ( .A1(n13441), .A2(n12460), .ZN(n12470) );
  NAND2_X1 U14958 ( .A1(n12462), .A2(n12461), .ZN(n12467) );
  INV_X1 U14959 ( .A(n12463), .ZN(n12464) );
  OR2_X1 U14960 ( .A1(n12465), .A2(n12464), .ZN(n12466) );
  INV_X1 U14961 ( .A(n13442), .ZN(n12468) );
  AOI21_X1 U14962 ( .B1(n12470), .B2(n12469), .A(n12468), .ZN(n12477) );
  INV_X1 U14963 ( .A(n14010), .ZN(n12471) );
  AOI22_X1 U14964 ( .A1(n13605), .A2(n12471), .B1(P2_REG3_REG_16__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12472) );
  OAI21_X1 U14965 ( .B1(n12473), .B2(n13607), .A(n12472), .ZN(n12474) );
  AOI21_X1 U14966 ( .B1(n12475), .B2(n13624), .A(n12474), .ZN(n12476) );
  OAI21_X1 U14967 ( .B1(n12477), .B2(n13627), .A(n12476), .ZN(P2_U3198) );
  INV_X1 U14968 ( .A(n12478), .ZN(n14889) );
  AOI22_X1 U14969 ( .A1(n12479), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n14080), .ZN(n12480) );
  OAI21_X1 U14970 ( .B1(n14889), .B2(n14075), .A(n12480), .ZN(P2_U3301) );
  NAND2_X1 U14971 ( .A1(n14279), .A2(n12635), .ZN(n12482) );
  NAND2_X1 U14972 ( .A1(n12621), .A2(n14492), .ZN(n12481) );
  NAND2_X1 U14973 ( .A1(n12482), .A2(n12481), .ZN(n12483) );
  XNOR2_X1 U14974 ( .A(n12483), .B(n12646), .ZN(n12497) );
  AOI22_X1 U14975 ( .A1(n14279), .A2(n12621), .B1(n10728), .B2(n14492), .ZN(
        n12498) );
  XNOR2_X1 U14976 ( .A(n12497), .B(n12498), .ZN(n12488) );
  NAND2_X1 U14977 ( .A1(n12485), .A2(n12484), .ZN(n12487) );
  OAI21_X1 U14978 ( .B1(n12488), .B2(n12487), .A(n12486), .ZN(n12489) );
  NAND2_X1 U14979 ( .A1(n12489), .A2(n15114), .ZN(n12496) );
  NAND2_X1 U14980 ( .A1(n15107), .A2(n15108), .ZN(n12491) );
  OAI211_X1 U14981 ( .C1(n12492), .C2(n15086), .A(n12491), .B(n12490), .ZN(
        n12493) );
  AOI21_X1 U14982 ( .B1(n12494), .B2(n14205), .A(n12493), .ZN(n12495) );
  OAI211_X1 U14983 ( .C1(n15181), .C2(n15111), .A(n12496), .B(n12495), .ZN(
        P1_U3236) );
  INV_X1 U14984 ( .A(n14917), .ZN(n14940) );
  INV_X1 U14985 ( .A(n12497), .ZN(n12499) );
  NAND2_X1 U14986 ( .A1(n12499), .A2(n12498), .ZN(n12502) );
  AND2_X1 U14987 ( .A1(n12486), .A2(n12502), .ZN(n12505) );
  NOR2_X1 U14988 ( .A1(n12644), .A2(n14946), .ZN(n12500) );
  AOI21_X1 U14989 ( .B1(n14917), .B2(n12621), .A(n12500), .ZN(n12535) );
  AOI22_X1 U14990 ( .A1(n14917), .A2(n12635), .B1(n12621), .B2(n15108), .ZN(
        n12501) );
  XNOR2_X1 U14991 ( .A(n12501), .B(n12646), .ZN(n12534) );
  XOR2_X1 U14992 ( .A(n12535), .B(n12534), .Z(n12504) );
  OAI211_X1 U14993 ( .C1(n12505), .C2(n12504), .A(n15114), .B(n12539), .ZN(
        n12508) );
  AOI22_X1 U14994 ( .A1(n14491), .A2(n15134), .B1(n14762), .B2(n14492), .ZN(
        n14925) );
  NAND2_X1 U14995 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3086), .ZN(n15254)
         );
  OAI21_X1 U14996 ( .B1(n14203), .B2(n14925), .A(n15254), .ZN(n12506) );
  AOI21_X1 U14997 ( .B1(n14930), .B2(n14205), .A(n12506), .ZN(n12507) );
  OAI211_X1 U14998 ( .C1(n14940), .C2(n15111), .A(n12508), .B(n12507), .ZN(
        P1_U3224) );
  XNOR2_X1 U14999 ( .A(n14441), .B(n12510), .ZN(n14848) );
  XNOR2_X1 U15000 ( .A(n14441), .B(n12511), .ZN(n12512) );
  NAND2_X1 U15001 ( .A1(n12512), .A2(n15160), .ZN(n14846) );
  INV_X1 U15002 ( .A(n14846), .ZN(n12513) );
  OAI22_X1 U15003 ( .A1(n14162), .A2(n14947), .B1(n14310), .B2(n15131), .ZN(
        n14844) );
  OAI21_X1 U15004 ( .B1(n12513), .B2(n14844), .A(n15143), .ZN(n12520) );
  INV_X1 U15005 ( .A(n12514), .ZN(n12516) );
  INV_X1 U15006 ( .A(n14757), .ZN(n12515) );
  AOI211_X1 U15007 ( .C1(n14845), .C2(n12516), .A(n14741), .B(n12515), .ZN(
        n14843) );
  AOI22_X1 U15008 ( .A1(n14931), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n14181), 
        .B2(n14929), .ZN(n12517) );
  OAI21_X1 U15009 ( .B1(n14323), .B2(n15141), .A(n12517), .ZN(n12518) );
  AOI21_X1 U15010 ( .B1(n14843), .B2(n15125), .A(n12518), .ZN(n12519) );
  OAI211_X1 U15011 ( .C1(n14848), .C2(n14750), .A(n12520), .B(n12519), .ZN(
        P1_U3275) );
  OAI22_X1 U15012 ( .A1(n14368), .A2(n14947), .B1(n14666), .B2(n15131), .ZN(
        n12524) );
  OR3_X1 U15013 ( .A1(n12521), .A2(n7476), .A3(n14446), .ZN(n12522) );
  AOI211_X1 U15014 ( .C1(n14786), .C2(n14649), .A(n14741), .B(n6702), .ZN(
        n14785) );
  AOI22_X1 U15015 ( .A1(n14088), .A2(n14929), .B1(P1_REG2_REG_27__SCAN_IN), 
        .B2(n14765), .ZN(n12526) );
  OAI21_X1 U15016 ( .B1(n14093), .B2(n15141), .A(n12526), .ZN(n12528) );
  NOR2_X1 U15017 ( .A1(n14789), .A2(n14921), .ZN(n12527) );
  AOI211_X1 U15018 ( .C1(n14785), .C2(n15125), .A(n12528), .B(n12527), .ZN(
        n12529) );
  OAI21_X1 U15019 ( .B1(n14788), .B2(n14765), .A(n12529), .ZN(P1_U3266) );
  INV_X1 U15020 ( .A(n12530), .ZN(n12532) );
  OAI222_X1 U15021 ( .A1(n14072), .A2(n12533), .B1(n14075), .B2(n12532), .C1(
        n12531), .C2(P2_U3088), .ZN(P2_U3305) );
  INV_X1 U15022 ( .A(n12534), .ZN(n12537) );
  NAND2_X1 U15023 ( .A1(n12537), .A2(n12536), .ZN(n12538) );
  OAI22_X1 U15024 ( .A1(n15112), .A2(n12648), .B1(n15087), .B2(n12645), .ZN(
        n12540) );
  XNOR2_X1 U15025 ( .A(n12540), .B(n12618), .ZN(n12548) );
  OR2_X1 U15026 ( .A1(n15112), .A2(n12645), .ZN(n12542) );
  NAND2_X1 U15027 ( .A1(n10728), .A2(n14491), .ZN(n12541) );
  AND2_X1 U15028 ( .A1(n12542), .A2(n12541), .ZN(n12547) );
  NAND2_X1 U15029 ( .A1(n12548), .A2(n12547), .ZN(n15103) );
  NAND2_X1 U15030 ( .A1(n15164), .A2(n12635), .ZN(n12544) );
  NAND2_X1 U15031 ( .A1(n15106), .A2(n12621), .ZN(n12543) );
  NAND2_X1 U15032 ( .A1(n12544), .A2(n12543), .ZN(n12545) );
  XNOR2_X1 U15033 ( .A(n12545), .B(n12618), .ZN(n12551) );
  NOR2_X1 U15034 ( .A1(n14948), .A2(n12644), .ZN(n12546) );
  AOI21_X1 U15035 ( .B1(n15164), .B2(n12621), .A(n12546), .ZN(n12550) );
  XNOR2_X1 U15036 ( .A(n12551), .B(n12550), .ZN(n15090) );
  NOR2_X1 U15037 ( .A1(n12548), .A2(n12547), .ZN(n15102) );
  NOR2_X1 U15038 ( .A1(n15090), .A2(n15102), .ZN(n12549) );
  NAND2_X1 U15039 ( .A1(n12552), .A2(n12635), .ZN(n12554) );
  OR2_X1 U15040 ( .A1(n15132), .A2(n12645), .ZN(n12553) );
  NAND2_X1 U15041 ( .A1(n12554), .A2(n12553), .ZN(n12555) );
  XNOR2_X1 U15042 ( .A(n12555), .B(n12646), .ZN(n12557) );
  OAI22_X1 U15043 ( .A1(n7512), .A2(n12645), .B1(n15132), .B2(n12644), .ZN(
        n14199) );
  INV_X1 U15044 ( .A(n12556), .ZN(n12558) );
  NAND2_X1 U15045 ( .A1(n12558), .A2(n12557), .ZN(n12559) );
  NAND2_X1 U15046 ( .A1(n14198), .A2(n12559), .ZN(n14132) );
  OAI22_X1 U15047 ( .A1(n15148), .A2(n12648), .B1(n14307), .B2(n12645), .ZN(
        n12560) );
  XNOR2_X1 U15048 ( .A(n12560), .B(n12646), .ZN(n12561) );
  OAI22_X1 U15049 ( .A1(n15148), .A2(n12645), .B1(n14307), .B2(n12644), .ZN(
        n12562) );
  XNOR2_X1 U15050 ( .A(n12561), .B(n12562), .ZN(n14133) );
  INV_X1 U15051 ( .A(n12561), .ZN(n12564) );
  INV_X1 U15052 ( .A(n12562), .ZN(n12563) );
  NAND2_X1 U15053 ( .A1(n12564), .A2(n12563), .ZN(n12565) );
  NAND2_X1 U15054 ( .A1(n14851), .A2(n12635), .ZN(n12567) );
  NAND2_X1 U15055 ( .A1(n15135), .A2(n12621), .ZN(n12566) );
  NAND2_X1 U15056 ( .A1(n12567), .A2(n12566), .ZN(n12568) );
  XNOR2_X1 U15057 ( .A(n12568), .B(n12646), .ZN(n14142) );
  NAND2_X1 U15058 ( .A1(n14851), .A2(n12621), .ZN(n12570) );
  NAND2_X1 U15059 ( .A1(n15135), .A2(n10728), .ZN(n12569) );
  NAND2_X1 U15060 ( .A1(n12570), .A2(n12569), .ZN(n14141) );
  NOR2_X1 U15061 ( .A1(n14142), .A2(n14141), .ZN(n12572) );
  NAND2_X1 U15062 ( .A1(n14142), .A2(n14141), .ZN(n12571) );
  OAI22_X1 U15063 ( .A1(n14323), .A2(n12648), .B1(n14324), .B2(n12645), .ZN(
        n12573) );
  XNOR2_X1 U15064 ( .A(n12573), .B(n12646), .ZN(n12579) );
  OAI22_X1 U15065 ( .A1(n14323), .A2(n12645), .B1(n14324), .B2(n12644), .ZN(
        n12578) );
  XNOR2_X1 U15066 ( .A(n12579), .B(n12578), .ZN(n14180) );
  NAND2_X1 U15067 ( .A1(n14758), .A2(n12635), .ZN(n12575) );
  NAND2_X1 U15068 ( .A1(n14488), .A2(n12621), .ZN(n12574) );
  NAND2_X1 U15069 ( .A1(n12575), .A2(n12574), .ZN(n12576) );
  XNOR2_X1 U15070 ( .A(n12576), .B(n12618), .ZN(n12582) );
  NOR2_X1 U15071 ( .A1(n14162), .A2(n12644), .ZN(n12577) );
  AOI21_X1 U15072 ( .B1(n14758), .B2(n12621), .A(n12577), .ZN(n12581) );
  XNOR2_X1 U15073 ( .A(n12582), .B(n12581), .ZN(n14103) );
  NOR2_X1 U15074 ( .A1(n12579), .A2(n12578), .ZN(n14104) );
  NOR2_X1 U15075 ( .A1(n14103), .A2(n14104), .ZN(n12580) );
  OAI22_X1 U15076 ( .A1(n14746), .A2(n12645), .B1(n14336), .B2(n12644), .ZN(
        n12584) );
  OAI22_X1 U15077 ( .A1(n14746), .A2(n12648), .B1(n14336), .B2(n12645), .ZN(
        n12583) );
  XNOR2_X1 U15078 ( .A(n12583), .B(n12646), .ZN(n12585) );
  XOR2_X1 U15079 ( .A(n12584), .B(n12585), .Z(n14161) );
  NAND2_X1 U15080 ( .A1(n12585), .A2(n12584), .ZN(n12586) );
  NAND2_X1 U15081 ( .A1(n14827), .A2(n12635), .ZN(n12589) );
  NAND2_X1 U15082 ( .A1(n14487), .A2(n12621), .ZN(n12588) );
  NAND2_X1 U15083 ( .A1(n12589), .A2(n12588), .ZN(n12590) );
  XNOR2_X1 U15084 ( .A(n12590), .B(n12618), .ZN(n12593) );
  AND2_X1 U15085 ( .A1(n14487), .A2(n10728), .ZN(n12591) );
  AOI21_X1 U15086 ( .B1(n14827), .B2(n12621), .A(n12591), .ZN(n12592) );
  NAND2_X1 U15087 ( .A1(n12593), .A2(n12592), .ZN(n14169) );
  OAI21_X1 U15088 ( .B1(n12593), .B2(n12592), .A(n14169), .ZN(n14113) );
  OAI22_X1 U15089 ( .A1(n14820), .A2(n12648), .B1(n14344), .B2(n12645), .ZN(
        n12594) );
  XNOR2_X1 U15090 ( .A(n12594), .B(n12646), .ZN(n12596) );
  OAI22_X1 U15091 ( .A1(n14820), .A2(n12645), .B1(n14344), .B2(n12644), .ZN(
        n12595) );
  NAND2_X1 U15092 ( .A1(n12596), .A2(n12595), .ZN(n12597) );
  NAND2_X1 U15093 ( .A1(n14812), .A2(n12635), .ZN(n12600) );
  NAND2_X1 U15094 ( .A1(n14485), .A2(n12621), .ZN(n12599) );
  NAND2_X1 U15095 ( .A1(n12600), .A2(n12599), .ZN(n12601) );
  XNOR2_X1 U15096 ( .A(n12601), .B(n12618), .ZN(n12603) );
  AND2_X1 U15097 ( .A1(n14485), .A2(n10728), .ZN(n12602) );
  AOI21_X1 U15098 ( .B1(n14812), .B2(n12621), .A(n12602), .ZN(n12604) );
  NAND2_X1 U15099 ( .A1(n12603), .A2(n12604), .ZN(n14151) );
  INV_X1 U15100 ( .A(n12603), .ZN(n12606) );
  INV_X1 U15101 ( .A(n12604), .ZN(n12605) );
  NAND2_X1 U15102 ( .A1(n12606), .A2(n12605), .ZN(n12607) );
  OAI22_X1 U15103 ( .A1(n14690), .A2(n12648), .B1(n14665), .B2(n12645), .ZN(
        n12608) );
  XNOR2_X1 U15104 ( .A(n12608), .B(n12618), .ZN(n12611) );
  INV_X1 U15105 ( .A(n14665), .ZN(n14484) );
  NAND2_X1 U15106 ( .A1(n14484), .A2(n10728), .ZN(n12609) );
  NAND2_X1 U15107 ( .A1(n12611), .A2(n12612), .ZN(n14120) );
  INV_X1 U15108 ( .A(n12611), .ZN(n12614) );
  INV_X1 U15109 ( .A(n12612), .ZN(n12613) );
  NAND2_X1 U15110 ( .A1(n12614), .A2(n12613), .ZN(n12615) );
  NAND2_X1 U15111 ( .A1(n14119), .A2(n14120), .ZN(n12627) );
  NAND2_X1 U15112 ( .A1(n14674), .A2(n12635), .ZN(n12617) );
  NAND2_X1 U15113 ( .A1(n14483), .A2(n12621), .ZN(n12616) );
  NAND2_X1 U15114 ( .A1(n12617), .A2(n12616), .ZN(n12619) );
  XNOR2_X1 U15115 ( .A(n12619), .B(n12618), .ZN(n12622) );
  AND2_X1 U15116 ( .A1(n14483), .A2(n10728), .ZN(n12620) );
  AOI21_X1 U15117 ( .B1(n14674), .B2(n12621), .A(n12620), .ZN(n12623) );
  NAND2_X1 U15118 ( .A1(n12622), .A2(n12623), .ZN(n12628) );
  INV_X1 U15119 ( .A(n12622), .ZN(n12625) );
  INV_X1 U15120 ( .A(n12623), .ZN(n12624) );
  NAND2_X1 U15121 ( .A1(n12625), .A2(n12624), .ZN(n12626) );
  NAND2_X1 U15122 ( .A1(n12627), .A2(n14121), .ZN(n14123) );
  OAI22_X1 U15123 ( .A1(n14656), .A2(n12648), .B1(n14666), .B2(n12645), .ZN(
        n12629) );
  XNOR2_X1 U15124 ( .A(n12629), .B(n12646), .ZN(n12633) );
  OR2_X1 U15125 ( .A1(n14656), .A2(n12645), .ZN(n12631) );
  INV_X1 U15126 ( .A(n14666), .ZN(n14482) );
  NAND2_X1 U15127 ( .A1(n14482), .A2(n10728), .ZN(n12630) );
  NAND2_X1 U15128 ( .A1(n12631), .A2(n12630), .ZN(n12632) );
  NOR2_X1 U15129 ( .A1(n12633), .A2(n12632), .ZN(n12634) );
  AOI21_X1 U15130 ( .B1(n12633), .B2(n12632), .A(n12634), .ZN(n14189) );
  NAND2_X1 U15131 ( .A1(n14786), .A2(n12635), .ZN(n12637) );
  NAND2_X1 U15132 ( .A1(n14481), .A2(n12621), .ZN(n12636) );
  NAND2_X1 U15133 ( .A1(n12637), .A2(n12636), .ZN(n12638) );
  XNOR2_X1 U15134 ( .A(n12638), .B(n12646), .ZN(n12642) );
  NAND2_X1 U15135 ( .A1(n14786), .A2(n12621), .ZN(n12640) );
  NAND2_X1 U15136 ( .A1(n14481), .A2(n10728), .ZN(n12639) );
  NAND2_X1 U15137 ( .A1(n12640), .A2(n12639), .ZN(n12641) );
  NOR2_X1 U15138 ( .A1(n12642), .A2(n12641), .ZN(n12643) );
  AOI21_X1 U15139 ( .B1(n12642), .B2(n12641), .A(n12643), .ZN(n14087) );
  OAI22_X1 U15140 ( .A1(n14780), .A2(n12645), .B1(n14368), .B2(n12644), .ZN(
        n12647) );
  XNOR2_X1 U15141 ( .A(n12647), .B(n12646), .ZN(n12650) );
  OAI22_X1 U15142 ( .A1(n14780), .A2(n12648), .B1(n14368), .B2(n12645), .ZN(
        n12649) );
  XNOR2_X1 U15143 ( .A(n12650), .B(n12649), .ZN(n12651) );
  XNOR2_X1 U15144 ( .A(n12652), .B(n12651), .ZN(n12658) );
  NAND2_X1 U15145 ( .A1(n14481), .A2(n14762), .ZN(n12653) );
  OAI21_X1 U15146 ( .B1(n14392), .B2(n14947), .A(n12653), .ZN(n14777) );
  OAI22_X1 U15147 ( .A1(n14641), .A2(n15119), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n12654), .ZN(n12656) );
  NOR2_X1 U15148 ( .A1(n14780), .A2(n15111), .ZN(n12655) );
  AOI211_X1 U15149 ( .C1(n14195), .C2(n14777), .A(n12656), .B(n12655), .ZN(
        n12657) );
  OAI21_X1 U15150 ( .B1(n12658), .B2(n15092), .A(n12657), .ZN(P1_U3220) );
  OAI222_X1 U15151 ( .A1(n14072), .A2(n12660), .B1(n14075), .B2(n12659), .C1(
        n8332), .C2(P2_U3088), .ZN(P2_U3306) );
  INV_X1 U15152 ( .A(n12661), .ZN(n14078) );
  OAI222_X1 U15153 ( .A1(n14891), .A2(n12663), .B1(n14885), .B2(n14078), .C1(
        P1_U3086), .C2(n12662), .ZN(P1_U3327) );
  INV_X1 U15154 ( .A(n12664), .ZN(n12665) );
  XNOR2_X1 U15155 ( .A(n13086), .B(n12669), .ZN(n12677) );
  INV_X1 U15156 ( .A(n12677), .ZN(n12670) );
  NAND2_X1 U15157 ( .A1(n12670), .A2(n12788), .ZN(n12683) );
  INV_X1 U15158 ( .A(n12671), .ZN(n12672) );
  NAND4_X1 U15159 ( .A1(n12682), .A2(n12788), .A3(n12672), .A4(n12677), .ZN(
        n12681) );
  NAND2_X1 U15160 ( .A1(n12673), .A2(n12794), .ZN(n12675) );
  AOI22_X1 U15161 ( .A1(n13096), .A2(n12790), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12674) );
  OAI211_X1 U15162 ( .C1(n13091), .C2(n12792), .A(n12675), .B(n12674), .ZN(
        n12679) );
  NOR4_X1 U15163 ( .A1(n12677), .A2(n12676), .A3(n12777), .A4(n13112), .ZN(
        n12678) );
  AOI211_X1 U15164 ( .C1(n9897), .C2(n13095), .A(n12679), .B(n12678), .ZN(
        n12680) );
  OAI211_X1 U15165 ( .C1(n12683), .C2(n12682), .A(n12681), .B(n12680), .ZN(
        P3_U3160) );
  INV_X1 U15166 ( .A(n12685), .ZN(n12686) );
  NAND2_X1 U15167 ( .A1(n14880), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n12688) );
  INV_X1 U15168 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n14070) );
  NAND2_X1 U15169 ( .A1(n14070), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n12801) );
  INV_X1 U15170 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n14877) );
  NAND2_X1 U15171 ( .A1(n14877), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n12690) );
  AND2_X1 U15172 ( .A1(n12801), .A2(n12690), .ZN(n12691) );
  INV_X1 U15173 ( .A(n12800), .ZN(n12693) );
  OAI222_X1 U15174 ( .A1(P3_U3151), .A2(n12684), .B1(n12666), .B2(n12693), 
        .C1(n10310), .C2(n13440), .ZN(P3_U3265) );
  INV_X1 U15175 ( .A(n12694), .ZN(n12750) );
  AOI21_X1 U15176 ( .B1(n13146), .B2(n12695), .A(n12750), .ZN(n12700) );
  AOI22_X1 U15177 ( .A1(n13159), .A2(n12770), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12697) );
  NAND2_X1 U15178 ( .A1(n13168), .A2(n12790), .ZN(n12696) );
  OAI211_X1 U15179 ( .C1(n12726), .C2(n12774), .A(n12697), .B(n12696), .ZN(
        n12698) );
  AOI21_X1 U15180 ( .B1(n13163), .B2(n9897), .A(n12698), .ZN(n12699) );
  OAI21_X1 U15181 ( .B1(n12700), .B2(n12777), .A(n12699), .ZN(P3_U3156) );
  XNOR2_X1 U15182 ( .A(n12702), .B(n12701), .ZN(n12707) );
  NAND2_X1 U15183 ( .A1(n6674), .A2(n12794), .ZN(n12703) );
  NAND2_X1 U15184 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n13043)
         );
  OAI211_X1 U15185 ( .C1(n12792), .C2(n13248), .A(n12703), .B(n13043), .ZN(
        n12704) );
  AOI21_X1 U15186 ( .B1(n13226), .B2(n12790), .A(n12704), .ZN(n12706) );
  NAND2_X1 U15187 ( .A1(n13225), .A2(n9897), .ZN(n12705) );
  OAI211_X1 U15188 ( .C1(n12707), .C2(n12777), .A(n12706), .B(n12705), .ZN(
        P3_U3159) );
  INV_X1 U15189 ( .A(n12708), .ZN(n13398) );
  AOI21_X1 U15190 ( .B1(n12710), .B2(n12709), .A(n12777), .ZN(n12712) );
  NAND2_X1 U15191 ( .A1(n12712), .A2(n12711), .ZN(n12716) );
  AOI22_X1 U15192 ( .A1(n13159), .A2(n12794), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12713) );
  OAI21_X1 U15193 ( .B1(n6673), .B2(n12792), .A(n12713), .ZN(n12714) );
  AOI21_X1 U15194 ( .B1(n13198), .B2(n12790), .A(n12714), .ZN(n12715) );
  OAI211_X1 U15195 ( .C1(n13398), .C2(n12797), .A(n12716), .B(n12715), .ZN(
        P3_U3163) );
  INV_X1 U15196 ( .A(n12721), .ZN(n12751) );
  INV_X1 U15197 ( .A(n12720), .ZN(n12719) );
  AND2_X1 U15198 ( .A1(n12718), .A2(n12717), .ZN(n12722) );
  NOR3_X1 U15199 ( .A1(n12751), .A2(n12719), .A3(n12722), .ZN(n12724) );
  NAND2_X1 U15200 ( .A1(n12721), .A2(n12720), .ZN(n12723) );
  OAI21_X1 U15201 ( .B1(n12724), .B2(n6759), .A(n12788), .ZN(n12729) );
  AOI22_X1 U15202 ( .A1(n13130), .A2(n12790), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12725) );
  OAI21_X1 U15203 ( .B1(n12726), .B2(n12792), .A(n12725), .ZN(n12727) );
  AOI21_X1 U15204 ( .B1(n12794), .B2(n13127), .A(n12727), .ZN(n12728) );
  OAI211_X1 U15205 ( .C1(n13385), .C2(n12797), .A(n12729), .B(n12728), .ZN(
        P3_U3165) );
  XNOR2_X1 U15206 ( .A(n12730), .B(n13277), .ZN(n12731) );
  XNOR2_X1 U15207 ( .A(n12732), .B(n12731), .ZN(n12738) );
  NAND2_X1 U15208 ( .A1(n12790), .A2(n13267), .ZN(n12735) );
  INV_X1 U15209 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n12733) );
  NOR2_X1 U15210 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12733), .ZN(n14991) );
  AOI21_X1 U15211 ( .B1(n12794), .B2(n13234), .A(n14991), .ZN(n12734) );
  OAI211_X1 U15212 ( .C1(n13262), .C2(n12792), .A(n12735), .B(n12734), .ZN(
        n12736) );
  AOI21_X1 U15213 ( .B1(n13266), .B2(n9897), .A(n12736), .ZN(n12737) );
  OAI21_X1 U15214 ( .B1(n12738), .B2(n12777), .A(n12737), .ZN(P3_U3166) );
  AOI21_X1 U15215 ( .B1(n12741), .B2(n12740), .A(n12739), .ZN(n12746) );
  NAND2_X1 U15216 ( .A1(n12790), .A2(n13252), .ZN(n12743) );
  AND2_X1 U15217 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n15020) );
  AOI21_X1 U15218 ( .B1(n12794), .B2(n13219), .A(n15020), .ZN(n12742) );
  OAI211_X1 U15219 ( .C1(n13277), .C2(n12792), .A(n12743), .B(n12742), .ZN(
        n12744) );
  AOI21_X1 U15220 ( .B1(n13251), .B2(n9897), .A(n12744), .ZN(n12745) );
  OAI21_X1 U15221 ( .B1(n12746), .B2(n12777), .A(n12745), .ZN(P3_U3168) );
  INV_X1 U15222 ( .A(n12747), .ZN(n12749) );
  NOR3_X1 U15223 ( .A1(n12750), .A2(n12749), .A3(n12748), .ZN(n12752) );
  OAI21_X1 U15224 ( .B1(n12752), .B2(n12751), .A(n12788), .ZN(n12757) );
  OAI22_X1 U15225 ( .A1(n13178), .A2(n12792), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12753), .ZN(n12755) );
  NOR2_X1 U15226 ( .A1(n13149), .A2(n12774), .ZN(n12754) );
  AOI211_X1 U15227 ( .C1(n13151), .C2(n12790), .A(n12755), .B(n12754), .ZN(
        n12756) );
  OAI211_X1 U15228 ( .C1(n12797), .C2(n13325), .A(n12757), .B(n12756), .ZN(
        P3_U3169) );
  INV_X1 U15229 ( .A(n12758), .ZN(n12759) );
  AOI21_X1 U15230 ( .B1(n12761), .B2(n12760), .A(n12759), .ZN(n12766) );
  AOI22_X1 U15231 ( .A1(n12771), .A2(n12794), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12762) );
  OAI21_X1 U15232 ( .B1(n13207), .B2(n12792), .A(n12762), .ZN(n12764) );
  NOR2_X1 U15233 ( .A1(n13402), .A2(n12797), .ZN(n12763) );
  AOI211_X1 U15234 ( .C1(n13210), .C2(n12790), .A(n12764), .B(n12763), .ZN(
        n12765) );
  OAI21_X1 U15235 ( .B1(n12766), .B2(n12777), .A(n12765), .ZN(P3_U3173) );
  INV_X1 U15236 ( .A(n12767), .ZN(n12768) );
  AOI21_X1 U15237 ( .B1(n13159), .B2(n12769), .A(n12768), .ZN(n12778) );
  AOI22_X1 U15238 ( .A1(n12771), .A2(n12770), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12773) );
  NAND2_X1 U15239 ( .A1(n12790), .A2(n13182), .ZN(n12772) );
  OAI211_X1 U15240 ( .C1(n13178), .C2(n12774), .A(n12773), .B(n12772), .ZN(
        n12775) );
  AOI21_X1 U15241 ( .B1(n13181), .B2(n9897), .A(n12775), .ZN(n12776) );
  OAI21_X1 U15242 ( .B1(n12778), .B2(n12777), .A(n12776), .ZN(P3_U3175) );
  INV_X1 U15243 ( .A(n13240), .ZN(n13350) );
  OAI211_X1 U15244 ( .C1(n12781), .C2(n12780), .A(n12779), .B(n12788), .ZN(
        n12785) );
  NAND2_X1 U15245 ( .A1(n12794), .A2(n13235), .ZN(n12782) );
  NAND2_X1 U15246 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n15037)
         );
  OAI211_X1 U15247 ( .C1(n12792), .C2(n13263), .A(n12782), .B(n15037), .ZN(
        n12783) );
  AOI21_X1 U15248 ( .B1(n13237), .B2(n12790), .A(n12783), .ZN(n12784) );
  OAI211_X1 U15249 ( .C1(n13350), .C2(n12797), .A(n12785), .B(n12784), .ZN(
        P3_U3178) );
  OAI21_X1 U15250 ( .B1(n12787), .B2(n6688), .A(n12786), .ZN(n12789) );
  NAND2_X1 U15251 ( .A1(n12789), .A2(n12788), .ZN(n12796) );
  AOI22_X1 U15252 ( .A1(n13117), .A2(n12790), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12791) );
  OAI21_X1 U15253 ( .B1(n13149), .B2(n12792), .A(n12791), .ZN(n12793) );
  AOI21_X1 U15254 ( .B1(n13112), .B2(n12794), .A(n12793), .ZN(n12795) );
  OAI211_X1 U15255 ( .C1(n13381), .C2(n12797), .A(n12796), .B(n12795), .ZN(
        P3_U3180) );
  INV_X1 U15256 ( .A(n12834), .ZN(n12974) );
  NOR2_X1 U15257 ( .A1(n12798), .A2(n12974), .ZN(n12814) );
  NAND2_X1 U15258 ( .A1(n12802), .A2(n12801), .ZN(n12804) );
  XNOR2_X1 U15259 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .ZN(n12803) );
  XNOR2_X1 U15260 ( .A(n12804), .B(n12803), .ZN(n13434) );
  NAND2_X1 U15261 ( .A1(n13434), .A2(n12805), .ZN(n12808) );
  OR2_X1 U15262 ( .A1(n12806), .A2(n13429), .ZN(n12807) );
  NOR2_X1 U15263 ( .A1(n12812), .A2(n13069), .ZN(n12980) );
  INV_X1 U15264 ( .A(n12809), .ZN(n12994) );
  OAI21_X1 U15265 ( .B1(n13373), .B2(n12994), .A(n12810), .ZN(n12977) );
  NOR2_X1 U15266 ( .A1(n12980), .A2(n12977), .ZN(n12816) );
  OAI21_X1 U15267 ( .B1(n13373), .B2(n12811), .A(n12816), .ZN(n12813) );
  AOI22_X1 U15268 ( .A1(n12812), .A2(n13069), .B1(n13373), .B2(n12994), .ZN(
        n12817) );
  OAI22_X1 U15269 ( .A1(n12814), .A2(n12813), .B1(n13370), .B2(n12817), .ZN(
        n12815) );
  XNOR2_X1 U15270 ( .A(n12815), .B(n7356), .ZN(n12986) );
  INV_X1 U15271 ( .A(n12839), .ZN(n12818) );
  INV_X1 U15272 ( .A(n12967), .ZN(n12836) );
  INV_X1 U15273 ( .A(n13164), .ZN(n13157) );
  OR2_X1 U15274 ( .A1(n13144), .A2(n13157), .ZN(n12958) );
  INV_X1 U15275 ( .A(n12958), .ZN(n12833) );
  INV_X1 U15276 ( .A(n13175), .ZN(n13179) );
  INV_X1 U15277 ( .A(n13280), .ZN(n13272) );
  NOR3_X1 U15278 ( .A1(n12819), .A2(n15702), .A3(n12857), .ZN(n12822) );
  NAND3_X1 U15279 ( .A1(n12822), .A2(n12821), .A3(n12820), .ZN(n12826) );
  INV_X1 U15280 ( .A(n12823), .ZN(n12824) );
  NAND4_X1 U15281 ( .A1(n12863), .A2(n6678), .A3(n12886), .A4(n12824), .ZN(
        n12825) );
  NOR4_X1 U15282 ( .A1(n12826), .A2(n12825), .A3(n15645), .A4(n12891), .ZN(
        n12827) );
  NAND4_X1 U15283 ( .A1(n7622), .A2(n8656), .A3(n12828), .A4(n12827), .ZN(
        n12829) );
  NOR4_X1 U15284 ( .A1(n13259), .A2(n13272), .A3(n13295), .A4(n12829), .ZN(
        n12830) );
  NAND4_X1 U15285 ( .A1(n13224), .A2(n12934), .A3(n13250), .A4(n12830), .ZN(
        n12831) );
  NOR4_X1 U15286 ( .A1(n13179), .A2(n13196), .A3(n13204), .A4(n12831), .ZN(
        n12832) );
  NAND4_X1 U15287 ( .A1(n12834), .A2(n13135), .A3(n12833), .A4(n12832), .ZN(
        n12835) );
  INV_X1 U15288 ( .A(n12837), .ZN(n12838) );
  MUX2_X1 U15289 ( .A(n12839), .B(n12838), .S(n12963), .Z(n12841) );
  NAND3_X1 U15290 ( .A1(n13104), .A2(n13112), .A3(n12975), .ZN(n12840) );
  OAI21_X1 U15291 ( .B1(n12842), .B2(n12841), .A(n12840), .ZN(n12969) );
  MUX2_X1 U15292 ( .A(n12844), .B(n12843), .S(n12975), .Z(n12949) );
  NAND2_X1 U15293 ( .A1(n12846), .A2(n12845), .ZN(n12847) );
  AND2_X1 U15294 ( .A1(n12847), .A2(n12850), .ZN(n12852) );
  NAND3_X1 U15295 ( .A1(n12850), .A2(n12849), .A3(n12848), .ZN(n12851) );
  MUX2_X1 U15296 ( .A(n12852), .B(n12851), .S(n12975), .Z(n12858) );
  NAND3_X1 U15297 ( .A1(n12853), .A2(n12864), .A3(n12854), .ZN(n12855) );
  NAND2_X1 U15298 ( .A1(n12855), .A2(n12975), .ZN(n12856) );
  OAI21_X1 U15299 ( .B1(n12858), .B2(n12857), .A(n12856), .ZN(n12862) );
  AOI21_X1 U15300 ( .B1(n12861), .B2(n12859), .A(n12975), .ZN(n12860) );
  AOI21_X1 U15301 ( .B1(n12862), .B2(n12861), .A(n12860), .ZN(n12866) );
  OAI21_X1 U15302 ( .B1(n12864), .B2(n12975), .A(n12863), .ZN(n12865) );
  OAI21_X1 U15303 ( .B1(n12866), .B2(n12865), .A(n6678), .ZN(n12875) );
  NAND2_X1 U15304 ( .A1(n12878), .A2(n12867), .ZN(n12870) );
  NAND2_X1 U15305 ( .A1(n12870), .A2(n12963), .ZN(n12874) );
  INV_X1 U15306 ( .A(n12868), .ZN(n12872) );
  NOR2_X1 U15307 ( .A1(n12870), .A2(n12869), .ZN(n12871) );
  MUX2_X1 U15308 ( .A(n12872), .B(n12871), .S(n12963), .Z(n12873) );
  AOI21_X1 U15309 ( .B1(n12875), .B2(n12874), .A(n12873), .ZN(n12882) );
  AOI21_X1 U15310 ( .B1(n12877), .B2(n12876), .A(n12963), .ZN(n12881) );
  MUX2_X1 U15311 ( .A(n12878), .B(n12877), .S(n12963), .Z(n12879) );
  OAI211_X1 U15312 ( .C1(n12882), .C2(n12881), .A(n12880), .B(n12879), .ZN(
        n12887) );
  MUX2_X1 U15313 ( .A(n12884), .B(n12883), .S(n12975), .Z(n12885) );
  NAND3_X1 U15314 ( .A1(n12887), .A2(n12886), .A3(n12885), .ZN(n12901) );
  MUX2_X1 U15315 ( .A(n12889), .B(n12888), .S(n12963), .Z(n12890) );
  INV_X1 U15316 ( .A(n12890), .ZN(n12892) );
  NOR3_X1 U15317 ( .A1(n12892), .A2(n12891), .A3(n15645), .ZN(n12900) );
  MUX2_X1 U15318 ( .A(n12894), .B(n12893), .S(n12975), .Z(n12898) );
  MUX2_X1 U15319 ( .A(n12896), .B(n12895), .S(n12975), .Z(n12897) );
  OAI211_X1 U15320 ( .C1(n12898), .C2(n15645), .A(n12897), .B(n8656), .ZN(
        n12899) );
  AOI21_X1 U15321 ( .B1(n12901), .B2(n12900), .A(n12899), .ZN(n12910) );
  NAND2_X1 U15322 ( .A1(n12907), .A2(n12902), .ZN(n12905) );
  NAND2_X1 U15323 ( .A1(n12906), .A2(n12903), .ZN(n12904) );
  MUX2_X1 U15324 ( .A(n12905), .B(n12904), .S(n12975), .Z(n12909) );
  MUX2_X1 U15325 ( .A(n12907), .B(n12906), .S(n12963), .Z(n12908) );
  OAI211_X1 U15326 ( .C1(n12910), .C2(n12909), .A(n7622), .B(n12908), .ZN(
        n12915) );
  INV_X1 U15327 ( .A(n13295), .ZN(n12914) );
  MUX2_X1 U15328 ( .A(n12912), .B(n12911), .S(n12963), .Z(n12913) );
  NAND3_X1 U15329 ( .A1(n12915), .A2(n12914), .A3(n12913), .ZN(n12919) );
  MUX2_X1 U15330 ( .A(n12917), .B(n12916), .S(n12963), .Z(n12918) );
  NAND2_X1 U15331 ( .A1(n12919), .A2(n12918), .ZN(n12923) );
  AOI21_X1 U15332 ( .B1(n12921), .B2(n12920), .A(n12963), .ZN(n12922) );
  AOI21_X1 U15333 ( .B1(n12923), .B2(n13280), .A(n12922), .ZN(n12927) );
  AND2_X1 U15334 ( .A1(n12925), .A2(n12924), .ZN(n12926) );
  OAI22_X1 U15335 ( .A1(n12927), .A2(n7380), .B1(n12926), .B2(n12975), .ZN(
        n12929) );
  OR3_X1 U15336 ( .A1(n13266), .A2(n13277), .A3(n12975), .ZN(n12928) );
  AOI211_X1 U15337 ( .C1(n12929), .C2(n12928), .A(n13245), .B(n13242), .ZN(
        n12943) );
  INV_X1 U15338 ( .A(n12935), .ZN(n12932) );
  OAI211_X1 U15339 ( .C1(n12932), .C2(n12931), .A(n12939), .B(n12930), .ZN(
        n12938) );
  NAND2_X1 U15340 ( .A1(n12934), .A2(n7379), .ZN(n12936) );
  NAND3_X1 U15341 ( .A1(n12936), .A2(n12940), .A3(n12935), .ZN(n12937) );
  MUX2_X1 U15342 ( .A(n12938), .B(n12937), .S(n12975), .Z(n12942) );
  MUX2_X1 U15343 ( .A(n12940), .B(n12939), .S(n12975), .Z(n12941) );
  OAI211_X1 U15344 ( .C1(n12943), .C2(n12942), .A(n8802), .B(n12941), .ZN(
        n12947) );
  MUX2_X1 U15345 ( .A(n12945), .B(n12944), .S(n12963), .Z(n12946) );
  NAND3_X1 U15346 ( .A1(n12947), .A2(n13193), .A3(n12946), .ZN(n12948) );
  NAND3_X1 U15347 ( .A1(n13175), .A2(n12949), .A3(n12948), .ZN(n12956) );
  NAND2_X1 U15348 ( .A1(n12956), .A2(n12950), .ZN(n12953) );
  NAND3_X1 U15349 ( .A1(n12951), .A2(n13178), .A3(n13163), .ZN(n12952) );
  OAI211_X1 U15350 ( .C1(n12958), .C2(n12953), .A(n12952), .B(n12954), .ZN(
        n12962) );
  INV_X1 U15351 ( .A(n12954), .ZN(n12959) );
  NAND2_X1 U15352 ( .A1(n12956), .A2(n12955), .ZN(n12957) );
  OAI22_X1 U15353 ( .A1(n12960), .A2(n12959), .B1(n12958), .B2(n12957), .ZN(
        n12961) );
  MUX2_X1 U15354 ( .A(n12962), .B(n12961), .S(n12975), .Z(n12968) );
  MUX2_X1 U15355 ( .A(n12965), .B(n12964), .S(n12963), .Z(n12966) );
  OAI21_X1 U15356 ( .B1(n12971), .B2(n12975), .A(n12970), .ZN(n12972) );
  NAND2_X1 U15357 ( .A1(n12973), .A2(n12972), .ZN(n12979) );
  AOI21_X1 U15358 ( .B1(n12976), .B2(n12975), .A(n12974), .ZN(n12978) );
  INV_X1 U15359 ( .A(n12980), .ZN(n12981) );
  AOI21_X1 U15360 ( .B1(n12986), .B2(n12985), .A(n12984), .ZN(n12993) );
  NAND2_X1 U15361 ( .A1(n12988), .A2(n12987), .ZN(n12989) );
  OAI211_X1 U15362 ( .C1(n12990), .C2(n12992), .A(n12989), .B(P3_B_REG_SCAN_IN), .ZN(n12991) );
  OAI21_X1 U15363 ( .B1(n12993), .B2(n12992), .A(n12991), .ZN(P3_U3296) );
  MUX2_X1 U15364 ( .A(P3_DATAO_REG_30__SCAN_IN), .B(n12994), .S(P3_U3897), .Z(
        P3_U3521) );
  MUX2_X1 U15365 ( .A(P3_DATAO_REG_26__SCAN_IN), .B(n13127), .S(P3_U3897), .Z(
        P3_U3517) );
  MUX2_X1 U15366 ( .A(P3_DATAO_REG_22__SCAN_IN), .B(n13159), .S(P3_U3897), .Z(
        P3_U3513) );
  MUX2_X1 U15367 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(n6674), .S(P3_U3897), .Z(
        P3_U3511) );
  MUX2_X1 U15368 ( .A(P3_DATAO_REG_17__SCAN_IN), .B(n13234), .S(P3_U3897), .Z(
        P3_U3508) );
  MUX2_X1 U15369 ( .A(P3_DATAO_REG_11__SCAN_IN), .B(n15640), .S(P3_U3897), .Z(
        P3_U3502) );
  MUX2_X1 U15370 ( .A(P3_DATAO_REG_10__SCAN_IN), .B(n15043), .S(P3_U3897), .Z(
        P3_U3501) );
  MUX2_X1 U15371 ( .A(P3_DATAO_REG_5__SCAN_IN), .B(n12995), .S(P3_U3897), .Z(
        P3_U3496) );
  MUX2_X1 U15372 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(n15681), .S(P3_U3897), .Z(
        P3_U3494) );
  MUX2_X1 U15373 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(n15698), .S(P3_U3897), .Z(
        P3_U3493) );
  MUX2_X1 U15374 ( .A(P3_DATAO_REG_0__SCAN_IN), .B(n15699), .S(P3_U3897), .Z(
        P3_U3491) );
  NAND2_X1 U15375 ( .A1(P3_REG2_REG_12__SCAN_IN), .A2(n15590), .ZN(n12999) );
  OAI21_X1 U15376 ( .B1(P3_REG2_REG_12__SCAN_IN), .B2(n15590), .A(n12999), 
        .ZN(n15584) );
  NOR2_X1 U15377 ( .A1(n13020), .A2(n13000), .ZN(n13001) );
  NOR2_X1 U15378 ( .A1(n8683), .A2(n15600), .ZN(n15599) );
  XNOR2_X1 U15379 ( .A(n15625), .B(P3_REG2_REG_14__SCAN_IN), .ZN(n15617) );
  NOR2_X1 U15380 ( .A1(n13058), .A2(n13002), .ZN(n13003) );
  AOI22_X1 U15381 ( .A1(P3_REG2_REG_16__SCAN_IN), .A2(n14990), .B1(n13047), 
        .B2(n13004), .ZN(n14985) );
  NOR2_X1 U15382 ( .A1(n13060), .A2(n13005), .ZN(n13006) );
  INV_X1 U15383 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n13007) );
  AOI22_X1 U15384 ( .A1(P3_REG2_REG_18__SCAN_IN), .A2(n15023), .B1(n13046), 
        .B2(n13007), .ZN(n15033) );
  XNOR2_X1 U15385 ( .A(n13037), .B(n13008), .ZN(n13038) );
  XNOR2_X1 U15386 ( .A(n13009), .B(n13038), .ZN(n13067) );
  MUX2_X1 U15387 ( .A(n13007), .B(n13063), .S(n13027), .Z(n15028) );
  MUX2_X1 U15388 ( .A(n15008), .B(n13353), .S(n13027), .Z(n13032) );
  NOR2_X1 U15389 ( .A1(n13060), .A2(n13032), .ZN(n13034) );
  MUX2_X1 U15390 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n13027), .Z(n13018) );
  INV_X1 U15391 ( .A(n13018), .ZN(n13019) );
  MUX2_X1 U15392 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n13027), .Z(n13016) );
  INV_X1 U15393 ( .A(n13016), .ZN(n13017) );
  MUX2_X1 U15394 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n13027), .Z(n13013) );
  INV_X1 U15395 ( .A(n13013), .ZN(n13014) );
  OAI21_X1 U15396 ( .B1(n13012), .B2(n13011), .A(n13010), .ZN(n15577) );
  XNOR2_X1 U15397 ( .A(n13013), .B(n13015), .ZN(n15576) );
  XNOR2_X1 U15398 ( .A(n13016), .B(n13048), .ZN(n15594) );
  NAND2_X1 U15399 ( .A1(n15595), .A2(n15594), .ZN(n15593) );
  OAI21_X1 U15400 ( .B1(n13048), .B2(n13017), .A(n15593), .ZN(n15609) );
  XNOR2_X1 U15401 ( .A(n13018), .B(n15605), .ZN(n15610) );
  NOR2_X1 U15402 ( .A1(n15609), .A2(n15610), .ZN(n15608) );
  INV_X1 U15403 ( .A(n15617), .ZN(n13023) );
  INV_X1 U15404 ( .A(n15625), .ZN(n13022) );
  NAND2_X1 U15405 ( .A1(n15625), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n13056) );
  INV_X1 U15406 ( .A(n13056), .ZN(n13021) );
  AOI21_X1 U15407 ( .B1(n13022), .B2(n13365), .A(n13021), .ZN(n15621) );
  MUX2_X1 U15408 ( .A(n13023), .B(n15621), .S(n13027), .Z(n15632) );
  NAND2_X1 U15409 ( .A1(n15633), .A2(n15632), .ZN(n15631) );
  NAND2_X1 U15410 ( .A1(n15625), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n13024) );
  MUX2_X1 U15411 ( .A(n13024), .B(n13056), .S(n13027), .Z(n13025) );
  NAND2_X1 U15412 ( .A1(n15631), .A2(n13025), .ZN(n13026) );
  INV_X1 U15413 ( .A(n13026), .ZN(n13028) );
  XNOR2_X1 U15414 ( .A(n13026), .B(n14974), .ZN(n14978) );
  MUX2_X1 U15415 ( .A(P3_REG2_REG_15__SCAN_IN), .B(P3_REG1_REG_15__SCAN_IN), 
        .S(n13027), .Z(n14979) );
  NOR2_X1 U15416 ( .A1(n14978), .A2(n14979), .ZN(n14977) );
  MUX2_X1 U15417 ( .A(P3_REG2_REG_16__SCAN_IN), .B(P3_REG1_REG_16__SCAN_IN), 
        .S(n13027), .Z(n13030) );
  AND2_X1 U15418 ( .A1(n13030), .A2(n13047), .ZN(n14998) );
  INV_X1 U15419 ( .A(n13030), .ZN(n13031) );
  NAND2_X1 U15420 ( .A1(n13031), .A2(n14990), .ZN(n14997) );
  OAI21_X1 U15421 ( .B1(n15002), .B2(n14998), .A(n14997), .ZN(n15013) );
  AOI21_X1 U15422 ( .B1(n13060), .B2(n13032), .A(n13034), .ZN(n13033) );
  INV_X1 U15423 ( .A(n13033), .ZN(n15014) );
  NOR2_X1 U15424 ( .A1(n15013), .A2(n15014), .ZN(n15012) );
  NOR2_X1 U15425 ( .A1(n13034), .A2(n15012), .ZN(n13035) );
  XNOR2_X1 U15426 ( .A(n13046), .B(n13035), .ZN(n15029) );
  NAND2_X1 U15427 ( .A1(n15028), .A2(n15029), .ZN(n15027) );
  NAND2_X1 U15428 ( .A1(n15023), .A2(n13035), .ZN(n13036) );
  NAND2_X1 U15429 ( .A1(n15027), .A2(n13036), .ZN(n13042) );
  XNOR2_X1 U15430 ( .A(n13037), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n13064) );
  INV_X1 U15431 ( .A(n13038), .ZN(n13040) );
  MUX2_X1 U15432 ( .A(n13064), .B(n13040), .S(n13039), .Z(n13041) );
  XNOR2_X1 U15433 ( .A(n13042), .B(n13041), .ZN(n13045) );
  NAND2_X1 U15434 ( .A1(n15623), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n13044) );
  OAI211_X1 U15435 ( .C1(n13045), .C2(n15611), .A(n13044), .B(n13043), .ZN(
        n13065) );
  AOI22_X1 U15436 ( .A1(P3_REG1_REG_18__SCAN_IN), .A2(n13046), .B1(n15023), 
        .B2(n13063), .ZN(n15026) );
  AOI22_X1 U15437 ( .A1(P3_REG1_REG_16__SCAN_IN), .A2(n13047), .B1(n14990), 
        .B2(n13357), .ZN(n14989) );
  NAND2_X1 U15438 ( .A1(P3_REG1_REG_12__SCAN_IN), .A2(n15590), .ZN(n13053) );
  AOI22_X1 U15439 ( .A1(P3_REG1_REG_12__SCAN_IN), .A2(n15590), .B1(n13048), 
        .B2(n8667), .ZN(n15587) );
  NAND2_X1 U15440 ( .A1(n15573), .A2(n13051), .ZN(n13052) );
  NAND2_X1 U15441 ( .A1(P3_REG1_REG_11__SCAN_IN), .A2(n15570), .ZN(n15569) );
  NAND2_X1 U15442 ( .A1(n15605), .A2(n13054), .ZN(n13055) );
  NAND2_X1 U15443 ( .A1(P3_REG1_REG_13__SCAN_IN), .A2(n15602), .ZN(n15601) );
  NAND2_X1 U15444 ( .A1(n13055), .A2(n15601), .ZN(n15620) );
  NAND2_X1 U15445 ( .A1(n15621), .A2(n15620), .ZN(n15619) );
  NAND2_X1 U15446 ( .A1(n13056), .A2(n15619), .ZN(n13057) );
  NAND2_X1 U15447 ( .A1(n14974), .A2(n13057), .ZN(n13059) );
  XNOR2_X1 U15448 ( .A(n13058), .B(n13057), .ZN(n14971) );
  NAND2_X1 U15449 ( .A1(P3_REG1_REG_15__SCAN_IN), .A2(n14971), .ZN(n14970) );
  NAND2_X1 U15450 ( .A1(n13059), .A2(n14970), .ZN(n14988) );
  NAND2_X1 U15451 ( .A1(n14989), .A2(n14988), .ZN(n14987) );
  OAI21_X1 U15452 ( .B1(n14990), .B2(n13357), .A(n14987), .ZN(n13061) );
  NAND2_X1 U15453 ( .A1(n15016), .A2(n13061), .ZN(n13062) );
  XNOR2_X1 U15454 ( .A(n13061), .B(n13060), .ZN(n15010) );
  NAND2_X1 U15455 ( .A1(P3_REG1_REG_17__SCAN_IN), .A2(n15010), .ZN(n15009) );
  NAND2_X1 U15456 ( .A1(n13062), .A2(n15009), .ZN(n15025) );
  NAND2_X1 U15457 ( .A1(n15026), .A2(n15025), .ZN(n15024) );
  OAI21_X1 U15458 ( .B1(n13067), .B2(n15636), .A(n13066), .ZN(P3_U3201) );
  NAND2_X1 U15459 ( .A1(n13070), .A2(n15710), .ZN(n13076) );
  AOI21_X1 U15460 ( .B1(n13368), .B2(n13076), .A(n13303), .ZN(n13072) );
  AOI21_X1 U15461 ( .B1(n15714), .B2(P3_REG2_REG_31__SCAN_IN), .A(n13072), 
        .ZN(n13071) );
  OAI21_X1 U15462 ( .B1(n13370), .B2(n13297), .A(n13071), .ZN(P3_U3202) );
  AOI21_X1 U15463 ( .B1(n15714), .B2(P3_REG2_REG_30__SCAN_IN), .A(n13072), 
        .ZN(n13073) );
  OAI21_X1 U15464 ( .B1(n13373), .B2(n13297), .A(n13073), .ZN(P3_U3203) );
  INV_X1 U15465 ( .A(n13074), .ZN(n13082) );
  NAND2_X1 U15466 ( .A1(n13075), .A2(n15693), .ZN(n13081) );
  OAI21_X1 U15467 ( .B1(n15693), .B2(n13077), .A(n13076), .ZN(n13078) );
  AOI21_X1 U15468 ( .B1(n13079), .B2(n15673), .A(n13078), .ZN(n13080) );
  OAI211_X1 U15469 ( .C1(n13082), .C2(n15054), .A(n13081), .B(n13080), .ZN(
        P3_U3204) );
  INV_X1 U15470 ( .A(n13083), .ZN(n13084) );
  NOR2_X1 U15471 ( .A1(n13085), .A2(n13084), .ZN(n13087) );
  XNOR2_X1 U15472 ( .A(n13087), .B(n13086), .ZN(n13309) );
  INV_X1 U15473 ( .A(n13309), .ZN(n13100) );
  AOI211_X1 U15474 ( .C1(n13090), .C2(n13089), .A(n15685), .B(n13088), .ZN(
        n13094) );
  OAI22_X1 U15475 ( .A1(n13092), .A2(n13278), .B1(n13091), .B2(n13276), .ZN(
        n13093) );
  OR2_X1 U15476 ( .A1(n13094), .A2(n13093), .ZN(n13308) );
  INV_X1 U15477 ( .A(n13095), .ZN(n13377) );
  AOI22_X1 U15478 ( .A1(n13096), .A2(n15710), .B1(n15714), .B2(
        P3_REG2_REG_28__SCAN_IN), .ZN(n13097) );
  OAI21_X1 U15479 ( .B1(n13377), .B2(n13297), .A(n13097), .ZN(n13098) );
  AOI21_X1 U15480 ( .B1(n13308), .B2(n15693), .A(n13098), .ZN(n13099) );
  OAI21_X1 U15481 ( .B1(n13100), .B2(n15054), .A(n13099), .ZN(P3_U3205) );
  INV_X1 U15482 ( .A(n13101), .ZN(n13108) );
  AOI22_X1 U15483 ( .A1(n13102), .A2(n15710), .B1(n13303), .B2(
        P3_REG2_REG_27__SCAN_IN), .ZN(n13103) );
  OAI21_X1 U15484 ( .B1(n13104), .B2(n13297), .A(n13103), .ZN(n13105) );
  AOI21_X1 U15485 ( .B1(n13106), .B2(n15711), .A(n13105), .ZN(n13107) );
  OAI21_X1 U15486 ( .B1(n13108), .B2(n13303), .A(n13107), .ZN(P3_U3206) );
  XOR2_X1 U15487 ( .A(n13111), .B(n13110), .Z(n13115) );
  NAND2_X1 U15488 ( .A1(n13112), .A2(n15697), .ZN(n13113) );
  OAI21_X1 U15489 ( .B1(n13149), .B2(n13276), .A(n13113), .ZN(n13114) );
  AOI21_X1 U15490 ( .B1(n13115), .B2(n15703), .A(n13114), .ZN(n13116) );
  OAI21_X1 U15491 ( .B1(n15707), .B2(n13312), .A(n13116), .ZN(n13313) );
  AOI22_X1 U15492 ( .A1(n13117), .A2(n15710), .B1(n15714), .B2(
        P3_REG2_REG_26__SCAN_IN), .ZN(n13120) );
  NAND2_X1 U15493 ( .A1(n13118), .A2(n15673), .ZN(n13119) );
  OAI211_X1 U15494 ( .C1(n13312), .C2(n13121), .A(n13120), .B(n13119), .ZN(
        n13122) );
  AOI21_X1 U15495 ( .B1(n13313), .B2(n15693), .A(n13122), .ZN(n13123) );
  INV_X1 U15496 ( .A(n13123), .ZN(P3_U3207) );
  OAI211_X1 U15497 ( .C1(n13126), .C2(n13125), .A(n13124), .B(n15703), .ZN(
        n13129) );
  AOI22_X1 U15498 ( .A1(n13127), .A2(n15697), .B1(n13160), .B2(n15700), .ZN(
        n13128) );
  INV_X1 U15499 ( .A(n13130), .ZN(n13132) );
  INV_X1 U15500 ( .A(P3_REG2_REG_25__SCAN_IN), .ZN(n13131) );
  OAI22_X1 U15501 ( .A1(n13132), .A2(n15675), .B1(n15693), .B2(n13131), .ZN(
        n13133) );
  AOI21_X1 U15502 ( .B1(n13134), .B2(n15673), .A(n13133), .ZN(n13138) );
  XNOR2_X1 U15503 ( .A(n13136), .B(n13135), .ZN(n13317) );
  NAND2_X1 U15504 ( .A1(n13317), .A2(n15649), .ZN(n13137) );
  OAI211_X1 U15505 ( .C1(n13319), .C2(n15714), .A(n13138), .B(n13137), .ZN(
        P3_U3208) );
  NAND2_X1 U15506 ( .A1(n13167), .A2(n13139), .ZN(n13140) );
  NAND2_X1 U15507 ( .A1(n13140), .A2(n13144), .ZN(n13142) );
  NAND2_X1 U15508 ( .A1(n13142), .A2(n13141), .ZN(n13322) );
  OAI211_X1 U15509 ( .C1(n13145), .C2(n13144), .A(n13143), .B(n15703), .ZN(
        n13148) );
  NAND2_X1 U15510 ( .A1(n13146), .A2(n15700), .ZN(n13147) );
  OAI211_X1 U15511 ( .C1(n13149), .C2(n13278), .A(n13148), .B(n13147), .ZN(
        n13150) );
  AOI21_X1 U15512 ( .B1(n15680), .B2(n13322), .A(n13150), .ZN(n13324) );
  AOI22_X1 U15513 ( .A1(n13151), .A2(n15710), .B1(n15714), .B2(
        P3_REG2_REG_24__SCAN_IN), .ZN(n13152) );
  OAI21_X1 U15514 ( .B1(n13325), .B2(n13297), .A(n13152), .ZN(n13153) );
  AOI21_X1 U15515 ( .B1(n13322), .B2(n15711), .A(n13153), .ZN(n13154) );
  OAI21_X1 U15516 ( .B1(n13324), .B2(n13303), .A(n13154), .ZN(P3_U3209) );
  INV_X1 U15517 ( .A(n13155), .ZN(n13158) );
  OAI211_X1 U15518 ( .C1(n13158), .C2(n13157), .A(n13156), .B(n15703), .ZN(
        n13162) );
  AOI22_X1 U15519 ( .A1(n13160), .A2(n15697), .B1(n15700), .B2(n13159), .ZN(
        n13161) );
  NAND2_X1 U15520 ( .A1(n13162), .A2(n13161), .ZN(n13326) );
  INV_X1 U15521 ( .A(n13163), .ZN(n13390) );
  OR2_X1 U15522 ( .A1(n13165), .A2(n13164), .ZN(n13166) );
  AND2_X1 U15523 ( .A1(n13167), .A2(n13166), .ZN(n13327) );
  NAND2_X1 U15524 ( .A1(n13327), .A2(n15649), .ZN(n13170) );
  AOI22_X1 U15525 ( .A1(n13303), .A2(P3_REG2_REG_23__SCAN_IN), .B1(n13168), 
        .B2(n15710), .ZN(n13169) );
  OAI211_X1 U15526 ( .C1(n13390), .C2(n13297), .A(n13170), .B(n13169), .ZN(
        n13171) );
  AOI21_X1 U15527 ( .B1(n13326), .B2(n15693), .A(n13171), .ZN(n13172) );
  INV_X1 U15528 ( .A(n13172), .ZN(P3_U3210) );
  NAND2_X1 U15529 ( .A1(n13216), .A2(n13173), .ZN(n13191) );
  NAND2_X1 U15530 ( .A1(n13191), .A2(n13174), .ZN(n13176) );
  XNOR2_X1 U15531 ( .A(n13176), .B(n13175), .ZN(n13177) );
  OAI222_X1 U15532 ( .A1(n13276), .A2(n13208), .B1(n13278), .B2(n13178), .C1(
        n15685), .C2(n13177), .ZN(n13330) );
  INV_X1 U15533 ( .A(n13330), .ZN(n13186) );
  XNOR2_X1 U15534 ( .A(n13180), .B(n13179), .ZN(n13331) );
  INV_X1 U15535 ( .A(n13181), .ZN(n13394) );
  AOI22_X1 U15536 ( .A1(n13303), .A2(P3_REG2_REG_22__SCAN_IN), .B1(n15710), 
        .B2(n13182), .ZN(n13183) );
  OAI21_X1 U15537 ( .B1(n13394), .B2(n13297), .A(n13183), .ZN(n13184) );
  AOI21_X1 U15538 ( .B1(n13331), .B2(n15649), .A(n13184), .ZN(n13185) );
  OAI21_X1 U15539 ( .B1(n13186), .B2(n15714), .A(n13185), .ZN(P3_U3211) );
  NAND2_X1 U15540 ( .A1(n13216), .A2(n13187), .ZN(n13189) );
  AND2_X1 U15541 ( .A1(n13189), .A2(n13188), .ZN(n13192) );
  AOI21_X1 U15542 ( .B1(n13193), .B2(n13192), .A(n7675), .ZN(n13194) );
  OAI222_X1 U15543 ( .A1(n13278), .A2(n13195), .B1(n13276), .B2(n6673), .C1(
        n15685), .C2(n13194), .ZN(n13334) );
  INV_X1 U15544 ( .A(n13334), .ZN(n13202) );
  XNOR2_X1 U15545 ( .A(n13197), .B(n13196), .ZN(n13335) );
  AOI22_X1 U15546 ( .A1(n13303), .A2(P3_REG2_REG_21__SCAN_IN), .B1(n15710), 
        .B2(n13198), .ZN(n13199) );
  OAI21_X1 U15547 ( .B1(n13398), .B2(n13297), .A(n13199), .ZN(n13200) );
  AOI21_X1 U15548 ( .B1(n13335), .B2(n15649), .A(n13200), .ZN(n13201) );
  OAI21_X1 U15549 ( .B1(n13202), .B2(n13303), .A(n13201), .ZN(P3_U3212) );
  NAND2_X1 U15550 ( .A1(n13216), .A2(n13203), .ZN(n13205) );
  XNOR2_X1 U15551 ( .A(n13205), .B(n13204), .ZN(n13206) );
  OAI222_X1 U15552 ( .A1(n13278), .A2(n13208), .B1(n13276), .B2(n13207), .C1(
        n13206), .C2(n15685), .ZN(n13338) );
  INV_X1 U15553 ( .A(n13338), .ZN(n13214) );
  XNOR2_X1 U15554 ( .A(n13209), .B(n8802), .ZN(n13339) );
  AOI22_X1 U15555 ( .A1(n13303), .A2(P3_REG2_REG_20__SCAN_IN), .B1(n15710), 
        .B2(n13210), .ZN(n13211) );
  OAI21_X1 U15556 ( .B1(n13402), .B2(n13297), .A(n13211), .ZN(n13212) );
  AOI21_X1 U15557 ( .B1(n13339), .B2(n15649), .A(n13212), .ZN(n13213) );
  OAI21_X1 U15558 ( .B1(n13214), .B2(n13303), .A(n13213), .ZN(P3_U3213) );
  INV_X1 U15559 ( .A(n13215), .ZN(n13218) );
  INV_X1 U15560 ( .A(n13224), .ZN(n13217) );
  OAI211_X1 U15561 ( .C1(n13218), .C2(n13217), .A(n15703), .B(n13216), .ZN(
        n13222) );
  AOI22_X1 U15562 ( .A1(n6674), .A2(n15697), .B1(n15700), .B2(n13219), .ZN(
        n13221) );
  NAND2_X1 U15563 ( .A1(n13222), .A2(n13221), .ZN(n13342) );
  INV_X1 U15564 ( .A(n13342), .ZN(n13230) );
  XOR2_X1 U15565 ( .A(n13223), .B(n13224), .Z(n13343) );
  INV_X1 U15566 ( .A(n13225), .ZN(n13406) );
  AOI22_X1 U15567 ( .A1(n13303), .A2(P3_REG2_REG_19__SCAN_IN), .B1(n15710), 
        .B2(n13226), .ZN(n13227) );
  OAI21_X1 U15568 ( .B1(n13406), .B2(n13297), .A(n13227), .ZN(n13228) );
  AOI21_X1 U15569 ( .B1(n13343), .B2(n15649), .A(n13228), .ZN(n13229) );
  OAI21_X1 U15570 ( .B1(n13230), .B2(n15714), .A(n13229), .ZN(P3_U3214) );
  INV_X1 U15571 ( .A(n13231), .ZN(n13233) );
  OAI21_X1 U15572 ( .B1(n13233), .B2(n13242), .A(n13232), .ZN(n13236) );
  AOI222_X1 U15573 ( .A1(n15703), .A2(n13236), .B1(n13235), .B2(n15697), .C1(
        n13234), .C2(n15700), .ZN(n13349) );
  INV_X1 U15574 ( .A(n13237), .ZN(n13238) );
  OAI22_X1 U15575 ( .A1(n15693), .A2(n13007), .B1(n13238), .B2(n15675), .ZN(
        n13239) );
  AOI21_X1 U15576 ( .B1(n13240), .B2(n15673), .A(n13239), .ZN(n13244) );
  NAND2_X1 U15577 ( .A1(n13241), .A2(n13242), .ZN(n13346) );
  NAND3_X1 U15578 ( .A1(n13347), .A2(n13346), .A3(n15649), .ZN(n13243) );
  OAI211_X1 U15579 ( .C1(n13349), .C2(n13303), .A(n13244), .B(n13243), .ZN(
        P3_U3215) );
  XNOR2_X1 U15580 ( .A(n13246), .B(n13245), .ZN(n13247) );
  OAI222_X1 U15581 ( .A1(n13278), .A2(n13248), .B1(n13276), .B2(n13277), .C1(
        n13247), .C2(n15685), .ZN(n13351) );
  INV_X1 U15582 ( .A(n13351), .ZN(n13256) );
  XNOR2_X1 U15583 ( .A(n13249), .B(n13250), .ZN(n13352) );
  INV_X1 U15584 ( .A(n13251), .ZN(n13411) );
  AOI22_X1 U15585 ( .A1(n13303), .A2(P3_REG2_REG_17__SCAN_IN), .B1(n15710), 
        .B2(n13252), .ZN(n13253) );
  OAI21_X1 U15586 ( .B1(n13411), .B2(n13297), .A(n13253), .ZN(n13254) );
  AOI21_X1 U15587 ( .B1(n13352), .B2(n15649), .A(n13254), .ZN(n13255) );
  OAI21_X1 U15588 ( .B1(n13256), .B2(n13303), .A(n13255), .ZN(P3_U3216) );
  NAND2_X1 U15589 ( .A1(n13258), .A2(n13257), .ZN(n13260) );
  XNOR2_X1 U15590 ( .A(n13260), .B(n13259), .ZN(n13261) );
  OAI222_X1 U15591 ( .A1(n13278), .A2(n13263), .B1(n13276), .B2(n13262), .C1(
        n13261), .C2(n15685), .ZN(n13355) );
  INV_X1 U15592 ( .A(n13355), .ZN(n13271) );
  XNOR2_X1 U15593 ( .A(n13265), .B(n13264), .ZN(n13356) );
  INV_X1 U15594 ( .A(n13266), .ZN(n13415) );
  AOI22_X1 U15595 ( .A1(n13303), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n15710), 
        .B2(n13267), .ZN(n13268) );
  OAI21_X1 U15596 ( .B1(n13415), .B2(n13297), .A(n13268), .ZN(n13269) );
  AOI21_X1 U15597 ( .B1(n13356), .B2(n15649), .A(n13269), .ZN(n13270) );
  OAI21_X1 U15598 ( .B1(n13271), .B2(n13303), .A(n13270), .ZN(P3_U3217) );
  XNOR2_X1 U15599 ( .A(n13273), .B(n13272), .ZN(n13274) );
  OAI222_X1 U15600 ( .A1(n13278), .A2(n13277), .B1(n13276), .B2(n13275), .C1(
        n13274), .C2(n15685), .ZN(n13359) );
  INV_X1 U15601 ( .A(n13359), .ZN(n13288) );
  OAI21_X1 U15602 ( .B1(n13281), .B2(n13280), .A(n13279), .ZN(n13360) );
  INV_X1 U15603 ( .A(n13282), .ZN(n13419) );
  INV_X1 U15604 ( .A(n13283), .ZN(n13284) );
  AOI22_X1 U15605 ( .A1(n13303), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n15710), 
        .B2(n13284), .ZN(n13285) );
  OAI21_X1 U15606 ( .B1(n13419), .B2(n13297), .A(n13285), .ZN(n13286) );
  AOI21_X1 U15607 ( .B1(n13360), .B2(n15649), .A(n13286), .ZN(n13287) );
  OAI21_X1 U15608 ( .B1(n13288), .B2(n15714), .A(n13287), .ZN(P3_U3218) );
  OAI211_X1 U15609 ( .C1(n13290), .C2(n13295), .A(n13289), .B(n15703), .ZN(
        n13294) );
  AOI22_X1 U15610 ( .A1(n15700), .A2(n13292), .B1(n13291), .B2(n15697), .ZN(
        n13293) );
  NAND2_X1 U15611 ( .A1(n13294), .A2(n13293), .ZN(n13363) );
  INV_X1 U15612 ( .A(n13363), .ZN(n13304) );
  XNOR2_X1 U15613 ( .A(n13296), .B(n13295), .ZN(n13364) );
  NOR2_X1 U15614 ( .A1(n13423), .A2(n13297), .ZN(n13301) );
  INV_X1 U15615 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n13299) );
  OAI22_X1 U15616 ( .A1(n15693), .A2(n13299), .B1(n13298), .B2(n15675), .ZN(
        n13300) );
  AOI211_X1 U15617 ( .C1(n13364), .C2(n15649), .A(n13301), .B(n13300), .ZN(
        n13302) );
  OAI21_X1 U15618 ( .B1(n13304), .B2(n13303), .A(n13302), .ZN(P3_U3219) );
  NOR2_X1 U15619 ( .A1(n13368), .A2(n15749), .ZN(n13306) );
  AOI21_X1 U15620 ( .B1(P3_REG1_REG_31__SCAN_IN), .B2(n15749), .A(n13306), 
        .ZN(n13305) );
  OAI21_X1 U15621 ( .B1(n13370), .B2(n13367), .A(n13305), .ZN(P3_U3490) );
  AOI21_X1 U15622 ( .B1(P3_REG1_REG_30__SCAN_IN), .B2(n15749), .A(n13306), 
        .ZN(n13307) );
  OAI21_X1 U15623 ( .B1(n13373), .B2(n13367), .A(n13307), .ZN(P3_U3489) );
  INV_X1 U15624 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n13310) );
  AOI21_X1 U15625 ( .B1(n13309), .B2(n15739), .A(n13308), .ZN(n13374) );
  MUX2_X1 U15626 ( .A(n13310), .B(n13374), .S(n15751), .Z(n13311) );
  OAI21_X1 U15627 ( .B1(n13377), .B2(n13367), .A(n13311), .ZN(P3_U3487) );
  INV_X1 U15628 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n13315) );
  INV_X1 U15629 ( .A(n13312), .ZN(n13314) );
  AOI21_X1 U15630 ( .B1(n15734), .B2(n13314), .A(n13313), .ZN(n13378) );
  MUX2_X1 U15631 ( .A(n13315), .B(n13378), .S(n15751), .Z(n13316) );
  OAI21_X1 U15632 ( .B1(n13381), .B2(n13367), .A(n13316), .ZN(P3_U3485) );
  INV_X1 U15633 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n13320) );
  NAND2_X1 U15634 ( .A1(n13317), .A2(n15739), .ZN(n13318) );
  MUX2_X1 U15635 ( .A(n13320), .B(n13382), .S(n15751), .Z(n13321) );
  OAI21_X1 U15636 ( .B1(n13385), .B2(n13367), .A(n13321), .ZN(P3_U3484) );
  NAND2_X1 U15637 ( .A1(n13322), .A2(n15734), .ZN(n13323) );
  OAI211_X1 U15638 ( .C1(n13325), .C2(n15730), .A(n13324), .B(n13323), .ZN(
        n13386) );
  MUX2_X1 U15639 ( .A(P3_REG1_REG_24__SCAN_IN), .B(n13386), .S(n15751), .Z(
        P3_U3483) );
  INV_X1 U15640 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n13328) );
  AOI21_X1 U15641 ( .B1(n13327), .B2(n15739), .A(n13326), .ZN(n13387) );
  MUX2_X1 U15642 ( .A(n13328), .B(n13387), .S(n15751), .Z(n13329) );
  OAI21_X1 U15643 ( .B1(n13390), .B2(n13367), .A(n13329), .ZN(P3_U3482) );
  INV_X1 U15644 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n13332) );
  AOI21_X1 U15645 ( .B1(n15739), .B2(n13331), .A(n13330), .ZN(n13391) );
  MUX2_X1 U15646 ( .A(n13332), .B(n13391), .S(n15751), .Z(n13333) );
  OAI21_X1 U15647 ( .B1(n13394), .B2(n13367), .A(n13333), .ZN(P3_U3481) );
  INV_X1 U15648 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n13336) );
  AOI21_X1 U15649 ( .B1(n15739), .B2(n13335), .A(n13334), .ZN(n13395) );
  MUX2_X1 U15650 ( .A(n13336), .B(n13395), .S(n15751), .Z(n13337) );
  OAI21_X1 U15651 ( .B1(n13398), .B2(n13367), .A(n13337), .ZN(P3_U3480) );
  INV_X1 U15652 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n13340) );
  AOI21_X1 U15653 ( .B1(n13339), .B2(n15739), .A(n13338), .ZN(n13399) );
  MUX2_X1 U15654 ( .A(n13340), .B(n13399), .S(n15751), .Z(n13341) );
  OAI21_X1 U15655 ( .B1(n13402), .B2(n13367), .A(n13341), .ZN(P3_U3479) );
  INV_X1 U15656 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n13344) );
  AOI21_X1 U15657 ( .B1(n15739), .B2(n13343), .A(n13342), .ZN(n13403) );
  MUX2_X1 U15658 ( .A(n13344), .B(n13403), .S(n15751), .Z(n13345) );
  OAI21_X1 U15659 ( .B1(n13406), .B2(n13367), .A(n13345), .ZN(P3_U3478) );
  NAND3_X1 U15660 ( .A1(n13347), .A2(n15739), .A3(n13346), .ZN(n13348) );
  OAI211_X1 U15661 ( .C1(n13350), .C2(n15730), .A(n13349), .B(n13348), .ZN(
        n13407) );
  MUX2_X1 U15662 ( .A(P3_REG1_REG_18__SCAN_IN), .B(n13407), .S(n15751), .Z(
        P3_U3477) );
  AOI21_X1 U15663 ( .B1(n13352), .B2(n15739), .A(n13351), .ZN(n13408) );
  MUX2_X1 U15664 ( .A(n13353), .B(n13408), .S(n15751), .Z(n13354) );
  OAI21_X1 U15665 ( .B1(n13411), .B2(n13367), .A(n13354), .ZN(P3_U3476) );
  AOI21_X1 U15666 ( .B1(n13356), .B2(n15739), .A(n13355), .ZN(n13412) );
  MUX2_X1 U15667 ( .A(n13357), .B(n13412), .S(n15751), .Z(n13358) );
  OAI21_X1 U15668 ( .B1(n13415), .B2(n13367), .A(n13358), .ZN(P3_U3475) );
  AOI21_X1 U15669 ( .B1(n15739), .B2(n13360), .A(n13359), .ZN(n13416) );
  MUX2_X1 U15670 ( .A(n13361), .B(n13416), .S(n15751), .Z(n13362) );
  OAI21_X1 U15671 ( .B1(n13419), .B2(n13367), .A(n13362), .ZN(P3_U3474) );
  AOI21_X1 U15672 ( .B1(n15739), .B2(n13364), .A(n13363), .ZN(n13420) );
  MUX2_X1 U15673 ( .A(n13365), .B(n13420), .S(n15751), .Z(n13366) );
  OAI21_X1 U15674 ( .B1(n13367), .B2(n13423), .A(n13366), .ZN(P3_U3473) );
  NOR2_X1 U15675 ( .A1(n13368), .A2(n15743), .ZN(n13371) );
  AOI21_X1 U15676 ( .B1(P3_REG0_REG_31__SCAN_IN), .B2(n15743), .A(n13371), 
        .ZN(n13369) );
  OAI21_X1 U15677 ( .B1(n13370), .B2(n13424), .A(n13369), .ZN(P3_U3458) );
  AOI21_X1 U15678 ( .B1(n15743), .B2(P3_REG0_REG_30__SCAN_IN), .A(n13371), 
        .ZN(n13372) );
  OAI21_X1 U15679 ( .B1(n13373), .B2(n13424), .A(n13372), .ZN(P3_U3457) );
  MUX2_X1 U15680 ( .A(n13375), .B(n13374), .S(n15741), .Z(n13376) );
  OAI21_X1 U15681 ( .B1(n13377), .B2(n13424), .A(n13376), .ZN(P3_U3455) );
  MUX2_X1 U15682 ( .A(n13379), .B(n13378), .S(n15741), .Z(n13380) );
  OAI21_X1 U15683 ( .B1(n13381), .B2(n13424), .A(n13380), .ZN(P3_U3453) );
  MUX2_X1 U15684 ( .A(n13383), .B(n13382), .S(n15741), .Z(n13384) );
  OAI21_X1 U15685 ( .B1(n13385), .B2(n13424), .A(n13384), .ZN(P3_U3452) );
  MUX2_X1 U15686 ( .A(P3_REG0_REG_24__SCAN_IN), .B(n13386), .S(n15741), .Z(
        P3_U3451) );
  MUX2_X1 U15687 ( .A(n13388), .B(n13387), .S(n15741), .Z(n13389) );
  OAI21_X1 U15688 ( .B1(n13390), .B2(n13424), .A(n13389), .ZN(P3_U3450) );
  MUX2_X1 U15689 ( .A(n13392), .B(n13391), .S(n15741), .Z(n13393) );
  OAI21_X1 U15690 ( .B1(n13394), .B2(n13424), .A(n13393), .ZN(P3_U3449) );
  MUX2_X1 U15691 ( .A(n13396), .B(n13395), .S(n15741), .Z(n13397) );
  OAI21_X1 U15692 ( .B1(n13398), .B2(n13424), .A(n13397), .ZN(P3_U3448) );
  INV_X1 U15693 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n13400) );
  MUX2_X1 U15694 ( .A(n13400), .B(n13399), .S(n15741), .Z(n13401) );
  OAI21_X1 U15695 ( .B1(n13402), .B2(n13424), .A(n13401), .ZN(P3_U3447) );
  INV_X1 U15696 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n13404) );
  MUX2_X1 U15697 ( .A(n13404), .B(n13403), .S(n15741), .Z(n13405) );
  OAI21_X1 U15698 ( .B1(n13406), .B2(n13424), .A(n13405), .ZN(P3_U3446) );
  MUX2_X1 U15699 ( .A(P3_REG0_REG_18__SCAN_IN), .B(n13407), .S(n15741), .Z(
        P3_U3444) );
  MUX2_X1 U15700 ( .A(n13409), .B(n13408), .S(n15741), .Z(n13410) );
  OAI21_X1 U15701 ( .B1(n13411), .B2(n13424), .A(n13410), .ZN(P3_U3441) );
  MUX2_X1 U15702 ( .A(n13413), .B(n13412), .S(n15741), .Z(n13414) );
  OAI21_X1 U15703 ( .B1(n13415), .B2(n13424), .A(n13414), .ZN(P3_U3438) );
  INV_X1 U15704 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n13417) );
  MUX2_X1 U15705 ( .A(n13417), .B(n13416), .S(n15741), .Z(n13418) );
  OAI21_X1 U15706 ( .B1(n13419), .B2(n13424), .A(n13418), .ZN(P3_U3435) );
  MUX2_X1 U15707 ( .A(n13421), .B(n13420), .S(n15741), .Z(n13422) );
  OAI21_X1 U15708 ( .B1(n13424), .B2(n13423), .A(n13422), .ZN(P3_U3432) );
  MUX2_X1 U15709 ( .A(P3_D_REG_1__SCAN_IN), .B(n13425), .S(n13426), .Z(
        P3_U3377) );
  MUX2_X1 U15710 ( .A(P3_D_REG_0__SCAN_IN), .B(n13427), .S(n13426), .Z(
        P3_U3376) );
  NAND3_X1 U15711 ( .A1(n6968), .A2(P3_IR_REG_31__SCAN_IN), .A3(
        P3_STATE_REG_SCAN_IN), .ZN(n13430) );
  OAI22_X1 U15712 ( .A1(n13431), .A2(n13430), .B1(n13429), .B2(n13440), .ZN(
        n13432) );
  AOI21_X1 U15713 ( .B1(n13434), .B2(n13433), .A(n13432), .ZN(n13435) );
  INV_X1 U15714 ( .A(n13435), .ZN(P3_U3264) );
  INV_X1 U15715 ( .A(n13436), .ZN(n13438) );
  OAI222_X1 U15716 ( .A1(n13440), .A2(n13439), .B1(n12666), .B2(n13438), .C1(
        n13437), .C2(P3_U3151), .ZN(P3_U3266) );
  XNOR2_X1 U15717 ( .A(n13443), .B(n13498), .ZN(n13444) );
  NAND2_X1 U15718 ( .A1(n13641), .A2(n13912), .ZN(n13445) );
  NAND2_X1 U15719 ( .A1(n13444), .A2(n13445), .ZN(n13449) );
  INV_X1 U15720 ( .A(n13444), .ZN(n13447) );
  INV_X1 U15721 ( .A(n13445), .ZN(n13446) );
  NAND2_X1 U15722 ( .A1(n13447), .A2(n13446), .ZN(n13448) );
  AND2_X1 U15723 ( .A1(n13449), .A2(n13448), .ZN(n13563) );
  INV_X1 U15724 ( .A(n13600), .ZN(n13455) );
  XNOR2_X1 U15725 ( .A(n14053), .B(n13498), .ZN(n13450) );
  NAND2_X1 U15726 ( .A1(n13640), .A2(n13912), .ZN(n13451) );
  XNOR2_X1 U15727 ( .A(n13450), .B(n13451), .ZN(n13599) );
  INV_X1 U15728 ( .A(n13450), .ZN(n13453) );
  INV_X1 U15729 ( .A(n13451), .ZN(n13452) );
  XNOR2_X1 U15730 ( .A(n13893), .B(n13498), .ZN(n13456) );
  NAND2_X1 U15731 ( .A1(n13639), .A2(n13912), .ZN(n13457) );
  NAND2_X1 U15732 ( .A1(n13456), .A2(n13457), .ZN(n13461) );
  INV_X1 U15733 ( .A(n13456), .ZN(n13459) );
  INV_X1 U15734 ( .A(n13457), .ZN(n13458) );
  NAND2_X1 U15735 ( .A1(n13459), .A2(n13458), .ZN(n13460) );
  AND2_X1 U15736 ( .A1(n13461), .A2(n13460), .ZN(n13521) );
  XNOR2_X1 U15737 ( .A(n13986), .B(n13498), .ZN(n13462) );
  NAND2_X1 U15738 ( .A1(n13638), .A2(n13912), .ZN(n13463) );
  NAND2_X1 U15739 ( .A1(n13462), .A2(n13463), .ZN(n13582) );
  INV_X1 U15740 ( .A(n13462), .ZN(n13465) );
  INV_X1 U15741 ( .A(n13463), .ZN(n13464) );
  NAND2_X1 U15742 ( .A1(n13465), .A2(n13464), .ZN(n13584) );
  XNOR2_X1 U15743 ( .A(n13859), .B(n13537), .ZN(n13468) );
  NAND2_X1 U15744 ( .A1(n13637), .A2(n13912), .ZN(n13466) );
  XNOR2_X1 U15745 ( .A(n13468), .B(n13466), .ZN(n13546) );
  NAND2_X1 U15746 ( .A1(n13545), .A2(n13546), .ZN(n13470) );
  INV_X1 U15747 ( .A(n13466), .ZN(n13467) );
  NAND2_X1 U15748 ( .A1(n13468), .A2(n13467), .ZN(n13469) );
  NAND2_X1 U15749 ( .A1(n13470), .A2(n13469), .ZN(n13473) );
  XNOR2_X1 U15750 ( .A(n13975), .B(n13498), .ZN(n13471) );
  NAND2_X1 U15751 ( .A1(n13636), .A2(n13912), .ZN(n13589) );
  NAND2_X1 U15752 ( .A1(n13590), .A2(n13589), .ZN(n13588) );
  INV_X1 U15753 ( .A(n13471), .ZN(n13472) );
  OR2_X1 U15754 ( .A1(n13473), .A2(n13472), .ZN(n13474) );
  XNOR2_X1 U15755 ( .A(n13970), .B(n13485), .ZN(n13475) );
  AND2_X1 U15756 ( .A1(n13635), .A2(n13912), .ZN(n13504) );
  NAND2_X1 U15757 ( .A1(n13503), .A2(n13504), .ZN(n13479) );
  INV_X1 U15758 ( .A(n13475), .ZN(n13476) );
  OR2_X1 U15759 ( .A1(n13477), .A2(n13476), .ZN(n13478) );
  XNOR2_X1 U15760 ( .A(n13965), .B(n13537), .ZN(n13482) );
  NAND2_X1 U15761 ( .A1(n13634), .A2(n13912), .ZN(n13480) );
  XNOR2_X1 U15762 ( .A(n13482), .B(n13480), .ZN(n13571) );
  NAND2_X1 U15763 ( .A1(n13570), .A2(n13571), .ZN(n13484) );
  INV_X1 U15764 ( .A(n13480), .ZN(n13481) );
  NAND2_X1 U15765 ( .A1(n13482), .A2(n13481), .ZN(n13483) );
  NAND2_X2 U15766 ( .A1(n13484), .A2(n13483), .ZN(n13554) );
  XNOR2_X1 U15767 ( .A(n14041), .B(n13485), .ZN(n13487) );
  NOR2_X1 U15768 ( .A1(n13486), .A2(n11777), .ZN(n13488) );
  XNOR2_X1 U15769 ( .A(n13487), .B(n13488), .ZN(n13553) );
  INV_X1 U15770 ( .A(n13487), .ZN(n13489) );
  NAND2_X1 U15771 ( .A1(n13489), .A2(n13488), .ZN(n13490) );
  XNOR2_X1 U15772 ( .A(n13778), .B(n13498), .ZN(n13492) );
  NAND2_X1 U15773 ( .A1(n13632), .A2(n13912), .ZN(n13493) );
  NAND2_X1 U15774 ( .A1(n13492), .A2(n13493), .ZN(n13497) );
  INV_X1 U15775 ( .A(n13492), .ZN(n13495) );
  INV_X1 U15776 ( .A(n13493), .ZN(n13494) );
  NAND2_X1 U15777 ( .A1(n13495), .A2(n13494), .ZN(n13496) );
  NAND2_X1 U15778 ( .A1(n13497), .A2(n13496), .ZN(n13613) );
  XNOR2_X1 U15779 ( .A(n13766), .B(n13498), .ZN(n13530) );
  NOR2_X1 U15780 ( .A1(n13616), .A2(n11777), .ZN(n13531) );
  XNOR2_X1 U15781 ( .A(n13530), .B(n13531), .ZN(n13534) );
  XNOR2_X1 U15782 ( .A(n13534), .B(n13535), .ZN(n13502) );
  AOI22_X1 U15783 ( .A1(n8388), .A2(n13602), .B1(n13617), .B2(n13632), .ZN(
        n13757) );
  AOI22_X1 U15784 ( .A1(n13764), .A2(n13623), .B1(P2_REG3_REG_27__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13499) );
  OAI21_X1 U15785 ( .B1(n13757), .B2(n13621), .A(n13499), .ZN(n13500) );
  AOI21_X1 U15786 ( .B1(n13948), .B2(n13624), .A(n13500), .ZN(n13501) );
  OAI21_X1 U15787 ( .B1(n13502), .B2(n13627), .A(n13501), .ZN(P2_U3186) );
  XNOR2_X1 U15788 ( .A(n13503), .B(n13504), .ZN(n13509) );
  OAI22_X1 U15789 ( .A1(n13555), .A2(n13615), .B1(n13505), .B2(n13577), .ZN(
        n13830) );
  AOI22_X1 U15790 ( .A1(n13830), .A2(n13605), .B1(P2_REG3_REG_23__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13506) );
  OAI21_X1 U15791 ( .B1(n13832), .B2(n13607), .A(n13506), .ZN(n13507) );
  AOI21_X1 U15792 ( .B1(n13970), .B2(n13624), .A(n13507), .ZN(n13508) );
  OAI21_X1 U15793 ( .B1(n13509), .B2(n13627), .A(n13508), .ZN(P2_U3188) );
  AOI21_X1 U15794 ( .B1(n13511), .B2(n13510), .A(n13627), .ZN(n13513) );
  NAND2_X1 U15795 ( .A1(n13513), .A2(n13512), .ZN(n13518) );
  AOI22_X1 U15796 ( .A1(n13515), .A2(n13624), .B1(n13605), .B2(n13514), .ZN(
        n13517) );
  MUX2_X1 U15797 ( .A(n13607), .B(P2_STATE_REG_SCAN_IN), .S(
        P2_REG3_REG_3__SCAN_IN), .Z(n13516) );
  NAND3_X1 U15798 ( .A1(n13518), .A2(n13517), .A3(n13516), .ZN(P2_U3190) );
  INV_X1 U15799 ( .A(n13893), .ZN(n13992) );
  OAI21_X1 U15800 ( .B1(n13522), .B2(n13521), .A(n13520), .ZN(n13523) );
  NAND2_X1 U15801 ( .A1(n13523), .A2(n13591), .ZN(n13529) );
  INV_X1 U15802 ( .A(n13888), .ZN(n13527) );
  NAND2_X1 U15803 ( .A1(n13638), .A2(n13602), .ZN(n13525) );
  NAND2_X1 U15804 ( .A1(n13640), .A2(n13617), .ZN(n13524) );
  AND2_X1 U15805 ( .A1(n13525), .A2(n13524), .ZN(n13990) );
  NAND2_X1 U15806 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n13720)
         );
  OAI21_X1 U15807 ( .B1(n13621), .B2(n13990), .A(n13720), .ZN(n13526) );
  AOI21_X1 U15808 ( .B1(n13527), .B2(n13623), .A(n13526), .ZN(n13528) );
  OAI211_X1 U15809 ( .C1(n13992), .C2(n13597), .A(n13529), .B(n13528), .ZN(
        P2_U3191) );
  INV_X1 U15810 ( .A(n13530), .ZN(n13533) );
  INV_X1 U15811 ( .A(n13531), .ZN(n13532) );
  NOR2_X1 U15812 ( .A1(n13536), .A2(n11777), .ZN(n13538) );
  XNOR2_X1 U15813 ( .A(n13538), .B(n13537), .ZN(n13539) );
  AOI22_X1 U15814 ( .A1(n13542), .A2(n13605), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13543) );
  OAI211_X1 U15815 ( .C1(n13750), .C2(n13607), .A(n13544), .B(n13543), .ZN(
        P2_U3192) );
  XNOR2_X1 U15816 ( .A(n13545), .B(n13546), .ZN(n13552) );
  AND2_X1 U15817 ( .A1(n13638), .A2(n13617), .ZN(n13547) );
  AOI21_X1 U15818 ( .B1(n13636), .B2(n13602), .A(n13547), .ZN(n13865) );
  OAI22_X1 U15819 ( .A1(n13621), .A2(n13865), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13548), .ZN(n13550) );
  NOR2_X1 U15820 ( .A1(n14048), .A2(n13597), .ZN(n13549) );
  AOI211_X1 U15821 ( .C1(n13623), .C2(n13855), .A(n13550), .B(n13549), .ZN(
        n13551) );
  OAI21_X1 U15822 ( .B1(n13552), .B2(n13627), .A(n13551), .ZN(P2_U3195) );
  XNOR2_X1 U15823 ( .A(n13554), .B(n13553), .ZN(n13560) );
  OAI22_X1 U15824 ( .A1(n13556), .A2(n13615), .B1(n13555), .B2(n13577), .ZN(
        n13788) );
  AOI22_X1 U15825 ( .A1(n13788), .A2(n13605), .B1(P2_REG3_REG_25__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13557) );
  OAI21_X1 U15826 ( .B1(n13795), .B2(n13607), .A(n13557), .ZN(n13558) );
  AOI21_X1 U15827 ( .B1(n13797), .B2(n13624), .A(n13558), .ZN(n13559) );
  OAI21_X1 U15828 ( .B1(n13560), .B2(n13627), .A(n13559), .ZN(P2_U3197) );
  OAI21_X1 U15829 ( .B1(n13563), .B2(n13562), .A(n13561), .ZN(n13564) );
  NAND2_X1 U15830 ( .A1(n13564), .A2(n13591), .ZN(n13569) );
  AND2_X1 U15831 ( .A1(P2_U3088), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n15447) );
  NOR2_X1 U15832 ( .A1(n13621), .A2(n13565), .ZN(n13566) );
  AOI211_X1 U15833 ( .C1(n13623), .C2(n13567), .A(n15447), .B(n13566), .ZN(
        n13568) );
  OAI211_X1 U15834 ( .C1(n14058), .C2(n13597), .A(n13569), .B(n13568), .ZN(
        P2_U3200) );
  XNOR2_X1 U15835 ( .A(n13570), .B(n13571), .ZN(n13576) );
  AOI22_X1 U15836 ( .A1(n13633), .A2(n13602), .B1(n13617), .B2(n13635), .ZN(
        n13805) );
  OAI22_X1 U15837 ( .A1(n13805), .A2(n13621), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13572), .ZN(n13573) );
  AOI21_X1 U15838 ( .B1(n13813), .B2(n13623), .A(n13573), .ZN(n13575) );
  NAND2_X1 U15839 ( .A1(n13965), .A2(n13624), .ZN(n13574) );
  OAI211_X1 U15840 ( .C1(n13576), .C2(n13627), .A(n13575), .B(n13574), .ZN(
        P2_U3201) );
  OAI22_X1 U15841 ( .A1(n13579), .A2(n13615), .B1(n13578), .B2(n13577), .ZN(
        n13875) );
  AOI22_X1 U15842 ( .A1(n13605), .A2(n13875), .B1(P2_REG3_REG_20__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13580) );
  OAI21_X1 U15843 ( .B1(n13877), .B2(n13607), .A(n13580), .ZN(n13586) );
  AOI21_X1 U15844 ( .B1(n13584), .B2(n13582), .A(n13581), .ZN(n13583) );
  AOI211_X1 U15845 ( .C1(n6734), .C2(n13584), .A(n13627), .B(n13583), .ZN(
        n13585) );
  AOI211_X1 U15846 ( .C1(n13986), .C2(n13624), .A(n13586), .B(n13585), .ZN(
        n13587) );
  INV_X1 U15847 ( .A(n13587), .ZN(P2_U3205) );
  INV_X1 U15848 ( .A(n13975), .ZN(n13598) );
  OAI21_X1 U15849 ( .B1(n13590), .B2(n13589), .A(n13588), .ZN(n13592) );
  NAND2_X1 U15850 ( .A1(n13592), .A2(n13591), .ZN(n13596) );
  AOI22_X1 U15851 ( .A1(n13635), .A2(n13602), .B1(n13617), .B2(n13637), .ZN(
        n13839) );
  OAI22_X1 U15852 ( .A1(n13621), .A2(n13839), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13593), .ZN(n13594) );
  AOI21_X1 U15853 ( .B1(n13843), .B2(n13623), .A(n13594), .ZN(n13595) );
  OAI211_X1 U15854 ( .C1(n13598), .C2(n13597), .A(n13596), .B(n13595), .ZN(
        P2_U3207) );
  XNOR2_X1 U15855 ( .A(n13600), .B(n13599), .ZN(n13610) );
  INV_X1 U15856 ( .A(n13601), .ZN(n13917) );
  NAND2_X1 U15857 ( .A1(P2_U3088), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n13684)
         );
  NAND2_X1 U15858 ( .A1(n13639), .A2(n13602), .ZN(n13604) );
  NAND2_X1 U15859 ( .A1(n13641), .A2(n13617), .ZN(n13603) );
  NAND2_X1 U15860 ( .A1(n13604), .A2(n13603), .ZN(n13905) );
  NAND2_X1 U15861 ( .A1(n13605), .A2(n13905), .ZN(n13606) );
  OAI211_X1 U15862 ( .C1(n13607), .C2(n13917), .A(n13684), .B(n13606), .ZN(
        n13608) );
  AOI21_X1 U15863 ( .B1(n14053), .B2(n13624), .A(n13608), .ZN(n13609) );
  OAI21_X1 U15864 ( .B1(n13610), .B2(n13627), .A(n13609), .ZN(P2_U3210) );
  INV_X1 U15865 ( .A(n13611), .ZN(n13612) );
  AOI21_X1 U15866 ( .B1(n13614), .B2(n13613), .A(n13612), .ZN(n13628) );
  OR2_X1 U15867 ( .A1(n13616), .A2(n13615), .ZN(n13619) );
  NAND2_X1 U15868 ( .A1(n13633), .A2(n13617), .ZN(n13618) );
  AND2_X1 U15869 ( .A1(n13619), .A2(n13618), .ZN(n13774) );
  OAI22_X1 U15870 ( .A1(n13774), .A2(n13621), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13620), .ZN(n13622) );
  AOI21_X1 U15871 ( .B1(n13779), .B2(n13623), .A(n13622), .ZN(n13626) );
  NAND2_X1 U15872 ( .A1(n13778), .A2(n13624), .ZN(n13625) );
  OAI211_X1 U15873 ( .C1(n13628), .C2(n13627), .A(n13626), .B(n13625), .ZN(
        P2_U3212) );
  INV_X2 U15874 ( .A(P2_U3947), .ZN(n13657) );
  MUX2_X1 U15875 ( .A(n13725), .B(P2_DATAO_REG_31__SCAN_IN), .S(n13657), .Z(
        P2_U3562) );
  MUX2_X1 U15876 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n13629), .S(P2_U3947), .Z(
        P2_U3561) );
  MUX2_X1 U15877 ( .A(n13630), .B(P2_DATAO_REG_29__SCAN_IN), .S(n13657), .Z(
        P2_U3560) );
  MUX2_X1 U15878 ( .A(n8388), .B(P2_DATAO_REG_28__SCAN_IN), .S(n13657), .Z(
        P2_U3559) );
  MUX2_X1 U15879 ( .A(n13631), .B(P2_DATAO_REG_27__SCAN_IN), .S(n13657), .Z(
        P2_U3558) );
  MUX2_X1 U15880 ( .A(n13632), .B(P2_DATAO_REG_26__SCAN_IN), .S(n13657), .Z(
        P2_U3557) );
  MUX2_X1 U15881 ( .A(n13633), .B(P2_DATAO_REG_25__SCAN_IN), .S(n13657), .Z(
        P2_U3556) );
  MUX2_X1 U15882 ( .A(n13634), .B(P2_DATAO_REG_24__SCAN_IN), .S(n13657), .Z(
        P2_U3555) );
  MUX2_X1 U15883 ( .A(n13635), .B(P2_DATAO_REG_23__SCAN_IN), .S(n13657), .Z(
        P2_U3554) );
  MUX2_X1 U15884 ( .A(n13636), .B(P2_DATAO_REG_22__SCAN_IN), .S(n13657), .Z(
        P2_U3553) );
  MUX2_X1 U15885 ( .A(n13637), .B(P2_DATAO_REG_21__SCAN_IN), .S(n13657), .Z(
        P2_U3552) );
  MUX2_X1 U15886 ( .A(n13638), .B(P2_DATAO_REG_20__SCAN_IN), .S(n13657), .Z(
        P2_U3551) );
  MUX2_X1 U15887 ( .A(n13639), .B(P2_DATAO_REG_19__SCAN_IN), .S(n13657), .Z(
        P2_U3550) );
  MUX2_X1 U15888 ( .A(n13640), .B(P2_DATAO_REG_18__SCAN_IN), .S(n13657), .Z(
        P2_U3549) );
  MUX2_X1 U15889 ( .A(n13641), .B(P2_DATAO_REG_17__SCAN_IN), .S(n13657), .Z(
        P2_U3548) );
  MUX2_X1 U15890 ( .A(n13642), .B(P2_DATAO_REG_16__SCAN_IN), .S(n13657), .Z(
        P2_U3547) );
  MUX2_X1 U15891 ( .A(n13643), .B(P2_DATAO_REG_15__SCAN_IN), .S(n13657), .Z(
        P2_U3546) );
  MUX2_X1 U15892 ( .A(n13644), .B(P2_DATAO_REG_14__SCAN_IN), .S(n13657), .Z(
        P2_U3545) );
  MUX2_X1 U15893 ( .A(n13645), .B(P2_DATAO_REG_13__SCAN_IN), .S(n13657), .Z(
        P2_U3544) );
  MUX2_X1 U15894 ( .A(n13646), .B(P2_DATAO_REG_12__SCAN_IN), .S(n13657), .Z(
        P2_U3543) );
  MUX2_X1 U15895 ( .A(n13647), .B(P2_DATAO_REG_11__SCAN_IN), .S(n13657), .Z(
        P2_U3542) );
  MUX2_X1 U15896 ( .A(n13648), .B(P2_DATAO_REG_10__SCAN_IN), .S(n13657), .Z(
        P2_U3541) );
  MUX2_X1 U15897 ( .A(n13649), .B(P2_DATAO_REG_9__SCAN_IN), .S(n13657), .Z(
        P2_U3540) );
  MUX2_X1 U15898 ( .A(n13650), .B(P2_DATAO_REG_8__SCAN_IN), .S(n13657), .Z(
        P2_U3539) );
  MUX2_X1 U15899 ( .A(n13651), .B(P2_DATAO_REG_7__SCAN_IN), .S(n13657), .Z(
        P2_U3538) );
  MUX2_X1 U15900 ( .A(n13652), .B(P2_DATAO_REG_6__SCAN_IN), .S(n13657), .Z(
        P2_U3537) );
  MUX2_X1 U15901 ( .A(n13653), .B(P2_DATAO_REG_5__SCAN_IN), .S(n13657), .Z(
        P2_U3536) );
  MUX2_X1 U15902 ( .A(n13654), .B(P2_DATAO_REG_4__SCAN_IN), .S(n13657), .Z(
        P2_U3535) );
  MUX2_X1 U15903 ( .A(n13655), .B(P2_DATAO_REG_3__SCAN_IN), .S(n13657), .Z(
        P2_U3534) );
  MUX2_X1 U15904 ( .A(n13656), .B(P2_DATAO_REG_2__SCAN_IN), .S(n13657), .Z(
        P2_U3533) );
  MUX2_X1 U15905 ( .A(n13658), .B(P2_DATAO_REG_1__SCAN_IN), .S(n13657), .Z(
        P2_U3532) );
  OR2_X1 U15906 ( .A1(n13665), .A2(n10712), .ZN(n13660) );
  AOI211_X1 U15907 ( .C1(n13661), .C2(n13660), .A(n13659), .B(n15407), .ZN(
        n13662) );
  AOI21_X1 U15908 ( .B1(n15453), .B2(n13663), .A(n13662), .ZN(n13670) );
  AOI22_X1 U15909 ( .A1(n15448), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3088), .ZN(n13669) );
  INV_X1 U15910 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n15525) );
  MUX2_X1 U15911 ( .A(n10510), .B(P2_REG1_REG_1__SCAN_IN), .S(n13663), .Z(
        n13664) );
  OAI21_X1 U15912 ( .B1(n15525), .B2(n13665), .A(n13664), .ZN(n13666) );
  NAND3_X1 U15913 ( .A1(n15456), .A2(n13667), .A3(n13666), .ZN(n13668) );
  NAND3_X1 U15914 ( .A1(n13670), .A2(n13669), .A3(n13668), .ZN(P2_U3215) );
  NAND2_X1 U15915 ( .A1(n15454), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n13681) );
  MUX2_X1 U15916 ( .A(n8062), .B(P2_REG2_REG_17__SCAN_IN), .S(n15454), .Z(
        n13671) );
  INV_X1 U15917 ( .A(n13671), .ZN(n15451) );
  NAND2_X1 U15918 ( .A1(n15436), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n13680) );
  MUX2_X1 U15919 ( .A(n12393), .B(P2_REG2_REG_16__SCAN_IN), .S(n15436), .Z(
        n13672) );
  INV_X1 U15920 ( .A(n13672), .ZN(n15438) );
  OAI21_X1 U15921 ( .B1(n13674), .B2(P2_REG2_REG_12__SCAN_IN), .A(n13673), 
        .ZN(n15409) );
  MUX2_X1 U15922 ( .A(n13675), .B(P2_REG2_REG_13__SCAN_IN), .S(n13689), .Z(
        n15408) );
  NAND2_X1 U15923 ( .A1(n15417), .A2(n13676), .ZN(n13677) );
  XNOR2_X1 U15924 ( .A(n13676), .B(n13691), .ZN(n15416) );
  NAND2_X1 U15925 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n15416), .ZN(n15415) );
  NAND2_X1 U15926 ( .A1(n13677), .A2(n15415), .ZN(n13678) );
  NAND2_X1 U15927 ( .A1(n15426), .A2(n13678), .ZN(n13679) );
  XOR2_X1 U15928 ( .A(n15426), .B(n13678), .Z(n15428) );
  NAND2_X1 U15929 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n15428), .ZN(n15427) );
  NAND2_X1 U15930 ( .A1(n13679), .A2(n15427), .ZN(n15439) );
  NAND2_X1 U15931 ( .A1(n15451), .A2(n15452), .ZN(n15449) );
  NAND2_X1 U15932 ( .A1(n13681), .A2(n15449), .ZN(n13705) );
  XNOR2_X1 U15933 ( .A(n13710), .B(n13705), .ZN(n13682) );
  NOR2_X1 U15934 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n13682), .ZN(n13707) );
  AOI21_X1 U15935 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n13682), .A(n13707), 
        .ZN(n13683) );
  OR2_X1 U15936 ( .A1(n13683), .A2(n15407), .ZN(n13704) );
  INV_X1 U15937 ( .A(n13684), .ZN(n13685) );
  AOI21_X1 U15938 ( .B1(n15448), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n13685), 
        .ZN(n13703) );
  NAND2_X1 U15939 ( .A1(n15453), .A2(n13710), .ZN(n13702) );
  XNOR2_X1 U15940 ( .A(n15454), .B(n14007), .ZN(n15458) );
  INV_X1 U15941 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n14014) );
  XNOR2_X1 U15942 ( .A(n15436), .B(n14014), .ZN(n15441) );
  AOI21_X1 U15943 ( .B1(n13688), .B2(n13687), .A(n13686), .ZN(n15406) );
  MUX2_X1 U15944 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n13690), .S(n13689), .Z(
        n15405) );
  NAND2_X1 U15945 ( .A1(n15406), .A2(n15405), .ZN(n15404) );
  OAI21_X1 U15946 ( .B1(n13690), .B2(n15400), .A(n15404), .ZN(n15420) );
  XNOR2_X1 U15947 ( .A(n13691), .B(P2_REG1_REG_14__SCAN_IN), .ZN(n15419) );
  NAND2_X1 U15948 ( .A1(n15420), .A2(n15419), .ZN(n15418) );
  OAI21_X1 U15949 ( .B1(n13692), .B2(n13691), .A(n15418), .ZN(n13693) );
  NAND2_X1 U15950 ( .A1(n15426), .A2(n13693), .ZN(n13695) );
  XNOR2_X1 U15951 ( .A(n13694), .B(n13693), .ZN(n15430) );
  NAND2_X1 U15952 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n15430), .ZN(n15429) );
  NAND2_X1 U15953 ( .A1(n13695), .A2(n15429), .ZN(n15442) );
  NAND2_X1 U15954 ( .A1(n15441), .A2(n15442), .ZN(n15440) );
  OAI21_X1 U15955 ( .B1(n13696), .B2(n14014), .A(n15440), .ZN(n15457) );
  NAND2_X1 U15956 ( .A1(n15458), .A2(n15457), .ZN(n15455) );
  OAI21_X1 U15957 ( .B1(n14007), .B2(n13697), .A(n15455), .ZN(n13709) );
  XNOR2_X1 U15958 ( .A(n13710), .B(n13709), .ZN(n13698) );
  INV_X1 U15959 ( .A(n13698), .ZN(n13700) );
  OAI211_X1 U15960 ( .C1(P2_REG1_REG_18__SCAN_IN), .C2(n13700), .A(n15456), 
        .B(n13711), .ZN(n13701) );
  NAND4_X1 U15961 ( .A1(n13704), .A2(n13703), .A3(n13702), .A4(n13701), .ZN(
        P2_U3232) );
  NOR2_X1 U15962 ( .A1(n13710), .A2(n13705), .ZN(n13706) );
  XOR2_X1 U15963 ( .A(n13708), .B(P2_REG2_REG_19__SCAN_IN), .Z(n13717) );
  INV_X1 U15964 ( .A(n13717), .ZN(n13715) );
  NAND2_X1 U15965 ( .A1(n13710), .A2(n13709), .ZN(n13712) );
  NAND2_X1 U15966 ( .A1(n13712), .A2(n13711), .ZN(n13713) );
  XOR2_X1 U15967 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n13713), .Z(n13716) );
  NOR2_X1 U15968 ( .A1(n13716), .A2(n15375), .ZN(n13714) );
  AOI22_X1 U15969 ( .A1(n13717), .A2(n15450), .B1(n15456), .B2(n13716), .ZN(
        n13719) );
  OAI211_X1 U15970 ( .C1(n7716), .C2(n13722), .A(n13721), .B(n13720), .ZN(
        P2_U3233) );
  NAND2_X1 U15971 ( .A1(n13732), .A2(n14029), .ZN(n13731) );
  NOR2_X1 U15972 ( .A1(n13919), .A2(n13724), .ZN(n13728) );
  INV_X1 U15973 ( .A(n13725), .ZN(n13726) );
  OR2_X1 U15974 ( .A1(n13727), .A2(n13726), .ZN(n13942) );
  NOR2_X1 U15975 ( .A1(n13926), .A2(n13942), .ZN(n13734) );
  AOI211_X1 U15976 ( .C1(n13729), .C2(n13933), .A(n13728), .B(n13734), .ZN(
        n13730) );
  OAI21_X1 U15977 ( .B1(n13939), .B2(n13922), .A(n13730), .ZN(P2_U3234) );
  OAI211_X1 U15978 ( .C1(n13732), .C2(n14029), .A(n11777), .B(n13731), .ZN(
        n13943) );
  NOR2_X1 U15979 ( .A1(n13919), .A2(n13733), .ZN(n13735) );
  AOI211_X1 U15980 ( .C1(n13736), .C2(n13933), .A(n13735), .B(n13734), .ZN(
        n13737) );
  OAI21_X1 U15981 ( .B1(n13943), .B2(n13922), .A(n13737), .ZN(P2_U3235) );
  NAND2_X1 U15982 ( .A1(n13738), .A2(n13924), .ZN(n13746) );
  OAI22_X1 U15983 ( .A1(n13740), .A2(n13916), .B1(n13739), .B2(n13919), .ZN(
        n13743) );
  NOR2_X1 U15984 ( .A1(n13741), .A2(n13922), .ZN(n13742) );
  AOI211_X1 U15985 ( .C1(n13933), .C2(n13744), .A(n13743), .B(n13742), .ZN(
        n13745) );
  OAI211_X1 U15986 ( .C1(n13747), .C2(n13926), .A(n13746), .B(n13745), .ZN(
        P2_U3236) );
  OAI22_X1 U15987 ( .A1(n14032), .A2(n13824), .B1(n13748), .B2(n13919), .ZN(
        n13749) );
  AOI21_X1 U15988 ( .B1(n7689), .B2(n13930), .A(n13749), .ZN(n13754) );
  NOR2_X1 U15989 ( .A1(n13750), .A2(n13916), .ZN(n13751) );
  OAI21_X1 U15990 ( .B1(n13752), .B2(n13751), .A(n13919), .ZN(n13753) );
  OAI211_X1 U15991 ( .C1(n13755), .C2(n13902), .A(n13754), .B(n13753), .ZN(
        P2_U3237) );
  XNOR2_X1 U15992 ( .A(n13756), .B(n13760), .ZN(n13759) );
  INV_X1 U15993 ( .A(n13757), .ZN(n13758) );
  AOI21_X1 U15994 ( .B1(n13759), .B2(n13906), .A(n13758), .ZN(n13951) );
  NAND2_X1 U15995 ( .A1(n13761), .A2(n13760), .ZN(n13946) );
  NAND3_X1 U15996 ( .A1(n13947), .A2(n13946), .A3(n13924), .ZN(n13770) );
  NOR2_X1 U15997 ( .A1(n13766), .A2(n13776), .ZN(n13762) );
  INV_X1 U15998 ( .A(n13950), .ZN(n13768) );
  AOI22_X1 U15999 ( .A1(n13764), .A2(n13931), .B1(P2_REG2_REG_27__SCAN_IN), 
        .B2(n13926), .ZN(n13765) );
  OAI21_X1 U16000 ( .B1(n13766), .B2(n13824), .A(n13765), .ZN(n13767) );
  AOI21_X1 U16001 ( .B1(n13768), .B2(n13930), .A(n13767), .ZN(n13769) );
  OAI211_X1 U16002 ( .C1(n13951), .C2(n13926), .A(n13770), .B(n13769), .ZN(
        P2_U3238) );
  XNOR2_X1 U16003 ( .A(n13771), .B(n13772), .ZN(n13955) );
  INV_X1 U16004 ( .A(n13955), .ZN(n13784) );
  XNOR2_X1 U16005 ( .A(n13773), .B(n13772), .ZN(n13775) );
  OAI21_X1 U16006 ( .B1(n13775), .B2(n13896), .A(n13774), .ZN(n13953) );
  INV_X1 U16007 ( .A(n13792), .ZN(n13777) );
  AOI211_X1 U16008 ( .C1(n13778), .C2(n13777), .A(n13912), .B(n13776), .ZN(
        n13954) );
  NAND2_X1 U16009 ( .A1(n13954), .A2(n13930), .ZN(n13781) );
  AOI22_X1 U16010 ( .A1(n13779), .A2(n13931), .B1(P2_REG2_REG_26__SCAN_IN), 
        .B2(n13926), .ZN(n13780) );
  OAI211_X1 U16011 ( .C1(n14037), .C2(n13824), .A(n13781), .B(n13780), .ZN(
        n13782) );
  AOI21_X1 U16012 ( .B1(n13919), .B2(n13953), .A(n13782), .ZN(n13783) );
  OAI21_X1 U16013 ( .B1(n13784), .B2(n13902), .A(n13783), .ZN(P2_U3239) );
  NAND3_X1 U16014 ( .A1(n13802), .A2(n7321), .A3(n13785), .ZN(n13786) );
  AOI21_X1 U16015 ( .B1(n13787), .B2(n13786), .A(n13896), .ZN(n13789) );
  INV_X1 U16016 ( .A(n13959), .ZN(n13801) );
  OAI21_X1 U16017 ( .B1(n13791), .B2(n7321), .A(n13790), .ZN(n13961) );
  NOR2_X1 U16018 ( .A1(n13812), .A2(n14041), .ZN(n13793) );
  OAI22_X1 U16019 ( .A1(n13795), .A2(n13916), .B1(n13919), .B2(n13794), .ZN(
        n13796) );
  AOI21_X1 U16020 ( .B1(n13797), .B2(n13933), .A(n13796), .ZN(n13798) );
  OAI21_X1 U16021 ( .B1(n13958), .B2(n13922), .A(n13798), .ZN(n13799) );
  AOI21_X1 U16022 ( .B1(n13961), .B2(n13924), .A(n13799), .ZN(n13800) );
  OAI21_X1 U16023 ( .B1(n13926), .B2(n13801), .A(n13800), .ZN(P2_U3240) );
  OAI21_X1 U16024 ( .B1(n13804), .B2(n13803), .A(n13802), .ZN(n13807) );
  INV_X1 U16025 ( .A(n13805), .ZN(n13806) );
  AOI21_X1 U16026 ( .B1(n13807), .B2(n13906), .A(n13806), .ZN(n13967) );
  OAI21_X1 U16027 ( .B1(n7691), .B2(n13809), .A(n13808), .ZN(n13968) );
  INV_X1 U16028 ( .A(n13968), .ZN(n13817) );
  NAND2_X1 U16029 ( .A1(n13822), .A2(n13965), .ZN(n13810) );
  NAND2_X1 U16030 ( .A1(n13810), .A2(n11777), .ZN(n13811) );
  NOR2_X1 U16031 ( .A1(n13812), .A2(n13811), .ZN(n13964) );
  NAND2_X1 U16032 ( .A1(n13964), .A2(n13930), .ZN(n13815) );
  AOI22_X1 U16033 ( .A1(n13926), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n13813), 
        .B2(n13931), .ZN(n13814) );
  OAI211_X1 U16034 ( .C1(n7164), .C2(n13824), .A(n13815), .B(n13814), .ZN(
        n13816) );
  AOI21_X1 U16035 ( .B1(n13817), .B2(n13924), .A(n13816), .ZN(n13818) );
  OAI21_X1 U16036 ( .B1(n13926), .B2(n13967), .A(n13818), .ZN(P2_U3241) );
  INV_X1 U16037 ( .A(n13819), .ZN(n13820) );
  AOI21_X1 U16038 ( .B1(n13828), .B2(n13821), .A(n13820), .ZN(n13973) );
  AOI211_X1 U16039 ( .C1(n13970), .C2(n13841), .A(n8410), .B(n7166), .ZN(
        n13969) );
  OAI22_X1 U16040 ( .A1(n7165), .A2(n13824), .B1(n13919), .B2(n13823), .ZN(
        n13825) );
  AOI21_X1 U16041 ( .B1(n13969), .B2(n13930), .A(n13825), .ZN(n13835) );
  AND2_X1 U16042 ( .A1(n13838), .A2(n13826), .ZN(n13829) );
  OAI21_X1 U16043 ( .B1(n13829), .B2(n13828), .A(n13827), .ZN(n13831) );
  AOI21_X1 U16044 ( .B1(n13831), .B2(n13906), .A(n13830), .ZN(n13972) );
  OAI21_X1 U16045 ( .B1(n13832), .B2(n13916), .A(n13972), .ZN(n13833) );
  NAND2_X1 U16046 ( .A1(n13833), .A2(n13919), .ZN(n13834) );
  OAI211_X1 U16047 ( .C1(n13973), .C2(n13902), .A(n13835), .B(n13834), .ZN(
        P2_U3242) );
  NAND2_X1 U16048 ( .A1(n13848), .A2(n13836), .ZN(n13837) );
  NAND3_X1 U16049 ( .A1(n13838), .A2(n13906), .A3(n13837), .ZN(n13840) );
  AOI21_X1 U16050 ( .B1(n13975), .B2(n13854), .A(n13912), .ZN(n13842) );
  AND2_X1 U16051 ( .A1(n13842), .A2(n13841), .ZN(n13974) );
  NAND2_X1 U16052 ( .A1(n13975), .A2(n13933), .ZN(n13845) );
  NAND2_X1 U16053 ( .A1(n13931), .A2(n13843), .ZN(n13844) );
  OAI211_X1 U16054 ( .C1(n13919), .C2(n13846), .A(n13845), .B(n13844), .ZN(
        n13851) );
  OAI21_X1 U16055 ( .B1(n13849), .B2(n13848), .A(n13847), .ZN(n13978) );
  NOR2_X1 U16056 ( .A1(n13978), .A2(n13902), .ZN(n13850) );
  AOI211_X1 U16057 ( .C1(n13974), .C2(n13930), .A(n13851), .B(n13850), .ZN(
        n13852) );
  OAI21_X1 U16058 ( .B1(n13926), .B2(n13977), .A(n13852), .ZN(P2_U3243) );
  XNOR2_X1 U16059 ( .A(n13853), .B(n13861), .ZN(n13979) );
  OAI211_X1 U16060 ( .C1(n13882), .C2(n14048), .A(n11777), .B(n13854), .ZN(
        n13980) );
  INV_X1 U16061 ( .A(n13855), .ZN(n13856) );
  OAI22_X1 U16062 ( .A1(n13919), .A2(n13857), .B1(n13856), .B2(n13916), .ZN(
        n13858) );
  AOI21_X1 U16063 ( .B1(n13859), .B2(n13933), .A(n13858), .ZN(n13860) );
  OAI21_X1 U16064 ( .B1(n13980), .B2(n13922), .A(n13860), .ZN(n13869) );
  OR2_X1 U16065 ( .A1(n13862), .A2(n13861), .ZN(n13863) );
  NAND2_X1 U16066 ( .A1(n13864), .A2(n13863), .ZN(n13867) );
  INV_X1 U16067 ( .A(n13865), .ZN(n13866) );
  AOI21_X1 U16068 ( .B1(n13867), .B2(n13906), .A(n13866), .ZN(n13981) );
  NOR2_X1 U16069 ( .A1(n13981), .A2(n13926), .ZN(n13868) );
  AOI211_X1 U16070 ( .C1(n13924), .C2(n13979), .A(n13869), .B(n13868), .ZN(
        n13870) );
  INV_X1 U16071 ( .A(n13870), .ZN(P2_U3244) );
  XNOR2_X1 U16072 ( .A(n13871), .B(n13874), .ZN(n13989) );
  OAI21_X1 U16073 ( .B1(n13874), .B2(n13873), .A(n13872), .ZN(n13876) );
  AOI21_X1 U16074 ( .B1(n13876), .B2(n13906), .A(n13875), .ZN(n13988) );
  OAI22_X1 U16075 ( .A1(n13919), .A2(n13878), .B1(n13877), .B2(n13916), .ZN(
        n13879) );
  AOI21_X1 U16076 ( .B1(n13986), .B2(n13933), .A(n13879), .ZN(n13884) );
  NAND2_X1 U16077 ( .A1(n6694), .A2(n13986), .ZN(n13880) );
  NAND2_X1 U16078 ( .A1(n13880), .A2(n11777), .ZN(n13881) );
  NOR2_X1 U16079 ( .A1(n13882), .A2(n13881), .ZN(n13985) );
  NAND2_X1 U16080 ( .A1(n13985), .A2(n13930), .ZN(n13883) );
  OAI211_X1 U16081 ( .C1(n13988), .C2(n13926), .A(n13884), .B(n13883), .ZN(
        n13885) );
  INV_X1 U16082 ( .A(n13885), .ZN(n13886) );
  OAI21_X1 U16083 ( .B1(n13989), .B2(n13902), .A(n13886), .ZN(P2_U3245) );
  XNOR2_X1 U16084 ( .A(n13887), .B(n13895), .ZN(n13995) );
  INV_X1 U16085 ( .A(n13995), .ZN(n13903) );
  OAI22_X1 U16086 ( .A1(n13919), .A2(n13889), .B1(n13888), .B2(n13916), .ZN(
        n13892) );
  AOI21_X1 U16087 ( .B1(n13893), .B2(n13914), .A(n13912), .ZN(n13890) );
  NAND2_X1 U16088 ( .A1(n13890), .A2(n6694), .ZN(n13991) );
  NOR2_X1 U16089 ( .A1(n13991), .A2(n13922), .ZN(n13891) );
  AOI211_X1 U16090 ( .C1(n13933), .C2(n13893), .A(n13892), .B(n13891), .ZN(
        n13901) );
  NAND2_X1 U16091 ( .A1(n13895), .A2(n13894), .ZN(n13897) );
  AOI21_X1 U16092 ( .B1(n13898), .B2(n13897), .A(n13896), .ZN(n13993) );
  INV_X1 U16093 ( .A(n13990), .ZN(n13899) );
  OAI21_X1 U16094 ( .B1(n13993), .B2(n13899), .A(n13919), .ZN(n13900) );
  OAI211_X1 U16095 ( .C1(n13903), .C2(n13902), .A(n13901), .B(n13900), .ZN(
        P2_U3246) );
  XNOR2_X1 U16096 ( .A(n13904), .B(n6793), .ZN(n13907) );
  AOI21_X1 U16097 ( .B1(n13907), .B2(n13906), .A(n13905), .ZN(n14000) );
  NAND2_X1 U16098 ( .A1(n13909), .A2(n13908), .ZN(n13910) );
  NAND2_X1 U16099 ( .A1(n13911), .A2(n13910), .ZN(n13997) );
  AOI21_X1 U16100 ( .B1(n14053), .B2(n13913), .A(n13912), .ZN(n13915) );
  NAND2_X1 U16101 ( .A1(n13915), .A2(n13914), .ZN(n13998) );
  OAI22_X1 U16102 ( .A1(n13919), .A2(n13918), .B1(n13917), .B2(n13916), .ZN(
        n13920) );
  AOI21_X1 U16103 ( .B1(n14053), .B2(n13933), .A(n13920), .ZN(n13921) );
  OAI21_X1 U16104 ( .B1(n13998), .B2(n13922), .A(n13921), .ZN(n13923) );
  AOI21_X1 U16105 ( .B1(n13997), .B2(n13924), .A(n13923), .ZN(n13925) );
  OAI21_X1 U16106 ( .B1(n14000), .B2(n13926), .A(n13925), .ZN(P2_U3247) );
  AOI22_X1 U16107 ( .A1(n13930), .A2(n13929), .B1(n13928), .B2(n13927), .ZN(
        n13938) );
  AOI22_X1 U16108 ( .A1(n13933), .A2(n13932), .B1(n13931), .B2(
        P2_REG3_REG_1__SCAN_IN), .ZN(n13937) );
  MUX2_X1 U16109 ( .A(n13935), .B(n13934), .S(n13919), .Z(n13936) );
  NAND3_X1 U16110 ( .A1(n13938), .A2(n13937), .A3(n13936), .ZN(P2_U3264) );
  INV_X1 U16111 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n13940) );
  OAI21_X1 U16112 ( .B1(n14025), .B2(n14016), .A(n13941), .ZN(P2_U3530) );
  AND2_X1 U16113 ( .A1(n13943), .A2(n13942), .ZN(n14026) );
  MUX2_X1 U16114 ( .A(n13944), .B(n14026), .S(n15539), .Z(n13945) );
  OAI21_X1 U16115 ( .B1(n14029), .B2(n14016), .A(n13945), .ZN(P2_U3529) );
  NAND3_X1 U16116 ( .A1(n13947), .A2(n15491), .A3(n13946), .ZN(n13952) );
  NAND2_X1 U16117 ( .A1(n13948), .A2(n15508), .ZN(n13949) );
  NAND4_X1 U16118 ( .A1(n13952), .A2(n13951), .A3(n13950), .A4(n13949), .ZN(
        n14033) );
  MUX2_X1 U16119 ( .A(n14033), .B(P2_REG1_REG_27__SCAN_IN), .S(n15536), .Z(
        P2_U3526) );
  INV_X1 U16120 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n13956) );
  AOI211_X1 U16121 ( .C1(n15491), .C2(n13955), .A(n13954), .B(n13953), .ZN(
        n14034) );
  MUX2_X1 U16122 ( .A(n13956), .B(n14034), .S(n15539), .Z(n13957) );
  OAI21_X1 U16123 ( .B1(n14037), .B2(n14016), .A(n13957), .ZN(P2_U3525) );
  INV_X1 U16124 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n13962) );
  INV_X1 U16125 ( .A(n13958), .ZN(n13960) );
  AOI211_X1 U16126 ( .C1(n13961), .C2(n15491), .A(n13960), .B(n13959), .ZN(
        n14038) );
  MUX2_X1 U16127 ( .A(n13962), .B(n14038), .S(n15539), .Z(n13963) );
  OAI21_X1 U16128 ( .B1(n14041), .B2(n14016), .A(n13963), .ZN(P2_U3524) );
  AOI21_X1 U16129 ( .B1(n15508), .B2(n13965), .A(n13964), .ZN(n13966) );
  OAI211_X1 U16130 ( .C1(n13968), .C2(n14022), .A(n13967), .B(n13966), .ZN(
        n14042) );
  MUX2_X1 U16131 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n14042), .S(n15539), .Z(
        P2_U3523) );
  AOI21_X1 U16132 ( .B1(n15508), .B2(n13970), .A(n13969), .ZN(n13971) );
  OAI211_X1 U16133 ( .C1(n13973), .C2(n14022), .A(n13972), .B(n13971), .ZN(
        n14043) );
  MUX2_X1 U16134 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n14043), .S(n15539), .Z(
        P2_U3522) );
  AOI21_X1 U16135 ( .B1(n15508), .B2(n13975), .A(n13974), .ZN(n13976) );
  OAI211_X1 U16136 ( .C1(n13978), .C2(n14022), .A(n13977), .B(n13976), .ZN(
        n14044) );
  MUX2_X1 U16137 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n14044), .S(n15539), .Z(
        P2_U3521) );
  NAND2_X1 U16138 ( .A1(n13979), .A2(n15491), .ZN(n13982) );
  NAND3_X1 U16139 ( .A1(n13982), .A2(n13981), .A3(n13980), .ZN(n14045) );
  MUX2_X1 U16140 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n14045), .S(n15539), .Z(
        n13983) );
  INV_X1 U16141 ( .A(n13983), .ZN(n13984) );
  OAI21_X1 U16142 ( .B1(n14048), .B2(n14016), .A(n13984), .ZN(P2_U3520) );
  AOI21_X1 U16143 ( .B1(n15508), .B2(n13986), .A(n13985), .ZN(n13987) );
  OAI211_X1 U16144 ( .C1(n13989), .C2(n14022), .A(n13988), .B(n13987), .ZN(
        n14049) );
  MUX2_X1 U16145 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n14049), .S(n15539), .Z(
        P2_U3519) );
  OAI211_X1 U16146 ( .C1(n13992), .C2(n15516), .A(n13991), .B(n13990), .ZN(
        n13994) );
  AOI211_X1 U16147 ( .C1(n15491), .C2(n13995), .A(n13994), .B(n13993), .ZN(
        n13996) );
  INV_X1 U16148 ( .A(n13996), .ZN(n14050) );
  MUX2_X1 U16149 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n14050), .S(n15539), .Z(
        P2_U3518) );
  NAND2_X1 U16150 ( .A1(n13997), .A2(n15491), .ZN(n13999) );
  NAND3_X1 U16151 ( .A1(n14000), .A2(n13999), .A3(n13998), .ZN(n14051) );
  MUX2_X1 U16152 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n14051), .S(n15539), .Z(
        n14001) );
  AOI21_X1 U16153 ( .B1(n14002), .B2(n14053), .A(n14001), .ZN(n14003) );
  INV_X1 U16154 ( .A(n14003), .ZN(P2_U3517) );
  AOI211_X1 U16155 ( .C1(n15491), .C2(n14006), .A(n14005), .B(n14004), .ZN(
        n14055) );
  MUX2_X1 U16156 ( .A(n14007), .B(n14055), .S(n15539), .Z(n14008) );
  OAI21_X1 U16157 ( .B1(n14058), .B2(n14016), .A(n14008), .ZN(P2_U3516) );
  NAND3_X1 U16158 ( .A1(n14011), .A2(n14010), .A3(n14009), .ZN(n14012) );
  AOI21_X1 U16159 ( .B1(n14013), .B2(n15491), .A(n14012), .ZN(n14059) );
  MUX2_X1 U16160 ( .A(n14014), .B(n14059), .S(n15539), .Z(n14015) );
  OAI21_X1 U16161 ( .B1(n14063), .B2(n14016), .A(n14015), .ZN(P2_U3515) );
  AOI211_X1 U16162 ( .C1(n15508), .C2(n14019), .A(n14018), .B(n14017), .ZN(
        n14020) );
  OAI21_X1 U16163 ( .B1(n14022), .B2(n14021), .A(n14020), .ZN(n14064) );
  MUX2_X1 U16164 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n14064), .S(n15539), .Z(
        P2_U3511) );
  INV_X1 U16165 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n14024) );
  MUX2_X1 U16166 ( .A(n14027), .B(n14026), .S(n15524), .Z(n14028) );
  OAI21_X1 U16167 ( .B1(n14029), .B2(n14062), .A(n14028), .ZN(P2_U3497) );
  OAI21_X1 U16168 ( .B1(n14032), .B2(n14062), .A(n14031), .ZN(P2_U3495) );
  MUX2_X1 U16169 ( .A(n14033), .B(P2_REG0_REG_27__SCAN_IN), .S(n15523), .Z(
        P2_U3494) );
  INV_X1 U16170 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n14035) );
  MUX2_X1 U16171 ( .A(n14035), .B(n14034), .S(n15524), .Z(n14036) );
  OAI21_X1 U16172 ( .B1(n14037), .B2(n14062), .A(n14036), .ZN(P2_U3493) );
  INV_X1 U16173 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n14039) );
  MUX2_X1 U16174 ( .A(n14039), .B(n14038), .S(n15524), .Z(n14040) );
  OAI21_X1 U16175 ( .B1(n14041), .B2(n14062), .A(n14040), .ZN(P2_U3492) );
  MUX2_X1 U16176 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n14042), .S(n15524), .Z(
        P2_U3491) );
  MUX2_X1 U16177 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n14043), .S(n15524), .Z(
        P2_U3490) );
  MUX2_X1 U16178 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n14044), .S(n15524), .Z(
        P2_U3489) );
  MUX2_X1 U16179 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n14045), .S(n15524), .Z(
        n14046) );
  INV_X1 U16180 ( .A(n14046), .ZN(n14047) );
  OAI21_X1 U16181 ( .B1(n14048), .B2(n14062), .A(n14047), .ZN(P2_U3488) );
  MUX2_X1 U16182 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n14049), .S(n15524), .Z(
        P2_U3487) );
  MUX2_X1 U16183 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n14050), .S(n15524), .Z(
        P2_U3486) );
  MUX2_X1 U16184 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n14051), .S(n15524), .Z(
        n14052) );
  AOI21_X1 U16185 ( .B1(n8423), .B2(n14053), .A(n14052), .ZN(n14054) );
  INV_X1 U16186 ( .A(n14054), .ZN(P2_U3484) );
  INV_X1 U16187 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n14056) );
  MUX2_X1 U16188 ( .A(n14056), .B(n14055), .S(n15524), .Z(n14057) );
  OAI21_X1 U16189 ( .B1(n14058), .B2(n14062), .A(n14057), .ZN(P2_U3481) );
  INV_X1 U16190 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n14060) );
  MUX2_X1 U16191 ( .A(n14060), .B(n14059), .S(n15524), .Z(n14061) );
  OAI21_X1 U16192 ( .B1(n14063), .B2(n14062), .A(n14061), .ZN(P2_U3478) );
  MUX2_X1 U16193 ( .A(P2_REG0_REG_12__SCAN_IN), .B(n14064), .S(n15524), .Z(
        P2_U3466) );
  INV_X1 U16194 ( .A(n14875), .ZN(n14068) );
  NOR4_X1 U16195 ( .A1(n7730), .A2(P2_IR_REG_30__SCAN_IN), .A3(n14065), .A4(
        P2_U3088), .ZN(n14066) );
  AOI21_X1 U16196 ( .B1(n14080), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n14066), 
        .ZN(n14067) );
  OAI21_X1 U16197 ( .B1(n14068), .B2(n14083), .A(n14067), .ZN(P2_U3296) );
  INV_X1 U16198 ( .A(n14372), .ZN(n14879) );
  OAI222_X1 U16199 ( .A1(n14075), .A2(n14879), .B1(P2_U3088), .B2(n14069), 
        .C1(n14070), .C2(n14072), .ZN(P2_U3297) );
  INV_X1 U16200 ( .A(n14071), .ZN(n14882) );
  INV_X1 U16201 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n14073) );
  OAI222_X1 U16202 ( .A1(n14075), .A2(n14882), .B1(P2_U3088), .B2(n14074), 
        .C1(n14073), .C2(n14072), .ZN(P2_U3298) );
  NAND2_X1 U16203 ( .A1(n14080), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n14076) );
  OAI211_X1 U16204 ( .C1(n14078), .C2(n14083), .A(n14077), .B(n14076), .ZN(
        P2_U3299) );
  INV_X1 U16205 ( .A(n14079), .ZN(n14884) );
  AOI22_X1 U16206 ( .A1(n14081), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_27__SCAN_IN), .B2(n14080), .ZN(n14082) );
  OAI21_X1 U16207 ( .B1(n14884), .B2(n14083), .A(n14082), .ZN(P2_U3300) );
  INV_X1 U16208 ( .A(n14084), .ZN(n14085) );
  MUX2_X1 U16209 ( .A(n14085), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  AOI22_X1 U16210 ( .A1(n14088), .A2(n14205), .B1(P1_REG3_REG_27__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14089) );
  OAI21_X1 U16211 ( .B1(n14666), .B2(n15086), .A(n14089), .ZN(n14090) );
  AOI21_X1 U16212 ( .B1(n14480), .B2(n15107), .A(n14090), .ZN(n14091) );
  OAI211_X1 U16213 ( .C1(n14093), .C2(n15111), .A(n14092), .B(n14091), .ZN(
        P1_U3214) );
  INV_X1 U16214 ( .A(n14812), .ZN(n14102) );
  INV_X1 U16215 ( .A(n14094), .ZN(n14172) );
  NOR3_X1 U16216 ( .A1(n14172), .A2(n7540), .A3(n14096), .ZN(n14097) );
  OAI21_X1 U16217 ( .B1(n14097), .B2(n6698), .A(n15114), .ZN(n14101) );
  OAI22_X1 U16218 ( .A1(n14665), .A2(n14947), .B1(n14344), .B2(n15131), .ZN(
        n14811) );
  OAI22_X1 U16219 ( .A1(n14699), .A2(n15119), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14098), .ZN(n14099) );
  AOI21_X1 U16220 ( .B1(n14811), .B2(n14195), .A(n14099), .ZN(n14100) );
  OAI211_X1 U16221 ( .C1(n14102), .C2(n15111), .A(n14101), .B(n14100), .ZN(
        P1_U3216) );
  INV_X1 U16222 ( .A(n14758), .ZN(n14838) );
  OAI21_X1 U16223 ( .B1(n6700), .B2(n14104), .A(n14103), .ZN(n14106) );
  NAND3_X1 U16224 ( .A1(n14106), .A2(n15114), .A3(n14105), .ZN(n14110) );
  NOR2_X1 U16225 ( .A1(n15119), .A2(n14764), .ZN(n14108) );
  INV_X1 U16226 ( .A(n15107), .ZN(n15088) );
  NAND2_X1 U16227 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n14622)
         );
  OAI21_X1 U16228 ( .B1(n15088), .B2(n14336), .A(n14622), .ZN(n14107) );
  AOI211_X1 U16229 ( .C1(n15109), .C2(n14761), .A(n14108), .B(n14107), .ZN(
        n14109) );
  OAI211_X1 U16230 ( .C1(n14838), .C2(n15111), .A(n14110), .B(n14109), .ZN(
        P1_U3219) );
  INV_X1 U16231 ( .A(n14111), .ZN(n14112) );
  AOI21_X1 U16232 ( .B1(n14114), .B2(n14113), .A(n14112), .ZN(n14118) );
  OAI22_X1 U16233 ( .A1(n14344), .A2(n14947), .B1(n14336), .B2(n15131), .ZN(
        n14724) );
  AOI22_X1 U16234 ( .A1(n14724), .A2(n14195), .B1(P1_REG3_REG_21__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14115) );
  OAI21_X1 U16235 ( .B1(n14730), .B2(n15119), .A(n14115), .ZN(n14116) );
  AOI21_X1 U16236 ( .B1(n14827), .B2(n15097), .A(n14116), .ZN(n14117) );
  OAI21_X1 U16237 ( .B1(n14118), .B2(n15092), .A(n14117), .ZN(P1_U3223) );
  INV_X1 U16238 ( .A(n14119), .ZN(n14153) );
  INV_X1 U16239 ( .A(n14120), .ZN(n14122) );
  NOR3_X1 U16240 ( .A1(n14153), .A2(n14122), .A3(n14121), .ZN(n14125) );
  INV_X1 U16241 ( .A(n14123), .ZN(n14124) );
  OAI21_X1 U16242 ( .B1(n14125), .B2(n14124), .A(n15114), .ZN(n14129) );
  AOI22_X1 U16243 ( .A1(n14484), .A2(n15109), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14126) );
  OAI21_X1 U16244 ( .B1(n14672), .B2(n15119), .A(n14126), .ZN(n14127) );
  AOI21_X1 U16245 ( .B1(n15107), .B2(n14482), .A(n14127), .ZN(n14128) );
  OAI211_X1 U16246 ( .C1(n14801), .C2(n15111), .A(n14129), .B(n14128), .ZN(
        P1_U3225) );
  INV_X1 U16247 ( .A(n14130), .ZN(n14131) );
  AOI21_X1 U16248 ( .B1(n14133), .B2(n14132), .A(n14131), .ZN(n14139) );
  NOR2_X1 U16249 ( .A1(n15119), .A2(n15137), .ZN(n14137) );
  NAND2_X1 U16250 ( .A1(n15107), .A2(n15135), .ZN(n14135) );
  OAI211_X1 U16251 ( .C1(n15132), .C2(n15086), .A(n14135), .B(n14134), .ZN(
        n14136) );
  AOI211_X1 U16252 ( .C1(n14309), .C2(n15097), .A(n14137), .B(n14136), .ZN(
        n14138) );
  OAI21_X1 U16253 ( .B1(n14139), .B2(n15092), .A(n14138), .ZN(P1_U3226) );
  XNOR2_X1 U16254 ( .A(n14142), .B(n14141), .ZN(n14143) );
  XNOR2_X1 U16255 ( .A(n14140), .B(n14143), .ZN(n14150) );
  OAI21_X1 U16256 ( .B1(n15086), .B2(n14307), .A(n14144), .ZN(n14145) );
  AOI21_X1 U16257 ( .B1(n15107), .B2(n14761), .A(n14145), .ZN(n14146) );
  OAI21_X1 U16258 ( .B1(n14147), .B2(n15119), .A(n14146), .ZN(n14148) );
  AOI21_X1 U16259 ( .B1(n14851), .B2(n15097), .A(n14148), .ZN(n14149) );
  OAI21_X1 U16260 ( .B1(n14150), .B2(n15092), .A(n14149), .ZN(P1_U3228) );
  NOR3_X1 U16261 ( .A1(n6698), .A2(n7539), .A3(n14152), .ZN(n14154) );
  OAI21_X1 U16262 ( .B1(n14154), .B2(n14153), .A(n15114), .ZN(n14159) );
  OAI22_X1 U16263 ( .A1(n14191), .A2(n14947), .B1(n14174), .B2(n15131), .ZN(
        n14679) );
  INV_X1 U16264 ( .A(n14687), .ZN(n14156) );
  OAI22_X1 U16265 ( .A1(n14156), .A2(n15119), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14155), .ZN(n14157) );
  AOI21_X1 U16266 ( .B1(n14679), .B2(n14195), .A(n14157), .ZN(n14158) );
  OAI211_X1 U16267 ( .C1(n14690), .C2(n15111), .A(n14159), .B(n14158), .ZN(
        P1_U3229) );
  XNOR2_X1 U16268 ( .A(n14160), .B(n14161), .ZN(n14168) );
  NOR2_X1 U16269 ( .A1(n14162), .A2(n15131), .ZN(n14163) );
  AOI21_X1 U16270 ( .B1(n14487), .B2(n15134), .A(n14163), .ZN(n14739) );
  OAI22_X1 U16271 ( .A1(n14739), .A2(n14203), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14164), .ZN(n14166) );
  NOR2_X1 U16272 ( .A1(n14746), .A2(n15111), .ZN(n14165) );
  AOI211_X1 U16273 ( .C1(n14205), .C2(n14744), .A(n14166), .B(n14165), .ZN(
        n14167) );
  OAI21_X1 U16274 ( .B1(n14168), .B2(n15092), .A(n14167), .ZN(P1_U3233) );
  INV_X1 U16275 ( .A(n14169), .ZN(n14170) );
  NOR2_X1 U16276 ( .A1(n14171), .A2(n14170), .ZN(n14173) );
  AOI21_X1 U16277 ( .B1(n14173), .B2(n14111), .A(n14172), .ZN(n14178) );
  OAI22_X1 U16278 ( .A1(n14174), .A2(n14947), .B1(n7453), .B2(n15131), .ZN(
        n14712) );
  AOI22_X1 U16279 ( .A1(n14712), .A2(n14195), .B1(P1_REG3_REG_22__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14175) );
  OAI21_X1 U16280 ( .B1(n14713), .B2(n15119), .A(n14175), .ZN(n14176) );
  AOI21_X1 U16281 ( .B1(n14718), .B2(n15097), .A(n14176), .ZN(n14177) );
  OAI21_X1 U16282 ( .B1(n14178), .B2(n15092), .A(n14177), .ZN(P1_U3235) );
  AOI21_X1 U16283 ( .B1(n14180), .B2(n14179), .A(n6700), .ZN(n14186) );
  INV_X1 U16284 ( .A(n14181), .ZN(n14183) );
  NAND2_X1 U16285 ( .A1(n14844), .A2(n14195), .ZN(n14182) );
  NAND2_X1 U16286 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n15268)
         );
  OAI211_X1 U16287 ( .C1(n15119), .C2(n14183), .A(n14182), .B(n15268), .ZN(
        n14184) );
  AOI21_X1 U16288 ( .B1(n14845), .B2(n15097), .A(n14184), .ZN(n14185) );
  OAI21_X1 U16289 ( .B1(n14186), .B2(n15092), .A(n14185), .ZN(P1_U3238) );
  OAI21_X1 U16290 ( .B1(n14189), .B2(n14188), .A(n14187), .ZN(n14190) );
  NAND2_X1 U16291 ( .A1(n14190), .A2(n15114), .ZN(n14197) );
  OAI22_X1 U16292 ( .A1(n14192), .A2(n14947), .B1(n14191), .B2(n15131), .ZN(
        n14792) );
  OAI22_X1 U16293 ( .A1(n14652), .A2(n15119), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14193), .ZN(n14194) );
  AOI21_X1 U16294 ( .B1(n14792), .B2(n14195), .A(n14194), .ZN(n14196) );
  OAI211_X1 U16295 ( .C1(n14656), .C2(n15111), .A(n14197), .B(n14196), .ZN(
        P1_U3240) );
  OAI211_X1 U16296 ( .C1(n14200), .C2(n14199), .A(n14198), .B(n15114), .ZN(
        n14208) );
  INV_X1 U16297 ( .A(n14201), .ZN(n14206) );
  OAI22_X1 U16298 ( .A1(n14203), .A2(n15153), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14202), .ZN(n14204) );
  AOI21_X1 U16299 ( .B1(n14206), .B2(n14205), .A(n14204), .ZN(n14207) );
  OAI211_X1 U16300 ( .C1(n7512), .C2(n15111), .A(n14208), .B(n14207), .ZN(
        P1_U3241) );
  NAND2_X1 U16301 ( .A1(n14212), .A2(n14211), .ZN(n14382) );
  INV_X1 U16302 ( .A(n14229), .ZN(n14335) );
  MUX2_X1 U16303 ( .A(n14656), .B(n14666), .S(n14335), .Z(n14361) );
  INV_X1 U16304 ( .A(n14229), .ZN(n14364) );
  MUX2_X1 U16305 ( .A(n15087), .B(n15112), .S(n14364), .Z(n14295) );
  INV_X1 U16306 ( .A(n14214), .ZN(n14215) );
  NAND2_X1 U16307 ( .A1(n14229), .A2(n14228), .ZN(n14231) );
  NAND2_X1 U16308 ( .A1(n14337), .A2(n6672), .ZN(n14230) );
  MUX2_X1 U16309 ( .A(n14231), .B(n14230), .S(n14500), .Z(n14232) );
  MUX2_X1 U16310 ( .A(n14233), .B(n14499), .S(n14337), .Z(n14237) );
  MUX2_X1 U16311 ( .A(n14499), .B(n14233), .S(n14411), .Z(n14234) );
  NAND2_X1 U16312 ( .A1(n14235), .A2(n14234), .ZN(n14241) );
  NAND2_X1 U16313 ( .A1(n14239), .A2(n14238), .ZN(n14240) );
  MUX2_X1 U16314 ( .A(n15293), .B(n14498), .S(n14390), .Z(n14245) );
  NAND2_X1 U16315 ( .A1(n14244), .A2(n14245), .ZN(n14243) );
  MUX2_X1 U16316 ( .A(n15293), .B(n14498), .S(n14364), .Z(n14242) );
  NAND2_X1 U16317 ( .A1(n14243), .A2(n14242), .ZN(n14249) );
  INV_X1 U16318 ( .A(n14244), .ZN(n14247) );
  INV_X1 U16319 ( .A(n14245), .ZN(n14246) );
  NAND2_X1 U16320 ( .A1(n14247), .A2(n14246), .ZN(n14248) );
  MUX2_X1 U16321 ( .A(n14250), .B(n14497), .S(n14364), .Z(n14252) );
  MUX2_X1 U16322 ( .A(n14497), .B(n14250), .S(n14411), .Z(n14251) );
  INV_X1 U16323 ( .A(n14252), .ZN(n14253) );
  MUX2_X1 U16324 ( .A(n15309), .B(n14496), .S(n14229), .Z(n14257) );
  NAND2_X1 U16325 ( .A1(n14256), .A2(n14257), .ZN(n14255) );
  MUX2_X1 U16326 ( .A(n15309), .B(n14496), .S(n14364), .Z(n14254) );
  NAND2_X1 U16327 ( .A1(n14255), .A2(n14254), .ZN(n14261) );
  INV_X1 U16328 ( .A(n14256), .ZN(n14259) );
  INV_X1 U16329 ( .A(n14257), .ZN(n14258) );
  NAND2_X1 U16330 ( .A1(n14259), .A2(n14258), .ZN(n14260) );
  MUX2_X1 U16331 ( .A(n14495), .B(n14262), .S(n14390), .Z(n14264) );
  MUX2_X1 U16332 ( .A(n14495), .B(n14262), .S(n14411), .Z(n14263) );
  INV_X1 U16333 ( .A(n14264), .ZN(n14265) );
  MUX2_X1 U16334 ( .A(n14494), .B(n14266), .S(n14335), .Z(n14270) );
  NAND2_X1 U16335 ( .A1(n14269), .A2(n14270), .ZN(n14268) );
  MUX2_X1 U16336 ( .A(n14494), .B(n14266), .S(n14229), .Z(n14267) );
  NAND2_X1 U16337 ( .A1(n14268), .A2(n14267), .ZN(n14274) );
  INV_X1 U16338 ( .A(n14269), .ZN(n14272) );
  INV_X1 U16339 ( .A(n14270), .ZN(n14271) );
  NAND2_X1 U16340 ( .A1(n14272), .A2(n14271), .ZN(n14273) );
  MUX2_X1 U16341 ( .A(n14493), .B(n14275), .S(n14390), .Z(n14277) );
  MUX2_X1 U16342 ( .A(n14493), .B(n14275), .S(n14337), .Z(n14276) );
  MUX2_X1 U16343 ( .A(n14492), .B(n14279), .S(n14335), .Z(n14283) );
  NAND2_X1 U16344 ( .A1(n14282), .A2(n14283), .ZN(n14281) );
  MUX2_X1 U16345 ( .A(n14492), .B(n14279), .S(n14229), .Z(n14280) );
  NAND2_X1 U16346 ( .A1(n14281), .A2(n14280), .ZN(n14287) );
  INV_X1 U16347 ( .A(n14282), .ZN(n14285) );
  INV_X1 U16348 ( .A(n14283), .ZN(n14284) );
  NAND2_X1 U16349 ( .A1(n14285), .A2(n14284), .ZN(n14286) );
  MUX2_X1 U16350 ( .A(n15108), .B(n14917), .S(n14390), .Z(n14289) );
  NAND2_X1 U16351 ( .A1(n14288), .A2(n14289), .ZN(n14293) );
  MUX2_X1 U16352 ( .A(n15108), .B(n14917), .S(n14335), .Z(n14292) );
  INV_X1 U16353 ( .A(n14288), .ZN(n14291) );
  INV_X1 U16354 ( .A(n14289), .ZN(n14290) );
  MUX2_X1 U16355 ( .A(n14491), .B(n15172), .S(n14229), .Z(n14294) );
  NAND2_X1 U16356 ( .A1(n14303), .A2(n14299), .ZN(n14302) );
  NAND2_X1 U16357 ( .A1(n14304), .A2(n14300), .ZN(n14301) );
  MUX2_X1 U16358 ( .A(n14302), .B(n14301), .S(n14335), .Z(n14306) );
  MUX2_X1 U16359 ( .A(n14304), .B(n14303), .S(n14411), .Z(n14305) );
  XOR2_X1 U16360 ( .A(n15135), .B(n14851), .Z(n14314) );
  MUX2_X1 U16361 ( .A(n14307), .B(n15148), .S(n14229), .Z(n14319) );
  AND2_X1 U16362 ( .A1(n14489), .A2(n14390), .ZN(n14308) );
  AOI21_X1 U16363 ( .B1(n14309), .B2(n14411), .A(n14308), .ZN(n14312) );
  NAND2_X1 U16364 ( .A1(n14851), .A2(n14310), .ZN(n14311) );
  NAND3_X1 U16365 ( .A1(n14313), .A2(n14312), .A3(n14311), .ZN(n14320) );
  OAI21_X1 U16366 ( .B1(n14314), .B2(n14319), .A(n14320), .ZN(n14315) );
  AND2_X1 U16367 ( .A1(n15135), .A2(n14335), .ZN(n14317) );
  OAI21_X1 U16368 ( .B1(n14335), .B2(n15135), .A(n14851), .ZN(n14316) );
  OAI21_X1 U16369 ( .B1(n14317), .B2(n14851), .A(n14316), .ZN(n14318) );
  OAI21_X1 U16370 ( .B1(n14320), .B2(n14319), .A(n14318), .ZN(n14321) );
  INV_X1 U16371 ( .A(n14321), .ZN(n14322) );
  INV_X1 U16372 ( .A(n14327), .ZN(n14330) );
  MUX2_X1 U16373 ( .A(n14324), .B(n14323), .S(n14335), .Z(n14325) );
  OAI211_X1 U16374 ( .C1(n14330), .C2(n14329), .A(n14755), .B(n14328), .ZN(
        n14334) );
  MUX2_X1 U16375 ( .A(n14332), .B(n14331), .S(n14411), .Z(n14333) );
  MUX2_X1 U16376 ( .A(n14746), .B(n14336), .S(n14335), .Z(n14339) );
  MUX2_X1 U16377 ( .A(n14763), .B(n14832), .S(n14337), .Z(n14338) );
  MUX2_X1 U16378 ( .A(n14827), .B(n14487), .S(n14364), .Z(n14343) );
  INV_X1 U16379 ( .A(n14341), .ZN(n14342) );
  INV_X1 U16380 ( .A(n14347), .ZN(n14350) );
  MUX2_X1 U16381 ( .A(n14820), .B(n14344), .S(n14335), .Z(n14346) );
  INV_X1 U16382 ( .A(n14346), .ZN(n14349) );
  INV_X1 U16383 ( .A(n14344), .ZN(n14486) );
  MUX2_X1 U16384 ( .A(n14486), .B(n14718), .S(n14335), .Z(n14345) );
  OAI21_X1 U16385 ( .B1(n14350), .B2(n14349), .A(n14348), .ZN(n14351) );
  MUX2_X1 U16386 ( .A(n14485), .B(n14812), .S(n14411), .Z(n14352) );
  MUX2_X1 U16387 ( .A(n14812), .B(n14485), .S(n14335), .Z(n14353) );
  MUX2_X1 U16388 ( .A(n14690), .B(n14665), .S(n14335), .Z(n14355) );
  MUX2_X1 U16389 ( .A(n14484), .B(n14806), .S(n14411), .Z(n14354) );
  MUX2_X1 U16390 ( .A(n14483), .B(n14674), .S(n14335), .Z(n14359) );
  NAND2_X1 U16391 ( .A1(n14358), .A2(n14359), .ZN(n14357) );
  MUX2_X1 U16392 ( .A(n14674), .B(n14483), .S(n14411), .Z(n14356) );
  MUX2_X1 U16393 ( .A(n14482), .B(n14793), .S(n14364), .Z(n14360) );
  MUX2_X1 U16394 ( .A(n14481), .B(n14786), .S(n14335), .Z(n14367) );
  MUX2_X1 U16395 ( .A(n14786), .B(n14481), .S(n14364), .Z(n14365) );
  MUX2_X1 U16396 ( .A(n14780), .B(n14368), .S(n14335), .Z(n14371) );
  MUX2_X1 U16397 ( .A(n14480), .B(n14369), .S(n14335), .Z(n14370) );
  NAND2_X1 U16398 ( .A1(n14372), .A2(n14407), .ZN(n14374) );
  OR2_X1 U16399 ( .A1(n14408), .A2(n14877), .ZN(n14373) );
  INV_X1 U16400 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n14379) );
  NAND2_X1 U16401 ( .A1(n14375), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n14378) );
  NAND2_X1 U16402 ( .A1(n14376), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n14377) );
  OAI211_X1 U16403 ( .C1(n14380), .C2(n14379), .A(n14378), .B(n14377), .ZN(
        n14477) );
  NAND2_X1 U16404 ( .A1(n14335), .A2(n14477), .ZN(n14385) );
  NAND2_X1 U16405 ( .A1(n14382), .A2(n14381), .ZN(n14384) );
  AOI21_X1 U16406 ( .B1(n14385), .B2(n14384), .A(n14383), .ZN(n14386) );
  AOI21_X1 U16407 ( .B1(n14417), .B2(n14229), .A(n14386), .ZN(n14402) );
  OAI21_X1 U16408 ( .B1(n14477), .B2(n14387), .A(n14478), .ZN(n14388) );
  INV_X1 U16409 ( .A(n14388), .ZN(n14389) );
  MUX2_X1 U16410 ( .A(n14389), .B(n14417), .S(n14411), .Z(n14399) );
  MUX2_X1 U16411 ( .A(n14392), .B(n14391), .S(n14390), .Z(n14396) );
  INV_X1 U16412 ( .A(n14392), .ZN(n14479) );
  MUX2_X1 U16413 ( .A(n14479), .B(n14393), .S(n14335), .Z(n14395) );
  AOI22_X1 U16414 ( .A1(n14402), .A2(n14399), .B1(n14396), .B2(n14395), .ZN(
        n14394) );
  INV_X1 U16415 ( .A(n14395), .ZN(n14398) );
  INV_X1 U16416 ( .A(n14396), .ZN(n14397) );
  INV_X1 U16417 ( .A(n14399), .ZN(n14400) );
  OAI21_X1 U16418 ( .B1(n14401), .B2(n14403), .A(n14400), .ZN(n14405) );
  NAND2_X1 U16419 ( .A1(n14875), .A2(n14407), .ZN(n14410) );
  INV_X1 U16420 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n14870) );
  OR2_X1 U16421 ( .A1(n14408), .A2(n14870), .ZN(n14409) );
  NAND2_X1 U16422 ( .A1(n14462), .A2(n14364), .ZN(n14465) );
  NOR2_X1 U16423 ( .A1(n14462), .A2(n14411), .ZN(n14457) );
  NAND2_X1 U16424 ( .A1(n14413), .A2(n14412), .ZN(n14415) );
  NAND2_X1 U16425 ( .A1(n14415), .A2(n14414), .ZN(n14464) );
  NAND2_X1 U16426 ( .A1(n14464), .A2(n14459), .ZN(n14461) );
  AOI21_X1 U16427 ( .B1(n14457), .B2(n14477), .A(n14461), .ZN(n14416) );
  OAI21_X1 U16428 ( .B1(n14477), .B2(n14465), .A(n14416), .ZN(n14452) );
  INV_X1 U16429 ( .A(n14477), .ZN(n14625) );
  XNOR2_X1 U16430 ( .A(n14462), .B(n14625), .ZN(n14454) );
  NOR2_X1 U16431 ( .A1(n14419), .A2(n14418), .ZN(n14423) );
  NAND4_X1 U16432 ( .A1(n14423), .A2(n14422), .A3(n6807), .A4(n14420), .ZN(
        n14424) );
  NOR2_X1 U16433 ( .A1(n14425), .A2(n14424), .ZN(n14428) );
  NAND4_X1 U16434 ( .A1(n14429), .A2(n14428), .A3(n14427), .A4(n14426), .ZN(
        n14430) );
  OR4_X1 U16435 ( .A1(n14433), .A2(n14432), .A3(n14431), .A4(n14430), .ZN(
        n14434) );
  NOR2_X1 U16436 ( .A1(n14923), .A2(n14434), .ZN(n14435) );
  AND2_X1 U16437 ( .A1(n14954), .A2(n14435), .ZN(n14436) );
  NAND4_X1 U16438 ( .A1(n14439), .A2(n14438), .A3(n14437), .A4(n14436), .ZN(
        n14440) );
  NOR4_X1 U16439 ( .A1(n14441), .A2(n7610), .A3(n15130), .A4(n14440), .ZN(
        n14443) );
  NAND4_X1 U16440 ( .A1(n14709), .A2(n14443), .A3(n14747), .A4(n14442), .ZN(
        n14444) );
  NOR4_X1 U16441 ( .A1(n14657), .A2(n14694), .A3(n14683), .A4(n14444), .ZN(
        n14447) );
  XOR2_X1 U16442 ( .A(n14619), .B(n14450), .Z(n14451) );
  OAI22_X1 U16443 ( .A1(n14453), .A2(n14452), .B1(n14459), .B2(n14451), .ZN(
        n14471) );
  INV_X1 U16444 ( .A(n14454), .ZN(n14456) );
  INV_X1 U16445 ( .A(n14464), .ZN(n14455) );
  NAND2_X1 U16446 ( .A1(n14456), .A2(n14455), .ZN(n14469) );
  INV_X1 U16447 ( .A(n14457), .ZN(n14458) );
  XNOR2_X1 U16448 ( .A(n14458), .B(n14464), .ZN(n14460) );
  NAND4_X1 U16449 ( .A1(n14460), .A2(n14772), .A3(n14459), .A4(n14477), .ZN(
        n14468) );
  INV_X1 U16450 ( .A(n14461), .ZN(n14463) );
  NAND4_X1 U16451 ( .A1(n14465), .A2(n14625), .A3(n14463), .A4(n14462), .ZN(
        n14467) );
  NOR3_X1 U16452 ( .A1(n14472), .A2(n6676), .A3(n15131), .ZN(n14474) );
  OAI21_X1 U16453 ( .B1(n14475), .B2(n9742), .A(P1_B_REG_SCAN_IN), .ZN(n14473)
         );
  MUX2_X1 U16454 ( .A(n14477), .B(P1_DATAO_REG_31__SCAN_IN), .S(n14501), .Z(
        P1_U3591) );
  MUX2_X1 U16455 ( .A(n14478), .B(P1_DATAO_REG_30__SCAN_IN), .S(n14501), .Z(
        P1_U3590) );
  INV_X1 U16456 ( .A(P1_U4016), .ZN(n14504) );
  MUX2_X1 U16457 ( .A(n14479), .B(P1_DATAO_REG_29__SCAN_IN), .S(n14504), .Z(
        P1_U3589) );
  MUX2_X1 U16458 ( .A(n14480), .B(P1_DATAO_REG_28__SCAN_IN), .S(n14501), .Z(
        P1_U3588) );
  MUX2_X1 U16459 ( .A(n14481), .B(P1_DATAO_REG_27__SCAN_IN), .S(n14504), .Z(
        P1_U3587) );
  MUX2_X1 U16460 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n14482), .S(P1_U4016), .Z(
        P1_U3586) );
  MUX2_X1 U16461 ( .A(n14483), .B(P1_DATAO_REG_25__SCAN_IN), .S(n14501), .Z(
        P1_U3585) );
  MUX2_X1 U16462 ( .A(n14484), .B(P1_DATAO_REG_24__SCAN_IN), .S(n14501), .Z(
        P1_U3584) );
  MUX2_X1 U16463 ( .A(n14485), .B(P1_DATAO_REG_23__SCAN_IN), .S(n14504), .Z(
        P1_U3583) );
  MUX2_X1 U16464 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n14486), .S(P1_U4016), .Z(
        P1_U3582) );
  MUX2_X1 U16465 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n14487), .S(P1_U4016), .Z(
        P1_U3581) );
  MUX2_X1 U16466 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n14763), .S(P1_U4016), .Z(
        P1_U3580) );
  MUX2_X1 U16467 ( .A(n14488), .B(P1_DATAO_REG_19__SCAN_IN), .S(n14501), .Z(
        P1_U3579) );
  MUX2_X1 U16468 ( .A(n14761), .B(P1_DATAO_REG_18__SCAN_IN), .S(n14501), .Z(
        P1_U3578) );
  MUX2_X1 U16469 ( .A(n15135), .B(P1_DATAO_REG_17__SCAN_IN), .S(n14504), .Z(
        P1_U3577) );
  MUX2_X1 U16470 ( .A(n14489), .B(P1_DATAO_REG_16__SCAN_IN), .S(n14504), .Z(
        P1_U3576) );
  MUX2_X1 U16471 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n14490), .S(P1_U4016), .Z(
        P1_U3575) );
  MUX2_X1 U16472 ( .A(n15106), .B(P1_DATAO_REG_14__SCAN_IN), .S(n14501), .Z(
        P1_U3574) );
  MUX2_X1 U16473 ( .A(n14491), .B(P1_DATAO_REG_13__SCAN_IN), .S(n14504), .Z(
        P1_U3573) );
  MUX2_X1 U16474 ( .A(n15108), .B(P1_DATAO_REG_12__SCAN_IN), .S(n14504), .Z(
        P1_U3572) );
  MUX2_X1 U16475 ( .A(n14492), .B(P1_DATAO_REG_11__SCAN_IN), .S(n14504), .Z(
        P1_U3571) );
  MUX2_X1 U16476 ( .A(n14493), .B(P1_DATAO_REG_10__SCAN_IN), .S(n14504), .Z(
        P1_U3570) );
  MUX2_X1 U16477 ( .A(n14494), .B(P1_DATAO_REG_9__SCAN_IN), .S(n14501), .Z(
        P1_U3569) );
  MUX2_X1 U16478 ( .A(n14495), .B(P1_DATAO_REG_8__SCAN_IN), .S(n14504), .Z(
        P1_U3568) );
  MUX2_X1 U16479 ( .A(n14496), .B(P1_DATAO_REG_7__SCAN_IN), .S(n14504), .Z(
        P1_U3567) );
  MUX2_X1 U16480 ( .A(n14497), .B(P1_DATAO_REG_6__SCAN_IN), .S(n14501), .Z(
        P1_U3566) );
  MUX2_X1 U16481 ( .A(n14498), .B(P1_DATAO_REG_5__SCAN_IN), .S(n14501), .Z(
        P1_U3565) );
  MUX2_X1 U16482 ( .A(n14499), .B(P1_DATAO_REG_4__SCAN_IN), .S(n14504), .Z(
        P1_U3564) );
  MUX2_X1 U16483 ( .A(n14500), .B(P1_DATAO_REG_3__SCAN_IN), .S(n14501), .Z(
        P1_U3563) );
  MUX2_X1 U16484 ( .A(n14502), .B(P1_DATAO_REG_2__SCAN_IN), .S(n14501), .Z(
        P1_U3562) );
  MUX2_X1 U16485 ( .A(n6847), .B(P1_DATAO_REG_1__SCAN_IN), .S(n14504), .Z(
        P1_U3561) );
  MUX2_X1 U16486 ( .A(n6808), .B(P1_DATAO_REG_0__SCAN_IN), .S(n14504), .Z(
        P1_U3560) );
  INV_X1 U16487 ( .A(n14512), .ZN(n14509) );
  OAI22_X1 U16488 ( .A1(n15270), .A2(n9900), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14506), .ZN(n14508) );
  AOI21_X1 U16489 ( .B1(n14509), .B2(n15232), .A(n14508), .ZN(n14517) );
  OAI211_X1 U16490 ( .C1(n14511), .C2(n14510), .A(n15261), .B(n14527), .ZN(
        n14516) );
  MUX2_X1 U16491 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n10571), .S(n14512), .Z(
        n14513) );
  INV_X1 U16492 ( .A(n14513), .ZN(n14514) );
  OAI211_X1 U16493 ( .C1(n14519), .C2(n14514), .A(n15258), .B(n14533), .ZN(
        n14515) );
  NAND3_X1 U16494 ( .A1(n14517), .A2(n14516), .A3(n14515), .ZN(P1_U3244) );
  MUX2_X1 U16495 ( .A(n14519), .B(n14518), .S(n6676), .Z(n14521) );
  NAND2_X1 U16496 ( .A1(n14521), .A2(n14520), .ZN(n14522) );
  OAI211_X1 U16497 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n14523), .A(n14522), .B(
        P1_U4016), .ZN(n15236) );
  OAI22_X1 U16498 ( .A1(n15270), .A2(n9901), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14524), .ZN(n14525) );
  AOI21_X1 U16499 ( .B1(n14530), .B2(n15232), .A(n14525), .ZN(n14538) );
  MUX2_X1 U16500 ( .A(n10550), .B(P1_REG1_REG_2__SCAN_IN), .S(n14530), .Z(
        n14528) );
  NAND3_X1 U16501 ( .A1(n14528), .A2(n14527), .A3(n14526), .ZN(n14529) );
  NAND3_X1 U16502 ( .A1(n15261), .A2(n14544), .A3(n14529), .ZN(n14537) );
  MUX2_X1 U16503 ( .A(n14531), .B(P1_REG2_REG_2__SCAN_IN), .S(n14530), .Z(
        n14534) );
  NAND3_X1 U16504 ( .A1(n14534), .A2(n14533), .A3(n14532), .ZN(n14535) );
  NAND3_X1 U16505 ( .A1(n15258), .A2(n14549), .A3(n14535), .ZN(n14536) );
  NAND4_X1 U16506 ( .A1(n15236), .A2(n14538), .A3(n14537), .A4(n14536), .ZN(
        P1_U3245) );
  INV_X1 U16507 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n14540) );
  OAI22_X1 U16508 ( .A1(n15270), .A2(n14540), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14539), .ZN(n14541) );
  AOI21_X1 U16509 ( .B1(n14546), .B2(n15232), .A(n14541), .ZN(n14553) );
  MUX2_X1 U16510 ( .A(n10554), .B(P1_REG1_REG_3__SCAN_IN), .S(n14546), .Z(
        n14543) );
  NAND3_X1 U16511 ( .A1(n14544), .A2(n14543), .A3(n14542), .ZN(n14545) );
  NAND3_X1 U16512 ( .A1(n15261), .A2(n15223), .A3(n14545), .ZN(n14552) );
  MUX2_X1 U16513 ( .A(n11140), .B(P1_REG2_REG_3__SCAN_IN), .S(n14546), .Z(
        n14548) );
  NAND3_X1 U16514 ( .A1(n14549), .A2(n14548), .A3(n14547), .ZN(n14550) );
  NAND3_X1 U16515 ( .A1(n15258), .A2(n15228), .A3(n14550), .ZN(n14551) );
  NAND3_X1 U16516 ( .A1(n14553), .A2(n14552), .A3(n14551), .ZN(P1_U3246) );
  OAI21_X1 U16517 ( .B1(n15270), .B2(n14555), .A(n14554), .ZN(n14556) );
  AOI21_X1 U16518 ( .B1(n14557), .B2(n15232), .A(n14556), .ZN(n14569) );
  OAI21_X1 U16519 ( .B1(n14560), .B2(n14559), .A(n14558), .ZN(n14561) );
  NAND2_X1 U16520 ( .A1(n15261), .A2(n14561), .ZN(n14568) );
  MUX2_X1 U16521 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n11470), .S(n14562), .Z(
        n14564) );
  NAND3_X1 U16522 ( .A1(n14564), .A2(n15230), .A3(n14563), .ZN(n14565) );
  NAND3_X1 U16523 ( .A1(n15258), .A2(n14566), .A3(n14565), .ZN(n14567) );
  NAND3_X1 U16524 ( .A1(n14569), .A2(n14568), .A3(n14567), .ZN(P1_U3248) );
  NOR2_X1 U16525 ( .A1(n14571), .A2(n14570), .ZN(n14572) );
  OAI21_X1 U16526 ( .B1(n14572), .B2(n14587), .A(n15261), .ZN(n14583) );
  OAI21_X1 U16527 ( .B1(n15270), .B2(n14574), .A(n14573), .ZN(n14575) );
  AOI21_X1 U16528 ( .B1(n14576), .B2(n15232), .A(n14575), .ZN(n14582) );
  MUX2_X1 U16529 ( .A(n10597), .B(P1_REG2_REG_8__SCAN_IN), .S(n14576), .Z(
        n14577) );
  NAND3_X1 U16530 ( .A1(n14579), .A2(n14578), .A3(n14577), .ZN(n14580) );
  NAND3_X1 U16531 ( .A1(n15258), .A2(n14597), .A3(n14580), .ZN(n14581) );
  NAND3_X1 U16532 ( .A1(n14583), .A2(n14582), .A3(n14581), .ZN(P1_U3251) );
  INV_X1 U16533 ( .A(n14584), .ZN(n14589) );
  NOR3_X1 U16534 ( .A1(n14587), .A2(n14586), .A3(n14585), .ZN(n14588) );
  OAI21_X1 U16535 ( .B1(n14589), .B2(n14588), .A(n15261), .ZN(n14602) );
  NOR2_X1 U16536 ( .A1(n15266), .A2(n14590), .ZN(n14591) );
  AOI211_X1 U16537 ( .C1(n14593), .C2(P1_ADDR_REG_9__SCAN_IN), .A(n14592), .B(
        n14591), .ZN(n14601) );
  MUX2_X1 U16538 ( .A(n10600), .B(P1_REG2_REG_9__SCAN_IN), .S(n14594), .Z(
        n14595) );
  NAND3_X1 U16539 ( .A1(n14597), .A2(n14596), .A3(n14595), .ZN(n14598) );
  NAND3_X1 U16540 ( .A1(n15258), .A2(n14599), .A3(n14598), .ZN(n14600) );
  NAND3_X1 U16541 ( .A1(n14602), .A2(n14601), .A3(n14600), .ZN(P1_U3252) );
  INV_X1 U16542 ( .A(n14603), .ZN(n14604) );
  AOI21_X1 U16543 ( .B1(n14605), .B2(P1_REG1_REG_17__SCAN_IN), .A(n14604), 
        .ZN(n14606) );
  XNOR2_X1 U16544 ( .A(n14606), .B(n14611), .ZN(n15262) );
  NAND2_X1 U16545 ( .A1(P1_REG1_REG_18__SCAN_IN), .A2(n15262), .ZN(n15260) );
  OR2_X1 U16546 ( .A1(n14606), .A2(n15265), .ZN(n14607) );
  NAND2_X1 U16547 ( .A1(n15260), .A2(n14607), .ZN(n14608) );
  XOR2_X1 U16548 ( .A(n14608), .B(P1_REG1_REG_19__SCAN_IN), .Z(n14618) );
  INV_X1 U16549 ( .A(n14618), .ZN(n14616) );
  NAND2_X1 U16550 ( .A1(n14610), .A2(n14609), .ZN(n14612) );
  XOR2_X1 U16551 ( .A(n14611), .B(n14612), .Z(n15259) );
  NAND2_X1 U16552 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n15259), .ZN(n15257) );
  NAND2_X1 U16553 ( .A1(n14612), .A2(n14611), .ZN(n14613) );
  NAND2_X1 U16554 ( .A1(n15257), .A2(n14613), .ZN(n14614) );
  XOR2_X1 U16555 ( .A(n14614), .B(P1_REG2_REG_19__SCAN_IN), .Z(n14617) );
  OAI21_X1 U16556 ( .B1(n14617), .B2(n15248), .A(n15266), .ZN(n14615) );
  AOI21_X1 U16557 ( .B1(n14616), .B2(n15261), .A(n14615), .ZN(n14621) );
  AOI22_X1 U16558 ( .A1(n14618), .A2(n15261), .B1(n15258), .B2(n14617), .ZN(
        n14620) );
  MUX2_X1 U16559 ( .A(n14621), .B(n14620), .S(n14619), .Z(n14623) );
  OAI211_X1 U16560 ( .C1(n7717), .C2(n15270), .A(n14623), .B(n14622), .ZN(
        P1_U3262) );
  NAND2_X1 U16561 ( .A1(n14630), .A2(n14775), .ZN(n14629) );
  XNOR2_X1 U16562 ( .A(n14629), .B(n14772), .ZN(n14624) );
  NAND2_X1 U16563 ( .A1(n14624), .A2(n15122), .ZN(n14771) );
  OR2_X1 U16564 ( .A1(n14626), .A2(n14625), .ZN(n14773) );
  NOR2_X1 U16565 ( .A1(n14765), .A2(n14773), .ZN(n14632) );
  NOR2_X1 U16566 ( .A1(n14772), .A2(n15141), .ZN(n14627) );
  AOI211_X1 U16567 ( .C1(n14765), .C2(P1_REG2_REG_31__SCAN_IN), .A(n14632), 
        .B(n14627), .ZN(n14628) );
  OAI21_X1 U16568 ( .B1(n14958), .B2(n14771), .A(n14628), .ZN(P1_U3263) );
  OAI211_X1 U16569 ( .C1(n14630), .C2(n14775), .A(n15122), .B(n14629), .ZN(
        n14774) );
  NOR2_X1 U16570 ( .A1(n14775), .A2(n15141), .ZN(n14631) );
  AOI211_X1 U16571 ( .C1(n14765), .C2(P1_REG2_REG_30__SCAN_IN), .A(n14632), 
        .B(n14631), .ZN(n14633) );
  OAI21_X1 U16572 ( .B1(n14958), .B2(n14774), .A(n14633), .ZN(P1_U3264) );
  XNOR2_X1 U16573 ( .A(n14634), .B(n14636), .ZN(n14784) );
  OAI21_X1 U16574 ( .B1(n14637), .B2(n14636), .A(n14635), .ZN(n14638) );
  INV_X1 U16575 ( .A(n14638), .ZN(n14782) );
  OAI211_X1 U16576 ( .C1(n14780), .C2(n6702), .A(n15122), .B(n14639), .ZN(
        n14779) );
  NOR2_X1 U16577 ( .A1(n14779), .A2(n14958), .ZN(n14645) );
  INV_X1 U16578 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n14640) );
  OAI22_X1 U16579 ( .A1(n14641), .A2(n15136), .B1(n14640), .B2(n15143), .ZN(
        n14642) );
  AOI21_X1 U16580 ( .B1(n14777), .B2(n15143), .A(n14642), .ZN(n14643) );
  OAI21_X1 U16581 ( .B1(n14780), .B2(n15141), .A(n14643), .ZN(n14644) );
  AOI211_X1 U16582 ( .C1(n14782), .C2(n15126), .A(n14645), .B(n14644), .ZN(
        n14646) );
  OAI21_X1 U16583 ( .B1(n14784), .B2(n14959), .A(n14646), .ZN(P1_U3265) );
  OAI21_X1 U16584 ( .B1(n14648), .B2(n14657), .A(n14647), .ZN(n14796) );
  INV_X1 U16585 ( .A(n14668), .ZN(n14651) );
  INV_X1 U16586 ( .A(n14649), .ZN(n14650) );
  AOI211_X1 U16587 ( .C1(n14793), .C2(n14651), .A(n14741), .B(n14650), .ZN(
        n14791) );
  INV_X1 U16588 ( .A(n14652), .ZN(n14653) );
  AOI22_X1 U16589 ( .A1(n14653), .A2(n14929), .B1(P1_REG2_REG_26__SCAN_IN), 
        .B2(n14765), .ZN(n14655) );
  NAND2_X1 U16590 ( .A1(n14792), .A2(n15143), .ZN(n14654) );
  OAI211_X1 U16591 ( .C1(n14656), .C2(n15141), .A(n14655), .B(n14654), .ZN(
        n14660) );
  AOI21_X1 U16592 ( .B1(n14658), .B2(n14657), .A(n12521), .ZN(n14790) );
  NOR2_X1 U16593 ( .A1(n14790), .A2(n14959), .ZN(n14659) );
  AOI211_X1 U16594 ( .C1(n14791), .C2(n15125), .A(n14660), .B(n14659), .ZN(
        n14661) );
  OAI21_X1 U16595 ( .B1(n14750), .B2(n14796), .A(n14661), .ZN(P1_U3267) );
  AOI21_X1 U16596 ( .B1(n14669), .B2(n14663), .A(n14662), .ZN(n14664) );
  OAI222_X1 U16597 ( .A1(n14947), .A2(n14666), .B1(n15131), .B2(n14665), .C1(
        n15175), .C2(n14664), .ZN(n14803) );
  AND2_X1 U16598 ( .A1(n14685), .A2(n14674), .ZN(n14667) );
  OR3_X1 U16599 ( .A1(n14668), .A2(n14667), .A3(n14741), .ZN(n14799) );
  OR2_X1 U16600 ( .A1(n14670), .A2(n14669), .ZN(n14798) );
  NAND3_X1 U16601 ( .A1(n14798), .A2(n15126), .A3(n14797), .ZN(n14676) );
  INV_X1 U16602 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n14671) );
  OAI22_X1 U16603 ( .A1(n14672), .A2(n15136), .B1(n14671), .B2(n15143), .ZN(
        n14673) );
  AOI21_X1 U16604 ( .B1(n14674), .B2(n14717), .A(n14673), .ZN(n14675) );
  OAI211_X1 U16605 ( .C1(n14799), .C2(n14958), .A(n14676), .B(n14675), .ZN(
        n14677) );
  AOI21_X1 U16606 ( .B1(n14803), .B2(n15143), .A(n14677), .ZN(n14678) );
  INV_X1 U16607 ( .A(n14678), .ZN(P1_U3268) );
  AOI21_X1 U16608 ( .B1(n6744), .B2(n14683), .A(n15175), .ZN(n14681) );
  AOI21_X1 U16609 ( .B1(n14681), .B2(n14680), .A(n14679), .ZN(n14808) );
  OAI21_X1 U16610 ( .B1(n14684), .B2(n14683), .A(n14682), .ZN(n14804) );
  AOI21_X1 U16611 ( .B1(n14806), .B2(n14696), .A(n14741), .ZN(n14686) );
  AND2_X1 U16612 ( .A1(n14686), .A2(n14685), .ZN(n14805) );
  NAND2_X1 U16613 ( .A1(n14805), .A2(n15125), .ZN(n14689) );
  AOI22_X1 U16614 ( .A1(n14687), .A2(n14929), .B1(P1_REG2_REG_24__SCAN_IN), 
        .B2(n14765), .ZN(n14688) );
  OAI211_X1 U16615 ( .C1(n14690), .C2(n15141), .A(n14689), .B(n14688), .ZN(
        n14691) );
  AOI21_X1 U16616 ( .B1(n14804), .B2(n15126), .A(n14691), .ZN(n14692) );
  OAI21_X1 U16617 ( .B1(n14808), .B2(n14765), .A(n14692), .ZN(P1_U3269) );
  AOI21_X1 U16618 ( .B1(n14695), .B2(n14694), .A(n14693), .ZN(n14817) );
  AOI21_X1 U16619 ( .B1(n14812), .B2(n14711), .A(n14741), .ZN(n14697) );
  AND2_X1 U16620 ( .A1(n14697), .A2(n14696), .ZN(n14810) );
  NAND2_X1 U16621 ( .A1(n14812), .A2(n14717), .ZN(n14702) );
  INV_X1 U16622 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n14698) );
  OAI22_X1 U16623 ( .A1(n14699), .A2(n15136), .B1(n14698), .B2(n15143), .ZN(
        n14700) );
  AOI21_X1 U16624 ( .B1(n14811), .B2(n15143), .A(n14700), .ZN(n14701) );
  NAND2_X1 U16625 ( .A1(n14702), .A2(n14701), .ZN(n14703) );
  AOI21_X1 U16626 ( .B1(n14810), .B2(n15125), .A(n14703), .ZN(n14707) );
  NAND2_X1 U16627 ( .A1(n14705), .A2(n14704), .ZN(n14813) );
  NAND3_X1 U16628 ( .A1(n14814), .A2(n14813), .A3(n15126), .ZN(n14706) );
  OAI211_X1 U16629 ( .C1(n14817), .C2(n14959), .A(n14707), .B(n14706), .ZN(
        P1_U3270) );
  XNOR2_X1 U16630 ( .A(n14708), .B(n14709), .ZN(n14824) );
  XNOR2_X1 U16631 ( .A(n14710), .B(n14709), .ZN(n14822) );
  OAI211_X1 U16632 ( .C1(n14820), .C2(n14729), .A(n15122), .B(n14711), .ZN(
        n14819) );
  INV_X1 U16633 ( .A(n14712), .ZN(n14818) );
  INV_X1 U16634 ( .A(n14713), .ZN(n14714) );
  AOI22_X1 U16635 ( .A1(n14714), .A2(n14929), .B1(P1_REG2_REG_22__SCAN_IN), 
        .B2(n14931), .ZN(n14715) );
  OAI21_X1 U16636 ( .B1(n14818), .B2(n14765), .A(n14715), .ZN(n14716) );
  AOI21_X1 U16637 ( .B1(n14718), .B2(n14717), .A(n14716), .ZN(n14719) );
  OAI21_X1 U16638 ( .B1(n14819), .B2(n14958), .A(n14719), .ZN(n14720) );
  AOI21_X1 U16639 ( .B1(n14822), .B2(n14721), .A(n14720), .ZN(n14722) );
  OAI21_X1 U16640 ( .B1(n14824), .B2(n14750), .A(n14722), .ZN(P1_U3271) );
  XNOR2_X1 U16641 ( .A(n14723), .B(n14727), .ZN(n14725) );
  AOI21_X1 U16642 ( .B1(n14725), .B2(n15160), .A(n14724), .ZN(n14829) );
  OAI21_X1 U16643 ( .B1(n14728), .B2(n14727), .A(n14726), .ZN(n14825) );
  AOI211_X1 U16644 ( .C1(n14827), .C2(n14742), .A(n14741), .B(n14729), .ZN(
        n14826) );
  NAND2_X1 U16645 ( .A1(n14826), .A2(n15125), .ZN(n14733) );
  INV_X1 U16646 ( .A(n14730), .ZN(n14731) );
  AOI22_X1 U16647 ( .A1(n14731), .A2(n14929), .B1(n14931), .B2(
        P1_REG2_REG_21__SCAN_IN), .ZN(n14732) );
  OAI211_X1 U16648 ( .C1(n14734), .C2(n15141), .A(n14733), .B(n14732), .ZN(
        n14735) );
  AOI21_X1 U16649 ( .B1(n15126), .B2(n14825), .A(n14735), .ZN(n14736) );
  OAI21_X1 U16650 ( .B1(n14829), .B2(n14765), .A(n14736), .ZN(P1_U3272) );
  OAI211_X1 U16651 ( .C1(n14738), .C2(n14747), .A(n14737), .B(n15160), .ZN(
        n14740) );
  AND2_X1 U16652 ( .A1(n14740), .A2(n14739), .ZN(n14834) );
  AOI21_X1 U16653 ( .B1(n14832), .B2(n14760), .A(n14741), .ZN(n14743) );
  AND2_X1 U16654 ( .A1(n14743), .A2(n14742), .ZN(n14831) );
  AOI22_X1 U16655 ( .A1(n14931), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n14744), 
        .B2(n14929), .ZN(n14745) );
  OAI21_X1 U16656 ( .B1(n14746), .B2(n15141), .A(n14745), .ZN(n14752) );
  INV_X1 U16657 ( .A(n14747), .ZN(n14749) );
  OAI21_X1 U16658 ( .B1(n14749), .B2(n6791), .A(n14748), .ZN(n14835) );
  NOR2_X1 U16659 ( .A1(n14835), .A2(n14750), .ZN(n14751) );
  AOI211_X1 U16660 ( .C1(n14831), .C2(n15125), .A(n14752), .B(n14751), .ZN(
        n14753) );
  OAI21_X1 U16661 ( .B1(n14765), .B2(n14834), .A(n14753), .ZN(P1_U3273) );
  XNOR2_X1 U16662 ( .A(n14754), .B(n7610), .ZN(n14842) );
  XNOR2_X1 U16663 ( .A(n14756), .B(n14755), .ZN(n14840) );
  NAND2_X1 U16664 ( .A1(n14758), .A2(n14757), .ZN(n14759) );
  NAND3_X1 U16665 ( .A1(n14760), .A2(n15122), .A3(n14759), .ZN(n14837) );
  AOI22_X1 U16666 ( .A1(n14763), .A2(n15134), .B1(n14762), .B2(n14761), .ZN(
        n14836) );
  OAI22_X1 U16667 ( .A1(n14836), .A2(n14765), .B1(n14764), .B2(n15136), .ZN(
        n14767) );
  NOR2_X1 U16668 ( .A1(n14838), .A2(n15141), .ZN(n14766) );
  AOI211_X1 U16669 ( .C1(n14931), .C2(P1_REG2_REG_19__SCAN_IN), .A(n14767), 
        .B(n14766), .ZN(n14768) );
  OAI21_X1 U16670 ( .B1(n14958), .B2(n14837), .A(n14768), .ZN(n14769) );
  AOI21_X1 U16671 ( .B1(n15126), .B2(n14840), .A(n14769), .ZN(n14770) );
  OAI21_X1 U16672 ( .B1(n14842), .B2(n14959), .A(n14770), .ZN(P1_U3274) );
  OAI211_X1 U16673 ( .C1(n14772), .C2(n15334), .A(n14771), .B(n14773), .ZN(
        n14855) );
  MUX2_X1 U16674 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n14855), .S(n15358), .Z(
        P1_U3559) );
  OAI211_X1 U16675 ( .C1(n14775), .C2(n15334), .A(n14774), .B(n14773), .ZN(
        n14856) );
  MUX2_X1 U16676 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n14856), .S(n15358), .Z(
        P1_U3558) );
  INV_X1 U16677 ( .A(n14777), .ZN(n14778) );
  OAI211_X1 U16678 ( .C1(n14780), .C2(n15334), .A(n14779), .B(n14778), .ZN(
        n14781) );
  OAI21_X1 U16679 ( .B1(n14784), .B2(n15175), .A(n14783), .ZN(n14857) );
  MUX2_X1 U16680 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n14857), .S(n15358), .Z(
        P1_U3556) );
  AOI21_X1 U16681 ( .B1(n15310), .B2(n14786), .A(n14785), .ZN(n14787) );
  OAI211_X1 U16682 ( .C1(n14789), .C2(n15313), .A(n14788), .B(n14787), .ZN(
        n14858) );
  MUX2_X1 U16683 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n14858), .S(n15358), .Z(
        P1_U3555) );
  OR2_X1 U16684 ( .A1(n14790), .A2(n15175), .ZN(n14795) );
  AOI211_X1 U16685 ( .C1(n15310), .C2(n14793), .A(n14792), .B(n14791), .ZN(
        n14794) );
  OAI211_X1 U16686 ( .C1(n15155), .C2(n14796), .A(n14795), .B(n14794), .ZN(
        n14859) );
  MUX2_X1 U16687 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n14859), .S(n15358), .Z(
        P1_U3554) );
  NAND3_X1 U16688 ( .A1(n14798), .A2(n15337), .A3(n14797), .ZN(n14800) );
  OAI211_X1 U16689 ( .C1(n14801), .C2(n15334), .A(n14800), .B(n14799), .ZN(
        n14802) );
  OR2_X1 U16690 ( .A1(n14803), .A2(n14802), .ZN(n14860) );
  MUX2_X1 U16691 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n14860), .S(n15358), .Z(
        P1_U3553) );
  INV_X1 U16692 ( .A(n14804), .ZN(n14809) );
  AOI21_X1 U16693 ( .B1(n15310), .B2(n14806), .A(n14805), .ZN(n14807) );
  OAI211_X1 U16694 ( .C1(n15155), .C2(n14809), .A(n14808), .B(n14807), .ZN(
        n14861) );
  MUX2_X1 U16695 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n14861), .S(n15358), .Z(
        P1_U3552) );
  AOI211_X1 U16696 ( .C1(n15310), .C2(n14812), .A(n14811), .B(n14810), .ZN(
        n14816) );
  NAND3_X1 U16697 ( .A1(n14814), .A2(n15337), .A3(n14813), .ZN(n14815) );
  OAI211_X1 U16698 ( .C1(n14817), .C2(n15175), .A(n14816), .B(n14815), .ZN(
        n14862) );
  MUX2_X1 U16699 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n14862), .S(n15358), .Z(
        P1_U3551) );
  OAI211_X1 U16700 ( .C1(n15334), .C2(n14820), .A(n14819), .B(n14818), .ZN(
        n14821) );
  AOI21_X1 U16701 ( .B1(n14822), .B2(n15160), .A(n14821), .ZN(n14823) );
  OAI21_X1 U16702 ( .B1(n15155), .B2(n14824), .A(n14823), .ZN(n14863) );
  MUX2_X1 U16703 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n14863), .S(n15358), .Z(
        P1_U3550) );
  INV_X1 U16704 ( .A(n14825), .ZN(n14830) );
  AOI21_X1 U16705 ( .B1(n15310), .B2(n14827), .A(n14826), .ZN(n14828) );
  OAI211_X1 U16706 ( .C1(n15155), .C2(n14830), .A(n14829), .B(n14828), .ZN(
        n14864) );
  MUX2_X1 U16707 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n14864), .S(n15358), .Z(
        P1_U3549) );
  AOI21_X1 U16708 ( .B1(n15310), .B2(n14832), .A(n14831), .ZN(n14833) );
  OAI211_X1 U16709 ( .C1(n15155), .C2(n14835), .A(n14834), .B(n14833), .ZN(
        n14865) );
  MUX2_X1 U16710 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n14865), .S(n15358), .Z(
        P1_U3548) );
  OAI211_X1 U16711 ( .C1(n14838), .C2(n15334), .A(n14837), .B(n14836), .ZN(
        n14839) );
  AOI21_X1 U16712 ( .B1(n14840), .B2(n15337), .A(n14839), .ZN(n14841) );
  OAI21_X1 U16713 ( .B1(n14842), .B2(n15175), .A(n14841), .ZN(n14866) );
  MUX2_X1 U16714 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n14866), .S(n15358), .Z(
        P1_U3547) );
  AOI211_X1 U16715 ( .C1(n15310), .C2(n14845), .A(n14844), .B(n14843), .ZN(
        n14847) );
  OAI211_X1 U16716 ( .C1(n15155), .C2(n14848), .A(n14847), .B(n14846), .ZN(
        n14867) );
  MUX2_X1 U16717 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n14867), .S(n15358), .Z(
        P1_U3546) );
  AOI211_X1 U16718 ( .C1(n15310), .C2(n14851), .A(n14850), .B(n14849), .ZN(
        n14852) );
  OAI21_X1 U16719 ( .B1(n15155), .B2(n14853), .A(n14852), .ZN(n14868) );
  MUX2_X1 U16720 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n14868), .S(n15358), .Z(
        P1_U3545) );
  MUX2_X1 U16721 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n14854), .S(n15358), .Z(
        P1_U3528) );
  MUX2_X1 U16722 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n14855), .S(n15341), .Z(
        P1_U3527) );
  MUX2_X1 U16723 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n14856), .S(n15341), .Z(
        P1_U3526) );
  MUX2_X1 U16724 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n14857), .S(n15341), .Z(
        P1_U3524) );
  MUX2_X1 U16725 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n14858), .S(n15341), .Z(
        P1_U3523) );
  MUX2_X1 U16726 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n14859), .S(n15341), .Z(
        P1_U3522) );
  MUX2_X1 U16727 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n14860), .S(n15341), .Z(
        P1_U3521) );
  MUX2_X1 U16728 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n14861), .S(n15341), .Z(
        P1_U3520) );
  MUX2_X1 U16729 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n14862), .S(n15341), .Z(
        P1_U3519) );
  MUX2_X1 U16730 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n14863), .S(n15341), .Z(
        P1_U3518) );
  MUX2_X1 U16731 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n14864), .S(n15341), .Z(
        P1_U3517) );
  MUX2_X1 U16732 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n14865), .S(n15341), .Z(
        P1_U3516) );
  MUX2_X1 U16733 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n14866), .S(n15341), .Z(
        P1_U3515) );
  MUX2_X1 U16734 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n14867), .S(n15341), .Z(
        P1_U3513) );
  MUX2_X1 U16735 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n14868), .S(n15341), .Z(
        P1_U3510) );
  NAND3_X1 U16736 ( .A1(n7402), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        P1_STATE_REG_SCAN_IN), .ZN(n14871) );
  OAI22_X1 U16737 ( .A1(n14872), .A2(n14871), .B1(n14870), .B2(n14869), .ZN(
        n14873) );
  AOI21_X1 U16738 ( .B1(n14875), .B2(n14874), .A(n14873), .ZN(n14876) );
  INV_X1 U16739 ( .A(n14876), .ZN(P1_U3324) );
  OAI222_X1 U16740 ( .A1(n14885), .A2(n14879), .B1(P1_U3086), .B2(n14878), 
        .C1(n14877), .C2(n14891), .ZN(P1_U3325) );
  OAI222_X1 U16741 ( .A1(n14885), .A2(n14882), .B1(P1_U3086), .B2(n14881), 
        .C1(n14880), .C2(n14891), .ZN(P1_U3326) );
  OAI222_X1 U16742 ( .A1(n14891), .A2(n14886), .B1(n14885), .B2(n14884), .C1(
        n6676), .C2(P1_U3086), .ZN(P1_U3328) );
  OAI222_X1 U16743 ( .A1(n14891), .A2(n14890), .B1(n14885), .B2(n14889), .C1(
        n14888), .C2(P1_U3086), .ZN(P1_U3329) );
  MUX2_X1 U16744 ( .A(n9742), .B(n14892), .S(P1_U3086), .Z(P1_U3333) );
  MUX2_X1 U16745 ( .A(n14893), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  AOI21_X1 U16746 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n14897) );
  OAI21_X1 U16747 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n14897), 
        .ZN(U28) );
  AOI21_X1 U16748 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n14898) );
  OAI21_X1 U16749 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n14898), 
        .ZN(U29) );
  OAI21_X1 U16750 ( .B1(n14901), .B2(n14900), .A(n14899), .ZN(n14902) );
  XNOR2_X1 U16751 ( .A(n14902), .B(P2_ADDR_REG_2__SCAN_IN), .ZN(SUB_1596_U61)
         );
  AOI21_X1 U16752 ( .B1(n14905), .B2(n14904), .A(n14903), .ZN(SUB_1596_U57) );
  OAI21_X1 U16753 ( .B1(n14908), .B2(n14907), .A(n14906), .ZN(SUB_1596_U55) );
  AOI21_X1 U16754 ( .B1(n14911), .B2(n14910), .A(n14909), .ZN(SUB_1596_U54) );
  AOI21_X1 U16755 ( .B1(n14914), .B2(n14913), .A(n14912), .ZN(n14915) );
  XOR2_X1 U16756 ( .A(P2_ADDR_REG_10__SCAN_IN), .B(n14915), .Z(SUB_1596_U70)
         );
  XNOR2_X1 U16757 ( .A(n14916), .B(n7593), .ZN(n14937) );
  NAND2_X1 U16758 ( .A1(n14918), .A2(n14917), .ZN(n14919) );
  NAND3_X1 U16759 ( .A1(n14920), .A2(n15122), .A3(n14919), .ZN(n14938) );
  OAI22_X1 U16760 ( .A1(n14937), .A2(n14921), .B1(n14958), .B2(n14938), .ZN(
        n14922) );
  INV_X1 U16761 ( .A(n14922), .ZN(n14936) );
  XNOR2_X1 U16762 ( .A(n14924), .B(n14923), .ZN(n14927) );
  INV_X1 U16763 ( .A(n14925), .ZN(n14926) );
  AOI21_X1 U16764 ( .B1(n14927), .B2(n15160), .A(n14926), .ZN(n14939) );
  OAI21_X1 U16765 ( .B1(n14928), .B2(n14937), .A(n14939), .ZN(n14934) );
  AOI22_X1 U16766 ( .A1(n14931), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n14930), 
        .B2(n14929), .ZN(n14932) );
  OAI21_X1 U16767 ( .B1(n14940), .B2(n15141), .A(n14932), .ZN(n14933) );
  AOI21_X1 U16768 ( .B1(n14934), .B2(n15143), .A(n14933), .ZN(n14935) );
  NAND2_X1 U16769 ( .A1(n14936), .A2(n14935), .ZN(P1_U3281) );
  INV_X1 U16770 ( .A(n14937), .ZN(n14942) );
  OAI211_X1 U16771 ( .C1(n14940), .C2(n15334), .A(n14939), .B(n14938), .ZN(
        n14941) );
  AOI21_X1 U16772 ( .B1(n14942), .B2(n15337), .A(n14941), .ZN(n14945) );
  INV_X1 U16773 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n14943) );
  AOI22_X1 U16774 ( .A1(n15341), .A2(n14945), .B1(n14943), .B2(n15339), .ZN(
        P1_U3495) );
  AOI22_X1 U16775 ( .A1(n15358), .A2(n14945), .B1(n14944), .B2(n15355), .ZN(
        P1_U3540) );
  OAI22_X1 U16776 ( .A1(n14948), .A2(n14947), .B1(n14946), .B2(n15131), .ZN(
        n15171) );
  INV_X1 U16777 ( .A(n15171), .ZN(n14949) );
  OAI211_X1 U16778 ( .C1(n15112), .C2(n14950), .A(n14949), .B(n15143), .ZN(
        n14951) );
  OAI21_X1 U16779 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n15143), .A(n14951), 
        .ZN(n14962) );
  XNOR2_X1 U16780 ( .A(n14953), .B(n14952), .ZN(n15178) );
  XNOR2_X1 U16781 ( .A(n14955), .B(n14954), .ZN(n15176) );
  OAI211_X1 U16782 ( .C1(n15112), .C2(n14957), .A(n15122), .B(n14956), .ZN(
        n15173) );
  OAI22_X1 U16783 ( .A1(n15176), .A2(n14959), .B1(n14958), .B2(n15173), .ZN(
        n14960) );
  AOI21_X1 U16784 ( .B1(n15126), .B2(n15178), .A(n14960), .ZN(n14961) );
  OAI211_X1 U16785 ( .C1(n15136), .C2(n15118), .A(n14962), .B(n14961), .ZN(
        P1_U3280) );
  AOI21_X1 U16786 ( .B1(n14965), .B2(n14964), .A(n14963), .ZN(n14966) );
  XOR2_X1 U16787 ( .A(P2_ADDR_REG_17__SCAN_IN), .B(n14966), .Z(SUB_1596_U63)
         );
  AOI21_X1 U16788 ( .B1(n14969), .B2(n14968), .A(n14967), .ZN(n14983) );
  OAI21_X1 U16789 ( .B1(P3_REG1_REG_15__SCAN_IN), .B2(n14971), .A(n14970), 
        .ZN(n14976) );
  AOI21_X1 U16790 ( .B1(n15623), .B2(P3_ADDR_REG_15__SCAN_IN), .A(n14972), 
        .ZN(n14973) );
  OAI21_X1 U16791 ( .B1(n15626), .B2(n14974), .A(n14973), .ZN(n14975) );
  AOI21_X1 U16792 ( .B1(n14976), .B2(n15628), .A(n14975), .ZN(n14982) );
  AOI21_X1 U16793 ( .B1(n14979), .B2(n14978), .A(n14977), .ZN(n14980) );
  OR2_X1 U16794 ( .A1(n14980), .A2(n15611), .ZN(n14981) );
  OAI211_X1 U16795 ( .C1(n14983), .C2(n15636), .A(n14982), .B(n14981), .ZN(
        P3_U3197) );
  AOI21_X1 U16796 ( .B1(n14986), .B2(n14985), .A(n14984), .ZN(n15005) );
  OAI21_X1 U16797 ( .B1(n14989), .B2(n14988), .A(n14987), .ZN(n14996) );
  NAND2_X1 U16798 ( .A1(n15540), .A2(n14990), .ZN(n14993) );
  INV_X1 U16799 ( .A(n14991), .ZN(n14992) );
  OAI211_X1 U16800 ( .C1(n14994), .C2(n15548), .A(n14993), .B(n14992), .ZN(
        n14995) );
  AOI21_X1 U16801 ( .B1(n14996), .B2(n15628), .A(n14995), .ZN(n15004) );
  INV_X1 U16802 ( .A(n14997), .ZN(n14999) );
  NOR2_X1 U16803 ( .A1(n14999), .A2(n14998), .ZN(n15001) );
  AOI21_X1 U16804 ( .B1(n15002), .B2(n15001), .A(n15611), .ZN(n15000) );
  OAI21_X1 U16805 ( .B1(n15002), .B2(n15001), .A(n15000), .ZN(n15003) );
  OAI211_X1 U16806 ( .C1(n15005), .C2(n15636), .A(n15004), .B(n15003), .ZN(
        P3_U3198) );
  AOI21_X1 U16807 ( .B1(n15008), .B2(n15007), .A(n15006), .ZN(n15022) );
  OAI21_X1 U16808 ( .B1(n15010), .B2(P3_REG1_REG_17__SCAN_IN), .A(n15009), 
        .ZN(n15011) );
  AND2_X1 U16809 ( .A1(n15011), .A2(n15628), .ZN(n15019) );
  AOI211_X1 U16810 ( .C1(n15014), .C2(n15013), .A(n15611), .B(n15012), .ZN(
        n15018) );
  OAI22_X1 U16811 ( .A1(n15626), .A2(n15016), .B1(n15015), .B2(n15548), .ZN(
        n15017) );
  NOR4_X1 U16812 ( .A1(n15020), .A2(n15019), .A3(n15018), .A4(n15017), .ZN(
        n15021) );
  OAI21_X1 U16813 ( .B1(n15022), .B2(n15636), .A(n15021), .ZN(P3_U3199) );
  AOI22_X1 U16814 ( .A1(n15540), .A2(n15023), .B1(n15623), .B2(
        P3_ADDR_REG_18__SCAN_IN), .ZN(n15039) );
  OAI21_X1 U16815 ( .B1(n15026), .B2(n15025), .A(n15024), .ZN(n15031) );
  OAI21_X1 U16816 ( .B1(n15029), .B2(n15028), .A(n15027), .ZN(n15030) );
  AOI22_X1 U16817 ( .A1(n15031), .A2(n15628), .B1(n15630), .B2(n15030), .ZN(
        n15038) );
  OAI221_X1 U16818 ( .B1(n15035), .B2(n15034), .C1(n15035), .C2(n15033), .A(
        n15032), .ZN(n15036) );
  NAND4_X1 U16819 ( .A1(n15039), .A2(n15038), .A3(n15037), .A4(n15036), .ZN(
        P3_U3200) );
  XNOR2_X1 U16820 ( .A(n15040), .B(n8656), .ZN(n15041) );
  NAND2_X1 U16821 ( .A1(n15041), .A2(n15703), .ZN(n15045) );
  AOI22_X1 U16822 ( .A1(n15700), .A2(n15043), .B1(n15042), .B2(n15697), .ZN(
        n15044) );
  NAND2_X1 U16823 ( .A1(n15045), .A2(n15044), .ZN(n15074) );
  OAI22_X1 U16824 ( .A1(n15693), .A2(n8651), .B1(n15675), .B2(n15046), .ZN(
        n15057) );
  NAND2_X1 U16825 ( .A1(n15048), .A2(n15047), .ZN(n15049) );
  NAND2_X1 U16826 ( .A1(n15050), .A2(n15049), .ZN(n15071) );
  INV_X1 U16827 ( .A(n15071), .ZN(n15055) );
  NOR2_X1 U16828 ( .A1(n15051), .A2(n15730), .ZN(n15072) );
  INV_X1 U16829 ( .A(n15072), .ZN(n15052) );
  OAI22_X1 U16830 ( .A1(n15055), .A2(n15054), .B1(n15053), .B2(n15052), .ZN(
        n15056) );
  AOI211_X1 U16831 ( .C1(n15693), .C2(n15074), .A(n15057), .B(n15056), .ZN(
        n15058) );
  INV_X1 U16832 ( .A(n15058), .ZN(P3_U3222) );
  INV_X1 U16833 ( .A(n15059), .ZN(n15062) );
  INV_X1 U16834 ( .A(n15060), .ZN(n15061) );
  AOI211_X1 U16835 ( .C1(n15063), .C2(n15739), .A(n15062), .B(n15061), .ZN(
        n15075) );
  INV_X1 U16836 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n15064) );
  AOI22_X1 U16837 ( .A1(n15751), .A2(n15075), .B1(n15064), .B2(n15749), .ZN(
        P3_U3472) );
  NOR2_X1 U16838 ( .A1(n15066), .A2(n15065), .ZN(n15068) );
  AOI211_X1 U16839 ( .C1(n15070), .C2(n15069), .A(n15068), .B(n15067), .ZN(
        n15077) );
  AOI22_X1 U16840 ( .A1(n15751), .A2(n15077), .B1(n8667), .B2(n15749), .ZN(
        P3_U3471) );
  AND2_X1 U16841 ( .A1(n15071), .A2(n15739), .ZN(n15073) );
  NOR3_X1 U16842 ( .A1(n15074), .A2(n15073), .A3(n15072), .ZN(n15079) );
  AOI22_X1 U16843 ( .A1(n15751), .A2(n15079), .B1(n8650), .B2(n15749), .ZN(
        P3_U3470) );
  INV_X1 U16844 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n15076) );
  AOI22_X1 U16845 ( .A1(n15743), .A2(n15076), .B1(n15075), .B2(n15741), .ZN(
        P3_U3429) );
  INV_X1 U16846 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n15078) );
  AOI22_X1 U16847 ( .A1(n15743), .A2(n15078), .B1(n15077), .B2(n15741), .ZN(
        P3_U3426) );
  INV_X1 U16848 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n15080) );
  AOI22_X1 U16849 ( .A1(n15743), .A2(n15080), .B1(n15079), .B2(n15741), .ZN(
        P3_U3423) );
  OAI21_X1 U16850 ( .B1(n7172), .B2(n15516), .A(n15081), .ZN(n15083) );
  AOI211_X1 U16851 ( .C1(n15084), .C2(n15491), .A(n15083), .B(n15082), .ZN(
        n15085) );
  AOI22_X1 U16852 ( .A1(n15539), .A2(n15085), .B1(n13690), .B2(n15536), .ZN(
        P2_U3512) );
  AOI22_X1 U16853 ( .A1(n15524), .A2(n15085), .B1(n7981), .B2(n15523), .ZN(
        P2_U3469) );
  OAI22_X1 U16854 ( .A1(n15088), .A2(n15132), .B1(n15087), .B2(n15086), .ZN(
        n15096) );
  INV_X1 U16855 ( .A(n15089), .ZN(n15091) );
  OAI21_X1 U16856 ( .B1(n15091), .B2(n15102), .A(n15090), .ZN(n15094) );
  AOI21_X1 U16857 ( .B1(n15094), .B2(n15093), .A(n15092), .ZN(n15095) );
  AOI211_X1 U16858 ( .C1(n15164), .C2(n15097), .A(n15096), .B(n15095), .ZN(
        n15099) );
  OAI211_X1 U16859 ( .C1(n15119), .C2(n15100), .A(n15099), .B(n15098), .ZN(
        P1_U3215) );
  INV_X1 U16860 ( .A(n15102), .ZN(n15104) );
  NAND2_X1 U16861 ( .A1(n15104), .A2(n15103), .ZN(n15105) );
  XNOR2_X1 U16862 ( .A(n15101), .B(n15105), .ZN(n15115) );
  AOI22_X1 U16863 ( .A1(n15109), .A2(n15108), .B1(n15107), .B2(n15106), .ZN(
        n15110) );
  OAI21_X1 U16864 ( .B1(n15112), .B2(n15111), .A(n15110), .ZN(n15113) );
  AOI21_X1 U16865 ( .B1(n15115), .B2(n15114), .A(n15113), .ZN(n15117) );
  OAI211_X1 U16866 ( .C1(n15119), .C2(n15118), .A(n15117), .B(n15116), .ZN(
        P1_U3234) );
  XNOR2_X1 U16867 ( .A(n15120), .B(n15130), .ZN(n15151) );
  INV_X1 U16868 ( .A(n15121), .ZN(n15123) );
  OAI211_X1 U16869 ( .C1(n15148), .C2(n15123), .A(n15122), .B(n6693), .ZN(
        n15147) );
  INV_X1 U16870 ( .A(n15147), .ZN(n15124) );
  AOI22_X1 U16871 ( .A1(n15151), .A2(n15126), .B1(n15125), .B2(n15124), .ZN(
        n15145) );
  INV_X1 U16872 ( .A(n15127), .ZN(n15128) );
  AOI21_X1 U16873 ( .B1(n15130), .B2(n15129), .A(n15128), .ZN(n15133) );
  OAI22_X1 U16874 ( .A1(n15133), .A2(n15175), .B1(n15132), .B2(n15131), .ZN(
        n15149) );
  NAND2_X1 U16875 ( .A1(n15135), .A2(n15134), .ZN(n15146) );
  INV_X1 U16876 ( .A(n15146), .ZN(n15139) );
  OAI22_X1 U16877 ( .A1(n15143), .A2(n12000), .B1(n15137), .B2(n15136), .ZN(
        n15138) );
  AOI21_X1 U16878 ( .B1(n15139), .B2(n15143), .A(n15138), .ZN(n15140) );
  OAI21_X1 U16879 ( .B1(n15148), .B2(n15141), .A(n15140), .ZN(n15142) );
  AOI21_X1 U16880 ( .B1(n15149), .B2(n15143), .A(n15142), .ZN(n15144) );
  NAND2_X1 U16881 ( .A1(n15145), .A2(n15144), .ZN(P1_U3277) );
  OAI211_X1 U16882 ( .C1(n15148), .C2(n15334), .A(n15147), .B(n15146), .ZN(
        n15150) );
  AOI211_X1 U16883 ( .C1(n15151), .C2(n15337), .A(n15150), .B(n15149), .ZN(
        n15187) );
  AOI22_X1 U16884 ( .A1(n15358), .A2(n15187), .B1(n15152), .B2(n15355), .ZN(
        P1_U3544) );
  OAI211_X1 U16885 ( .C1(n7512), .C2(n15334), .A(n15154), .B(n15153), .ZN(
        n15158) );
  NOR2_X1 U16886 ( .A1(n15156), .A2(n15155), .ZN(n15157) );
  AOI211_X1 U16887 ( .C1(n15160), .C2(n15159), .A(n15158), .B(n15157), .ZN(
        n15189) );
  INV_X1 U16888 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n15161) );
  AOI22_X1 U16889 ( .A1(n15358), .A2(n15189), .B1(n15161), .B2(n15355), .ZN(
        P1_U3543) );
  NAND3_X1 U16890 ( .A1(n15163), .A2(n15162), .A3(n15337), .ZN(n15167) );
  NAND2_X1 U16891 ( .A1(n15164), .A2(n15310), .ZN(n15165) );
  AND3_X1 U16892 ( .A1(n15167), .A2(n15166), .A3(n15165), .ZN(n15168) );
  AND2_X1 U16893 ( .A1(n15169), .A2(n15168), .ZN(n15191) );
  AOI22_X1 U16894 ( .A1(n15358), .A2(n15191), .B1(n15170), .B2(n15355), .ZN(
        P1_U3542) );
  AOI21_X1 U16895 ( .B1(n15172), .B2(n15310), .A(n15171), .ZN(n15174) );
  OAI211_X1 U16896 ( .C1(n15176), .C2(n15175), .A(n15174), .B(n15173), .ZN(
        n15177) );
  AOI21_X1 U16897 ( .B1(n15178), .B2(n15337), .A(n15177), .ZN(n15193) );
  AOI22_X1 U16898 ( .A1(n15358), .A2(n15193), .B1(n10893), .B2(n15355), .ZN(
        P1_U3541) );
  AND2_X1 U16899 ( .A1(n15179), .A2(n15337), .ZN(n15183) );
  OAI21_X1 U16900 ( .B1(n15181), .B2(n15334), .A(n15180), .ZN(n15182) );
  NOR3_X1 U16901 ( .A1(n15184), .A2(n15183), .A3(n15182), .ZN(n15195) );
  AOI22_X1 U16902 ( .A1(n15358), .A2(n15195), .B1(n15185), .B2(n15355), .ZN(
        P1_U3539) );
  INV_X1 U16903 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n15186) );
  AOI22_X1 U16904 ( .A1(n15341), .A2(n15187), .B1(n15186), .B2(n15339), .ZN(
        P1_U3507) );
  INV_X1 U16905 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n15188) );
  AOI22_X1 U16906 ( .A1(n15341), .A2(n15189), .B1(n15188), .B2(n15339), .ZN(
        P1_U3504) );
  INV_X1 U16907 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n15190) );
  AOI22_X1 U16908 ( .A1(n15341), .A2(n15191), .B1(n15190), .B2(n15339), .ZN(
        P1_U3501) );
  INV_X1 U16909 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n15192) );
  AOI22_X1 U16910 ( .A1(n15341), .A2(n15193), .B1(n15192), .B2(n15339), .ZN(
        P1_U3498) );
  INV_X1 U16911 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n15194) );
  AOI22_X1 U16912 ( .A1(n15341), .A2(n15195), .B1(n15194), .B2(n15339), .ZN(
        P1_U3492) );
  AOI21_X1 U16913 ( .B1(n15198), .B2(n15197), .A(n15196), .ZN(n15199) );
  XOR2_X1 U16914 ( .A(P2_ADDR_REG_11__SCAN_IN), .B(n15199), .Z(SUB_1596_U69)
         );
  OAI21_X1 U16915 ( .B1(n15202), .B2(n15201), .A(n15200), .ZN(n15203) );
  XNOR2_X1 U16916 ( .A(n15203), .B(P2_ADDR_REG_12__SCAN_IN), .ZN(SUB_1596_U68)
         );
  OAI222_X1 U16917 ( .A1(n15208), .A2(n15207), .B1(n15208), .B2(n15206), .C1(
        n15205), .C2(n15204), .ZN(SUB_1596_U67) );
  OAI21_X1 U16918 ( .B1(n15211), .B2(n15210), .A(n15209), .ZN(n15212) );
  XNOR2_X1 U16919 ( .A(n15212), .B(P2_ADDR_REG_14__SCAN_IN), .ZN(SUB_1596_U66)
         );
  AOI21_X1 U16920 ( .B1(n15215), .B2(n15214), .A(n15213), .ZN(n15216) );
  XOR2_X1 U16921 ( .A(P2_ADDR_REG_15__SCAN_IN), .B(n15216), .Z(SUB_1596_U65)
         );
  AOI21_X1 U16922 ( .B1(n15219), .B2(n15218), .A(n15217), .ZN(n15220) );
  XOR2_X1 U16923 ( .A(P2_ADDR_REG_16__SCAN_IN), .B(n15220), .Z(SUB_1596_U64)
         );
  MUX2_X1 U16924 ( .A(n10557), .B(P1_REG1_REG_4__SCAN_IN), .S(n15231), .Z(
        n15221) );
  NAND3_X1 U16925 ( .A1(n15223), .A2(n15222), .A3(n15221), .ZN(n15224) );
  NAND3_X1 U16926 ( .A1(n15261), .A2(n15225), .A3(n15224), .ZN(n15235) );
  MUX2_X1 U16927 ( .A(n10577), .B(P1_REG2_REG_4__SCAN_IN), .S(n15231), .Z(
        n15226) );
  NAND3_X1 U16928 ( .A1(n15228), .A2(n15227), .A3(n15226), .ZN(n15229) );
  NAND3_X1 U16929 ( .A1(n15258), .A2(n15230), .A3(n15229), .ZN(n15234) );
  NAND2_X1 U16930 ( .A1(n15232), .A2(n15231), .ZN(n15233) );
  AND4_X1 U16931 ( .A1(n15236), .A2(n15235), .A3(n15234), .A4(n15233), .ZN(
        n15238) );
  OAI211_X1 U16932 ( .C1(n15270), .C2(n15239), .A(n15238), .B(n15237), .ZN(
        P1_U3247) );
  AOI21_X1 U16933 ( .B1(n15242), .B2(n15241), .A(n15240), .ZN(n15244) );
  OR2_X1 U16934 ( .A1(n15244), .A2(n15243), .ZN(n15251) );
  AOI21_X1 U16935 ( .B1(n15247), .B2(n15246), .A(n15245), .ZN(n15249) );
  OR2_X1 U16936 ( .A1(n15249), .A2(n15248), .ZN(n15250) );
  OAI211_X1 U16937 ( .C1(n15266), .C2(n15252), .A(n15251), .B(n15250), .ZN(
        n15253) );
  INV_X1 U16938 ( .A(n15253), .ZN(n15255) );
  OAI211_X1 U16939 ( .C1(n15256), .C2(n15270), .A(n15255), .B(n15254), .ZN(
        P1_U3255) );
  OAI211_X1 U16940 ( .C1(n15259), .C2(P1_REG2_REG_18__SCAN_IN), .A(n15258), 
        .B(n15257), .ZN(n15264) );
  OAI211_X1 U16941 ( .C1(P1_REG1_REG_18__SCAN_IN), .C2(n15262), .A(n15261), 
        .B(n15260), .ZN(n15263) );
  OAI211_X1 U16942 ( .C1(n15266), .C2(n15265), .A(n15264), .B(n15263), .ZN(
        n15267) );
  INV_X1 U16943 ( .A(n15267), .ZN(n15269) );
  OAI211_X1 U16944 ( .C1(n15271), .C2(n15270), .A(n15269), .B(n15268), .ZN(
        P1_U3261) );
  AND2_X1 U16945 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n15272), .ZN(P1_U3294) );
  AND2_X1 U16946 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n15272), .ZN(P1_U3295) );
  AND2_X1 U16947 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n15272), .ZN(P1_U3296) );
  AND2_X1 U16948 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n15272), .ZN(P1_U3297) );
  AND2_X1 U16949 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n15272), .ZN(P1_U3298) );
  AND2_X1 U16950 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n15272), .ZN(P1_U3299) );
  AND2_X1 U16951 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n15272), .ZN(P1_U3300) );
  AND2_X1 U16952 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n15272), .ZN(P1_U3301) );
  AND2_X1 U16953 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n15272), .ZN(P1_U3302) );
  AND2_X1 U16954 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n15272), .ZN(P1_U3303) );
  AND2_X1 U16955 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n15272), .ZN(P1_U3304) );
  AND2_X1 U16956 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n15272), .ZN(P1_U3305) );
  AND2_X1 U16957 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n15272), .ZN(P1_U3306) );
  AND2_X1 U16958 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n15272), .ZN(P1_U3307) );
  AND2_X1 U16959 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n15272), .ZN(P1_U3308) );
  AND2_X1 U16960 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n15272), .ZN(P1_U3309) );
  AND2_X1 U16961 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n15272), .ZN(P1_U3310) );
  AND2_X1 U16962 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n15272), .ZN(P1_U3311) );
  AND2_X1 U16963 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n15272), .ZN(P1_U3312) );
  AND2_X1 U16964 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n15272), .ZN(P1_U3313) );
  AND2_X1 U16965 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n15272), .ZN(P1_U3314) );
  AND2_X1 U16966 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n15272), .ZN(P1_U3315) );
  AND2_X1 U16967 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n15272), .ZN(P1_U3316) );
  AND2_X1 U16968 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n15272), .ZN(P1_U3317) );
  AND2_X1 U16969 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n15272), .ZN(P1_U3318) );
  AND2_X1 U16970 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n15272), .ZN(P1_U3319) );
  AND2_X1 U16971 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n15272), .ZN(P1_U3320) );
  AND2_X1 U16972 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n15272), .ZN(P1_U3321) );
  AND2_X1 U16973 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n15272), .ZN(P1_U3322) );
  AND2_X1 U16974 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n15272), .ZN(P1_U3323) );
  INV_X1 U16975 ( .A(n15313), .ZN(n15331) );
  INV_X1 U16976 ( .A(n15273), .ZN(n15274) );
  OAI21_X1 U16977 ( .B1(n10815), .B2(n15334), .A(n15274), .ZN(n15277) );
  INV_X1 U16978 ( .A(n15275), .ZN(n15276) );
  AOI211_X1 U16979 ( .C1(n15331), .C2(n15278), .A(n15277), .B(n15276), .ZN(
        n15342) );
  INV_X1 U16980 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n15279) );
  AOI22_X1 U16981 ( .A1(n15341), .A2(n15342), .B1(n15279), .B2(n15339), .ZN(
        P1_U3462) );
  OAI21_X1 U16982 ( .B1(n15281), .B2(n15334), .A(n15280), .ZN(n15284) );
  INV_X1 U16983 ( .A(n15282), .ZN(n15283) );
  AOI211_X1 U16984 ( .C1(n15331), .C2(n15285), .A(n15284), .B(n15283), .ZN(
        n15343) );
  INV_X1 U16985 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n15286) );
  AOI22_X1 U16986 ( .A1(n15341), .A2(n15343), .B1(n15286), .B2(n15339), .ZN(
        P1_U3465) );
  OAI21_X1 U16987 ( .B1(n15288), .B2(n15334), .A(n15287), .ZN(n15290) );
  AOI211_X1 U16988 ( .C1(n15291), .C2(n15337), .A(n15290), .B(n15289), .ZN(
        n15344) );
  INV_X1 U16989 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n15292) );
  AOI22_X1 U16990 ( .A1(n15341), .A2(n15344), .B1(n15292), .B2(n15339), .ZN(
        P1_U3471) );
  NAND2_X1 U16991 ( .A1(n15299), .A2(n15331), .ZN(n15296) );
  NAND2_X1 U16992 ( .A1(n15293), .A2(n15310), .ZN(n15294) );
  NAND4_X1 U16993 ( .A1(n15297), .A2(n15296), .A3(n15295), .A4(n15294), .ZN(
        n15298) );
  AOI21_X1 U16994 ( .B1(n15317), .B2(n15299), .A(n15298), .ZN(n15346) );
  INV_X1 U16995 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n15300) );
  AOI22_X1 U16996 ( .A1(n15341), .A2(n15346), .B1(n15300), .B2(n15339), .ZN(
        P1_U3474) );
  INV_X1 U16997 ( .A(n15301), .ZN(n15306) );
  OAI21_X1 U16998 ( .B1(n15303), .B2(n15334), .A(n15302), .ZN(n15305) );
  AOI211_X1 U16999 ( .C1(n15331), .C2(n15306), .A(n15305), .B(n15304), .ZN(
        n15348) );
  INV_X1 U17000 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n15307) );
  AOI22_X1 U17001 ( .A1(n15341), .A2(n15348), .B1(n15307), .B2(n15339), .ZN(
        P1_U3477) );
  INV_X1 U17002 ( .A(n15314), .ZN(n15316) );
  AOI21_X1 U17003 ( .B1(n15310), .B2(n15309), .A(n15308), .ZN(n15311) );
  OAI211_X1 U17004 ( .C1(n15314), .C2(n15313), .A(n15312), .B(n15311), .ZN(
        n15315) );
  AOI21_X1 U17005 ( .B1(n15317), .B2(n15316), .A(n15315), .ZN(n15350) );
  INV_X1 U17006 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n15318) );
  AOI22_X1 U17007 ( .A1(n15341), .A2(n15350), .B1(n15318), .B2(n15339), .ZN(
        P1_U3480) );
  OAI21_X1 U17008 ( .B1(n15320), .B2(n15334), .A(n15319), .ZN(n15322) );
  AOI211_X1 U17009 ( .C1(n15323), .C2(n15337), .A(n15322), .B(n15321), .ZN(
        n15352) );
  INV_X1 U17010 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n15324) );
  AOI22_X1 U17011 ( .A1(n15341), .A2(n15352), .B1(n15324), .B2(n15339), .ZN(
        P1_U3483) );
  INV_X1 U17012 ( .A(n15325), .ZN(n15330) );
  OAI21_X1 U17013 ( .B1(n15327), .B2(n15334), .A(n15326), .ZN(n15329) );
  AOI211_X1 U17014 ( .C1(n15331), .C2(n15330), .A(n15329), .B(n15328), .ZN(
        n15354) );
  INV_X1 U17015 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n15332) );
  AOI22_X1 U17016 ( .A1(n15341), .A2(n15354), .B1(n15332), .B2(n15339), .ZN(
        P1_U3486) );
  OAI21_X1 U17017 ( .B1(n7465), .B2(n15334), .A(n15333), .ZN(n15336) );
  AOI211_X1 U17018 ( .C1(n15338), .C2(n15337), .A(n15336), .B(n15335), .ZN(
        n15357) );
  INV_X1 U17019 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n15340) );
  AOI22_X1 U17020 ( .A1(n15341), .A2(n15357), .B1(n15340), .B2(n15339), .ZN(
        P1_U3489) );
  AOI22_X1 U17021 ( .A1(n15358), .A2(n15342), .B1(n10551), .B2(n15355), .ZN(
        P1_U3529) );
  AOI22_X1 U17022 ( .A1(n15358), .A2(n15343), .B1(n10550), .B2(n15355), .ZN(
        P1_U3530) );
  AOI22_X1 U17023 ( .A1(n15358), .A2(n15344), .B1(n10557), .B2(n15355), .ZN(
        P1_U3532) );
  AOI22_X1 U17024 ( .A1(n15358), .A2(n15346), .B1(n15345), .B2(n15355), .ZN(
        P1_U3533) );
  AOI22_X1 U17025 ( .A1(n15358), .A2(n15348), .B1(n15347), .B2(n15355), .ZN(
        P1_U3534) );
  AOI22_X1 U17026 ( .A1(n15358), .A2(n15350), .B1(n15349), .B2(n15355), .ZN(
        P1_U3535) );
  AOI22_X1 U17027 ( .A1(n15358), .A2(n15352), .B1(n15351), .B2(n15355), .ZN(
        P1_U3536) );
  AOI22_X1 U17028 ( .A1(n15358), .A2(n15354), .B1(n15353), .B2(n15355), .ZN(
        P1_U3537) );
  AOI22_X1 U17029 ( .A1(n15358), .A2(n15357), .B1(n15356), .B2(n15355), .ZN(
        P1_U3538) );
  NOR2_X1 U17030 ( .A1(n15448), .A2(P2_U3947), .ZN(P2_U3087) );
  OR2_X1 U17031 ( .A1(n15359), .A2(P2_U3088), .ZN(n15389) );
  NAND2_X1 U17032 ( .A1(n15360), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15361) );
  OAI211_X1 U17033 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(P2_STATE_REG_SCAN_IN), 
        .A(n15389), .B(n15361), .ZN(n15372) );
  OAI211_X1 U17034 ( .C1(n15364), .C2(n15363), .A(n15450), .B(n15362), .ZN(
        n15371) );
  AOI211_X1 U17035 ( .C1(n15367), .C2(n15366), .A(n15365), .B(n15375), .ZN(
        n15368) );
  INV_X1 U17036 ( .A(n15368), .ZN(n15370) );
  NAND2_X1 U17037 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(n15448), .ZN(n15369) );
  NAND4_X1 U17038 ( .A1(n15372), .A2(n15371), .A3(n15370), .A4(n15369), .ZN(
        P2_U3217) );
  NAND2_X1 U17039 ( .A1(n15373), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15374) );
  OAI211_X1 U17040 ( .C1(P2_REG3_REG_4__SCAN_IN), .C2(P2_STATE_REG_SCAN_IN), 
        .A(n15389), .B(n15374), .ZN(n15386) );
  AOI211_X1 U17041 ( .C1(n15378), .C2(n15377), .A(n15376), .B(n15375), .ZN(
        n15379) );
  INV_X1 U17042 ( .A(n15379), .ZN(n15385) );
  NAND2_X1 U17043 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(n15448), .ZN(n15384) );
  OAI211_X1 U17044 ( .C1(n15382), .C2(n15381), .A(n15450), .B(n15380), .ZN(
        n15383) );
  NAND4_X1 U17045 ( .A1(n15386), .A2(n15385), .A3(n15384), .A4(n15383), .ZN(
        P2_U3218) );
  NAND2_X1 U17046 ( .A1(n15387), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15388) );
  OAI211_X1 U17047 ( .C1(P2_REG3_REG_10__SCAN_IN), .C2(P2_STATE_REG_SCAN_IN), 
        .A(n15389), .B(n15388), .ZN(n15399) );
  OAI211_X1 U17048 ( .C1(n15392), .C2(n15391), .A(n15390), .B(n15456), .ZN(
        n15398) );
  OAI211_X1 U17049 ( .C1(n15395), .C2(n15394), .A(n15393), .B(n15450), .ZN(
        n15397) );
  NAND2_X1 U17050 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(n15448), .ZN(n15396) );
  NAND4_X1 U17051 ( .A1(n15399), .A2(n15398), .A3(n15397), .A4(n15396), .ZN(
        P2_U3224) );
  NOR2_X1 U17052 ( .A1(n15401), .A2(n15400), .ZN(n15402) );
  AOI211_X1 U17053 ( .C1(n15448), .C2(P2_ADDR_REG_13__SCAN_IN), .A(n15403), 
        .B(n15402), .ZN(n15414) );
  OAI211_X1 U17054 ( .C1(n15406), .C2(n15405), .A(n15404), .B(n15456), .ZN(
        n15413) );
  AOI21_X1 U17055 ( .B1(n15409), .B2(n15408), .A(n15407), .ZN(n15411) );
  NAND2_X1 U17056 ( .A1(n15411), .A2(n15410), .ZN(n15412) );
  NAND3_X1 U17057 ( .A1(n15414), .A2(n15413), .A3(n15412), .ZN(P2_U3227) );
  AOI22_X1 U17058 ( .A1(n15448), .A2(P2_ADDR_REG_14__SCAN_IN), .B1(
        P2_REG3_REG_14__SCAN_IN), .B2(P2_U3088), .ZN(n15424) );
  OAI211_X1 U17059 ( .C1(n15416), .C2(P2_REG2_REG_14__SCAN_IN), .A(n15450), 
        .B(n15415), .ZN(n15423) );
  NAND2_X1 U17060 ( .A1(n15453), .A2(n15417), .ZN(n15422) );
  OAI211_X1 U17061 ( .C1(n15420), .C2(n15419), .A(n15418), .B(n15456), .ZN(
        n15421) );
  NAND4_X1 U17062 ( .A1(n15424), .A2(n15423), .A3(n15422), .A4(n15421), .ZN(
        P2_U3228) );
  AOI21_X1 U17063 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(n15448), .A(n15425), 
        .ZN(n15434) );
  NAND2_X1 U17064 ( .A1(n15453), .A2(n15426), .ZN(n15433) );
  OAI211_X1 U17065 ( .C1(n15428), .C2(P2_REG2_REG_15__SCAN_IN), .A(n15450), 
        .B(n15427), .ZN(n15432) );
  OAI211_X1 U17066 ( .C1(P2_REG1_REG_15__SCAN_IN), .C2(n15430), .A(n15456), 
        .B(n15429), .ZN(n15431) );
  NAND4_X1 U17067 ( .A1(n15434), .A2(n15433), .A3(n15432), .A4(n15431), .ZN(
        P2_U3229) );
  AOI22_X1 U17068 ( .A1(n15448), .A2(P2_ADDR_REG_16__SCAN_IN), .B1(
        P2_REG3_REG_16__SCAN_IN), .B2(P2_U3088), .ZN(n15446) );
  NAND2_X1 U17069 ( .A1(n15453), .A2(n15436), .ZN(n15445) );
  OAI211_X1 U17070 ( .C1(n15439), .C2(n15438), .A(n15450), .B(n15437), .ZN(
        n15444) );
  OAI211_X1 U17071 ( .C1(n15442), .C2(n15441), .A(n15456), .B(n15440), .ZN(
        n15443) );
  NAND4_X1 U17072 ( .A1(n15446), .A2(n15445), .A3(n15444), .A4(n15443), .ZN(
        P2_U3230) );
  AOI21_X1 U17073 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(n15448), .A(n15447), 
        .ZN(n15462) );
  OAI211_X1 U17074 ( .C1(n15452), .C2(n15451), .A(n15450), .B(n15449), .ZN(
        n15461) );
  NAND2_X1 U17075 ( .A1(n15454), .A2(n15453), .ZN(n15460) );
  OAI211_X1 U17076 ( .C1(n15458), .C2(n15457), .A(n15456), .B(n15455), .ZN(
        n15459) );
  NAND4_X1 U17077 ( .A1(n15462), .A2(n15461), .A3(n15460), .A4(n15459), .ZN(
        P2_U3231) );
  AND2_X1 U17078 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n15464), .ZN(P2_U3266) );
  AND2_X1 U17079 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n15464), .ZN(P2_U3267) );
  AND2_X1 U17080 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n15464), .ZN(P2_U3268) );
  AND2_X1 U17081 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n15464), .ZN(P2_U3269) );
  AND2_X1 U17082 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n15464), .ZN(P2_U3270) );
  AND2_X1 U17083 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n15464), .ZN(P2_U3271) );
  AND2_X1 U17084 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n15464), .ZN(P2_U3272) );
  AND2_X1 U17085 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n15464), .ZN(P2_U3273) );
  AND2_X1 U17086 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n15464), .ZN(P2_U3274) );
  AND2_X1 U17087 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n15464), .ZN(P2_U3275) );
  AND2_X1 U17088 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n15464), .ZN(P2_U3276) );
  AND2_X1 U17089 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n15464), .ZN(P2_U3277) );
  AND2_X1 U17090 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n15464), .ZN(P2_U3278) );
  AND2_X1 U17091 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n15464), .ZN(P2_U3279) );
  AND2_X1 U17092 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n15464), .ZN(P2_U3280) );
  AND2_X1 U17093 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n15464), .ZN(P2_U3281) );
  AND2_X1 U17094 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n15464), .ZN(P2_U3282) );
  AND2_X1 U17095 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n15464), .ZN(P2_U3283) );
  AND2_X1 U17096 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n15464), .ZN(P2_U3284) );
  AND2_X1 U17097 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n15464), .ZN(P2_U3285) );
  AND2_X1 U17098 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n15464), .ZN(P2_U3286) );
  AND2_X1 U17099 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n15464), .ZN(P2_U3287) );
  AND2_X1 U17100 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n15464), .ZN(P2_U3288) );
  AND2_X1 U17101 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n15464), .ZN(P2_U3289) );
  AND2_X1 U17102 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n15464), .ZN(P2_U3290) );
  AND2_X1 U17103 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n15464), .ZN(P2_U3291) );
  AND2_X1 U17104 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n15464), .ZN(P2_U3292) );
  AND2_X1 U17105 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n15464), .ZN(P2_U3293) );
  AND2_X1 U17106 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n15464), .ZN(P2_U3294) );
  AND2_X1 U17107 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n15464), .ZN(P2_U3295) );
  OAI21_X1 U17108 ( .B1(n15470), .B2(n15466), .A(n15465), .ZN(P2_U3416) );
  INV_X1 U17109 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n15468) );
  AOI22_X1 U17110 ( .A1(n15470), .A2(n15469), .B1(n15468), .B2(n15467), .ZN(
        P2_U3417) );
  INV_X1 U17111 ( .A(n15511), .ZN(n15519) );
  INV_X1 U17112 ( .A(n15471), .ZN(n15472) );
  AOI211_X1 U17113 ( .C1(n15519), .C2(n15474), .A(n15473), .B(n15472), .ZN(
        n15526) );
  AOI22_X1 U17114 ( .A1(n15524), .A2(n15526), .B1(n7752), .B2(n15523), .ZN(
        P2_U3430) );
  OAI21_X1 U17115 ( .B1(n15476), .B2(n15516), .A(n15475), .ZN(n15478) );
  AOI211_X1 U17116 ( .C1(n15479), .C2(n15491), .A(n15478), .B(n15477), .ZN(
        n15527) );
  AOI22_X1 U17117 ( .A1(n15524), .A2(n15527), .B1(n7805), .B2(n15523), .ZN(
        P2_U3445) );
  NOR2_X1 U17118 ( .A1(n15480), .A2(n15511), .ZN(n15486) );
  NOR2_X1 U17119 ( .A1(n15480), .A2(n11052), .ZN(n15485) );
  OAI21_X1 U17120 ( .B1(n15482), .B2(n15516), .A(n15481), .ZN(n15484) );
  NOR4_X1 U17121 ( .A1(n15486), .A2(n15485), .A3(n15484), .A4(n15483), .ZN(
        n15529) );
  AOI22_X1 U17122 ( .A1(n15524), .A2(n15529), .B1(n7841), .B2(n15523), .ZN(
        P2_U3448) );
  OAI21_X1 U17123 ( .B1(n15488), .B2(n15516), .A(n15487), .ZN(n15490) );
  AOI211_X1 U17124 ( .C1(n15492), .C2(n15491), .A(n15490), .B(n15489), .ZN(
        n15530) );
  AOI22_X1 U17125 ( .A1(n15524), .A2(n15530), .B1(n7862), .B2(n15523), .ZN(
        P2_U3451) );
  OAI21_X1 U17126 ( .B1(n7159), .B2(n15516), .A(n15493), .ZN(n15494) );
  AOI21_X1 U17127 ( .B1(n15496), .B2(n15519), .A(n15494), .ZN(n15498) );
  AOI21_X1 U17128 ( .B1(n15496), .B2(n15514), .A(n15495), .ZN(n15497) );
  AND2_X1 U17129 ( .A1(n15498), .A2(n15497), .ZN(n15532) );
  AOI22_X1 U17130 ( .A1(n15524), .A2(n15532), .B1(n7881), .B2(n15523), .ZN(
        P2_U3454) );
  AOI21_X1 U17131 ( .B1(n11052), .B2(n15511), .A(n15499), .ZN(n15504) );
  NOR2_X1 U17132 ( .A1(n15500), .A2(n15516), .ZN(n15503) );
  NOR4_X1 U17133 ( .A1(n15504), .A2(n15503), .A3(n15502), .A4(n15501), .ZN(
        n15534) );
  AOI22_X1 U17134 ( .A1(n15524), .A2(n15534), .B1(n7898), .B2(n15523), .ZN(
        P2_U3457) );
  INV_X1 U17135 ( .A(n15510), .ZN(n15513) );
  AOI211_X1 U17136 ( .C1(n15508), .C2(n15507), .A(n15506), .B(n15505), .ZN(
        n15509) );
  OAI21_X1 U17137 ( .B1(n15511), .B2(n15510), .A(n15509), .ZN(n15512) );
  AOI21_X1 U17138 ( .B1(n15514), .B2(n15513), .A(n15512), .ZN(n15535) );
  AOI22_X1 U17139 ( .A1(n15524), .A2(n15535), .B1(n7923), .B2(n15523), .ZN(
        P2_U3460) );
  OAI21_X1 U17140 ( .B1(n15517), .B2(n15516), .A(n15515), .ZN(n15518) );
  AOI21_X1 U17141 ( .B1(n15520), .B2(n15519), .A(n15518), .ZN(n15521) );
  AND2_X1 U17142 ( .A1(n15522), .A2(n15521), .ZN(n15538) );
  AOI22_X1 U17143 ( .A1(n15524), .A2(n15538), .B1(n7939), .B2(n15523), .ZN(
        P2_U3463) );
  AOI22_X1 U17144 ( .A1(n15539), .A2(n15526), .B1(n15525), .B2(n15536), .ZN(
        P2_U3499) );
  AOI22_X1 U17145 ( .A1(n15539), .A2(n15527), .B1(n10516), .B2(n15536), .ZN(
        P2_U3504) );
  AOI22_X1 U17146 ( .A1(n15539), .A2(n15529), .B1(n15528), .B2(n15536), .ZN(
        P2_U3505) );
  AOI22_X1 U17147 ( .A1(n15539), .A2(n15530), .B1(n10534), .B2(n15536), .ZN(
        P2_U3506) );
  AOI22_X1 U17148 ( .A1(n15539), .A2(n15532), .B1(n15531), .B2(n15536), .ZN(
        P2_U3507) );
  AOI22_X1 U17149 ( .A1(n15539), .A2(n15534), .B1(n15533), .B2(n15536), .ZN(
        P2_U3508) );
  AOI22_X1 U17150 ( .A1(n15539), .A2(n15535), .B1(n11071), .B2(n15536), .ZN(
        P2_U3509) );
  AOI22_X1 U17151 ( .A1(n15539), .A2(n15538), .B1(n15537), .B2(n15536), .ZN(
        P2_U3510) );
  NOR2_X1 U17152 ( .A1(P3_U3897), .A2(n15623), .ZN(P3_U3150) );
  AOI22_X1 U17153 ( .A1(n15540), .A2(P3_IR_REG_0__SCAN_IN), .B1(
        P3_REG3_REG_0__SCAN_IN), .B2(P3_U3151), .ZN(n15547) );
  NAND3_X1 U17154 ( .A1(n15636), .A2(n15541), .A3(n15611), .ZN(n15545) );
  OAI21_X1 U17155 ( .B1(P3_IR_REG_0__SCAN_IN), .B2(n15543), .A(n15542), .ZN(
        n15544) );
  NAND2_X1 U17156 ( .A1(n15545), .A2(n15544), .ZN(n15546) );
  OAI211_X1 U17157 ( .C1(n15549), .C2(n15548), .A(n15547), .B(n15546), .ZN(
        P3_U3182) );
  AOI21_X1 U17158 ( .B1(n15552), .B2(n15551), .A(n15550), .ZN(n15566) );
  NAND2_X1 U17159 ( .A1(n15554), .A2(n15553), .ZN(n15555) );
  XNOR2_X1 U17160 ( .A(n15556), .B(n15555), .ZN(n15558) );
  OAI22_X1 U17161 ( .A1(n15558), .A2(n15611), .B1(n15557), .B2(n15626), .ZN(
        n15559) );
  AOI211_X1 U17162 ( .C1(P3_ADDR_REG_9__SCAN_IN), .C2(n15623), .A(n15560), .B(
        n15559), .ZN(n15565) );
  OAI21_X1 U17163 ( .B1(P3_REG1_REG_9__SCAN_IN), .B2(n15562), .A(n15561), .ZN(
        n15563) );
  NAND2_X1 U17164 ( .A1(n15563), .A2(n15628), .ZN(n15564) );
  OAI211_X1 U17165 ( .C1(n15566), .C2(n15636), .A(n15565), .B(n15564), .ZN(
        P3_U3191) );
  AOI21_X1 U17166 ( .B1(n8651), .B2(n15568), .A(n15567), .ZN(n15582) );
  OAI21_X1 U17167 ( .B1(P3_REG1_REG_11__SCAN_IN), .B2(n15570), .A(n15569), 
        .ZN(n15575) );
  AOI21_X1 U17168 ( .B1(n15623), .B2(P3_ADDR_REG_11__SCAN_IN), .A(n15571), 
        .ZN(n15572) );
  OAI21_X1 U17169 ( .B1(n15626), .B2(n15573), .A(n15572), .ZN(n15574) );
  AOI21_X1 U17170 ( .B1(n15575), .B2(n15628), .A(n15574), .ZN(n15581) );
  NOR2_X1 U17171 ( .A1(n15577), .A2(n15576), .ZN(n15579) );
  OAI21_X1 U17172 ( .B1(n15579), .B2(n15578), .A(n15630), .ZN(n15580) );
  OAI211_X1 U17173 ( .C1(n15582), .C2(n15636), .A(n15581), .B(n15580), .ZN(
        P3_U3193) );
  AOI21_X1 U17174 ( .B1(n6786), .B2(n15584), .A(n15583), .ZN(n15598) );
  OAI21_X1 U17175 ( .B1(n15587), .B2(n15586), .A(n15585), .ZN(n15592) );
  AOI21_X1 U17176 ( .B1(n15623), .B2(P3_ADDR_REG_12__SCAN_IN), .A(n15588), 
        .ZN(n15589) );
  OAI21_X1 U17177 ( .B1(n15626), .B2(n15590), .A(n15589), .ZN(n15591) );
  AOI21_X1 U17178 ( .B1(n15592), .B2(n15628), .A(n15591), .ZN(n15597) );
  OAI211_X1 U17179 ( .C1(n15595), .C2(n15594), .A(n15593), .B(n15630), .ZN(
        n15596) );
  OAI211_X1 U17180 ( .C1(n15598), .C2(n15636), .A(n15597), .B(n15596), .ZN(
        P3_U3194) );
  AOI21_X1 U17181 ( .B1(n8683), .B2(n15600), .A(n15599), .ZN(n15615) );
  OAI21_X1 U17182 ( .B1(P3_REG1_REG_13__SCAN_IN), .B2(n15602), .A(n15601), 
        .ZN(n15607) );
  AOI21_X1 U17183 ( .B1(n15623), .B2(P3_ADDR_REG_13__SCAN_IN), .A(n15603), 
        .ZN(n15604) );
  OAI21_X1 U17184 ( .B1(n15626), .B2(n15605), .A(n15604), .ZN(n15606) );
  AOI21_X1 U17185 ( .B1(n15607), .B2(n15628), .A(n15606), .ZN(n15614) );
  AOI21_X1 U17186 ( .B1(n15610), .B2(n15609), .A(n15608), .ZN(n15612) );
  OR2_X1 U17187 ( .A1(n15612), .A2(n15611), .ZN(n15613) );
  OAI211_X1 U17188 ( .C1(n15615), .C2(n15636), .A(n15614), .B(n15613), .ZN(
        P3_U3195) );
  AOI21_X1 U17189 ( .B1(n15618), .B2(n15617), .A(n15616), .ZN(n15637) );
  OAI21_X1 U17190 ( .B1(n15621), .B2(n15620), .A(n15619), .ZN(n15629) );
  AOI21_X1 U17191 ( .B1(n15623), .B2(P3_ADDR_REG_14__SCAN_IN), .A(n15622), 
        .ZN(n15624) );
  OAI21_X1 U17192 ( .B1(n15626), .B2(n15625), .A(n15624), .ZN(n15627) );
  AOI21_X1 U17193 ( .B1(n15629), .B2(n15628), .A(n15627), .ZN(n15635) );
  OAI211_X1 U17194 ( .C1(n15633), .C2(n15632), .A(n15631), .B(n15630), .ZN(
        n15634) );
  OAI211_X1 U17195 ( .C1(n15637), .C2(n15636), .A(n15635), .B(n15634), .ZN(
        P3_U3196) );
  XOR2_X1 U17196 ( .A(n15638), .B(n15645), .Z(n15641) );
  AOI222_X1 U17197 ( .A1(n15703), .A2(n15641), .B1(n15640), .B2(n15697), .C1(
        n15639), .C2(n15700), .ZN(n15736) );
  AOI22_X1 U17198 ( .A1(P3_REG2_REG_10__SCAN_IN), .A2(n15714), .B1(n15710), 
        .B2(n15642), .ZN(n15651) );
  INV_X1 U17199 ( .A(n15643), .ZN(n15644) );
  AOI21_X1 U17200 ( .B1(n15646), .B2(n15645), .A(n15644), .ZN(n15740) );
  NOR2_X1 U17201 ( .A1(n15647), .A2(n15730), .ZN(n15738) );
  AOI22_X1 U17202 ( .A1(n15740), .A2(n15649), .B1(n15648), .B2(n15738), .ZN(
        n15650) );
  OAI211_X1 U17203 ( .C1(n15714), .C2(n15736), .A(n15651), .B(n15650), .ZN(
        P3_U3223) );
  INV_X1 U17204 ( .A(n15652), .ZN(n15668) );
  OAI21_X1 U17205 ( .B1(n15668), .B2(n15654), .A(n15653), .ZN(n15655) );
  MUX2_X1 U17206 ( .A(n15655), .B(P3_REG2_REG_7__SCAN_IN), .S(n15714), .Z(
        n15656) );
  AOI21_X1 U17207 ( .B1(n15673), .B2(n15657), .A(n15656), .ZN(n15658) );
  OAI21_X1 U17208 ( .B1(n15659), .B2(n15675), .A(n15658), .ZN(P3_U3226) );
  OAI21_X1 U17209 ( .B1(n15668), .B2(n15661), .A(n15660), .ZN(n15662) );
  MUX2_X1 U17210 ( .A(n15662), .B(P3_REG2_REG_6__SCAN_IN), .S(n15714), .Z(
        n15663) );
  AOI21_X1 U17211 ( .B1(n15673), .B2(n15664), .A(n15663), .ZN(n15665) );
  OAI21_X1 U17212 ( .B1(n15666), .B2(n15675), .A(n15665), .ZN(P3_U3227) );
  OAI21_X1 U17213 ( .B1(n15669), .B2(n15668), .A(n15667), .ZN(n15670) );
  MUX2_X1 U17214 ( .A(P3_REG2_REG_4__SCAN_IN), .B(n15670), .S(n15693), .Z(
        n15671) );
  AOI21_X1 U17215 ( .B1(n15673), .B2(n15672), .A(n15671), .ZN(n15674) );
  OAI21_X1 U17216 ( .B1(n15676), .B2(n15675), .A(n15674), .ZN(P3_U3229) );
  XNOR2_X1 U17217 ( .A(n15677), .B(n15678), .ZN(n15686) );
  OAI21_X1 U17218 ( .B1(n15679), .B2(n15678), .A(n12853), .ZN(n15720) );
  NAND2_X1 U17219 ( .A1(n15720), .A2(n15680), .ZN(n15684) );
  AOI22_X1 U17220 ( .A1(n15700), .A2(n15682), .B1(n15681), .B2(n15697), .ZN(
        n15683) );
  OAI211_X1 U17221 ( .C1(n15686), .C2(n15685), .A(n15684), .B(n15683), .ZN(
        n15718) );
  INV_X1 U17222 ( .A(n15720), .ZN(n15691) );
  NOR2_X1 U17223 ( .A1(n15687), .A2(n15730), .ZN(n15719) );
  INV_X1 U17224 ( .A(n15719), .ZN(n15688) );
  OAI22_X1 U17225 ( .A1(n15691), .A2(n15690), .B1(n15689), .B2(n15688), .ZN(
        n15692) );
  AOI211_X1 U17226 ( .C1(P3_REG3_REG_2__SCAN_IN), .C2(n15710), .A(n15718), .B(
        n15692), .ZN(n15694) );
  AOI22_X1 U17227 ( .A1(n15714), .A2(n8481), .B1(n15694), .B2(n15693), .ZN(
        P3_U3231) );
  NOR2_X1 U17228 ( .A1(n15695), .A2(n15730), .ZN(n15716) );
  XNOR2_X1 U17229 ( .A(n15702), .B(n15696), .ZN(n15709) );
  AOI22_X1 U17230 ( .A1(n15700), .A2(n15699), .B1(n15698), .B2(n15697), .ZN(
        n15706) );
  XNOR2_X1 U17231 ( .A(n15702), .B(n15701), .ZN(n15704) );
  NAND2_X1 U17232 ( .A1(n15704), .A2(n15703), .ZN(n15705) );
  OAI211_X1 U17233 ( .C1(n15709), .C2(n15707), .A(n15706), .B(n15705), .ZN(
        n15715) );
  AOI21_X1 U17234 ( .B1(n15716), .B2(n15708), .A(n15715), .ZN(n15713) );
  INV_X1 U17235 ( .A(n15709), .ZN(n15717) );
  AOI22_X1 U17236 ( .A1(n15717), .A2(n15711), .B1(P3_REG3_REG_1__SCAN_IN), 
        .B2(n15710), .ZN(n15712) );
  OAI221_X1 U17237 ( .B1(n15714), .B2(n15713), .C1(n15693), .C2(n8469), .A(
        n15712), .ZN(P3_U3232) );
  AOI211_X1 U17238 ( .C1(n15734), .C2(n15717), .A(n15716), .B(n15715), .ZN(
        n15744) );
  AOI22_X1 U17239 ( .A1(n15743), .A2(n8470), .B1(n15744), .B2(n15741), .ZN(
        P3_U3393) );
  AOI211_X1 U17240 ( .C1(n15734), .C2(n15720), .A(n15719), .B(n15718), .ZN(
        n15745) );
  AOI22_X1 U17241 ( .A1(n15743), .A2(n8479), .B1(n15745), .B2(n15741), .ZN(
        P3_U3396) );
  INV_X1 U17242 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n15725) );
  AOI21_X1 U17243 ( .B1(n15722), .B2(n15734), .A(n15721), .ZN(n15723) );
  AND2_X1 U17244 ( .A1(n15724), .A2(n15723), .ZN(n15746) );
  AOI22_X1 U17245 ( .A1(n15743), .A2(n15725), .B1(n15746), .B2(n15741), .ZN(
        P3_U3405) );
  INV_X1 U17246 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n15729) );
  AOI211_X1 U17247 ( .C1(n15734), .C2(n15728), .A(n15727), .B(n15726), .ZN(
        n15747) );
  AOI22_X1 U17248 ( .A1(n15743), .A2(n15729), .B1(n15747), .B2(n15741), .ZN(
        P3_U3414) );
  NOR2_X1 U17249 ( .A1(n15731), .A2(n15730), .ZN(n15733) );
  AOI211_X1 U17250 ( .C1(n15735), .C2(n15734), .A(n15733), .B(n15732), .ZN(
        n15748) );
  AOI22_X1 U17251 ( .A1(n15743), .A2(n8599), .B1(n15748), .B2(n15741), .ZN(
        P3_U3417) );
  INV_X1 U17252 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n15742) );
  INV_X1 U17253 ( .A(n15736), .ZN(n15737) );
  AOI211_X1 U17254 ( .C1(n15740), .C2(n15739), .A(n15738), .B(n15737), .ZN(
        n15750) );
  AOI22_X1 U17255 ( .A1(n15743), .A2(n15742), .B1(n15750), .B2(n15741), .ZN(
        P3_U3420) );
  AOI22_X1 U17256 ( .A1(n15751), .A2(n15744), .B1(n11297), .B2(n15749), .ZN(
        P3_U3460) );
  AOI22_X1 U17257 ( .A1(n15751), .A2(n15745), .B1(n10923), .B2(n15749), .ZN(
        P3_U3461) );
  AOI22_X1 U17258 ( .A1(n15751), .A2(n15746), .B1(n8525), .B2(n15749), .ZN(
        P3_U3464) );
  AOI22_X1 U17259 ( .A1(n15751), .A2(n15747), .B1(n8579), .B2(n15749), .ZN(
        P3_U3467) );
  AOI22_X1 U17260 ( .A1(n15751), .A2(n15748), .B1(n8595), .B2(n15749), .ZN(
        P3_U3468) );
  AOI22_X1 U17261 ( .A1(n15751), .A2(n15750), .B1(n8617), .B2(n15749), .ZN(
        P3_U3469) );
  OAI21_X1 U17262 ( .B1(n15754), .B2(n15753), .A(n15752), .ZN(SUB_1596_U59) );
  OAI21_X1 U17263 ( .B1(n15757), .B2(n15756), .A(n15755), .ZN(SUB_1596_U58) );
  XOR2_X1 U17264 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(n15758), .Z(SUB_1596_U53) );
  OAI21_X1 U17265 ( .B1(n15761), .B2(n15760), .A(n15759), .ZN(SUB_1596_U56) );
  AOI21_X1 U17266 ( .B1(n15764), .B2(n15763), .A(n15762), .ZN(n15765) );
  XOR2_X1 U17267 ( .A(P2_ADDR_REG_3__SCAN_IN), .B(n15765), .Z(SUB_1596_U60) );
  AOI21_X1 U17268 ( .B1(n15768), .B2(n15767), .A(n15766), .ZN(SUB_1596_U5) );
  CLKBUF_X1 U7432 ( .A(n13537), .Z(n13485) );
  CLKBUF_X1 U7439 ( .A(n8465), .Z(n6852) );
  CLKBUF_X1 U7478 ( .A(n7775), .Z(n8403) );
  CLKBUF_X1 U7483 ( .A(n11014), .Z(n12644) );
  CLKBUF_X1 U7692 ( .A(n7868), .Z(n6854) );
  XNOR2_X1 U8758 ( .A(n9970), .B(n7222), .ZN(n14908) );
endmodule

