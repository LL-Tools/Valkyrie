

module b14_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, U3352, U3351, U3350, U3349, 
        U3348, U3347, U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, 
        U3338, U3337, U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, 
        U3328, U3327, U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, 
        U3320, U3319, U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, 
        U3310, U3309, U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, 
        U3300, U3299, U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, 
        U3467, U3469, U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, 
        U3487, U3489, U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, 
        U3506, U3507, U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, 
        U3516, U3517, U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, 
        U3526, U3527, U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, 
        U3536, U3537, U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, 
        U3546, U3547, U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, 
        U3284, U3283, U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, 
        U3274, U3273, U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, 
        U3264, U3263, U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, 
        U3255, U3254, U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, 
        U3245, U3244, U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, 
        U3554, U3555, U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, 
        U3564, U3565, U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, 
        U3574, U3575, U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, 
        U3237, U3236, U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, 
        U3227, U3226, U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, 
        U3217, U3216, U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, 
        U4043, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, 
        keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, 
        keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, 
        keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, 
        keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, 
        keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, 
        keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, 
        keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, 
        keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, 
        keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, 
        keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, 
        keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, 
        keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, 
        keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, 
        keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, 
        keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, 
        keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, 
        keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, 
        keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, 
        keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, 
        keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, 
        keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, 
        keyinput125, keyinput126, keyinput127 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148,
         n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158,
         n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168,
         n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178,
         n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188,
         n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198,
         n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208,
         n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218,
         n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228,
         n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238,
         n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248,
         n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258,
         n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268,
         n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278,
         n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288,
         n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298,
         n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308,
         n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318,
         n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328,
         n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338,
         n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348,
         n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358,
         n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368,
         n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378,
         n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388,
         n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398,
         n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408,
         n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418,
         n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428,
         n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438,
         n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448,
         n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458,
         n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468,
         n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478,
         n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488,
         n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498,
         n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508,
         n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518,
         n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528,
         n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538,
         n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548,
         n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558,
         n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568,
         n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578,
         n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588,
         n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598,
         n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608,
         n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618,
         n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628,
         n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638,
         n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648,
         n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658,
         n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668,
         n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678,
         n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688,
         n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698,
         n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708,
         n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718,
         n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728,
         n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738,
         n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748,
         n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758,
         n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768,
         n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778,
         n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788,
         n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798,
         n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808,
         n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818,
         n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828,
         n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838,
         n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848,
         n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858,
         n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868,
         n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878,
         n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888,
         n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898,
         n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908,
         n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918,
         n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928,
         n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938,
         n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948,
         n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958,
         n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968,
         n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978,
         n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988,
         n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998,
         n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008,
         n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018,
         n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028,
         n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038,
         n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048,
         n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058,
         n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068,
         n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078,
         n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088,
         n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098,
         n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108,
         n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118,
         n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128,
         n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138,
         n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148,
         n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158,
         n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168,
         n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178,
         n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188,
         n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
         n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
         n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
         n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
         n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
         n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
         n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258,
         n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268,
         n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278,
         n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288,
         n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298,
         n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308,
         n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318,
         n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328,
         n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338,
         n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348,
         n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358,
         n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368,
         n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378,
         n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388,
         n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398,
         n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408,
         n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418,
         n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428,
         n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438,
         n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448,
         n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458,
         n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468,
         n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478,
         n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488,
         n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498,
         n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508,
         n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518,
         n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528,
         n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538,
         n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548,
         n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558,
         n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568,
         n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578,
         n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588,
         n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598,
         n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608,
         n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618,
         n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628,
         n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638,
         n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648,
         n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658,
         n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668,
         n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678,
         n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688,
         n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698,
         n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708,
         n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718,
         n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728,
         n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738,
         n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748,
         n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758,
         n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768,
         n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778,
         n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788,
         n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798,
         n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808,
         n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818,
         n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828,
         n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838,
         n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848,
         n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858,
         n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868,
         n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878,
         n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888,
         n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898,
         n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908,
         n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918,
         n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928,
         n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938,
         n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948,
         n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958,
         n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968,
         n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978,
         n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988,
         n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
         n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008,
         n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018,
         n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028,
         n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038,
         n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048,
         n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058,
         n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068,
         n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078,
         n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088,
         n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098,
         n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108,
         n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118,
         n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128,
         n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138,
         n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148,
         n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158,
         n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168,
         n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178,
         n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188,
         n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198,
         n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208,
         n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218,
         n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228,
         n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238,
         n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248,
         n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258,
         n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268,
         n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278,
         n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288,
         n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
         n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
         n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
         n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
         n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
         n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
         n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
         n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
         n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
         n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
         n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
         n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
         n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
         n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
         n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
         n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
         n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
         n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
         n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
         n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
         n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
         n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808,
         n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
         n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
         n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838,
         n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
         n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858,
         n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868,
         n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878,
         n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888,
         n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898,
         n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908,
         n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918,
         n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928,
         n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938,
         n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948,
         n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958,
         n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968,
         n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978,
         n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988,
         n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998,
         n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008,
         n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018,
         n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028,
         n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038,
         n5039, n5040, n5041, n5042, n5043;

  INV_X1 U2381 ( .A(n3754), .ZN(n3658) );
  NAND2_X1 U2382 ( .A1(n3358), .A2(n4460), .ZN(n3966) );
  INV_X1 U2383 ( .A(n3327), .ZN(n3403) );
  AND4_X2 U2384 ( .A1(n2714), .A2(n2713), .A3(n2712), .A4(n2711), .ZN(n3354)
         );
  CLKBUF_X2 U2385 ( .A(n2680), .Z(n2860) );
  INV_X1 U2386 ( .A(n3269), .ZN(n3279) );
  NOR2_X1 U2387 ( .A1(n2631), .A2(n2630), .ZN(n2633) );
  INV_X1 U2388 ( .A(n3174), .ZN(n3731) );
  OR2_X1 U2389 ( .A1(n2471), .A2(n3054), .ZN(n2472) );
  NAND2_X1 U2390 ( .A1(n2957), .A2(n4082), .ZN(n3162) );
  INV_X1 U2391 ( .A(n2808), .ZN(n2891) );
  NAND2_X1 U2392 ( .A1(n3015), .A2(n2559), .ZN(n3212) );
  INV_X1 U2394 ( .A(n2765), .ZN(n2335) );
  AND2_X1 U2395 ( .A1(n3614), .A2(n3656), .ZN(n4403) );
  INV_X1 U2396 ( .A(n3354), .ZN(n4460) );
  INV_X1 U2397 ( .A(n4599), .ZN(n3726) );
  XNOR2_X2 U2398 ( .A(n2241), .B(n3195), .ZN(n3192) );
  INV_X2 U2399 ( .A(IR_REG_7__SCAN_IN), .ZN(n2486) );
  NOR3_X2 U2400 ( .A1(n3470), .A2(n2426), .A3(n2425), .ZN(n2424) );
  XNOR2_X2 U2401 ( .A(n2490), .B(n3263), .ZN(n3259) );
  NAND2_X2 U2402 ( .A1(n4339), .A2(n2837), .ZN(n2838) );
  NAND2_X2 U2403 ( .A1(n4355), .A2(n2826), .ZN(n4339) );
  NAND2_X2 U2404 ( .A1(n3279), .A2(n4105), .ZN(n3953) );
  OR2_X2 U2405 ( .A1(n2635), .A2(n2549), .ZN(n2636) );
  NAND3_X2 U2406 ( .A1(n2686), .A2(n2685), .A3(n2684), .ZN(n2909) );
  AND2_X1 U2407 ( .A1(n2683), .A2(n2682), .ZN(n2684) );
  INV_X1 U2408 ( .A(n4565), .ZN(n4381) );
  NAND2_X1 U2409 ( .A1(n4521), .A2(n2359), .ZN(n4248) );
  NAND2_X1 U2410 ( .A1(n2354), .A2(n2353), .ZN(n3573) );
  AND2_X1 U2411 ( .A1(n2790), .A2(n2789), .ZN(n4565) );
  AND2_X1 U2412 ( .A1(n2179), .A2(n2236), .ZN(n3057) );
  INV_X2 U2413 ( .A(n2909), .ZN(n3272) );
  AOI21_X1 U2414 ( .B1(n2967), .B2(n5040), .A(n2962), .ZN(n2963) );
  OR2_X1 U2415 ( .A1(n3628), .A2(n2256), .ZN(n2967) );
  AOI21_X1 U2416 ( .B1(n4498), .B2(n4596), .A(n2211), .ZN(n4875) );
  XNOR2_X1 U2417 ( .A(n4179), .B(n4051), .ZN(n4498) );
  INV_X1 U2418 ( .A(n2240), .ZN(n4985) );
  OAI211_X1 U2419 ( .C1(n3793), .C2(n4441), .A(n3792), .B(n3791), .ZN(n4175)
         );
  NAND2_X1 U2420 ( .A1(n2213), .A2(n2212), .ZN(n2211) );
  XNOR2_X1 U2421 ( .A(n2291), .B(n3789), .ZN(n3793) );
  OR2_X1 U2422 ( .A1(n4154), .A2(n2276), .ZN(n2275) );
  NAND2_X1 U2423 ( .A1(n2316), .A2(n2314), .ZN(n2512) );
  OR2_X1 U2424 ( .A1(n2798), .A2(n4396), .ZN(n2802) );
  NAND2_X1 U2425 ( .A1(n3425), .A2(n2734), .ZN(n2736) );
  NAND2_X1 U2426 ( .A1(n2238), .A2(n2237), .ZN(n3367) );
  NOR2_X1 U2427 ( .A1(n4420), .A2(n4561), .ZN(n3614) );
  OR2_X1 U2428 ( .A1(n3471), .A2(n3480), .ZN(n3470) );
  OR2_X1 U2429 ( .A1(n2481), .A2(n3195), .ZN(n2482) );
  AOI21_X1 U2430 ( .B1(n3447), .B2(n3959), .A(n2253), .ZN(n2252) );
  NAND2_X1 U2431 ( .A1(n2364), .A2(n2180), .ZN(n2360) );
  OAI21_X1 U2432 ( .B1(n2143), .B2(n2365), .A(n3967), .ZN(n2364) );
  OR2_X1 U2433 ( .A1(n3410), .A2(n3320), .ZN(n3413) );
  NAND2_X1 U2434 ( .A1(n3203), .A2(n4599), .ZN(n3941) );
  NAND3_X1 U2435 ( .A1(n2231), .A2(n2233), .A3(n2234), .ZN(n2236) );
  INV_X1 U2436 ( .A(n2723), .ZN(n3341) );
  AND4_X1 U2437 ( .A1(n2702), .A2(n2701), .A3(n2700), .A4(n2699), .ZN(n3327)
         );
  AND4_X1 U2438 ( .A1(n2721), .A2(n2205), .A3(n2722), .A4(n2720), .ZN(n2723)
         );
  NAND2_X1 U2439 ( .A1(n2658), .A2(n2657), .ZN(n4599) );
  AND2_X1 U2440 ( .A1(n2232), .A2(REG1_REG_4__SCAN_IN), .ZN(n2231) );
  NAND2_X1 U2441 ( .A1(n2139), .A2(DATAI_0_), .ZN(n2658) );
  NAND2_X2 U2442 ( .A1(n3162), .A2(n3161), .ZN(n3754) );
  OR2_X1 U2443 ( .A1(n2680), .A2(n4607), .ZN(n2660) );
  AND2_X1 U2444 ( .A1(n2558), .A2(n2567), .ZN(n2996) );
  XNOR2_X1 U2445 ( .A(n2546), .B(IR_REG_25__SCAN_IN), .ZN(n3015) );
  OR2_X1 U2446 ( .A1(n3105), .A2(n2311), .ZN(n2310) );
  XNOR2_X1 U2447 ( .A(n2387), .B(IR_REG_21__SCAN_IN), .ZN(n4082) );
  NAND2_X1 U2448 ( .A1(n2991), .A2(IR_REG_31__SCAN_IN), .ZN(n2206) );
  NAND2_X1 U2449 ( .A1(n2468), .A2(n2463), .ZN(n3110) );
  NAND3_X1 U2450 ( .A1(n4782), .A2(n2447), .A3(n2466), .ZN(n2474) );
  INV_X1 U2451 ( .A(IR_REG_23__SCAN_IN), .ZN(n2561) );
  NOR2_X2 U2452 ( .A1(IR_REG_0__SCAN_IN), .A2(IR_REG_1__SCAN_IN), .ZN(n2466)
         );
  INV_X2 U2453 ( .A(IR_REG_31__SCAN_IN), .ZN(n2549) );
  INV_X1 U2454 ( .A(IR_REG_22__SCAN_IN), .ZN(n4606) );
  NOR2_X1 U2455 ( .A1(IR_REG_19__SCAN_IN), .A2(IR_REG_13__SCAN_IN), .ZN(n2541)
         );
  NOR2_X1 U2456 ( .A1(IR_REG_15__SCAN_IN), .A2(IR_REG_17__SCAN_IN), .ZN(n2540)
         );
  NOR2_X1 U2457 ( .A1(IR_REG_20__SCAN_IN), .A2(IR_REG_16__SCAN_IN), .ZN(n2539)
         );
  NOR2_X1 U2458 ( .A1(IR_REG_4__SCAN_IN), .A2(IR_REG_11__SCAN_IN), .ZN(n2448)
         );
  NOR2_X1 U2459 ( .A1(IR_REG_9__SCAN_IN), .A2(IR_REG_8__SCAN_IN), .ZN(n2450)
         );
  INV_X1 U2460 ( .A(IR_REG_6__SCAN_IN), .ZN(n4624) );
  NOR2_X1 U2461 ( .A1(IR_REG_10__SCAN_IN), .A2(IR_REG_12__SCAN_IN), .ZN(n2449)
         );
  NAND2_X1 U2462 ( .A1(n2194), .A2(n2192), .ZN(n4279) );
  OR2_X1 U2463 ( .A1(n2907), .A2(n3941), .ZN(n3127) );
  INV_X4 U2464 ( .A(IR_REG_5__SCAN_IN), .ZN(n4781) );
  CLKBUF_X1 U2465 ( .A(n2664), .Z(n4602) );
  NAND2_X2 U2466 ( .A1(n3953), .A2(n3951), .ZN(n3271) );
  NAND2_X2 U2467 ( .A1(n3210), .A2(n3269), .ZN(n3951) );
  INV_X1 U2468 ( .A(n2765), .ZN(n2139) );
  XNOR2_X2 U2469 ( .A(n2523), .B(n2791), .ZN(n4969) );
  NAND2_X2 U2470 ( .A1(n2906), .A2(n3942), .ZN(n2907) );
  NAND2_X2 U2471 ( .A1(n2984), .A2(n4477), .ZN(n2906) );
  OAI21_X2 U2472 ( .B1(n4151), .B2(n4759), .A(n2520), .ZN(n4961) );
  XNOR2_X2 U2473 ( .A(n2519), .B(n4938), .ZN(n4151) );
  NAND2_X2 U2474 ( .A1(n2245), .A2(n2244), .ZN(n2519) );
  AOI21_X1 U2475 ( .B1(n4412), .B2(n2804), .A(n2436), .ZN(n2816) );
  OAI22_X2 U2476 ( .A1(n3787), .A2(n4052), .B1(n4495), .B2(n3786), .ZN(n3788)
         );
  BUF_X1 U2477 ( .A(n2708), .Z(n2140) );
  BUF_X2 U2478 ( .A(n2708), .Z(n2141) );
  NAND2_X1 U2479 ( .A1(n3001), .A2(n2639), .ZN(n2708) );
  OR2_X2 U2480 ( .A1(n4229), .A2(n2341), .ZN(n2340) );
  XNOR2_X1 U2481 ( .A(n4945), .B(REG1_REG_1__SCAN_IN), .ZN(n4107) );
  NAND2_X1 U2482 ( .A1(n3199), .A2(n4268), .ZN(n2359) );
  AND2_X1 U2483 ( .A1(n3826), .A2(n2393), .ZN(n2392) );
  NAND2_X1 U2484 ( .A1(n2394), .A2(n3894), .ZN(n2393) );
  INV_X1 U2485 ( .A(n2396), .ZN(n2394) );
  OR2_X1 U2486 ( .A1(n3071), .A2(n4087), .ZN(n3161) );
  INV_X1 U2487 ( .A(n3001), .ZN(n2637) );
  AND2_X1 U2488 ( .A1(n4944), .A2(REG1_REG_2__SCAN_IN), .ZN(n2311) );
  OAI21_X1 U2489 ( .B1(n4140), .B2(n2601), .A(n2602), .ZN(n2604) );
  NAND2_X1 U2490 ( .A1(n4506), .A2(n4208), .ZN(n2351) );
  OR2_X1 U2491 ( .A1(n2483), .A2(IR_REG_6__SCAN_IN), .ZN(n2493) );
  NAND2_X1 U2492 ( .A1(n2466), .A2(n2447), .ZN(n2463) );
  AND2_X1 U2493 ( .A1(n3511), .A2(n2439), .ZN(n2227) );
  INV_X1 U2494 ( .A(n3593), .ZN(n2223) );
  INV_X1 U2495 ( .A(n3162), .ZN(n3070) );
  NAND2_X1 U2496 ( .A1(n2367), .A2(n2366), .ZN(n2368) );
  NAND2_X1 U2497 ( .A1(n2567), .A2(n2165), .ZN(n2367) );
  AND2_X1 U2498 ( .A1(n2227), .A2(n2157), .ZN(n2226) );
  NAND2_X1 U2499 ( .A1(n2144), .A2(n2157), .ZN(n2225) );
  NAND2_X1 U2502 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n2324) );
  NAND2_X1 U2503 ( .A1(n2171), .A2(n3046), .ZN(n2234) );
  NAND2_X1 U2504 ( .A1(n2242), .A2(n2315), .ZN(n2314) );
  NOR2_X1 U2505 ( .A1(n2319), .A2(n2320), .ZN(n2315) );
  OAI21_X1 U2506 ( .B1(n2595), .B2(n2267), .A(n2597), .ZN(n2260) );
  NAND2_X1 U2507 ( .A1(n2275), .A2(n2274), .ZN(n2273) );
  INV_X1 U2508 ( .A(n4956), .ZN(n2274) );
  AND2_X1 U2509 ( .A1(n2890), .A2(n4172), .ZN(n3762) );
  NAND2_X1 U2510 ( .A1(n2286), .A2(REG3_REG_25__SCAN_IN), .ZN(n2874) );
  NAND2_X1 U2511 ( .A1(n2873), .A2(REG3_REG_26__SCAN_IN), .ZN(n2889) );
  INV_X1 U2512 ( .A(n2874), .ZN(n2873) );
  OAI21_X1 U2513 ( .B1(n2193), .B2(n2181), .A(n2199), .ZN(n2192) );
  NAND2_X1 U2514 ( .A1(n2838), .A2(n2190), .ZN(n2194) );
  NAND2_X1 U2515 ( .A1(n2173), .A2(n2756), .ZN(n2353) );
  INV_X1 U2516 ( .A(n2385), .ZN(n2384) );
  AOI21_X1 U2517 ( .B1(n2385), .B2(n2383), .A(n2382), .ZN(n2381) );
  AND2_X1 U2518 ( .A1(n2386), .A2(n3958), .ZN(n2385) );
  OAI21_X1 U2519 ( .B1(n4198), .B2(n4070), .A(n3935), .ZN(n4180) );
  NAND2_X1 U2520 ( .A1(n2505), .A2(IR_REG_31__SCAN_IN), .ZN(n2509) );
  AOI21_X1 U2521 ( .B1(n3294), .B2(n2399), .A(n2398), .ZN(n3356) );
  OAI21_X1 U2522 ( .B1(n2402), .B2(n2184), .A(n2403), .ZN(n2398) );
  NOR2_X1 U2523 ( .A1(n2401), .A2(n2184), .ZN(n2399) );
  INV_X1 U2524 ( .A(n3351), .ZN(n2403) );
  INV_X1 U2525 ( .A(n4272), .ZN(n4099) );
  INV_X1 U2526 ( .A(n3678), .ZN(n3681) );
  INV_X1 U2527 ( .A(IR_REG_2__SCAN_IN), .ZN(n2447) );
  OR2_X1 U2528 ( .A1(n3390), .A2(n3389), .ZN(n2439) );
  NOR2_X1 U2529 ( .A1(n2646), .A2(n3886), .ZN(n2287) );
  AND2_X1 U2530 ( .A1(n3501), .A2(n3500), .ZN(n3525) );
  NAND2_X1 U2531 ( .A1(n2371), .A2(n4008), .ZN(n2369) );
  NOR2_X1 U2532 ( .A1(n2373), .A2(n2372), .ZN(n2371) );
  INV_X1 U2533 ( .A(n2376), .ZN(n2373) );
  INV_X1 U2534 ( .A(n2350), .ZN(n2348) );
  NAND2_X1 U2535 ( .A1(n4237), .A2(n4503), .ZN(n2352) );
  NOR2_X1 U2536 ( .A1(n3988), .A2(n2379), .ZN(n2378) );
  INV_X1 U2537 ( .A(n4055), .ZN(n2379) );
  INV_X1 U2538 ( .A(n2203), .ZN(n2202) );
  OAI21_X1 U2539 ( .B1(n4024), .B2(n2204), .A(n2772), .ZN(n2203) );
  INV_X1 U2540 ( .A(n2764), .ZN(n2204) );
  AND2_X1 U2541 ( .A1(n3338), .A2(n2724), .ZN(n2725) );
  NAND2_X1 U2542 ( .A1(n2723), .A2(n3411), .ZN(n2724) );
  INV_X1 U2543 ( .A(n2717), .ZN(n2622) );
  NOR2_X1 U2544 ( .A1(n2429), .A2(n4503), .ZN(n2428) );
  INV_X1 U2545 ( .A(n2430), .ZN(n2429) );
  AND2_X1 U2546 ( .A1(n2434), .A2(n4341), .ZN(n2433) );
  NOR2_X1 U2547 ( .A1(n4349), .A2(n4380), .ZN(n2434) );
  INV_X1 U2548 ( .A(n4405), .ZN(n3656) );
  NAND2_X1 U2549 ( .A1(n3576), .A2(n4445), .ZN(n2426) );
  INV_X1 U2550 ( .A(n4477), .ZN(n3164) );
  NOR2_X1 U2551 ( .A1(n3203), .A2(n3726), .ZN(n3126) );
  NAND2_X1 U2552 ( .A1(n3126), .A2(n2907), .ZN(n3125) );
  INV_X1 U2553 ( .A(IR_REG_21__SCAN_IN), .ZN(n2543) );
  AND2_X1 U2554 ( .A1(n2419), .A2(n2175), .ZN(n2216) );
  AND2_X1 U2555 ( .A1(n2174), .A2(n3873), .ZN(n2419) );
  NAND2_X1 U2556 ( .A1(n2626), .A2(n2295), .ZN(n2839) );
  INV_X1 U2557 ( .A(n3751), .ZN(n2415) );
  NAND2_X1 U2558 ( .A1(n3232), .A2(n4473), .ZN(n3088) );
  AND2_X1 U2559 ( .A1(n2295), .A2(REG3_REG_20__SCAN_IN), .ZN(n2294) );
  OR2_X1 U2560 ( .A1(n2841), .A2(n3835), .ZN(n2646) );
  NAND2_X1 U2561 ( .A1(n3818), .A2(n3705), .ZN(n3861) );
  AND2_X1 U2562 ( .A1(n3707), .A2(n3708), .ZN(n3705) );
  NAND2_X1 U2563 ( .A1(n2287), .A2(REG3_REG_23__SCAN_IN), .ZN(n2855) );
  OR2_X1 U2564 ( .A1(n3597), .A2(n3777), .ZN(n2409) );
  NAND2_X1 U2565 ( .A1(n3597), .A2(n3777), .ZN(n2408) );
  NOR2_X1 U2566 ( .A1(n3008), .A2(n2940), .ZN(n2559) );
  AND3_X1 U2567 ( .A1(n3069), .A2(n3068), .A3(n3067), .ZN(n3082) );
  OAI21_X1 U2568 ( .B1(n3667), .B2(n3666), .A(n2445), .ZN(n3671) );
  NAND2_X1 U2569 ( .A1(n3657), .A2(n3663), .ZN(n3666) );
  INV_X1 U2570 ( .A(n2437), .ZN(n2404) );
  OR2_X1 U2571 ( .A1(n2437), .A2(n3315), .ZN(n2402) );
  INV_X1 U2572 ( .A(n3728), .ZN(n2416) );
  AND2_X1 U2573 ( .A1(n3652), .A2(n3651), .ZN(n3918) );
  INV_X1 U2574 ( .A(IR_REG_19__SCAN_IN), .ZN(n2532) );
  NOR2_X1 U2575 ( .A1(n3753), .A2(n3073), .ZN(n4089) );
  AND2_X1 U2576 ( .A1(n2863), .A2(n2862), .ZN(n3820) );
  NAND2_X1 U2577 ( .A1(n2575), .A2(n2574), .ZN(n4111) );
  OR2_X1 U2578 ( .A1(n4945), .A2(n2573), .ZN(n2575) );
  NAND2_X1 U2579 ( .A1(n3101), .A2(n2577), .ZN(n2578) );
  INV_X1 U2580 ( .A(n2584), .ZN(n2271) );
  NAND2_X1 U2581 ( .A1(n2583), .A2(n2582), .ZN(n3059) );
  INV_X1 U2582 ( .A(n3060), .ZN(n2269) );
  NAND2_X1 U2583 ( .A1(n3192), .A2(REG1_REG_6__SCAN_IN), .ZN(n3191) );
  INV_X1 U2584 ( .A(n4118), .ZN(n2319) );
  INV_X1 U2585 ( .A(REG1_REG_10__SCAN_IN), .ZN(n2320) );
  NAND2_X1 U2586 ( .A1(n2594), .A2(n3465), .ZN(n2595) );
  XNOR2_X1 U2587 ( .A(n2604), .B(n2603), .ZN(n4155) );
  NAND2_X1 U2588 ( .A1(n2273), .A2(n2185), .ZN(n2298) );
  NAND2_X1 U2589 ( .A1(n4980), .A2(n2283), .ZN(n4991) );
  OR2_X1 U2590 ( .A1(n2609), .A2(REG2_REG_17__SCAN_IN), .ZN(n2283) );
  INV_X1 U2591 ( .A(n2328), .ZN(n2327) );
  INV_X1 U2592 ( .A(n2338), .ZN(n2337) );
  OAI21_X1 U2593 ( .B1(n2343), .B2(n2339), .A(n2162), .ZN(n2338) );
  AND2_X1 U2594 ( .A1(n3999), .A2(n3934), .ZN(n4052) );
  AND2_X1 U2595 ( .A1(n2352), .A2(n2864), .ZN(n2350) );
  NAND2_X1 U2596 ( .A1(n2198), .A2(n2151), .ZN(n2197) );
  OR2_X1 U2597 ( .A1(n4352), .A2(n4341), .ZN(n2837) );
  NAND2_X1 U2598 ( .A1(n2288), .A2(REG3_REG_17__SCAN_IN), .ZN(n2817) );
  INV_X1 U2599 ( .A(n2806), .ZN(n2288) );
  NAND2_X1 U2600 ( .A1(n2626), .A2(REG3_REG_18__SCAN_IN), .ZN(n2828) );
  OR2_X1 U2601 ( .A1(n2801), .A2(n2800), .ZN(n4370) );
  AND2_X1 U2602 ( .A1(n4058), .A2(n4055), .ZN(n4399) );
  NAND2_X1 U2603 ( .A1(n2290), .A2(REG3_REG_15__SCAN_IN), .ZN(n2794) );
  INV_X1 U2604 ( .A(n2792), .ZN(n2290) );
  NAND2_X1 U2605 ( .A1(n2284), .A2(REG3_REG_13__SCAN_IN), .ZN(n2780) );
  INV_X1 U2606 ( .A(n2773), .ZN(n2284) );
  NAND2_X1 U2607 ( .A1(n3573), .A2(n4024), .ZN(n3572) );
  NAND2_X1 U2608 ( .A1(n2624), .A2(REG3_REG_10__SCAN_IN), .ZN(n2758) );
  INV_X1 U2609 ( .A(n2749), .ZN(n2624) );
  NOR2_X1 U2610 ( .A1(n2746), .A2(n2358), .ZN(n2357) );
  INV_X1 U2611 ( .A(n2735), .ZN(n2358) );
  AND2_X1 U2612 ( .A1(n4359), .A2(n3346), .ZN(n3091) );
  NAND2_X1 U2613 ( .A1(n2360), .A2(n2361), .ZN(n2247) );
  NAND2_X1 U2614 ( .A1(n3246), .A2(n2360), .ZN(n2248) );
  NAND2_X1 U2615 ( .A1(n3940), .A2(n3071), .ZN(n2959) );
  AND2_X1 U2616 ( .A1(n4203), .A2(n4584), .ZN(n2258) );
  NOR2_X1 U2617 ( .A1(n2959), .A2(n2958), .ZN(n4359) );
  NAND2_X1 U2618 ( .A1(n4418), .A2(n3571), .ZN(n4596) );
  NAND2_X1 U2619 ( .A1(n2567), .A2(IR_REG_31__SCAN_IN), .ZN(n2571) );
  INV_X1 U2620 ( .A(n2631), .ZN(n2420) );
  INV_X1 U2621 ( .A(IR_REG_11__SCAN_IN), .ZN(n2508) );
  INV_X1 U2622 ( .A(IR_REG_9__SCAN_IN), .ZN(n2498) );
  INV_X1 U2623 ( .A(IR_REG_10__SCAN_IN), .ZN(n4794) );
  XNOR2_X1 U2624 ( .A(n2494), .B(IR_REG_9__SCAN_IN), .ZN(n3364) );
  INV_X1 U2625 ( .A(IR_REG_8__SCAN_IN), .ZN(n2491) );
  INV_X1 U2626 ( .A(IR_REG_1__SCAN_IN), .ZN(n2322) );
  INV_X1 U2627 ( .A(IR_REG_0__SCAN_IN), .ZN(n2323) );
  NAND2_X1 U2628 ( .A1(n3223), .A2(n3224), .ZN(n3236) );
  OAI21_X1 U2629 ( .B1(n3391), .B2(n2222), .A(n2219), .ZN(n3776) );
  AOI21_X1 U2630 ( .B1(n2221), .B2(n2220), .A(n2183), .ZN(n2219) );
  INV_X1 U2631 ( .A(n2226), .ZN(n2220) );
  AND2_X1 U2632 ( .A1(n2874), .A2(n2867), .ZN(n4220) );
  NAND2_X1 U2633 ( .A1(n3236), .A2(n3235), .ZN(n3294) );
  AND2_X1 U2634 ( .A1(n3237), .A2(n3234), .ZN(n3235) );
  INV_X1 U2635 ( .A(n3499), .ZN(n3535) );
  INV_X1 U2636 ( .A(n4269), .ZN(n4313) );
  INV_X1 U2637 ( .A(n3923), .ZN(n3906) );
  OAI21_X1 U2638 ( .B1(n4172), .B2(n2808), .A(n2905), .ZN(n4097) );
  NAND2_X1 U2639 ( .A1(n2880), .A2(n2879), .ZN(n4493) );
  OR2_X1 U2640 ( .A1(n4209), .A2(n2681), .ZN(n2880) );
  NOR2_X1 U2641 ( .A1(n4106), .A2(n2442), .ZN(n3107) );
  NAND2_X1 U2642 ( .A1(n3046), .A2(n2472), .ZN(n2473) );
  NAND2_X1 U2643 ( .A1(n2490), .A2(n2590), .ZN(n2237) );
  NAND2_X1 U2644 ( .A1(n3259), .A2(REG1_REG_8__SCAN_IN), .ZN(n2238) );
  NAND2_X1 U2645 ( .A1(n2600), .A2(n2599), .ZN(n4140) );
  XNOR2_X1 U2646 ( .A(n2298), .B(n5024), .ZN(n4967) );
  NAND2_X1 U2647 ( .A1(n4967), .A2(n4966), .ZN(n4965) );
  OR2_X1 U2648 ( .A1(n4953), .A2(n3182), .ZN(n5000) );
  INV_X1 U2649 ( .A(n4984), .ZN(n2239) );
  INV_X1 U2650 ( .A(n4970), .ZN(n4996) );
  NOR2_X1 U2651 ( .A1(n4991), .A2(n4992), .ZN(n4990) );
  NAND2_X1 U2652 ( .A1(n2301), .A2(n4974), .ZN(n2300) );
  NAND2_X1 U2653 ( .A1(n4991), .A2(n4992), .ZN(n2301) );
  OAI21_X1 U2654 ( .B1(n5000), .B2(n5021), .A(n2304), .ZN(n2303) );
  AOI21_X1 U2655 ( .B1(n4994), .B2(ADDR_REG_18__SCAN_IN), .A(n4993), .ZN(n2304) );
  OR2_X1 U2656 ( .A1(n4953), .A2(n4950), .ZN(n4970) );
  AND2_X1 U2657 ( .A1(n2935), .A2(n4595), .ZN(n3628) );
  XNOR2_X1 U2658 ( .A(n2249), .B(n4052), .ZN(n2935) );
  NAND2_X1 U2659 ( .A1(n2250), .A2(n2374), .ZN(n2249) );
  INV_X1 U2660 ( .A(n2293), .ZN(n2374) );
  INV_X1 U2661 ( .A(n3997), .ZN(n4203) );
  AND2_X1 U2662 ( .A1(n2898), .A2(n2897), .ZN(n4495) );
  NAND2_X1 U2663 ( .A1(n2336), .A2(n2343), .ZN(n4179) );
  XNOR2_X1 U2664 ( .A(n2476), .B(n4781), .ZN(n3063) );
  INV_X1 U2665 ( .A(n3369), .ZN(n2280) );
  NOR2_X1 U2666 ( .A1(n2280), .A2(n4463), .ZN(n2278) );
  INV_X1 U2667 ( .A(n3953), .ZN(n2365) );
  NOR2_X1 U2668 ( .A1(n2827), .A2(n2296), .ZN(n2295) );
  OAI21_X1 U2669 ( .B1(n2390), .B2(n2217), .A(n2216), .ZN(n2418) );
  AOI21_X1 U2670 ( .B1(n2392), .B2(n2395), .A(n2170), .ZN(n2389) );
  INV_X1 U2671 ( .A(n3894), .ZN(n2395) );
  INV_X1 U2672 ( .A(n3679), .ZN(n3680) );
  INV_X1 U2673 ( .A(n3289), .ZN(n3735) );
  NOR2_X1 U2674 ( .A1(n2267), .A2(n2747), .ZN(n2265) );
  INV_X1 U2675 ( .A(n4143), .ZN(n2307) );
  NOR2_X1 U2676 ( .A1(n2307), .A2(n4792), .ZN(n2243) );
  INV_X1 U2677 ( .A(n2886), .ZN(n2339) );
  NAND2_X1 U2678 ( .A1(n2342), .A2(n2886), .ZN(n2341) );
  INV_X1 U2679 ( .A(n2345), .ZN(n2342) );
  NOR2_X1 U2680 ( .A1(n4181), .A2(n2377), .ZN(n2376) );
  INV_X1 U2681 ( .A(n3935), .ZN(n2377) );
  OR2_X1 U2682 ( .A1(n4237), .A2(n4222), .ZN(n4196) );
  NOR2_X1 U2683 ( .A1(n2195), .A2(n2197), .ZN(n2190) );
  INV_X1 U2684 ( .A(n2199), .ZN(n2195) );
  INV_X1 U2685 ( .A(n2152), .ZN(n2193) );
  INV_X1 U2686 ( .A(n2817), .ZN(n2626) );
  AND2_X1 U2687 ( .A1(n2357), .A2(n2756), .ZN(n2355) );
  INV_X1 U2688 ( .A(n3974), .ZN(n2253) );
  NAND2_X1 U2689 ( .A1(n2911), .A2(n3966), .ZN(n2386) );
  INV_X1 U2690 ( .A(n3969), .ZN(n2382) );
  NAND2_X1 U2691 ( .A1(n2180), .A2(n2362), .ZN(n2361) );
  INV_X1 U2692 ( .A(n2365), .ZN(n2362) );
  NOR2_X1 U2693 ( .A1(n4240), .A2(n2431), .ZN(n2430) );
  INV_X1 U2694 ( .A(IR_REG_27__SCAN_IN), .ZN(n2628) );
  INV_X1 U2695 ( .A(IR_REG_24__SCAN_IN), .ZN(n2545) );
  INV_X1 U2696 ( .A(IR_REG_15__SCAN_IN), .ZN(n2460) );
  INV_X1 U2697 ( .A(IR_REG_13__SCAN_IN), .ZN(n4627) );
  OR2_X1 U2698 ( .A1(n2493), .A2(n2492), .ZN(n2497) );
  INV_X1 U2699 ( .A(n2153), .ZN(n2401) );
  INV_X1 U2700 ( .A(n2287), .ZN(n2847) );
  NOR2_X1 U2701 ( .A1(n3893), .A2(n2397), .ZN(n2396) );
  INV_X1 U2702 ( .A(n3670), .ZN(n2397) );
  INV_X1 U2703 ( .A(REG3_REG_19__SCAN_IN), .ZN(n2827) );
  NAND2_X1 U2704 ( .A1(n2622), .A2(n2163), .ZN(n2749) );
  AND2_X1 U2705 ( .A1(REG3_REG_8__SCAN_IN), .A2(REG3_REG_9__SCAN_IN), .ZN(
        n2623) );
  NAND2_X1 U2706 ( .A1(n2622), .A2(n2155), .ZN(n2739) );
  NAND2_X1 U2707 ( .A1(n2390), .A2(n2389), .ZN(n3870) );
  NAND2_X1 U2708 ( .A1(n3870), .A2(n3871), .ZN(n3869) );
  AND2_X1 U2709 ( .A1(n3177), .A2(n3176), .ZN(n3178) );
  NAND2_X1 U2710 ( .A1(n2625), .A2(REG3_REG_14__SCAN_IN), .ZN(n2792) );
  INV_X1 U2711 ( .A(n2780), .ZN(n2625) );
  OR2_X1 U2712 ( .A1(n3840), .A2(n3841), .ZN(n3915) );
  AND2_X1 U2713 ( .A1(n3840), .A2(n3841), .ZN(n3916) );
  OR2_X1 U2714 ( .A1(n2141), .A2(n3116), .ZN(n2678) );
  INV_X1 U2715 ( .A(n4124), .ZN(n2267) );
  AND2_X1 U2716 ( .A1(n2605), .A2(n4938), .ZN(n2276) );
  NAND2_X1 U2717 ( .A1(n4998), .A2(n2329), .ZN(n2328) );
  INV_X1 U2718 ( .A(n2526), .ZN(n2329) );
  NAND2_X1 U2719 ( .A1(n2292), .A2(n2164), .ZN(n2291) );
  OR2_X1 U2720 ( .A1(n2369), .A2(n4215), .ZN(n2292) );
  NAND2_X1 U2721 ( .A1(n3934), .A2(n2293), .ZN(n2370) );
  OAI21_X1 U2722 ( .B1(n4181), .B2(n2375), .A(n3998), .ZN(n2293) );
  NAND2_X1 U2723 ( .A1(n4070), .A2(n3935), .ZN(n2375) );
  NAND2_X1 U2724 ( .A1(n4198), .A2(n2376), .ZN(n2250) );
  AND2_X1 U2725 ( .A1(n2885), .A2(n2884), .ZN(n3997) );
  NAND2_X1 U2726 ( .A1(n2349), .A2(n2351), .ZN(n2345) );
  OR2_X1 U2727 ( .A1(n2347), .A2(n2344), .ZN(n2343) );
  INV_X1 U2728 ( .A(n2351), .ZN(n2344) );
  AOI21_X1 U2729 ( .B1(n2348), .B2(n2349), .A(n2159), .ZN(n2347) );
  NAND2_X1 U2730 ( .A1(n2380), .A2(n2378), .ZN(n4328) );
  NAND2_X1 U2731 ( .A1(n2289), .A2(REG3_REG_16__SCAN_IN), .ZN(n2806) );
  INV_X1 U2732 ( .A(n2794), .ZN(n2289) );
  NAND2_X1 U2733 ( .A1(n2920), .A2(n3983), .ZN(n4413) );
  NAND2_X1 U2734 ( .A1(n2285), .A2(REG3_REG_12__SCAN_IN), .ZN(n2773) );
  INV_X1 U2735 ( .A(n2766), .ZN(n2285) );
  AOI21_X1 U2736 ( .B1(n2202), .B2(n2204), .A(n2166), .ZN(n2200) );
  INV_X1 U2737 ( .A(REG3_REG_11__SCAN_IN), .ZN(n4850) );
  OR2_X1 U2738 ( .A1(n2758), .A2(n4850), .ZN(n2766) );
  AND4_X1 U2739 ( .A1(n2755), .A2(n2754), .A3(n2753), .A4(n2752), .ZN(n3509)
         );
  NAND2_X1 U2740 ( .A1(n2621), .A2(REG3_REG_5__SCAN_IN), .ZN(n2717) );
  OAI21_X1 U2741 ( .B1(n3246), .B2(n2361), .A(n2360), .ZN(n3402) );
  OR2_X1 U2742 ( .A1(n2141), .A2(n2715), .ZN(n2205) );
  NAND2_X1 U2743 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n2696) );
  NAND2_X1 U2744 ( .A1(n3246), .A2(n3950), .ZN(n3277) );
  NAND2_X1 U2745 ( .A1(n3125), .A2(n2665), .ZN(n2968) );
  NAND2_X1 U2746 ( .A1(n3127), .A2(n2906), .ZN(n2972) );
  AOI21_X1 U2747 ( .B1(n2952), .B2(n3027), .A(n3026), .ZN(n3068) );
  NAND2_X1 U2748 ( .A1(n2335), .A2(DATAI_31_), .ZN(n4078) );
  OR2_X1 U2749 ( .A1(n4183), .A2(n3761), .ZN(n3795) );
  NOR2_X1 U2750 ( .A1(n3795), .A2(n3932), .ZN(n4162) );
  NAND2_X1 U2751 ( .A1(n2335), .A2(DATAI_27_), .ZN(n4185) );
  AND2_X1 U2752 ( .A1(n4275), .A2(n2187), .ZN(n4206) );
  INV_X1 U2753 ( .A(n4222), .ZN(n4503) );
  NAND2_X1 U2754 ( .A1(n4275), .A2(n2430), .ZN(n4242) );
  NAND2_X1 U2755 ( .A1(n4275), .A2(n4258), .ZN(n4257) );
  AND2_X1 U2756 ( .A1(n2335), .A2(DATAI_21_), .ZN(n4524) );
  AND2_X1 U2757 ( .A1(n4403), .A2(n2150), .ZN(n4318) );
  NAND2_X1 U2758 ( .A1(n4403), .A2(n2433), .ZN(n4340) );
  NAND2_X1 U2759 ( .A1(n4403), .A2(n2434), .ZN(n4358) );
  NAND2_X1 U2760 ( .A1(n4403), .A2(n4546), .ZN(n4376) );
  NAND2_X1 U2761 ( .A1(n3596), .A2(n4573), .ZN(n2425) );
  NOR3_X1 U2762 ( .A1(n3470), .A2(n4583), .A3(n2955), .ZN(n4446) );
  NOR2_X1 U2763 ( .A1(n3470), .A2(n2955), .ZN(n3568) );
  OR2_X1 U2764 ( .A1(n3413), .A2(n3345), .ZN(n3430) );
  NOR2_X1 U2765 ( .A1(n3430), .A2(n4458), .ZN(n3451) );
  AND2_X1 U2766 ( .A1(n3726), .A2(n3306), .ZN(n2421) );
  NOR2_X1 U2767 ( .A1(n2422), .A2(n2423), .ZN(n3307) );
  NAND2_X1 U2768 ( .A1(n2954), .A2(n3164), .ZN(n2422) );
  NAND2_X1 U2769 ( .A1(n3252), .A2(n2954), .ZN(n3268) );
  AND2_X1 U2770 ( .A1(n3164), .A2(n3726), .ZN(n3252) );
  OR2_X1 U2771 ( .A1(n3076), .A2(n4947), .ZN(n4547) );
  INV_X1 U2772 ( .A(n4564), .ZN(n4601) );
  NAND2_X1 U2773 ( .A1(n2939), .A2(n2996), .ZN(n2977) );
  NAND2_X1 U2774 ( .A1(n3212), .A2(n5018), .ZN(n3086) );
  NOR2_X1 U2775 ( .A1(n2452), .A2(IR_REG_26__SCAN_IN), .ZN(n2330) );
  XNOR2_X1 U2776 ( .A(n2564), .B(n4606), .ZN(n3071) );
  INV_X1 U2777 ( .A(IR_REG_20__SCAN_IN), .ZN(n2900) );
  NAND2_X1 U2778 ( .A1(n2899), .A2(IR_REG_31__SCAN_IN), .ZN(n2388) );
  INV_X1 U2779 ( .A(IR_REG_4__SCAN_IN), .ZN(n2475) );
  NAND2_X1 U2780 ( .A1(n2463), .A2(IR_REG_31__SCAN_IN), .ZN(n2470) );
  INV_X1 U2781 ( .A(n2467), .ZN(n2468) );
  OAI22_X1 U2782 ( .A1(n2305), .A2(n2466), .B1(IR_REG_31__SCAN_IN), .B2(
        IR_REG_2__SCAN_IN), .ZN(n2467) );
  NAND2_X1 U2783 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_2__SCAN_IN), .ZN(n2305)
         );
  NAND2_X1 U2784 ( .A1(n2412), .A2(n3904), .ZN(n3752) );
  NAND2_X1 U2785 ( .A1(n2417), .A2(n2413), .ZN(n2412) );
  INV_X1 U2786 ( .A(n2406), .ZN(n2405) );
  OAI21_X1 U2787 ( .B1(n2409), .B2(n2147), .A(n3641), .ZN(n2406) );
  NAND2_X1 U2788 ( .A1(n3701), .A2(n3871), .ZN(n2215) );
  OR2_X1 U2789 ( .A1(n2216), .A2(n2218), .ZN(n2214) );
  AOI21_X1 U2790 ( .B1(n3391), .B2(n2227), .A(n2144), .ZN(n3558) );
  NAND2_X1 U2791 ( .A1(n2391), .A2(n3894), .ZN(n3825) );
  NAND2_X1 U2792 ( .A1(n3671), .A2(n2396), .ZN(n2391) );
  OAI21_X1 U2793 ( .B1(n3730), .B2(n2414), .A(n2148), .ZN(n3775) );
  NAND2_X1 U2794 ( .A1(n2413), .A2(n2411), .ZN(n2410) );
  INV_X1 U2795 ( .A(REG3_REG_21__SCAN_IN), .ZN(n3835) );
  NAND2_X1 U2796 ( .A1(n3869), .A2(n3873), .ZN(n3813) );
  AND2_X1 U2797 ( .A1(n2813), .A2(n2812), .ZN(n4391) );
  NAND2_X1 U2798 ( .A1(n3294), .A2(n3293), .ZN(n3316) );
  OR2_X1 U2799 ( .A1(n4363), .A2(n2808), .ZN(n2824) );
  AND2_X1 U2800 ( .A1(n2872), .A2(n2871), .ZN(n4201) );
  AND2_X1 U2801 ( .A1(n2866), .A2(n2856), .ZN(n4243) );
  AND4_X1 U2802 ( .A1(n2733), .A2(n2732), .A3(n2731), .A4(n2730), .ZN(n3534)
         );
  NAND2_X1 U2803 ( .A1(n2407), .A2(n2408), .ZN(n3642) );
  NAND2_X1 U2804 ( .A1(n3776), .A2(n2409), .ZN(n2407) );
  AND2_X1 U2805 ( .A1(n2853), .A2(n2852), .ZN(n4272) );
  NAND2_X1 U2806 ( .A1(n3216), .A2(n3215), .ZN(n3889) );
  NAND2_X1 U2807 ( .A1(n2224), .A2(n2225), .ZN(n3594) );
  NAND2_X1 U2808 ( .A1(n3391), .A2(n2226), .ZN(n2224) );
  AND2_X1 U2809 ( .A1(n2835), .A2(n2834), .ZN(n4352) );
  OR2_X1 U2810 ( .A1(n3184), .A2(n3084), .ZN(n3898) );
  NAND2_X1 U2811 ( .A1(n3671), .A2(n3670), .ZN(n3892) );
  NAND2_X1 U2812 ( .A1(n2400), .A2(n2402), .ZN(n3352) );
  NAND2_X1 U2813 ( .A1(n3294), .A2(n2153), .ZN(n2400) );
  INV_X1 U2814 ( .A(n3908), .ZN(n3925) );
  OR2_X1 U2815 ( .A1(n3184), .A2(n3183), .ZN(n3923) );
  INV_X1 U2816 ( .A(n3913), .ZN(n3920) );
  INV_X1 U2817 ( .A(n3898), .ZN(n3927) );
  INV_X1 U2818 ( .A(n3889), .ZN(n3931) );
  AND2_X1 U2819 ( .A1(n2534), .A2(n2899), .ZN(n4087) );
  INV_X1 U2820 ( .A(n4495), .ZN(n4098) );
  INV_X1 U2821 ( .A(n4201), .ZN(n4237) );
  INV_X1 U2822 ( .A(n3820), .ZN(n4504) );
  NAND2_X1 U2823 ( .A1(n2651), .A2(n2650), .ZN(n4269) );
  NAND2_X1 U2824 ( .A1(n2846), .A2(n2845), .ZN(n4525) );
  INV_X1 U2825 ( .A(n4352), .ZN(n4311) );
  INV_X1 U2826 ( .A(n4391), .ZN(n4350) );
  OAI211_X1 U2827 ( .C1(n2860), .C2(n4922), .A(n2796), .B(n2795), .ZN(n4570)
         );
  OR2_X1 U2828 ( .A1(n2778), .A2(n2777), .ZN(n4586) );
  INV_X1 U2829 ( .A(n4100), .ZN(n4103) );
  INV_X1 U2830 ( .A(n3534), .ZN(n4104) );
  NOR2_X1 U2831 ( .A1(n3107), .A2(n3106), .ZN(n3105) );
  XNOR2_X1 U2832 ( .A(n2578), .B(n3054), .ZN(n3045) );
  INV_X1 U2833 ( .A(n2308), .ZN(n3048) );
  AOI21_X1 U2834 ( .B1(n3059), .B2(n2146), .A(n2167), .ZN(n2272) );
  INV_X1 U2835 ( .A(n2241), .ZN(n2481) );
  NAND2_X1 U2836 ( .A1(n2279), .A2(n2592), .ZN(n3368) );
  NAND2_X1 U2837 ( .A1(n3260), .A2(REG2_REG_8__SCAN_IN), .ZN(n2279) );
  NAND2_X1 U2838 ( .A1(n3367), .A2(n2496), .ZN(n3365) );
  NAND2_X1 U2839 ( .A1(n2318), .A2(n2502), .ZN(n4119) );
  INV_X1 U2840 ( .A(n2502), .ZN(n2313) );
  AOI21_X1 U2841 ( .B1(n2502), .B2(n2320), .A(n2319), .ZN(n2312) );
  NAND2_X1 U2842 ( .A1(n2266), .A2(n2595), .ZN(n4125) );
  NAND2_X1 U2843 ( .A1(n3461), .A2(REG2_REG_10__SCAN_IN), .ZN(n2266) );
  OAI21_X1 U2844 ( .B1(n3461), .B2(n2262), .A(n2261), .ZN(n4123) );
  INV_X1 U2845 ( .A(n2595), .ZN(n2262) );
  AOI21_X1 U2846 ( .B1(n2595), .B2(n2747), .A(n2267), .ZN(n2261) );
  NAND2_X1 U2847 ( .A1(n2514), .A2(n2513), .ZN(n4144) );
  NAND2_X1 U2848 ( .A1(n4129), .A2(REG1_REG_12__SCAN_IN), .ZN(n2514) );
  NAND2_X1 U2849 ( .A1(n4144), .A2(n4143), .ZN(n4142) );
  NAND2_X1 U2850 ( .A1(n4961), .A2(n4962), .ZN(n4960) );
  INV_X1 U2851 ( .A(n2273), .ZN(n4955) );
  INV_X1 U2852 ( .A(n2275), .ZN(n4957) );
  INV_X1 U2853 ( .A(n2298), .ZN(n2607) );
  AOI21_X1 U2854 ( .B1(n2327), .B2(n4984), .A(n2186), .ZN(n2326) );
  OR2_X1 U2855 ( .A1(n2889), .A2(n2888), .ZN(n4172) );
  INV_X1 U2856 ( .A(n2213), .ZN(n4497) );
  NAND2_X1 U2857 ( .A1(n2346), .A2(n2349), .ZN(n4195) );
  NAND2_X1 U2858 ( .A1(n4229), .A2(n2350), .ZN(n2346) );
  INV_X1 U2859 ( .A(n4524), .ZN(n4300) );
  NAND2_X1 U2860 ( .A1(n2191), .A2(n2152), .ZN(n4284) );
  OR2_X1 U2861 ( .A1(n2196), .A2(n2197), .ZN(n2191) );
  INV_X1 U2862 ( .A(n2838), .ZN(n2196) );
  NAND2_X1 U2863 ( .A1(n2380), .A2(n4055), .ZN(n4367) );
  NAND2_X1 U2864 ( .A1(n3572), .A2(n2764), .ZN(n3547) );
  INV_X1 U2865 ( .A(n4585), .ZN(n3781) );
  NAND2_X1 U2866 ( .A1(n2356), .A2(n2745), .ZN(n3468) );
  NAND2_X1 U2867 ( .A1(n2736), .A2(n2357), .ZN(n2356) );
  OAI21_X1 U2868 ( .B1(n3448), .B2(n3447), .A(n3959), .ZN(n3469) );
  NAND2_X1 U2869 ( .A1(n4484), .A2(n3091), .ZN(n4449) );
  NAND2_X1 U2870 ( .A1(n2363), .A2(n3953), .ZN(n3303) );
  NAND2_X1 U2871 ( .A1(n3246), .A2(n2143), .ZN(n2363) );
  INV_X1 U2872 ( .A(n4449), .ZN(n4480) );
  OR2_X1 U2873 ( .A1(n3086), .A2(n2982), .ZN(n4461) );
  OR2_X1 U2874 ( .A1(n2141), .A2(n2469), .ZN(n2654) );
  INV_X1 U2875 ( .A(n3379), .ZN(n4475) );
  AND2_X1 U2876 ( .A1(n4484), .A2(n3337), .ZN(n4467) );
  INV_X1 U2877 ( .A(n2959), .ZN(n4600) );
  AND2_X1 U2878 ( .A1(n5043), .A2(n4359), .ZN(n4559) );
  OAI21_X1 U2879 ( .B1(n3630), .B2(n4543), .A(n2257), .ZN(n2256) );
  NOR2_X1 U2880 ( .A1(n2936), .A2(n2258), .ZN(n2257) );
  INV_X1 U2881 ( .A(n4496), .ZN(n2212) );
  AND2_X1 U2882 ( .A1(n5040), .A2(n4359), .ZN(n4918) );
  INV_X1 U2883 ( .A(IR_REG_30__SCAN_IN), .ZN(n2992) );
  NAND2_X1 U2884 ( .A1(n2440), .A2(IR_REG_31__SCAN_IN), .ZN(n2546) );
  INV_X1 U2885 ( .A(n2957), .ZN(n2958) );
  INV_X1 U2886 ( .A(n4087), .ZN(n3346) );
  XNOR2_X1 U2887 ( .A(n2515), .B(IR_REG_13__SCAN_IN), .ZN(n4939) );
  XNOR2_X1 U2888 ( .A(n2511), .B(IR_REG_12__SCAN_IN), .ZN(n4940) );
  XNOR2_X1 U2889 ( .A(n2509), .B(n2508), .ZN(n4120) );
  XNOR2_X1 U2890 ( .A(n2500), .B(n4794), .ZN(n3018) );
  XNOR2_X1 U2891 ( .A(n2489), .B(n2491), .ZN(n3263) );
  XNOR2_X1 U2892 ( .A(n2487), .B(IR_REG_7__SCAN_IN), .ZN(n4941) );
  NAND2_X1 U2893 ( .A1(n2323), .A2(IR_REG_1__SCAN_IN), .ZN(n2228) );
  INV_X1 U2894 ( .A(n2321), .ZN(n3055) );
  INV_X1 U2895 ( .A(n2303), .ZN(n2302) );
  OR2_X1 U2896 ( .A1(n2300), .A2(n4990), .ZN(n2299) );
  NAND2_X1 U2897 ( .A1(n2255), .A2(n2254), .ZN(U3546) );
  NOR2_X1 U2898 ( .A1(n2154), .A2(n2966), .ZN(n2254) );
  NAND2_X1 U2899 ( .A1(n2967), .A2(n5043), .ZN(n2255) );
  NOR2_X1 U2900 ( .A1(n5043), .A2(n2965), .ZN(n2966) );
  OAI21_X1 U2901 ( .B1(n4875), .B2(n2210), .A(n2207), .ZN(U3545) );
  AND2_X1 U2902 ( .A1(n2209), .A2(n2208), .ZN(n2207) );
  NAND2_X1 U2903 ( .A1(n2210), .A2(REG1_REG_27__SCAN_IN), .ZN(n2208) );
  OR2_X1 U2904 ( .A1(n4878), .A2(n4594), .ZN(n2209) );
  AND2_X1 U2905 ( .A1(n3950), .A2(n3951), .ZN(n2143) );
  INV_X1 U2906 ( .A(n3753), .ZN(n3232) );
  NAND2_X1 U2907 ( .A1(n2446), .A2(n3510), .ZN(n2144) );
  AND2_X1 U2908 ( .A1(n3820), .A2(n4235), .ZN(n2145) );
  NOR2_X1 U2909 ( .A1(n4942), .A2(n2269), .ZN(n2146) );
  INV_X1 U2910 ( .A(n2474), .ZN(n2331) );
  NAND2_X1 U2911 ( .A1(n2408), .A2(n2182), .ZN(n2147) );
  AND2_X1 U2912 ( .A1(n2169), .A2(n2410), .ZN(n2148) );
  AND2_X1 U2913 ( .A1(n2378), .A2(n2259), .ZN(n2149) );
  NAND2_X1 U2914 ( .A1(n2172), .A2(n2352), .ZN(n2349) );
  INV_X1 U2915 ( .A(n3701), .ZN(n2218) );
  OR2_X1 U2916 ( .A1(n2156), .A2(n3815), .ZN(n3701) );
  AND2_X1 U2917 ( .A1(n2644), .A2(n2643), .ZN(n4527) );
  AND2_X1 U2918 ( .A1(n2433), .A2(n4320), .ZN(n2150) );
  AND2_X1 U2919 ( .A1(n3945), .A2(n3948), .ZN(n2908) );
  NAND2_X1 U2920 ( .A1(n4388), .A2(n4399), .ZN(n2380) );
  OR2_X1 U2921 ( .A1(n4311), .A2(n4040), .ZN(n2151) );
  NAND3_X1 U2922 ( .A1(n2420), .A2(n2331), .A3(n2330), .ZN(n2567) );
  XNOR2_X1 U2923 ( .A(n2388), .B(n2900), .ZN(n2957) );
  XNOR2_X1 U2924 ( .A(n4203), .B(n4185), .ZN(n4181) );
  OR2_X1 U2925 ( .A1(n4037), .A2(n4036), .ZN(n2152) );
  AND2_X1 U2926 ( .A1(n2404), .A2(n3293), .ZN(n2153) );
  NOR2_X1 U2927 ( .A1(n3626), .A2(n4594), .ZN(n2154) );
  AND2_X1 U2928 ( .A1(REG3_REG_6__SCAN_IN), .A2(REG3_REG_7__SCAN_IN), .ZN(
        n2155) );
  CLKBUF_X3 U2929 ( .A(n2681), .Z(n2808) );
  INV_X1 U2930 ( .A(n3054), .ZN(n2309) );
  OR2_X1 U2931 ( .A1(n3816), .A2(n3817), .ZN(n2156) );
  NAND2_X1 U2932 ( .A1(n3513), .A2(n3512), .ZN(n2157) );
  INV_X1 U2933 ( .A(IR_REG_29__SCAN_IN), .ZN(n2634) );
  INV_X1 U2934 ( .A(IR_REG_28__SCAN_IN), .ZN(n2568) );
  MUX2_X1 U2935 ( .A(DATAI_4_), .B(n4943), .S(n2765), .Z(n3269) );
  NAND2_X1 U2936 ( .A1(n2420), .A2(n2632), .ZN(n2557) );
  INV_X1 U2937 ( .A(n3576), .ZN(n2955) );
  AND2_X1 U2938 ( .A1(n4201), .A2(n4222), .ZN(n2158) );
  AND2_X1 U2939 ( .A1(n4493), .A2(n3907), .ZN(n2159) );
  NAND2_X1 U2940 ( .A1(n3509), .A2(n3562), .ZN(n2160) );
  NAND2_X1 U2941 ( .A1(n2477), .A2(REG1_REG_5__SCAN_IN), .ZN(n2161) );
  OR2_X1 U2942 ( .A1(n3997), .A2(n4185), .ZN(n2162) );
  AND2_X1 U2943 ( .A1(n2155), .A2(n2623), .ZN(n2163) );
  AND2_X1 U2944 ( .A1(n2370), .A2(n3999), .ZN(n2164) );
  AND2_X1 U2945 ( .A1(IR_REG_28__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .ZN(n2165)
         );
  AND2_X1 U2946 ( .A1(n3596), .A2(n4436), .ZN(n2166) );
  INV_X1 U2947 ( .A(REG3_REG_13__SCAN_IN), .ZN(n3607) );
  NOR2_X1 U2948 ( .A1(n4942), .A2(n2584), .ZN(n2167) );
  NAND2_X1 U2949 ( .A1(n2380), .A2(n2149), .ZN(n2168) );
  NAND2_X1 U2950 ( .A1(n4275), .A2(n2428), .ZN(n2432) );
  INV_X1 U2951 ( .A(n4583), .ZN(n3596) );
  INV_X1 U2952 ( .A(n2222), .ZN(n2221) );
  NAND2_X1 U2953 ( .A1(n2225), .A2(n2223), .ZN(n2222) );
  INV_X1 U2954 ( .A(n3934), .ZN(n2372) );
  AND2_X1 U2955 ( .A1(n2415), .A2(n3904), .ZN(n2169) );
  AND2_X1 U2956 ( .A1(n3681), .A2(n3680), .ZN(n2170) );
  INV_X1 U2957 ( .A(n2286), .ZN(n2866) );
  NOR2_X1 U2958 ( .A1(n2855), .A2(n4822), .ZN(n2286) );
  AND2_X1 U2959 ( .A1(n2472), .A2(n3119), .ZN(n2171) );
  OR2_X1 U2960 ( .A1(n2158), .A2(n2145), .ZN(n2172) );
  NAND2_X1 U2961 ( .A1(n2745), .A2(n2160), .ZN(n2173) );
  INV_X1 U2962 ( .A(IR_REG_3__SCAN_IN), .ZN(n4782) );
  NOR2_X1 U2963 ( .A1(n3814), .A2(n2156), .ZN(n2174) );
  OR2_X1 U2964 ( .A1(n2389), .A2(n2217), .ZN(n2175) );
  AND2_X1 U2965 ( .A1(n2149), .A2(n4056), .ZN(n2176) );
  NAND2_X1 U2966 ( .A1(n2622), .A2(REG3_REG_6__SCAN_IN), .ZN(n2177) );
  AND2_X1 U2967 ( .A1(n3701), .A2(n3707), .ZN(n2178) );
  NAND2_X1 U2968 ( .A1(n2473), .A2(n4943), .ZN(n2179) );
  INV_X1 U2969 ( .A(n5043), .ZN(n2210) );
  INV_X1 U2970 ( .A(n3987), .ZN(n2259) );
  NAND2_X1 U2971 ( .A1(n3306), .A2(n3403), .ZN(n2180) );
  INV_X1 U2972 ( .A(n3966), .ZN(n2383) );
  INV_X1 U2973 ( .A(n3729), .ZN(n2411) );
  AND2_X1 U2974 ( .A1(n3391), .A2(n2439), .ZN(n3526) );
  INV_X1 U2975 ( .A(n2427), .ZN(n4448) );
  NOR3_X1 U2976 ( .A1(n3470), .A2(n2426), .A3(n4583), .ZN(n2427) );
  INV_X1 U2977 ( .A(n3871), .ZN(n2217) );
  INV_X1 U2978 ( .A(n4334), .ZN(n4549) );
  AND2_X1 U2979 ( .A1(n2824), .A2(n2823), .ZN(n4334) );
  AND2_X1 U2980 ( .A1(n4269), .A2(n4524), .ZN(n2181) );
  INV_X1 U2981 ( .A(REG3_REG_15__SCAN_IN), .ZN(n3922) );
  INV_X1 U2982 ( .A(n2414), .ZN(n2413) );
  NAND2_X1 U2983 ( .A1(n3903), .A2(n2416), .ZN(n2414) );
  INV_X1 U2984 ( .A(n4341), .ZN(n4040) );
  NAND2_X1 U2985 ( .A1(n2201), .A2(n2200), .ZN(n4443) );
  INV_X1 U2986 ( .A(REG3_REG_18__SCAN_IN), .ZN(n2296) );
  INV_X1 U2987 ( .A(REG3_REG_20__SCAN_IN), .ZN(n2297) );
  AND2_X2 U2988 ( .A1(n2981), .A2(n2964), .ZN(n5040) );
  NAND2_X1 U2989 ( .A1(n2335), .A2(DATAI_23_), .ZN(n4258) );
  INV_X1 U2990 ( .A(n4258), .ZN(n2431) );
  OR2_X1 U2991 ( .A1(n3602), .A2(n3601), .ZN(n2182) );
  AND2_X1 U2992 ( .A1(n3516), .A2(n3515), .ZN(n2183) );
  AND2_X1 U2993 ( .A1(n3322), .A2(n3321), .ZN(n2184) );
  AND2_X1 U2994 ( .A1(n2335), .A2(DATAI_20_), .ZN(n4310) );
  INV_X1 U2995 ( .A(n4268), .ZN(n4273) );
  INV_X1 U2996 ( .A(n3907), .ZN(n4208) );
  AND2_X1 U2997 ( .A1(n2335), .A2(DATAI_26_), .ZN(n3907) );
  NAND2_X1 U2998 ( .A1(n2797), .A2(REG2_REG_15__SCAN_IN), .ZN(n2185) );
  INV_X1 U2999 ( .A(REG3_REG_23__SCAN_IN), .ZN(n4668) );
  NOR2_X1 U3000 ( .A1(n5021), .A2(n2821), .ZN(n2186) );
  AND2_X1 U3001 ( .A1(n2428), .A2(n4208), .ZN(n2187) );
  INV_X1 U3002 ( .A(DATAI_1_), .ZN(n2333) );
  OAI21_X2 U3003 ( .B1(n3152), .B2(REG1_REG_7__SCAN_IN), .A(n4941), .ZN(n2485)
         );
  INV_X1 U3004 ( .A(n2310), .ZN(n2471) );
  NAND2_X1 U3005 ( .A1(n2235), .A2(n4943), .ZN(n2232) );
  NOR2_X1 U3006 ( .A1(n4986), .A2(n2526), .ZN(n4997) );
  OAI21_X1 U3007 ( .B1(n2502), .B2(n2319), .A(n2507), .ZN(n2317) );
  NAND2_X1 U3008 ( .A1(n4965), .A2(n2608), .ZN(n4979) );
  NAND2_X1 U3009 ( .A1(n3153), .A2(n2589), .ZN(n2591) );
  NOR2_X1 U3010 ( .A1(n4155), .A2(n4772), .ZN(n4154) );
  NOR2_X1 U3011 ( .A1(n4990), .A2(n2282), .ZN(n2281) );
  XNOR2_X1 U3012 ( .A(n2281), .B(n2610), .ZN(n2618) );
  INV_X1 U3013 ( .A(n2189), .ZN(n2188) );
  OR2_X2 U3014 ( .A1(n4182), .A2(n4441), .ZN(n2213) );
  NAND3_X2 U3015 ( .A1(n2656), .A2(n2655), .A3(n2654), .ZN(n4473) );
  NAND2_X2 U3016 ( .A1(n3191), .A2(n2482), .ZN(n3152) );
  NOR2_X1 U3017 ( .A1(n4969), .A2(REG1_REG_16__SCAN_IN), .ZN(n4968) );
  INV_X1 U3018 ( .A(n2317), .ZN(n2316) );
  NAND2_X2 U3019 ( .A1(n2485), .A2(n2484), .ZN(n2490) );
  NAND2_X2 U3020 ( .A1(n3365), .A2(n2438), .ZN(n2501) );
  NAND2_X1 U3021 ( .A1(n2268), .A2(n2272), .ZN(n3190) );
  NAND2_X1 U3022 ( .A1(n4111), .A2(n4112), .ZN(n4110) );
  NAND2_X1 U3023 ( .A1(n2264), .A2(n2263), .ZN(n2598) );
  NAND2_X1 U3024 ( .A1(n2277), .A2(n2188), .ZN(n2594) );
  OAI21_X1 U3025 ( .B1(n2592), .B2(n2280), .A(n2593), .ZN(n2189) );
  NAND2_X1 U3026 ( .A1(n2838), .A2(n2151), .ZN(n4306) );
  INV_X1 U3027 ( .A(n4037), .ZN(n2198) );
  NAND2_X1 U3028 ( .A1(n4313), .A2(n4300), .ZN(n2199) );
  NAND2_X1 U3029 ( .A1(n3573), .A2(n2202), .ZN(n2201) );
  INV_X2 U3030 ( .A(n2140), .ZN(n2659) );
  XNOR2_X2 U3031 ( .A(n2206), .B(n2992), .ZN(n2639) );
  XNOR2_X2 U3032 ( .A(n2636), .B(IR_REG_29__SCAN_IN), .ZN(n3001) );
  NOR2_X4 U3033 ( .A1(n2474), .A2(n2452), .ZN(n2632) );
  OAI21_X2 U3034 ( .B1(n2390), .B2(n2215), .A(n2214), .ZN(n3818) );
  INV_X2 U3035 ( .A(n4473), .ZN(n3203) );
  INV_X2 U3036 ( .A(n2680), .ZN(n3037) );
  NAND2_X2 U3037 ( .A1(n2637), .A2(n2639), .ZN(n2680) );
  NOR2_X1 U3038 ( .A1(n4107), .A2(n2324), .ZN(n4106) );
  NAND3_X2 U3039 ( .A1(n2230), .A2(n2229), .A3(n2228), .ZN(n4945) );
  NAND3_X1 U3040 ( .A1(n2322), .A2(IR_REG_31__SCAN_IN), .A3(IR_REG_0__SCAN_IN), 
        .ZN(n2229) );
  NAND2_X1 U3041 ( .A1(n2549), .A2(IR_REG_1__SCAN_IN), .ZN(n2230) );
  INV_X1 U3042 ( .A(n2472), .ZN(n2235) );
  OR2_X2 U3043 ( .A1(n3046), .A2(n3119), .ZN(n2233) );
  NAND3_X1 U3044 ( .A1(n2234), .A2(n2233), .A3(n2232), .ZN(n3117) );
  INV_X1 U3045 ( .A(n2236), .ZN(n3115) );
  AND2_X2 U3046 ( .A1(n2240), .A2(n2239), .ZN(n4986) );
  OR2_X2 U3047 ( .A1(n4968), .A2(n2524), .ZN(n2240) );
  XNOR2_X2 U3048 ( .A(n2310), .B(n3054), .ZN(n2308) );
  NAND2_X2 U3049 ( .A1(n2321), .A2(n2161), .ZN(n2241) );
  NAND2_X1 U3050 ( .A1(n2242), .A2(REG1_REG_10__SCAN_IN), .ZN(n2318) );
  OAI21_X1 U3051 ( .B1(n2313), .B2(n2242), .A(n2312), .ZN(n4117) );
  XNOR2_X1 U3052 ( .A(n2242), .B(REG1_REG_10__SCAN_IN), .ZN(n3467) );
  XNOR2_X2 U3053 ( .A(n2501), .B(n3018), .ZN(n2242) );
  NAND2_X1 U3054 ( .A1(n4129), .A2(n2243), .ZN(n2245) );
  INV_X1 U3055 ( .A(n2306), .ZN(n2244) );
  NAND2_X2 U3056 ( .A1(n2246), .A2(n3955), .ZN(n3339) );
  NAND3_X1 U3057 ( .A1(n2248), .A2(n2247), .A3(n3968), .ZN(n2246) );
  NAND2_X2 U3058 ( .A1(n3247), .A2(n4014), .ZN(n3246) );
  NOR2_X2 U3059 ( .A1(n4215), .A2(n3937), .ZN(n4198) );
  NAND2_X1 U3060 ( .A1(n3448), .A2(n3959), .ZN(n2251) );
  NAND2_X1 U3061 ( .A1(n2251), .A2(n2252), .ZN(n2913) );
  AND2_X1 U3062 ( .A1(n2632), .A2(n2633), .ZN(n2635) );
  NAND3_X1 U3063 ( .A1(n2632), .A2(n2633), .A3(n2634), .ZN(n2991) );
  NAND2_X1 U3064 ( .A1(n2380), .A2(n2176), .ZN(n4288) );
  NAND2_X1 U3065 ( .A1(n3461), .A2(n2265), .ZN(n2264) );
  INV_X1 U3066 ( .A(n2260), .ZN(n2263) );
  NAND2_X1 U3067 ( .A1(n3059), .A2(n3060), .ZN(n3058) );
  NAND2_X1 U3068 ( .A1(n3058), .A2(n2270), .ZN(n2268) );
  NAND2_X1 U3069 ( .A1(n3058), .A2(n2584), .ZN(n2585) );
  NAND2_X1 U3070 ( .A1(n3190), .A2(REG2_REG_6__SCAN_IN), .ZN(n2587) );
  NOR2_X1 U3071 ( .A1(n3195), .A2(n2271), .ZN(n2270) );
  NAND2_X1 U3072 ( .A1(n3260), .A2(n2278), .ZN(n2277) );
  AND2_X1 U3073 ( .A1(n2825), .A2(REG2_REG_18__SCAN_IN), .ZN(n2282) );
  NAND2_X1 U3074 ( .A1(n2626), .A2(n2294), .ZN(n2841) );
  XNOR2_X2 U3075 ( .A(n2591), .B(n3263), .ZN(n3260) );
  NAND2_X1 U3076 ( .A1(n3155), .A2(n3154), .ZN(n3153) );
  NAND3_X1 U3077 ( .A1(n4999), .A2(n2302), .A3(n2299), .ZN(U3258) );
  NAND2_X2 U3078 ( .A1(n4960), .A2(n2522), .ZN(n2523) );
  OAI21_X1 U3079 ( .B1(n2513), .B2(n2307), .A(n2516), .ZN(n2306) );
  NAND2_X2 U3080 ( .A1(n2308), .A2(REG1_REG_3__SCAN_IN), .ZN(n3046) );
  OR2_X2 U3081 ( .A1(n3057), .A2(n3056), .ZN(n2321) );
  NAND2_X1 U3082 ( .A1(n4985), .A2(n2327), .ZN(n2325) );
  NAND2_X1 U3083 ( .A1(n2325), .A2(n2326), .ZN(n2538) );
  OR2_X2 U3084 ( .A1(n4986), .A2(n2328), .ZN(n4995) );
  XNOR2_X2 U3085 ( .A(n2594), .B(n3018), .ZN(n3461) );
  NAND3_X1 U3086 ( .A1(n2968), .A2(n2690), .A3(n3243), .ZN(n2693) );
  AND2_X1 U3087 ( .A1(n2688), .A2(n3271), .ZN(n2690) );
  OAI21_X2 U3088 ( .B1(n2765), .B2(n2333), .A(n2332), .ZN(n4477) );
  NAND2_X1 U3089 ( .A1(n2765), .A2(n4945), .ZN(n2332) );
  OAI21_X1 U3090 ( .B1(n2765), .B2(DATAI_2_), .A(n2334), .ZN(n3251) );
  NAND2_X1 U3091 ( .A1(n2765), .A2(n3110), .ZN(n2334) );
  MUX2_X1 U3092 ( .A(n2687), .B(n3054), .S(n2765), .Z(n3378) );
  MUX2_X1 U3093 ( .A(DATAI_6_), .B(n4942), .S(n2765), .Z(n3320) );
  MUX2_X1 U3094 ( .A(n2703), .B(n3063), .S(n2765), .Z(n3306) );
  MUX2_X1 U3095 ( .A(n2797), .B(DATAI_15_), .S(n2335), .Z(n4561) );
  MUX2_X1 U3096 ( .A(n4941), .B(DATAI_7_), .S(n2335), .Z(n3345) );
  MUX2_X1 U3097 ( .A(n2836), .B(n3346), .S(n2765), .Z(n4341) );
  MUX2_X1 U3098 ( .A(n2791), .B(DATAI_16_), .S(n2335), .Z(n4405) );
  MUX2_X1 U3099 ( .A(n3364), .B(DATAI_9_), .S(n2335), .Z(n3499) );
  MUX2_X1 U3100 ( .A(n3263), .B(n3010), .S(n2335), .Z(n3428) );
  MUX2_X1 U3101 ( .A(n5022), .B(n2814), .S(n2335), .Z(n4546) );
  MUX2_X1 U3102 ( .A(n3018), .B(n3019), .S(n2335), .Z(n3562) );
  AND2_X4 U3103 ( .A1(n2368), .A2(n2569), .ZN(n2765) );
  OR2_X1 U3104 ( .A1(n4229), .A2(n2345), .ZN(n2336) );
  AOI21_X1 U3105 ( .B1(n4229), .B2(n2864), .A(n2145), .ZN(n4214) );
  AND2_X2 U3106 ( .A1(n2340), .A2(n2337), .ZN(n3787) );
  NAND2_X1 U3107 ( .A1(n2736), .A2(n2355), .ZN(n2354) );
  NAND2_X1 U3108 ( .A1(n2736), .A2(n2735), .ZN(n3450) );
  NAND2_X2 U3109 ( .A1(n4279), .A2(n4278), .ZN(n4521) );
  NAND2_X1 U3110 ( .A1(n2571), .A2(n2628), .ZN(n2366) );
  OAI21_X1 U3111 ( .B1(n3339), .B2(n2384), .A(n2381), .ZN(n3448) );
  OAI21_X1 U3112 ( .B1(n3339), .B2(n2911), .A(n3966), .ZN(n3424) );
  OAI21_X1 U3113 ( .B1(n2566), .B2(n2565), .A(IR_REG_31__SCAN_IN), .ZN(n2387)
         );
  NAND2_X1 U3114 ( .A1(n2533), .A2(n2532), .ZN(n2899) );
  NAND2_X1 U3115 ( .A1(n3671), .A2(n2392), .ZN(n2390) );
  NAND2_X2 U3116 ( .A1(n3356), .A2(n3355), .ZN(n3391) );
  OAI21_X2 U3117 ( .B1(n3776), .B2(n2147), .A(n2405), .ZN(n3805) );
  NAND2_X1 U3118 ( .A1(n3805), .A2(n3644), .ZN(n3646) );
  NAND2_X1 U3119 ( .A1(n3730), .A2(n3729), .ZN(n2417) );
  AND2_X1 U3120 ( .A1(n2417), .A2(n2416), .ZN(n3902) );
  NAND2_X1 U3121 ( .A1(n2418), .A2(n2178), .ZN(n3710) );
  NAND2_X1 U3122 ( .A1(n3279), .A2(n3726), .ZN(n2423) );
  NAND4_X1 U3123 ( .A1(n2954), .A2(n3164), .A3(n3279), .A4(n2421), .ZN(n3410)
         );
  INV_X1 U3124 ( .A(n2424), .ZN(n4420) );
  INV_X1 U3125 ( .A(n2432), .ZN(n4218) );
  OR2_X1 U3126 ( .A1(n3753), .A2(n3379), .ZN(n3173) );
  AND2_X1 U3127 ( .A1(n3008), .A2(n2940), .ZN(n3026) );
  XOR2_X1 U3128 ( .A(n4078), .B(n4161), .Z(n3640) );
  NAND2_X4 U3129 ( .A1(n3070), .A2(n3212), .ZN(n3753) );
  NAND2_X1 U3130 ( .A1(n2552), .A2(n2440), .ZN(n3008) );
  NAND2_X1 U3131 ( .A1(n4206), .A2(n4185), .ZN(n4183) );
  INV_X2 U3132 ( .A(n2664), .ZN(n2984) );
  NAND4_X2 U3133 ( .A1(n2663), .A2(n2662), .A3(n2661), .A4(n2660), .ZN(n2664)
         );
  OAI21_X1 U3134 ( .B1(n4162), .B2(n4164), .A(n4161), .ZN(n4874) );
  NAND2_X1 U3135 ( .A1(n4162), .A2(n4164), .ZN(n4161) );
  AOI22_X2 U3136 ( .A1(n4248), .A2(n2854), .B1(n2431), .B2(n4099), .ZN(n4229)
         );
  AOI21_X2 U3137 ( .B1(n2779), .B2(n2444), .A(n2443), .ZN(n4412) );
  INV_X1 U3138 ( .A(n4484), .ZN(n4386) );
  AND2_X1 U3139 ( .A1(n2545), .A2(n2561), .ZN(n2435) );
  NOR2_X1 U3140 ( .A1(n2803), .A2(n4369), .ZN(n2436) );
  AND2_X1 U3141 ( .A1(n3314), .A2(n3313), .ZN(n2437) );
  OR2_X1 U3142 ( .A1(n3375), .A2(n4838), .ZN(n2438) );
  NAND2_X1 U3143 ( .A1(n2547), .A2(n2435), .ZN(n2440) );
  INV_X1 U3144 ( .A(n3015), .ZN(n2937) );
  INV_X1 U3145 ( .A(IR_REG_25__SCAN_IN), .ZN(n2553) );
  INV_X1 U3146 ( .A(n3988), .ZN(n2925) );
  INV_X1 U3147 ( .A(REG2_REG_1__SCAN_IN), .ZN(n2573) );
  AND4_X1 U31480 ( .A1(n2554), .A2(n4606), .A3(n2561), .A4(n2553), .ZN(n2441)
         );
  AND2_X1 U31490 ( .A1(n4945), .A2(REG1_REG_1__SCAN_IN), .ZN(n2442) );
  AND2_X1 U3150 ( .A1(n4439), .A2(n4586), .ZN(n2443) );
  OR2_X1 U3151 ( .A1(n4439), .A2(n4586), .ZN(n2444) );
  AND3_X1 U3152 ( .A1(n3665), .A2(n3850), .A3(n3664), .ZN(n2445) );
  AND2_X1 U3153 ( .A1(n3506), .A2(n3505), .ZN(n2446) );
  INV_X1 U3154 ( .A(n3918), .ZN(n3653) );
  INV_X1 U3155 ( .A(IR_REG_26__SCAN_IN), .ZN(n2629) );
  NAND2_X1 U3156 ( .A1(n3654), .A2(n3653), .ZN(n3657) );
  AND2_X1 U3157 ( .A1(n2543), .A2(n2555), .ZN(n2544) );
  INV_X1 U3158 ( .A(n3559), .ZN(n3510) );
  INV_X1 U3159 ( .A(n3853), .ZN(n3668) );
  INV_X1 U3160 ( .A(n3753), .ZN(n3647) );
  NAND2_X1 U3161 ( .A1(n3669), .A2(n3668), .ZN(n3670) );
  INV_X1 U3162 ( .A(REG3_REG_16__SCAN_IN), .ZN(n4734) );
  OR2_X1 U3163 ( .A1(n3885), .A2(n2808), .ZN(n2644) );
  NAND2_X1 U3164 ( .A1(n3152), .A2(REG1_REG_7__SCAN_IN), .ZN(n2484) );
  INV_X1 U3165 ( .A(n4240), .ZN(n4235) );
  NAND2_X1 U3166 ( .A1(n4334), .A2(n4360), .ZN(n2826) );
  OR2_X1 U3167 ( .A1(n4377), .A2(n2681), .ZN(n2813) );
  AND2_X1 U3168 ( .A1(n4092), .A2(n4082), .ZN(n2941) );
  AND2_X1 U3169 ( .A1(n2335), .A2(DATAI_28_), .ZN(n3761) );
  AND2_X1 U3170 ( .A1(n2335), .A2(DATAI_22_), .ZN(n4268) );
  OR2_X1 U3171 ( .A1(n3604), .A2(n3603), .ZN(n3641) );
  INV_X1 U3172 ( .A(n4459), .ZN(n3478) );
  INV_X1 U3173 ( .A(n3526), .ZN(n3392) );
  INV_X1 U3174 ( .A(n4101), .ZN(n4436) );
  AND3_X1 U3175 ( .A1(n2784), .A2(n2783), .A3(n2782), .ZN(n4437) );
  INV_X1 U3176 ( .A(n2495), .ZN(n2496) );
  AND2_X1 U3177 ( .A1(n4013), .A2(n4250), .ZN(n4285) );
  AND2_X1 U3178 ( .A1(n3950), .A2(n3947), .ZN(n4014) );
  INV_X1 U3179 ( .A(n4547), .ZN(n4584) );
  INV_X1 U3180 ( .A(n2977), .ZN(n2952) );
  AND2_X1 U3181 ( .A1(n2335), .A2(DATAI_24_), .ZN(n4240) );
  INV_X1 U3182 ( .A(n4439), .ZN(n4445) );
  INV_X1 U3183 ( .A(n3562), .ZN(n3480) );
  AND2_X1 U3184 ( .A1(n2934), .A2(n2933), .ZN(n4441) );
  INV_X1 U3185 ( .A(n4582), .ZN(n4572) );
  NAND2_X1 U3186 ( .A1(n3083), .A2(n4461), .ZN(n3908) );
  INV_X1 U3187 ( .A(n3082), .ZN(n3184) );
  INV_X1 U3188 ( .A(n4989), .ZN(n4974) );
  INV_X1 U3189 ( .A(n3428), .ZN(n4458) );
  INV_X1 U3190 ( .A(n4295), .ZN(n4476) );
  NAND2_X1 U3191 ( .A1(n3451), .A2(n3535), .ZN(n3471) );
  NAND2_X1 U3192 ( .A1(n2961), .A2(n2960), .ZN(n2962) );
  INV_X1 U3193 ( .A(n4441), .ZN(n4595) );
  AND3_X1 U3194 ( .A1(n3066), .A2(n2953), .A3(n3067), .ZN(n2964) );
  INV_X1 U3195 ( .A(n2996), .ZN(n2940) );
  INV_X1 U3196 ( .A(n3071), .ZN(n4092) );
  AND2_X1 U3197 ( .A1(n2615), .A2(n2614), .ZN(n4994) );
  OR2_X1 U3198 ( .A1(n3184), .A2(n3087), .ZN(n3913) );
  NAND2_X1 U3199 ( .A1(n3092), .A2(n5018), .ZN(n4100) );
  INV_X1 U3200 ( .A(n3509), .ZN(n4102) );
  OR2_X1 U3201 ( .A1(n4953), .A2(n4090), .ZN(n4989) );
  INV_X1 U3202 ( .A(n4994), .ZN(n4978) );
  XNOR2_X1 U3203 ( .A(n2538), .B(n2537), .ZN(n2620) );
  INV_X1 U3204 ( .A(n4467), .ZN(n4304) );
  INV_X1 U3205 ( .A(n4484), .ZN(n4454) );
  INV_X1 U3206 ( .A(n4559), .ZN(n4594) );
  AND2_X2 U3207 ( .A1(n2964), .A2(n3068), .ZN(n5043) );
  INV_X1 U3208 ( .A(n4918), .ZN(n4936) );
  INV_X1 U3209 ( .A(n5040), .ZN(n5039) );
  INV_X1 U32100 ( .A(n5012), .ZN(n5017) );
  NAND2_X1 U32110 ( .A1(n2977), .A2(n2976), .ZN(n5012) );
  AND2_X1 U32120 ( .A1(n3211), .A2(STATE_REG_SCAN_IN), .ZN(n5018) );
  INV_X1 U32130 ( .A(n2609), .ZN(n5022) );
  INV_X2 U32140 ( .A(n4100), .ZN(U4043) );
  INV_X1 U32150 ( .A(n2963), .ZN(U3514) );
  INV_X2 U32160 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  INV_X1 U32170 ( .A(REG1_REG_18__SCAN_IN), .ZN(n2821) );
  AND3_X2 U32180 ( .A1(n4624), .A2(n2486), .A3(n4781), .ZN(n2451) );
  NAND4_X2 U32190 ( .A1(n2451), .A2(n2450), .A3(n2449), .A4(n2448), .ZN(n2452)
         );
  AND2_X1 U32200 ( .A1(n2632), .A2(n4627), .ZN(n2517) );
  INV_X1 U32210 ( .A(IR_REG_16__SCAN_IN), .ZN(n2453) );
  NAND2_X1 U32220 ( .A1(n2460), .A2(n2453), .ZN(n2527) );
  NOR2_X1 U32230 ( .A1(n2527), .A2(IR_REG_14__SCAN_IN), .ZN(n2454) );
  NAND2_X1 U32240 ( .A1(n2517), .A2(n2454), .ZN(n2456) );
  OAI21_X1 U32250 ( .B1(n2456), .B2(IR_REG_17__SCAN_IN), .A(IR_REG_31__SCAN_IN), .ZN(n2455) );
  XNOR2_X1 U32260 ( .A(n2455), .B(IR_REG_18__SCAN_IN), .ZN(n2825) );
  INV_X1 U32270 ( .A(n2825), .ZN(n5021) );
  AOI22_X1 U32280 ( .A1(REG1_REG_18__SCAN_IN), .A2(n2825), .B1(n5021), .B2(
        n2821), .ZN(n4998) );
  NAND2_X1 U32290 ( .A1(n2456), .A2(IR_REG_31__SCAN_IN), .ZN(n2457) );
  XNOR2_X1 U32300 ( .A(n2457), .B(IR_REG_17__SCAN_IN), .ZN(n2609) );
  NOR2_X1 U32310 ( .A1(n2609), .A2(REG1_REG_17__SCAN_IN), .ZN(n2526) );
  INV_X1 U32320 ( .A(IR_REG_14__SCAN_IN), .ZN(n2458) );
  NAND2_X1 U32330 ( .A1(n2517), .A2(n2458), .ZN(n2459) );
  NAND2_X1 U32340 ( .A1(n2459), .A2(IR_REG_31__SCAN_IN), .ZN(n2521) );
  NAND2_X1 U32350 ( .A1(n2521), .A2(n2460), .ZN(n2461) );
  NAND2_X1 U32360 ( .A1(n2461), .A2(IR_REG_31__SCAN_IN), .ZN(n2462) );
  XNOR2_X1 U32370 ( .A(n2462), .B(IR_REG_16__SCAN_IN), .ZN(n2791) );
  NAND2_X1 U32380 ( .A1(n2470), .A2(n4782), .ZN(n2464) );
  NAND2_X1 U32390 ( .A1(n2464), .A2(IR_REG_31__SCAN_IN), .ZN(n2465) );
  XNOR2_X1 U32400 ( .A(n2465), .B(IR_REG_4__SCAN_IN), .ZN(n4943) );
  INV_X1 U32410 ( .A(n3110), .ZN(n4944) );
  INV_X1 U32420 ( .A(REG1_REG_0__SCAN_IN), .ZN(n2469) );
  XOR2_X1 U32430 ( .A(REG1_REG_2__SCAN_IN), .B(n3110), .Z(n3106) );
  XNOR2_X1 U32440 ( .A(n2470), .B(n4782), .ZN(n3054) );
  INV_X1 U32450 ( .A(REG1_REG_3__SCAN_IN), .ZN(n3049) );
  INV_X1 U32460 ( .A(REG1_REG_4__SCAN_IN), .ZN(n3116) );
  NAND2_X1 U32470 ( .A1(n2331), .A2(n2475), .ZN(n2478) );
  NAND2_X1 U32480 ( .A1(n2478), .A2(IR_REG_31__SCAN_IN), .ZN(n2476) );
  XOR2_X1 U32490 ( .A(REG1_REG_5__SCAN_IN), .B(n3063), .Z(n3056) );
  INV_X1 U32500 ( .A(n3063), .ZN(n2477) );
  INV_X1 U32510 ( .A(n2478), .ZN(n2479) );
  NAND2_X1 U32520 ( .A1(n2479), .A2(n4781), .ZN(n2483) );
  NAND2_X1 U32530 ( .A1(n2483), .A2(IR_REG_31__SCAN_IN), .ZN(n2480) );
  XNOR2_X1 U32540 ( .A(n2480), .B(IR_REG_6__SCAN_IN), .ZN(n4942) );
  INV_X1 U32550 ( .A(n4942), .ZN(n3195) );
  NAND2_X1 U32560 ( .A1(n2493), .A2(IR_REG_31__SCAN_IN), .ZN(n2487) );
  INV_X1 U32570 ( .A(REG1_REG_7__SCAN_IN), .ZN(n2707) );
  NAND2_X1 U32580 ( .A1(n2487), .A2(n2486), .ZN(n2488) );
  NAND2_X1 U32590 ( .A1(n2488), .A2(IR_REG_31__SCAN_IN), .ZN(n2489) );
  INV_X1 U32600 ( .A(n3263), .ZN(n2590) );
  INV_X1 U32610 ( .A(REG1_REG_9__SCAN_IN), .ZN(n4838) );
  NAND2_X1 U32620 ( .A1(n2486), .A2(n2491), .ZN(n2492) );
  NAND2_X1 U32630 ( .A1(n2497), .A2(IR_REG_31__SCAN_IN), .ZN(n2494) );
  MUX2_X1 U32640 ( .A(n4838), .B(REG1_REG_9__SCAN_IN), .S(n3364), .Z(n2495) );
  INV_X1 U32650 ( .A(n3364), .ZN(n3375) );
  INV_X1 U32660 ( .A(n2497), .ZN(n2499) );
  NAND2_X1 U32670 ( .A1(n2499), .A2(n2498), .ZN(n2503) );
  NAND2_X1 U32680 ( .A1(n2503), .A2(IR_REG_31__SCAN_IN), .ZN(n2500) );
  INV_X1 U32690 ( .A(n3018), .ZN(n3465) );
  NAND2_X1 U32700 ( .A1(n2501), .A2(n3465), .ZN(n2502) );
  INV_X1 U32710 ( .A(REG1_REG_11__SCAN_IN), .ZN(n3584) );
  INV_X1 U32720 ( .A(n2503), .ZN(n2504) );
  NAND2_X1 U32730 ( .A1(n2504), .A2(n4794), .ZN(n2505) );
  MUX2_X1 U32740 ( .A(n3584), .B(REG1_REG_11__SCAN_IN), .S(n4120), .Z(n4118)
         );
  INV_X1 U32750 ( .A(n4120), .ZN(n2506) );
  NAND2_X1 U32760 ( .A1(n2506), .A2(REG1_REG_11__SCAN_IN), .ZN(n2507) );
  NAND2_X1 U32770 ( .A1(n2509), .A2(n2508), .ZN(n2510) );
  NAND2_X1 U32780 ( .A1(n2510), .A2(IR_REG_31__SCAN_IN), .ZN(n2511) );
  INV_X1 U32790 ( .A(n4940), .ZN(n4134) );
  XNOR2_X2 U32800 ( .A(n2512), .B(n4134), .ZN(n4129) );
  NAND2_X1 U32810 ( .A1(n2512), .A2(n4940), .ZN(n2513) );
  INV_X1 U32820 ( .A(REG1_REG_13__SCAN_IN), .ZN(n4580) );
  OR2_X1 U32830 ( .A1(n2632), .A2(n2549), .ZN(n2515) );
  MUX2_X1 U32840 ( .A(REG1_REG_13__SCAN_IN), .B(n4580), .S(n4939), .Z(n4143)
         );
  NAND2_X1 U32850 ( .A1(n4939), .A2(REG1_REG_13__SCAN_IN), .ZN(n2516) );
  OR2_X1 U32860 ( .A1(n2517), .A2(n2549), .ZN(n2518) );
  XNOR2_X1 U32870 ( .A(n2518), .B(IR_REG_14__SCAN_IN), .ZN(n4938) );
  INV_X1 U32880 ( .A(REG1_REG_14__SCAN_IN), .ZN(n4759) );
  NAND2_X1 U32890 ( .A1(n2519), .A2(n4938), .ZN(n2520) );
  XNOR2_X1 U32900 ( .A(n2521), .B(IR_REG_15__SCAN_IN), .ZN(n2797) );
  INV_X1 U32910 ( .A(n2797), .ZN(n5026) );
  INV_X1 U32920 ( .A(REG1_REG_15__SCAN_IN), .ZN(n4840) );
  AOI22_X1 U32930 ( .A1(REG1_REG_15__SCAN_IN), .A2(n2797), .B1(n5026), .B2(
        n4840), .ZN(n4962) );
  NAND2_X1 U32940 ( .A1(REG1_REG_15__SCAN_IN), .A2(n2797), .ZN(n2522) );
  NOR2_X1 U32950 ( .A1(n2791), .A2(n2523), .ZN(n2524) );
  INV_X1 U32960 ( .A(REG1_REG_17__SCAN_IN), .ZN(n2525) );
  AOI22_X1 U32970 ( .A1(n2609), .A2(n2525), .B1(REG1_REG_17__SCAN_IN), .B2(
        n5022), .ZN(n4984) );
  INV_X1 U32980 ( .A(REG1_REG_19__SCAN_IN), .ZN(n2535) );
  INV_X1 U32990 ( .A(n2632), .ZN(n2566) );
  NOR2_X2 U33000 ( .A1(IR_REG_18__SCAN_IN), .A2(IR_REG_14__SCAN_IN), .ZN(n2542) );
  INV_X1 U33010 ( .A(n2527), .ZN(n2529) );
  INV_X1 U33020 ( .A(IR_REG_17__SCAN_IN), .ZN(n2528) );
  NAND4_X1 U33030 ( .A1(n2542), .A2(n2529), .A3(n4627), .A4(n2528), .ZN(n2530)
         );
  OAI21_X2 U33040 ( .B1(n2566), .B2(n2530), .A(IR_REG_31__SCAN_IN), .ZN(n2533)
         );
  INV_X1 U33050 ( .A(n2533), .ZN(n2531) );
  NAND2_X1 U33060 ( .A1(n2531), .A2(IR_REG_19__SCAN_IN), .ZN(n2534) );
  MUX2_X1 U33070 ( .A(n2535), .B(REG1_REG_19__SCAN_IN), .S(n4087), .Z(n2536)
         );
  INV_X1 U33080 ( .A(n2536), .ZN(n2537) );
  NAND4_X1 U33090 ( .A1(n2542), .A2(n2541), .A3(n2540), .A4(n2539), .ZN(n2565)
         );
  INV_X1 U33100 ( .A(n2565), .ZN(n2555) );
  NAND2_X1 U33110 ( .A1(n2544), .A2(n2632), .ZN(n2563) );
  NOR2_X2 U33120 ( .A1(n2563), .A2(IR_REG_22__SCAN_IN), .ZN(n2547) );
  INV_X1 U33130 ( .A(n2547), .ZN(n2560) );
  AND2_X1 U33140 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_24__SCAN_IN), .ZN(n2551) );
  NAND2_X1 U33150 ( .A1(IR_REG_23__SCAN_IN), .A2(IR_REG_24__SCAN_IN), .ZN(
        n2548) );
  AOI22_X1 U33160 ( .A1(IR_REG_24__SCAN_IN), .A2(n2549), .B1(n2548), .B2(
        IR_REG_31__SCAN_IN), .ZN(n2550) );
  AOI21_X1 U33170 ( .B1(n2560), .B2(n2551), .A(n2550), .ZN(n2552) );
  NOR2_X1 U33180 ( .A1(IR_REG_21__SCAN_IN), .A2(IR_REG_24__SCAN_IN), .ZN(n2554) );
  NAND2_X1 U33190 ( .A1(n2555), .A2(n2441), .ZN(n2631) );
  NAND2_X1 U33200 ( .A1(n2557), .A2(IR_REG_31__SCAN_IN), .ZN(n2556) );
  MUX2_X1 U33210 ( .A(IR_REG_31__SCAN_IN), .B(n2556), .S(IR_REG_26__SCAN_IN), 
        .Z(n2558) );
  NAND2_X1 U33220 ( .A1(n2560), .A2(IR_REG_31__SCAN_IN), .ZN(n2562) );
  XNOR2_X1 U33230 ( .A(n2562), .B(n2561), .ZN(n3211) );
  OR2_X1 U33240 ( .A1(n3211), .A2(U3149), .ZN(n4095) );
  NAND2_X1 U33250 ( .A1(n3086), .A2(n4095), .ZN(n2615) );
  NAND2_X1 U33260 ( .A1(n2563), .A2(IR_REG_31__SCAN_IN), .ZN(n2564) );
  NAND2_X1 U33270 ( .A1(n2941), .A2(n3211), .ZN(n2570) );
  NAND2_X1 U33280 ( .A1(n2628), .A2(IR_REG_28__SCAN_IN), .ZN(n2569) );
  AND2_X1 U33290 ( .A1(n2570), .A2(n2335), .ZN(n2613) );
  NAND2_X1 U33300 ( .A1(n2615), .A2(n2613), .ZN(n4953) );
  XNOR2_X1 U33310 ( .A(n2571), .B(IR_REG_27__SCAN_IN), .ZN(n4950) );
  INV_X1 U33320 ( .A(REG2_REG_18__SCAN_IN), .ZN(n4820) );
  AOI22_X1 U33330 ( .A1(REG2_REG_18__SCAN_IN), .A2(n5021), .B1(n2825), .B2(
        n4820), .ZN(n4992) );
  NOR2_X1 U33340 ( .A1(n2609), .A2(REG2_REG_17__SCAN_IN), .ZN(n2572) );
  AOI21_X1 U33350 ( .B1(REG2_REG_17__SCAN_IN), .B2(n2609), .A(n2572), .ZN(
        n4981) );
  INV_X1 U33360 ( .A(REG2_REG_2__SCAN_IN), .ZN(n2667) );
  MUX2_X1 U33370 ( .A(n2667), .B(REG2_REG_2__SCAN_IN), .S(n3110), .Z(n3103) );
  NAND2_X1 U33380 ( .A1(n4945), .A2(n2573), .ZN(n2574) );
  AND2_X1 U33390 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n4112) );
  NAND2_X1 U33400 ( .A1(n4945), .A2(REG2_REG_1__SCAN_IN), .ZN(n2576) );
  NAND2_X1 U33410 ( .A1(n4110), .A2(n2576), .ZN(n3102) );
  NAND2_X1 U33420 ( .A1(n3103), .A2(n3102), .ZN(n3101) );
  OR2_X1 U33430 ( .A1(n3110), .A2(n2667), .ZN(n2577) );
  NAND2_X1 U33440 ( .A1(n3045), .A2(REG2_REG_3__SCAN_IN), .ZN(n2580) );
  NAND2_X1 U33450 ( .A1(n2578), .A2(n2309), .ZN(n2579) );
  NAND2_X1 U33460 ( .A1(n2580), .A2(n2579), .ZN(n2581) );
  INV_X1 U33470 ( .A(n4943), .ZN(n3119) );
  XNOR2_X1 U33480 ( .A(n2581), .B(n3119), .ZN(n3114) );
  NAND2_X1 U33490 ( .A1(n3114), .A2(REG2_REG_4__SCAN_IN), .ZN(n2583) );
  NAND2_X1 U33500 ( .A1(n2581), .A2(n4943), .ZN(n2582) );
  INV_X1 U33510 ( .A(REG2_REG_5__SCAN_IN), .ZN(n2694) );
  MUX2_X1 U33520 ( .A(n2694), .B(REG2_REG_5__SCAN_IN), .S(n3063), .Z(n3060) );
  OR2_X1 U3353 ( .A1(n3063), .A2(n2694), .ZN(n2584) );
  NAND2_X1 U33540 ( .A1(n2585), .A2(n4942), .ZN(n2586) );
  NAND2_X1 U3355 ( .A1(n2587), .A2(n2586), .ZN(n3155) );
  INV_X1 U3356 ( .A(REG2_REG_7__SCAN_IN), .ZN(n2588) );
  MUX2_X1 U3357 ( .A(REG2_REG_7__SCAN_IN), .B(n2588), .S(n4941), .Z(n3154) );
  NAND2_X1 U3358 ( .A1(n4941), .A2(REG2_REG_7__SCAN_IN), .ZN(n2589) );
  NAND2_X1 U3359 ( .A1(n2591), .A2(n2590), .ZN(n2592) );
  INV_X1 U3360 ( .A(REG2_REG_9__SCAN_IN), .ZN(n3453) );
  XNOR2_X1 U3361 ( .A(n3364), .B(n3453), .ZN(n3369) );
  NAND2_X1 U3362 ( .A1(n3364), .A2(REG2_REG_9__SCAN_IN), .ZN(n2593) );
  INV_X1 U3363 ( .A(REG2_REG_11__SCAN_IN), .ZN(n2596) );
  MUX2_X1 U3364 ( .A(n2596), .B(REG2_REG_11__SCAN_IN), .S(n4120), .Z(n4124) );
  OR2_X1 U3365 ( .A1(n4120), .A2(n2596), .ZN(n2597) );
  XNOR2_X1 U3366 ( .A(n2598), .B(n4134), .ZN(n4130) );
  NAND2_X1 U3367 ( .A1(n4130), .A2(REG2_REG_12__SCAN_IN), .ZN(n2600) );
  NAND2_X1 U3368 ( .A1(n2598), .A2(n4940), .ZN(n2599) );
  AND2_X1 U3369 ( .A1(n4939), .A2(REG2_REG_13__SCAN_IN), .ZN(n2601) );
  OR2_X1 U3370 ( .A1(n4939), .A2(REG2_REG_13__SCAN_IN), .ZN(n2602) );
  INV_X1 U3371 ( .A(n2604), .ZN(n2605) );
  INV_X1 U3372 ( .A(n4938), .ZN(n2603) );
  INV_X1 U3373 ( .A(REG2_REG_14__SCAN_IN), .ZN(n4772) );
  NAND2_X1 U3374 ( .A1(REG2_REG_15__SCAN_IN), .A2(n2797), .ZN(n2606) );
  OAI21_X1 U3375 ( .B1(REG2_REG_15__SCAN_IN), .B2(n2797), .A(n2606), .ZN(n4956) );
  INV_X1 U3376 ( .A(n2791), .ZN(n5024) );
  NAND2_X1 U3377 ( .A1(n2607), .A2(n5024), .ZN(n2608) );
  INV_X1 U3378 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4966) );
  NAND2_X1 U3379 ( .A1(n4981), .A2(n4979), .ZN(n4980) );
  MUX2_X1 U3380 ( .A(REG2_REG_19__SCAN_IN), .B(n2832), .S(n4087), .Z(n2610) );
  INV_X1 U3381 ( .A(n4950), .ZN(n2612) );
  OAI21_X1 U3382 ( .B1(n2567), .B2(IR_REG_27__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2611) );
  XNOR2_X1 U3383 ( .A(n2611), .B(n2568), .ZN(n4947) );
  OR2_X1 U3384 ( .A1(n2612), .A2(n4947), .ZN(n4090) );
  INV_X1 U3385 ( .A(n4947), .ZN(n3182) );
  NAND2_X1 U3386 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n3827) );
  INV_X1 U3387 ( .A(n2613), .ZN(n2614) );
  NAND2_X1 U3388 ( .A1(n4994), .A2(ADDR_REG_19__SCAN_IN), .ZN(n2616) );
  OAI211_X1 U3389 ( .C1(n5000), .C2(n3346), .A(n3827), .B(n2616), .ZN(n2617)
         );
  AOI21_X1 U3390 ( .B1(n2618), .B2(n4974), .A(n2617), .ZN(n2619) );
  OAI21_X1 U3391 ( .B1(n2620), .B2(n4970), .A(n2619), .ZN(U3259) );
  INV_X1 U3392 ( .A(n2696), .ZN(n2621) );
  INV_X1 U3393 ( .A(REG3_REG_22__SCAN_IN), .ZN(n3886) );
  NAND2_X1 U3394 ( .A1(n2646), .A2(n3886), .ZN(n2627) );
  NAND2_X1 U3395 ( .A1(n2847), .A2(n2627), .ZN(n3885) );
  NAND3_X1 U3396 ( .A1(n2629), .A2(n2628), .A3(n2568), .ZN(n2630) );
  INV_X2 U3397 ( .A(n2639), .ZN(n3004) );
  NAND2_X2 U3398 ( .A1(n3001), .A2(n3004), .ZN(n2681) );
  INV_X1 U3399 ( .A(REG0_REG_22__SCAN_IN), .ZN(n4896) );
  NAND2_X2 U3400 ( .A1(n2637), .A2(n3004), .ZN(n2672) );
  INV_X1 U3401 ( .A(REG2_REG_22__SCAN_IN), .ZN(n2638) );
  OR2_X1 U3402 ( .A1(n3040), .A2(n2638), .ZN(n2641) );
  INV_X1 U3403 ( .A(REG1_REG_22__SCAN_IN), .ZN(n4659) );
  OR2_X1 U3404 ( .A1(n2141), .A2(n4659), .ZN(n2640) );
  OAI211_X1 U3405 ( .C1(n2860), .C2(n4896), .A(n2641), .B(n2640), .ZN(n2642)
         );
  INV_X1 U3406 ( .A(n2642), .ZN(n2643) );
  NAND2_X1 U3407 ( .A1(n2841), .A2(n3835), .ZN(n2645) );
  AND2_X1 U3408 ( .A1(n2646), .A2(n2645), .ZN(n4297) );
  NAND2_X1 U3409 ( .A1(n4297), .A2(n2891), .ZN(n2651) );
  INV_X1 U3410 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4531) );
  INV_X2 U3411 ( .A(n2672), .ZN(n2892) );
  NAND2_X1 U3412 ( .A1(n2892), .A2(REG2_REG_21__SCAN_IN), .ZN(n2648) );
  NAND2_X1 U3413 ( .A1(n3037), .A2(REG0_REG_21__SCAN_IN), .ZN(n2647) );
  OAI211_X1 U3414 ( .C1(n2142), .C2(n4531), .A(n2648), .B(n2647), .ZN(n2649)
         );
  INV_X1 U3415 ( .A(n2649), .ZN(n2650) );
  NAND2_X1 U3416 ( .A1(n3037), .A2(REG0_REG_0__SCAN_IN), .ZN(n2656) );
  INV_X1 U3417 ( .A(REG2_REG_0__SCAN_IN), .ZN(n4617) );
  OR2_X1 U3418 ( .A1(n2672), .A2(n4617), .ZN(n2653) );
  INV_X1 U3419 ( .A(REG3_REG_0__SCAN_IN), .ZN(n3722) );
  OR2_X1 U3420 ( .A1(n2681), .A2(n3722), .ZN(n2652) );
  AND2_X2 U3421 ( .A1(n2653), .A2(n2652), .ZN(n2655) );
  NAND2_X1 U3422 ( .A1(n2765), .A2(IR_REG_0__SCAN_IN), .ZN(n2657) );
  OR2_X1 U3423 ( .A1(n2672), .A2(n2573), .ZN(n2663) );
  NAND2_X1 U3424 ( .A1(n2659), .A2(REG1_REG_1__SCAN_IN), .ZN(n2662) );
  INV_X1 U3425 ( .A(REG3_REG_1__SCAN_IN), .ZN(n3204) );
  OR2_X1 U3426 ( .A1(n2681), .A2(n3204), .ZN(n2661) );
  INV_X1 U3427 ( .A(REG0_REG_1__SCAN_IN), .ZN(n4607) );
  NAND2_X1 U3428 ( .A1(n3164), .A2(n2664), .ZN(n3942) );
  NAND2_X1 U3429 ( .A1(n4477), .A2(n4602), .ZN(n2665) );
  NAND2_X1 U3430 ( .A1(n2659), .A2(REG1_REG_2__SCAN_IN), .ZN(n2671) );
  INV_X1 U3431 ( .A(REG0_REG_2__SCAN_IN), .ZN(n2666) );
  OR2_X1 U3432 ( .A1(n2680), .A2(n2666), .ZN(n2670) );
  INV_X1 U3433 ( .A(REG3_REG_2__SCAN_IN), .ZN(n3189) );
  OR2_X1 U3434 ( .A1(n2681), .A2(n3189), .ZN(n2669) );
  OR2_X1 U3435 ( .A1(n2672), .A2(n2667), .ZN(n2668) );
  AND4_X2 U3436 ( .A1(n2671), .A2(n2670), .A3(n2669), .A4(n2668), .ZN(n3379)
         );
  NAND2_X1 U3437 ( .A1(n3379), .A2(n3251), .ZN(n3243) );
  INV_X1 U3438 ( .A(n2672), .ZN(n2673) );
  NAND2_X1 U3439 ( .A1(n2673), .A2(REG2_REG_4__SCAN_IN), .ZN(n2677) );
  OAI21_X1 U3440 ( .B1(REG3_REG_3__SCAN_IN), .B2(REG3_REG_4__SCAN_IN), .A(
        n2696), .ZN(n3270) );
  OR2_X1 U3441 ( .A1(n2681), .A2(n3270), .ZN(n2676) );
  INV_X1 U3442 ( .A(REG0_REG_4__SCAN_IN), .ZN(n2674) );
  OR2_X1 U3443 ( .A1(n2680), .A2(n2674), .ZN(n2675) );
  NAND4_X2 U3444 ( .A1(n2677), .A2(n2678), .A3(n2676), .A4(n2675), .ZN(n4105)
         );
  AND4_X2 U3445 ( .A1(n2678), .A2(n2677), .A3(n2676), .A4(n2675), .ZN(n3210)
         );
  NAND2_X1 U3446 ( .A1(n2892), .A2(REG2_REG_3__SCAN_IN), .ZN(n2686) );
  OR2_X1 U3447 ( .A1(n2141), .A2(n3049), .ZN(n2685) );
  INV_X1 U3448 ( .A(REG0_REG_3__SCAN_IN), .ZN(n2679) );
  OR2_X1 U3449 ( .A1(n2680), .A2(n2679), .ZN(n2683) );
  OR2_X1 U3450 ( .A1(n2681), .A2(REG3_REG_3__SCAN_IN), .ZN(n2682) );
  INV_X1 U3451 ( .A(DATAI_3_), .ZN(n2687) );
  NAND2_X1 U3452 ( .A1(n3272), .A2(n3378), .ZN(n2688) );
  INV_X1 U3453 ( .A(n3378), .ZN(n3253) );
  AND2_X1 U3454 ( .A1(n3253), .A2(n2909), .ZN(n2689) );
  AOI22_X1 U3455 ( .A1(n3271), .A2(n2689), .B1(n3269), .B2(n4105), .ZN(n2692)
         );
  INV_X1 U3456 ( .A(n3251), .ZN(n3186) );
  NAND2_X1 U3457 ( .A1(n3379), .A2(n3186), .ZN(n3945) );
  NAND2_X1 U34580 ( .A1(n3251), .A2(n4475), .ZN(n3948) );
  NAND3_X1 U34590 ( .A1(n2690), .A2(n2908), .A3(n3243), .ZN(n2691) );
  NAND3_X1 U3460 ( .A1(n2693), .A2(n2692), .A3(n2691), .ZN(n3301) );
  NAND2_X1 U3461 ( .A1(n3036), .A2(REG1_REG_5__SCAN_IN), .ZN(n2702) );
  OR2_X1 U3462 ( .A1(n3040), .A2(n2694), .ZN(n2701) );
  INV_X1 U3463 ( .A(REG3_REG_5__SCAN_IN), .ZN(n2695) );
  NAND2_X1 U3464 ( .A1(n2696), .A2(n2695), .ZN(n2697) );
  NAND2_X1 U3465 ( .A1(n2717), .A2(n2697), .ZN(n3436) );
  OR2_X1 U3466 ( .A1(n2808), .A2(n3436), .ZN(n2700) );
  INV_X1 U34670 ( .A(REG0_REG_5__SCAN_IN), .ZN(n2698) );
  OR2_X1 U3468 ( .A1(n2860), .A2(n2698), .ZN(n2699) );
  INV_X1 U34690 ( .A(DATAI_5_), .ZN(n2703) );
  NAND2_X1 U3470 ( .A1(n3327), .A2(n3306), .ZN(n2704) );
  NAND2_X1 U34710 ( .A1(n3301), .A2(n2704), .ZN(n2706) );
  INV_X1 U3472 ( .A(n3306), .ZN(n3435) );
  NAND2_X1 U34730 ( .A1(n3435), .A2(n3403), .ZN(n2705) );
  NAND2_X1 U3474 ( .A1(n2706), .A2(n2705), .ZN(n3332) );
  NAND2_X1 U34750 ( .A1(n2892), .A2(REG2_REG_7__SCAN_IN), .ZN(n2714) );
  OR2_X1 U3476 ( .A1(n2141), .A2(n2707), .ZN(n2713) );
  INV_X1 U34770 ( .A(REG3_REG_7__SCAN_IN), .ZN(n4628) );
  NAND2_X1 U3478 ( .A1(n2177), .A2(n4628), .ZN(n2709) );
  NAND2_X1 U34790 ( .A1(n2739), .A2(n2709), .ZN(n3363) );
  OR2_X1 U3480 ( .A1(n2808), .A2(n3363), .ZN(n2712) );
  INV_X1 U34810 ( .A(REG0_REG_7__SCAN_IN), .ZN(n2710) );
  OR2_X1 U3482 ( .A1(n2860), .A2(n2710), .ZN(n2711) );
  NAND2_X1 U34830 ( .A1(n3354), .A2(n3345), .ZN(n2910) );
  INV_X1 U3484 ( .A(n3345), .ZN(n3358) );
  NAND2_X1 U34850 ( .A1(n2910), .A2(n3966), .ZN(n3338) );
  NAND2_X1 U3486 ( .A1(n2892), .A2(REG2_REG_6__SCAN_IN), .ZN(n2722) );
  INV_X1 U34870 ( .A(REG1_REG_6__SCAN_IN), .ZN(n2715) );
  INV_X1 U3488 ( .A(REG3_REG_6__SCAN_IN), .ZN(n2716) );
  NAND2_X1 U34890 ( .A1(n2717), .A2(n2716), .ZN(n2718) );
  NAND2_X1 U3490 ( .A1(n2177), .A2(n2718), .ZN(n3408) );
  OR2_X1 U34910 ( .A1(n2808), .A2(n3408), .ZN(n2721) );
  INV_X1 U3492 ( .A(REG0_REG_6__SCAN_IN), .ZN(n2719) );
  OR2_X1 U34930 ( .A1(n2860), .A2(n2719), .ZN(n2720) );
  NAND2_X1 U3494 ( .A1(n3332), .A2(n2725), .ZN(n2728) );
  AND2_X1 U34950 ( .A1(n3320), .A2(n3341), .ZN(n2726) );
  AOI22_X1 U3496 ( .A1(n3338), .A2(n2726), .B1(n3345), .B2(n4460), .ZN(n2727)
         );
  NAND2_X1 U34970 ( .A1(n2728), .A2(n2727), .ZN(n3425) );
  NAND2_X1 U3498 ( .A1(n3036), .A2(REG1_REG_8__SCAN_IN), .ZN(n2733) );
  INV_X1 U34990 ( .A(REG2_REG_8__SCAN_IN), .ZN(n4463) );
  OR2_X1 U3500 ( .A1(n3040), .A2(n4463), .ZN(n2732) );
  INV_X1 U35010 ( .A(REG3_REG_8__SCAN_IN), .ZN(n2738) );
  XNOR2_X1 U3502 ( .A(n2739), .B(n2738), .ZN(n4462) );
  OR2_X1 U35030 ( .A1(n2808), .A2(n4462), .ZN(n2731) );
  INV_X1 U3504 ( .A(REG0_REG_8__SCAN_IN), .ZN(n2729) );
  OR2_X1 U35050 ( .A1(n2860), .A2(n2729), .ZN(n2730) );
  INV_X1 U35060 ( .A(DATAI_8_), .ZN(n3010) );
  NAND2_X1 U35070 ( .A1(n3534), .A2(n3428), .ZN(n2734) );
  NAND2_X1 U35080 ( .A1(n4458), .A2(n4104), .ZN(n2735) );
  NAND2_X1 U35090 ( .A1(n2892), .A2(REG2_REG_9__SCAN_IN), .ZN(n2744) );
  OR2_X1 U35100 ( .A1(n2141), .A2(n4838), .ZN(n2743) );
  INV_X1 U35110 ( .A(REG3_REG_9__SCAN_IN), .ZN(n2737) );
  OAI21_X1 U35120 ( .B1(n2739), .B2(n2738), .A(n2737), .ZN(n2740) );
  NAND2_X1 U35130 ( .A1(n2740), .A2(n2749), .ZN(n3540) );
  OR2_X1 U35140 ( .A1(n2808), .A2(n3540), .ZN(n2742) );
  INV_X1 U35150 ( .A(REG0_REG_9__SCAN_IN), .ZN(n3493) );
  OR2_X1 U35160 ( .A1(n2860), .A2(n3493), .ZN(n2741) );
  NAND4_X1 U35170 ( .A1(n2744), .A2(n2743), .A3(n2742), .A4(n2741), .ZN(n4459)
         );
  AND2_X1 U35180 ( .A1(n3499), .A2(n4459), .ZN(n2746) );
  NAND2_X1 U35190 ( .A1(n3478), .A2(n3535), .ZN(n2745) );
  NAND2_X1 U35200 ( .A1(n3036), .A2(REG1_REG_10__SCAN_IN), .ZN(n2755) );
  INV_X1 U35210 ( .A(REG2_REG_10__SCAN_IN), .ZN(n2747) );
  OR2_X1 U35220 ( .A1(n3040), .A2(n2747), .ZN(n2754) );
  INV_X1 U35230 ( .A(REG3_REG_10__SCAN_IN), .ZN(n2748) );
  NAND2_X1 U35240 ( .A1(n2749), .A2(n2748), .ZN(n2750) );
  NAND2_X1 U35250 ( .A1(n2758), .A2(n2750), .ZN(n3567) );
  OR2_X1 U35260 ( .A1(n2808), .A2(n3567), .ZN(n2753) );
  INV_X1 U35270 ( .A(REG0_REG_10__SCAN_IN), .ZN(n2751) );
  OR2_X1 U35280 ( .A1(n2860), .A2(n2751), .ZN(n2752) );
  INV_X1 U35290 ( .A(DATAI_10_), .ZN(n3019) );
  NAND2_X1 U35300 ( .A1(n3480), .A2(n4102), .ZN(n2756) );
  INV_X1 U35310 ( .A(DATAI_11_), .ZN(n2757) );
  MUX2_X1 U35320 ( .A(n2757), .B(n4120), .S(n2765), .Z(n3576) );
  NAND2_X1 U35330 ( .A1(n2892), .A2(REG2_REG_11__SCAN_IN), .ZN(n2763) );
  OR2_X1 U35340 ( .A1(n2142), .A2(n3584), .ZN(n2762) );
  NAND2_X1 U35350 ( .A1(n2758), .A2(n4850), .ZN(n2759) );
  NAND2_X1 U35360 ( .A1(n2766), .A2(n2759), .ZN(n3586) );
  OR2_X1 U35370 ( .A1(n2808), .A2(n3586), .ZN(n2761) );
  INV_X1 U35380 ( .A(REG0_REG_11__SCAN_IN), .ZN(n3581) );
  OR2_X1 U35390 ( .A1(n2860), .A2(n3581), .ZN(n2760) );
  NAND4_X1 U35400 ( .A1(n2763), .A2(n2762), .A3(n2761), .A4(n2760), .ZN(n4585)
         );
  NAND2_X1 U35410 ( .A1(n3576), .A2(n4585), .ZN(n3543) );
  NAND2_X1 U35420 ( .A1(n2955), .A2(n3781), .ZN(n3541) );
  NAND2_X1 U35430 ( .A1(n3543), .A2(n3541), .ZN(n4024) );
  NAND2_X1 U35440 ( .A1(n3576), .A2(n3781), .ZN(n2764) );
  MUX2_X1 U35450 ( .A(DATAI_12_), .B(n4940), .S(n2765), .Z(n4583) );
  NAND2_X1 U35460 ( .A1(n2892), .A2(REG2_REG_12__SCAN_IN), .ZN(n2771) );
  INV_X1 U35470 ( .A(REG1_REG_12__SCAN_IN), .ZN(n4792) );
  OR2_X1 U35480 ( .A1(n2142), .A2(n4792), .ZN(n2770) );
  INV_X1 U35490 ( .A(REG3_REG_12__SCAN_IN), .ZN(n4714) );
  NAND2_X1 U35500 ( .A1(n2766), .A2(n4714), .ZN(n2767) );
  NAND2_X1 U35510 ( .A1(n2773), .A2(n2767), .ZN(n3548) );
  OR2_X1 U35520 ( .A1(n2808), .A2(n3548), .ZN(n2769) );
  INV_X1 U35530 ( .A(REG0_REG_12__SCAN_IN), .ZN(n4933) );
  OR2_X1 U35540 ( .A1(n2860), .A2(n4933), .ZN(n2768) );
  NAND4_X1 U35550 ( .A1(n2771), .A2(n2770), .A3(n2769), .A4(n2768), .ZN(n4101)
         );
  NAND2_X1 U35560 ( .A1(n4583), .A2(n4101), .ZN(n2772) );
  INV_X1 U35570 ( .A(n4443), .ZN(n2779) );
  MUX2_X1 U35580 ( .A(n4939), .B(DATAI_13_), .S(n2335), .Z(n4439) );
  NAND2_X1 U35590 ( .A1(n2773), .A2(n3607), .ZN(n2774) );
  NAND2_X1 U35600 ( .A1(n2780), .A2(n2774), .ZN(n4450) );
  NAND2_X1 U35610 ( .A1(n3037), .A2(REG0_REG_13__SCAN_IN), .ZN(n2775) );
  OAI21_X1 U35620 ( .B1(n4450), .B2(n2808), .A(n2775), .ZN(n2778) );
  NAND2_X1 U35630 ( .A1(n2892), .A2(REG2_REG_13__SCAN_IN), .ZN(n2776) );
  OAI21_X1 U35640 ( .B1(n2141), .B2(n4580), .A(n2776), .ZN(n2777) );
  INV_X1 U35650 ( .A(REG3_REG_14__SCAN_IN), .ZN(n4833) );
  NAND2_X1 U35660 ( .A1(n2780), .A2(n4833), .ZN(n2781) );
  NAND2_X1 U35670 ( .A1(n2792), .A2(n2781), .ZN(n3806) );
  OR2_X1 U35680 ( .A1(n3806), .A2(n2808), .ZN(n2784) );
  AOI22_X1 U35690 ( .A1(n2892), .A2(REG2_REG_14__SCAN_IN), .B1(n2659), .B2(
        REG1_REG_14__SCAN_IN), .ZN(n2783) );
  NAND2_X1 U35700 ( .A1(n3037), .A2(REG0_REG_14__SCAN_IN), .ZN(n2782) );
  MUX2_X1 U35710 ( .A(n4938), .B(DATAI_14_), .S(n2335), .Z(n3807) );
  NAND2_X1 U35720 ( .A1(n4437), .A2(n3807), .ZN(n3979) );
  INV_X1 U35730 ( .A(n4437), .ZN(n4562) );
  INV_X1 U35740 ( .A(n3807), .ZN(n4573) );
  NAND2_X1 U35750 ( .A1(n4562), .A2(n4573), .ZN(n3961) );
  NAND2_X1 U35760 ( .A1(n3979), .A2(n3961), .ZN(n4416) );
  NAND2_X1 U35770 ( .A1(n2794), .A2(n4734), .ZN(n2785) );
  AND2_X1 U35780 ( .A1(n2806), .A2(n2785), .ZN(n4406) );
  NAND2_X1 U35790 ( .A1(n4406), .A2(n2891), .ZN(n2790) );
  INV_X1 U35800 ( .A(REG1_REG_16__SCAN_IN), .ZN(n4656) );
  NAND2_X1 U35810 ( .A1(n2892), .A2(REG2_REG_16__SCAN_IN), .ZN(n2787) );
  NAND2_X1 U3582 ( .A1(n3037), .A2(REG0_REG_16__SCAN_IN), .ZN(n2786) );
  OAI211_X1 U3583 ( .C1(n2142), .C2(n4656), .A(n2787), .B(n2786), .ZN(n2788)
         );
  INV_X1 U3584 ( .A(n2788), .ZN(n2789) );
  NAND2_X1 U3585 ( .A1(n4381), .A2(n4405), .ZN(n2799) );
  INV_X1 U3586 ( .A(n2799), .ZN(n2798) );
  NAND2_X1 U3587 ( .A1(n4565), .A2(n4405), .ZN(n4058) );
  NAND2_X1 U3588 ( .A1(n4381), .A2(n3656), .ZN(n4055) );
  INV_X1 U3589 ( .A(n4399), .ZN(n4387) );
  INV_X1 U3590 ( .A(REG0_REG_15__SCAN_IN), .ZN(n4922) );
  NAND2_X1 U3591 ( .A1(n2792), .A2(n3922), .ZN(n2793) );
  NAND2_X1 U3592 ( .A1(n2794), .A2(n2793), .ZN(n3930) );
  OR2_X1 U3593 ( .A1(n3930), .A2(n2808), .ZN(n2796) );
  AOI22_X1 U3594 ( .A1(n2892), .A2(REG2_REG_15__SCAN_IN), .B1(n3036), .B2(
        REG1_REG_15__SCAN_IN), .ZN(n2795) );
  INV_X1 U3595 ( .A(n4570), .ZN(n2921) );
  INV_X1 U3596 ( .A(n4561), .ZN(n3924) );
  NAND2_X1 U3597 ( .A1(n2921), .A2(n3924), .ZN(n4397) );
  AND2_X1 U3598 ( .A1(n4387), .A2(n4397), .ZN(n4396) );
  INV_X1 U3599 ( .A(n2802), .ZN(n2801) );
  NAND2_X1 U3600 ( .A1(n4570), .A2(n4561), .ZN(n4394) );
  AND2_X1 U3601 ( .A1(n4394), .A2(n2799), .ZN(n2800) );
  AND2_X1 U3602 ( .A1(n4416), .A2(n4370), .ZN(n2804) );
  INV_X1 U3603 ( .A(n4370), .ZN(n2803) );
  NAND2_X1 U3604 ( .A1(n4437), .A2(n4573), .ZN(n3613) );
  AND2_X1 U3605 ( .A1(n3613), .A2(n2802), .ZN(n4369) );
  INV_X1 U3606 ( .A(REG3_REG_17__SCAN_IN), .ZN(n2805) );
  NAND2_X1 U3607 ( .A1(n2806), .A2(n2805), .ZN(n2807) );
  NAND2_X1 U3608 ( .A1(n2817), .A2(n2807), .ZN(n4377) );
  INV_X1 U3609 ( .A(REG2_REG_17__SCAN_IN), .ZN(n4378) );
  NAND2_X1 U3610 ( .A1(n3037), .A2(REG0_REG_17__SCAN_IN), .ZN(n2810) );
  OR2_X1 U3611 ( .A1(n2141), .A2(n2525), .ZN(n2809) );
  OAI211_X1 U3612 ( .C1(n3040), .C2(n4378), .A(n2810), .B(n2809), .ZN(n2811)
         );
  INV_X1 U3613 ( .A(n2811), .ZN(n2812) );
  INV_X1 U3614 ( .A(DATAI_17_), .ZN(n2814) );
  NAND2_X1 U3615 ( .A1(n4391), .A2(n4546), .ZN(n2815) );
  INV_X1 U3616 ( .A(n4546), .ZN(n4380) );
  AOI22_X1 U3617 ( .A1(n2816), .A2(n2815), .B1(n4380), .B2(n4350), .ZN(n4357)
         );
  NAND2_X1 U3618 ( .A1(n2817), .A2(n2296), .ZN(n2818) );
  NAND2_X1 U3619 ( .A1(n2828), .A2(n2818), .ZN(n4363) );
  NAND2_X1 U3620 ( .A1(n2892), .A2(REG2_REG_18__SCAN_IN), .ZN(n2820) );
  NAND2_X1 U3621 ( .A1(n3037), .A2(REG0_REG_18__SCAN_IN), .ZN(n2819) );
  OAI211_X1 U3622 ( .C1(n2142), .C2(n2821), .A(n2820), .B(n2819), .ZN(n2822)
         );
  INV_X1 U3623 ( .A(n2822), .ZN(n2823) );
  MUX2_X1 U3624 ( .A(n2825), .B(DATAI_18_), .S(n2335), .Z(n4349) );
  NAND2_X1 U3625 ( .A1(n4334), .A2(n4349), .ZN(n4329) );
  INV_X1 U3626 ( .A(n4349), .ZN(n4360) );
  NAND2_X1 U3627 ( .A1(n4549), .A2(n4360), .ZN(n4330) );
  NAND2_X1 U3628 ( .A1(n4329), .A2(n4330), .ZN(n4356) );
  NAND2_X1 U3629 ( .A1(n4357), .A2(n4356), .ZN(n4355) );
  NAND2_X1 U3630 ( .A1(n2828), .A2(n2827), .ZN(n2829) );
  AND2_X1 U3631 ( .A1(n2839), .A2(n2829), .ZN(n4343) );
  NAND2_X1 U3632 ( .A1(n4343), .A2(n2891), .ZN(n2835) );
  INV_X1 U3633 ( .A(REG2_REG_19__SCAN_IN), .ZN(n2832) );
  NAND2_X1 U3634 ( .A1(n3037), .A2(REG0_REG_19__SCAN_IN), .ZN(n2831) );
  OR2_X1 U3635 ( .A1(n2142), .A2(n2535), .ZN(n2830) );
  OAI211_X1 U3636 ( .C1(n3040), .C2(n2832), .A(n2831), .B(n2830), .ZN(n2833)
         );
  INV_X1 U3637 ( .A(n2833), .ZN(n2834) );
  INV_X1 U3638 ( .A(DATAI_19_), .ZN(n2836) );
  NAND2_X1 U3639 ( .A1(n2839), .A2(n2297), .ZN(n2840) );
  NAND2_X1 U3640 ( .A1(n2841), .A2(n2840), .ZN(n3875) );
  OR2_X1 U3641 ( .A1(n3875), .A2(n2808), .ZN(n2846) );
  INV_X1 U3642 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4904) );
  NAND2_X1 U3643 ( .A1(n2892), .A2(REG2_REG_20__SCAN_IN), .ZN(n2843) );
  NAND2_X1 U3644 ( .A1(n3036), .A2(REG1_REG_20__SCAN_IN), .ZN(n2842) );
  OAI211_X1 U3645 ( .C1(n4904), .C2(n2860), .A(n2843), .B(n2842), .ZN(n2844)
         );
  INV_X1 U3646 ( .A(n2844), .ZN(n2845) );
  NAND2_X1 U3647 ( .A1(n4525), .A2(n4310), .ZN(n4036) );
  NOR2_X1 U3648 ( .A1(n4525), .A2(n4310), .ZN(n4037) );
  NAND2_X1 U3649 ( .A1(n4527), .A2(n4268), .ZN(n4251) );
  INV_X1 U3650 ( .A(n4527), .ZN(n3199) );
  NAND2_X1 U3651 ( .A1(n3199), .A2(n4273), .ZN(n2932) );
  NAND2_X1 U3652 ( .A1(n4251), .A2(n2932), .ZN(n4278) );
  NAND2_X1 U3653 ( .A1(n2847), .A2(n4668), .ZN(n2848) );
  AND2_X1 U3654 ( .A1(n2855), .A2(n2848), .ZN(n4259) );
  NAND2_X1 U3655 ( .A1(n4259), .A2(n2891), .ZN(n2853) );
  INV_X1 U3656 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4517) );
  NAND2_X1 U3657 ( .A1(n2892), .A2(REG2_REG_23__SCAN_IN), .ZN(n2850) );
  NAND2_X1 U3658 ( .A1(n3037), .A2(REG0_REG_23__SCAN_IN), .ZN(n2849) );
  OAI211_X1 U3659 ( .C1(n2142), .C2(n4517), .A(n2850), .B(n2849), .ZN(n2851)
         );
  INV_X1 U3660 ( .A(n2851), .ZN(n2852) );
  NAND2_X1 U3661 ( .A1(n4272), .A2(n4258), .ZN(n2854) );
  INV_X1 U3662 ( .A(REG3_REG_24__SCAN_IN), .ZN(n4822) );
  NAND2_X1 U3663 ( .A1(n2855), .A2(n4822), .ZN(n2856) );
  NAND2_X1 U3664 ( .A1(n4243), .A2(n2891), .ZN(n2863) );
  INV_X1 U3665 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4888) );
  INV_X1 U3666 ( .A(REG2_REG_24__SCAN_IN), .ZN(n2857) );
  OR2_X1 U3667 ( .A1(n3040), .A2(n2857), .ZN(n2859) );
  INV_X1 U3668 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4666) );
  OR2_X1 U3669 ( .A1(n2141), .A2(n4666), .ZN(n2858) );
  OAI211_X1 U3670 ( .C1(n2860), .C2(n4888), .A(n2859), .B(n2858), .ZN(n2861)
         );
  INV_X1 U3671 ( .A(n2861), .ZN(n2862) );
  NAND2_X1 U3672 ( .A1(n4504), .A2(n4240), .ZN(n2864) );
  INV_X1 U3673 ( .A(REG3_REG_25__SCAN_IN), .ZN(n2865) );
  NAND2_X1 U3674 ( .A1(n2866), .A2(n2865), .ZN(n2867) );
  NAND2_X1 U3675 ( .A1(n4220), .A2(n2891), .ZN(n2872) );
  INV_X1 U3676 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4884) );
  NAND2_X1 U3677 ( .A1(n2892), .A2(REG2_REG_25__SCAN_IN), .ZN(n2869) );
  INV_X1 U3678 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4510) );
  OR2_X1 U3679 ( .A1(n2141), .A2(n4510), .ZN(n2868) );
  OAI211_X1 U3680 ( .C1(n4884), .C2(n2860), .A(n2869), .B(n2868), .ZN(n2870)
         );
  INV_X1 U3681 ( .A(n2870), .ZN(n2871) );
  NAND2_X1 U3682 ( .A1(n2335), .A2(DATAI_25_), .ZN(n4222) );
  INV_X1 U3683 ( .A(REG3_REG_26__SCAN_IN), .ZN(n4824) );
  NAND2_X1 U3684 ( .A1(n2874), .A2(n4824), .ZN(n2875) );
  NAND2_X1 U3685 ( .A1(n2889), .A2(n2875), .ZN(n4209) );
  NAND2_X1 U3686 ( .A1(n3037), .A2(REG0_REG_26__SCAN_IN), .ZN(n2877) );
  NAND2_X1 U3687 ( .A1(n3036), .A2(REG1_REG_26__SCAN_IN), .ZN(n2876) );
  OAI211_X1 U3688 ( .C1(n3040), .C2(n4809), .A(n2877), .B(n2876), .ZN(n2878)
         );
  INV_X1 U3689 ( .A(n2878), .ZN(n2879) );
  INV_X1 U3690 ( .A(n4493), .ZN(n4506) );
  XNOR2_X1 U3691 ( .A(n2889), .B(REG3_REG_27__SCAN_IN), .ZN(n4187) );
  NAND2_X1 U3692 ( .A1(n4187), .A2(n2891), .ZN(n2885) );
  INV_X1 U3693 ( .A(REG2_REG_27__SCAN_IN), .ZN(n4184) );
  NAND2_X1 U3694 ( .A1(n3037), .A2(REG0_REG_27__SCAN_IN), .ZN(n2882) );
  NAND2_X1 U3695 ( .A1(n3036), .A2(REG1_REG_27__SCAN_IN), .ZN(n2881) );
  OAI211_X1 U3696 ( .C1(n3040), .C2(n4184), .A(n2882), .B(n2881), .ZN(n2883)
         );
  INV_X1 U3697 ( .A(n2883), .ZN(n2884) );
  NAND2_X1 U3698 ( .A1(n3997), .A2(n4185), .ZN(n2886) );
  INV_X1 U3699 ( .A(REG3_REG_27__SCAN_IN), .ZN(n3744) );
  INV_X1 U3700 ( .A(REG3_REG_28__SCAN_IN), .ZN(n2887) );
  OAI21_X1 U3701 ( .B1(n2889), .B2(n3744), .A(n2887), .ZN(n2890) );
  NAND2_X1 U3702 ( .A1(REG3_REG_27__SCAN_IN), .A2(REG3_REG_28__SCAN_IN), .ZN(
        n2888) );
  NAND2_X1 U3703 ( .A1(n3762), .A2(n2891), .ZN(n2898) );
  INV_X1 U3704 ( .A(REG0_REG_28__SCAN_IN), .ZN(n2895) );
  NAND2_X1 U3705 ( .A1(n2892), .A2(REG2_REG_28__SCAN_IN), .ZN(n2894) );
  NAND2_X1 U3706 ( .A1(n3036), .A2(REG1_REG_28__SCAN_IN), .ZN(n2893) );
  OAI211_X1 U3707 ( .C1(n2895), .C2(n2860), .A(n2894), .B(n2893), .ZN(n2896)
         );
  INV_X1 U3708 ( .A(n2896), .ZN(n2897) );
  NAND2_X1 U3709 ( .A1(n4495), .A2(n3761), .ZN(n3999) );
  INV_X1 U3710 ( .A(n3761), .ZN(n3786) );
  NAND2_X1 U3711 ( .A1(n4098), .A2(n3786), .ZN(n3934) );
  XNOR2_X1 U3712 ( .A(n3787), .B(n4052), .ZN(n3630) );
  XNOR2_X1 U3713 ( .A(n3162), .B(n4092), .ZN(n2901) );
  NAND2_X1 U3714 ( .A1(n2901), .A2(n3346), .ZN(n4418) );
  NAND3_X1 U3715 ( .A1(n2957), .A2(n3071), .A3(n4087), .ZN(n3571) );
  INV_X1 U3716 ( .A(n4596), .ZN(n4543) );
  INV_X1 U3717 ( .A(n2941), .ZN(n3076) );
  INV_X1 U3718 ( .A(REG2_REG_29__SCAN_IN), .ZN(n4178) );
  NAND2_X1 U3719 ( .A1(n3037), .A2(REG0_REG_29__SCAN_IN), .ZN(n2903) );
  NAND2_X1 U3720 ( .A1(n3036), .A2(REG1_REG_29__SCAN_IN), .ZN(n2902) );
  OAI211_X1 U3721 ( .C1(n3040), .C2(n4178), .A(n2903), .B(n2902), .ZN(n2904)
         );
  INV_X1 U3722 ( .A(n2904), .ZN(n2905) );
  INV_X1 U3723 ( .A(n4097), .ZN(n3765) );
  NAND2_X1 U3724 ( .A1(n2941), .A2(n4947), .ZN(n4564) );
  INV_X1 U3725 ( .A(n4082), .ZN(n3940) );
  AND2_X1 U3726 ( .A1(n4600), .A2(n2958), .ZN(n4582) );
  OAI22_X1 U3727 ( .A1(n3765), .A2(n4564), .B1(n4572), .B2(n3786), .ZN(n2936)
         );
  NAND2_X1 U3728 ( .A1(n2972), .A2(n2908), .ZN(n2971) );
  NAND2_X1 U3729 ( .A1(n2971), .A2(n3945), .ZN(n3247) );
  NAND2_X1 U3730 ( .A1(n3272), .A2(n3253), .ZN(n3950) );
  NAND2_X1 U3731 ( .A1(n3378), .A2(n2909), .ZN(n3947) );
  NAND2_X1 U3732 ( .A1(n3327), .A2(n3435), .ZN(n3967) );
  INV_X1 U3733 ( .A(n3320), .ZN(n3411) );
  NAND2_X1 U3734 ( .A1(n3411), .A2(n3341), .ZN(n3968) );
  NAND2_X1 U3735 ( .A1(n2723), .A2(n3320), .ZN(n3955) );
  INV_X1 U3736 ( .A(n2910), .ZN(n2911) );
  NAND2_X1 U3737 ( .A1(n3534), .A2(n4458), .ZN(n3958) );
  NAND2_X1 U3738 ( .A1(n3428), .A2(n4104), .ZN(n3969) );
  AND2_X1 U3739 ( .A1(n3535), .A2(n4459), .ZN(n3447) );
  INV_X1 U3740 ( .A(n3447), .ZN(n2912) );
  NAND2_X1 U3741 ( .A1(n3478), .A2(n3499), .ZN(n3959) );
  NAND2_X1 U3742 ( .A1(n3562), .A2(n4102), .ZN(n3974) );
  NAND2_X1 U3743 ( .A1(n3480), .A2(n3509), .ZN(n3971) );
  NAND2_X1 U3744 ( .A1(n2913), .A2(n3971), .ZN(n3574) );
  NAND2_X1 U3745 ( .A1(n3596), .A2(n4101), .ZN(n4431) );
  NAND2_X1 U3746 ( .A1(n4445), .A2(n4586), .ZN(n2914) );
  NAND2_X1 U3747 ( .A1(n4431), .A2(n2914), .ZN(n2916) );
  INV_X1 U3748 ( .A(n3543), .ZN(n2915) );
  NOR2_X1 U3749 ( .A1(n2916), .A2(n2915), .ZN(n3975) );
  NAND2_X1 U3750 ( .A1(n3574), .A2(n3975), .ZN(n2920) );
  INV_X1 U3751 ( .A(n2916), .ZN(n2919) );
  NAND2_X1 U3752 ( .A1(n4583), .A2(n4436), .ZN(n4433) );
  NAND2_X1 U3753 ( .A1(n4433), .A2(n3541), .ZN(n2918) );
  NOR2_X1 U3754 ( .A1(n4445), .A2(n4586), .ZN(n2917) );
  AOI21_X1 U3755 ( .B1(n2919), .B2(n2918), .A(n2917), .ZN(n3983) );
  INV_X1 U3756 ( .A(n4416), .ZN(n4021) );
  NAND2_X1 U3757 ( .A1(n4413), .A2(n4021), .ZN(n4414) );
  NAND2_X1 U3758 ( .A1(n2921), .A2(n4561), .ZN(n3980) );
  NAND2_X1 U3759 ( .A1(n4570), .A2(n3924), .ZN(n3962) );
  NAND2_X1 U3760 ( .A1(n3980), .A2(n3962), .ZN(n4018) );
  INV_X1 U3761 ( .A(n3979), .ZN(n2922) );
  NOR2_X1 U3762 ( .A1(n4018), .A2(n2922), .ZN(n2923) );
  NAND2_X1 U3763 ( .A1(n4414), .A2(n2923), .ZN(n2924) );
  NAND2_X1 U3764 ( .A1(n2924), .A2(n3962), .ZN(n4388) );
  AND2_X1 U3765 ( .A1(n4350), .A2(n4546), .ZN(n3988) );
  NAND2_X1 U3766 ( .A1(n4311), .A2(n4341), .ZN(n2926) );
  NAND2_X1 U3767 ( .A1(n2926), .A2(n4330), .ZN(n3987) );
  INV_X1 U3768 ( .A(n4310), .ZN(n4320) );
  NAND2_X1 U3769 ( .A1(n4525), .A2(n4320), .ZN(n4056) );
  NAND2_X1 U3770 ( .A1(n4313), .A2(n4524), .ZN(n4250) );
  NAND2_X1 U3771 ( .A1(n4251), .A2(n4250), .ZN(n3991) );
  NAND2_X1 U3772 ( .A1(n4391), .A2(n4380), .ZN(n4327) );
  AND2_X1 U3773 ( .A1(n4329), .A2(n4327), .ZN(n2927) );
  OR2_X1 U3774 ( .A1(n2927), .A2(n3987), .ZN(n2929) );
  NAND2_X1 U3775 ( .A1(n4352), .A2(n4040), .ZN(n2928) );
  AND2_X1 U3776 ( .A1(n2929), .A2(n2928), .ZN(n4307) );
  INV_X1 U3777 ( .A(n4525), .ZN(n4294) );
  NAND2_X1 U3778 ( .A1(n4294), .A2(n4310), .ZN(n2930) );
  NAND2_X1 U3779 ( .A1(n4307), .A2(n2930), .ZN(n2931) );
  AND2_X1 U3780 ( .A1(n2931), .A2(n4056), .ZN(n3939) );
  NOR2_X1 U3781 ( .A1(n3991), .A2(n3939), .ZN(n4060) );
  AND2_X1 U3782 ( .A1(n4269), .A2(n4300), .ZN(n4012) );
  AND2_X1 U3783 ( .A1(n4251), .A2(n4012), .ZN(n4061) );
  NAND2_X1 U3784 ( .A1(n4099), .A2(n4258), .ZN(n4011) );
  NAND2_X1 U3785 ( .A1(n4011), .A2(n2932), .ZN(n3936) );
  AOI211_X2 U3786 ( .C1(n4288), .C2(n4060), .A(n4061), .B(n3936), .ZN(n4232)
         );
  OR2_X1 U3787 ( .A1(n4504), .A2(n4235), .ZN(n4009) );
  OR2_X1 U3788 ( .A1(n4099), .A2(n4258), .ZN(n4230) );
  NAND2_X1 U3789 ( .A1(n4009), .A2(n4230), .ZN(n4065) );
  NAND2_X1 U3790 ( .A1(n4504), .A2(n4235), .ZN(n4010) );
  OAI21_X1 U3791 ( .B1(n4232), .B2(n4065), .A(n4010), .ZN(n4215) );
  AND2_X1 U3792 ( .A1(n4237), .A2(n4222), .ZN(n3937) );
  OAI21_X1 U3793 ( .B1(n4493), .B2(n4208), .A(n4196), .ZN(n4070) );
  NAND2_X1 U3794 ( .A1(n4493), .A2(n4208), .ZN(n3935) );
  OR2_X1 U3795 ( .A1(n4203), .A2(n4185), .ZN(n3998) );
  NAND2_X1 U3796 ( .A1(n2958), .A2(n4082), .ZN(n2934) );
  NAND2_X1 U3797 ( .A1(n4092), .A2(n4087), .ZN(n2933) );
  NAND2_X1 U3798 ( .A1(n2937), .A2(n3008), .ZN(n2938) );
  MUX2_X1 U3799 ( .A(n3008), .B(n2938), .S(B_REG_SCAN_IN), .Z(n2939) );
  INV_X1 U3800 ( .A(D_REG_0__SCAN_IN), .ZN(n3027) );
  INV_X1 U3801 ( .A(n3068), .ZN(n2981) );
  NAND2_X1 U3802 ( .A1(n2937), .A2(n2940), .ZN(n3024) );
  OAI21_X1 U3803 ( .B1(n2977), .B2(D_REG_1__SCAN_IN), .A(n3024), .ZN(n3066) );
  OR2_X1 U3804 ( .A1(n3571), .A2(n4082), .ZN(n2982) );
  NAND2_X1 U3805 ( .A1(n2957), .A2(n3346), .ZN(n3074) );
  NAND2_X1 U3806 ( .A1(n2941), .A2(n3074), .ZN(n3078) );
  NAND2_X1 U3807 ( .A1(n2982), .A2(n3078), .ZN(n2942) );
  NOR2_X1 U3808 ( .A1(n3086), .A2(n2942), .ZN(n2953) );
  NOR3_X1 U3809 ( .A1(D_REG_11__SCAN_IN), .A2(D_REG_30__SCAN_IN), .A3(
        D_REG_28__SCAN_IN), .ZN(n2944) );
  NOR4_X1 U3810 ( .A1(D_REG_2__SCAN_IN), .A2(D_REG_15__SCAN_IN), .A3(
        D_REG_27__SCAN_IN), .A4(D_REG_5__SCAN_IN), .ZN(n2943) );
  INV_X1 U3811 ( .A(D_REG_3__SCAN_IN), .ZN(n5015) );
  INV_X1 U3812 ( .A(D_REG_19__SCAN_IN), .ZN(n5006) );
  NAND4_X1 U3813 ( .A1(n2944), .A2(n2943), .A3(n5015), .A4(n5006), .ZN(n4632)
         );
  OR4_X1 U3814 ( .A1(D_REG_26__SCAN_IN), .A2(D_REG_31__SCAN_IN), .A3(
        D_REG_9__SCAN_IN), .A4(D_REG_13__SCAN_IN), .ZN(n2950) );
  NOR4_X1 U3815 ( .A1(D_REG_21__SCAN_IN), .A2(D_REG_7__SCAN_IN), .A3(
        D_REG_6__SCAN_IN), .A4(D_REG_8__SCAN_IN), .ZN(n2948) );
  NOR4_X1 U3816 ( .A1(D_REG_17__SCAN_IN), .A2(D_REG_29__SCAN_IN), .A3(
        D_REG_14__SCAN_IN), .A4(D_REG_4__SCAN_IN), .ZN(n2947) );
  NOR4_X1 U3817 ( .A1(D_REG_23__SCAN_IN), .A2(D_REG_20__SCAN_IN), .A3(
        D_REG_22__SCAN_IN), .A4(D_REG_24__SCAN_IN), .ZN(n2946) );
  NOR4_X1 U3818 ( .A1(D_REG_10__SCAN_IN), .A2(D_REG_18__SCAN_IN), .A3(
        D_REG_12__SCAN_IN), .A4(D_REG_16__SCAN_IN), .ZN(n2945) );
  NAND4_X1 U3819 ( .A1(n2948), .A2(n2947), .A3(n2946), .A4(n2945), .ZN(n2949)
         );
  OR4_X1 U3820 ( .A1(D_REG_25__SCAN_IN), .A2(n4632), .A3(n2950), .A4(n2949), 
        .ZN(n2951) );
  NAND2_X1 U3821 ( .A1(n2952), .A2(n2951), .ZN(n3067) );
  AND2_X1 U3822 ( .A1(n3251), .A2(n3378), .ZN(n2954) );
  AND2_X2 U3823 ( .A1(n4318), .A2(n4300), .ZN(n4291) );
  AND2_X2 U3824 ( .A1(n4291), .A2(n4273), .ZN(n4275) );
  NAND2_X1 U3825 ( .A1(n4183), .A2(n3761), .ZN(n2956) );
  NAND2_X1 U3826 ( .A1(n3795), .A2(n2956), .ZN(n3626) );
  OR2_X1 U3827 ( .A1(n3626), .A2(n4936), .ZN(n2961) );
  NAND2_X1 U3828 ( .A1(n5039), .A2(REG0_REG_28__SCAN_IN), .ZN(n2960) );
  INV_X1 U3829 ( .A(REG1_REG_28__SCAN_IN), .ZN(n2965) );
  INV_X1 U3830 ( .A(n3212), .ZN(n3092) );
  OR2_X1 U3831 ( .A1(n2968), .A2(n2908), .ZN(n3244) );
  NAND2_X1 U3832 ( .A1(n2968), .A2(n2908), .ZN(n2969) );
  AND2_X1 U3833 ( .A1(n3244), .A2(n2969), .ZN(n3143) );
  INV_X1 U3834 ( .A(n3143), .ZN(n2970) );
  INV_X1 U3835 ( .A(n4418), .ZN(n3578) );
  NAND2_X1 U3836 ( .A1(n2970), .A2(n3578), .ZN(n2975) );
  OAI21_X1 U3837 ( .B1(n2908), .B2(n2972), .A(n2971), .ZN(n2973) );
  NAND2_X1 U3838 ( .A1(n2973), .A2(n4595), .ZN(n2974) );
  NAND2_X1 U3839 ( .A1(n2975), .A2(n2974), .ZN(n3144) );
  AND3_X1 U3840 ( .A1(n3067), .A2(n3024), .A3(n3078), .ZN(n2980) );
  INV_X1 U3841 ( .A(D_REG_1__SCAN_IN), .ZN(n2978) );
  INV_X1 U3842 ( .A(n3086), .ZN(n2976) );
  OAI21_X1 U3843 ( .B1(n3086), .B2(n2978), .A(n5012), .ZN(n2979) );
  NAND3_X1 U3844 ( .A1(n2981), .A2(n2980), .A3(n2979), .ZN(n2983) );
  NAND2_X2 U3845 ( .A1(n2983), .A2(n4461), .ZN(n4484) );
  MUX2_X1 U3846 ( .A(REG2_REG_2__SCAN_IN), .B(n3144), .S(n4484), .Z(n2989) );
  AND2_X1 U3847 ( .A1(n4484), .A2(n4584), .ZN(n4474) );
  INV_X1 U3848 ( .A(n4474), .ZN(n4293) );
  NAND2_X1 U3849 ( .A1(n4484), .A2(n4601), .ZN(n4295) );
  OAI22_X1 U3850 ( .A1(n4293), .A2(n2984), .B1(n3272), .B2(n4295), .ZN(n2988)
         );
  OR2_X1 U3851 ( .A1(n3162), .A2(n3346), .ZN(n3336) );
  INV_X1 U3852 ( .A(n3336), .ZN(n2985) );
  AND2_X1 U3853 ( .A1(n4484), .A2(n2985), .ZN(n4483) );
  INV_X1 U3854 ( .A(n4483), .ZN(n4429) );
  OAI22_X1 U3855 ( .A1(n4429), .A2(n3143), .B1(n3189), .B2(n4461), .ZN(n2987)
         );
  AND2_X1 U3856 ( .A1(n4484), .A2(n4582), .ZN(n4478) );
  INV_X1 U3857 ( .A(n4478), .ZN(n4424) );
  XNOR2_X1 U3858 ( .A(n3252), .B(n3251), .ZN(n3146) );
  OAI22_X1 U3859 ( .A1(n4424), .A2(n3251), .B1(n3146), .B2(n4449), .ZN(n2986)
         );
  OR4_X1 U3860 ( .A1(n2989), .A2(n2988), .A3(n2987), .A4(n2986), .ZN(U3288) );
  MUX2_X1 U3861 ( .A(n2687), .B(n3054), .S(STATE_REG_SCAN_IN), .Z(n2990) );
  INV_X1 U3862 ( .A(n2990), .ZN(U3349) );
  NAND3_X1 U3863 ( .A1(n2992), .A2(IR_REG_31__SCAN_IN), .A3(STATE_REG_SCAN_IN), 
        .ZN(n2994) );
  INV_X1 U3864 ( .A(DATAI_31_), .ZN(n2993) );
  OAI22_X1 U3865 ( .A1(n2991), .A2(n2994), .B1(STATE_REG_SCAN_IN), .B2(n2993), 
        .ZN(U3321) );
  MUX2_X1 U3866 ( .A(n2703), .B(n3063), .S(STATE_REG_SCAN_IN), .Z(n2995) );
  INV_X1 U3867 ( .A(n2995), .ZN(U3347) );
  INV_X1 U3868 ( .A(DATAI_26_), .ZN(n2998) );
  NAND2_X1 U3869 ( .A1(n2996), .A2(STATE_REG_SCAN_IN), .ZN(n2997) );
  OAI21_X1 U3870 ( .B1(STATE_REG_SCAN_IN), .B2(n2998), .A(n2997), .ZN(U3326)
         );
  INV_X1 U3871 ( .A(DATAI_22_), .ZN(n3000) );
  NAND2_X1 U3872 ( .A1(n4092), .A2(STATE_REG_SCAN_IN), .ZN(n2999) );
  OAI21_X1 U3873 ( .B1(STATE_REG_SCAN_IN), .B2(n3000), .A(n2999), .ZN(U3330)
         );
  INV_X1 U3874 ( .A(DATAI_29_), .ZN(n4723) );
  NAND2_X1 U3875 ( .A1(n3001), .A2(STATE_REG_SCAN_IN), .ZN(n3002) );
  OAI21_X1 U3876 ( .B1(STATE_REG_SCAN_IN), .B2(n4723), .A(n3002), .ZN(U3323)
         );
  INV_X1 U3877 ( .A(DATAI_21_), .ZN(n4813) );
  NAND2_X1 U3878 ( .A1(n4082), .A2(STATE_REG_SCAN_IN), .ZN(n3003) );
  OAI21_X1 U3879 ( .B1(STATE_REG_SCAN_IN), .B2(n4813), .A(n3003), .ZN(U3331)
         );
  INV_X1 U3880 ( .A(DATAI_30_), .ZN(n3006) );
  NAND2_X1 U3881 ( .A1(n3004), .A2(STATE_REG_SCAN_IN), .ZN(n3005) );
  OAI21_X1 U3882 ( .B1(STATE_REG_SCAN_IN), .B2(n3006), .A(n3005), .ZN(U3322)
         );
  INV_X1 U3883 ( .A(DATAI_24_), .ZN(n3007) );
  MUX2_X1 U3884 ( .A(n3008), .B(n3007), .S(U3149), .Z(n3009) );
  INV_X1 U3885 ( .A(n3009), .ZN(U3328) );
  MUX2_X1 U3886 ( .A(n3010), .B(n3263), .S(STATE_REG_SCAN_IN), .Z(n3011) );
  INV_X1 U3887 ( .A(n3011), .ZN(U3344) );
  INV_X1 U3888 ( .A(DATAI_20_), .ZN(n3013) );
  NAND2_X1 U3889 ( .A1(n2958), .A2(STATE_REG_SCAN_IN), .ZN(n3012) );
  OAI21_X1 U3890 ( .B1(STATE_REG_SCAN_IN), .B2(n3013), .A(n3012), .ZN(U3332)
         );
  MUX2_X1 U3891 ( .A(n3346), .B(n2836), .S(U3149), .Z(n3014) );
  INV_X1 U3892 ( .A(n3014), .ZN(U3333) );
  INV_X1 U3893 ( .A(DATAI_25_), .ZN(n3017) );
  NAND2_X1 U3894 ( .A1(n3015), .A2(STATE_REG_SCAN_IN), .ZN(n3016) );
  OAI21_X1 U3895 ( .B1(STATE_REG_SCAN_IN), .B2(n3017), .A(n3016), .ZN(U3327)
         );
  MUX2_X1 U3896 ( .A(n3019), .B(n3018), .S(STATE_REG_SCAN_IN), .Z(n3020) );
  INV_X1 U3897 ( .A(n3020), .ZN(U3342) );
  INV_X1 U3898 ( .A(DATAI_9_), .ZN(n3021) );
  MUX2_X1 U3899 ( .A(n3375), .B(n3021), .S(U3149), .Z(n3022) );
  INV_X1 U3900 ( .A(n3022), .ZN(U3343) );
  MUX2_X1 U3901 ( .A(n2757), .B(n4120), .S(STATE_REG_SCAN_IN), .Z(n3023) );
  INV_X1 U3902 ( .A(n3023), .ZN(U3341) );
  INV_X1 U3903 ( .A(n3024), .ZN(n3025) );
  AOI22_X1 U3904 ( .A1(n5012), .A2(n2978), .B1(n3025), .B2(n5018), .ZN(U3459)
         );
  AOI22_X1 U3905 ( .A1(n5012), .A2(n3027), .B1(n5018), .B2(n3026), .ZN(U3458)
         );
  NOR2_X1 U3906 ( .A1(n4994), .A2(n4103), .ZN(U3148) );
  INV_X1 U3907 ( .A(DATAO_REG_31__SCAN_IN), .ZN(n4748) );
  INV_X1 U3908 ( .A(REG0_REG_31__SCAN_IN), .ZN(n3636) );
  INV_X1 U3909 ( .A(REG2_REG_31__SCAN_IN), .ZN(n3028) );
  OR2_X1 U3910 ( .A1(n3040), .A2(n3028), .ZN(n3030) );
  NAND2_X1 U3911 ( .A1(n3036), .A2(REG1_REG_31__SCAN_IN), .ZN(n3029) );
  OAI211_X1 U3912 ( .C1(n2860), .C2(n3636), .A(n3030), .B(n3029), .ZN(n4004)
         );
  NAND2_X1 U3913 ( .A1(U4043), .A2(n4004), .ZN(n3031) );
  OAI21_X1 U3914 ( .B1(n4103), .B2(n4748), .A(n3031), .ZN(U3581) );
  INV_X1 U3915 ( .A(DATAO_REG_7__SCAN_IN), .ZN(n4722) );
  NAND2_X1 U3916 ( .A1(U4043), .A2(n4460), .ZN(n3032) );
  OAI21_X1 U3917 ( .B1(U4043), .B2(n4722), .A(n3032), .ZN(U3557) );
  INV_X1 U3918 ( .A(DATAO_REG_0__SCAN_IN), .ZN(n4694) );
  NAND2_X1 U3919 ( .A1(U4043), .A2(n4473), .ZN(n3033) );
  OAI21_X1 U3920 ( .B1(U4043), .B2(n4694), .A(n3033), .ZN(U3550) );
  INV_X1 U3921 ( .A(DATAO_REG_5__SCAN_IN), .ZN(n4735) );
  NAND2_X1 U3922 ( .A1(U4043), .A2(n3403), .ZN(n3034) );
  OAI21_X1 U3923 ( .B1(U4043), .B2(n4735), .A(n3034), .ZN(U3555) );
  INV_X1 U3924 ( .A(DATAO_REG_6__SCAN_IN), .ZN(n4708) );
  NAND2_X1 U3925 ( .A1(U4043), .A2(n3341), .ZN(n3035) );
  OAI21_X1 U3926 ( .B1(U4043), .B2(n4708), .A(n3035), .ZN(U3556) );
  INV_X1 U3927 ( .A(DATAO_REG_30__SCAN_IN), .ZN(n4691) );
  INV_X1 U3928 ( .A(REG2_REG_30__SCAN_IN), .ZN(n4811) );
  NAND2_X1 U3929 ( .A1(n3036), .A2(REG1_REG_30__SCAN_IN), .ZN(n3039) );
  NAND2_X1 U3930 ( .A1(n3037), .A2(REG0_REG_30__SCAN_IN), .ZN(n3038) );
  OAI211_X1 U3931 ( .C1(n3040), .C2(n4811), .A(n3039), .B(n3038), .ZN(n4005)
         );
  NAND2_X1 U3932 ( .A1(U4043), .A2(n4005), .ZN(n3041) );
  OAI21_X1 U3933 ( .B1(U4043), .B2(n4691), .A(n3041), .ZN(U3580) );
  INV_X1 U3934 ( .A(DATAO_REG_15__SCAN_IN), .ZN(n4706) );
  NAND2_X1 U3935 ( .A1(n4570), .A2(n4103), .ZN(n3042) );
  OAI21_X1 U3936 ( .B1(U4043), .B2(n4706), .A(n3042), .ZN(U3565) );
  INV_X1 U3937 ( .A(DATAO_REG_14__SCAN_IN), .ZN(n4743) );
  NAND2_X1 U3938 ( .A1(n4562), .A2(n4103), .ZN(n3043) );
  OAI21_X1 U3939 ( .B1(U4043), .B2(n4743), .A(n3043), .ZN(U3564) );
  INV_X1 U3940 ( .A(DATAO_REG_17__SCAN_IN), .ZN(n4732) );
  NAND2_X1 U3941 ( .A1(n4350), .A2(n4103), .ZN(n3044) );
  OAI21_X1 U3942 ( .B1(n4103), .B2(n4732), .A(n3044), .ZN(U3567) );
  INV_X1 U3943 ( .A(REG2_REG_3__SCAN_IN), .ZN(n3377) );
  XNOR2_X1 U3944 ( .A(n3045), .B(n3377), .ZN(n3051) );
  INV_X1 U3945 ( .A(n3046), .ZN(n3047) );
  AOI211_X1 U3946 ( .C1(n3049), .C2(n3048), .A(n4970), .B(n3047), .ZN(n3050)
         );
  AOI21_X1 U3947 ( .B1(n4974), .B2(n3051), .A(n3050), .ZN(n3053) );
  AOI22_X1 U3948 ( .A1(n4994), .A2(ADDR_REG_3__SCAN_IN), .B1(
        REG3_REG_3__SCAN_IN), .B2(U3149), .ZN(n3052) );
  OAI211_X1 U3949 ( .C1(n3054), .C2(n5000), .A(n3053), .B(n3052), .ZN(U3243)
         );
  AOI211_X1 U3950 ( .C1(n3057), .C2(n3056), .A(n4970), .B(n3055), .ZN(n3065)
         );
  OAI211_X1 U3951 ( .C1(n3060), .C2(n3059), .A(n4974), .B(n3058), .ZN(n3062)
         );
  AND2_X1 U3952 ( .A1(U3149), .A2(REG3_REG_5__SCAN_IN), .ZN(n3297) );
  AOI21_X1 U3953 ( .B1(n4994), .B2(ADDR_REG_5__SCAN_IN), .A(n3297), .ZN(n3061)
         );
  OAI211_X1 U3954 ( .C1(n5000), .C2(n3063), .A(n3062), .B(n3061), .ZN(n3064)
         );
  OR2_X1 U3955 ( .A1(n3065), .A2(n3064), .ZN(U3245) );
  INV_X1 U3956 ( .A(n3066), .ZN(n3069) );
  INV_X1 U3957 ( .A(n3161), .ZN(n3072) );
  NAND2_X1 U3958 ( .A1(n5018), .A2(n3072), .ZN(n3073) );
  NAND2_X1 U3959 ( .A1(n3184), .A2(n4089), .ZN(n3215) );
  INV_X1 U3960 ( .A(n3215), .ZN(n3080) );
  NAND2_X1 U3961 ( .A1(n4600), .A2(n3074), .ZN(n3075) );
  NAND2_X1 U3962 ( .A1(n3076), .A2(n3075), .ZN(n3085) );
  NAND2_X1 U3963 ( .A1(n4572), .A2(n3085), .ZN(n3077) );
  NAND2_X1 U3964 ( .A1(n3184), .A2(n3077), .ZN(n3079) );
  NAND2_X1 U3965 ( .A1(n3079), .A2(n3078), .ZN(n3214) );
  NOR3_X1 U3966 ( .A1(n3080), .A2(n3214), .A3(n3086), .ZN(n3205) );
  NOR2_X1 U3967 ( .A1(n3086), .A2(n4572), .ZN(n3081) );
  NAND2_X1 U3968 ( .A1(n3082), .A2(n3081), .ZN(n3083) );
  NAND2_X1 U3969 ( .A1(n4089), .A2(n4947), .ZN(n3084) );
  OR2_X1 U3970 ( .A1(n3086), .A2(n3085), .ZN(n3087) );
  NAND2_X2 U3971 ( .A1(n3162), .A2(n3212), .ZN(n3174) );
  NAND2_X1 U3972 ( .A1(n3731), .A2(n4599), .ZN(n3089) );
  NAND2_X1 U3973 ( .A1(n3089), .A2(n3088), .ZN(n3165) );
  NOR2_X1 U3974 ( .A1(n3212), .A2(n2469), .ZN(n3090) );
  OR2_X2 U3975 ( .A1(n3165), .A2(n3090), .ZN(n3167) );
  OR2_X2 U3976 ( .A1(n3174), .A2(n3091), .ZN(n3289) );
  AOI22_X1 U3977 ( .A1(n3647), .A2(n4599), .B1(n3092), .B2(IR_REG_0__SCAN_IN), 
        .ZN(n3093) );
  OAI21_X1 U3978 ( .B1(n3289), .B2(n3203), .A(n3093), .ZN(n3168) );
  XNOR2_X1 U3979 ( .A(n3167), .B(n3168), .ZN(n3100) );
  OAI22_X1 U3980 ( .A1(n2984), .A2(n3898), .B1(n3913), .B2(n3100), .ZN(n3094)
         );
  AOI21_X1 U3981 ( .B1(n4599), .B2(n3908), .A(n3094), .ZN(n3095) );
  OAI21_X1 U3982 ( .B1(n3205), .B2(n3722), .A(n3095), .ZN(U3229) );
  NOR2_X1 U3983 ( .A1(n4947), .A2(n4950), .ZN(n3099) );
  AND2_X1 U3984 ( .A1(n4950), .A2(n4617), .ZN(n3096) );
  OR2_X1 U3985 ( .A1(n3096), .A2(n4947), .ZN(n4948) );
  NOR2_X1 U3986 ( .A1(n4090), .A2(n4617), .ZN(n3097) );
  MUX2_X1 U3987 ( .A(n4948), .B(n3097), .S(IR_REG_0__SCAN_IN), .Z(n3098) );
  AOI211_X1 U3988 ( .C1(n3100), .C2(n3099), .A(n3098), .B(n4100), .ZN(n3121)
         );
  OAI211_X1 U3989 ( .C1(n3103), .C2(n3102), .A(n4974), .B(n3101), .ZN(n3104)
         );
  INV_X1 U3990 ( .A(n3104), .ZN(n3113) );
  AOI211_X1 U3991 ( .C1(n3107), .C2(n3106), .A(n3105), .B(n4970), .ZN(n3112)
         );
  NOR2_X1 U3992 ( .A1(n3189), .A2(STATE_REG_SCAN_IN), .ZN(n3108) );
  AOI21_X1 U3993 ( .B1(n4994), .B2(ADDR_REG_2__SCAN_IN), .A(n3108), .ZN(n3109)
         );
  OAI21_X1 U3994 ( .B1(n5000), .B2(n3110), .A(n3109), .ZN(n3111) );
  OR4_X1 U3995 ( .A1(n3121), .A2(n3113), .A3(n3112), .A4(n3111), .ZN(U3242) );
  XNOR2_X1 U3996 ( .A(n3114), .B(REG2_REG_4__SCAN_IN), .ZN(n3124) );
  AOI211_X1 U3997 ( .C1(n3117), .C2(n3116), .A(n4970), .B(n3115), .ZN(n3122)
         );
  AND2_X1 U3998 ( .A1(U3149), .A2(REG3_REG_4__SCAN_IN), .ZN(n3240) );
  AOI21_X1 U3999 ( .B1(n4994), .B2(ADDR_REG_4__SCAN_IN), .A(n3240), .ZN(n3118)
         );
  OAI21_X1 U4000 ( .B1(n5000), .B2(n3119), .A(n3118), .ZN(n3120) );
  NOR3_X1 U4001 ( .A1(n3122), .A2(n3121), .A3(n3120), .ZN(n3123) );
  OAI21_X1 U4002 ( .B1(n3124), .B2(n4989), .A(n3123), .ZN(U3244) );
  INV_X1 U4003 ( .A(REG1_REG_1__SCAN_IN), .ZN(n3136) );
  OAI21_X1 U4004 ( .B1(n2907), .B2(n3126), .A(n3125), .ZN(n3132) );
  INV_X1 U4005 ( .A(n3132), .ZN(n4482) );
  INV_X1 U4006 ( .A(n2907), .ZN(n4015) );
  INV_X1 U4007 ( .A(n3941), .ZN(n3128) );
  OAI21_X1 U4008 ( .B1(n4015), .B2(n3128), .A(n3127), .ZN(n3129) );
  AOI22_X1 U4009 ( .A1(n4482), .A2(n3578), .B1(n3129), .B2(n4595), .ZN(n4485)
         );
  OAI22_X1 U4010 ( .A1(n3203), .A2(n4547), .B1(n3379), .B2(n4564), .ZN(n3130)
         );
  AOI21_X1 U4011 ( .B1(n4477), .B2(n4582), .A(n3130), .ZN(n3131) );
  OAI211_X1 U4012 ( .C1(n3571), .C2(n3132), .A(n4485), .B(n3131), .ZN(n3137)
         );
  NAND2_X1 U4013 ( .A1(n3137), .A2(n5043), .ZN(n3135) );
  AND2_X1 U4014 ( .A1(n4477), .A2(n4599), .ZN(n3133) );
  NOR2_X1 U4015 ( .A1(n3252), .A2(n3133), .ZN(n4479) );
  NAND2_X1 U4016 ( .A1(n4559), .A2(n4479), .ZN(n3134) );
  OAI211_X1 U4017 ( .C1(n5043), .C2(n3136), .A(n3135), .B(n3134), .ZN(U3519)
         );
  NAND2_X1 U4018 ( .A1(n3137), .A2(n5040), .ZN(n3139) );
  NAND2_X1 U4019 ( .A1(n4918), .A2(n4479), .ZN(n3138) );
  OAI211_X1 U4020 ( .C1(n5040), .C2(n4607), .A(n3139), .B(n3138), .ZN(U3469)
         );
  INV_X1 U4021 ( .A(DATAO_REG_21__SCAN_IN), .ZN(n4745) );
  NAND2_X1 U4022 ( .A1(n4269), .A2(n4103), .ZN(n3140) );
  OAI21_X1 U4023 ( .B1(n4103), .B2(n4745), .A(n3140), .ZN(U3571) );
  OAI22_X1 U4024 ( .A1(n3272), .A2(n4564), .B1(n2984), .B2(n4547), .ZN(n3141)
         );
  AOI21_X1 U4025 ( .B1(n3186), .B2(n4582), .A(n3141), .ZN(n3142) );
  OAI21_X1 U4026 ( .B1(n3143), .B2(n3571), .A(n3142), .ZN(n3145) );
  NOR2_X1 U4027 ( .A1(n3145), .A2(n3144), .ZN(n3150) );
  INV_X1 U4028 ( .A(n3146), .ZN(n3148) );
  AOI22_X1 U4029 ( .A1(n4559), .A2(n3148), .B1(n2210), .B2(REG1_REG_2__SCAN_IN), .ZN(n3147) );
  OAI21_X1 U4030 ( .B1(n3150), .B2(n2210), .A(n3147), .ZN(U3520) );
  AOI22_X1 U4031 ( .A1(n4918), .A2(n3148), .B1(n5039), .B2(REG0_REG_2__SCAN_IN), .ZN(n3149) );
  OAI21_X1 U4032 ( .B1(n3150), .B2(n5039), .A(n3149), .ZN(U3471) );
  XOR2_X1 U4033 ( .A(REG1_REG_7__SCAN_IN), .B(n4941), .Z(n3151) );
  XNOR2_X1 U4034 ( .A(n3152), .B(n3151), .ZN(n3159) );
  INV_X1 U4035 ( .A(n5000), .ZN(n4158) );
  INV_X1 U4036 ( .A(ADDR_REG_7__SCAN_IN), .ZN(n4854) );
  NAND2_X1 U4037 ( .A1(REG3_REG_7__SCAN_IN), .A2(U3149), .ZN(n3357) );
  OAI211_X1 U4038 ( .C1(n3155), .C2(n3154), .A(n3153), .B(n4974), .ZN(n3156)
         );
  OAI211_X1 U4039 ( .C1(n4978), .C2(n4854), .A(n3357), .B(n3156), .ZN(n3157)
         );
  AOI21_X1 U4040 ( .B1(n4158), .B2(n4941), .A(n3157), .ZN(n3158) );
  OAI21_X1 U4041 ( .B1(n3159), .B2(n4970), .A(n3158), .ZN(U3247) );
  NAND2_X1 U4042 ( .A1(n3731), .A2(n4477), .ZN(n3160) );
  OAI21_X1 U40430 ( .B1(n2984), .B2(n3753), .A(n3160), .ZN(n3163) );
  XNOR2_X1 U4044 ( .A(n3163), .B(n3754), .ZN(n3169) );
  OAI22_X1 U4045 ( .A1(n2984), .A2(n3289), .B1(n3164), .B2(n3753), .ZN(n3170)
         );
  XNOR2_X1 U4046 ( .A(n3169), .B(n3170), .ZN(n3202) );
  INV_X1 U4047 ( .A(n3165), .ZN(n3166) );
  AOI22_X1 U4048 ( .A1(n3168), .A2(n3167), .B1(n3658), .B2(n3166), .ZN(n3201)
         );
  NOR2_X1 U4049 ( .A1(n3202), .A2(n3201), .ZN(n3172) );
  AND2_X1 U4050 ( .A1(n3170), .A2(n3169), .ZN(n3171) );
  NOR2_X2 U4051 ( .A1(n3172), .A2(n3171), .ZN(n3180) );
  OAI21_X1 U4052 ( .B1(n3174), .B2(n3251), .A(n3173), .ZN(n3175) );
  XNOR2_X1 U4053 ( .A(n3175), .B(n3754), .ZN(n3177) );
  OAI22_X1 U4054 ( .A1(n3289), .A2(n3379), .B1(n3251), .B2(n3753), .ZN(n3176)
         );
  NOR2_X1 U4055 ( .A1(n3177), .A2(n3176), .ZN(n3220) );
  NOR2_X1 U4056 ( .A1(n3220), .A2(n3178), .ZN(n3179) );
  NAND2_X1 U4057 ( .A1(n3180), .A2(n3179), .ZN(n3222) );
  OAI21_X1 U4058 ( .B1(n3180), .B2(n3179), .A(n3222), .ZN(n3181) );
  NAND2_X1 U4059 ( .A1(n3181), .A2(n3920), .ZN(n3188) );
  NAND2_X1 U4060 ( .A1(n4089), .A2(n3182), .ZN(n3183) );
  OAI22_X1 U4061 ( .A1(n3272), .A2(n3898), .B1(n3923), .B2(n2984), .ZN(n3185)
         );
  AOI21_X1 U4062 ( .B1(n3186), .B2(n3908), .A(n3185), .ZN(n3187) );
  OAI211_X1 U4063 ( .C1(n3205), .C2(n3189), .A(n3188), .B(n3187), .ZN(U3234)
         );
  INV_X1 U4064 ( .A(REG2_REG_6__SCAN_IN), .ZN(n3409) );
  XNOR2_X1 U4065 ( .A(n3190), .B(n3409), .ZN(n3197) );
  OAI211_X1 U4066 ( .C1(n3192), .C2(REG1_REG_6__SCAN_IN), .A(n3191), .B(n4996), 
        .ZN(n3194) );
  AND2_X1 U4067 ( .A1(U3149), .A2(REG3_REG_6__SCAN_IN), .ZN(n3329) );
  AOI21_X1 U4068 ( .B1(n4994), .B2(ADDR_REG_6__SCAN_IN), .A(n3329), .ZN(n3193)
         );
  OAI211_X1 U4069 ( .C1(n5000), .C2(n3195), .A(n3194), .B(n3193), .ZN(n3196)
         );
  AOI21_X1 U4070 ( .B1(n4974), .B2(n3197), .A(n3196), .ZN(n3198) );
  INV_X1 U4071 ( .A(n3198), .ZN(U3246) );
  INV_X1 U4072 ( .A(DATAO_REG_22__SCAN_IN), .ZN(n4730) );
  NAND2_X1 U4073 ( .A1(n3199), .A2(n4103), .ZN(n3200) );
  OAI21_X1 U4074 ( .B1(U4043), .B2(n4730), .A(n3200), .ZN(U3572) );
  XNOR2_X1 U4075 ( .A(n3202), .B(n3201), .ZN(n3209) );
  OAI22_X1 U4076 ( .A1(n3379), .A2(n3898), .B1(n3923), .B2(n3203), .ZN(n3207)
         );
  NOR2_X1 U4077 ( .A1(n3205), .A2(n3204), .ZN(n3206) );
  AOI211_X1 U4078 ( .C1(n4477), .C2(n3908), .A(n3207), .B(n3206), .ZN(n3208)
         );
  OAI21_X1 U4079 ( .B1(n3209), .B2(n3913), .A(n3208), .ZN(U3219) );
  OAI22_X1 U4080 ( .A1(n3210), .A2(n3898), .B1(n3923), .B2(n3379), .ZN(n3218)
         );
  NAND2_X1 U4081 ( .A1(n3212), .A2(n3211), .ZN(n3213) );
  OAI21_X1 U4082 ( .B1(n3214), .B2(n3213), .A(STATE_REG_SCAN_IN), .ZN(n3216)
         );
  MUX2_X1 U4083 ( .A(n3889), .B(U3149), .S(REG3_REG_3__SCAN_IN), .Z(n3217) );
  AOI211_X1 U4084 ( .C1(n3253), .C2(n3908), .A(n3218), .B(n3217), .ZN(n3227)
         );
  OAI22_X1 U4085 ( .A1(n3289), .A2(n3272), .B1(n3378), .B2(n3753), .ZN(n3228)
         );
  OAI22_X1 U4086 ( .A1(n3272), .A2(n3753), .B1(n3378), .B2(n3174), .ZN(n3219)
         );
  XNOR2_X1 U4087 ( .A(n3219), .B(n3754), .ZN(n3229) );
  XOR2_X1 U4088 ( .A(n3228), .B(n3229), .Z(n3224) );
  INV_X1 U4089 ( .A(n3220), .ZN(n3221) );
  NAND2_X1 U4090 ( .A1(n3222), .A2(n3221), .ZN(n3223) );
  OAI21_X1 U4091 ( .B1(n3224), .B2(n3223), .A(n3236), .ZN(n3225) );
  NAND2_X1 U4092 ( .A1(n3225), .A2(n3920), .ZN(n3226) );
  NAND2_X1 U4093 ( .A1(n3227), .A2(n3226), .ZN(U3215) );
  OR2_X1 U4094 ( .A1(n3229), .A2(n3228), .ZN(n3234) );
  AND2_X1 U4095 ( .A1(n3236), .A2(n3234), .ZN(n3238) );
  NAND2_X1 U4096 ( .A1(n3731), .A2(n3269), .ZN(n3230) );
  OAI21_X1 U4097 ( .B1(n3210), .B2(n3753), .A(n3230), .ZN(n3231) );
  XNOR2_X1 U4098 ( .A(n3231), .B(n3658), .ZN(n3290) );
  NAND2_X1 U4099 ( .A1(n3647), .A2(n3269), .ZN(n3233) );
  OAI21_X1 U4100 ( .B1(n3289), .B2(n3210), .A(n3233), .ZN(n3291) );
  XNOR2_X1 U4101 ( .A(n3290), .B(n3291), .ZN(n3237) );
  OAI211_X1 U4102 ( .C1(n3238), .C2(n3237), .A(n3920), .B(n3294), .ZN(n3242)
         );
  OAI22_X1 U4103 ( .A1(n3925), .A2(n3279), .B1(n3272), .B2(n3923), .ZN(n3239)
         );
  AOI211_X1 U4104 ( .C1(n3927), .C2(n3403), .A(n3240), .B(n3239), .ZN(n3241)
         );
  OAI211_X1 U4105 ( .C1(n3931), .C2(n3270), .A(n3242), .B(n3241), .ZN(U3227)
         );
  NAND2_X1 U4106 ( .A1(n3244), .A2(n3243), .ZN(n3273) );
  INV_X1 U4107 ( .A(n4014), .ZN(n3245) );
  XNOR2_X1 U4108 ( .A(n3273), .B(n3245), .ZN(n3383) );
  OAI22_X1 U4109 ( .A1(n3379), .A2(n4547), .B1(n3378), .B2(n4572), .ZN(n3250)
         );
  OAI21_X1 U4110 ( .B1(n4014), .B2(n3247), .A(n3246), .ZN(n3248) );
  AOI22_X1 U4111 ( .A1(n3248), .A2(n4595), .B1(n4601), .B2(n4105), .ZN(n3386)
         );
  INV_X1 U4112 ( .A(n3386), .ZN(n3249) );
  AOI211_X1 U4113 ( .C1(n4596), .C2(n3383), .A(n3250), .B(n3249), .ZN(n3258)
         );
  NAND2_X1 U4114 ( .A1(n3252), .A2(n3251), .ZN(n3254) );
  NAND2_X1 U4115 ( .A1(n3254), .A2(n3253), .ZN(n3255) );
  AND2_X1 U4116 ( .A1(n3255), .A2(n3268), .ZN(n3382) );
  AOI22_X1 U4117 ( .A1(n4559), .A2(n3382), .B1(n2210), .B2(REG1_REG_3__SCAN_IN), .ZN(n3256) );
  OAI21_X1 U4118 ( .B1(n3258), .B2(n2210), .A(n3256), .ZN(U3521) );
  AOI22_X1 U4119 ( .A1(n4918), .A2(n3382), .B1(n5039), .B2(REG0_REG_3__SCAN_IN), .ZN(n3257) );
  OAI21_X1 U4120 ( .B1(n3258), .B2(n5039), .A(n3257), .ZN(U3473) );
  XNOR2_X1 U4121 ( .A(n3259), .B(REG1_REG_8__SCAN_IN), .ZN(n3267) );
  XOR2_X1 U4122 ( .A(n3260), .B(REG2_REG_8__SCAN_IN), .Z(n3261) );
  NAND2_X1 U4123 ( .A1(n4974), .A2(n3261), .ZN(n3262) );
  NAND2_X1 U4124 ( .A1(REG3_REG_8__SCAN_IN), .A2(U3149), .ZN(n3396) );
  NAND2_X1 U4125 ( .A1(n3262), .A2(n3396), .ZN(n3265) );
  NOR2_X1 U4126 ( .A1(n5000), .A2(n3263), .ZN(n3264) );
  AOI211_X1 U4127 ( .C1(n4994), .C2(ADDR_REG_8__SCAN_IN), .A(n3265), .B(n3264), 
        .ZN(n3266) );
  OAI21_X1 U4128 ( .B1(n3267), .B2(n4970), .A(n3266), .ZN(U3248) );
  INV_X1 U4129 ( .A(n4359), .ZN(n5032) );
  AOI211_X1 U4130 ( .C1(n3269), .C2(n3268), .A(n5032), .B(n3307), .ZN(n5030)
         );
  NOR2_X1 U4131 ( .A1(n4461), .A2(n3270), .ZN(n3283) );
  INV_X1 U4132 ( .A(n3273), .ZN(n3275) );
  OAI21_X1 U4133 ( .B1(n3273), .B2(n3272), .A(n3378), .ZN(n3274) );
  OAI21_X1 U4134 ( .B1(n3275), .B2(n2909), .A(n3274), .ZN(n3276) );
  XOR2_X1 U4135 ( .A(n3271), .B(n3276), .Z(n3284) );
  XOR2_X1 U4136 ( .A(n3271), .B(n3277), .Z(n3281) );
  AOI22_X1 U4137 ( .A1(n4601), .A2(n3403), .B1(n2909), .B2(n4584), .ZN(n3278)
         );
  OAI21_X1 U4138 ( .B1(n3279), .B2(n4572), .A(n3278), .ZN(n3280) );
  AOI21_X1 U4139 ( .B1(n3281), .B2(n4595), .A(n3280), .ZN(n3282) );
  OAI21_X1 U4140 ( .B1(n3284), .B2(n4418), .A(n3282), .ZN(n5029) );
  AOI211_X1 U4141 ( .C1(n5030), .C2(n3346), .A(n3283), .B(n5029), .ZN(n3286)
         );
  INV_X1 U4142 ( .A(n3284), .ZN(n5031) );
  AOI22_X1 U4143 ( .A1(n5031), .A2(n4483), .B1(REG2_REG_4__SCAN_IN), .B2(n4454), .ZN(n3285) );
  OAI21_X1 U4144 ( .B1(n3286), .B2(n4454), .A(n3285), .ZN(U3286) );
  OR2_X1 U4145 ( .A1(n3753), .A2(n3327), .ZN(n3287) );
  OAI21_X1 U4146 ( .B1(n3174), .B2(n3306), .A(n3287), .ZN(n3288) );
  XNOR2_X1 U4147 ( .A(n3288), .B(n3658), .ZN(n3312) );
  OAI22_X1 U4148 ( .A1(n3289), .A2(n3327), .B1(n3753), .B2(n3306), .ZN(n3313)
         );
  XNOR2_X1 U4149 ( .A(n3312), .B(n3313), .ZN(n3315) );
  INV_X1 U4150 ( .A(n3290), .ZN(n3292) );
  NAND2_X1 U4151 ( .A1(n3292), .A2(n3291), .ZN(n3293) );
  XOR2_X1 U4152 ( .A(n3315), .B(n3316), .Z(n3295) );
  NAND2_X1 U4153 ( .A1(n3295), .A2(n3920), .ZN(n3299) );
  OAI22_X1 U4154 ( .A1(n3925), .A2(n3306), .B1(n3210), .B2(n3923), .ZN(n3296)
         );
  AOI211_X1 U4155 ( .C1(n3927), .C2(n3341), .A(n3297), .B(n3296), .ZN(n3298)
         );
  OAI211_X1 U4156 ( .C1(n3931), .C2(n3436), .A(n3299), .B(n3298), .ZN(U3224)
         );
  INV_X1 U4157 ( .A(DATAO_REG_24__SCAN_IN), .ZN(n4715) );
  NAND2_X1 U4158 ( .A1(n4504), .A2(n4103), .ZN(n3300) );
  OAI21_X1 U4159 ( .B1(U4043), .B2(n4715), .A(n3300), .ZN(U3574) );
  AND2_X1 U4160 ( .A1(n2180), .A2(n3967), .ZN(n4016) );
  XNOR2_X1 U4161 ( .A(n3301), .B(n4016), .ZN(n3439) );
  AOI22_X1 U4162 ( .A1(n4105), .A2(n4584), .B1(n4601), .B2(n3341), .ZN(n3302)
         );
  OAI21_X1 U4163 ( .B1(n3306), .B2(n4572), .A(n3302), .ZN(n3305) );
  XNOR2_X1 U4164 ( .A(n3303), .B(n4016), .ZN(n3304) );
  NOR2_X1 U4165 ( .A1(n3304), .A2(n4441), .ZN(n3445) );
  AOI211_X1 U4166 ( .C1(n3439), .C2(n4596), .A(n3305), .B(n3445), .ZN(n3311)
         );
  OR2_X1 U4167 ( .A1(n3307), .A2(n3306), .ZN(n3308) );
  AND2_X1 U4168 ( .A1(n3410), .A2(n3308), .ZN(n3438) );
  AOI22_X1 U4169 ( .A1(n4918), .A2(n3438), .B1(n5039), .B2(REG0_REG_5__SCAN_IN), .ZN(n3309) );
  OAI21_X1 U4170 ( .B1(n3311), .B2(n5039), .A(n3309), .ZN(U3477) );
  AOI22_X1 U4171 ( .A1(n4559), .A2(n3438), .B1(n2210), .B2(REG1_REG_5__SCAN_IN), .ZN(n3310) );
  OAI21_X1 U4172 ( .B1(n3311), .B2(n2210), .A(n3310), .ZN(U3523) );
  INV_X1 U4173 ( .A(n3312), .ZN(n3314) );
  NAND2_X1 U4174 ( .A1(n3731), .A2(n3320), .ZN(n3318) );
  NAND2_X1 U4175 ( .A1(n3647), .A2(n3341), .ZN(n3317) );
  NAND2_X1 U4176 ( .A1(n3318), .A2(n3317), .ZN(n3319) );
  XNOR2_X1 U4177 ( .A(n3319), .B(n3658), .ZN(n3323) );
  INV_X1 U4178 ( .A(n3323), .ZN(n3322) );
  AOI22_X1 U4179 ( .A1(n3735), .A2(n3341), .B1(n3232), .B2(n3320), .ZN(n3324)
         );
  INV_X1 U4180 ( .A(n3324), .ZN(n3321) );
  AND2_X1 U4181 ( .A1(n3324), .A2(n3323), .ZN(n3351) );
  NOR2_X1 U4182 ( .A1(n2184), .A2(n3351), .ZN(n3325) );
  XNOR2_X1 U4183 ( .A(n3352), .B(n3325), .ZN(n3326) );
  NAND2_X1 U4184 ( .A1(n3326), .A2(n3920), .ZN(n3331) );
  OAI22_X1 U4185 ( .A1(n3925), .A2(n3411), .B1(n3327), .B2(n3923), .ZN(n3328)
         );
  AOI211_X1 U4186 ( .C1(n3927), .C2(n4460), .A(n3329), .B(n3328), .ZN(n3330)
         );
  OAI211_X1 U4187 ( .C1(n3931), .C2(n3408), .A(n3331), .B(n3330), .ZN(U3236)
         );
  INV_X1 U4188 ( .A(n3332), .ZN(n3333) );
  OAI21_X1 U4189 ( .B1(n3333), .B2(n2723), .A(n3411), .ZN(n3334) );
  OAI21_X1 U4190 ( .B1(n3341), .B2(n3332), .A(n3334), .ZN(n3335) );
  XNOR2_X1 U4191 ( .A(n3335), .B(n3338), .ZN(n3420) );
  INV_X1 U4192 ( .A(n3420), .ZN(n3350) );
  NAND2_X1 U4193 ( .A1(n4418), .A2(n3336), .ZN(n3337) );
  INV_X1 U4194 ( .A(n3338), .ZN(n4020) );
  XNOR2_X1 U4195 ( .A(n3339), .B(n4020), .ZN(n3340) );
  NAND2_X1 U4196 ( .A1(n3340), .A2(n4595), .ZN(n3343) );
  AOI22_X1 U4197 ( .A1(n4104), .A2(n4601), .B1(n4584), .B2(n3341), .ZN(n3342)
         );
  OAI211_X1 U4198 ( .C1(n4572), .C2(n3358), .A(n3343), .B(n3342), .ZN(n3418)
         );
  NAND2_X1 U4199 ( .A1(n3418), .A2(n4484), .ZN(n3349) );
  INV_X1 U4200 ( .A(n3430), .ZN(n3344) );
  AOI211_X1 U4201 ( .C1(n3345), .C2(n3413), .A(n5032), .B(n3344), .ZN(n3419)
         );
  NAND2_X1 U4202 ( .A1(n4484), .A2(n3346), .ZN(n4362) );
  INV_X1 U4203 ( .A(n4362), .ZN(n3721) );
  OAI22_X1 U4204 ( .A1(n4484), .A2(n2588), .B1(n3363), .B2(n4461), .ZN(n3347)
         );
  AOI21_X1 U4205 ( .B1(n3419), .B2(n3721), .A(n3347), .ZN(n3348) );
  OAI211_X1 U4206 ( .C1(n3350), .C2(n4304), .A(n3349), .B(n3348), .ZN(U3283)
         );
  OAI22_X1 U4207 ( .A1(n3358), .A2(n3174), .B1(n3354), .B2(n3753), .ZN(n3353)
         );
  XNOR2_X1 U4208 ( .A(n3353), .B(n3754), .ZN(n3388) );
  OAI22_X1 U4209 ( .A1(n3354), .A2(n3289), .B1(n3358), .B2(n3753), .ZN(n3387)
         );
  XOR2_X1 U4210 ( .A(n3388), .B(n3387), .Z(n3355) );
  OAI211_X1 U4211 ( .C1(n3356), .C2(n3355), .A(n3391), .B(n3920), .ZN(n3362)
         );
  INV_X1 U4212 ( .A(n3357), .ZN(n3360) );
  OAI22_X1 U4213 ( .A1(n3925), .A2(n3358), .B1(n2723), .B2(n3923), .ZN(n3359)
         );
  AOI211_X1 U4214 ( .C1(n3927), .C2(n4104), .A(n3360), .B(n3359), .ZN(n3361)
         );
  OAI211_X1 U4215 ( .C1(n3931), .C2(n3363), .A(n3362), .B(n3361), .ZN(U3210)
         );
  MUX2_X1 U4216 ( .A(REG1_REG_9__SCAN_IN), .B(n4838), .S(n3364), .Z(n3366) );
  OAI211_X1 U4217 ( .C1(n3367), .C2(n3366), .A(n4996), .B(n3365), .ZN(n3374)
         );
  NOR2_X1 U4218 ( .A1(STATE_REG_SCAN_IN), .A2(n2737), .ZN(n3537) );
  INV_X1 U4219 ( .A(ADDR_REG_9__SCAN_IN), .ZN(n4852) );
  XOR2_X1 U4220 ( .A(n3369), .B(n3368), .Z(n3370) );
  NAND2_X1 U4221 ( .A1(n3370), .A2(n4974), .ZN(n3371) );
  OAI21_X1 U4222 ( .B1(n4978), .B2(n4852), .A(n3371), .ZN(n3372) );
  NOR2_X1 U4223 ( .A1(n3537), .A2(n3372), .ZN(n3373) );
  OAI211_X1 U4224 ( .C1(n5000), .C2(n3375), .A(n3374), .B(n3373), .ZN(U3249)
         );
  INV_X1 U4225 ( .A(DATAO_REG_25__SCAN_IN), .ZN(n4729) );
  NAND2_X1 U4226 ( .A1(n4237), .A2(n4103), .ZN(n3376) );
  OAI21_X1 U4227 ( .B1(U4043), .B2(n4729), .A(n3376), .ZN(U3575) );
  OAI22_X1 U4228 ( .A1(n4484), .A2(n3377), .B1(REG3_REG_3__SCAN_IN), .B2(n4461), .ZN(n3381) );
  OAI22_X1 U4229 ( .A1(n3379), .A2(n4293), .B1(n4424), .B2(n3378), .ZN(n3380)
         );
  AOI211_X1 U4230 ( .C1(n4480), .C2(n3382), .A(n3381), .B(n3380), .ZN(n3385)
         );
  NAND2_X1 U4231 ( .A1(n4467), .A2(n3383), .ZN(n3384) );
  OAI211_X1 U4232 ( .C1(n4386), .C2(n3386), .A(n3385), .B(n3384), .ZN(U3287)
         );
  INV_X1 U4233 ( .A(n3387), .ZN(n3390) );
  INV_X1 U4234 ( .A(n3388), .ZN(n3389) );
  OR2_X1 U4235 ( .A1(n3753), .A2(n3534), .ZN(n3393) );
  OAI21_X1 U4236 ( .B1(n3174), .B2(n3428), .A(n3393), .ZN(n3394) );
  XNOR2_X1 U4237 ( .A(n3394), .B(n3754), .ZN(n3503) );
  OAI22_X1 U4238 ( .A1(n3289), .A2(n3534), .B1(n3428), .B2(n3753), .ZN(n3530)
         );
  INV_X1 U4239 ( .A(n3530), .ZN(n3528) );
  XNOR2_X1 U4240 ( .A(n3503), .B(n3528), .ZN(n3395) );
  XNOR2_X1 U4241 ( .A(n3392), .B(n3395), .ZN(n3401) );
  INV_X1 U4242 ( .A(n4462), .ZN(n3399) );
  AOI22_X1 U4243 ( .A1(n4458), .A2(n3908), .B1(n3906), .B2(n4460), .ZN(n3397)
         );
  OAI211_X1 U4244 ( .C1(n3478), .C2(n3898), .A(n3397), .B(n3396), .ZN(n3398)
         );
  AOI21_X1 U4245 ( .B1(n3399), .B2(n3889), .A(n3398), .ZN(n3400) );
  OAI21_X1 U4246 ( .B1(n3401), .B2(n3913), .A(n3400), .ZN(U3218) );
  AND2_X1 U4247 ( .A1(n3955), .A2(n3968), .ZN(n4019) );
  XOR2_X1 U4248 ( .A(n4019), .B(n3402), .Z(n3407) );
  XNOR2_X1 U4249 ( .A(n3332), .B(n4019), .ZN(n5038) );
  AOI22_X1 U4250 ( .A1(n4601), .A2(n4460), .B1(n3403), .B2(n4584), .ZN(n3404)
         );
  OAI21_X1 U4251 ( .B1(n3411), .B2(n4572), .A(n3404), .ZN(n3405) );
  AOI21_X1 U4252 ( .B1(n5038), .B2(n3578), .A(n3405), .ZN(n3406) );
  OAI21_X1 U4253 ( .B1(n3407), .B2(n4441), .A(n3406), .ZN(n5035) );
  INV_X1 U4254 ( .A(n5035), .ZN(n3417) );
  OAI22_X1 U4255 ( .A1(n4484), .A2(n3409), .B1(n3408), .B2(n4461), .ZN(n3415)
         );
  INV_X1 U4256 ( .A(n3410), .ZN(n3412) );
  NOR2_X1 U4257 ( .A1(n3412), .A2(n3411), .ZN(n5034) );
  INV_X1 U4258 ( .A(n3413), .ZN(n5033) );
  NOR3_X1 U4259 ( .A1(n5034), .A2(n4449), .A3(n5033), .ZN(n3414) );
  AOI211_X1 U4260 ( .C1(n5038), .C2(n4483), .A(n3415), .B(n3414), .ZN(n3416)
         );
  OAI21_X1 U4261 ( .B1(n3417), .B2(n4454), .A(n3416), .ZN(U3284) );
  AOI211_X1 U4262 ( .C1(n4596), .C2(n3420), .A(n3419), .B(n3418), .ZN(n3423)
         );
  NAND2_X1 U4263 ( .A1(n2210), .A2(REG1_REG_7__SCAN_IN), .ZN(n3421) );
  OAI21_X1 U4264 ( .B1(n3423), .B2(n2210), .A(n3421), .ZN(U3525) );
  NAND2_X1 U4265 ( .A1(n5039), .A2(REG0_REG_7__SCAN_IN), .ZN(n3422) );
  OAI21_X1 U4266 ( .B1(n3423), .B2(n5039), .A(n3422), .ZN(U3481) );
  AND2_X1 U4267 ( .A1(n3958), .A2(n3969), .ZN(n4029) );
  XOR2_X1 U4268 ( .A(n3424), .B(n4029), .Z(n4457) );
  XNOR2_X1 U4269 ( .A(n3425), .B(n4029), .ZN(n4468) );
  NAND2_X1 U4270 ( .A1(n4468), .A2(n4596), .ZN(n3427) );
  AOI22_X1 U4271 ( .A1(n4460), .A2(n4584), .B1(n4601), .B2(n4459), .ZN(n3426)
         );
  OAI211_X1 U4272 ( .C1(n4572), .C2(n3428), .A(n3427), .B(n3426), .ZN(n3429)
         );
  AOI21_X1 U4273 ( .B1(n4457), .B2(n4595), .A(n3429), .ZN(n3434) );
  AND2_X1 U4274 ( .A1(n3430), .A2(n4458), .ZN(n3431) );
  NOR2_X1 U4275 ( .A1(n3451), .A2(n3431), .ZN(n4466) );
  AOI22_X1 U4276 ( .A1(n4466), .A2(n4559), .B1(REG1_REG_8__SCAN_IN), .B2(n2210), .ZN(n3432) );
  OAI21_X1 U4277 ( .B1(n3434), .B2(n2210), .A(n3432), .ZN(U3526) );
  AOI22_X1 U4278 ( .A1(n4466), .A2(n4918), .B1(REG0_REG_8__SCAN_IN), .B2(n5039), .ZN(n3433) );
  OAI21_X1 U4279 ( .B1(n3434), .B2(n5039), .A(n3433), .ZN(U3483) );
  AOI22_X1 U4280 ( .A1(n4478), .A2(n3435), .B1(n4474), .B2(n4105), .ZN(n3443)
         );
  OAI22_X1 U4281 ( .A1(n4484), .A2(n2694), .B1(n3436), .B2(n4461), .ZN(n3437)
         );
  AOI21_X1 U4282 ( .B1(n4480), .B2(n3438), .A(n3437), .ZN(n3442) );
  OR2_X1 U4283 ( .A1(n4295), .A2(n2723), .ZN(n3441) );
  NAND2_X1 U4284 ( .A1(n3439), .A2(n4467), .ZN(n3440) );
  NAND4_X1 U4285 ( .A1(n3443), .A2(n3442), .A3(n3441), .A4(n3440), .ZN(n3444)
         );
  AOI21_X1 U4286 ( .B1(n3445), .B2(n4484), .A(n3444), .ZN(n3446) );
  INV_X1 U4287 ( .A(n3446), .ZN(U3285) );
  AND2_X1 U4288 ( .A1(n2912), .A2(n3959), .ZN(n4030) );
  XNOR2_X1 U4289 ( .A(n3448), .B(n4030), .ZN(n3449) );
  NOR2_X1 U4290 ( .A1(n3449), .A2(n4441), .ZN(n3490) );
  INV_X1 U4291 ( .A(n3490), .ZN(n3459) );
  XNOR2_X1 U4292 ( .A(n3450), .B(n4030), .ZN(n3492) );
  OR2_X1 U4293 ( .A1(n3451), .A2(n3535), .ZN(n3452) );
  NAND2_X1 U4294 ( .A1(n3471), .A2(n3452), .ZN(n3524) );
  OAI22_X1 U4295 ( .A1(n4484), .A2(n3453), .B1(n3540), .B2(n4461), .ZN(n3455)
         );
  OAI22_X1 U4296 ( .A1(n4293), .A2(n3534), .B1(n3509), .B2(n4295), .ZN(n3454)
         );
  AOI211_X1 U4297 ( .C1(n3499), .C2(n4478), .A(n3455), .B(n3454), .ZN(n3456)
         );
  OAI21_X1 U4298 ( .B1(n4449), .B2(n3524), .A(n3456), .ZN(n3457) );
  AOI21_X1 U4299 ( .B1(n4467), .B2(n3492), .A(n3457), .ZN(n3458) );
  OAI21_X1 U4300 ( .B1(n3459), .B2(n4454), .A(n3458), .ZN(U3281) );
  INV_X1 U4301 ( .A(DATAO_REG_27__SCAN_IN), .ZN(n4686) );
  NAND2_X1 U4302 ( .A1(n4203), .A2(n4103), .ZN(n3460) );
  OAI21_X1 U4303 ( .B1(U4043), .B2(n4686), .A(n3460), .ZN(U3577) );
  AND2_X1 U4304 ( .A1(U3149), .A2(REG3_REG_10__SCAN_IN), .ZN(n3564) );
  INV_X1 U4305 ( .A(ADDR_REG_10__SCAN_IN), .ZN(n4836) );
  XOR2_X1 U4306 ( .A(REG2_REG_10__SCAN_IN), .B(n3461), .Z(n3462) );
  NAND2_X1 U4307 ( .A1(n3462), .A2(n4974), .ZN(n3463) );
  OAI21_X1 U4308 ( .B1(n4978), .B2(n4836), .A(n3463), .ZN(n3464) );
  AOI211_X1 U4309 ( .C1(n4158), .C2(n3465), .A(n3564), .B(n3464), .ZN(n3466)
         );
  OAI21_X1 U4310 ( .B1(n3467), .B2(n4970), .A(n3466), .ZN(U3250) );
  AND2_X1 U4311 ( .A1(n3971), .A2(n3974), .ZN(n4031) );
  XNOR2_X1 U4312 ( .A(n3468), .B(n4031), .ZN(n3482) );
  XNOR2_X1 U4313 ( .A(n3469), .B(n4031), .ZN(n3484) );
  NOR2_X1 U4314 ( .A1(n4454), .A2(n4441), .ZN(n4456) );
  NAND2_X1 U4315 ( .A1(n3484), .A2(n4456), .ZN(n3477) );
  INV_X1 U4316 ( .A(n3470), .ZN(n3570) );
  AOI21_X1 U4317 ( .B1(n3480), .B2(n3471), .A(n3570), .ZN(n3486) );
  AOI22_X1 U4318 ( .A1(n3480), .A2(n4478), .B1(n4474), .B2(n4459), .ZN(n3474)
         );
  INV_X1 U4319 ( .A(n3567), .ZN(n3472) );
  INV_X1 U4320 ( .A(n4461), .ZN(n4481) );
  AOI22_X1 U4321 ( .A1(n4454), .A2(REG2_REG_10__SCAN_IN), .B1(n3472), .B2(
        n4481), .ZN(n3473) );
  OAI211_X1 U4322 ( .C1(n3781), .C2(n4295), .A(n3474), .B(n3473), .ZN(n3475)
         );
  AOI21_X1 U4323 ( .B1(n3486), .B2(n4480), .A(n3475), .ZN(n3476) );
  OAI211_X1 U4324 ( .C1(n4304), .C2(n3482), .A(n3477), .B(n3476), .ZN(U3280)
         );
  OAI22_X1 U4325 ( .A1(n3478), .A2(n4547), .B1(n3781), .B2(n4564), .ZN(n3479)
         );
  AOI21_X1 U4326 ( .B1(n3480), .B2(n4582), .A(n3479), .ZN(n3481) );
  OAI21_X1 U4327 ( .B1(n3482), .B2(n4543), .A(n3481), .ZN(n3483) );
  AOI21_X1 U4328 ( .B1(n3484), .B2(n4595), .A(n3483), .ZN(n3488) );
  AOI22_X1 U4329 ( .A1(n3486), .A2(n4559), .B1(REG1_REG_10__SCAN_IN), .B2(
        n2210), .ZN(n3485) );
  OAI21_X1 U4330 ( .B1(n3488), .B2(n2210), .A(n3485), .ZN(U3528) );
  AOI22_X1 U4331 ( .A1(n3486), .A2(n4918), .B1(REG0_REG_10__SCAN_IN), .B2(
        n5039), .ZN(n3487) );
  OAI21_X1 U4332 ( .B1(n3488), .B2(n5039), .A(n3487), .ZN(U3487) );
  AOI22_X1 U4333 ( .A1(n4584), .A2(n4104), .B1(n4102), .B2(n4601), .ZN(n3489)
         );
  OAI21_X1 U4334 ( .B1(n3535), .B2(n4572), .A(n3489), .ZN(n3491) );
  AOI211_X1 U4335 ( .C1(n3492), .C2(n4596), .A(n3491), .B(n3490), .ZN(n3522)
         );
  OAI22_X1 U4336 ( .A1(n3524), .A2(n4936), .B1(n5040), .B2(n3493), .ZN(n3494)
         );
  INV_X1 U4337 ( .A(n3494), .ZN(n3495) );
  OAI21_X1 U4338 ( .B1(n3522), .B2(n5039), .A(n3495), .ZN(U3485) );
  NAND2_X1 U4339 ( .A1(n3731), .A2(n3499), .ZN(n3497) );
  NAND2_X1 U4340 ( .A1(n3647), .A2(n4459), .ZN(n3496) );
  NAND2_X1 U4341 ( .A1(n3497), .A2(n3496), .ZN(n3498) );
  XNOR2_X1 U4342 ( .A(n3498), .B(n3754), .ZN(n3557) );
  NAND2_X1 U4343 ( .A1(n3735), .A2(n4459), .ZN(n3501) );
  NAND2_X1 U4344 ( .A1(n3647), .A2(n3499), .ZN(n3500) );
  INV_X1 U4345 ( .A(n3525), .ZN(n3556) );
  AOI22_X1 U4346 ( .A1(n3503), .A2(n3530), .B1(n3557), .B2(n3556), .ZN(n3511)
         );
  OAI21_X1 U4347 ( .B1(n3503), .B2(n3530), .A(n3557), .ZN(n3502) );
  NAND2_X1 U4348 ( .A1(n3502), .A2(n3525), .ZN(n3506) );
  INV_X1 U4349 ( .A(n3503), .ZN(n3527) );
  INV_X1 U4350 ( .A(n3557), .ZN(n3504) );
  NAND3_X1 U4351 ( .A1(n3527), .A2(n3528), .A3(n3504), .ZN(n3505) );
  OR2_X1 U4352 ( .A1(n3753), .A2(n3509), .ZN(n3507) );
  OAI21_X1 U4353 ( .B1(n3562), .B2(n3174), .A(n3507), .ZN(n3508) );
  XNOR2_X1 U4354 ( .A(n3508), .B(n3754), .ZN(n3513) );
  OAI22_X1 U4355 ( .A1(n3289), .A2(n3509), .B1(n3753), .B2(n3562), .ZN(n3512)
         );
  XNOR2_X1 U4356 ( .A(n3513), .B(n3512), .ZN(n3559) );
  OAI22_X1 U4357 ( .A1(n3576), .A2(n3174), .B1(n3781), .B2(n3753), .ZN(n3514)
         );
  XNOR2_X1 U4358 ( .A(n3514), .B(n3754), .ZN(n3516) );
  OAI22_X1 U4359 ( .A1(n3753), .A2(n3576), .B1(n3289), .B2(n3781), .ZN(n3515)
         );
  NOR2_X1 U4360 ( .A1(n3516), .A2(n3515), .ZN(n3593) );
  NOR2_X1 U4361 ( .A1(n3593), .A2(n2183), .ZN(n3517) );
  XNOR2_X1 U4362 ( .A(n3594), .B(n3517), .ZN(n3518) );
  NAND2_X1 U4363 ( .A1(n3518), .A2(n3920), .ZN(n3521) );
  NOR2_X1 U4364 ( .A1(n4850), .A2(STATE_REG_SCAN_IN), .ZN(n4122) );
  OAI22_X1 U4365 ( .A1(n3925), .A2(n3576), .B1(n4436), .B2(n3898), .ZN(n3519)
         );
  AOI211_X1 U4366 ( .C1(n3906), .C2(n4102), .A(n4122), .B(n3519), .ZN(n3520)
         );
  OAI211_X1 U4367 ( .C1(n3931), .C2(n3586), .A(n3521), .B(n3520), .ZN(U3233)
         );
  MUX2_X1 U4368 ( .A(n4838), .B(n3522), .S(n5043), .Z(n3523) );
  OAI21_X1 U4369 ( .B1(n4594), .B2(n3524), .A(n3523), .ZN(U3527) );
  XNOR2_X1 U4370 ( .A(n3525), .B(n3557), .ZN(n3532) );
  AOI21_X1 U4371 ( .B1(n3526), .B2(n3528), .A(n3527), .ZN(n3529) );
  AOI21_X1 U4372 ( .B1(n3392), .B2(n3530), .A(n3529), .ZN(n3531) );
  NAND2_X1 U4373 ( .A1(n3531), .A2(n3532), .ZN(n3555) );
  OAI21_X1 U4374 ( .B1(n3532), .B2(n3531), .A(n3555), .ZN(n3533) );
  NAND2_X1 U4375 ( .A1(n3533), .A2(n3920), .ZN(n3539) );
  OAI22_X1 U4376 ( .A1(n3925), .A2(n3535), .B1(n3534), .B2(n3923), .ZN(n3536)
         );
  AOI211_X1 U4377 ( .C1(n3927), .C2(n4102), .A(n3537), .B(n3536), .ZN(n3538)
         );
  OAI211_X1 U4378 ( .C1(n3931), .C2(n3540), .A(n3539), .B(n3538), .ZN(U3228)
         );
  INV_X1 U4379 ( .A(n3541), .ZN(n3542) );
  OR2_X1 U4380 ( .A1(n3574), .A2(n3542), .ZN(n3544) );
  NAND2_X1 U4381 ( .A1(n3544), .A2(n3543), .ZN(n4434) );
  AND2_X1 U4382 ( .A1(n4431), .A2(n4433), .ZN(n4039) );
  INV_X1 U4383 ( .A(n4039), .ZN(n3546) );
  XNOR2_X1 U4384 ( .A(n4434), .B(n3546), .ZN(n3545) );
  NAND2_X1 U4385 ( .A1(n3545), .A2(n4595), .ZN(n4592) );
  XNOR2_X1 U4386 ( .A(n3547), .B(n3546), .ZN(n4590) );
  AOI22_X1 U4387 ( .A1(n4476), .A2(n4586), .B1(n4474), .B2(n4585), .ZN(n3550)
         );
  INV_X1 U4388 ( .A(n3548), .ZN(n3783) );
  AOI22_X1 U4389 ( .A1(n4454), .A2(REG2_REG_12__SCAN_IN), .B1(n3783), .B2(
        n4481), .ZN(n3549) );
  OAI211_X1 U4390 ( .C1(n3596), .C2(n4424), .A(n3550), .B(n3549), .ZN(n3553)
         );
  INV_X1 U4391 ( .A(n4446), .ZN(n3551) );
  OAI21_X1 U4392 ( .B1(n3568), .B2(n3596), .A(n3551), .ZN(n4937) );
  NOR2_X1 U4393 ( .A1(n4937), .A2(n4449), .ZN(n3552) );
  AOI211_X1 U4394 ( .C1(n4467), .C2(n4590), .A(n3553), .B(n3552), .ZN(n3554)
         );
  OAI21_X1 U4395 ( .B1(n4592), .B2(n4454), .A(n3554), .ZN(U3278) );
  OAI21_X1 U4396 ( .B1(n3557), .B2(n3556), .A(n3555), .ZN(n3560) );
  AOI211_X1 U4397 ( .C1(n3560), .C2(n3559), .A(n3558), .B(n3913), .ZN(n3561)
         );
  INV_X1 U4398 ( .A(n3561), .ZN(n3566) );
  OAI22_X1 U4399 ( .A1(n3925), .A2(n3562), .B1(n3781), .B2(n3898), .ZN(n3563)
         );
  AOI211_X1 U4400 ( .C1(n3906), .C2(n4459), .A(n3564), .B(n3563), .ZN(n3565)
         );
  OAI211_X1 U4401 ( .C1(n3931), .C2(n3567), .A(n3566), .B(n3565), .ZN(U3214)
         );
  INV_X1 U4402 ( .A(n3568), .ZN(n3569) );
  OAI21_X1 U4403 ( .B1(n3570), .B2(n3576), .A(n3569), .ZN(n3587) );
  INV_X1 U4404 ( .A(n3571), .ZN(n5037) );
  OAI21_X1 U4405 ( .B1(n3573), .B2(n4024), .A(n3572), .ZN(n3591) );
  XNOR2_X1 U4406 ( .A(n3574), .B(n4024), .ZN(n3580) );
  AOI22_X1 U4407 ( .A1(n4102), .A2(n4584), .B1(n4601), .B2(n4101), .ZN(n3575)
         );
  OAI21_X1 U4408 ( .B1(n3576), .B2(n4572), .A(n3575), .ZN(n3577) );
  AOI21_X1 U4409 ( .B1(n3591), .B2(n3578), .A(n3577), .ZN(n3579) );
  OAI21_X1 U4410 ( .B1(n3580), .B2(n4441), .A(n3579), .ZN(n3588) );
  AOI21_X1 U4411 ( .B1(n5037), .B2(n3591), .A(n3588), .ZN(n3583) );
  MUX2_X1 U4412 ( .A(n3581), .B(n3583), .S(n5040), .Z(n3582) );
  OAI21_X1 U4413 ( .B1(n3587), .B2(n4936), .A(n3582), .ZN(U3489) );
  MUX2_X1 U4414 ( .A(n3584), .B(n3583), .S(n5043), .Z(n3585) );
  OAI21_X1 U4415 ( .B1(n4594), .B2(n3587), .A(n3585), .ZN(U3529) );
  OAI22_X1 U4416 ( .A1(n3587), .A2(n4449), .B1(n3586), .B2(n4461), .ZN(n3590)
         );
  MUX2_X1 U4417 ( .A(n3588), .B(REG2_REG_11__SCAN_IN), .S(n4386), .Z(n3589) );
  AOI211_X1 U4418 ( .C1(n4483), .C2(n3591), .A(n3590), .B(n3589), .ZN(n3592)
         );
  INV_X1 U4419 ( .A(n3592), .ZN(U3279) );
  OAI22_X1 U4420 ( .A1(n3596), .A2(n3174), .B1(n4436), .B2(n3753), .ZN(n3595)
         );
  XNOR2_X1 U4421 ( .A(n3595), .B(n3754), .ZN(n3597) );
  INV_X1 U4422 ( .A(n3597), .ZN(n3778) );
  OAI22_X1 U4423 ( .A1(n3596), .A2(n3753), .B1(n4436), .B2(n3289), .ZN(n3777)
         );
  AOI22_X1 U4424 ( .A1(n3735), .A2(n4586), .B1(n4439), .B2(n3232), .ZN(n3602)
         );
  NAND2_X1 U4425 ( .A1(n3731), .A2(n4439), .ZN(n3599) );
  NAND2_X1 U4426 ( .A1(n3647), .A2(n4586), .ZN(n3598) );
  NAND2_X1 U4427 ( .A1(n3599), .A2(n3598), .ZN(n3600) );
  XNOR2_X1 U4428 ( .A(n3600), .B(n3658), .ZN(n3601) );
  INV_X1 U4429 ( .A(n3601), .ZN(n3604) );
  INV_X1 U4430 ( .A(n3602), .ZN(n3603) );
  NAND2_X1 U4431 ( .A1(n2182), .A2(n3641), .ZN(n3605) );
  XNOR2_X1 U4432 ( .A(n3642), .B(n3605), .ZN(n3606) );
  NAND2_X1 U4433 ( .A1(n3606), .A2(n3920), .ZN(n3610) );
  NOR2_X1 U4434 ( .A1(n3607), .A2(STATE_REG_SCAN_IN), .ZN(n4147) );
  OAI22_X1 U4435 ( .A1(n3925), .A2(n4445), .B1(n4437), .B2(n3898), .ZN(n3608)
         );
  AOI211_X1 U4436 ( .C1(n3906), .C2(n4101), .A(n4147), .B(n3608), .ZN(n3609)
         );
  OAI211_X1 U4437 ( .C1(n3931), .C2(n4450), .A(n3610), .B(n3609), .ZN(U3231)
         );
  NAND2_X1 U4438 ( .A1(n4414), .A2(n3979), .ZN(n3611) );
  XNOR2_X1 U4439 ( .A(n3611), .B(n4018), .ZN(n3612) );
  NOR2_X1 U4440 ( .A1(n3612), .A2(n4441), .ZN(n4566) );
  INV_X1 U4441 ( .A(n4566), .ZN(n3621) );
  NAND2_X1 U4442 ( .A1(n4412), .A2(n4416), .ZN(n4411) );
  NAND2_X1 U4443 ( .A1(n4411), .A2(n3613), .ZN(n4395) );
  XNOR2_X1 U4444 ( .A(n4395), .B(n4018), .ZN(n4568) );
  INV_X1 U4445 ( .A(n3614), .ZN(n4404) );
  OAI21_X1 U4446 ( .B1(n2424), .B2(n3924), .A(n4404), .ZN(n4924) );
  INV_X1 U4447 ( .A(REG2_REG_15__SCAN_IN), .ZN(n3615) );
  OAI22_X1 U4448 ( .A1(n4484), .A2(n3615), .B1(n3930), .B2(n4461), .ZN(n3617)
         );
  OAI22_X1 U4449 ( .A1(n4293), .A2(n4437), .B1(n4565), .B2(n4295), .ZN(n3616)
         );
  AOI211_X1 U4450 ( .C1(n4561), .C2(n4478), .A(n3617), .B(n3616), .ZN(n3618)
         );
  OAI21_X1 U4451 ( .B1(n4924), .B2(n4449), .A(n3618), .ZN(n3619) );
  AOI21_X1 U4452 ( .B1(n4568), .B2(n4467), .A(n3619), .ZN(n3620) );
  OAI21_X1 U4453 ( .B1(n3621), .B2(n4454), .A(n3620), .ZN(U3275) );
  AOI22_X1 U4454 ( .A1(n4478), .A2(n3761), .B1(n4454), .B2(
        REG2_REG_28__SCAN_IN), .ZN(n3623) );
  NAND2_X1 U4455 ( .A1(n3762), .A2(n4481), .ZN(n3622) );
  OAI211_X1 U4456 ( .C1(n3765), .C2(n4295), .A(n3623), .B(n3622), .ZN(n3624)
         );
  AOI21_X1 U4457 ( .B1(n4474), .B2(n4203), .A(n3624), .ZN(n3625) );
  OAI21_X1 U4458 ( .B1(n3626), .B2(n4449), .A(n3625), .ZN(n3627) );
  AOI21_X1 U4459 ( .B1(n3628), .B2(n4484), .A(n3627), .ZN(n3629) );
  OAI21_X1 U4460 ( .B1(n3630), .B2(n4304), .A(n3629), .ZN(U3262) );
  AND2_X1 U4461 ( .A1(n2335), .A2(DATAI_29_), .ZN(n3932) );
  NAND2_X1 U4462 ( .A1(n2335), .A2(DATAI_30_), .ZN(n4164) );
  AND2_X1 U4463 ( .A1(n4950), .A2(B_REG_SCAN_IN), .ZN(n3631) );
  NOR2_X1 U4464 ( .A1(n4564), .A2(n3631), .ZN(n3790) );
  NAND2_X1 U4465 ( .A1(n3790), .A2(n4004), .ZN(n4167) );
  OAI21_X1 U4466 ( .B1(n4078), .B2(n4572), .A(n4167), .ZN(n3638) );
  NAND2_X1 U4467 ( .A1(n4484), .A2(n3638), .ZN(n3633) );
  NAND2_X1 U4468 ( .A1(n4454), .A2(REG2_REG_31__SCAN_IN), .ZN(n3632) );
  OAI211_X1 U4469 ( .C1(n3640), .C2(n4449), .A(n3633), .B(n3632), .ZN(U3260)
         );
  NAND2_X1 U4470 ( .A1(n5043), .A2(n3638), .ZN(n3635) );
  NAND2_X1 U4471 ( .A1(n2210), .A2(REG1_REG_31__SCAN_IN), .ZN(n3634) );
  OAI211_X1 U4472 ( .C1(n3640), .C2(n4594), .A(n3635), .B(n3634), .ZN(U3549)
         );
  NOR2_X1 U4473 ( .A1(n5040), .A2(n3636), .ZN(n3637) );
  AOI21_X1 U4474 ( .B1(n5040), .B2(n3638), .A(n3637), .ZN(n3639) );
  OAI21_X1 U4475 ( .B1(n3640), .B2(n4936), .A(n3639), .ZN(U3517) );
  OAI22_X1 U4476 ( .A1(n4437), .A2(n3753), .B1(n4573), .B2(n3174), .ZN(n3643)
         );
  XOR2_X1 U4477 ( .A(n3754), .B(n3643), .Z(n3644) );
  OAI22_X1 U4478 ( .A1(n4437), .A2(n3289), .B1(n4573), .B2(n3753), .ZN(n3802)
         );
  INV_X1 U4479 ( .A(n3805), .ZN(n3645) );
  INV_X1 U4480 ( .A(n3644), .ZN(n3803) );
  AOI22_X1 U4481 ( .A1(n3646), .A2(n3802), .B1(n3645), .B2(n3803), .ZN(n3840)
         );
  INV_X1 U4482 ( .A(n3840), .ZN(n3667) );
  NAND2_X1 U4483 ( .A1(n4570), .A2(n3647), .ZN(n3649) );
  NAND2_X1 U4484 ( .A1(n3731), .A2(n4561), .ZN(n3648) );
  NAND2_X1 U4485 ( .A1(n3649), .A2(n3648), .ZN(n3650) );
  XNOR2_X1 U4486 ( .A(n3650), .B(n3658), .ZN(n3841) );
  INV_X1 U4487 ( .A(n3841), .ZN(n3654) );
  NAND2_X1 U4488 ( .A1(n4570), .A2(n3735), .ZN(n3652) );
  NAND2_X1 U4489 ( .A1(n3232), .A2(n4561), .ZN(n3651) );
  OAI22_X1 U4490 ( .A1(n4565), .A2(n3753), .B1(n3174), .B2(n3656), .ZN(n3655)
         );
  XNOR2_X1 U4491 ( .A(n3655), .B(n3754), .ZN(n3843) );
  OAI22_X1 U4492 ( .A1(n4565), .A2(n3289), .B1(n3753), .B2(n3656), .ZN(n3661)
         );
  NAND2_X1 U4493 ( .A1(n3843), .A2(n3661), .ZN(n3663) );
  OAI22_X1 U4494 ( .A1(n4391), .A2(n3753), .B1(n4546), .B2(n3174), .ZN(n3659)
         );
  XNOR2_X1 U4495 ( .A(n3659), .B(n3658), .ZN(n3852) );
  NOR2_X1 U4496 ( .A1(n4546), .A2(n3753), .ZN(n3660) );
  AOI21_X1 U4497 ( .B1(n4350), .B2(n3735), .A(n3660), .ZN(n3853) );
  NAND2_X1 U4498 ( .A1(n3852), .A2(n3853), .ZN(n3665) );
  INV_X1 U4499 ( .A(n3843), .ZN(n3662) );
  INV_X1 U4500 ( .A(n3661), .ZN(n3842) );
  NAND2_X1 U4501 ( .A1(n3662), .A2(n3842), .ZN(n3850) );
  NAND3_X1 U4502 ( .A1(n3663), .A2(n3918), .A3(n3841), .ZN(n3664) );
  INV_X1 U4503 ( .A(n3852), .ZN(n3669) );
  OAI22_X1 U4504 ( .A1(n4334), .A2(n3753), .B1(n3174), .B2(n4360), .ZN(n3672)
         );
  XNOR2_X1 U4505 ( .A(n3672), .B(n3754), .ZN(n3673) );
  OAI22_X1 U4506 ( .A1(n4334), .A2(n3289), .B1(n3753), .B2(n4360), .ZN(n3674)
         );
  AND2_X1 U4507 ( .A1(n3673), .A2(n3674), .ZN(n3893) );
  INV_X1 U4508 ( .A(n3673), .ZN(n3676) );
  INV_X1 U4509 ( .A(n3674), .ZN(n3675) );
  NAND2_X1 U4510 ( .A1(n3676), .A2(n3675), .ZN(n3894) );
  OAI22_X1 U4511 ( .A1(n4352), .A2(n3289), .B1(n3753), .B2(n4341), .ZN(n3679)
         );
  OAI22_X1 U4512 ( .A1(n4352), .A2(n3753), .B1(n3174), .B2(n4341), .ZN(n3677)
         );
  XNOR2_X1 U4513 ( .A(n3677), .B(n3754), .ZN(n3678) );
  XOR2_X1 U4514 ( .A(n3679), .B(n3678), .Z(n3826) );
  NAND2_X1 U4515 ( .A1(n4525), .A2(n3232), .ZN(n3683) );
  NAND2_X1 U4516 ( .A1(n3731), .A2(n4310), .ZN(n3682) );
  NAND2_X1 U4517 ( .A1(n3683), .A2(n3682), .ZN(n3684) );
  XNOR2_X1 U4518 ( .A(n3684), .B(n3754), .ZN(n3687) );
  NAND2_X1 U4519 ( .A1(n4525), .A2(n3735), .ZN(n3686) );
  NAND2_X1 U4520 ( .A1(n3647), .A2(n4310), .ZN(n3685) );
  NAND2_X1 U4521 ( .A1(n3686), .A2(n3685), .ZN(n3688) );
  NAND2_X1 U4522 ( .A1(n3687), .A2(n3688), .ZN(n3871) );
  INV_X1 U4523 ( .A(n3687), .ZN(n3690) );
  INV_X1 U4524 ( .A(n3688), .ZN(n3689) );
  NAND2_X1 U4525 ( .A1(n3690), .A2(n3689), .ZN(n3873) );
  NAND2_X1 U4526 ( .A1(n4269), .A2(n3647), .ZN(n3692) );
  NAND2_X1 U4527 ( .A1(n3731), .A2(n4524), .ZN(n3691) );
  NAND2_X1 U4528 ( .A1(n3692), .A2(n3691), .ZN(n3693) );
  XNOR2_X1 U4529 ( .A(n3693), .B(n3754), .ZN(n3833) );
  NAND2_X1 U4530 ( .A1(n4269), .A2(n3735), .ZN(n3695) );
  NAND2_X1 U4531 ( .A1(n3647), .A2(n4524), .ZN(n3694) );
  NAND2_X1 U4532 ( .A1(n3695), .A2(n3694), .ZN(n3832) );
  NOR2_X1 U4533 ( .A1(n3833), .A2(n3832), .ZN(n3814) );
  OAI22_X1 U4534 ( .A1(n4272), .A2(n3753), .B1(n4258), .B2(n3174), .ZN(n3696)
         );
  XNOR2_X1 U4535 ( .A(n3696), .B(n3754), .ZN(n3703) );
  OAI22_X1 U4536 ( .A1(n4272), .A2(n3289), .B1(n4258), .B2(n3753), .ZN(n3702)
         );
  XNOR2_X1 U4537 ( .A(n3703), .B(n3702), .ZN(n3816) );
  OAI22_X1 U4538 ( .A1(n4527), .A2(n3753), .B1(n4273), .B2(n3174), .ZN(n3697)
         );
  XNOR2_X1 U4539 ( .A(n3697), .B(n3754), .ZN(n3699) );
  OAI22_X1 U4540 ( .A1(n4527), .A2(n3289), .B1(n4273), .B2(n3753), .ZN(n3698)
         );
  NOR2_X1 U4541 ( .A1(n3699), .A2(n3698), .ZN(n3817) );
  XNOR2_X1 U4542 ( .A(n3699), .B(n3698), .ZN(n3884) );
  INV_X1 U4543 ( .A(n3884), .ZN(n3700) );
  NAND2_X1 U4544 ( .A1(n3833), .A2(n3832), .ZN(n3880) );
  AND2_X1 U4545 ( .A1(n3700), .A2(n3880), .ZN(n3815) );
  NAND2_X1 U4546 ( .A1(n3703), .A2(n3702), .ZN(n3707) );
  NOR2_X1 U4547 ( .A1(n3753), .A2(n4235), .ZN(n3704) );
  AOI21_X1 U4548 ( .B1(n4504), .B2(n3735), .A(n3704), .ZN(n3708) );
  OAI22_X1 U4549 ( .A1(n3820), .A2(n3753), .B1(n4235), .B2(n3174), .ZN(n3706)
         );
  XNOR2_X1 U4550 ( .A(n3706), .B(n3754), .ZN(n3863) );
  NAND2_X1 U4551 ( .A1(n3861), .A2(n3863), .ZN(n3711) );
  INV_X1 U4552 ( .A(n3708), .ZN(n3709) );
  NAND2_X1 U4553 ( .A1(n3710), .A2(n3709), .ZN(n3860) );
  NAND2_X1 U4554 ( .A1(n3711), .A2(n3860), .ZN(n3730) );
  OAI22_X1 U4555 ( .A1(n4201), .A2(n3753), .B1(n3174), .B2(n4222), .ZN(n3712)
         );
  XNOR2_X1 U4556 ( .A(n3712), .B(n3754), .ZN(n3714) );
  OAI22_X1 U4557 ( .A1(n4201), .A2(n3289), .B1(n3753), .B2(n4222), .ZN(n3713)
         );
  OR2_X1 U4558 ( .A1(n3714), .A2(n3713), .ZN(n3729) );
  AND2_X1 U4559 ( .A1(n3714), .A2(n3713), .ZN(n3728) );
  NOR2_X1 U4560 ( .A1(n2411), .A2(n3728), .ZN(n3715) );
  XNOR2_X1 U4561 ( .A(n3730), .B(n3715), .ZN(n3720) );
  AOI22_X1 U4562 ( .A1(n4504), .A2(n3906), .B1(REG3_REG_25__SCAN_IN), .B2(
        U3149), .ZN(n3717) );
  NAND2_X1 U4563 ( .A1(n3908), .A2(n4503), .ZN(n3716) );
  OAI211_X1 U4564 ( .C1(n4506), .C2(n3898), .A(n3717), .B(n3716), .ZN(n3718)
         );
  AOI21_X1 U4565 ( .B1(n4220), .B2(n3889), .A(n3718), .ZN(n3719) );
  OAI21_X1 U4566 ( .B1(n3720), .B2(n3913), .A(n3719), .ZN(U3222) );
  AOI21_X1 U4567 ( .B1(n4600), .B2(n3721), .A(n4478), .ZN(n3727) );
  NAND2_X1 U4568 ( .A1(n3726), .A2(n4473), .ZN(n3943) );
  NAND2_X1 U4569 ( .A1(n3943), .A2(n3941), .ZN(n4598) );
  OAI21_X1 U4570 ( .B1(n4456), .B2(n4467), .A(n4598), .ZN(n3725) );
  OAI22_X1 U4571 ( .A1(n4484), .A2(n4617), .B1(n3722), .B2(n4461), .ZN(n3723)
         );
  AOI21_X1 U4572 ( .B1(n4476), .B2(n4602), .A(n3723), .ZN(n3724) );
  OAI211_X1 U4573 ( .C1(n3727), .C2(n3726), .A(n3725), .B(n3724), .ZN(U3290)
         );
  NAND2_X1 U4574 ( .A1(n4493), .A2(n3647), .ZN(n3733) );
  NAND2_X1 U4575 ( .A1(n3731), .A2(n3907), .ZN(n3732) );
  NAND2_X1 U4576 ( .A1(n3733), .A2(n3732), .ZN(n3734) );
  XNOR2_X1 U4577 ( .A(n3734), .B(n3754), .ZN(n3738) );
  NAND2_X1 U4578 ( .A1(n4493), .A2(n3735), .ZN(n3737) );
  NAND2_X1 U4579 ( .A1(n3232), .A2(n3907), .ZN(n3736) );
  NAND2_X1 U4580 ( .A1(n3737), .A2(n3736), .ZN(n3739) );
  NAND2_X1 U4581 ( .A1(n3738), .A2(n3739), .ZN(n3903) );
  INV_X1 U4582 ( .A(n3738), .ZN(n3741) );
  INV_X1 U4583 ( .A(n3739), .ZN(n3740) );
  NAND2_X1 U4584 ( .A1(n3741), .A2(n3740), .ZN(n3904) );
  OAI22_X1 U4585 ( .A1(n3997), .A2(n3753), .B1(n4185), .B2(n3174), .ZN(n3742)
         );
  XNOR2_X1 U4586 ( .A(n3742), .B(n3754), .ZN(n3759) );
  OAI22_X1 U4587 ( .A1(n3997), .A2(n3289), .B1(n4185), .B2(n3753), .ZN(n3758)
         );
  XNOR2_X1 U4588 ( .A(n3759), .B(n3758), .ZN(n3751) );
  XNOR2_X1 U4589 ( .A(n3752), .B(n3751), .ZN(n3750) );
  INV_X1 U4590 ( .A(n4185), .ZN(n4492) );
  NAND2_X1 U4591 ( .A1(n3908), .A2(n4492), .ZN(n3743) );
  OAI21_X1 U4592 ( .B1(STATE_REG_SCAN_IN), .B2(n3744), .A(n3743), .ZN(n3745)
         );
  AOI21_X1 U4593 ( .B1(n4493), .B2(n3906), .A(n3745), .ZN(n3747) );
  NAND2_X1 U4594 ( .A1(n4187), .A2(n3889), .ZN(n3746) );
  OAI211_X1 U4595 ( .C1(n4495), .C2(n3898), .A(n3747), .B(n3746), .ZN(n3748)
         );
  INV_X1 U4596 ( .A(n3748), .ZN(n3749) );
  OAI21_X1 U4597 ( .B1(n3750), .B2(n3913), .A(n3749), .ZN(U3211) );
  OAI22_X1 U4598 ( .A1(n4495), .A2(n3289), .B1(n3753), .B2(n3786), .ZN(n3755)
         );
  XNOR2_X1 U4599 ( .A(n3755), .B(n3754), .ZN(n3757) );
  OAI22_X1 U4600 ( .A1(n4495), .A2(n3753), .B1(n3174), .B2(n3786), .ZN(n3756)
         );
  XNOR2_X1 U4601 ( .A(n3757), .B(n3756), .ZN(n3766) );
  NAND2_X1 U4602 ( .A1(n3766), .A2(n3920), .ZN(n3774) );
  AND2_X1 U4603 ( .A1(n3759), .A2(n3758), .ZN(n3767) );
  NOR3_X1 U4604 ( .A1(n3766), .A2(n3767), .A3(n3913), .ZN(n3760) );
  NAND2_X1 U4605 ( .A1(n3775), .A2(n3760), .ZN(n3773) );
  AOI22_X1 U4606 ( .A1(n3908), .A2(n3761), .B1(REG3_REG_28__SCAN_IN), .B2(
        U3149), .ZN(n3764) );
  NAND2_X1 U4607 ( .A1(n3762), .A2(n3889), .ZN(n3763) );
  OAI211_X1 U4608 ( .C1(n3765), .C2(n3898), .A(n3764), .B(n3763), .ZN(n3771)
         );
  INV_X1 U4609 ( .A(n3766), .ZN(n3769) );
  INV_X1 U4610 ( .A(n3767), .ZN(n3768) );
  NOR3_X1 U4611 ( .A1(n3769), .A2(n3913), .A3(n3768), .ZN(n3770) );
  AOI211_X1 U4612 ( .C1(n3906), .C2(n4203), .A(n3771), .B(n3770), .ZN(n3772)
         );
  OAI211_X1 U4613 ( .C1(n3775), .C2(n3774), .A(n3773), .B(n3772), .ZN(U3217)
         );
  XNOR2_X1 U4614 ( .A(n3778), .B(n3777), .ZN(n3779) );
  XNOR2_X1 U4615 ( .A(n3776), .B(n3779), .ZN(n3785) );
  AOI22_X1 U4616 ( .A1(n4583), .A2(n3908), .B1(n3927), .B2(n4586), .ZN(n3780)
         );
  NAND2_X1 U4617 ( .A1(U3149), .A2(REG3_REG_12__SCAN_IN), .ZN(n4132) );
  OAI211_X1 U4618 ( .C1(n3781), .C2(n3923), .A(n3780), .B(n4132), .ZN(n3782)
         );
  AOI21_X1 U4619 ( .B1(n3783), .B2(n3889), .A(n3782), .ZN(n3784) );
  OAI21_X1 U4620 ( .B1(n3785), .B2(n3913), .A(n3784), .ZN(U3221) );
  INV_X1 U4621 ( .A(REG1_REG_29__SCAN_IN), .ZN(n3794) );
  XNOR2_X1 U4622 ( .A(n4097), .B(n3932), .ZN(n4048) );
  XNOR2_X1 U4623 ( .A(n3788), .B(n4048), .ZN(n4170) );
  INV_X1 U4624 ( .A(n4048), .ZN(n3789) );
  AOI22_X1 U4625 ( .A1(n3790), .A2(n4005), .B1(n3932), .B2(n4582), .ZN(n3792)
         );
  NAND2_X1 U4626 ( .A1(n4098), .A2(n4584), .ZN(n3791) );
  AOI21_X1 U4627 ( .B1(n4170), .B2(n4596), .A(n4175), .ZN(n3798) );
  MUX2_X1 U4628 ( .A(n3794), .B(n3798), .S(n5043), .Z(n3797) );
  AOI21_X1 U4629 ( .B1(n3932), .B2(n3795), .A(n4162), .ZN(n4171) );
  NAND2_X1 U4630 ( .A1(n4171), .A2(n4559), .ZN(n3796) );
  NAND2_X1 U4631 ( .A1(n3797), .A2(n3796), .ZN(U3547) );
  INV_X1 U4632 ( .A(REG0_REG_29__SCAN_IN), .ZN(n3799) );
  MUX2_X1 U4633 ( .A(n3799), .B(n3798), .S(n5040), .Z(n3801) );
  NAND2_X1 U4634 ( .A1(n4171), .A2(n4918), .ZN(n3800) );
  NAND2_X1 U4635 ( .A1(n3801), .A2(n3800), .ZN(U3515) );
  XNOR2_X1 U4636 ( .A(n3803), .B(n3802), .ZN(n3804) );
  XNOR2_X1 U4637 ( .A(n3805), .B(n3804), .ZN(n3812) );
  INV_X1 U4638 ( .A(n3806), .ZN(n4421) );
  INV_X1 U4639 ( .A(n4586), .ZN(n3809) );
  AOI22_X1 U4640 ( .A1(n3807), .A2(n3908), .B1(n3927), .B2(n4570), .ZN(n3808)
         );
  NAND2_X1 U4641 ( .A1(U3149), .A2(REG3_REG_14__SCAN_IN), .ZN(n4152) );
  OAI211_X1 U4642 ( .C1(n3809), .C2(n3923), .A(n3808), .B(n4152), .ZN(n3810)
         );
  AOI21_X1 U4643 ( .B1(n4421), .B2(n3889), .A(n3810), .ZN(n3811) );
  OAI21_X1 U4644 ( .B1(n3812), .B2(n3913), .A(n3811), .ZN(U3212) );
  OR2_X1 U4645 ( .A1(n3813), .A2(n3814), .ZN(n3881) );
  AND2_X1 U4646 ( .A1(n3881), .A2(n3815), .ZN(n3882) );
  OAI21_X1 U4647 ( .B1(n3882), .B2(n3817), .A(n3816), .ZN(n3819) );
  NAND3_X1 U4648 ( .A1(n3819), .A2(n3920), .A3(n3818), .ZN(n3824) );
  OAI22_X1 U4649 ( .A1(n4527), .A2(n3923), .B1(STATE_REG_SCAN_IN), .B2(n4668), 
        .ZN(n3822) );
  OAI22_X1 U4650 ( .A1(n3820), .A2(n3898), .B1(n3925), .B2(n4258), .ZN(n3821)
         );
  AOI211_X1 U4651 ( .C1(n4259), .C2(n3889), .A(n3822), .B(n3821), .ZN(n3823)
         );
  NAND2_X1 U4652 ( .A1(n3824), .A2(n3823), .ZN(U3213) );
  XOR2_X1 U4653 ( .A(n3826), .B(n3825), .Z(n3831) );
  AOI22_X1 U4654 ( .A1(n4040), .A2(n3908), .B1(n3906), .B2(n4549), .ZN(n3828)
         );
  OAI211_X1 U4655 ( .C1(n4294), .C2(n3898), .A(n3828), .B(n3827), .ZN(n3829)
         );
  AOI21_X1 U4656 ( .B1(n4343), .B2(n3889), .A(n3829), .ZN(n3830) );
  OAI21_X1 U4657 ( .B1(n3831), .B2(n3913), .A(n3830), .ZN(U3216) );
  XNOR2_X1 U4658 ( .A(n3833), .B(n3832), .ZN(n3834) );
  XNOR2_X1 U4659 ( .A(n3813), .B(n3834), .ZN(n3839) );
  OAI22_X1 U4660 ( .A1(n4294), .A2(n3923), .B1(n3925), .B2(n4300), .ZN(n3837)
         );
  OAI22_X1 U4661 ( .A1(n4527), .A2(n3898), .B1(STATE_REG_SCAN_IN), .B2(n3835), 
        .ZN(n3836) );
  AOI211_X1 U4662 ( .C1(n4297), .C2(n3889), .A(n3837), .B(n3836), .ZN(n3838)
         );
  OAI21_X1 U4663 ( .B1(n3839), .B2(n3913), .A(n3838), .ZN(U3220) );
  AOI21_X1 U4664 ( .B1(n3918), .B2(n3915), .A(n3916), .ZN(n3844) );
  XNOR2_X1 U4665 ( .A(n3843), .B(n3842), .ZN(n3849) );
  XNOR2_X1 U4666 ( .A(n3844), .B(n3849), .ZN(n3848) );
  AOI22_X1 U4667 ( .A1(n4405), .A2(n3908), .B1(n3906), .B2(n4570), .ZN(n3845)
         );
  NAND2_X1 U4668 ( .A1(U3149), .A2(REG3_REG_16__SCAN_IN), .ZN(n4975) );
  OAI211_X1 U4669 ( .C1(n4391), .C2(n3898), .A(n3845), .B(n4975), .ZN(n3846)
         );
  AOI21_X1 U4670 ( .B1(n4406), .B2(n3889), .A(n3846), .ZN(n3847) );
  OAI21_X1 U4671 ( .B1(n3848), .B2(n3913), .A(n3847), .ZN(U3223) );
  OAI211_X1 U4672 ( .C1(n3916), .C2(n3918), .A(n3849), .B(n3915), .ZN(n3851)
         );
  NAND2_X1 U4673 ( .A1(n3851), .A2(n3850), .ZN(n3855) );
  XOR2_X1 U4674 ( .A(n3853), .B(n3852), .Z(n3854) );
  XNOR2_X1 U4675 ( .A(n3855), .B(n3854), .ZN(n3856) );
  NAND2_X1 U4676 ( .A1(n3856), .A2(n3920), .ZN(n3859) );
  AND2_X1 U4677 ( .A1(U3149), .A2(REG3_REG_17__SCAN_IN), .ZN(n4983) );
  OAI22_X1 U4678 ( .A1(n3925), .A2(n4546), .B1(n4334), .B2(n3898), .ZN(n3857)
         );
  AOI211_X1 U4679 ( .C1(n3906), .C2(n4381), .A(n4983), .B(n3857), .ZN(n3858)
         );
  OAI211_X1 U4680 ( .C1(n3931), .C2(n4377), .A(n3859), .B(n3858), .ZN(U3225)
         );
  NAND2_X1 U4681 ( .A1(n3860), .A2(n3861), .ZN(n3862) );
  XOR2_X1 U4682 ( .A(n3863), .B(n3862), .Z(n3868) );
  OAI22_X1 U4683 ( .A1(n4272), .A2(n3923), .B1(STATE_REG_SCAN_IN), .B2(n4822), 
        .ZN(n3864) );
  AOI21_X1 U4684 ( .B1(n4240), .B2(n3908), .A(n3864), .ZN(n3865) );
  OAI21_X1 U4685 ( .B1(n4201), .B2(n3898), .A(n3865), .ZN(n3866) );
  AOI21_X1 U4686 ( .B1(n4243), .B2(n3889), .A(n3866), .ZN(n3867) );
  OAI21_X1 U4687 ( .B1(n3868), .B2(n3913), .A(n3867), .ZN(U3226) );
  INV_X1 U4688 ( .A(n3869), .ZN(n3874) );
  AOI21_X1 U4689 ( .B1(n3873), .B2(n3871), .A(n3870), .ZN(n3872) );
  AOI21_X1 U4690 ( .B1(n3874), .B2(n3873), .A(n3872), .ZN(n3879) );
  INV_X1 U4691 ( .A(n3875), .ZN(n4322) );
  OAI22_X1 U4692 ( .A1(n3925), .A2(n4320), .B1(n4352), .B2(n3923), .ZN(n3877)
         );
  OAI22_X1 U4693 ( .A1(n4313), .A2(n3898), .B1(STATE_REG_SCAN_IN), .B2(n2297), 
        .ZN(n3876) );
  AOI211_X1 U4694 ( .C1(n4322), .C2(n3889), .A(n3877), .B(n3876), .ZN(n3878)
         );
  OAI21_X1 U4695 ( .B1(n3879), .B2(n3913), .A(n3878), .ZN(U3230) );
  NAND2_X1 U4696 ( .A1(n3881), .A2(n3880), .ZN(n3883) );
  AOI21_X1 U4697 ( .B1(n3884), .B2(n3883), .A(n3882), .ZN(n3891) );
  INV_X1 U4698 ( .A(n3885), .ZN(n4276) );
  OAI22_X1 U4699 ( .A1(n4313), .A2(n3923), .B1(n3925), .B2(n4273), .ZN(n3888)
         );
  OAI22_X1 U4700 ( .A1(n4272), .A2(n3898), .B1(STATE_REG_SCAN_IN), .B2(n3886), 
        .ZN(n3887) );
  AOI211_X1 U4701 ( .C1(n4276), .C2(n3889), .A(n3888), .B(n3887), .ZN(n3890)
         );
  OAI21_X1 U4702 ( .B1(n3891), .B2(n3913), .A(n3890), .ZN(U3232) );
  INV_X1 U4703 ( .A(n3893), .ZN(n3895) );
  NAND2_X1 U4704 ( .A1(n3895), .A2(n3894), .ZN(n3896) );
  XNOR2_X1 U4705 ( .A(n3892), .B(n3896), .ZN(n3897) );
  NAND2_X1 U4706 ( .A1(n3897), .A2(n3920), .ZN(n3901) );
  NOR2_X1 U4707 ( .A1(n2296), .A2(STATE_REG_SCAN_IN), .ZN(n4993) );
  OAI22_X1 U4708 ( .A1(n3925), .A2(n4360), .B1(n4352), .B2(n3898), .ZN(n3899)
         );
  AOI211_X1 U4709 ( .C1(n3906), .C2(n4350), .A(n4993), .B(n3899), .ZN(n3900)
         );
  OAI211_X1 U4710 ( .C1(n3931), .C2(n4363), .A(n3901), .B(n3900), .ZN(U3235)
         );
  NAND2_X1 U4711 ( .A1(n3904), .A2(n3903), .ZN(n3905) );
  XNOR2_X1 U4712 ( .A(n3902), .B(n3905), .ZN(n3914) );
  NAND2_X1 U4713 ( .A1(n4237), .A2(n3906), .ZN(n3910) );
  AOI22_X1 U4714 ( .A1(n3908), .A2(n3907), .B1(REG3_REG_26__SCAN_IN), .B2(
        U3149), .ZN(n3909) );
  OAI211_X1 U4715 ( .C1(n3931), .C2(n4209), .A(n3910), .B(n3909), .ZN(n3911)
         );
  AOI21_X1 U4716 ( .B1(n3927), .B2(n4203), .A(n3911), .ZN(n3912) );
  OAI21_X1 U4717 ( .B1(n3914), .B2(n3913), .A(n3912), .ZN(U3237) );
  INV_X1 U4718 ( .A(n3915), .ZN(n3917) );
  NOR2_X1 U4719 ( .A1(n3917), .A2(n3916), .ZN(n3919) );
  XNOR2_X1 U4720 ( .A(n3919), .B(n3918), .ZN(n3921) );
  NAND2_X1 U4721 ( .A1(n3921), .A2(n3920), .ZN(n3929) );
  NOR2_X1 U4722 ( .A1(n3922), .A2(STATE_REG_SCAN_IN), .ZN(n4959) );
  OAI22_X1 U4723 ( .A1(n3925), .A2(n3924), .B1(n4437), .B2(n3923), .ZN(n3926)
         );
  AOI211_X1 U4724 ( .C1(n3927), .C2(n4381), .A(n4959), .B(n3926), .ZN(n3928)
         );
  OAI211_X1 U4725 ( .C1(n3931), .C2(n3930), .A(n3929), .B(n3928), .ZN(U3238)
         );
  INV_X1 U4726 ( .A(n3932), .ZN(n4000) );
  NAND2_X1 U4727 ( .A1(n4097), .A2(n4000), .ZN(n3933) );
  AND2_X1 U4728 ( .A1(n3934), .A2(n3933), .ZN(n4003) );
  NAND2_X1 U4729 ( .A1(n4003), .A2(n3935), .ZN(n4074) );
  INV_X1 U4730 ( .A(n4074), .ZN(n3996) );
  INV_X1 U4731 ( .A(n3936), .ZN(n3938) );
  INV_X1 U4732 ( .A(n3937), .ZN(n4008) );
  OAI211_X1 U4733 ( .C1(n3938), .C2(n4065), .A(n4008), .B(n4010), .ZN(n4066)
         );
  INV_X1 U4734 ( .A(n3939), .ZN(n4287) );
  NAND2_X1 U4735 ( .A1(n3941), .A2(n3940), .ZN(n3944) );
  NAND3_X1 U4736 ( .A1(n3944), .A2(n3943), .A3(n3942), .ZN(n3946) );
  NAND3_X1 U4737 ( .A1(n3946), .A2(n2906), .A3(n3945), .ZN(n3949) );
  NAND3_X1 U4738 ( .A1(n3949), .A2(n3948), .A3(n3947), .ZN(n3952) );
  NAND3_X1 U4739 ( .A1(n3952), .A2(n3951), .A3(n3950), .ZN(n3954) );
  NAND4_X1 U4740 ( .A1(n3954), .A2(n3953), .A3(n3968), .A4(n2180), .ZN(n3956)
         );
  NAND3_X1 U4741 ( .A1(n3956), .A2(n4020), .A3(n3955), .ZN(n3957) );
  NAND3_X1 U4742 ( .A1(n3957), .A2(n3966), .A3(n3969), .ZN(n3960) );
  NAND3_X1 U4743 ( .A1(n3960), .A2(n3959), .A3(n3958), .ZN(n3964) );
  NAND2_X1 U4744 ( .A1(n3962), .A2(n3961), .ZN(n3965) );
  INV_X1 U4745 ( .A(n3965), .ZN(n3963) );
  NAND3_X1 U4746 ( .A1(n3964), .A2(n3963), .A3(n2912), .ZN(n3978) );
  NAND2_X1 U4747 ( .A1(n3965), .A2(n3980), .ZN(n4053) );
  NOR2_X1 U4748 ( .A1(n2383), .A2(n3967), .ZN(n3970) );
  NAND4_X1 U4749 ( .A1(n3970), .A2(n2912), .A3(n3969), .A4(n3968), .ZN(n3972)
         );
  NAND2_X1 U4750 ( .A1(n3972), .A2(n3971), .ZN(n3973) );
  NAND2_X1 U4751 ( .A1(n4053), .A2(n3973), .ZN(n3977) );
  NAND2_X1 U4752 ( .A1(n3975), .A2(n3974), .ZN(n3976) );
  AOI21_X1 U4753 ( .B1(n3978), .B2(n3977), .A(n3976), .ZN(n3985) );
  NAND2_X1 U4754 ( .A1(n3980), .A2(n3979), .ZN(n4054) );
  INV_X1 U4755 ( .A(n4054), .ZN(n3982) );
  INV_X1 U4756 ( .A(n4053), .ZN(n3981) );
  AOI21_X1 U4757 ( .B1(n3983), .B2(n3982), .A(n3981), .ZN(n3984) );
  OAI21_X1 U4758 ( .B1(n3985), .B2(n3984), .A(n4055), .ZN(n3986) );
  NAND2_X1 U4759 ( .A1(n3986), .A2(n4058), .ZN(n3989) );
  NAND4_X1 U4760 ( .A1(n3989), .A2(n2259), .A3(n4056), .A4(n2925), .ZN(n3990)
         );
  AOI21_X1 U4761 ( .B1(n4287), .B2(n3990), .A(n4012), .ZN(n3992) );
  NOR3_X1 U4762 ( .A1(n4065), .A2(n3992), .A3(n3991), .ZN(n3994) );
  INV_X1 U4763 ( .A(n4070), .ZN(n3993) );
  OAI21_X1 U4764 ( .B1(n4066), .B2(n3994), .A(n3993), .ZN(n3995) );
  OAI211_X1 U4765 ( .C1(n4492), .C2(n3997), .A(n3996), .B(n3995), .ZN(n4007)
         );
  NAND2_X1 U4766 ( .A1(n3999), .A2(n3998), .ZN(n4071) );
  OR2_X1 U4767 ( .A1(n4097), .A2(n4000), .ZN(n4002) );
  NAND2_X1 U4768 ( .A1(n4004), .A2(n4078), .ZN(n4006) );
  OR2_X1 U4769 ( .A1(n4005), .A2(n4164), .ZN(n4001) );
  AND2_X1 U4770 ( .A1(n4006), .A2(n4001), .ZN(n4025) );
  NAND2_X1 U4771 ( .A1(n4002), .A2(n4025), .ZN(n4069) );
  AOI21_X1 U4772 ( .B1(n4071), .B2(n4003), .A(n4069), .ZN(n4073) );
  OR2_X1 U4773 ( .A1(n4004), .A2(n4078), .ZN(n4075) );
  NAND2_X1 U4774 ( .A1(n4005), .A2(n4164), .ZN(n4077) );
  NAND2_X1 U4775 ( .A1(n4075), .A2(n4077), .ZN(n4027) );
  AOI22_X1 U4776 ( .A1(n4007), .A2(n4073), .B1(n4006), .B2(n4027), .ZN(n4086)
         );
  INV_X1 U4777 ( .A(n4181), .ZN(n4051) );
  NAND2_X1 U4778 ( .A1(n4008), .A2(n4196), .ZN(n4216) );
  NAND2_X1 U4779 ( .A1(n4010), .A2(n4009), .ZN(n4234) );
  INV_X1 U4780 ( .A(n4234), .ZN(n4046) );
  NAND2_X1 U4781 ( .A1(n4230), .A2(n4011), .ZN(n4252) );
  INV_X1 U4782 ( .A(n4252), .ZN(n4045) );
  INV_X1 U4783 ( .A(n4012), .ZN(n4013) );
  NAND2_X1 U4784 ( .A1(n2925), .A2(n4327), .ZN(n4372) );
  NAND4_X1 U4785 ( .A1(n4016), .A2(n4015), .A3(n2908), .A4(n4014), .ZN(n4017)
         );
  NOR4_X1 U4786 ( .A1(n4372), .A2(n3271), .A3(n4017), .A4(n4598), .ZN(n4035)
         );
  INV_X1 U4787 ( .A(n4018), .ZN(n4022) );
  NAND4_X1 U4788 ( .A1(n4022), .A2(n4021), .A3(n4020), .A4(n4019), .ZN(n4023)
         );
  NOR3_X1 U4789 ( .A1(n4356), .A2(n4024), .A3(n4023), .ZN(n4034) );
  XNOR2_X1 U4790 ( .A(n4439), .B(n4586), .ZN(n4444) );
  INV_X1 U4791 ( .A(n4025), .ZN(n4026) );
  NOR2_X1 U4792 ( .A1(n4027), .A2(n4026), .ZN(n4028) );
  AND4_X1 U4793 ( .A1(n4030), .A2(n4444), .A3(n4029), .A4(n4028), .ZN(n4033)
         );
  AND2_X1 U4794 ( .A1(n4399), .A2(n4031), .ZN(n4032) );
  AND4_X1 U4795 ( .A1(n4035), .A2(n4034), .A3(n4033), .A4(n4032), .ZN(n4042)
         );
  INV_X1 U4796 ( .A(n4036), .ZN(n4038) );
  OR2_X1 U4797 ( .A1(n4038), .A2(n4037), .ZN(n4308) );
  AND2_X1 U4798 ( .A1(n4308), .A2(n4039), .ZN(n4041) );
  XNOR2_X1 U4799 ( .A(n4352), .B(n4040), .ZN(n4338) );
  INV_X1 U4800 ( .A(n4338), .ZN(n4332) );
  NAND4_X1 U4801 ( .A1(n4285), .A2(n4042), .A3(n4041), .A4(n4332), .ZN(n4043)
         );
  NOR2_X1 U4802 ( .A1(n4043), .A2(n4278), .ZN(n4044) );
  NAND3_X1 U4803 ( .A1(n4046), .A2(n4045), .A3(n4044), .ZN(n4047) );
  NOR2_X1 U4804 ( .A1(n4216), .A2(n4047), .ZN(n4050) );
  XNOR2_X1 U4805 ( .A(n4493), .B(n4208), .ZN(n4194) );
  INV_X1 U4806 ( .A(n4194), .ZN(n4199) );
  AND2_X1 U4807 ( .A1(n4199), .A2(n4048), .ZN(n4049) );
  AND4_X1 U4808 ( .A1(n4052), .A2(n4051), .A3(n4050), .A4(n4049), .ZN(n4084)
         );
  OAI21_X1 U4809 ( .B1(n4413), .B2(n4054), .A(n4053), .ZN(n4059) );
  NAND4_X1 U4810 ( .A1(n2259), .A2(n4056), .A3(n4055), .A4(n2925), .ZN(n4057)
         );
  AOI21_X1 U4811 ( .B1(n4059), .B2(n4058), .A(n4057), .ZN(n4064) );
  INV_X1 U4812 ( .A(n4060), .ZN(n4063) );
  INV_X1 U4813 ( .A(n4061), .ZN(n4062) );
  OAI21_X1 U4814 ( .B1(n4064), .B2(n4063), .A(n4062), .ZN(n4068) );
  INV_X1 U4815 ( .A(n4065), .ZN(n4067) );
  AOI21_X1 U4816 ( .B1(n4068), .B2(n4067), .A(n4066), .ZN(n4072) );
  NOR4_X1 U4817 ( .A1(n4072), .A2(n4071), .A3(n4070), .A4(n4069), .ZN(n4081)
         );
  OAI21_X1 U4818 ( .B1(n4181), .B2(n4074), .A(n4073), .ZN(n4076) );
  OAI211_X1 U4819 ( .C1(n4078), .C2(n4077), .A(n4076), .B(n4075), .ZN(n4080)
         );
  INV_X1 U4820 ( .A(n4078), .ZN(n4079) );
  OAI22_X1 U4821 ( .A1(n4081), .A2(n4080), .B1(n4079), .B2(n4164), .ZN(n4083)
         );
  MUX2_X1 U4822 ( .A(n4084), .B(n4083), .S(n4082), .Z(n4085) );
  MUX2_X1 U4823 ( .A(n4086), .B(n4085), .S(n2958), .Z(n4088) );
  XNOR2_X1 U4824 ( .A(n4088), .B(n4087), .ZN(n4096) );
  INV_X1 U4825 ( .A(n4089), .ZN(n4091) );
  NOR2_X1 U4826 ( .A1(n4091), .A2(n4090), .ZN(n4094) );
  OAI21_X1 U4827 ( .B1(n4095), .B2(n4092), .A(B_REG_SCAN_IN), .ZN(n4093) );
  OAI22_X1 U4828 ( .A1(n4096), .A2(n4095), .B1(n4094), .B2(n4093), .ZN(U3239)
         );
  MUX2_X1 U4829 ( .A(DATAO_REG_29__SCAN_IN), .B(n4097), .S(U4043), .Z(U3579)
         );
  MUX2_X1 U4830 ( .A(DATAO_REG_28__SCAN_IN), .B(n4098), .S(U4043), .Z(U3578)
         );
  MUX2_X1 U4831 ( .A(DATAO_REG_26__SCAN_IN), .B(n4493), .S(U4043), .Z(U3576)
         );
  MUX2_X1 U4832 ( .A(DATAO_REG_23__SCAN_IN), .B(n4099), .S(n4103), .Z(U3573)
         );
  MUX2_X1 U4833 ( .A(DATAO_REG_20__SCAN_IN), .B(n4525), .S(U4043), .Z(U3570)
         );
  MUX2_X1 U4834 ( .A(DATAO_REG_19__SCAN_IN), .B(n4311), .S(U4043), .Z(U3569)
         );
  MUX2_X1 U4835 ( .A(DATAO_REG_18__SCAN_IN), .B(n4549), .S(U4043), .Z(U3568)
         );
  MUX2_X1 U4836 ( .A(n4381), .B(DATAO_REG_16__SCAN_IN), .S(n4100), .Z(U3566)
         );
  MUX2_X1 U4837 ( .A(DATAO_REG_13__SCAN_IN), .B(n4586), .S(n4103), .Z(U3563)
         );
  MUX2_X1 U4838 ( .A(DATAO_REG_12__SCAN_IN), .B(n4101), .S(U4043), .Z(U3562)
         );
  MUX2_X1 U4839 ( .A(DATAO_REG_11__SCAN_IN), .B(n4585), .S(U4043), .Z(U3561)
         );
  MUX2_X1 U4840 ( .A(DATAO_REG_10__SCAN_IN), .B(n4102), .S(U4043), .Z(U3560)
         );
  MUX2_X1 U4841 ( .A(DATAO_REG_9__SCAN_IN), .B(n4459), .S(n4103), .Z(U3559) );
  MUX2_X1 U4842 ( .A(DATAO_REG_8__SCAN_IN), .B(n4104), .S(U4043), .Z(U3558) );
  MUX2_X1 U4843 ( .A(DATAO_REG_4__SCAN_IN), .B(n4105), .S(U4043), .Z(U3554) );
  MUX2_X1 U4844 ( .A(DATAO_REG_3__SCAN_IN), .B(n2909), .S(U4043), .Z(U3553) );
  MUX2_X1 U4845 ( .A(DATAO_REG_2__SCAN_IN), .B(n4475), .S(U4043), .Z(U3552) );
  MUX2_X1 U4846 ( .A(DATAO_REG_1__SCAN_IN), .B(n4602), .S(U4043), .Z(U3551) );
  NAND2_X1 U4847 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n4108) );
  AOI211_X1 U4848 ( .C1(n4108), .C2(n4107), .A(n4106), .B(n4970), .ZN(n4109)
         );
  INV_X1 U4849 ( .A(n4109), .ZN(n4116) );
  AOI22_X1 U4850 ( .A1(n4994), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n4115) );
  NAND2_X1 U4851 ( .A1(n4158), .A2(n4945), .ZN(n4114) );
  OAI211_X1 U4852 ( .C1(n4112), .C2(n4111), .A(n4974), .B(n4110), .ZN(n4113)
         );
  NAND4_X1 U4853 ( .A1(n4116), .A2(n4115), .A3(n4114), .A4(n4113), .ZN(U3241)
         );
  OAI211_X1 U4854 ( .C1(n4119), .C2(n4118), .A(n4117), .B(n4996), .ZN(n4128)
         );
  NOR2_X1 U4855 ( .A1(n5000), .A2(n4120), .ZN(n4121) );
  AOI211_X1 U4856 ( .C1(n4994), .C2(ADDR_REG_11__SCAN_IN), .A(n4122), .B(n4121), .ZN(n4127) );
  OAI211_X1 U4857 ( .C1(n4125), .C2(n4124), .A(n4123), .B(n4974), .ZN(n4126)
         );
  NAND3_X1 U4858 ( .A1(n4128), .A2(n4127), .A3(n4126), .ZN(U3251) );
  XNOR2_X1 U4859 ( .A(n4129), .B(REG1_REG_12__SCAN_IN), .ZN(n4138) );
  XOR2_X1 U4860 ( .A(REG2_REG_12__SCAN_IN), .B(n4130), .Z(n4131) );
  NAND2_X1 U4861 ( .A1(n4974), .A2(n4131), .ZN(n4133) );
  NAND2_X1 U4862 ( .A1(n4133), .A2(n4132), .ZN(n4136) );
  NOR2_X1 U4863 ( .A1(n5000), .A2(n4134), .ZN(n4135) );
  AOI211_X1 U4864 ( .C1(n4994), .C2(ADDR_REG_12__SCAN_IN), .A(n4136), .B(n4135), .ZN(n4137) );
  OAI21_X1 U4865 ( .B1(n4138), .B2(n4970), .A(n4137), .ZN(U3252) );
  INV_X1 U4866 ( .A(REG2_REG_13__SCAN_IN), .ZN(n4139) );
  MUX2_X1 U4867 ( .A(n4139), .B(REG2_REG_13__SCAN_IN), .S(n4939), .Z(n4141) );
  XOR2_X1 U4868 ( .A(n4141), .B(n4140), .Z(n4150) );
  OAI211_X1 U4869 ( .C1(n4144), .C2(n4143), .A(n4142), .B(n4996), .ZN(n4149)
         );
  INV_X1 U4870 ( .A(n4939), .ZN(n4145) );
  NOR2_X1 U4871 ( .A1(n5000), .A2(n4145), .ZN(n4146) );
  AOI211_X1 U4872 ( .C1(n4994), .C2(ADDR_REG_13__SCAN_IN), .A(n4147), .B(n4146), .ZN(n4148) );
  OAI211_X1 U4873 ( .C1(n4989), .C2(n4150), .A(n4149), .B(n4148), .ZN(U3253)
         );
  XOR2_X1 U4874 ( .A(REG1_REG_14__SCAN_IN), .B(n4151), .Z(n4160) );
  INV_X1 U4875 ( .A(ADDR_REG_14__SCAN_IN), .ZN(n4153) );
  OAI21_X1 U4876 ( .B1(n4978), .B2(n4153), .A(n4152), .ZN(n4157) );
  AOI211_X1 U4877 ( .C1(n4772), .C2(n4155), .A(n4989), .B(n4154), .ZN(n4156)
         );
  AOI211_X1 U4878 ( .C1(n4158), .C2(n4938), .A(n4157), .B(n4156), .ZN(n4159)
         );
  OAI21_X1 U4879 ( .B1(n4160), .B2(n4970), .A(n4159), .ZN(U3254) );
  INV_X1 U4880 ( .A(n4874), .ZN(n4163) );
  NAND2_X1 U4881 ( .A1(n4163), .A2(n4480), .ZN(n4169) );
  INV_X1 U4882 ( .A(n4164), .ZN(n4165) );
  NAND2_X1 U4883 ( .A1(n4165), .A2(n4582), .ZN(n4166) );
  NAND2_X1 U4884 ( .A1(n4167), .A2(n4166), .ZN(n4871) );
  NAND2_X1 U4885 ( .A1(n4484), .A2(n4871), .ZN(n4168) );
  OAI211_X1 U4886 ( .C1(n4484), .C2(n4811), .A(n4169), .B(n4168), .ZN(U3261)
         );
  NAND2_X1 U4887 ( .A1(n4170), .A2(n4467), .ZN(n4177) );
  INV_X1 U4888 ( .A(n4171), .ZN(n4173) );
  OAI22_X1 U4889 ( .A1(n4173), .A2(n4449), .B1(n4172), .B2(n4461), .ZN(n4174)
         );
  OAI21_X1 U4890 ( .B1(n4175), .B2(n4174), .A(n4484), .ZN(n4176) );
  OAI211_X1 U4891 ( .C1(n4484), .C2(n4178), .A(n4177), .B(n4176), .ZN(U3354)
         );
  INV_X1 U4892 ( .A(n4498), .ZN(n4193) );
  XOR2_X1 U4893 ( .A(n4181), .B(n4180), .Z(n4182) );
  OAI21_X1 U4894 ( .B1(n4206), .B2(n4185), .A(n4183), .ZN(n4878) );
  NOR2_X1 U4895 ( .A1(n4878), .A2(n4449), .ZN(n4191) );
  OAI22_X1 U4896 ( .A1(n4424), .A2(n4185), .B1(n4184), .B2(n4484), .ZN(n4186)
         );
  AOI21_X1 U4897 ( .B1(n4493), .B2(n4474), .A(n4186), .ZN(n4189) );
  NAND2_X1 U4898 ( .A1(n4187), .A2(n4481), .ZN(n4188) );
  OAI211_X1 U4899 ( .C1(n4495), .C2(n4295), .A(n4189), .B(n4188), .ZN(n4190)
         );
  AOI211_X1 U4900 ( .C1(n4497), .C2(n4484), .A(n4191), .B(n4190), .ZN(n4192)
         );
  OAI21_X1 U4901 ( .B1(n4193), .B2(n4304), .A(n4192), .ZN(U3263) );
  XNOR2_X1 U4902 ( .A(n4195), .B(n4194), .ZN(n4500) );
  INV_X1 U4903 ( .A(n4500), .ZN(n4213) );
  INV_X1 U4904 ( .A(n4196), .ZN(n4197) );
  NOR2_X1 U4905 ( .A1(n4198), .A2(n4197), .ZN(n4200) );
  XNOR2_X1 U4906 ( .A(n4200), .B(n4199), .ZN(n4205) );
  OAI22_X1 U4907 ( .A1(n4201), .A2(n4547), .B1(n4208), .B2(n4572), .ZN(n4202)
         );
  AOI21_X1 U4908 ( .B1(n4203), .B2(n4601), .A(n4202), .ZN(n4204) );
  OAI21_X1 U4909 ( .B1(n4205), .B2(n4441), .A(n4204), .ZN(n4499) );
  INV_X1 U4910 ( .A(n4206), .ZN(n4207) );
  OAI21_X1 U4911 ( .B1(n4218), .B2(n4208), .A(n4207), .ZN(n4882) );
  NOR2_X1 U4912 ( .A1(n4882), .A2(n4449), .ZN(n4211) );
  OAI22_X1 U4913 ( .A1(n4209), .A2(n4461), .B1(n4809), .B2(n4484), .ZN(n4210)
         );
  AOI211_X1 U4914 ( .C1(n4499), .C2(n4484), .A(n4211), .B(n4210), .ZN(n4212)
         );
  OAI21_X1 U4915 ( .B1(n4213), .B2(n4304), .A(n4212), .ZN(U3264) );
  XOR2_X1 U4916 ( .A(n4216), .B(n4214), .Z(n4509) );
  INV_X1 U4917 ( .A(n4509), .ZN(n4228) );
  XOR2_X1 U4918 ( .A(n4216), .B(n4215), .Z(n4217) );
  NOR2_X1 U4919 ( .A1(n4217), .A2(n4441), .ZN(n4508) );
  NAND2_X1 U4920 ( .A1(n4242), .A2(n4503), .ZN(n4219) );
  NAND2_X1 U4921 ( .A1(n2432), .A2(n4219), .ZN(n4886) );
  AOI22_X1 U4922 ( .A1(n4220), .A2(n4481), .B1(REG2_REG_25__SCAN_IN), .B2(
        n4454), .ZN(n4221) );
  OAI21_X1 U4923 ( .B1(n4222), .B2(n4424), .A(n4221), .ZN(n4224) );
  NOR2_X1 U4924 ( .A1(n4506), .A2(n4295), .ZN(n4223) );
  AOI211_X1 U4925 ( .C1(n4474), .C2(n4504), .A(n4224), .B(n4223), .ZN(n4225)
         );
  OAI21_X1 U4926 ( .B1(n4886), .B2(n4449), .A(n4225), .ZN(n4226) );
  AOI21_X1 U4927 ( .B1(n4508), .B2(n4484), .A(n4226), .ZN(n4227) );
  OAI21_X1 U4928 ( .B1(n4228), .B2(n4304), .A(n4227), .ZN(U3265) );
  XNOR2_X1 U4929 ( .A(n4229), .B(n4234), .ZN(n4513) );
  INV_X1 U4930 ( .A(n4513), .ZN(n4247) );
  INV_X1 U4931 ( .A(n4230), .ZN(n4231) );
  NOR2_X1 U4932 ( .A1(n4232), .A2(n4231), .ZN(n4233) );
  XOR2_X1 U4933 ( .A(n4234), .B(n4233), .Z(n4239) );
  OAI22_X1 U4934 ( .A1(n4272), .A2(n4547), .B1(n4235), .B2(n4572), .ZN(n4236)
         );
  AOI21_X1 U4935 ( .B1(n4237), .B2(n4601), .A(n4236), .ZN(n4238) );
  OAI21_X1 U4936 ( .B1(n4239), .B2(n4441), .A(n4238), .ZN(n4512) );
  NAND2_X1 U4937 ( .A1(n4257), .A2(n4240), .ZN(n4241) );
  NAND2_X1 U4938 ( .A1(n4242), .A2(n4241), .ZN(n4890) );
  AOI22_X1 U4939 ( .A1(n4243), .A2(n4481), .B1(REG2_REG_24__SCAN_IN), .B2(
        n4454), .ZN(n4244) );
  OAI21_X1 U4940 ( .B1(n4890), .B2(n4449), .A(n4244), .ZN(n4245) );
  AOI21_X1 U4941 ( .B1(n4512), .B2(n4484), .A(n4245), .ZN(n4246) );
  OAI21_X1 U4942 ( .B1(n4247), .B2(n4304), .A(n4246), .ZN(U3266) );
  XOR2_X1 U4943 ( .A(n4252), .B(n4248), .Z(n4516) );
  INV_X1 U4944 ( .A(n4516), .ZN(n4263) );
  NAND2_X1 U4945 ( .A1(n4288), .A2(n4287), .ZN(n4249) );
  NAND2_X1 U4946 ( .A1(n4249), .A2(n4285), .ZN(n4290) );
  NAND2_X1 U4947 ( .A1(n4290), .A2(n4250), .ZN(n4265) );
  INV_X1 U4948 ( .A(n4278), .ZN(n4266) );
  NAND2_X1 U4949 ( .A1(n4265), .A2(n4266), .ZN(n4264) );
  NAND2_X1 U4950 ( .A1(n4264), .A2(n4251), .ZN(n4253) );
  XNOR2_X1 U4951 ( .A(n4253), .B(n4252), .ZN(n4256) );
  OAI22_X1 U4952 ( .A1(n4527), .A2(n4547), .B1(n4572), .B2(n4258), .ZN(n4254)
         );
  AOI21_X1 U4953 ( .B1(n4504), .B2(n4601), .A(n4254), .ZN(n4255) );
  OAI21_X1 U4954 ( .B1(n4256), .B2(n4441), .A(n4255), .ZN(n4515) );
  OAI21_X1 U4955 ( .B1(n4275), .B2(n4258), .A(n4257), .ZN(n4894) );
  AOI22_X1 U4956 ( .A1(n4259), .A2(n4481), .B1(REG2_REG_23__SCAN_IN), .B2(
        n4454), .ZN(n4260) );
  OAI21_X1 U4957 ( .B1(n4894), .B2(n4449), .A(n4260), .ZN(n4261) );
  AOI21_X1 U4958 ( .B1(n4515), .B2(n4484), .A(n4261), .ZN(n4262) );
  OAI21_X1 U4959 ( .B1(n4263), .B2(n4304), .A(n4262), .ZN(U3267) );
  OAI21_X1 U4960 ( .B1(n4266), .B2(n4265), .A(n4264), .ZN(n4267) );
  NAND2_X1 U4961 ( .A1(n4267), .A2(n4595), .ZN(n4271) );
  AOI22_X1 U4962 ( .A1(n4269), .A2(n4584), .B1(n4268), .B2(n4582), .ZN(n4270)
         );
  OAI211_X1 U4963 ( .C1(n4272), .C2(n4564), .A(n4271), .B(n4270), .ZN(n4520)
         );
  NOR2_X1 U4964 ( .A1(n4291), .A2(n4273), .ZN(n4274) );
  OR2_X1 U4965 ( .A1(n4275), .A2(n4274), .ZN(n4898) );
  AOI22_X1 U4966 ( .A1(n4276), .A2(n4481), .B1(REG2_REG_22__SCAN_IN), .B2(
        n4454), .ZN(n4277) );
  OAI21_X1 U4967 ( .B1(n4898), .B2(n4449), .A(n4277), .ZN(n4282) );
  NOR2_X1 U4968 ( .A1(n4279), .A2(n4278), .ZN(n4519) );
  INV_X1 U4969 ( .A(n4521), .ZN(n4280) );
  NOR3_X1 U4970 ( .A1(n4519), .A2(n4280), .A3(n4304), .ZN(n4281) );
  AOI211_X1 U4971 ( .C1(n4484), .C2(n4520), .A(n4282), .B(n4281), .ZN(n4283)
         );
  INV_X1 U4972 ( .A(n4283), .ZN(U3268) );
  XNOR2_X1 U4973 ( .A(n4284), .B(n4285), .ZN(n4530) );
  INV_X1 U4974 ( .A(n4530), .ZN(n4305) );
  INV_X1 U4975 ( .A(n4285), .ZN(n4286) );
  NAND3_X1 U4976 ( .A1(n4288), .A2(n4287), .A3(n4286), .ZN(n4289) );
  AOI21_X1 U4977 ( .B1(n4290), .B2(n4289), .A(n4441), .ZN(n4529) );
  INV_X1 U4978 ( .A(n4291), .ZN(n4292) );
  OAI21_X1 U4979 ( .B1(n4318), .B2(n4300), .A(n4292), .ZN(n4902) );
  NOR2_X1 U4980 ( .A1(n4902), .A2(n4449), .ZN(n4302) );
  OAI22_X1 U4981 ( .A1(n4527), .A2(n4295), .B1(n4294), .B2(n4293), .ZN(n4296)
         );
  INV_X1 U4982 ( .A(n4296), .ZN(n4299) );
  AOI22_X1 U4983 ( .A1(n4297), .A2(n4481), .B1(n4386), .B2(
        REG2_REG_21__SCAN_IN), .ZN(n4298) );
  OAI211_X1 U4984 ( .C1(n4300), .C2(n4424), .A(n4299), .B(n4298), .ZN(n4301)
         );
  AOI211_X1 U4985 ( .C1(n4529), .C2(n4484), .A(n4302), .B(n4301), .ZN(n4303)
         );
  OAI21_X1 U4986 ( .B1(n4305), .B2(n4304), .A(n4303), .ZN(U3269) );
  XNOR2_X1 U4987 ( .A(n4306), .B(n4308), .ZN(n4317) );
  NAND2_X1 U4988 ( .A1(n2168), .A2(n4307), .ZN(n4309) );
  XNOR2_X1 U4989 ( .A(n4309), .B(n4308), .ZN(n4315) );
  AOI22_X1 U4990 ( .A1(n4311), .A2(n4584), .B1(n4310), .B2(n4582), .ZN(n4312)
         );
  OAI21_X1 U4991 ( .B1(n4313), .B2(n4564), .A(n4312), .ZN(n4314) );
  AOI21_X1 U4992 ( .B1(n4315), .B2(n4595), .A(n4314), .ZN(n4316) );
  OAI21_X1 U4993 ( .B1(n4317), .B2(n4418), .A(n4316), .ZN(n4533) );
  INV_X1 U4994 ( .A(n4533), .ZN(n4326) );
  INV_X1 U4995 ( .A(n4317), .ZN(n4534) );
  INV_X1 U4996 ( .A(n4340), .ZN(n4321) );
  INV_X1 U4997 ( .A(n4318), .ZN(n4319) );
  OAI21_X1 U4998 ( .B1(n4321), .B2(n4320), .A(n4319), .ZN(n4906) );
  AOI22_X1 U4999 ( .A1(REG2_REG_20__SCAN_IN), .A2(n4454), .B1(n4322), .B2(
        n4481), .ZN(n4323) );
  OAI21_X1 U5000 ( .B1(n4906), .B2(n4449), .A(n4323), .ZN(n4324) );
  AOI21_X1 U5001 ( .B1(n4534), .B2(n4483), .A(n4324), .ZN(n4325) );
  OAI21_X1 U5002 ( .B1(n4326), .B2(n4386), .A(n4325), .ZN(U3270) );
  NAND2_X1 U5003 ( .A1(n4328), .A2(n4327), .ZN(n4348) );
  INV_X1 U5004 ( .A(n4329), .ZN(n4331) );
  OAI21_X1 U5005 ( .B1(n4348), .B2(n4331), .A(n4330), .ZN(n4333) );
  XNOR2_X1 U5006 ( .A(n4333), .B(n4332), .ZN(n4337) );
  OAI22_X1 U5007 ( .A1(n4334), .A2(n4547), .B1(n4572), .B2(n4341), .ZN(n4335)
         );
  AOI21_X1 U5008 ( .B1(n4525), .B2(n4601), .A(n4335), .ZN(n4336) );
  OAI21_X1 U5009 ( .B1(n4337), .B2(n4441), .A(n4336), .ZN(n4537) );
  INV_X1 U5010 ( .A(n4537), .ZN(n4347) );
  XNOR2_X1 U5011 ( .A(n4339), .B(n4338), .ZN(n4538) );
  INV_X1 U5012 ( .A(n4358), .ZN(n4342) );
  OAI21_X1 U5013 ( .B1(n4342), .B2(n4341), .A(n4340), .ZN(n4910) );
  AOI22_X1 U5014 ( .A1(n4454), .A2(REG2_REG_19__SCAN_IN), .B1(n4343), .B2(
        n4481), .ZN(n4344) );
  OAI21_X1 U5015 ( .B1(n4910), .B2(n4449), .A(n4344), .ZN(n4345) );
  AOI21_X1 U5016 ( .B1(n4538), .B2(n4467), .A(n4345), .ZN(n4346) );
  OAI21_X1 U5017 ( .B1(n4347), .B2(n4386), .A(n4346), .ZN(U3271) );
  XOR2_X1 U5018 ( .A(n4356), .B(n4348), .Z(n4354) );
  AOI22_X1 U5019 ( .A1(n4350), .A2(n4584), .B1(n4349), .B2(n4582), .ZN(n4351)
         );
  OAI21_X1 U5020 ( .B1(n4352), .B2(n4564), .A(n4351), .ZN(n4353) );
  AOI21_X1 U5021 ( .B1(n4354), .B2(n4595), .A(n4353), .ZN(n4542) );
  OAI21_X1 U5022 ( .B1(n4357), .B2(n4356), .A(n4355), .ZN(n4540) );
  INV_X1 U5023 ( .A(n4376), .ZN(n4361) );
  OAI211_X1 U5024 ( .C1(n4361), .C2(n4360), .A(n4359), .B(n4358), .ZN(n4541)
         );
  NOR2_X1 U5025 ( .A1(n4541), .A2(n4362), .ZN(n4365) );
  OAI22_X1 U5026 ( .A1(n4484), .A2(n4820), .B1(n4363), .B2(n4461), .ZN(n4364)
         );
  AOI211_X1 U5027 ( .C1(n4540), .C2(n4467), .A(n4365), .B(n4364), .ZN(n4366)
         );
  OAI21_X1 U5028 ( .B1(n4542), .B2(n4386), .A(n4366), .ZN(U3272) );
  XNOR2_X1 U5029 ( .A(n4367), .B(n4372), .ZN(n4368) );
  NAND2_X1 U5030 ( .A1(n4368), .A2(n4595), .ZN(n4550) );
  NAND2_X1 U5031 ( .A1(n4411), .A2(n4369), .ZN(n4371) );
  NAND2_X1 U5032 ( .A1(n4371), .A2(n4370), .ZN(n4374) );
  INV_X1 U5033 ( .A(n4372), .ZN(n4373) );
  XNOR2_X1 U5034 ( .A(n4374), .B(n4373), .ZN(n4545) );
  OR2_X1 U5035 ( .A1(n4403), .A2(n4546), .ZN(n4375) );
  NAND2_X1 U5036 ( .A1(n4376), .A2(n4375), .ZN(n4915) );
  OAI22_X1 U5037 ( .A1(n4484), .A2(n4378), .B1(n4377), .B2(n4461), .ZN(n4379)
         );
  AOI21_X1 U5038 ( .B1(n4380), .B2(n4478), .A(n4379), .ZN(n4383) );
  AOI22_X1 U5039 ( .A1(n4476), .A2(n4549), .B1(n4474), .B2(n4381), .ZN(n4382)
         );
  OAI211_X1 U5040 ( .C1(n4915), .C2(n4449), .A(n4383), .B(n4382), .ZN(n4384)
         );
  AOI21_X1 U5041 ( .B1(n4545), .B2(n4467), .A(n4384), .ZN(n4385) );
  OAI21_X1 U5042 ( .B1(n4386), .B2(n4550), .A(n4385), .ZN(U3273) );
  XNOR2_X1 U5043 ( .A(n4388), .B(n4387), .ZN(n4393) );
  NAND2_X1 U5044 ( .A1(n4570), .A2(n4584), .ZN(n4390) );
  NAND2_X1 U5045 ( .A1(n4405), .A2(n4582), .ZN(n4389) );
  OAI211_X1 U5046 ( .C1(n4391), .C2(n4564), .A(n4390), .B(n4389), .ZN(n4392)
         );
  AOI21_X1 U5047 ( .B1(n4393), .B2(n4595), .A(n4392), .ZN(n4557) );
  NAND2_X1 U5048 ( .A1(n4395), .A2(n4394), .ZN(n4398) );
  NAND2_X1 U5049 ( .A1(n4398), .A2(n4396), .ZN(n4402) );
  NAND2_X1 U5050 ( .A1(n4398), .A2(n4397), .ZN(n4400) );
  NAND2_X1 U5051 ( .A1(n4400), .A2(n4399), .ZN(n4401) );
  AND2_X1 U5052 ( .A1(n4402), .A2(n4401), .ZN(n4555) );
  AOI21_X1 U5053 ( .B1(n4405), .B2(n4404), .A(n4403), .ZN(n4919) );
  INV_X1 U5054 ( .A(n4919), .ZN(n4408) );
  AOI22_X1 U5055 ( .A1(n4454), .A2(REG2_REG_16__SCAN_IN), .B1(n4406), .B2(
        n4481), .ZN(n4407) );
  OAI21_X1 U5056 ( .B1(n4408), .B2(n4449), .A(n4407), .ZN(n4409) );
  AOI21_X1 U5057 ( .B1(n4555), .B2(n4467), .A(n4409), .ZN(n4410) );
  OAI21_X1 U5058 ( .B1(n4557), .B2(n4454), .A(n4410), .ZN(U3274) );
  OAI21_X1 U5059 ( .B1(n4412), .B2(n4416), .A(n4411), .ZN(n4576) );
  INV_X1 U5060 ( .A(n4576), .ZN(n4430) );
  INV_X1 U5061 ( .A(n4413), .ZN(n4417) );
  INV_X1 U5062 ( .A(n4414), .ZN(n4415) );
  AOI21_X1 U5063 ( .B1(n4417), .B2(n4416), .A(n4415), .ZN(n4419) );
  OAI22_X1 U5064 ( .A1(n4419), .A2(n4441), .B1(n4430), .B2(n4418), .ZN(n4574)
         );
  NAND2_X1 U5065 ( .A1(n4574), .A2(n4484), .ZN(n4428) );
  OAI21_X1 U5066 ( .B1(n2427), .B2(n4573), .A(n4420), .ZN(n4928) );
  INV_X1 U5067 ( .A(n4928), .ZN(n4426) );
  AOI22_X1 U5068 ( .A1(n4476), .A2(n4570), .B1(n4474), .B2(n4586), .ZN(n4423)
         );
  AOI22_X1 U5069 ( .A1(n4454), .A2(REG2_REG_14__SCAN_IN), .B1(n4421), .B2(
        n4481), .ZN(n4422) );
  OAI211_X1 U5070 ( .C1(n4573), .C2(n4424), .A(n4423), .B(n4422), .ZN(n4425)
         );
  AOI21_X1 U5071 ( .B1(n4426), .B2(n4480), .A(n4425), .ZN(n4427) );
  OAI211_X1 U5072 ( .C1(n4430), .C2(n4429), .A(n4428), .B(n4427), .ZN(U3276)
         );
  INV_X1 U5073 ( .A(n4431), .ZN(n4432) );
  AOI21_X1 U5074 ( .B1(n4434), .B2(n4433), .A(n4432), .ZN(n4435) );
  XOR2_X1 U5075 ( .A(n4444), .B(n4435), .Z(n4442) );
  OAI22_X1 U5076 ( .A1(n4437), .A2(n4564), .B1(n4436), .B2(n4547), .ZN(n4438)
         );
  AOI21_X1 U5077 ( .B1(n4439), .B2(n4582), .A(n4438), .ZN(n4440) );
  OAI21_X1 U5078 ( .B1(n4442), .B2(n4441), .A(n4440), .ZN(n4578) );
  INV_X1 U5079 ( .A(n4578), .ZN(n4455) );
  XOR2_X1 U5080 ( .A(n4444), .B(n4443), .Z(n4579) );
  OR2_X1 U5081 ( .A1(n4446), .A2(n4445), .ZN(n4447) );
  NAND2_X1 U5082 ( .A1(n4448), .A2(n4447), .ZN(n4932) );
  NOR2_X1 U5083 ( .A1(n4932), .A2(n4449), .ZN(n4452) );
  OAI22_X1 U5084 ( .A1(n4484), .A2(n4139), .B1(n4450), .B2(n4461), .ZN(n4451)
         );
  AOI211_X1 U5085 ( .C1(n4579), .C2(n4467), .A(n4452), .B(n4451), .ZN(n4453)
         );
  OAI21_X1 U5086 ( .B1(n4455), .B2(n4454), .A(n4453), .ZN(U3277) );
  NAND2_X1 U5087 ( .A1(n4457), .A2(n4456), .ZN(n4472) );
  AOI22_X1 U5088 ( .A1(n4476), .A2(n4459), .B1(n4478), .B2(n4458), .ZN(n4471)
         );
  AND2_X1 U5089 ( .A1(n4474), .A2(n4460), .ZN(n4465) );
  OAI22_X1 U5090 ( .A1(n4484), .A2(n4463), .B1(n4462), .B2(n4461), .ZN(n4464)
         );
  AOI211_X1 U5091 ( .C1(n4466), .C2(n4480), .A(n4465), .B(n4464), .ZN(n4470)
         );
  NAND2_X1 U5092 ( .A1(n4468), .A2(n4467), .ZN(n4469) );
  NAND4_X1 U5093 ( .A1(n4472), .A2(n4471), .A3(n4470), .A4(n4469), .ZN(U3282)
         );
  AOI22_X1 U5094 ( .A1(n4476), .A2(n4475), .B1(n4474), .B2(n4473), .ZN(n4489)
         );
  AOI22_X1 U5095 ( .A1(n4480), .A2(n4479), .B1(n4478), .B2(n4477), .ZN(n4488)
         );
  AOI22_X1 U5096 ( .A1(n4483), .A2(n4482), .B1(REG3_REG_1__SCAN_IN), .B2(n4481), .ZN(n4487) );
  MUX2_X1 U5097 ( .A(n2573), .B(n4485), .S(n4484), .Z(n4486) );
  NAND4_X1 U5098 ( .A1(n4489), .A2(n4488), .A3(n4487), .A4(n4486), .ZN(U3289)
         );
  NAND2_X1 U5099 ( .A1(n5043), .A2(n4871), .ZN(n4491) );
  NAND2_X1 U5100 ( .A1(n2210), .A2(REG1_REG_30__SCAN_IN), .ZN(n4490) );
  OAI211_X1 U5101 ( .C1(n4874), .C2(n4594), .A(n4491), .B(n4490), .ZN(U3548)
         );
  AOI22_X1 U5102 ( .A1(n4493), .A2(n4584), .B1(n4492), .B2(n4582), .ZN(n4494)
         );
  OAI21_X1 U5103 ( .B1(n4495), .B2(n4564), .A(n4494), .ZN(n4496) );
  INV_X1 U5104 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4501) );
  AOI21_X1 U5105 ( .B1(n4500), .B2(n4596), .A(n4499), .ZN(n4879) );
  MUX2_X1 U5106 ( .A(n4501), .B(n4879), .S(n5043), .Z(n4502) );
  OAI21_X1 U5107 ( .B1(n4594), .B2(n4882), .A(n4502), .ZN(U3544) );
  AOI22_X1 U5108 ( .A1(n4504), .A2(n4584), .B1(n4503), .B2(n4582), .ZN(n4505)
         );
  OAI21_X1 U5109 ( .B1(n4506), .B2(n4564), .A(n4505), .ZN(n4507) );
  AOI211_X1 U5110 ( .C1(n4509), .C2(n4596), .A(n4508), .B(n4507), .ZN(n4883)
         );
  MUX2_X1 U5111 ( .A(n4510), .B(n4883), .S(n5043), .Z(n4511) );
  OAI21_X1 U5112 ( .B1(n4594), .B2(n4886), .A(n4511), .ZN(U3543) );
  AOI21_X1 U5113 ( .B1(n4513), .B2(n4596), .A(n4512), .ZN(n4887) );
  MUX2_X1 U5114 ( .A(n4666), .B(n4887), .S(n5043), .Z(n4514) );
  OAI21_X1 U5115 ( .B1(n4594), .B2(n4890), .A(n4514), .ZN(U3542) );
  AOI21_X1 U5116 ( .B1(n4516), .B2(n4596), .A(n4515), .ZN(n4891) );
  MUX2_X1 U5117 ( .A(n4517), .B(n4891), .S(n5043), .Z(n4518) );
  OAI21_X1 U5118 ( .B1(n4594), .B2(n4894), .A(n4518), .ZN(U3541) );
  NOR2_X1 U5119 ( .A1(n4519), .A2(n4543), .ZN(n4522) );
  AOI21_X1 U5120 ( .B1(n4522), .B2(n4521), .A(n4520), .ZN(n4895) );
  MUX2_X1 U5121 ( .A(n4659), .B(n4895), .S(n5043), .Z(n4523) );
  OAI21_X1 U5122 ( .B1(n4594), .B2(n4898), .A(n4523), .ZN(U3540) );
  AOI22_X1 U5123 ( .A1(n4525), .A2(n4584), .B1(n4582), .B2(n4524), .ZN(n4526)
         );
  OAI21_X1 U5124 ( .B1(n4527), .B2(n4564), .A(n4526), .ZN(n4528) );
  AOI211_X1 U5125 ( .C1(n4530), .C2(n4596), .A(n4529), .B(n4528), .ZN(n4899)
         );
  MUX2_X1 U5126 ( .A(n4531), .B(n4899), .S(n5043), .Z(n4532) );
  OAI21_X1 U5127 ( .B1(n4594), .B2(n4902), .A(n4532), .ZN(U3539) );
  INV_X1 U5128 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4535) );
  AOI21_X1 U5129 ( .B1(n5037), .B2(n4534), .A(n4533), .ZN(n4903) );
  MUX2_X1 U5130 ( .A(n4535), .B(n4903), .S(n5043), .Z(n4536) );
  OAI21_X1 U5131 ( .B1(n4594), .B2(n4906), .A(n4536), .ZN(U3538) );
  AOI21_X1 U5132 ( .B1(n4596), .B2(n4538), .A(n4537), .ZN(n4907) );
  MUX2_X1 U5133 ( .A(n2535), .B(n4907), .S(n5043), .Z(n4539) );
  OAI21_X1 U5134 ( .B1(n4594), .B2(n4910), .A(n4539), .ZN(U3537) );
  INV_X1 U5135 ( .A(n4540), .ZN(n4544) );
  OAI211_X1 U5136 ( .C1(n4544), .C2(n4543), .A(n4542), .B(n4541), .ZN(n4911)
         );
  MUX2_X1 U5137 ( .A(REG1_REG_18__SCAN_IN), .B(n4911), .S(n5043), .Z(U3536) );
  NAND2_X1 U5138 ( .A1(n4545), .A2(n4596), .ZN(n4552) );
  OAI22_X1 U5139 ( .A1(n4565), .A2(n4547), .B1(n4572), .B2(n4546), .ZN(n4548)
         );
  AOI21_X1 U5140 ( .B1(n4549), .B2(n4601), .A(n4548), .ZN(n4551) );
  NAND3_X1 U5141 ( .A1(n4552), .A2(n4551), .A3(n4550), .ZN(n4912) );
  MUX2_X1 U5142 ( .A(n4912), .B(REG1_REG_17__SCAN_IN), .S(n2210), .Z(n4553) );
  INV_X1 U5143 ( .A(n4553), .ZN(n4554) );
  OAI21_X1 U5144 ( .B1(n4594), .B2(n4915), .A(n4554), .ZN(U3535) );
  NAND2_X1 U5145 ( .A1(n4555), .A2(n4596), .ZN(n4556) );
  NAND2_X1 U5146 ( .A1(n4557), .A2(n4556), .ZN(n4916) );
  MUX2_X1 U5147 ( .A(n4916), .B(REG1_REG_16__SCAN_IN), .S(n2210), .Z(n4558) );
  AOI21_X1 U5148 ( .B1(n4559), .B2(n4919), .A(n4558), .ZN(n4560) );
  INV_X1 U5149 ( .A(n4560), .ZN(U3534) );
  AOI22_X1 U5150 ( .A1(n4562), .A2(n4584), .B1(n4582), .B2(n4561), .ZN(n4563)
         );
  OAI21_X1 U5151 ( .B1(n4565), .B2(n4564), .A(n4563), .ZN(n4567) );
  AOI211_X1 U5152 ( .C1(n4596), .C2(n4568), .A(n4567), .B(n4566), .ZN(n4921)
         );
  MUX2_X1 U5153 ( .A(n4840), .B(n4921), .S(n5043), .Z(n4569) );
  OAI21_X1 U5154 ( .B1(n4594), .B2(n4924), .A(n4569), .ZN(U3533) );
  AOI22_X1 U5155 ( .A1(n4570), .A2(n4601), .B1(n4584), .B2(n4586), .ZN(n4571)
         );
  OAI21_X1 U5156 ( .B1(n4573), .B2(n4572), .A(n4571), .ZN(n4575) );
  AOI211_X1 U5157 ( .C1(n5037), .C2(n4576), .A(n4575), .B(n4574), .ZN(n4925)
         );
  MUX2_X1 U5158 ( .A(n4759), .B(n4925), .S(n5043), .Z(n4577) );
  OAI21_X1 U5159 ( .B1(n4594), .B2(n4928), .A(n4577), .ZN(U3532) );
  AOI21_X1 U5160 ( .B1(n4596), .B2(n4579), .A(n4578), .ZN(n4929) );
  MUX2_X1 U5161 ( .A(n4580), .B(n4929), .S(n5043), .Z(n4581) );
  OAI21_X1 U5162 ( .B1(n4594), .B2(n4932), .A(n4581), .ZN(U3531) );
  NAND2_X1 U5163 ( .A1(n4583), .A2(n4582), .ZN(n4588) );
  AOI22_X1 U5164 ( .A1(n4586), .A2(n4601), .B1(n4585), .B2(n4584), .ZN(n4587)
         );
  NAND2_X1 U5165 ( .A1(n4588), .A2(n4587), .ZN(n4589) );
  AOI21_X1 U5166 ( .B1(n4590), .B2(n4596), .A(n4589), .ZN(n4591) );
  AND2_X1 U5167 ( .A1(n4592), .A2(n4591), .ZN(n4934) );
  MUX2_X1 U5168 ( .A(n4792), .B(n4934), .S(n5043), .Z(n4593) );
  OAI21_X1 U5169 ( .B1(n4594), .B2(n4937), .A(n4593), .ZN(U3530) );
  OR2_X1 U5170 ( .A1(n4596), .A2(n4595), .ZN(n4597) );
  NAND2_X1 U5171 ( .A1(n4598), .A2(n4597), .ZN(n4604) );
  AOI22_X1 U5172 ( .A1(n4602), .A2(n4601), .B1(n4600), .B2(n4599), .ZN(n4603)
         );
  NAND2_X1 U5173 ( .A1(n4604), .A2(n4603), .ZN(n5028) );
  MUX2_X1 U5174 ( .A(REG1_REG_0__SCAN_IN), .B(n5028), .S(n5043), .Z(n4870) );
  NOR4_X1 U5175 ( .A1(REG3_REG_18__SCAN_IN), .A2(REG1_REG_21__SCAN_IN), .A3(
        REG1_REG_16__SCAN_IN), .A4(REG0_REG_11__SCAN_IN), .ZN(n4614) );
  NOR4_X1 U5176 ( .A1(IR_REG_5__SCAN_IN), .A2(REG3_REG_9__SCAN_IN), .A3(
        REG3_REG_4__SCAN_IN), .A4(n2757), .ZN(n4613) );
  NAND4_X1 U5177 ( .A1(D_REG_17__SCAN_IN), .A2(D_REG_29__SCAN_IN), .A3(
        D_REG_14__SCAN_IN), .A4(D_REG_4__SCAN_IN), .ZN(n4611) );
  INV_X1 U5178 ( .A(REG1_REG_31__SCAN_IN), .ZN(n4669) );
  AND4_X1 U5179 ( .A1(ADDR_REG_5__SCAN_IN), .A2(ADDR_REG_1__SCAN_IN), .A3(
        n4686), .A4(n4691), .ZN(n4605) );
  NAND4_X1 U5180 ( .A1(n4606), .A2(n2629), .A3(n4669), .A4(n4605), .ZN(n4610)
         );
  NAND4_X1 U5181 ( .A1(n4607), .A2(IR_REG_28__SCAN_IN), .A3(
        REG1_REG_29__SCAN_IN), .A4(D_REG_13__SCAN_IN), .ZN(n4609) );
  INV_X1 U5182 ( .A(D_REG_9__SCAN_IN), .ZN(n4608) );
  NOR4_X1 U5183 ( .A1(n4611), .A2(n4610), .A3(n4609), .A4(n4608), .ZN(n4612)
         );
  NAND3_X1 U5184 ( .A1(n4614), .A2(n4613), .A3(n4612), .ZN(n4635) );
  NOR2_X1 U5185 ( .A1(D_REG_1__SCAN_IN), .A2(n2545), .ZN(n4616) );
  INV_X1 U5186 ( .A(D_REG_21__SCAN_IN), .ZN(n5005) );
  NOR4_X1 U5187 ( .A1(DATAO_REG_6__SCAN_IN), .A2(DATAO_REG_15__SCAN_IN), .A3(
        DATAO_REG_24__SCAN_IN), .A4(n5005), .ZN(n4615) );
  NAND4_X1 U5188 ( .A1(DATAI_13_), .A2(DATAO_REG_0__SCAN_IN), .A3(n4616), .A4(
        n4615), .ZN(n4634) );
  NOR4_X1 U5189 ( .A1(n4617), .A2(DATAI_7_), .A3(DATAI_4_), .A4(DATAI_6_), 
        .ZN(n4626) );
  INV_X1 U5190 ( .A(IR_REG_18__SCAN_IN), .ZN(n4763) );
  NOR4_X1 U5191 ( .A1(REG2_REG_11__SCAN_IN), .A2(REG2_REG_14__SCAN_IN), .A3(
        REG2_REG_7__SCAN_IN), .A4(n4763), .ZN(n4618) );
  NAND3_X1 U5192 ( .A1(REG2_REG_5__SCAN_IN), .A2(REG2_REG_13__SCAN_IN), .A3(
        n4618), .ZN(n4623) );
  AND4_X1 U5193 ( .A1(REG1_REG_23__SCAN_IN), .A2(n4668), .A3(n4659), .A4(n4896), .ZN(n4621) );
  AND4_X1 U5194 ( .A1(REG0_REG_25__SCAN_IN), .A2(REG1_REG_25__SCAN_IN), .A3(
        n4666), .A4(n4888), .ZN(n4620) );
  INV_X1 U5195 ( .A(DATAI_14_), .ZN(n4762) );
  INV_X1 U5196 ( .A(DATAI_12_), .ZN(n4761) );
  NOR4_X1 U5197 ( .A1(IR_REG_12__SCAN_IN), .A2(n4762), .A3(n4759), .A4(n4761), 
        .ZN(n4619) );
  NAND4_X1 U5198 ( .A1(REG1_REG_5__SCAN_IN), .A2(n4621), .A3(n4620), .A4(n4619), .ZN(n4622) );
  NOR4_X1 U5199 ( .A1(n4624), .A2(DATAO_REG_25__SCAN_IN), .A3(n4623), .A4(
        n4622), .ZN(n4625) );
  NAND4_X1 U5200 ( .A1(n4626), .A2(DATAI_1_), .A3(n4625), .A4(n4735), .ZN(
        n4631) );
  NAND4_X1 U5201 ( .A1(n4627), .A2(IR_REG_10__SCAN_IN), .A3(IR_REG_3__SCAN_IN), 
        .A4(IR_REG_4__SCAN_IN), .ZN(n4630) );
  NAND4_X1 U5202 ( .A1(n4628), .A2(n4792), .A3(IR_REG_27__SCAN_IN), .A4(
        DATAI_10_), .ZN(n4629) );
  OR4_X1 U5203 ( .A1(n4631), .A2(n4730), .A3(n4630), .A4(n4629), .ZN(n4633) );
  NOR4_X1 U5204 ( .A1(n4635), .A2(n4634), .A3(n4633), .A4(n4632), .ZN(n4642)
         );
  NOR4_X1 U5205 ( .A1(REG1_REG_9__SCAN_IN), .A2(REG1_REG_13__SCAN_IN), .A3(
        REG1_REG_2__SCAN_IN), .A4(n4840), .ZN(n4641) );
  NOR4_X1 U5206 ( .A1(DATAO_REG_14__SCAN_IN), .A2(ADDR_REG_14__SCAN_IN), .A3(
        DATAO_REG_21__SCAN_IN), .A4(n2561), .ZN(n4639) );
  NOR4_X1 U5207 ( .A1(REG3_REG_16__SCAN_IN), .A2(DATAO_REG_7__SCAN_IN), .A3(
        DATAO_REG_17__SCAN_IN), .A4(n4723), .ZN(n4638) );
  NOR4_X1 U5208 ( .A1(IR_REG_17__SCAN_IN), .A2(IR_REG_15__SCAN_IN), .A3(
        REG0_REG_15__SCAN_IN), .A4(n2458), .ZN(n4637) );
  INV_X1 U5209 ( .A(ADDR_REG_13__SCAN_IN), .ZN(n4720) );
  INV_X1 U5210 ( .A(ADDR_REG_3__SCAN_IN), .ZN(n4718) );
  NOR4_X1 U5211 ( .A1(REG3_REG_12__SCAN_IN), .A2(ADDR_REG_0__SCAN_IN), .A3(
        n4720), .A4(n4718), .ZN(n4636) );
  AND4_X1 U5212 ( .A1(n4639), .A2(n4638), .A3(n4637), .A4(n4636), .ZN(n4640)
         );
  NAND3_X1 U5213 ( .A1(n4642), .A2(n4641), .A3(n4640), .ZN(n4653) );
  NOR4_X1 U5214 ( .A1(REG2_REG_29__SCAN_IN), .A2(REG2_REG_27__SCAN_IN), .A3(
        n3377), .A4(n4820), .ZN(n4651) );
  NOR4_X1 U5215 ( .A1(ADDR_REG_9__SCAN_IN), .A2(ADDR_REG_7__SCAN_IN), .A3(
        ADDR_REG_10__SCAN_IN), .A4(n2747), .ZN(n4643) );
  NAND3_X1 U5216 ( .A1(ADDR_REG_17__SCAN_IN), .A2(ADDR_REG_16__SCAN_IN), .A3(
        n4643), .ZN(n4649) );
  INV_X1 U5217 ( .A(REG2_REG_26__SCAN_IN), .ZN(n4809) );
  NOR4_X1 U5218 ( .A1(REG2_REG_24__SCAN_IN), .A2(REG2_REG_22__SCAN_IN), .A3(
        n4809), .A4(n4811), .ZN(n4647) );
  NOR4_X1 U5219 ( .A1(REG3_REG_28__SCAN_IN), .A2(REG3_REG_26__SCAN_IN), .A3(
        REG3_REG_24__SCAN_IN), .A4(REG2_REG_31__SCAN_IN), .ZN(n4646) );
  INV_X1 U5220 ( .A(REG2_REG_4__SCAN_IN), .ZN(n4847) );
  NOR4_X1 U5221 ( .A1(REG1_REG_6__SCAN_IN), .A2(REG2_REG_6__SCAN_IN), .A3(
        ADDR_REG_2__SCAN_IN), .A4(n4847), .ZN(n4645) );
  NOR4_X1 U5222 ( .A1(DATAI_23_), .A2(n4850), .A3(n4813), .A4(n2814), .ZN(
        n4644) );
  NAND4_X1 U5223 ( .A1(n4647), .A2(n4646), .A3(n4645), .A4(n4644), .ZN(n4648)
         );
  NOR4_X1 U5224 ( .A1(REG3_REG_14__SCAN_IN), .A2(ADDR_REG_12__SCAN_IN), .A3(
        n4649), .A4(n4648), .ZN(n4650) );
  NAND4_X1 U5225 ( .A1(DATAI_16_), .A2(DATAO_REG_31__SCAN_IN), .A3(n4651), 
        .A4(n4650), .ZN(n4652) );
  OAI21_X1 U5226 ( .B1(n4653), .B2(n4652), .A(IR_REG_25__SCAN_IN), .ZN(n4868)
         );
  AOI22_X1 U5227 ( .A1(n2757), .A2(keyinput36), .B1(n3581), .B2(keyinput48), 
        .ZN(n4654) );
  OAI221_X1 U5228 ( .B1(n2757), .B2(keyinput36), .C1(n3581), .C2(keyinput48), 
        .A(n4654), .ZN(n4663) );
  AOI22_X1 U5229 ( .A1(n4656), .A2(keyinput87), .B1(n2296), .B2(keyinput80), 
        .ZN(n4655) );
  OAI221_X1 U5230 ( .B1(n4656), .B2(keyinput87), .C1(n2296), .C2(keyinput80), 
        .A(n4655), .ZN(n4662) );
  AOI22_X1 U5231 ( .A1(n4531), .A2(keyinput70), .B1(n4896), .B2(keyinput23), 
        .ZN(n4657) );
  OAI221_X1 U5232 ( .B1(n4531), .B2(keyinput70), .C1(n4896), .C2(keyinput23), 
        .A(n4657), .ZN(n4661) );
  AOI22_X1 U5233 ( .A1(n4659), .A2(keyinput52), .B1(n4517), .B2(keyinput24), 
        .ZN(n4658) );
  OAI221_X1 U5234 ( .B1(n4659), .B2(keyinput52), .C1(n4517), .C2(keyinput24), 
        .A(n4658), .ZN(n4660) );
  NOR4_X1 U5235 ( .A1(n4663), .A2(n4662), .A3(n4661), .A4(n4660), .ZN(n4702)
         );
  AOI22_X1 U5236 ( .A1(n4510), .A2(keyinput77), .B1(n3794), .B2(keyinput8), 
        .ZN(n4664) );
  OAI221_X1 U5237 ( .B1(n4510), .B2(keyinput77), .C1(n3794), .C2(keyinput8), 
        .A(n4664), .ZN(n4675) );
  AOI22_X1 U5238 ( .A1(n4666), .A2(keyinput58), .B1(n4884), .B2(keyinput78), 
        .ZN(n4665) );
  OAI221_X1 U5239 ( .B1(n4666), .B2(keyinput58), .C1(n4884), .C2(keyinput78), 
        .A(n4665), .ZN(n4674) );
  AOI22_X1 U5240 ( .A1(n4668), .A2(keyinput103), .B1(keyinput106), .B2(n4888), 
        .ZN(n4667) );
  OAI221_X1 U5241 ( .B1(n4668), .B2(keyinput103), .C1(n4888), .C2(keyinput106), 
        .A(n4667), .ZN(n4673) );
  XOR2_X1 U5242 ( .A(n4669), .B(keyinput11), .Z(n4671) );
  XNOR2_X1 U5243 ( .A(IR_REG_28__SCAN_IN), .B(keyinput59), .ZN(n4670) );
  NAND2_X1 U5244 ( .A1(n4671), .A2(n4670), .ZN(n4672) );
  NOR4_X1 U5245 ( .A1(n4675), .A2(n4674), .A3(n4673), .A4(n4672), .ZN(n4701)
         );
  INV_X1 U5246 ( .A(D_REG_13__SCAN_IN), .ZN(n5010) );
  INV_X1 U5247 ( .A(D_REG_17__SCAN_IN), .ZN(n5007) );
  AOI22_X1 U5248 ( .A1(n5010), .A2(keyinput43), .B1(keyinput72), .B2(n5007), 
        .ZN(n4676) );
  OAI221_X1 U5249 ( .B1(n5010), .B2(keyinput43), .C1(n5007), .C2(keyinput72), 
        .A(n4676), .ZN(n4684) );
  INV_X1 U5250 ( .A(D_REG_29__SCAN_IN), .ZN(n5002) );
  INV_X1 U5251 ( .A(D_REG_14__SCAN_IN), .ZN(n5009) );
  AOI22_X1 U5252 ( .A1(n5002), .A2(keyinput110), .B1(keyinput93), .B2(n5009), 
        .ZN(n4677) );
  OAI221_X1 U5253 ( .B1(n5002), .B2(keyinput110), .C1(n5009), .C2(keyinput93), 
        .A(n4677), .ZN(n4683) );
  XOR2_X1 U5254 ( .A(n2629), .B(keyinput1), .Z(n4681) );
  XOR2_X1 U5255 ( .A(n4608), .B(keyinput10), .Z(n4680) );
  XNOR2_X1 U5256 ( .A(REG0_REG_1__SCAN_IN), .B(keyinput31), .ZN(n4679) );
  XNOR2_X1 U5257 ( .A(IR_REG_22__SCAN_IN), .B(keyinput69), .ZN(n4678) );
  NAND4_X1 U5258 ( .A1(n4681), .A2(n4680), .A3(n4679), .A4(n4678), .ZN(n4682)
         );
  NOR3_X1 U5259 ( .A1(n4684), .A2(n4683), .A3(n4682), .ZN(n4700) );
  INV_X1 U5260 ( .A(D_REG_4__SCAN_IN), .ZN(n5014) );
  AOI22_X1 U5261 ( .A1(n5014), .A2(keyinput68), .B1(keyinput35), .B2(n4686), 
        .ZN(n4685) );
  OAI221_X1 U5262 ( .B1(n5014), .B2(keyinput68), .C1(n4686), .C2(keyinput35), 
        .A(n4685), .ZN(n4698) );
  INV_X1 U5263 ( .A(D_REG_11__SCAN_IN), .ZN(n5011) );
  INV_X1 U5264 ( .A(ADDR_REG_5__SCAN_IN), .ZN(n4688) );
  AOI22_X1 U5265 ( .A1(n5011), .A2(keyinput107), .B1(keyinput91), .B2(n4688), 
        .ZN(n4687) );
  OAI221_X1 U5266 ( .B1(n5011), .B2(keyinput107), .C1(n4688), .C2(keyinput91), 
        .A(n4687), .ZN(n4697) );
  INV_X1 U5267 ( .A(ADDR_REG_1__SCAN_IN), .ZN(n4690) );
  AOI22_X1 U5268 ( .A1(n4691), .A2(keyinput99), .B1(keyinput119), .B2(n4690), 
        .ZN(n4689) );
  OAI221_X1 U5269 ( .B1(n4691), .B2(keyinput99), .C1(n4690), .C2(keyinput119), 
        .A(n4689), .ZN(n4696) );
  INV_X1 U5270 ( .A(DATAI_13_), .ZN(n4693) );
  AOI22_X1 U5271 ( .A1(n4694), .A2(keyinput55), .B1(n4693), .B2(keyinput71), 
        .ZN(n4692) );
  OAI221_X1 U5272 ( .B1(n4694), .B2(keyinput55), .C1(n4693), .C2(keyinput71), 
        .A(n4692), .ZN(n4695) );
  NOR4_X1 U5273 ( .A1(n4698), .A2(n4697), .A3(n4696), .A4(n4695), .ZN(n4699)
         );
  NAND4_X1 U5274 ( .A1(n4702), .A2(n4701), .A3(n4700), .A4(n4699), .ZN(n4866)
         );
  AOI22_X1 U5275 ( .A1(n2978), .A2(keyinput22), .B1(n2545), .B2(keyinput38), 
        .ZN(n4703) );
  OAI221_X1 U5276 ( .B1(n2978), .B2(keyinput22), .C1(n2545), .C2(keyinput38), 
        .A(n4703), .ZN(n4712) );
  INV_X1 U5277 ( .A(D_REG_30__SCAN_IN), .ZN(n5001) );
  AOI22_X1 U5278 ( .A1(n5001), .A2(keyinput41), .B1(keyinput33), .B2(n5005), 
        .ZN(n4704) );
  OAI221_X1 U5279 ( .B1(n5001), .B2(keyinput41), .C1(n5005), .C2(keyinput33), 
        .A(n4704), .ZN(n4711) );
  AOI22_X1 U5280 ( .A1(n5015), .A2(keyinput34), .B1(keyinput6), .B2(n4706), 
        .ZN(n4705) );
  OAI221_X1 U5281 ( .B1(n5015), .B2(keyinput34), .C1(n4706), .C2(keyinput6), 
        .A(n4705), .ZN(n4710) );
  AOI22_X1 U5282 ( .A1(n5006), .A2(keyinput17), .B1(keyinput13), .B2(n4708), 
        .ZN(n4707) );
  OAI221_X1 U5283 ( .B1(n5006), .B2(keyinput17), .C1(n4708), .C2(keyinput13), 
        .A(n4707), .ZN(n4709) );
  NOR4_X1 U5284 ( .A1(n4712), .A2(n4711), .A3(n4710), .A4(n4709), .ZN(n4756)
         );
  AOI22_X1 U5285 ( .A1(n4715), .A2(keyinput124), .B1(n4714), .B2(keyinput126), 
        .ZN(n4713) );
  OAI221_X1 U5286 ( .B1(n4715), .B2(keyinput124), .C1(n4714), .C2(keyinput126), 
        .A(n4713), .ZN(n4727) );
  INV_X1 U5287 ( .A(ADDR_REG_0__SCAN_IN), .ZN(n4717) );
  AOI22_X1 U5288 ( .A1(n4718), .A2(keyinput116), .B1(keyinput114), .B2(n4717), 
        .ZN(n4716) );
  OAI221_X1 U5289 ( .B1(n4718), .B2(keyinput116), .C1(n4717), .C2(keyinput114), 
        .A(n4716), .ZN(n4726) );
  INV_X1 U5290 ( .A(D_REG_2__SCAN_IN), .ZN(n5016) );
  AOI22_X1 U5291 ( .A1(n4720), .A2(keyinput117), .B1(n5016), .B2(keyinput112), 
        .ZN(n4719) );
  OAI221_X1 U5292 ( .B1(n4720), .B2(keyinput117), .C1(n5016), .C2(keyinput112), 
        .A(n4719), .ZN(n4725) );
  AOI22_X1 U5293 ( .A1(n4723), .A2(keyinput105), .B1(keyinput104), .B2(n4722), 
        .ZN(n4721) );
  OAI221_X1 U5294 ( .B1(n4723), .B2(keyinput105), .C1(n4722), .C2(keyinput104), 
        .A(n4721), .ZN(n4724) );
  NOR4_X1 U5295 ( .A1(n4727), .A2(n4726), .A3(n4725), .A4(n4724), .ZN(n4755)
         );
  AOI22_X1 U5296 ( .A1(n4730), .A2(keyinput84), .B1(keyinput85), .B2(n4729), 
        .ZN(n4728) );
  OAI221_X1 U5297 ( .B1(n4730), .B2(keyinput84), .C1(n4729), .C2(keyinput85), 
        .A(n4728), .ZN(n4741) );
  INV_X1 U5298 ( .A(D_REG_27__SCAN_IN), .ZN(n5004) );
  AOI22_X1 U5299 ( .A1(n4732), .A2(keyinput90), .B1(n5004), .B2(keyinput88), 
        .ZN(n4731) );
  OAI221_X1 U5300 ( .B1(n4732), .B2(keyinput90), .C1(n5004), .C2(keyinput88), 
        .A(n4731), .ZN(n4740) );
  INV_X1 U5301 ( .A(D_REG_15__SCAN_IN), .ZN(n5008) );
  AOI22_X1 U5302 ( .A1(n5008), .A2(keyinput100), .B1(keyinput94), .B2(n4734), 
        .ZN(n4733) );
  OAI221_X1 U5303 ( .B1(n5008), .B2(keyinput100), .C1(n4734), .C2(keyinput94), 
        .A(n4733), .ZN(n4739) );
  XOR2_X1 U5304 ( .A(n4735), .B(keyinput81), .Z(n4737) );
  XNOR2_X1 U5305 ( .A(REG2_REG_0__SCAN_IN), .B(keyinput76), .ZN(n4736) );
  NAND2_X1 U5306 ( .A1(n4737), .A2(n4736), .ZN(n4738) );
  NOR4_X1 U5307 ( .A1(n4741), .A2(n4740), .A3(n4739), .A4(n4738), .ZN(n4754)
         );
  INV_X1 U5308 ( .A(D_REG_5__SCAN_IN), .ZN(n5013) );
  AOI22_X1 U5309 ( .A1(n5013), .A2(keyinput74), .B1(keyinput73), .B2(n4743), 
        .ZN(n4742) );
  OAI221_X1 U5310 ( .B1(n5013), .B2(keyinput74), .C1(n4743), .C2(keyinput73), 
        .A(n4742), .ZN(n4752) );
  INV_X1 U5311 ( .A(D_REG_28__SCAN_IN), .ZN(n5003) );
  AOI22_X1 U5312 ( .A1(n5003), .A2(keyinput66), .B1(keyinput65), .B2(n4745), 
        .ZN(n4744) );
  OAI221_X1 U5313 ( .B1(n5003), .B2(keyinput66), .C1(n4745), .C2(keyinput65), 
        .A(n4744), .ZN(n4751) );
  AOI22_X1 U5314 ( .A1(n4153), .A2(keyinput61), .B1(n2561), .B2(keyinput57), 
        .ZN(n4746) );
  OAI221_X1 U5315 ( .B1(n4153), .B2(keyinput61), .C1(n2561), .C2(keyinput57), 
        .A(n4746), .ZN(n4750) );
  INV_X1 U5316 ( .A(DATAI_16_), .ZN(n5023) );
  AOI22_X1 U5317 ( .A1(n4748), .A2(keyinput54), .B1(n5023), .B2(keyinput45), 
        .ZN(n4747) );
  OAI221_X1 U5318 ( .B1(n4748), .B2(keyinput54), .C1(n5023), .C2(keyinput45), 
        .A(n4747), .ZN(n4749) );
  NOR4_X1 U5319 ( .A1(n4752), .A2(n4751), .A3(n4750), .A4(n4749), .ZN(n4753)
         );
  NAND4_X1 U5320 ( .A1(n4756), .A2(n4755), .A3(n4754), .A4(n4753), .ZN(n4865)
         );
  AOI22_X1 U5321 ( .A1(n2460), .A2(keyinput44), .B1(keyinput56), .B2(n2458), 
        .ZN(n4757) );
  OAI221_X1 U5322 ( .B1(n2460), .B2(keyinput44), .C1(n2458), .C2(keyinput56), 
        .A(n4757), .ZN(n4769) );
  AOI22_X1 U5323 ( .A1(n4922), .A2(keyinput83), .B1(keyinput127), .B2(n4759), 
        .ZN(n4758) );
  OAI221_X1 U5324 ( .B1(n4922), .B2(keyinput83), .C1(n4759), .C2(keyinput127), 
        .A(n4758), .ZN(n4768) );
  AOI22_X1 U5325 ( .A1(n4762), .A2(keyinput14), .B1(keyinput20), .B2(n4761), 
        .ZN(n4760) );
  OAI221_X1 U5326 ( .B1(n4762), .B2(keyinput14), .C1(n4761), .C2(keyinput20), 
        .A(n4760), .ZN(n4767) );
  XOR2_X1 U5327 ( .A(n4763), .B(keyinput67), .Z(n4765) );
  XNOR2_X1 U5328 ( .A(IR_REG_17__SCAN_IN), .B(keyinput50), .ZN(n4764) );
  NAND2_X1 U5329 ( .A1(n4765), .A2(n4764), .ZN(n4766) );
  NOR4_X1 U5330 ( .A1(n4769), .A2(n4768), .A3(n4767), .A4(n4766), .ZN(n4807)
         );
  AOI22_X1 U5331 ( .A1(n2694), .A2(keyinput30), .B1(keyinput18), .B2(n2588), 
        .ZN(n4770) );
  OAI221_X1 U5332 ( .B1(n2694), .B2(keyinput30), .C1(n2588), .C2(keyinput18), 
        .A(n4770), .ZN(n4779) );
  AOI22_X1 U5333 ( .A1(n2596), .A2(keyinput96), .B1(n4772), .B2(keyinput25), 
        .ZN(n4771) );
  OAI221_X1 U5334 ( .B1(n2596), .B2(keyinput96), .C1(n4772), .C2(keyinput25), 
        .A(n4771), .ZN(n4778) );
  XNOR2_X1 U5335 ( .A(IR_REG_27__SCAN_IN), .B(keyinput46), .ZN(n4776) );
  XNOR2_X1 U5336 ( .A(REG1_REG_2__SCAN_IN), .B(keyinput39), .ZN(n4775) );
  XNOR2_X1 U5337 ( .A(keyinput64), .B(REG2_REG_13__SCAN_IN), .ZN(n4774) );
  XNOR2_X1 U5338 ( .A(keyinput79), .B(REG1_REG_5__SCAN_IN), .ZN(n4773) );
  NAND4_X1 U5339 ( .A1(n4776), .A2(n4775), .A3(n4774), .A4(n4773), .ZN(n4777)
         );
  NOR3_X1 U5340 ( .A1(n4779), .A2(n4778), .A3(n4777), .ZN(n4806) );
  AOI22_X1 U5341 ( .A1(n4781), .A2(keyinput5), .B1(keyinput51), .B2(n2737), 
        .ZN(n4780) );
  OAI221_X1 U5342 ( .B1(n4781), .B2(keyinput5), .C1(n2737), .C2(keyinput51), 
        .A(n4780), .ZN(n4790) );
  XNOR2_X1 U5343 ( .A(n4782), .B(keyinput37), .ZN(n4789) );
  XNOR2_X1 U5344 ( .A(keyinput82), .B(n2333), .ZN(n4788) );
  XNOR2_X1 U5345 ( .A(IR_REG_4__SCAN_IN), .B(keyinput115), .ZN(n4786) );
  XNOR2_X1 U5346 ( .A(DATAI_4_), .B(keyinput60), .ZN(n4785) );
  XNOR2_X1 U5347 ( .A(REG3_REG_4__SCAN_IN), .B(keyinput125), .ZN(n4784) );
  XNOR2_X1 U5348 ( .A(IR_REG_6__SCAN_IN), .B(keyinput121), .ZN(n4783) );
  NAND4_X1 U5349 ( .A1(n4786), .A2(n4785), .A3(n4784), .A4(n4783), .ZN(n4787)
         );
  NOR4_X1 U5350 ( .A1(n4790), .A2(n4789), .A3(n4788), .A4(n4787), .ZN(n4805)
         );
  INV_X1 U5351 ( .A(IR_REG_12__SCAN_IN), .ZN(n4793) );
  AOI22_X1 U5352 ( .A1(n4793), .A2(keyinput21), .B1(keyinput7), .B2(n4792), 
        .ZN(n4791) );
  OAI221_X1 U5353 ( .B1(n4793), .B2(keyinput21), .C1(n4792), .C2(keyinput7), 
        .A(n4791), .ZN(n4803) );
  XNOR2_X1 U5354 ( .A(n4794), .B(keyinput49), .ZN(n4802) );
  XNOR2_X1 U5355 ( .A(IR_REG_13__SCAN_IN), .B(keyinput122), .ZN(n4798) );
  XNOR2_X1 U5356 ( .A(DATAI_10_), .B(keyinput26), .ZN(n4797) );
  XNOR2_X1 U5357 ( .A(REG3_REG_7__SCAN_IN), .B(keyinput101), .ZN(n4796) );
  XNOR2_X1 U5358 ( .A(DATAI_6_), .B(keyinput89), .ZN(n4795) );
  NAND4_X1 U5359 ( .A1(n4798), .A2(n4797), .A3(n4796), .A4(n4795), .ZN(n4801)
         );
  INV_X1 U5360 ( .A(DATAI_7_), .ZN(n4799) );
  XNOR2_X1 U5361 ( .A(keyinput108), .B(n4799), .ZN(n4800) );
  NOR4_X1 U5362 ( .A1(n4803), .A2(n4802), .A3(n4801), .A4(n4800), .ZN(n4804)
         );
  NAND4_X1 U5363 ( .A1(n4807), .A2(n4806), .A3(n4805), .A4(n4804), .ZN(n4864)
         );
  AOI22_X1 U5364 ( .A1(n4809), .A2(keyinput3), .B1(keyinput53), .B2(n2857), 
        .ZN(n4808) );
  OAI221_X1 U5365 ( .B1(n4809), .B2(keyinput3), .C1(n2857), .C2(keyinput53), 
        .A(n4808), .ZN(n4818) );
  AOI22_X1 U5366 ( .A1(n3028), .A2(keyinput16), .B1(n4811), .B2(keyinput62), 
        .ZN(n4810) );
  OAI221_X1 U5367 ( .B1(n3028), .B2(keyinput16), .C1(n4811), .C2(keyinput62), 
        .A(n4810), .ZN(n4817) );
  AOI22_X1 U5368 ( .A1(n4813), .A2(keyinput4), .B1(keyinput118), .B2(n2814), 
        .ZN(n4812) );
  OAI221_X1 U5369 ( .B1(n4813), .B2(keyinput4), .C1(n2814), .C2(keyinput118), 
        .A(n4812), .ZN(n4816) );
  INV_X1 U5370 ( .A(DATAI_23_), .ZN(n5019) );
  AOI22_X1 U5371 ( .A1(n2638), .A2(keyinput0), .B1(n5019), .B2(keyinput12), 
        .ZN(n4814) );
  OAI221_X1 U5372 ( .B1(n2638), .B2(keyinput0), .C1(n5019), .C2(keyinput12), 
        .A(n4814), .ZN(n4815) );
  NOR4_X1 U5373 ( .A1(n4818), .A2(n4817), .A3(n4816), .A4(n4815), .ZN(n4862)
         );
  AOI22_X1 U5374 ( .A1(n4184), .A2(keyinput15), .B1(keyinput97), .B2(n4820), 
        .ZN(n4819) );
  OAI221_X1 U5375 ( .B1(n4184), .B2(keyinput15), .C1(n4820), .C2(keyinput97), 
        .A(n4819), .ZN(n4831) );
  AOI22_X1 U5376 ( .A1(n2887), .A2(keyinput120), .B1(keyinput9), .B2(n4822), 
        .ZN(n4821) );
  OAI221_X1 U5377 ( .B1(n2887), .B2(keyinput120), .C1(n4822), .C2(keyinput9), 
        .A(n4821), .ZN(n4830) );
  AOI22_X1 U5378 ( .A1(n4178), .A2(keyinput86), .B1(keyinput75), .B2(n4824), 
        .ZN(n4823) );
  OAI221_X1 U5379 ( .B1(n4178), .B2(keyinput86), .C1(n4824), .C2(keyinput75), 
        .A(n4823), .ZN(n4829) );
  INV_X1 U5380 ( .A(keyinput123), .ZN(n4825) );
  NAND2_X1 U5381 ( .A1(n4825), .A2(IR_REG_25__SCAN_IN), .ZN(n4827) );
  NAND2_X1 U5382 ( .A1(n3377), .A2(keyinput113), .ZN(n4826) );
  OAI211_X1 U5383 ( .C1(keyinput113), .C2(n3377), .A(n4827), .B(n4826), .ZN(
        n4828) );
  NOR4_X1 U5384 ( .A1(n4831), .A2(n4830), .A3(n4829), .A4(n4828), .ZN(n4861)
         );
  INV_X1 U5385 ( .A(ADDR_REG_16__SCAN_IN), .ZN(n4977) );
  AOI22_X1 U5386 ( .A1(n4833), .A2(keyinput29), .B1(keyinput28), .B2(n4977), 
        .ZN(n4832) );
  OAI221_X1 U5387 ( .B1(n4833), .B2(keyinput29), .C1(n4977), .C2(keyinput28), 
        .A(n4832), .ZN(n4845) );
  INV_X1 U5388 ( .A(ADDR_REG_12__SCAN_IN), .ZN(n4835) );
  AOI22_X1 U5389 ( .A1(n4836), .A2(keyinput111), .B1(n4835), .B2(keyinput42), 
        .ZN(n4834) );
  OAI221_X1 U5390 ( .B1(n4836), .B2(keyinput111), .C1(n4835), .C2(keyinput42), 
        .A(n4834), .ZN(n4844) );
  AOI22_X1 U5391 ( .A1(n4580), .A2(keyinput32), .B1(keyinput27), .B2(n4838), 
        .ZN(n4837) );
  OAI221_X1 U5392 ( .B1(n4580), .B2(keyinput32), .C1(n4838), .C2(keyinput27), 
        .A(n4837), .ZN(n4843) );
  INV_X1 U5393 ( .A(ADDR_REG_17__SCAN_IN), .ZN(n4841) );
  AOI22_X1 U5394 ( .A1(n4841), .A2(keyinput63), .B1(n4840), .B2(keyinput98), 
        .ZN(n4839) );
  OAI221_X1 U5395 ( .B1(n4841), .B2(keyinput63), .C1(n4840), .C2(keyinput98), 
        .A(n4839), .ZN(n4842) );
  NOR4_X1 U5396 ( .A1(n4845), .A2(n4844), .A3(n4843), .A4(n4842), .ZN(n4860)
         );
  AOI22_X1 U5397 ( .A1(n4847), .A2(keyinput19), .B1(n3409), .B2(keyinput102), 
        .ZN(n4846) );
  OAI221_X1 U5398 ( .B1(n4847), .B2(keyinput19), .C1(n3409), .C2(keyinput102), 
        .A(n4846), .ZN(n4858) );
  INV_X1 U5399 ( .A(ADDR_REG_2__SCAN_IN), .ZN(n4849) );
  AOI22_X1 U5400 ( .A1(n4850), .A2(keyinput2), .B1(keyinput92), .B2(n4849), 
        .ZN(n4848) );
  OAI221_X1 U5401 ( .B1(n4850), .B2(keyinput2), .C1(n4849), .C2(keyinput92), 
        .A(n4848), .ZN(n4857) );
  AOI22_X1 U5402 ( .A1(n4852), .A2(keyinput109), .B1(n2747), .B2(keyinput47), 
        .ZN(n4851) );
  OAI221_X1 U5403 ( .B1(n4852), .B2(keyinput109), .C1(n2747), .C2(keyinput47), 
        .A(n4851), .ZN(n4856) );
  AOI22_X1 U5404 ( .A1(n2715), .A2(keyinput40), .B1(keyinput95), .B2(n4854), 
        .ZN(n4853) );
  OAI221_X1 U5405 ( .B1(n2715), .B2(keyinput40), .C1(n4854), .C2(keyinput95), 
        .A(n4853), .ZN(n4855) );
  NOR4_X1 U5406 ( .A1(n4858), .A2(n4857), .A3(n4856), .A4(n4855), .ZN(n4859)
         );
  NAND4_X1 U5407 ( .A1(n4862), .A2(n4861), .A3(n4860), .A4(n4859), .ZN(n4863)
         );
  OR4_X1 U5408 ( .A1(n4866), .A2(n4865), .A3(n4864), .A4(n4863), .ZN(n4867) );
  AOI21_X1 U5409 ( .B1(keyinput123), .B2(n4868), .A(n4867), .ZN(n4869) );
  XOR2_X1 U5410 ( .A(n4870), .B(n4869), .Z(U3518) );
  NAND2_X1 U5411 ( .A1(n5040), .A2(n4871), .ZN(n4873) );
  NAND2_X1 U5412 ( .A1(n5039), .A2(REG0_REG_30__SCAN_IN), .ZN(n4872) );
  OAI211_X1 U5413 ( .C1(n4874), .C2(n4936), .A(n4873), .B(n4872), .ZN(U3516)
         );
  INV_X1 U5414 ( .A(REG0_REG_27__SCAN_IN), .ZN(n4876) );
  MUX2_X1 U5415 ( .A(n4876), .B(n4875), .S(n5040), .Z(n4877) );
  OAI21_X1 U5416 ( .B1(n4878), .B2(n4936), .A(n4877), .ZN(U3513) );
  INV_X1 U5417 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4880) );
  MUX2_X1 U5418 ( .A(n4880), .B(n4879), .S(n5040), .Z(n4881) );
  OAI21_X1 U5419 ( .B1(n4882), .B2(n4936), .A(n4881), .ZN(U3512) );
  MUX2_X1 U5420 ( .A(n4884), .B(n4883), .S(n5040), .Z(n4885) );
  OAI21_X1 U5421 ( .B1(n4886), .B2(n4936), .A(n4885), .ZN(U3511) );
  MUX2_X1 U5422 ( .A(n4888), .B(n4887), .S(n5040), .Z(n4889) );
  OAI21_X1 U5423 ( .B1(n4890), .B2(n4936), .A(n4889), .ZN(U3510) );
  INV_X1 U5424 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4892) );
  MUX2_X1 U5425 ( .A(n4892), .B(n4891), .S(n5040), .Z(n4893) );
  OAI21_X1 U5426 ( .B1(n4894), .B2(n4936), .A(n4893), .ZN(U3509) );
  MUX2_X1 U5427 ( .A(n4896), .B(n4895), .S(n5040), .Z(n4897) );
  OAI21_X1 U5428 ( .B1(n4898), .B2(n4936), .A(n4897), .ZN(U3508) );
  INV_X1 U5429 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4900) );
  MUX2_X1 U5430 ( .A(n4900), .B(n4899), .S(n5040), .Z(n4901) );
  OAI21_X1 U5431 ( .B1(n4902), .B2(n4936), .A(n4901), .ZN(U3507) );
  MUX2_X1 U5432 ( .A(n4904), .B(n4903), .S(n5040), .Z(n4905) );
  OAI21_X1 U5433 ( .B1(n4906), .B2(n4936), .A(n4905), .ZN(U3506) );
  INV_X1 U5434 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4908) );
  MUX2_X1 U5435 ( .A(n4908), .B(n4907), .S(n5040), .Z(n4909) );
  OAI21_X1 U5436 ( .B1(n4910), .B2(n4936), .A(n4909), .ZN(U3505) );
  MUX2_X1 U5437 ( .A(REG0_REG_18__SCAN_IN), .B(n4911), .S(n5040), .Z(U3503) );
  MUX2_X1 U5438 ( .A(REG0_REG_17__SCAN_IN), .B(n4912), .S(n5040), .Z(n4913) );
  INV_X1 U5439 ( .A(n4913), .ZN(n4914) );
  OAI21_X1 U5440 ( .B1(n4915), .B2(n4936), .A(n4914), .ZN(U3501) );
  MUX2_X1 U5441 ( .A(n4916), .B(REG0_REG_16__SCAN_IN), .S(n5039), .Z(n4917) );
  AOI21_X1 U5442 ( .B1(n4919), .B2(n4918), .A(n4917), .ZN(n4920) );
  INV_X1 U5443 ( .A(n4920), .ZN(U3499) );
  MUX2_X1 U5444 ( .A(n4922), .B(n4921), .S(n5040), .Z(n4923) );
  OAI21_X1 U5445 ( .B1(n4924), .B2(n4936), .A(n4923), .ZN(U3497) );
  INV_X1 U5446 ( .A(REG0_REG_14__SCAN_IN), .ZN(n4926) );
  MUX2_X1 U5447 ( .A(n4926), .B(n4925), .S(n5040), .Z(n4927) );
  OAI21_X1 U5448 ( .B1(n4928), .B2(n4936), .A(n4927), .ZN(U3495) );
  INV_X1 U5449 ( .A(REG0_REG_13__SCAN_IN), .ZN(n4930) );
  MUX2_X1 U5450 ( .A(n4930), .B(n4929), .S(n5040), .Z(n4931) );
  OAI21_X1 U5451 ( .B1(n4932), .B2(n4936), .A(n4931), .ZN(U3493) );
  MUX2_X1 U5452 ( .A(n4934), .B(n4933), .S(n5039), .Z(n4935) );
  OAI21_X1 U5453 ( .B1(n4937), .B2(n4936), .A(n4935), .ZN(U3491) );
  MUX2_X1 U5454 ( .A(n4950), .B(DATAI_27_), .S(U3149), .Z(U3325) );
  MUX2_X1 U5455 ( .A(n4938), .B(DATAI_14_), .S(U3149), .Z(U3338) );
  MUX2_X1 U5456 ( .A(n4939), .B(DATAI_13_), .S(U3149), .Z(U3339) );
  MUX2_X1 U5457 ( .A(DATAI_12_), .B(n4940), .S(STATE_REG_SCAN_IN), .Z(U3340)
         );
  MUX2_X1 U5458 ( .A(n4941), .B(DATAI_7_), .S(U3149), .Z(U3345) );
  MUX2_X1 U5459 ( .A(DATAI_6_), .B(n4942), .S(STATE_REG_SCAN_IN), .Z(U3346) );
  MUX2_X1 U5460 ( .A(DATAI_4_), .B(n4943), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U5461 ( .A(DATAI_2_), .B(n4944), .S(STATE_REG_SCAN_IN), .Z(U3350) );
  MUX2_X1 U5462 ( .A(n4945), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  INV_X1 U5463 ( .A(DATAI_28_), .ZN(n4946) );
  AOI22_X1 U5464 ( .A1(STATE_REG_SCAN_IN), .A2(n4947), .B1(n4946), .B2(U3149), 
        .ZN(U3324) );
  INV_X1 U5465 ( .A(n4948), .ZN(n4949) );
  OAI21_X1 U5466 ( .B1(REG1_REG_0__SCAN_IN), .B2(n4950), .A(n4949), .ZN(n4951)
         );
  XOR2_X1 U5467 ( .A(n4951), .B(IR_REG_0__SCAN_IN), .Z(n4954) );
  AOI22_X1 U5468 ( .A1(ADDR_REG_0__SCAN_IN), .A2(n4994), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n4952) );
  OAI21_X1 U5469 ( .B1(n4954), .B2(n4953), .A(n4952), .ZN(U3240) );
  AOI211_X1 U5470 ( .C1(n4957), .C2(n4956), .A(n4955), .B(n4989), .ZN(n4958)
         );
  AOI211_X1 U5471 ( .C1(n4994), .C2(ADDR_REG_15__SCAN_IN), .A(n4959), .B(n4958), .ZN(n4964) );
  OAI211_X1 U5472 ( .C1(n4962), .C2(n4961), .A(n4996), .B(n4960), .ZN(n4963)
         );
  OAI211_X1 U5473 ( .C1(n5000), .C2(n5026), .A(n4964), .B(n4963), .ZN(U3255)
         );
  OAI21_X1 U5474 ( .B1(n4967), .B2(n4966), .A(n4965), .ZN(n4973) );
  AOI21_X1 U5475 ( .B1(REG1_REG_16__SCAN_IN), .B2(n4969), .A(n4968), .ZN(n4971) );
  OAI22_X1 U5476 ( .A1(n4971), .A2(n4970), .B1(n5024), .B2(n5000), .ZN(n4972)
         );
  AOI21_X1 U5477 ( .B1(n4974), .B2(n4973), .A(n4972), .ZN(n4976) );
  OAI211_X1 U5478 ( .C1(n4978), .C2(n4977), .A(n4976), .B(n4975), .ZN(U3256)
         );
  AOI221_X1 U5479 ( .B1(n4981), .B2(n4980), .C1(n4979), .C2(n4980), .A(n4989), 
        .ZN(n4982) );
  AOI211_X1 U5480 ( .C1(n4994), .C2(ADDR_REG_17__SCAN_IN), .A(n4983), .B(n4982), .ZN(n4988) );
  OAI221_X1 U5481 ( .B1(n4986), .B2(n4985), .C1(n4986), .C2(n4984), .A(n4996), 
        .ZN(n4987) );
  OAI211_X1 U5482 ( .C1(n5000), .C2(n5022), .A(n4988), .B(n4987), .ZN(U3257)
         );
  OAI211_X1 U5483 ( .C1(n4998), .C2(n4997), .A(n4996), .B(n4995), .ZN(n4999)
         );
  AND2_X1 U5484 ( .A1(D_REG_31__SCAN_IN), .A2(n5012), .ZN(U3291) );
  NOR2_X1 U5485 ( .A1(n5017), .A2(n5001), .ZN(U3292) );
  NOR2_X1 U5486 ( .A1(n5017), .A2(n5002), .ZN(U3293) );
  NOR2_X1 U5487 ( .A1(n5017), .A2(n5003), .ZN(U3294) );
  NOR2_X1 U5488 ( .A1(n5017), .A2(n5004), .ZN(U3295) );
  AND2_X1 U5489 ( .A1(D_REG_26__SCAN_IN), .A2(n5012), .ZN(U3296) );
  AND2_X1 U5490 ( .A1(D_REG_25__SCAN_IN), .A2(n5012), .ZN(U3297) );
  AND2_X1 U5491 ( .A1(D_REG_24__SCAN_IN), .A2(n5012), .ZN(U3298) );
  AND2_X1 U5492 ( .A1(D_REG_23__SCAN_IN), .A2(n5012), .ZN(U3299) );
  AND2_X1 U5493 ( .A1(D_REG_22__SCAN_IN), .A2(n5012), .ZN(U3300) );
  NOR2_X1 U5494 ( .A1(n5017), .A2(n5005), .ZN(U3301) );
  AND2_X1 U5495 ( .A1(D_REG_20__SCAN_IN), .A2(n5012), .ZN(U3302) );
  NOR2_X1 U5496 ( .A1(n5017), .A2(n5006), .ZN(U3303) );
  AND2_X1 U5497 ( .A1(D_REG_18__SCAN_IN), .A2(n5012), .ZN(U3304) );
  NOR2_X1 U5498 ( .A1(n5017), .A2(n5007), .ZN(U3305) );
  AND2_X1 U5499 ( .A1(D_REG_16__SCAN_IN), .A2(n5012), .ZN(U3306) );
  NOR2_X1 U5500 ( .A1(n5017), .A2(n5008), .ZN(U3307) );
  NOR2_X1 U5501 ( .A1(n5017), .A2(n5009), .ZN(U3308) );
  NOR2_X1 U5502 ( .A1(n5017), .A2(n5010), .ZN(U3309) );
  AND2_X1 U5503 ( .A1(D_REG_12__SCAN_IN), .A2(n5012), .ZN(U3310) );
  NOR2_X1 U5504 ( .A1(n5017), .A2(n5011), .ZN(U3311) );
  AND2_X1 U5505 ( .A1(D_REG_10__SCAN_IN), .A2(n5012), .ZN(U3312) );
  NOR2_X1 U5506 ( .A1(n5017), .A2(n4608), .ZN(U3313) );
  AND2_X1 U5507 ( .A1(D_REG_8__SCAN_IN), .A2(n5012), .ZN(U3314) );
  AND2_X1 U5508 ( .A1(D_REG_7__SCAN_IN), .A2(n5012), .ZN(U3315) );
  AND2_X1 U5509 ( .A1(D_REG_6__SCAN_IN), .A2(n5012), .ZN(U3316) );
  NOR2_X1 U5510 ( .A1(n5017), .A2(n5013), .ZN(U3317) );
  NOR2_X1 U5511 ( .A1(n5017), .A2(n5014), .ZN(U3318) );
  NOR2_X1 U5512 ( .A1(n5017), .A2(n5015), .ZN(U3319) );
  NOR2_X1 U5513 ( .A1(n5017), .A2(n5016), .ZN(U3320) );
  AOI21_X1 U5514 ( .B1(U3149), .B2(n5019), .A(n5018), .ZN(U3329) );
  INV_X1 U5515 ( .A(DATAI_18_), .ZN(n5020) );
  AOI22_X1 U5516 ( .A1(STATE_REG_SCAN_IN), .A2(n5021), .B1(n5020), .B2(U3149), 
        .ZN(U3334) );
  AOI22_X1 U5517 ( .A1(STATE_REG_SCAN_IN), .A2(n5022), .B1(n2814), .B2(U3149), 
        .ZN(U3335) );
  AOI22_X1 U5518 ( .A1(STATE_REG_SCAN_IN), .A2(n5024), .B1(n5023), .B2(U3149), 
        .ZN(U3336) );
  INV_X1 U5519 ( .A(DATAI_15_), .ZN(n5025) );
  AOI22_X1 U5520 ( .A1(STATE_REG_SCAN_IN), .A2(n5026), .B1(n5025), .B2(U3149), 
        .ZN(U3337) );
  INV_X1 U5521 ( .A(DATAI_0_), .ZN(n5027) );
  AOI22_X1 U5522 ( .A1(STATE_REG_SCAN_IN), .A2(n2323), .B1(n5027), .B2(U3149), 
        .ZN(U3352) );
  MUX2_X1 U5523 ( .A(REG0_REG_0__SCAN_IN), .B(n5028), .S(n5040), .Z(U3467) );
  AOI211_X1 U5524 ( .C1(n5037), .C2(n5031), .A(n5030), .B(n5029), .ZN(n5041)
         );
  AOI22_X1 U5525 ( .A1(n5040), .A2(n5041), .B1(n2674), .B2(n5039), .ZN(U3475)
         );
  NOR3_X1 U5526 ( .A1(n5034), .A2(n5033), .A3(n5032), .ZN(n5036) );
  AOI211_X1 U5527 ( .C1(n5038), .C2(n5037), .A(n5036), .B(n5035), .ZN(n5042)
         );
  AOI22_X1 U5528 ( .A1(n5040), .A2(n5042), .B1(n2719), .B2(n5039), .ZN(U3479)
         );
  AOI22_X1 U5529 ( .A1(n5043), .A2(n5041), .B1(n3116), .B2(n2210), .ZN(U3522)
         );
  AOI22_X1 U5530 ( .A1(n5043), .A2(n5042), .B1(n2715), .B2(n2210), .ZN(U3524)
         );
  CLKBUF_X1 U2393 ( .A(n2659), .Z(n3036) );
  CLKBUF_X1 U2500 ( .A(n2672), .Z(n3040) );
  CLKBUF_X1 U2501 ( .A(n2708), .Z(n2142) );
endmodule

