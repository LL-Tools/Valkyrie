

module b14_C_gen_AntiSAT_k_256_9 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, keyinput_f0, keyinput_f1, 
        keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, 
        keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, 
        keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, 
        keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, 
        keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, 
        keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, 
        keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, 
        keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, 
        keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, 
        keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, 
        keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, 
        keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, 
        keyinput_f62, keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66, 
        keyinput_f67, keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71, 
        keyinput_f72, keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76, 
        keyinput_f77, keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81, 
        keyinput_f82, keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86, 
        keyinput_f87, keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91, 
        keyinput_f92, keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96, 
        keyinput_f97, keyinput_f98, keyinput_f99, keyinput_f100, keyinput_f101, 
        keyinput_f102, keyinput_f103, keyinput_f104, keyinput_f105, 
        keyinput_f106, keyinput_f107, keyinput_f108, keyinput_f109, 
        keyinput_f110, keyinput_f111, keyinput_f112, keyinput_f113, 
        keyinput_f114, keyinput_f115, keyinput_f116, keyinput_f117, 
        keyinput_f118, keyinput_f119, keyinput_f120, keyinput_f121, 
        keyinput_f122, keyinput_f123, keyinput_f124, keyinput_f125, 
        keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, keyinput_g2, 
        keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, 
        keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, 
        keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, 
        keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, 
        keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, 
        keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, 
        keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, 
        keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, 
        keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, 
        keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, 
        keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, 
        keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, 
        keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, keyinput_g67, 
        keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, keyinput_g72, 
        keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, keyinput_g77, 
        keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, keyinput_g82, 
        keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, keyinput_g87, 
        keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, keyinput_g92, 
        keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, keyinput_g97, 
        keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101, 
        keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105, 
        keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109, 
        keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113, 
        keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117, 
        keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121, 
        keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125, 
        keyinput_g126, keyinput_g127, U3352, U3351, U3350, U3349, U3348, U3347, 
        U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, U3338, U3337, 
        U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, U3328, U3327, 
        U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, U3320, U3319, 
        U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, U3310, U3309, 
        U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, U3300, U3299, 
        U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, U3467, U3469, 
        U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, U3487, U3489, 
        U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, U3506, U3507, 
        U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, U3516, U3517, 
        U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, U3526, U3527, 
        U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, U3536, U3537, 
        U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, U3546, U3547, 
        U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, U3284, U3283, 
        U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, U3274, U3273, 
        U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, U3264, U3263, 
        U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, U3255, U3254, 
        U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, U3245, U3244, 
        U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, U3554, U3555, 
        U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, U3564, U3565, 
        U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, U3574, U3575, 
        U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, U3237, U3236, 
        U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, U3227, U3226, 
        U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, U3217, U3216, 
        U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, U4043 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66, keyinput_f67,
         keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71, keyinput_f72,
         keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76, keyinput_f77,
         keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81, keyinput_f82,
         keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86, keyinput_f87,
         keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91, keyinput_f92,
         keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96, keyinput_f97,
         keyinput_f98, keyinput_f99, keyinput_f100, keyinput_f101,
         keyinput_f102, keyinput_f103, keyinput_f104, keyinput_f105,
         keyinput_f106, keyinput_f107, keyinput_f108, keyinput_f109,
         keyinput_f110, keyinput_f111, keyinput_f112, keyinput_f113,
         keyinput_f114, keyinput_f115, keyinput_f116, keyinput_f117,
         keyinput_f118, keyinput_f119, keyinput_f120, keyinput_f121,
         keyinput_f122, keyinput_f123, keyinput_f124, keyinput_f125,
         keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, keyinput_g2,
         keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7,
         keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12,
         keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17,
         keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22,
         keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27,
         keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32,
         keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37,
         keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42,
         keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47,
         keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52,
         keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57,
         keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62,
         keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, keyinput_g67,
         keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, keyinput_g72,
         keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, keyinput_g77,
         keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, keyinput_g82,
         keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, keyinput_g87,
         keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, keyinput_g92,
         keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, keyinput_g97,
         keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101,
         keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105,
         keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109,
         keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113,
         keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117,
         keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121,
         keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125,
         keyinput_g126, keyinput_g127;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2232, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503,
         n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513,
         n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523,
         n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533,
         n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543,
         n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
         n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563,
         n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573,
         n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
         n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
         n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603,
         n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613,
         n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623,
         n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633,
         n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643,
         n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653,
         n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663,
         n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673,
         n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683,
         n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693,
         n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703,
         n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713,
         n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723,
         n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733,
         n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743,
         n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753,
         n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763,
         n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773,
         n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783,
         n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793,
         n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803,
         n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813,
         n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823,
         n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833,
         n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843,
         n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853,
         n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863,
         n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873,
         n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883,
         n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893,
         n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903,
         n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913,
         n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923,
         n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933,
         n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943,
         n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953,
         n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963,
         n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973,
         n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983,
         n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993,
         n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003,
         n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013,
         n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023,
         n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033,
         n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043,
         n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053,
         n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063,
         n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073,
         n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083,
         n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093,
         n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103,
         n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113,
         n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123,
         n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133,
         n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143,
         n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153,
         n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163,
         n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173,
         n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183,
         n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193,
         n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203,
         n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213,
         n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223,
         n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233,
         n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243,
         n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253,
         n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263,
         n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273,
         n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283,
         n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293,
         n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303,
         n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313,
         n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323,
         n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333,
         n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
         n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353,
         n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363,
         n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373,
         n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383,
         n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393,
         n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403,
         n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413,
         n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423,
         n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433,
         n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443,
         n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453,
         n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463,
         n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473,
         n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483,
         n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493,
         n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503,
         n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513,
         n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523,
         n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533,
         n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543,
         n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553,
         n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563,
         n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
         n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
         n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593,
         n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
         n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
         n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
         n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
         n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
         n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
         n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
         n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
         n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
         n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
         n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
         n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713,
         n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723,
         n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733,
         n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743,
         n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753,
         n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763,
         n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773,
         n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783,
         n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793,
         n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803,
         n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813,
         n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823,
         n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833,
         n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843,
         n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853,
         n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863,
         n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873,
         n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883,
         n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893,
         n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903,
         n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913,
         n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923,
         n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933,
         n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943,
         n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953,
         n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963,
         n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973,
         n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3983, n3984,
         n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
         n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004,
         n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014,
         n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024,
         n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034,
         n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044,
         n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
         n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
         n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
         n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084,
         n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094,
         n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104,
         n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114,
         n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124,
         n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134,
         n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144,
         n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
         n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164,
         n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
         n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184,
         n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194,
         n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204,
         n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214,
         n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224,
         n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234,
         n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244,
         n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254,
         n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264,
         n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
         n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
         n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
         n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
         n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097;

  INV_X1 U2474 ( .A(n3675), .ZN(n3661) );
  AND2_X1 U2477 ( .A1(n2505), .A2(n2504), .ZN(n2741) );
  NAND2_X1 U2478 ( .A1(n2869), .A2(IR_REG_31__SCAN_IN), .ZN(n2861) );
  INV_X1 U2479 ( .A(IR_REG_31__SCAN_IN), .ZN(n2863) );
  AOI211_X1 U2480 ( .C1(n4101), .C2(n4100), .A(n2257), .B(n4630), .ZN(n4102)
         );
  INV_X1 U2481 ( .A(n3197), .ZN(n3191) );
  OAI22_X2 U2482 ( .A1(n4091), .A2(n4090), .B1(n4521), .B2(
        REG2_REG_13__SCAN_IN), .ZN(n4092) );
  NOR2_X2 U2483 ( .A1(IR_REG_5__SCAN_IN), .A2(IR_REG_9__SCAN_IN), .ZN(n2669)
         );
  NAND2_X1 U2484 ( .A1(n2924), .A2(n2923), .ZN(n3675) );
  AND2_X4 U2485 ( .A1(n4517), .A2(n2516), .ZN(n2537) );
  XNOR2_X2 U2486 ( .A(n2861), .B(IR_REG_24__SCAN_IN), .ZN(n2868) );
  NOR2_X1 U2487 ( .A1(n4603), .A2(n4094), .ZN(n4613) );
  NOR2_X1 U2488 ( .A1(n4604), .A2(n3437), .ZN(n4603) );
  NAND2_X1 U2489 ( .A1(n3237), .A2(n3236), .ZN(n3235) );
  NAND2_X1 U2490 ( .A1(n4052), .A2(REG2_REG_12__SCAN_IN), .ZN(n4059) );
  AND4_X1 U2491 ( .A1(n2531), .A2(n2532), .A3(n2533), .A4(n2530), .ZN(n2928)
         );
  AND2_X2 U2492 ( .A1(n3031), .A2(n4517), .ZN(n2529) );
  AOI211_X1 U2493 ( .C1(n3800), .C2(n4554), .A(n3799), .B(n3798), .ZN(n3801)
         );
  AOI21_X1 U2494 ( .B1(n3555), .B2(n3554), .A(n3553), .ZN(n3576) );
  NOR2_X1 U2495 ( .A1(n4182), .A2(n4166), .ZN(n4160) );
  AND2_X1 U2496 ( .A1(n2456), .A2(n2454), .ZN(n3522) );
  OR2_X1 U2497 ( .A1(n2816), .A2(n2301), .ZN(n2297) );
  AND2_X1 U2498 ( .A1(n4592), .A2(n2360), .ZN(n4060) );
  AND2_X1 U2499 ( .A1(n2457), .A2(n2455), .ZN(n2454) );
  OR2_X1 U2500 ( .A1(n2347), .A2(n2236), .ZN(n2344) );
  OR2_X1 U2501 ( .A1(n3181), .A2(n2306), .ZN(n2305) );
  OR2_X1 U2502 ( .A1(n2459), .A2(n2246), .ZN(n2457) );
  AOI21_X1 U2503 ( .B1(n2469), .B2(n2473), .A(n2348), .ZN(n2347) );
  OAI22_X1 U2504 ( .A1(n4047), .A2(n4653), .B1(n4046), .B2(n2355), .ZN(n4573)
         );
  XNOR2_X1 U2505 ( .A(n2356), .B(n3161), .ZN(n4047) );
  AND2_X1 U2506 ( .A1(n2277), .A2(n2276), .ZN(n3192) );
  NAND2_X2 U2507 ( .A1(n2868), .A2(n2867), .ZN(n2921) );
  INV_X1 U2508 ( .A(n2923), .ZN(n3124) );
  AND4_X1 U2509 ( .A1(n2548), .A2(n2547), .A3(n2546), .A4(n2545), .ZN(n3228)
         );
  OAI21_X1 U2510 ( .B1(n2234), .B2(n2376), .A(n2375), .ZN(n3197) );
  NAND2_X1 U2511 ( .A1(n4518), .A2(n3963), .ZN(n2923) );
  INV_X1 U2512 ( .A(n3866), .ZN(n4518) );
  INV_X2 U2513 ( .A(n2536), .ZN(n2528) );
  NAND2_X1 U2514 ( .A1(n2799), .A2(n2804), .ZN(n3866) );
  MUX2_X1 U2515 ( .A(IR_REG_31__SCAN_IN), .B(n2797), .S(IR_REG_21__SCAN_IN), 
        .Z(n2799) );
  NAND2_X1 U2516 ( .A1(n2513), .A2(n2512), .ZN(n2515) );
  OR2_X1 U2517 ( .A1(n2859), .A2(n2858), .ZN(n3015) );
  OR2_X1 U2518 ( .A1(n3022), .A2(n2863), .ZN(n2514) );
  AND2_X1 U2519 ( .A1(n2475), .A2(n2437), .ZN(n3022) );
  NAND2_X1 U2520 ( .A1(n2507), .A2(IR_REG_31__SCAN_IN), .ZN(n2904) );
  AND2_X1 U2521 ( .A1(n2439), .A2(n2509), .ZN(n2438) );
  AND2_X1 U2522 ( .A1(n2484), .A2(n2477), .ZN(n2475) );
  AND2_X1 U2523 ( .A1(n4806), .A2(n2258), .ZN(n2439) );
  INV_X1 U2524 ( .A(IR_REG_6__SCAN_IN), .ZN(n4826) );
  NOR2_X1 U2525 ( .A1(IR_REG_0__SCAN_IN), .A2(IR_REG_1__SCAN_IN), .ZN(n2549)
         );
  NOR2_X1 U2526 ( .A1(IR_REG_3__SCAN_IN), .A2(IR_REG_4__SCAN_IN), .ZN(n2493)
         );
  INV_X1 U2527 ( .A(IR_REG_11__SCAN_IN), .ZN(n4866) );
  NOR2_X1 U2528 ( .A1(IR_REG_21__SCAN_IN), .A2(IR_REG_24__SCAN_IN), .ZN(n2501)
         );
  INV_X1 U2529 ( .A(IR_REG_12__SCAN_IN), .ZN(n2668) );
  AND2_X2 U2530 ( .A1(n2666), .A2(n2353), .ZN(n2673) );
  AOI21_X2 U2531 ( .B1(n3524), .B2(n3523), .A(n3522), .ZN(n3555) );
  INV_X1 U2532 ( .A(n2741), .ZN(n2234) );
  INV_X2 U2533 ( .A(n2741), .ZN(n2235) );
  AND3_X1 U2534 ( .A1(n2475), .A2(n2439), .A3(n2673), .ZN(n2850) );
  NAND2_X1 U2535 ( .A1(n2399), .A2(n2398), .ZN(n2602) );
  AOI21_X1 U2536 ( .B1(n2402), .B2(n2404), .A(n2261), .ZN(n2398) );
  NAND2_X1 U2537 ( .A1(n2921), .A2(n4666), .ZN(n3118) );
  NAND2_X1 U2538 ( .A1(n3730), .A2(n3775), .ZN(n2468) );
  NOR2_X1 U2539 ( .A1(n2776), .A2(n3694), .ZN(n2785) );
  AND2_X1 U2540 ( .A1(n4286), .A2(n2832), .ZN(n4234) );
  NOR2_X1 U2541 ( .A1(n2421), .A2(n2649), .ZN(n2420) );
  INV_X1 U2542 ( .A(n2424), .ZN(n2421) );
  NOR2_X1 U2543 ( .A1(n2582), .A2(n2406), .ZN(n2405) );
  OR2_X1 U2544 ( .A1(n3035), .A2(D_REG_1__SCAN_IN), .ZN(n2984) );
  NOR2_X1 U2545 ( .A1(n2387), .A2(n2385), .ZN(n2484) );
  NAND2_X1 U2546 ( .A1(n2501), .A2(n2502), .ZN(n2387) );
  AND2_X1 U2547 ( .A1(n2733), .A2(n4983), .ZN(n2734) );
  AND2_X1 U2548 ( .A1(n2497), .A2(n2453), .ZN(n2451) );
  OAI22_X1 U2549 ( .A1(n3228), .A2(n3674), .B1(n3663), .B2(n4360), .ZN(n2944)
         );
  OAI22_X1 U2550 ( .A1(n3228), .A2(n3678), .B1(n3677), .B2(n4360), .ZN(n2942)
         );
  OR2_X1 U2551 ( .A1(n2750), .A2(n4973), .ZN(n2767) );
  NAND3_X1 U2552 ( .A1(n3121), .A2(n2985), .A3(n2984), .ZN(n3005) );
  INV_X1 U2553 ( .A(n2529), .ZN(n2843) );
  OR2_X1 U2554 ( .A1(n3089), .A2(n3088), .ZN(n2327) );
  NAND2_X1 U2555 ( .A1(n2362), .A2(n2361), .ZN(n2368) );
  NAND2_X1 U2556 ( .A1(n2364), .A2(REG2_REG_4__SCAN_IN), .ZN(n2361) );
  NAND2_X1 U2557 ( .A1(n2364), .A2(n4526), .ZN(n2363) );
  XNOR2_X1 U2558 ( .A(n3098), .B(n2325), .ZN(n3065) );
  NAND2_X1 U2559 ( .A1(n4616), .A2(n4080), .ZN(n4081) );
  AND2_X1 U2560 ( .A1(n4268), .A2(n4257), .ZN(n2436) );
  NAND2_X1 U2561 ( .A1(n2407), .A2(n2245), .ZN(n2404) );
  AND2_X1 U2562 ( .A1(n2922), .A2(n3866), .ZN(n3126) );
  AND2_X1 U2563 ( .A1(n2983), .A2(n3036), .ZN(n3121) );
  NAND2_X1 U2564 ( .A1(n2511), .A2(n2510), .ZN(n2513) );
  NAND2_X1 U2565 ( .A1(n2509), .A2(IR_REG_31__SCAN_IN), .ZN(n2510) );
  NOR2_X1 U2566 ( .A1(n2866), .A2(n3015), .ZN(n2867) );
  XNOR2_X1 U2567 ( .A(n4081), .B(n4668), .ZN(n4625) );
  INV_X1 U2568 ( .A(n2308), .ZN(n2306) );
  INV_X1 U2569 ( .A(n2310), .ZN(n2304) );
  AND2_X1 U2570 ( .A1(n3757), .A2(n4538), .ZN(n2339) );
  NAND2_X1 U2571 ( .A1(n2448), .A2(n4548), .ZN(n2337) );
  NAND2_X1 U2572 ( .A1(n4019), .A2(n2445), .ZN(n2444) );
  NAND2_X1 U2573 ( .A1(n4022), .A2(REG1_REG_2__SCAN_IN), .ZN(n2445) );
  OR2_X1 U2574 ( .A1(n3163), .A2(n2357), .ZN(n2356) );
  AND2_X1 U2575 ( .A1(n4523), .A2(REG2_REG_7__SCAN_IN), .ZN(n2357) );
  AND2_X1 U2576 ( .A1(n2359), .A2(n2358), .ZN(n4097) );
  NAND2_X1 U2577 ( .A1(n4096), .A2(REG2_REG_15__SCAN_IN), .ZN(n2358) );
  NAND2_X1 U2578 ( .A1(n2237), .A2(n2840), .ZN(n2318) );
  NOR2_X1 U2579 ( .A1(n2430), .A2(n2756), .ZN(n2429) );
  INV_X1 U2580 ( .A(n2432), .ZN(n2430) );
  INV_X1 U2581 ( .A(n2241), .ZN(n2427) );
  INV_X1 U2582 ( .A(n2411), .ZN(n2410) );
  OAI21_X1 U2583 ( .B1(n4337), .B2(n2412), .A(n2736), .ZN(n2411) );
  INV_X1 U2584 ( .A(n2725), .ZN(n2412) );
  OR2_X1 U2585 ( .A1(n2699), .A2(n2397), .ZN(n2396) );
  INV_X1 U2586 ( .A(n2689), .ZN(n2397) );
  AOI21_X1 U2587 ( .B1(n2425), .B2(n2612), .A(n2250), .ZN(n2424) );
  NAND2_X1 U2588 ( .A1(n2391), .A2(n4356), .ZN(n2389) );
  NAND2_X1 U2589 ( .A1(n2928), .A2(n3197), .ZN(n3901) );
  NOR2_X1 U2590 ( .A1(n4218), .A2(n2284), .ZN(n2283) );
  INV_X1 U2591 ( .A(IR_REG_26__SCAN_IN), .ZN(n4806) );
  INV_X1 U2592 ( .A(IR_REG_23__SCAN_IN), .ZN(n2871) );
  INV_X1 U2593 ( .A(n2556), .ZN(n2452) );
  NOR2_X1 U2594 ( .A1(n2991), .A2(n2460), .ZN(n2459) );
  INV_X1 U2595 ( .A(n2982), .ZN(n2460) );
  OAI22_X1 U2596 ( .A1(n3677), .A2(n3191), .B1(n2928), .B2(n3618), .ZN(n2927)
         );
  OAI22_X1 U2597 ( .A1(n2928), .A2(n3674), .B1(n3618), .B2(n3191), .ZN(n2940)
         );
  NAND2_X1 U2598 ( .A1(n2462), .A2(n2248), .ZN(n3765) );
  NOR2_X1 U2599 ( .A1(n3650), .A2(n3651), .ZN(n2466) );
  OAI21_X1 U2600 ( .B1(n3714), .B2(n3650), .A(n3651), .ZN(n3766) );
  NAND2_X1 U2601 ( .A1(n2349), .A2(n2272), .ZN(n2343) );
  NAND3_X1 U2602 ( .A1(n2345), .A2(n2344), .A3(n2349), .ZN(n2342) );
  OR2_X1 U2603 ( .A1(n2921), .A2(n2935), .ZN(n2488) );
  NAND2_X1 U2604 ( .A1(n2468), .A2(n2467), .ZN(n2465) );
  XNOR2_X1 U2605 ( .A(n3418), .B(n2232), .ZN(n3523) );
  AND2_X1 U2606 ( .A1(n2338), .A2(n2337), .ZN(n4553) );
  NAND2_X1 U2607 ( .A1(n3743), .A2(n3744), .ZN(n2481) );
  INV_X1 U2608 ( .A(n3589), .ZN(n3590) );
  OR2_X1 U2609 ( .A1(n2777), .A2(n2785), .ZN(n3693) );
  NAND2_X1 U2610 ( .A1(n4021), .A2(n4020), .ZN(n4019) );
  XNOR2_X1 U2611 ( .A(n2444), .B(n4527), .ZN(n3052) );
  NOR2_X1 U2612 ( .A1(n3052), .A2(n3207), .ZN(n3063) );
  XNOR2_X1 U2613 ( .A(n3064), .B(n2371), .ZN(n3074) );
  OAI22_X1 U2614 ( .A1(n3070), .A2(n2365), .B1(n2251), .B2(n2368), .ZN(n3101)
         );
  NAND2_X1 U2615 ( .A1(n2367), .A2(n2366), .ZN(n2365) );
  INV_X1 U2616 ( .A(n2251), .ZN(n2366) );
  NAND2_X1 U2617 ( .A1(n4525), .A2(REG1_REG_5__SCAN_IN), .ZN(n2326) );
  NAND2_X1 U2618 ( .A1(n2321), .A2(n2442), .ZN(n3162) );
  NAND2_X1 U2619 ( .A1(n4523), .A2(REG1_REG_7__SCAN_IN), .ZN(n2442) );
  OR2_X1 U2620 ( .A1(n3159), .A2(n2267), .ZN(n2321) );
  NAND2_X1 U2621 ( .A1(n4589), .A2(n2323), .ZN(n4063) );
  NAND2_X1 U2622 ( .A1(n4522), .A2(REG1_REG_11__SCAN_IN), .ZN(n2323) );
  OR2_X1 U2623 ( .A1(n4613), .A2(n4612), .ZN(n2359) );
  AOI22_X1 U2624 ( .A1(n4171), .A2(n2775), .B1(n4385), .B2(n4183), .ZN(n4153)
         );
  AOI21_X1 U2625 ( .B1(n4173), .B2(n3961), .A(n3852), .ZN(n4155) );
  AOI21_X1 U2626 ( .B1(n2290), .B2(n3950), .A(n2288), .ZN(n2287) );
  AND2_X1 U2627 ( .A1(n2433), .A2(n2435), .ZN(n2432) );
  NAND2_X1 U2628 ( .A1(n3984), .A2(n4240), .ZN(n2435) );
  NAND2_X1 U2629 ( .A1(n2241), .A2(n2436), .ZN(n2433) );
  NOR2_X1 U2630 ( .A1(n4252), .A2(n4255), .ZN(n4251) );
  AND2_X1 U2631 ( .A1(n4236), .A2(n2835), .ZN(n4255) );
  AOI22_X1 U2632 ( .A1(n3544), .A2(n2717), .B1(n4557), .B2(n3598), .ZN(n4335)
         );
  NAND2_X1 U2633 ( .A1(n4335), .A2(n4337), .ZN(n4334) );
  OR2_X1 U2634 ( .A1(n2700), .A2(n5067), .ZN(n2709) );
  OAI21_X1 U2635 ( .B1(n3487), .B2(n2677), .A(n2676), .ZN(n3429) );
  INV_X1 U2636 ( .A(n2420), .ZN(n2419) );
  AOI21_X1 U2637 ( .B1(n2420), .B2(n2418), .A(n2249), .ZN(n2417) );
  INV_X1 U2638 ( .A(n2425), .ZN(n2418) );
  AOI21_X1 U2639 ( .B1(n3918), .B2(n2300), .A(n2299), .ZN(n2298) );
  INV_X1 U2640 ( .A(n3916), .ZN(n2300) );
  INV_X1 U2641 ( .A(n3915), .ZN(n2299) );
  INV_X1 U2642 ( .A(n3992), .ZN(n3390) );
  INV_X1 U2643 ( .A(n2403), .ZN(n2402) );
  OAI21_X1 U2644 ( .B1(n2405), .B2(n2404), .A(n2590), .ZN(n2403) );
  NOR2_X1 U2645 ( .A1(n3245), .A2(n2311), .ZN(n2310) );
  INV_X1 U2646 ( .A(n3911), .ZN(n2311) );
  AOI21_X1 U2647 ( .B1(n2310), .B2(n2812), .A(n2309), .ZN(n2308) );
  INV_X1 U2648 ( .A(n3923), .ZN(n2309) );
  INV_X1 U2649 ( .A(n4357), .ZN(n2393) );
  INV_X1 U2650 ( .A(n4366), .ZN(n4342) );
  NAND2_X1 U2651 ( .A1(n2235), .A2(DATAI_0_), .ZN(n2276) );
  NAND2_X1 U2652 ( .A1(n2741), .A2(IR_REG_0__SCAN_IN), .ZN(n2277) );
  INV_X1 U2653 ( .A(n2807), .ZN(n3859) );
  AND2_X1 U2654 ( .A1(n4160), .A2(n3686), .ZN(n2914) );
  AND4_X1 U2655 ( .A1(n2684), .A2(n2683), .A3(n2682), .A4(n2681), .ZN(n3579)
         );
  NAND2_X1 U2656 ( .A1(n3126), .A2(n3850), .ZN(n4433) );
  AND3_X1 U2657 ( .A1(n2886), .A2(n2885), .A3(n2983), .ZN(n2893) );
  NAND2_X1 U2658 ( .A1(n2865), .A2(n3016), .ZN(n3035) );
  NOR2_X1 U2659 ( .A1(n2479), .A2(IR_REG_25__SCAN_IN), .ZN(n2477) );
  NAND2_X1 U2660 ( .A1(n2869), .A2(n2872), .ZN(n3041) );
  OR2_X1 U2661 ( .A1(n2870), .A2(n2871), .ZN(n2872) );
  NAND2_X1 U2662 ( .A1(n2804), .A2(IR_REG_31__SCAN_IN), .ZN(n2805) );
  NOR2_X1 U2663 ( .A1(n2667), .A2(n2500), .ZN(n2353) );
  INV_X1 U2664 ( .A(IR_REG_13__SCAN_IN), .ZN(n2498) );
  INV_X1 U2665 ( .A(IR_REG_9__SCAN_IN), .ZN(n2624) );
  OR3_X1 U2666 ( .A1(n2620), .A2(IR_REG_7__SCAN_IN), .A3(IR_REG_8__SCAN_IN), 
        .ZN(n2623) );
  INV_X1 U2667 ( .A(n4194), .ZN(n4385) );
  AND4_X1 U2668 ( .A1(n2596), .A2(n2595), .A3(n2594), .A4(n2593), .ZN(n3368)
         );
  INV_X1 U2669 ( .A(n3192), .ZN(n3127) );
  OR2_X1 U2670 ( .A1(n3005), .A2(n3000), .ZN(n4528) );
  INV_X1 U2671 ( .A(n4531), .ZN(n4559) );
  OR2_X1 U2672 ( .A1(n3005), .A2(n2989), .ZN(n3813) );
  OAI21_X1 U2673 ( .B1(n4261), .B2(n2843), .A(n2527), .ZN(n4268) );
  INV_X1 U2674 ( .A(n3368), .ZN(n3995) );
  INV_X1 U2675 ( .A(n3305), .ZN(n3999) );
  NOR2_X1 U2676 ( .A1(n3105), .A2(n3104), .ZN(n3163) );
  OAI21_X1 U2677 ( .B1(n4625), .B2(n2331), .A(n2329), .ZN(n4639) );
  OR2_X1 U2678 ( .A1(n4638), .A2(REG1_REG_16__SCAN_IN), .ZN(n2331) );
  INV_X1 U2679 ( .A(n4638), .ZN(n2330) );
  NAND2_X1 U2680 ( .A1(n2295), .A2(n2293), .ZN(n2916) );
  INV_X1 U2681 ( .A(n4137), .ZN(n2295) );
  AND2_X1 U2682 ( .A1(n2909), .A2(n2294), .ZN(n2293) );
  INV_X1 U2683 ( .A(n2908), .ZN(n2294) );
  OR2_X1 U2684 ( .A1(n2916), .A2(n4702), .ZN(n2912) );
  NAND2_X1 U2685 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2534)
         );
  NOR2_X1 U2686 ( .A1(n2560), .A2(n2392), .ZN(n2391) );
  INV_X1 U2687 ( .A(n2551), .ZN(n2392) );
  NOR2_X1 U2688 ( .A1(IR_REG_22__SCAN_IN), .A2(IR_REG_23__SCAN_IN), .ZN(n2386)
         );
  NOR2_X1 U2689 ( .A1(IR_REG_19__SCAN_IN), .A2(IR_REG_18__SCAN_IN), .ZN(n2502)
         );
  NAND2_X1 U2690 ( .A1(n2351), .A2(n2798), .ZN(n2350) );
  INV_X1 U2691 ( .A(n2795), .ZN(n2351) );
  INV_X1 U2692 ( .A(IR_REG_14__SCAN_IN), .ZN(n4982) );
  INV_X1 U2693 ( .A(IR_REG_18__SCAN_IN), .ZN(n4983) );
  NAND2_X1 U2694 ( .A1(n2240), .A2(n3638), .ZN(n2463) );
  NAND2_X1 U2695 ( .A1(n2468), .A2(n2247), .ZN(n2462) );
  INV_X1 U2696 ( .A(n3365), .ZN(n2349) );
  NAND2_X1 U2697 ( .A1(n3701), .A2(n3699), .ZN(n3582) );
  INV_X1 U2698 ( .A(REG3_REG_12__SCAN_IN), .ZN(n2650) );
  INV_X1 U2699 ( .A(n3091), .ZN(n2364) );
  INV_X1 U2700 ( .A(n3952), .ZN(n2288) );
  INV_X1 U2701 ( .A(REG3_REG_14__SCAN_IN), .ZN(n2678) );
  OR2_X1 U2702 ( .A1(n2651), .A2(n2650), .ZN(n2660) );
  AND2_X1 U2703 ( .A1(n2611), .A2(n2256), .ZN(n2425) );
  OR2_X1 U2704 ( .A1(n2603), .A2(n5057), .ZN(n2614) );
  NAND2_X1 U2705 ( .A1(n2305), .A2(n2302), .ZN(n2813) );
  AOI21_X1 U2706 ( .B1(n2308), .B2(n2304), .A(n2303), .ZN(n2302) );
  XNOR2_X1 U2707 ( .A(n2514), .B(n3021), .ZN(n2516) );
  INV_X1 U2708 ( .A(n2313), .ZN(n2899) );
  AOI21_X1 U2709 ( .B1(n4173), .B2(n2244), .A(n2314), .ZN(n2313) );
  INV_X1 U2710 ( .A(n2318), .ZN(n2314) );
  AND2_X1 U2711 ( .A1(n2234), .A2(DATAI_20_), .ZN(n4290) );
  NAND2_X1 U2712 ( .A1(n4434), .A2(n4530), .ZN(n2279) );
  NAND2_X1 U2713 ( .A1(n3342), .A2(n2263), .ZN(n2282) );
  NOR2_X1 U2714 ( .A1(n3347), .A2(n2890), .ZN(n2281) );
  NAND2_X1 U2715 ( .A1(n3859), .A2(n2286), .ZN(n2808) );
  NAND2_X1 U2716 ( .A1(n4291), .A2(n2543), .ZN(n2388) );
  OR2_X1 U2717 ( .A1(n3035), .A2(n2884), .ZN(n2983) );
  INV_X1 U2718 ( .A(IR_REG_22__SCAN_IN), .ZN(n5023) );
  NOR2_X1 U2719 ( .A1(IR_REG_16__SCAN_IN), .A2(IR_REG_17__SCAN_IN), .ZN(n2733)
         );
  INV_X1 U2720 ( .A(IR_REG_8__SCAN_IN), .ZN(n2499) );
  NAND2_X1 U2721 ( .A1(n2462), .A2(n2463), .ZN(n3714) );
  NOR2_X1 U2722 ( .A1(n2614), .A2(n2613), .ZN(n2627) );
  CLKBUF_X1 U2723 ( .A(n2536), .Z(n2562) );
  NAND2_X1 U2724 ( .A1(n2338), .A2(n2265), .ZN(n3723) );
  NAND2_X1 U2725 ( .A1(n3235), .A2(n2346), .ZN(n2345) );
  NOR2_X1 U2726 ( .A1(n2470), .A2(n2236), .ZN(n2346) );
  AOI21_X1 U2727 ( .B1(n3594), .B2(n3593), .A(n3595), .ZN(n4538) );
  NAND2_X1 U2728 ( .A1(n2748), .A2(REG3_REG_23__SCAN_IN), .ZN(n2750) );
  NAND2_X1 U2729 ( .A1(n2342), .A2(n2340), .ZN(n2456) );
  NOR2_X1 U2730 ( .A1(n2458), .A2(n2341), .ZN(n2340) );
  OR2_X1 U2731 ( .A1(n3376), .A2(n2246), .ZN(n2458) );
  INV_X1 U2732 ( .A(n2343), .ZN(n2341) );
  AND2_X1 U2733 ( .A1(n2939), .A2(n2940), .ZN(n2941) );
  INV_X1 U2734 ( .A(n2944), .ZN(n2943) );
  INV_X1 U2735 ( .A(REG3_REG_6__SCAN_IN), .ZN(n3060) );
  NAND2_X1 U2736 ( .A1(n2961), .A2(n2962), .ZN(n2963) );
  INV_X1 U2737 ( .A(n4546), .ZN(n3805) );
  NOR2_X1 U2738 ( .A1(n2679), .A2(n2678), .ZN(n2690) );
  NOR2_X1 U2739 ( .A1(n3062), .A2(n2441), .ZN(n2322) );
  INV_X1 U2740 ( .A(n2444), .ZN(n3062) );
  NOR2_X1 U2741 ( .A1(n3074), .A2(n4709), .ZN(n3073) );
  INV_X1 U2742 ( .A(n2367), .ZN(n2369) );
  OAI21_X1 U2743 ( .B1(n4037), .B2(n3338), .A(n4036), .ZN(n4570) );
  INV_X1 U2744 ( .A(n2356), .ZN(n2355) );
  NAND2_X1 U2745 ( .A1(n4065), .A2(n4066), .ZN(n4069) );
  NAND2_X1 U2746 ( .A1(n4522), .A2(REG2_REG_11__SCAN_IN), .ZN(n2360) );
  NAND2_X1 U2747 ( .A1(n4667), .A2(n2384), .ZN(n2383) );
  INV_X1 U2748 ( .A(REG2_REG_17__SCAN_IN), .ZN(n2384) );
  INV_X1 U2749 ( .A(n2383), .ZN(n2381) );
  NAND2_X1 U2750 ( .A1(n4520), .A2(REG2_REG_18__SCAN_IN), .ZN(n2382) );
  OAI21_X1 U2751 ( .B1(n4173), .B2(n2317), .A(n2315), .ZN(n2320) );
  AOI21_X1 U2752 ( .B1(n2318), .B2(n2316), .A(n3839), .ZN(n2315) );
  NAND2_X1 U2753 ( .A1(n2318), .A2(n3836), .ZN(n2317) );
  NOR2_X1 U2754 ( .A1(n2244), .A2(n3835), .ZN(n2316) );
  AND2_X1 U2755 ( .A1(n2793), .A2(n2792), .ZN(n4131) );
  NOR2_X1 U2756 ( .A1(n3839), .A2(n3835), .ZN(n3895) );
  AOI21_X1 U2757 ( .B1(n4153), .B2(n2784), .A(n2783), .ZN(n2897) );
  AND2_X1 U2758 ( .A1(n2839), .A2(n2840), .ZN(n4154) );
  AOI21_X1 U2759 ( .B1(n2429), .B2(n2427), .A(n2254), .ZN(n2426) );
  INV_X1 U2760 ( .A(n2429), .ZN(n2428) );
  AND2_X1 U2761 ( .A1(n3827), .A2(n2291), .ZN(n2290) );
  NAND2_X1 U2762 ( .A1(n2834), .A2(n2292), .ZN(n2291) );
  INV_X1 U2763 ( .A(n3823), .ZN(n2292) );
  AND2_X1 U2764 ( .A1(n2521), .A2(n2520), .ZN(n4243) );
  AND2_X1 U2765 ( .A1(n2743), .A2(REG3_REG_22__SCAN_IN), .ZN(n2748) );
  AND2_X1 U2766 ( .A1(n3882), .A2(n4235), .ZN(n4270) );
  AOI21_X1 U2767 ( .B1(n2410), .B2(n2412), .A(n2262), .ZN(n2409) );
  NAND2_X1 U2768 ( .A1(n2728), .A2(REG3_REG_19__SCAN_IN), .ZN(n2737) );
  OR2_X1 U2769 ( .A1(n2737), .A2(n4815), .ZN(n2742) );
  AND2_X1 U2770 ( .A1(n2718), .A2(REG3_REG_18__SCAN_IN), .ZN(n2728) );
  AND2_X1 U2771 ( .A1(n4312), .A2(n4229), .ZN(n3867) );
  OAI21_X1 U2772 ( .B1(n3429), .B2(n2396), .A(n2394), .ZN(n3503) );
  INV_X1 U2773 ( .A(n2395), .ZN(n2394) );
  OAI21_X1 U2774 ( .B1(n3428), .B2(n2396), .A(n2698), .ZN(n2395) );
  NAND2_X1 U2775 ( .A1(n3503), .A2(n3502), .ZN(n3501) );
  AND2_X1 U2776 ( .A1(n2712), .A2(n2711), .ZN(n4533) );
  NAND2_X1 U2777 ( .A1(n2416), .A2(n2414), .ZN(n3487) );
  AOI21_X1 U2778 ( .B1(n2253), .B2(n2417), .A(n2415), .ZN(n2414) );
  NOR2_X1 U2779 ( .A1(n2821), .A2(n3537), .ZN(n2415) );
  NAND2_X1 U2780 ( .A1(n2422), .A2(n2424), .ZN(n3444) );
  NAND2_X1 U2781 ( .A1(n3324), .A2(n2425), .ZN(n2422) );
  NAND2_X1 U2782 ( .A1(n2816), .A2(n3916), .ZN(n3325) );
  AND3_X1 U2783 ( .A1(n2492), .A2(n2555), .A3(n2554), .ZN(n2947) );
  OR2_X1 U2784 ( .A1(n2904), .A2(n2494), .ZN(n2505) );
  NAND2_X1 U2785 ( .A1(n2904), .A2(n2503), .ZN(n2504) );
  AND2_X1 U2786 ( .A1(IR_REG_28__SCAN_IN), .A2(IR_REG_27__SCAN_IN), .ZN(n2494)
         );
  NAND2_X1 U2787 ( .A1(n3191), .A2(n3192), .ZN(n4370) );
  NOR2_X1 U2788 ( .A1(n4377), .A2(n4381), .ZN(n4376) );
  INV_X1 U2789 ( .A(n4121), .ZN(n4381) );
  INV_X1 U2790 ( .A(n4133), .ZN(n2913) );
  AND2_X1 U2791 ( .A1(n2235), .A2(DATAI_28_), .ZN(n4143) );
  INV_X1 U2792 ( .A(n4143), .ZN(n3686) );
  NAND2_X1 U2793 ( .A1(n4223), .A2(n2239), .ZN(n4182) );
  NAND2_X1 U2794 ( .A1(n4223), .A2(n2283), .ZN(n4199) );
  AND2_X1 U2795 ( .A1(n4223), .A2(n4399), .ZN(n4212) );
  NOR2_X1 U2796 ( .A1(n4250), .A2(n4240), .ZN(n4223) );
  INV_X1 U2797 ( .A(n3787), .ZN(n4257) );
  OR2_X1 U2798 ( .A1(n4278), .A2(n4257), .ZN(n4250) );
  NOR2_X1 U2799 ( .A1(n4326), .A2(n4290), .ZN(n4299) );
  OR2_X1 U2800 ( .A1(n4345), .A2(n3875), .ZN(n4326) );
  AND2_X1 U2801 ( .A1(n2705), .A2(n2704), .ZN(n4436) );
  NOR3_X1 U2802 ( .A1(n4449), .A2(n3584), .A3(n3496), .ZN(n3546) );
  NOR2_X1 U2803 ( .A1(n4449), .A2(n3584), .ZN(n3504) );
  NOR2_X1 U2804 ( .A1(n2282), .A2(n3525), .ZN(n3489) );
  NAND2_X1 U2805 ( .A1(n3342), .A2(n2281), .ZN(n3442) );
  NAND2_X1 U2806 ( .A1(n3342), .A2(n3379), .ZN(n3441) );
  OR2_X1 U2807 ( .A1(n3290), .A2(n3291), .ZN(n3331) );
  NOR2_X1 U2808 ( .A1(n3331), .A2(n3332), .ZN(n3342) );
  NAND2_X1 U2809 ( .A1(n4298), .A2(n4696), .ZN(n4694) );
  OR2_X1 U2810 ( .A1(n3263), .A2(n3272), .ZN(n3290) );
  INV_X1 U2811 ( .A(n2400), .ZN(n3259) );
  AOI21_X1 U2812 ( .B1(n2570), .B2(n2405), .A(n2401), .ZN(n2400) );
  INV_X1 U2813 ( .A(n2407), .ZN(n2401) );
  NOR2_X1 U2814 ( .A1(n4683), .A2(n3231), .ZN(n3178) );
  INV_X1 U2815 ( .A(n4433), .ZN(n4380) );
  INV_X1 U2816 ( .A(n4694), .ZN(n4441) );
  INV_X1 U2817 ( .A(n4678), .ZN(n4701) );
  INV_X1 U2818 ( .A(n2985), .ZN(n3122) );
  NAND2_X1 U2819 ( .A1(n2852), .A2(n2851), .ZN(n3046) );
  AND2_X1 U2820 ( .A1(n2484), .A2(n2478), .ZN(n2476) );
  XNOR2_X1 U2821 ( .A(n2803), .B(n2802), .ZN(n3963) );
  NAND2_X1 U2822 ( .A1(n2796), .A2(IR_REG_31__SCAN_IN), .ZN(n2800) );
  AND2_X1 U2823 ( .A1(n2706), .A2(n2697), .ZN(n4096) );
  INV_X1 U2824 ( .A(IR_REG_3__SCAN_IN), .ZN(n2557) );
  NOR2_X1 U2825 ( .A1(n2965), .A2(n3314), .ZN(n2473) );
  XNOR2_X1 U2826 ( .A(n3671), .B(n3670), .ZN(n3692) );
  INV_X1 U2827 ( .A(n3989), .ZN(n3704) );
  INV_X1 U2828 ( .A(n3993), .ZN(n3447) );
  NAND2_X1 U2829 ( .A1(n2461), .A2(n2982), .ZN(n2990) );
  OR2_X1 U2830 ( .A1(n3375), .A2(n3376), .ZN(n2461) );
  NAND2_X1 U2831 ( .A1(n2235), .A2(DATAI_21_), .ZN(n4415) );
  AND4_X1 U2832 ( .A1(n2640), .A2(n2639), .A3(n2638), .A4(n2637), .ZN(n3538)
         );
  INV_X1 U2833 ( .A(n2465), .ZN(n3783) );
  INV_X1 U2834 ( .A(n3638), .ZN(n2464) );
  OAI22_X1 U2835 ( .A1(n4546), .A2(n2947), .B1(n2928), .B2(n4528), .ZN(n3145)
         );
  NAND2_X1 U2836 ( .A1(n2336), .A2(n2447), .ZN(n4550) );
  INV_X1 U2837 ( .A(n4528), .ZN(n4556) );
  XNOR2_X1 U2838 ( .A(n2354), .B(n3794), .ZN(n3800) );
  INV_X1 U2839 ( .A(n3813), .ZN(n4554) );
  AND2_X1 U2840 ( .A1(n3003), .A2(n4651), .ZN(n4531) );
  INV_X1 U2841 ( .A(n4563), .ZN(n3811) );
  NOR2_X1 U2842 ( .A1(n3663), .A2(n2997), .ZN(n3974) );
  OAI21_X1 U2843 ( .B1(n3693), .B2(n2843), .A(n2782), .ZN(n4177) );
  NAND2_X1 U2844 ( .A1(n2774), .A2(n2773), .ZN(n4194) );
  NAND2_X1 U2845 ( .A1(n2762), .A2(n2761), .ZN(n4178) );
  INV_X1 U2846 ( .A(n4243), .ZN(n3983) );
  INV_X1 U2847 ( .A(n4533), .ZN(n4557) );
  INV_X1 U2848 ( .A(n4436), .ZN(n3986) );
  INV_X1 U2849 ( .A(n3538), .ZN(n3991) );
  CLKBUF_X1 U2850 ( .A(U4043), .Z(n3996) );
  INV_X1 U2851 ( .A(n2947), .ZN(n4363) );
  INV_X1 U2852 ( .A(n3228), .ZN(n4000) );
  AND2_X1 U2853 ( .A1(n3045), .A2(n3044), .ZN(n4006) );
  AND2_X1 U2854 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n4013)
         );
  OAI21_X1 U2855 ( .B1(n2372), .B2(n3047), .A(n2324), .ZN(n4010) );
  NAND2_X1 U2856 ( .A1(n2372), .A2(n3047), .ZN(n2324) );
  NOR2_X1 U2857 ( .A1(n3073), .A2(n2440), .ZN(n3089) );
  NOR2_X1 U2858 ( .A1(n3064), .A2(n2371), .ZN(n2440) );
  INV_X1 U2859 ( .A(n2327), .ZN(n3087) );
  OAI21_X1 U2860 ( .B1(n2369), .B2(n3070), .A(n2368), .ZN(n2370) );
  AOI21_X1 U2861 ( .B1(n3070), .B2(REG2_REG_4__SCAN_IN), .A(n2369), .ZN(n3092)
         );
  NOR2_X1 U2862 ( .A1(n3098), .A2(n2325), .ZN(n2443) );
  XNOR2_X1 U2863 ( .A(n4063), .B(n4043), .ZN(n4044) );
  NAND2_X1 U2864 ( .A1(n4044), .A2(REG1_REG_12__SCAN_IN), .ZN(n4065) );
  AND2_X1 U2865 ( .A1(n4006), .A2(n3973), .ZN(n4593) );
  INV_X1 U2866 ( .A(n2359), .ZN(n4611) );
  OR2_X1 U2867 ( .A1(n4625), .A2(REG1_REG_16__SCAN_IN), .ZN(n2332) );
  INV_X1 U2868 ( .A(n4082), .ZN(n2328) );
  NOR2_X1 U2869 ( .A1(n4639), .A2(n4084), .ZN(n4111) );
  NAND2_X1 U2870 ( .A1(n4632), .A2(n2383), .ZN(n4100) );
  NAND2_X1 U2871 ( .A1(n2378), .A2(n2377), .ZN(n4107) );
  NAND2_X1 U2872 ( .A1(n2380), .A2(n2382), .ZN(n2377) );
  NAND2_X1 U2873 ( .A1(n2431), .A2(n2432), .ZN(n4205) );
  NAND2_X1 U2874 ( .A1(n4251), .A2(n2241), .ZN(n2431) );
  NOR2_X1 U2875 ( .A1(n4251), .A2(n2436), .ZN(n4228) );
  NAND2_X1 U2876 ( .A1(n4334), .A2(n2725), .ZN(n4311) );
  NAND2_X1 U2877 ( .A1(n3427), .A2(n2689), .ZN(n3458) );
  OR2_X1 U2878 ( .A1(n3488), .A2(n3435), .ZN(n4449) );
  NAND2_X1 U2879 ( .A1(n2413), .A2(n2417), .ZN(n3404) );
  OR2_X1 U2880 ( .A1(n3324), .A2(n2419), .ZN(n2413) );
  NAND2_X1 U2881 ( .A1(n2297), .A2(n2298), .ZN(n3339) );
  OR2_X1 U2882 ( .A1(n3324), .A2(n2612), .ZN(n2423) );
  OR2_X1 U2883 ( .A1(n3118), .A2(n3002), .ZN(n4651) );
  OAI21_X1 U2884 ( .B1(n2570), .B2(n2404), .A(n2402), .ZN(n3282) );
  NAND2_X1 U2885 ( .A1(n2307), .A2(n2308), .ZN(n3260) );
  NAND2_X1 U2886 ( .A1(n3181), .A2(n2310), .ZN(n2307) );
  AND4_X1 U2887 ( .A1(n2566), .A2(n2565), .A3(n2564), .A4(n2563), .ZN(n3305)
         );
  NAND2_X1 U2888 ( .A1(n2312), .A2(n3911), .ZN(n3246) );
  OR2_X1 U2889 ( .A1(n3181), .A2(n2812), .ZN(n2312) );
  NAND2_X1 U2890 ( .A1(n4355), .A2(n2551), .ZN(n3133) );
  AND2_X1 U2891 ( .A1(n4654), .A2(n4380), .ZN(n4282) );
  NAND2_X1 U2892 ( .A1(n2275), .A2(n4360), .ZN(n4683) );
  INV_X1 U2893 ( .A(n4370), .ZN(n2275) );
  INV_X1 U2894 ( .A(n4328), .ZN(n4657) );
  XNOR2_X1 U2895 ( .A(n2807), .B(n3898), .ZN(n3201) );
  NAND2_X1 U2896 ( .A1(n3859), .A2(n2285), .ZN(n3194) );
  INV_X1 U2897 ( .A(n3193), .ZN(n2285) );
  INV_X1 U2898 ( .A(n4651), .ZN(n4643) );
  NAND2_X1 U2899 ( .A1(n3035), .A2(n3034), .ZN(n4664) );
  AND2_X1 U2900 ( .A1(n2673), .A2(n2438), .ZN(n2437) );
  INV_X1 U2901 ( .A(n3046), .ZN(n3083) );
  XNOR2_X1 U2902 ( .A(n2864), .B(IR_REG_26__SCAN_IN), .ZN(n3016) );
  OR2_X1 U2903 ( .A1(n2858), .A2(n2863), .ZN(n2864) );
  AND2_X1 U2904 ( .A1(n3041), .A2(STATE_REG_SCAN_IN), .ZN(n4666) );
  INV_X1 U2905 ( .A(n2922), .ZN(n3976) );
  XNOR2_X1 U2906 ( .A(n2800), .B(IR_REG_19__SCAN_IN), .ZN(n4519) );
  NOR2_X1 U2907 ( .A1(n2626), .A2(n2641), .ZN(n4567) );
  AND2_X1 U2908 ( .A1(n2609), .A2(n2600), .ZN(n4523) );
  AND2_X1 U2909 ( .A1(n2581), .A2(n2580), .ZN(n4525) );
  OAI22_X1 U2910 ( .A1(n4546), .A2(n2928), .B1(n3813), .B2(n3114), .ZN(n3115)
         );
  OAI21_X1 U2911 ( .B1(n2916), .B2(n4713), .A(n2918), .ZN(n2919) );
  NAND2_X1 U2912 ( .A1(n4702), .A2(n2910), .ZN(n2911) );
  NAND2_X1 U2913 ( .A1(n2374), .A2(n2373), .ZN(U3351) );
  NAND2_X1 U2914 ( .A1(U3149), .A2(DATAI_1_), .ZN(n2373) );
  AND2_X4 U2915 ( .A1(n2516), .A2(n2515), .ZN(n2538) );
  NAND2_X1 U2916 ( .A1(n2452), .A2(n2493), .ZN(n2577) );
  NAND2_X1 U2917 ( .A1(n4982), .A2(n2480), .ZN(n2479) );
  AND2_X1 U2918 ( .A1(n2968), .A2(n2967), .ZN(n2236) );
  INV_X1 U2919 ( .A(n3984), .ZN(n4400) );
  NAND2_X1 U2920 ( .A1(n2755), .A2(n2754), .ZN(n3984) );
  NAND2_X1 U2921 ( .A1(n4154), .A2(n2319), .ZN(n2237) );
  AND2_X1 U2922 ( .A1(n2298), .A2(n2296), .ZN(n2238) );
  AND2_X1 U2923 ( .A1(n2235), .A2(DATAI_24_), .ZN(n4218) );
  AND2_X1 U2924 ( .A1(n2283), .A2(n4183), .ZN(n2239) );
  AND2_X1 U2925 ( .A1(n2657), .A2(n2644), .ZN(n4522) );
  NOR2_X1 U2926 ( .A1(n3713), .A2(n3712), .ZN(n2240) );
  OR2_X1 U2927 ( .A1(n3984), .A2(n4240), .ZN(n2241) );
  AND2_X1 U2928 ( .A1(n2475), .A2(n2673), .ZN(n2858) );
  AND2_X1 U2929 ( .A1(n2465), .A2(n2464), .ZN(n2242) );
  OR2_X1 U2930 ( .A1(n3990), .A2(n3525), .ZN(n2243) );
  AND2_X1 U2931 ( .A1(n2840), .A2(n3961), .ZN(n2244) );
  NAND4_X1 U2932 ( .A1(n2542), .A2(n2541), .A3(n2540), .A4(n2539), .ZN(n2933)
         );
  OR2_X1 U2933 ( .A1(n3997), .A2(n3272), .ZN(n2245) );
  AND2_X1 U2934 ( .A1(n3416), .A2(n3415), .ZN(n2246) );
  AND2_X1 U2935 ( .A1(n4157), .A2(n3686), .ZN(n3835) );
  NOR2_X1 U2936 ( .A1(n3063), .A2(n2322), .ZN(n3064) );
  AND2_X1 U2937 ( .A1(n2240), .A2(n2467), .ZN(n2247) );
  INV_X1 U2938 ( .A(n2470), .ZN(n2469) );
  OAI21_X1 U2939 ( .B1(n2474), .B2(n2472), .A(n2471), .ZN(n2470) );
  AND2_X1 U2940 ( .A1(n2463), .A2(n2466), .ZN(n2248) );
  NOR2_X1 U2941 ( .A1(n2648), .A2(n2647), .ZN(n2249) );
  NOR2_X1 U2942 ( .A1(n3447), .A2(n3379), .ZN(n2250) );
  AND2_X1 U2943 ( .A1(n4525), .A2(REG2_REG_5__SCAN_IN), .ZN(n2251) );
  AND2_X1 U2944 ( .A1(n2327), .A2(n2326), .ZN(n3098) );
  NAND2_X1 U2945 ( .A1(n2549), .A2(n2497), .ZN(n2556) );
  OR2_X1 U2946 ( .A1(n2796), .A2(n2795), .ZN(n2252) );
  AND2_X1 U2947 ( .A1(n2419), .A2(n2243), .ZN(n2253) );
  AND2_X1 U2948 ( .A1(n4243), .A2(n4399), .ZN(n2254) );
  AND2_X1 U2949 ( .A1(n2417), .A2(n2243), .ZN(n2255) );
  OR2_X1 U2950 ( .A1(n3993), .A2(n3347), .ZN(n2256) );
  AND2_X1 U2951 ( .A1(n4632), .A2(n2379), .ZN(n2257) );
  INV_X1 U2952 ( .A(n4325), .ZN(n3985) );
  AND2_X1 U2953 ( .A1(n2722), .A2(n2721), .ZN(n4325) );
  AND2_X1 U2954 ( .A1(n2508), .A2(n2482), .ZN(n2258) );
  INV_X1 U2955 ( .A(n2479), .ZN(n2478) );
  AND2_X1 U2956 ( .A1(n2332), .A2(n2328), .ZN(n2259) );
  NAND2_X1 U2957 ( .A1(n4363), .A2(n3231), .ZN(n2260) );
  INV_X1 U2958 ( .A(IR_REG_20__SCAN_IN), .ZN(n2802) );
  INV_X1 U2959 ( .A(n3618), .ZN(n3636) );
  INV_X2 U2960 ( .A(n3585), .ZN(n3663) );
  INV_X1 U2961 ( .A(n4524), .ZN(n2325) );
  AND2_X1 U2962 ( .A1(n2814), .A2(n3916), .ZN(n2261) );
  AND2_X1 U2963 ( .A1(n2673), .A2(n2478), .ZN(n2735) );
  INV_X1 U2964 ( .A(n3525), .ZN(n3537) );
  NAND2_X1 U2965 ( .A1(n2673), .A2(n4982), .ZN(n2687) );
  AND2_X1 U2966 ( .A1(n2334), .A2(n2333), .ZN(n3701) );
  INV_X1 U2967 ( .A(IR_REG_10__SCAN_IN), .ZN(n2453) );
  NAND2_X1 U2968 ( .A1(n2450), .A2(n3596), .ZN(n3755) );
  INV_X1 U2969 ( .A(n3898), .ZN(n2286) );
  AND2_X1 U2970 ( .A1(n4545), .A2(n4327), .ZN(n2262) );
  XOR2_X1 U2971 ( .A(n2232), .B(n3556), .Z(n3575) );
  INV_X1 U2972 ( .A(n3575), .ZN(n2335) );
  INV_X1 U2973 ( .A(n3852), .ZN(n2319) );
  INV_X1 U2974 ( .A(n3347), .ZN(n3379) );
  AND2_X1 U2975 ( .A1(n2281), .A2(n3422), .ZN(n2263) );
  INV_X1 U2976 ( .A(n3918), .ZN(n2301) );
  AND3_X1 U2977 ( .A1(n2451), .A2(n2493), .A3(n2549), .ZN(n2666) );
  OR2_X1 U2978 ( .A1(n3667), .A2(n3666), .ZN(n2264) );
  AND2_X1 U2979 ( .A1(n2337), .A2(n4549), .ZN(n2265) );
  INV_X1 U2980 ( .A(n2448), .ZN(n2447) );
  OAI21_X1 U2981 ( .B1(n3596), .B2(n2449), .A(n3756), .ZN(n2448) );
  INV_X1 U2982 ( .A(IR_REG_27__SCAN_IN), .ZN(n2482) );
  NAND2_X1 U2983 ( .A1(n2352), .A2(IR_REG_31__SCAN_IN), .ZN(n2870) );
  AND2_X1 U2984 ( .A1(n2339), .A2(n4548), .ZN(n2266) );
  AND2_X1 U2985 ( .A1(n3160), .A2(n4711), .ZN(n2267) );
  INV_X1 U2986 ( .A(n3757), .ZN(n2449) );
  AND2_X1 U2987 ( .A1(n2264), .A2(n3745), .ZN(n2268) );
  INV_X1 U2988 ( .A(IR_REG_28__SCAN_IN), .ZN(n2508) );
  INV_X1 U2989 ( .A(IR_REG_15__SCAN_IN), .ZN(n2480) );
  NAND2_X1 U2990 ( .A1(n2870), .A2(n2871), .ZN(n2869) );
  NAND2_X1 U2991 ( .A1(n2342), .A2(n2343), .ZN(n3375) );
  NAND2_X1 U2992 ( .A1(n2423), .A2(n2611), .ZN(n3341) );
  INV_X1 U2993 ( .A(n3921), .ZN(n2303) );
  NAND2_X1 U2994 ( .A1(n2345), .A2(n2344), .ZN(n3364) );
  NAND2_X1 U2995 ( .A1(n3235), .A2(n2963), .ZN(n3312) );
  NAND2_X1 U2996 ( .A1(n2235), .A2(DATAI_23_), .ZN(n4225) );
  INV_X1 U2997 ( .A(n4225), .ZN(n4240) );
  OR2_X1 U2998 ( .A1(n3584), .A2(n4558), .ZN(n2269) );
  NAND2_X1 U2999 ( .A1(n3429), .A2(n3428), .ZN(n3427) );
  XNOR2_X1 U3000 ( .A(n2805), .B(n5023), .ZN(n2922) );
  NOR3_X1 U3001 ( .A1(n4449), .A2(n2279), .A3(n2269), .ZN(n2280) );
  AND2_X1 U3002 ( .A1(n2461), .A2(n2459), .ZN(n2270) );
  INV_X1 U3003 ( .A(n3496), .ZN(n4530) );
  INV_X1 U3004 ( .A(n2278), .ZN(n4344) );
  NOR3_X1 U3005 ( .A1(n4449), .A2(n2279), .A3(n3584), .ZN(n2278) );
  OR2_X1 U3006 ( .A1(n2507), .A2(IR_REG_27__SCAN_IN), .ZN(n2271) );
  INV_X1 U3007 ( .A(n3930), .ZN(n2296) );
  INV_X1 U3008 ( .A(n3520), .ZN(n2455) );
  AND2_X1 U3009 ( .A1(n2716), .A2(n2723), .ZN(n4099) );
  INV_X1 U3010 ( .A(n4099), .ZN(n4667) );
  INV_X1 U3011 ( .A(n2928), .ZN(n2543) );
  NAND2_X1 U3012 ( .A1(n2235), .A2(DATAI_25_), .ZN(n4197) );
  INV_X1 U3013 ( .A(n4197), .ZN(n2284) );
  AND2_X1 U3014 ( .A1(n2974), .A2(n2973), .ZN(n2272) );
  AND2_X1 U3015 ( .A1(n4364), .A2(n2388), .ZN(n2273) );
  NAND2_X1 U3016 ( .A1(n2393), .A2(n2809), .ZN(n4355) );
  INV_X1 U3017 ( .A(n4183), .ZN(n4176) );
  NAND2_X1 U3018 ( .A1(n2234), .A2(DATAI_26_), .ZN(n4183) );
  AND2_X1 U3019 ( .A1(n4633), .A2(n2382), .ZN(n2274) );
  INV_X1 U3020 ( .A(n2380), .ZN(n2379) );
  OR2_X1 U3021 ( .A1(n4101), .A2(n2381), .ZN(n2380) );
  XNOR2_X1 U3022 ( .A(n2568), .B(IR_REG_4__SCAN_IN), .ZN(n4526) );
  XNOR2_X1 U3023 ( .A(n2514), .B(IR_REG_30__SCAN_IN), .ZN(n3031) );
  AND2_X1 U3024 ( .A1(n2567), .A2(n2559), .ZN(n4527) );
  INV_X1 U3025 ( .A(n4527), .ZN(n2441) );
  INV_X1 U3026 ( .A(n2280), .ZN(n4345) );
  INV_X1 U3027 ( .A(n2282), .ZN(n3405) );
  NAND3_X1 U3028 ( .A1(n2475), .A2(n4806), .A3(n2673), .ZN(n2507) );
  OAI21_X1 U3029 ( .B1(n2833), .B2(n3950), .A(n2290), .ZN(n4207) );
  NAND2_X1 U3030 ( .A1(n2289), .A2(n2287), .ZN(n2838) );
  NAND2_X1 U3031 ( .A1(n2833), .A2(n2290), .ZN(n2289) );
  NAND2_X1 U3032 ( .A1(n2297), .A2(n2238), .ZN(n2817) );
  XNOR2_X1 U3033 ( .A(n2320), .B(n2900), .ZN(n2907) );
  NAND2_X1 U3034 ( .A1(n3162), .A2(n3161), .ZN(n4036) );
  NOR2_X1 U3035 ( .A1(n3099), .A2(n2443), .ZN(n3159) );
  XNOR2_X2 U3036 ( .A(n2534), .B(IR_REG_1__SCAN_IN), .ZN(n2372) );
  NAND2_X1 U3037 ( .A1(n4082), .A2(n2330), .ZN(n2329) );
  INV_X1 U3038 ( .A(n2332), .ZN(n4626) );
  NAND2_X1 U3039 ( .A1(n3576), .A2(n2335), .ZN(n2333) );
  OAI21_X1 U3040 ( .B1(n3576), .B2(n2335), .A(n3577), .ZN(n2334) );
  NAND3_X1 U3041 ( .A1(n2446), .A2(n3802), .A3(n2339), .ZN(n2336) );
  NAND3_X1 U3042 ( .A1(n2446), .A2(n3802), .A3(n2266), .ZN(n2338) );
  NAND3_X1 U3043 ( .A1(n2446), .A2(n3802), .A3(n4538), .ZN(n2450) );
  OAI21_X1 U3044 ( .B1(n3235), .B2(n2473), .A(n2469), .ZN(n3566) );
  INV_X1 U3045 ( .A(n3565), .ZN(n2348) );
  NOR2_X1 U3046 ( .A1(n2796), .A2(n2350), .ZN(n2860) );
  NAND2_X1 U3047 ( .A1(n2860), .A2(n5023), .ZN(n2352) );
  NAND2_X1 U3048 ( .A1(n2481), .A2(n3745), .ZN(n2354) );
  XNOR2_X2 U3049 ( .A(n4060), .B(n4064), .ZN(n4052) );
  OR2_X1 U3050 ( .A1(n3059), .A2(n2363), .ZN(n2362) );
  OR2_X1 U3051 ( .A1(n3059), .A2(n2371), .ZN(n2367) );
  XNOR2_X1 U3052 ( .A(n3059), .B(n4526), .ZN(n3070) );
  INV_X1 U3053 ( .A(n2370), .ZN(n3090) );
  INV_X1 U3054 ( .A(n4526), .ZN(n2371) );
  NAND2_X1 U3055 ( .A1(n2372), .A2(REG2_REG_1__SCAN_IN), .ZN(n4024) );
  NAND2_X1 U3056 ( .A1(n2372), .A2(REG1_REG_1__SCAN_IN), .ZN(n3051) );
  NAND2_X1 U3057 ( .A1(n2372), .A2(STATE_REG_SCAN_IN), .ZN(n2374) );
  XNOR2_X1 U3058 ( .A(n2372), .B(n3050), .ZN(n4014) );
  NAND2_X1 U3059 ( .A1(n2234), .A2(DATAI_1_), .ZN(n2375) );
  INV_X1 U3060 ( .A(n2372), .ZN(n2376) );
  NAND2_X1 U3061 ( .A1(n4045), .A2(n2372), .ZN(n4018) );
  NAND2_X1 U3062 ( .A1(n4631), .A2(n2274), .ZN(n2378) );
  NAND2_X1 U3063 ( .A1(n4631), .A2(n4633), .ZN(n4632) );
  NAND4_X1 U3064 ( .A1(n2386), .A2(n2802), .A3(n4844), .A4(n2713), .ZN(n2385)
         );
  NAND3_X1 U3065 ( .A1(n2390), .A2(n2389), .A3(n2260), .ZN(n3179) );
  NAND2_X1 U3066 ( .A1(n2391), .A2(n4357), .ZN(n2390) );
  NAND2_X1 U3067 ( .A1(n2570), .A2(n2402), .ZN(n2399) );
  NAND2_X1 U3068 ( .A1(n2570), .A2(n2569), .ZN(n3244) );
  INV_X1 U3069 ( .A(n2569), .ZN(n2406) );
  OR2_X1 U3070 ( .A1(n3998), .A2(n3303), .ZN(n2407) );
  NAND2_X1 U3071 ( .A1(n2408), .A2(n2409), .ZN(n4285) );
  NAND2_X1 U3072 ( .A1(n4335), .A2(n2410), .ZN(n2408) );
  NAND2_X1 U3073 ( .A1(n3324), .A2(n2255), .ZN(n2416) );
  OAI21_X1 U3074 ( .B1(n4251), .B2(n2428), .A(n2426), .ZN(n2434) );
  INV_X1 U3075 ( .A(n2434), .ZN(n4190) );
  NOR2_X1 U3076 ( .A1(n3151), .A2(n3149), .ZN(n3150) );
  XNOR2_X1 U3077 ( .A(n2939), .B(n2940), .ZN(n3149) );
  NAND2_X1 U3078 ( .A1(n3803), .A2(n4536), .ZN(n2446) );
  NAND2_X1 U3079 ( .A1(n2456), .A2(n2457), .ZN(n3521) );
  INV_X1 U3080 ( .A(n3633), .ZN(n2467) );
  OR2_X1 U3081 ( .A1(n2963), .A2(n3313), .ZN(n2471) );
  INV_X1 U3082 ( .A(n3314), .ZN(n2472) );
  AND2_X1 U3083 ( .A1(n2963), .A2(n3313), .ZN(n2474) );
  AND2_X1 U3084 ( .A1(n2673), .A2(n2476), .ZN(n2856) );
  NAND2_X1 U3085 ( .A1(n2481), .A2(n2268), .ZN(n3668) );
  NAND2_X1 U3086 ( .A1(n3668), .A2(n3793), .ZN(n3691) );
  NAND2_X1 U3087 ( .A1(n3031), .A2(n2515), .ZN(n2536) );
  OR2_X1 U3088 ( .A1(n2536), .A2(n2535), .ZN(n2541) );
  NAND2_X1 U3089 ( .A1(n2955), .A2(n2956), .ZN(n2957) );
  AOI21_X1 U3090 ( .B1(n4285), .B2(n3862), .A(n3864), .ZN(n4271) );
  AOI21_X1 U3091 ( .B1(n4190), .B2(n2764), .A(n2763), .ZN(n4171) );
  AND2_X1 U3092 ( .A1(n2953), .A2(n2952), .ZN(n2483) );
  OR2_X1 U3093 ( .A1(n4135), .A2(n4515), .ZN(n2485) );
  OR2_X1 U3094 ( .A1(n4141), .A2(n4515), .ZN(n2486) );
  AND2_X2 U3095 ( .A1(n2893), .A2(n3122), .ZN(n4704) );
  NAND2_X1 U3096 ( .A1(n2893), .A2(n2985), .ZN(n4713) );
  AND3_X1 U3097 ( .A1(n2732), .A2(n2731), .A3(n2730), .ZN(n4545) );
  OR2_X1 U3098 ( .A1(n4436), .A2(n4530), .ZN(n2487) );
  OR2_X1 U3099 ( .A1(n4141), .A2(n4458), .ZN(n2489) );
  INV_X1 U3100 ( .A(REG3_REG_13__SCAN_IN), .ZN(n2659) );
  INV_X1 U3101 ( .A(REG3_REG_9__SCAN_IN), .ZN(n2613) );
  OR2_X1 U3102 ( .A1(n4131), .A2(n3686), .ZN(n2490) );
  OR2_X1 U3103 ( .A1(n4135), .A2(n4458), .ZN(n2491) );
  AND2_X1 U3104 ( .A1(n2553), .A2(n2552), .ZN(n2492) );
  INV_X1 U3105 ( .A(n3016), .ZN(n2866) );
  INV_X1 U3106 ( .A(n4327), .ZN(n3875) );
  NOR2_X2 U3107 ( .A1(n2921), .A2(n2920), .ZN(U4043) );
  INV_X1 U3108 ( .A(n2809), .ZN(n4356) );
  NAND2_X1 U3109 ( .A1(n3905), .A2(n3902), .ZN(n2809) );
  INV_X1 U3110 ( .A(IR_REG_19__SCAN_IN), .ZN(n2794) );
  OR2_X1 U3111 ( .A1(n4510), .A2(n4509), .ZN(U3499) );
  AND2_X1 U3112 ( .A1(n2937), .A2(n2488), .ZN(n2496) );
  INV_X1 U3113 ( .A(n3628), .ZN(n3678) );
  NAND2_X1 U3114 ( .A1(n2794), .A2(n2802), .ZN(n2795) );
  INV_X1 U3115 ( .A(IR_REG_16__SCAN_IN), .ZN(n2713) );
  INV_X1 U3116 ( .A(IR_REG_17__SCAN_IN), .ZN(n4844) );
  INV_X1 U3117 ( .A(REG3_REG_24__SCAN_IN), .ZN(n4973) );
  NAND2_X1 U3118 ( .A1(n2936), .A2(n2496), .ZN(n3079) );
  AND2_X1 U3119 ( .A1(n3178), .A2(n3215), .ZN(n3250) );
  OAI22_X1 U3120 ( .A1(n2947), .A2(n3678), .B1(n3677), .B2(n2949), .ZN(n2948)
         );
  INV_X1 U3121 ( .A(REG3_REG_8__SCAN_IN), .ZN(n5057) );
  OR2_X1 U3122 ( .A1(n2660), .A2(n2659), .ZN(n2679) );
  INV_X1 U3123 ( .A(REG3_REG_17__SCAN_IN), .ZN(n2708) );
  INV_X1 U3124 ( .A(n3674), .ZN(n3665) );
  OR2_X1 U3125 ( .A1(n2767), .A2(n2765), .ZN(n2776) );
  INV_X1 U3126 ( .A(n3078), .ZN(n3082) );
  NAND2_X1 U3127 ( .A1(n4325), .A2(n4346), .ZN(n2725) );
  INV_X1 U3128 ( .A(n4384), .ZN(n4166) );
  AND2_X1 U3129 ( .A1(n2627), .A2(REG3_REG_10__SCAN_IN), .ZN(n2635) );
  OAI22_X1 U3130 ( .A1(n3691), .A2(n3692), .B1(n3673), .B2(n3672), .ZN(n3682)
         );
  INV_X1 U3131 ( .A(REG3_REG_21__SCAN_IN), .ZN(n3737) );
  INV_X1 U3132 ( .A(n3303), .ZN(n3249) );
  INV_X1 U3133 ( .A(n3182), .ZN(n3215) );
  INV_X1 U3134 ( .A(REG3_REG_20__SCAN_IN), .ZN(n4815) );
  NOR2_X1 U3135 ( .A1(n2709), .A2(n2708), .ZN(n2718) );
  AND2_X1 U3136 ( .A1(n2776), .A2(n2768), .ZN(n4185) );
  INV_X1 U3137 ( .A(n4064), .ZN(n4043) );
  INV_X1 U3138 ( .A(REG3_REG_16__SCAN_IN), .ZN(n5067) );
  INV_X1 U3139 ( .A(n4177), .ZN(n4146) );
  AND2_X1 U3140 ( .A1(n4131), .A2(n4143), .ZN(n3839) );
  INV_X1 U3141 ( .A(n4178), .ZN(n4210) );
  AND2_X1 U3142 ( .A1(n3931), .A2(n3933), .ZN(n3856) );
  AND2_X1 U3143 ( .A1(n4518), .A2(n3976), .ZN(n3042) );
  OR2_X1 U3144 ( .A1(n3035), .A2(D_REG_0__SCAN_IN), .ZN(n2888) );
  INV_X1 U3145 ( .A(REG0_REG_29__SCAN_IN), .ZN(n2910) );
  INV_X1 U3146 ( .A(n4362), .ZN(n4293) );
  NAND2_X1 U3147 ( .A1(n3042), .A2(n3083), .ZN(n4435) );
  AND2_X1 U31480 ( .A1(n2842), .A2(n3845), .ZN(n4366) );
  NAND2_X1 U31490 ( .A1(n2806), .A2(n4116), .ZN(n4298) );
  INV_X1 U3150 ( .A(IR_REG_7__SCAN_IN), .ZN(n2598) );
  OR2_X1 U3151 ( .A1(n3005), .A2(n3004), .ZN(n4546) );
  NOR2_X1 U3152 ( .A1(n2742), .A2(n3737), .ZN(n2743) );
  AND2_X1 U3153 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n2571) );
  INV_X1 U3154 ( .A(n4519), .ZN(n4116) );
  INV_X1 U3155 ( .A(n4666), .ZN(n2920) );
  XNOR2_X1 U3156 ( .A(n2658), .B(IR_REG_12__SCAN_IN), .ZN(n4064) );
  INV_X1 U3157 ( .A(n4521), .ZN(n4073) );
  AND2_X1 U3158 ( .A1(n4006), .A2(n4001), .ZN(n4637) );
  AND2_X1 U3159 ( .A1(n2235), .A2(DATAI_29_), .ZN(n4133) );
  INV_X1 U3160 ( .A(n4435), .ZN(n4291) );
  INV_X1 U3161 ( .A(n4353), .ZN(n4273) );
  AND2_X1 U3162 ( .A1(n3042), .A2(n3046), .ZN(n4362) );
  NAND2_X1 U3163 ( .A1(n3126), .A2(n3963), .ZN(n4678) );
  AND2_X1 U3164 ( .A1(n2888), .A2(n3038), .ZN(n2985) );
  NAND2_X1 U3165 ( .A1(n2235), .A2(DATAI_27_), .ZN(n4384) );
  INV_X1 U3166 ( .A(n4218), .ZN(n4399) );
  INV_X1 U3167 ( .A(n3478), .ZN(n3560) );
  INV_X1 U3168 ( .A(n2890), .ZN(n3446) );
  AND2_X1 U3169 ( .A1(n3129), .A2(n2922), .ZN(n4690) );
  INV_X1 U3170 ( .A(n3118), .ZN(n3034) );
  INV_X1 U3171 ( .A(n2633), .ZN(n2641) );
  AND2_X1 U3172 ( .A1(n3045), .A2(n3043), .ZN(n4636) );
  AND2_X1 U3173 ( .A1(n2998), .A2(n3111), .ZN(n4563) );
  INV_X1 U3174 ( .A(n4131), .ZN(n4157) );
  INV_X1 U3175 ( .A(n4545), .ZN(n4339) );
  NAND2_X1 U3176 ( .A1(n4006), .A2(n3046), .ZN(n4642) );
  INV_X1 U3177 ( .A(n4593), .ZN(n4630) );
  NAND2_X1 U3178 ( .A1(n4654), .A2(n3223), .ZN(n4353) );
  AND2_X2 U3179 ( .A1(n3123), .A2(n4651), .ZN(n4663) );
  OR2_X1 U3180 ( .A1(n4347), .A2(n4678), .ZN(n4328) );
  NAND2_X1 U3181 ( .A1(n4716), .A2(n4701), .ZN(n4458) );
  INV_X2 U3182 ( .A(n4713), .ZN(n4716) );
  NAND2_X1 U3183 ( .A1(n4701), .A2(n4704), .ZN(n4515) );
  INV_X1 U3184 ( .A(n4704), .ZN(n4702) );
  INV_X1 U3185 ( .A(n4664), .ZN(n4665) );
  AND2_X1 U3186 ( .A1(n2675), .A2(n2674), .ZN(n4521) );
  INV_X1 U3187 ( .A(IR_REG_2__SCAN_IN), .ZN(n2497) );
  NAND3_X1 U3188 ( .A1(n2669), .A2(n2498), .A3(n2668), .ZN(n2500) );
  NAND4_X1 U3189 ( .A1(n2598), .A2(n4826), .A3(n4866), .A4(n2499), .ZN(n2667)
         );
  NAND2_X1 U3190 ( .A1(n2508), .A2(n2482), .ZN(n2503) );
  NAND2_X1 U3191 ( .A1(n2571), .A2(REG3_REG_5__SCAN_IN), .ZN(n2583) );
  NOR2_X1 U3192 ( .A1(n2583), .A2(n3060), .ZN(n2591) );
  NAND2_X1 U3193 ( .A1(n2591), .A2(REG3_REG_7__SCAN_IN), .ZN(n2603) );
  NAND2_X1 U3194 ( .A1(n2635), .A2(REG3_REG_11__SCAN_IN), .ZN(n2651) );
  NAND2_X1 U3195 ( .A1(n2690), .A2(REG3_REG_15__SCAN_IN), .ZN(n2700) );
  NAND2_X1 U3196 ( .A1(n2750), .A2(n4973), .ZN(n2506) );
  NAND2_X1 U3197 ( .A1(n2767), .A2(n2506), .ZN(n4214) );
  INV_X1 U3198 ( .A(IR_REG_29__SCAN_IN), .ZN(n2509) );
  OAI21_X1 U3199 ( .B1(n2850), .B2(n2863), .A(IR_REG_29__SCAN_IN), .ZN(n2511)
         );
  INV_X1 U3200 ( .A(n3022), .ZN(n2512) );
  INV_X1 U3201 ( .A(n2515), .ZN(n4517) );
  OR2_X1 U3202 ( .A1(n4214), .A2(n2843), .ZN(n2521) );
  INV_X1 U3203 ( .A(REG2_REG_24__SCAN_IN), .ZN(n4215) );
  NAND2_X1 U3204 ( .A1(n2538), .A2(REG0_REG_24__SCAN_IN), .ZN(n2518) );
  NAND2_X1 U3205 ( .A1(n2537), .A2(REG1_REG_24__SCAN_IN), .ZN(n2517) );
  OAI211_X1 U3206 ( .C1(n4215), .C2(n2562), .A(n2518), .B(n2517), .ZN(n2519)
         );
  INV_X1 U3207 ( .A(n2519), .ZN(n2520) );
  AND2_X1 U3208 ( .A1(n4218), .A2(n3983), .ZN(n2756) );
  NAND2_X1 U3209 ( .A1(n2234), .A2(DATAI_22_), .ZN(n3787) );
  NOR2_X1 U32100 ( .A1(n2743), .A2(REG3_REG_22__SCAN_IN), .ZN(n2522) );
  OR2_X1 U32110 ( .A1(n2748), .A2(n2522), .ZN(n4261) );
  INV_X1 U32120 ( .A(REG2_REG_22__SCAN_IN), .ZN(n2525) );
  NAND2_X1 U32130 ( .A1(n2538), .A2(REG0_REG_22__SCAN_IN), .ZN(n2524) );
  NAND2_X1 U32140 ( .A1(n2537), .A2(REG1_REG_22__SCAN_IN), .ZN(n2523) );
  OAI211_X1 U32150 ( .C1(n2525), .C2(n2562), .A(n2524), .B(n2523), .ZN(n2526)
         );
  INV_X1 U32160 ( .A(n2526), .ZN(n2527) );
  NAND2_X1 U32170 ( .A1(n2528), .A2(REG2_REG_1__SCAN_IN), .ZN(n2533) );
  NAND2_X1 U32180 ( .A1(n2529), .A2(REG3_REG_1__SCAN_IN), .ZN(n2532) );
  NAND2_X1 U32190 ( .A1(n2537), .A2(REG1_REG_1__SCAN_IN), .ZN(n2531) );
  NAND2_X1 U32200 ( .A1(n2538), .A2(REG0_REG_1__SCAN_IN), .ZN(n2530) );
  NAND2_X1 U32210 ( .A1(n2543), .A2(n3191), .ZN(n3899) );
  NAND2_X1 U32220 ( .A1(n3899), .A2(n3901), .ZN(n2807) );
  NAND2_X1 U32230 ( .A1(n2529), .A2(REG3_REG_0__SCAN_IN), .ZN(n2542) );
  INV_X1 U32240 ( .A(REG2_REG_0__SCAN_IN), .ZN(n2535) );
  NAND2_X1 U32250 ( .A1(n2537), .A2(REG1_REG_0__SCAN_IN), .ZN(n2540) );
  NAND2_X1 U32260 ( .A1(n2538), .A2(REG0_REG_0__SCAN_IN), .ZN(n2539) );
  INV_X1 U32270 ( .A(n2933), .ZN(n3153) );
  AND2_X1 U32280 ( .A1(n2933), .A2(n3127), .ZN(n3193) );
  NAND2_X1 U32290 ( .A1(n2807), .A2(n3193), .ZN(n3195) );
  NAND2_X1 U32300 ( .A1(n2543), .A2(n3197), .ZN(n2544) );
  NAND2_X1 U32310 ( .A1(n3195), .A2(n2544), .ZN(n4357) );
  NAND2_X1 U32320 ( .A1(n2529), .A2(REG3_REG_2__SCAN_IN), .ZN(n2548) );
  NAND2_X1 U32330 ( .A1(n2528), .A2(REG2_REG_2__SCAN_IN), .ZN(n2547) );
  NAND2_X1 U32340 ( .A1(n2537), .A2(REG1_REG_2__SCAN_IN), .ZN(n2546) );
  NAND2_X1 U32350 ( .A1(n2538), .A2(REG0_REG_2__SCAN_IN), .ZN(n2545) );
  OR2_X1 U32360 ( .A1(n2549), .A2(n2863), .ZN(n2550) );
  XNOR2_X2 U32370 ( .A(n2550), .B(IR_REG_2__SCAN_IN), .ZN(n4022) );
  MUX2_X1 U32380 ( .A(n4022), .B(DATAI_2_), .S(n2234), .Z(n4369) );
  INV_X1 U32390 ( .A(n4369), .ZN(n4360) );
  NAND2_X1 U32400 ( .A1(n4000), .A2(n4360), .ZN(n3905) );
  NAND2_X1 U32410 ( .A1(n3228), .A2(n4369), .ZN(n3902) );
  NAND2_X1 U32420 ( .A1(n3228), .A2(n4360), .ZN(n2551) );
  NAND2_X1 U32430 ( .A1(n2538), .A2(REG0_REG_3__SCAN_IN), .ZN(n2553) );
  NAND2_X1 U32440 ( .A1(n2528), .A2(REG2_REG_3__SCAN_IN), .ZN(n2552) );
  NAND2_X1 U32450 ( .A1(n2537), .A2(REG1_REG_3__SCAN_IN), .ZN(n2555) );
  INV_X1 U32460 ( .A(REG3_REG_3__SCAN_IN), .ZN(n4828) );
  NAND2_X1 U32470 ( .A1(n2529), .A2(n4828), .ZN(n2554) );
  NAND2_X1 U32480 ( .A1(n2556), .A2(IR_REG_31__SCAN_IN), .ZN(n2558) );
  NAND2_X1 U32490 ( .A1(n2558), .A2(n2557), .ZN(n2567) );
  OR2_X1 U32500 ( .A1(n2558), .A2(n2557), .ZN(n2559) );
  MUX2_X1 U32510 ( .A(n4527), .B(DATAI_3_), .S(n2235), .Z(n3231) );
  NOR2_X1 U32520 ( .A1(n4363), .A2(n3231), .ZN(n2560) );
  NOR2_X1 U32530 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n2561) );
  NOR2_X1 U32540 ( .A1(n2571), .A2(n2561), .ZN(n3211) );
  NAND2_X1 U32550 ( .A1(n2529), .A2(n3211), .ZN(n2566) );
  NAND2_X1 U32560 ( .A1(n2528), .A2(REG2_REG_4__SCAN_IN), .ZN(n2565) );
  NAND2_X1 U32570 ( .A1(n2538), .A2(REG0_REG_4__SCAN_IN), .ZN(n2564) );
  NAND2_X1 U32580 ( .A1(n2537), .A2(REG1_REG_4__SCAN_IN), .ZN(n2563) );
  NAND2_X1 U32590 ( .A1(n2567), .A2(IR_REG_31__SCAN_IN), .ZN(n2568) );
  MUX2_X1 U32600 ( .A(n4526), .B(DATAI_4_), .S(n2235), .Z(n3182) );
  NAND2_X1 U32610 ( .A1(n3305), .A2(n3182), .ZN(n3908) );
  NAND2_X1 U32620 ( .A1(n3999), .A2(n3215), .ZN(n3911) );
  NAND2_X1 U32630 ( .A1(n3908), .A2(n3911), .ZN(n3180) );
  NAND2_X1 U32640 ( .A1(n3179), .A2(n3180), .ZN(n2570) );
  NAND2_X1 U32650 ( .A1(n3999), .A2(n3182), .ZN(n2569) );
  OAI21_X1 U32660 ( .B1(n2571), .B2(REG3_REG_5__SCAN_IN), .A(n2583), .ZN(n3300) );
  INV_X1 U32670 ( .A(n3300), .ZN(n2572) );
  NAND2_X1 U32680 ( .A1(n2529), .A2(n2572), .ZN(n2576) );
  NAND2_X1 U32690 ( .A1(n2528), .A2(REG2_REG_5__SCAN_IN), .ZN(n2575) );
  NAND2_X1 U32700 ( .A1(n2538), .A2(REG0_REG_5__SCAN_IN), .ZN(n2574) );
  NAND2_X1 U32710 ( .A1(n2537), .A2(REG1_REG_5__SCAN_IN), .ZN(n2573) );
  NAND4_X1 U32720 ( .A1(n2576), .A2(n2575), .A3(n2574), .A4(n2573), .ZN(n3998)
         );
  NAND2_X1 U32730 ( .A1(n2577), .A2(IR_REG_31__SCAN_IN), .ZN(n2579) );
  INV_X1 U32740 ( .A(IR_REG_5__SCAN_IN), .ZN(n2578) );
  MUX2_X1 U32750 ( .A(n2579), .B(IR_REG_31__SCAN_IN), .S(n2578), .Z(n2581) );
  NOR2_X1 U32760 ( .A1(n2577), .A2(IR_REG_5__SCAN_IN), .ZN(n2597) );
  INV_X1 U32770 ( .A(n2597), .ZN(n2580) );
  MUX2_X1 U32780 ( .A(n4525), .B(DATAI_5_), .S(n2235), .Z(n3303) );
  AND2_X1 U32790 ( .A1(n3998), .A2(n3303), .ZN(n2582) );
  AND2_X1 U32800 ( .A1(n2583), .A2(n3060), .ZN(n2584) );
  NOR2_X1 U32810 ( .A1(n2591), .A2(n2584), .ZN(n3321) );
  NAND2_X1 U32820 ( .A1(n2529), .A2(n3321), .ZN(n2588) );
  NAND2_X1 U32830 ( .A1(n2528), .A2(REG2_REG_6__SCAN_IN), .ZN(n2587) );
  NAND2_X1 U32840 ( .A1(n2538), .A2(REG0_REG_6__SCAN_IN), .ZN(n2586) );
  NAND2_X1 U32850 ( .A1(n2537), .A2(REG1_REG_6__SCAN_IN), .ZN(n2585) );
  NAND4_X1 U32860 ( .A1(n2588), .A2(n2587), .A3(n2586), .A4(n2585), .ZN(n3997)
         );
  OR2_X1 U32870 ( .A1(n2597), .A2(n2863), .ZN(n2589) );
  XNOR2_X1 U32880 ( .A(n2589), .B(IR_REG_6__SCAN_IN), .ZN(n4524) );
  MUX2_X1 U32890 ( .A(n4524), .B(DATAI_6_), .S(n2235), .Z(n3272) );
  NAND2_X1 U32900 ( .A1(n3997), .A2(n3272), .ZN(n2590) );
  OR2_X1 U32910 ( .A1(n2591), .A2(REG3_REG_7__SCAN_IN), .ZN(n2592) );
  AND2_X1 U32920 ( .A1(n2603), .A2(n2592), .ZN(n3572) );
  NAND2_X1 U32930 ( .A1(n2529), .A2(n3572), .ZN(n2596) );
  NAND2_X1 U32940 ( .A1(n2528), .A2(REG2_REG_7__SCAN_IN), .ZN(n2595) );
  NAND2_X1 U32950 ( .A1(n2538), .A2(REG0_REG_7__SCAN_IN), .ZN(n2594) );
  NAND2_X1 U32960 ( .A1(n2537), .A2(REG1_REG_7__SCAN_IN), .ZN(n2593) );
  NAND2_X1 U32970 ( .A1(n2597), .A2(n4826), .ZN(n2620) );
  NAND2_X1 U32980 ( .A1(n2620), .A2(IR_REG_31__SCAN_IN), .ZN(n2599) );
  NAND2_X1 U32990 ( .A1(n2599), .A2(n2598), .ZN(n2609) );
  OR2_X1 U33000 ( .A1(n2599), .A2(n2598), .ZN(n2600) );
  MUX2_X1 U33010 ( .A(n4523), .B(DATAI_7_), .S(n2235), .Z(n3291) );
  NAND2_X1 U33020 ( .A1(n3368), .A2(n3291), .ZN(n2814) );
  INV_X1 U33030 ( .A(n3291), .ZN(n3570) );
  NAND2_X1 U33040 ( .A1(n3995), .A2(n3570), .ZN(n3916) );
  NAND2_X1 U33050 ( .A1(n3995), .A2(n3291), .ZN(n2601) );
  NAND2_X1 U33060 ( .A1(n2602), .A2(n2601), .ZN(n3324) );
  NAND2_X1 U33070 ( .A1(n2603), .A2(n5057), .ZN(n2604) );
  AND2_X1 U33080 ( .A1(n2614), .A2(n2604), .ZN(n3363) );
  NAND2_X1 U33090 ( .A1(n2529), .A2(n3363), .ZN(n2608) );
  NAND2_X1 U33100 ( .A1(n2528), .A2(REG2_REG_8__SCAN_IN), .ZN(n2607) );
  NAND2_X1 U33110 ( .A1(n2538), .A2(REG0_REG_8__SCAN_IN), .ZN(n2606) );
  NAND2_X1 U33120 ( .A1(n2537), .A2(REG1_REG_8__SCAN_IN), .ZN(n2605) );
  NAND4_X1 U33130 ( .A1(n2608), .A2(n2607), .A3(n2606), .A4(n2605), .ZN(n3994)
         );
  NAND2_X1 U33140 ( .A1(n2609), .A2(IR_REG_31__SCAN_IN), .ZN(n2610) );
  XNOR2_X1 U33150 ( .A(n2610), .B(IR_REG_8__SCAN_IN), .ZN(n3161) );
  MUX2_X1 U33160 ( .A(n3161), .B(DATAI_8_), .S(n2235), .Z(n3332) );
  AND2_X1 U33170 ( .A1(n3994), .A2(n3332), .ZN(n2612) );
  INV_X1 U33180 ( .A(n3994), .ZN(n3353) );
  INV_X1 U33190 ( .A(n3332), .ZN(n3369) );
  NAND2_X1 U33200 ( .A1(n3353), .A2(n3369), .ZN(n2611) );
  AND2_X1 U33210 ( .A1(n2614), .A2(n2613), .ZN(n2615) );
  OR2_X1 U33220 ( .A1(n2615), .A2(n2627), .ZN(n3345) );
  INV_X1 U33230 ( .A(n3345), .ZN(n3381) );
  NAND2_X1 U33240 ( .A1(n2529), .A2(n3381), .ZN(n2619) );
  NAND2_X1 U33250 ( .A1(n2528), .A2(REG2_REG_9__SCAN_IN), .ZN(n2618) );
  NAND2_X1 U33260 ( .A1(n2537), .A2(REG1_REG_9__SCAN_IN), .ZN(n2617) );
  NAND2_X1 U33270 ( .A1(n2538), .A2(REG0_REG_9__SCAN_IN), .ZN(n2616) );
  NAND4_X1 U33280 ( .A1(n2619), .A2(n2618), .A3(n2617), .A4(n2616), .ZN(n3993)
         );
  NAND2_X1 U33290 ( .A1(n2623), .A2(IR_REG_31__SCAN_IN), .ZN(n2621) );
  MUX2_X1 U33300 ( .A(n2621), .B(IR_REG_31__SCAN_IN), .S(n2624), .Z(n2622) );
  INV_X1 U33310 ( .A(n2622), .ZN(n2626) );
  INV_X1 U33320 ( .A(n2623), .ZN(n2625) );
  NAND2_X1 U33330 ( .A1(n2625), .A2(n2624), .ZN(n2633) );
  MUX2_X1 U33340 ( .A(n4567), .B(DATAI_9_), .S(n2235), .Z(n3347) );
  NOR2_X1 U33350 ( .A1(n2627), .A2(REG3_REG_10__SCAN_IN), .ZN(n2628) );
  OR2_X1 U33360 ( .A1(n2635), .A2(n2628), .ZN(n2999) );
  INV_X1 U33370 ( .A(n2999), .ZN(n4644) );
  NAND2_X1 U33380 ( .A1(n2529), .A2(n4644), .ZN(n2632) );
  NAND2_X1 U33390 ( .A1(n2528), .A2(REG2_REG_10__SCAN_IN), .ZN(n2631) );
  NAND2_X1 U33400 ( .A1(n2537), .A2(REG1_REG_10__SCAN_IN), .ZN(n2630) );
  NAND2_X1 U33410 ( .A1(n2538), .A2(REG0_REG_10__SCAN_IN), .ZN(n2629) );
  NAND4_X1 U33420 ( .A1(n2632), .A2(n2631), .A3(n2630), .A4(n2629), .ZN(n3992)
         );
  NAND2_X1 U33430 ( .A1(n2633), .A2(IR_REG_31__SCAN_IN), .ZN(n2634) );
  XNOR2_X1 U33440 ( .A(n2634), .B(IR_REG_10__SCAN_IN), .ZN(n4049) );
  MUX2_X1 U33450 ( .A(n4049), .B(DATAI_10_), .S(n2235), .Z(n2890) );
  AND2_X1 U33460 ( .A1(n3992), .A2(n2890), .ZN(n3384) );
  OR2_X1 U33470 ( .A1(n2635), .A2(REG3_REG_11__SCAN_IN), .ZN(n2636) );
  AND2_X1 U33480 ( .A1(n2651), .A2(n2636), .ZN(n3424) );
  NAND2_X1 U33490 ( .A1(n2529), .A2(n3424), .ZN(n2640) );
  NAND2_X1 U33500 ( .A1(n2528), .A2(REG2_REG_11__SCAN_IN), .ZN(n2639) );
  NAND2_X1 U33510 ( .A1(n2538), .A2(REG0_REG_11__SCAN_IN), .ZN(n2638) );
  NAND2_X1 U33520 ( .A1(n2537), .A2(REG1_REG_11__SCAN_IN), .ZN(n2637) );
  NAND2_X1 U3353 ( .A1(n2641), .A2(n2453), .ZN(n2642) );
  NAND2_X1 U33540 ( .A1(n2642), .A2(IR_REG_31__SCAN_IN), .ZN(n2643) );
  NAND2_X1 U3355 ( .A1(n2643), .A2(n4866), .ZN(n2657) );
  OR2_X1 U3356 ( .A1(n2643), .A2(n4866), .ZN(n2644) );
  MUX2_X1 U3357 ( .A(n4522), .B(DATAI_11_), .S(n2235), .Z(n3417) );
  INV_X1 U3358 ( .A(n3417), .ZN(n3422) );
  NAND2_X1 U3359 ( .A1(n3538), .A2(n3422), .ZN(n2646) );
  INV_X1 U3360 ( .A(n2646), .ZN(n2645) );
  NAND2_X1 U3361 ( .A1(n3538), .A2(n3417), .ZN(n3399) );
  NAND2_X1 U3362 ( .A1(n3991), .A2(n3422), .ZN(n3401) );
  NAND2_X1 U3363 ( .A1(n3399), .A2(n3401), .ZN(n3387) );
  NOR2_X1 U3364 ( .A1(n2645), .A2(n3387), .ZN(n2648) );
  OR2_X1 U3365 ( .A1(n3384), .A2(n2648), .ZN(n2649) );
  NAND2_X1 U3366 ( .A1(n3390), .A2(n3446), .ZN(n3385) );
  AND2_X1 U3367 ( .A1(n3385), .A2(n2646), .ZN(n2647) );
  NAND2_X1 U3368 ( .A1(n2651), .A2(n2650), .ZN(n2652) );
  AND2_X1 U3369 ( .A1(n2660), .A2(n2652), .ZN(n3407) );
  NAND2_X1 U3370 ( .A1(n2529), .A2(n3407), .ZN(n2656) );
  NAND2_X1 U3371 ( .A1(n2528), .A2(REG2_REG_12__SCAN_IN), .ZN(n2655) );
  NAND2_X1 U3372 ( .A1(n2538), .A2(REG0_REG_12__SCAN_IN), .ZN(n2654) );
  NAND2_X1 U3373 ( .A1(n2537), .A2(REG1_REG_12__SCAN_IN), .ZN(n2653) );
  NAND4_X1 U3374 ( .A1(n2656), .A2(n2655), .A3(n2654), .A4(n2653), .ZN(n3990)
         );
  NAND2_X1 U3375 ( .A1(n2657), .A2(IR_REG_31__SCAN_IN), .ZN(n2658) );
  MUX2_X1 U3376 ( .A(n4064), .B(DATAI_12_), .S(n2234), .Z(n3525) );
  INV_X1 U3377 ( .A(n3990), .ZN(n2821) );
  NAND2_X1 U3378 ( .A1(n2660), .A2(n2659), .ZN(n2661) );
  NAND2_X1 U3379 ( .A1(n2679), .A2(n2661), .ZN(n3490) );
  INV_X1 U3380 ( .A(n3490), .ZN(n3562) );
  NAND2_X1 U3381 ( .A1(n2529), .A2(n3562), .ZN(n2665) );
  NAND2_X1 U3382 ( .A1(n2528), .A2(REG2_REG_13__SCAN_IN), .ZN(n2664) );
  NAND2_X1 U3383 ( .A1(n2537), .A2(REG1_REG_13__SCAN_IN), .ZN(n2663) );
  NAND2_X1 U3384 ( .A1(n2538), .A2(REG0_REG_13__SCAN_IN), .ZN(n2662) );
  NAND4_X1 U3385 ( .A1(n2665), .A2(n2664), .A3(n2663), .A4(n2662), .ZN(n3989)
         );
  INV_X1 U3386 ( .A(n2667), .ZN(n2670) );
  NAND4_X1 U3387 ( .A1(n2666), .A2(n2670), .A3(n2669), .A4(n2668), .ZN(n2671)
         );
  NAND2_X1 U3388 ( .A1(n2671), .A2(IR_REG_31__SCAN_IN), .ZN(n2672) );
  MUX2_X1 U3389 ( .A(IR_REG_31__SCAN_IN), .B(n2672), .S(IR_REG_13__SCAN_IN), 
        .Z(n2675) );
  INV_X1 U3390 ( .A(n2673), .ZN(n2674) );
  MUX2_X1 U3391 ( .A(n4521), .B(DATAI_13_), .S(n2235), .Z(n3478) );
  AND2_X1 U3392 ( .A1(n3989), .A2(n3478), .ZN(n2677) );
  NAND2_X1 U3393 ( .A1(n3704), .A2(n3560), .ZN(n2676) );
  AND2_X1 U3394 ( .A1(n2679), .A2(n2678), .ZN(n2680) );
  NOR2_X1 U3395 ( .A1(n2690), .A2(n2680), .ZN(n3436) );
  NAND2_X1 U3396 ( .A1(n2529), .A2(n3436), .ZN(n2684) );
  NAND2_X1 U3397 ( .A1(n2528), .A2(REG2_REG_14__SCAN_IN), .ZN(n2683) );
  NAND2_X1 U3398 ( .A1(n2538), .A2(REG0_REG_14__SCAN_IN), .ZN(n2682) );
  NAND2_X1 U3399 ( .A1(n2537), .A2(REG1_REG_14__SCAN_IN), .ZN(n2681) );
  NOR2_X1 U3400 ( .A1(n2673), .A2(n2863), .ZN(n2685) );
  MUX2_X1 U3401 ( .A(n2863), .B(n2685), .S(IR_REG_14__SCAN_IN), .Z(n2686) );
  INV_X1 U3402 ( .A(n2686), .ZN(n2688) );
  AND2_X1 U3403 ( .A1(n2688), .A2(n2687), .ZN(n4093) );
  MUX2_X1 U3404 ( .A(n4093), .B(DATAI_14_), .S(n2235), .Z(n3435) );
  NAND2_X1 U3405 ( .A1(n3579), .A2(n3435), .ZN(n3816) );
  INV_X1 U3406 ( .A(n3579), .ZN(n3988) );
  INV_X1 U3407 ( .A(n3435), .ZN(n3705) );
  NAND2_X1 U3408 ( .A1(n3988), .A2(n3705), .ZN(n3817) );
  NAND2_X1 U3409 ( .A1(n3816), .A2(n3817), .ZN(n3428) );
  NAND2_X1 U3410 ( .A1(n3579), .A2(n3705), .ZN(n2689) );
  OR2_X1 U3411 ( .A1(n2690), .A2(REG3_REG_15__SCAN_IN), .ZN(n2691) );
  AND2_X1 U3412 ( .A1(n2691), .A2(n2700), .ZN(n3810) );
  NAND2_X1 U3413 ( .A1(n2529), .A2(n3810), .ZN(n2695) );
  NAND2_X1 U3414 ( .A1(n2528), .A2(REG2_REG_15__SCAN_IN), .ZN(n2694) );
  NAND2_X1 U3415 ( .A1(n2538), .A2(REG0_REG_15__SCAN_IN), .ZN(n2693) );
  NAND2_X1 U3416 ( .A1(n2537), .A2(REG1_REG_15__SCAN_IN), .ZN(n2692) );
  NAND4_X1 U3417 ( .A1(n2695), .A2(n2694), .A3(n2693), .A4(n2692), .ZN(n3987)
         );
  NAND2_X1 U3418 ( .A1(n2687), .A2(IR_REG_31__SCAN_IN), .ZN(n2696) );
  NAND2_X1 U3419 ( .A1(n2696), .A2(n2480), .ZN(n2706) );
  OR2_X1 U3420 ( .A1(n2696), .A2(n2480), .ZN(n2697) );
  MUX2_X1 U3421 ( .A(n4096), .B(DATAI_15_), .S(n2235), .Z(n3584) );
  NOR2_X1 U3422 ( .A1(n3987), .A2(n3584), .ZN(n2699) );
  NAND2_X1 U3423 ( .A1(n3987), .A2(n3584), .ZN(n2698) );
  AOI22_X1 U3424 ( .A1(n2528), .A2(REG2_REG_16__SCAN_IN), .B1(n2538), .B2(
        REG0_REG_16__SCAN_IN), .ZN(n2705) );
  NAND2_X1 U3425 ( .A1(n2700), .A2(n5067), .ZN(n2701) );
  NAND2_X1 U3426 ( .A1(n2709), .A2(n2701), .ZN(n4543) );
  NAND2_X1 U3427 ( .A1(n2537), .A2(REG1_REG_16__SCAN_IN), .ZN(n2702) );
  OAI21_X1 U3428 ( .B1(n4543), .B2(n2843), .A(n2702), .ZN(n2703) );
  INV_X1 U3429 ( .A(n2703), .ZN(n2704) );
  NAND2_X1 U3430 ( .A1(n2706), .A2(IR_REG_31__SCAN_IN), .ZN(n2707) );
  XNOR2_X1 U3431 ( .A(n2707), .B(IR_REG_16__SCAN_IN), .ZN(n4668) );
  MUX2_X1 U3432 ( .A(n4668), .B(DATAI_16_), .S(n2235), .Z(n3496) );
  NAND2_X1 U3433 ( .A1(n4436), .A2(n3496), .ZN(n3943) );
  NAND2_X1 U3434 ( .A1(n3986), .A2(n4530), .ZN(n3821) );
  NAND2_X1 U3435 ( .A1(n3943), .A2(n3821), .ZN(n3502) );
  NAND2_X1 U3436 ( .A1(n3501), .A2(n2487), .ZN(n3544) );
  AND2_X1 U3437 ( .A1(n2709), .A2(n2708), .ZN(n2710) );
  NOR2_X1 U3438 ( .A1(n2718), .A2(n2710), .ZN(n3762) );
  AOI22_X1 U3439 ( .A1(n2529), .A2(n3762), .B1(n2537), .B2(
        REG1_REG_17__SCAN_IN), .ZN(n2712) );
  AOI22_X1 U3440 ( .A1(n2528), .A2(REG2_REG_17__SCAN_IN), .B1(n2538), .B2(
        REG0_REG_17__SCAN_IN), .ZN(n2711) );
  NAND2_X1 U3441 ( .A1(n2735), .A2(n2713), .ZN(n2714) );
  NAND2_X1 U3442 ( .A1(n2714), .A2(IR_REG_31__SCAN_IN), .ZN(n2715) );
  MUX2_X1 U3443 ( .A(IR_REG_31__SCAN_IN), .B(n2715), .S(IR_REG_17__SCAN_IN), 
        .Z(n2716) );
  NAND2_X1 U3444 ( .A1(n2735), .A2(n2733), .ZN(n2723) );
  INV_X1 U3445 ( .A(DATAI_17_), .ZN(n4794) );
  MUX2_X1 U3446 ( .A(n4667), .B(n4794), .S(n2235), .Z(n4434) );
  NAND2_X1 U3447 ( .A1(n4533), .A2(n4434), .ZN(n2717) );
  INV_X1 U3448 ( .A(n4434), .ZN(n3598) );
  NOR2_X1 U3449 ( .A1(n2718), .A2(REG3_REG_18__SCAN_IN), .ZN(n2719) );
  OR2_X1 U3450 ( .A1(n2728), .A2(n2719), .ZN(n4562) );
  INV_X1 U3451 ( .A(REG2_REG_18__SCAN_IN), .ZN(n4348) );
  OAI22_X1 U3452 ( .A1(n2843), .A2(n4562), .B1(n2562), .B2(n4348), .ZN(n2720)
         );
  INV_X1 U3453 ( .A(n2720), .ZN(n2722) );
  AOI22_X1 U3454 ( .A1(n2537), .A2(REG1_REG_18__SCAN_IN), .B1(n2538), .B2(
        REG0_REG_18__SCAN_IN), .ZN(n2721) );
  NAND2_X1 U3455 ( .A1(n2723), .A2(IR_REG_31__SCAN_IN), .ZN(n2724) );
  XNOR2_X1 U3456 ( .A(n2724), .B(IR_REG_18__SCAN_IN), .ZN(n4520) );
  MUX2_X1 U3457 ( .A(n4520), .B(DATAI_18_), .S(n2235), .Z(n4558) );
  NAND2_X1 U34580 ( .A1(n4325), .A2(n4558), .ZN(n4317) );
  INV_X1 U34590 ( .A(n4558), .ZN(n4346) );
  NAND2_X1 U3460 ( .A1(n3985), .A2(n4346), .ZN(n4315) );
  NAND2_X1 U3461 ( .A1(n4317), .A2(n4315), .ZN(n4337) );
  NAND2_X1 U3462 ( .A1(n2538), .A2(REG0_REG_19__SCAN_IN), .ZN(n2727) );
  NAND2_X1 U3463 ( .A1(n2537), .A2(REG1_REG_19__SCAN_IN), .ZN(n2726) );
  AND2_X1 U3464 ( .A1(n2727), .A2(n2726), .ZN(n2732) );
  OR2_X1 U3465 ( .A1(n2728), .A2(REG3_REG_19__SCAN_IN), .ZN(n2729) );
  AND2_X1 U3466 ( .A1(n2737), .A2(n2729), .ZN(n3721) );
  NAND2_X1 U34670 ( .A1(n3721), .A2(n2529), .ZN(n2731) );
  NAND2_X1 U3468 ( .A1(n2528), .A2(REG2_REG_19__SCAN_IN), .ZN(n2730) );
  NAND2_X1 U34690 ( .A1(n2735), .A2(n2734), .ZN(n2796) );
  INV_X1 U3470 ( .A(DATAI_19_), .ZN(n4854) );
  MUX2_X1 U34710 ( .A(n4116), .B(n4854), .S(n2235), .Z(n4327) );
  OR2_X1 U3472 ( .A1(n4545), .A2(n4327), .ZN(n2736) );
  NAND2_X1 U34730 ( .A1(n2737), .A2(n4815), .ZN(n2738) );
  NAND2_X1 U3474 ( .A1(n2742), .A2(n2738), .ZN(n4303) );
  AOI22_X1 U34750 ( .A1(n2537), .A2(REG1_REG_20__SCAN_IN), .B1(n2538), .B2(
        REG0_REG_20__SCAN_IN), .ZN(n2740) );
  NAND2_X1 U3476 ( .A1(n2528), .A2(REG2_REG_20__SCAN_IN), .ZN(n2739) );
  OAI211_X1 U34770 ( .C1(n4303), .C2(n2843), .A(n2740), .B(n2739), .ZN(n4322)
         );
  NAND2_X1 U3478 ( .A1(n4322), .A2(n4290), .ZN(n3862) );
  NOR2_X1 U34790 ( .A1(n4322), .A2(n4290), .ZN(n3864) );
  AND2_X1 U3480 ( .A1(n2742), .A2(n3737), .ZN(n2744) );
  OR2_X1 U34810 ( .A1(n2744), .A2(n2743), .ZN(n4274) );
  AOI22_X1 U3482 ( .A1(n2537), .A2(REG1_REG_21__SCAN_IN), .B1(n2538), .B2(
        REG0_REG_21__SCAN_IN), .ZN(n2746) );
  NAND2_X1 U34830 ( .A1(n2528), .A2(REG2_REG_21__SCAN_IN), .ZN(n2745) );
  OAI211_X1 U3484 ( .C1(n4274), .C2(n2843), .A(n2746), .B(n2745), .ZN(n4258)
         );
  INV_X1 U34850 ( .A(n4258), .ZN(n4294) );
  NOR2_X1 U3486 ( .A1(n4294), .A2(n4415), .ZN(n2747) );
  INV_X1 U34870 ( .A(n4415), .ZN(n4281) );
  OAI22_X1 U3488 ( .A1(n4271), .A2(n2747), .B1(n4281), .B2(n4258), .ZN(n4252)
         );
  OR2_X1 U34890 ( .A1(n4268), .A2(n3787), .ZN(n4236) );
  NAND2_X1 U3490 ( .A1(n4268), .A2(n3787), .ZN(n2835) );
  OR2_X1 U34910 ( .A1(n2748), .A2(REG3_REG_23__SCAN_IN), .ZN(n2749) );
  AND2_X1 U3492 ( .A1(n2750), .A2(n2749), .ZN(n3711) );
  NAND2_X1 U34930 ( .A1(n3711), .A2(n2529), .ZN(n2755) );
  INV_X1 U3494 ( .A(REG2_REG_23__SCAN_IN), .ZN(n4245) );
  NAND2_X1 U34950 ( .A1(n2537), .A2(REG1_REG_23__SCAN_IN), .ZN(n2752) );
  NAND2_X1 U3496 ( .A1(n2538), .A2(REG0_REG_23__SCAN_IN), .ZN(n2751) );
  OAI211_X1 U34970 ( .C1(n4245), .C2(n2562), .A(n2752), .B(n2751), .ZN(n2753)
         );
  INV_X1 U3498 ( .A(n2753), .ZN(n2754) );
  XNOR2_X1 U34990 ( .A(n2767), .B(REG3_REG_25__SCAN_IN), .ZN(n4200) );
  NAND2_X1 U3500 ( .A1(n4200), .A2(n2529), .ZN(n2762) );
  INV_X1 U35010 ( .A(REG2_REG_25__SCAN_IN), .ZN(n2759) );
  NAND2_X1 U3502 ( .A1(n2537), .A2(REG1_REG_25__SCAN_IN), .ZN(n2758) );
  NAND2_X1 U35030 ( .A1(n2538), .A2(REG0_REG_25__SCAN_IN), .ZN(n2757) );
  OAI211_X1 U3504 ( .C1(n2759), .C2(n2562), .A(n2758), .B(n2757), .ZN(n2760)
         );
  INV_X1 U35050 ( .A(n2760), .ZN(n2761) );
  NAND2_X1 U35060 ( .A1(n4210), .A2(n4197), .ZN(n2764) );
  NOR2_X1 U35070 ( .A1(n4210), .A2(n4197), .ZN(n2763) );
  NAND2_X1 U35080 ( .A1(REG3_REG_25__SCAN_IN), .A2(REG3_REG_26__SCAN_IN), .ZN(
        n2765) );
  INV_X1 U35090 ( .A(REG3_REG_25__SCAN_IN), .ZN(n3747) );
  INV_X1 U35100 ( .A(REG3_REG_26__SCAN_IN), .ZN(n2766) );
  OAI21_X1 U35110 ( .B1(n2767), .B2(n3747), .A(n2766), .ZN(n2768) );
  NAND2_X1 U35120 ( .A1(n4185), .A2(n2529), .ZN(n2774) );
  INV_X1 U35130 ( .A(REG2_REG_26__SCAN_IN), .ZN(n2771) );
  NAND2_X1 U35140 ( .A1(n2538), .A2(REG0_REG_26__SCAN_IN), .ZN(n2770) );
  NAND2_X1 U35150 ( .A1(n2537), .A2(REG1_REG_26__SCAN_IN), .ZN(n2769) );
  OAI211_X1 U35160 ( .C1(n2771), .C2(n2562), .A(n2770), .B(n2769), .ZN(n2772)
         );
  INV_X1 U35170 ( .A(n2772), .ZN(n2773) );
  NAND2_X1 U35180 ( .A1(n4194), .A2(n4176), .ZN(n2775) );
  INV_X1 U35190 ( .A(REG3_REG_27__SCAN_IN), .ZN(n3694) );
  AND2_X1 U35200 ( .A1(n2776), .A2(n3694), .ZN(n2777) );
  INV_X1 U35210 ( .A(REG2_REG_27__SCAN_IN), .ZN(n2780) );
  NAND2_X1 U35220 ( .A1(n2537), .A2(REG1_REG_27__SCAN_IN), .ZN(n2779) );
  NAND2_X1 U35230 ( .A1(n2538), .A2(REG0_REG_27__SCAN_IN), .ZN(n2778) );
  OAI211_X1 U35240 ( .C1(n2780), .C2(n2562), .A(n2779), .B(n2778), .ZN(n2781)
         );
  INV_X1 U35250 ( .A(n2781), .ZN(n2782) );
  NAND2_X1 U35260 ( .A1(n4146), .A2(n4384), .ZN(n2784) );
  NOR2_X1 U35270 ( .A1(n4146), .A2(n4384), .ZN(n2783) );
  NAND2_X1 U35280 ( .A1(n2785), .A2(REG3_REG_28__SCAN_IN), .ZN(n4134) );
  INV_X1 U35290 ( .A(n2785), .ZN(n2786) );
  INV_X1 U35300 ( .A(REG3_REG_28__SCAN_IN), .ZN(n3685) );
  NAND2_X1 U35310 ( .A1(n2786), .A2(n3685), .ZN(n2787) );
  NAND2_X1 U35320 ( .A1(n4134), .A2(n2787), .ZN(n3684) );
  OR2_X1 U35330 ( .A1(n3684), .A2(n2843), .ZN(n2793) );
  INV_X1 U35340 ( .A(REG2_REG_28__SCAN_IN), .ZN(n2790) );
  NAND2_X1 U35350 ( .A1(n2537), .A2(REG1_REG_28__SCAN_IN), .ZN(n2789) );
  NAND2_X1 U35360 ( .A1(n2538), .A2(REG0_REG_28__SCAN_IN), .ZN(n2788) );
  OAI211_X1 U35370 ( .C1(n2790), .C2(n2562), .A(n2789), .B(n2788), .ZN(n2791)
         );
  INV_X1 U35380 ( .A(n2791), .ZN(n2792) );
  XNOR2_X1 U35390 ( .A(n2897), .B(n3895), .ZN(n4152) );
  NAND2_X1 U35400 ( .A1(n2252), .A2(IR_REG_31__SCAN_IN), .ZN(n2797) );
  INV_X1 U35410 ( .A(IR_REG_21__SCAN_IN), .ZN(n2798) );
  INV_X1 U35420 ( .A(n2860), .ZN(n2804) );
  NAND2_X1 U35430 ( .A1(n2800), .A2(n2794), .ZN(n2801) );
  NAND2_X1 U35440 ( .A1(n2801), .A2(IR_REG_31__SCAN_IN), .ZN(n2803) );
  XNOR2_X1 U35450 ( .A(n2923), .B(n3976), .ZN(n2806) );
  AND2_X1 U35460 ( .A1(n3963), .A2(n4519), .ZN(n3129) );
  INV_X1 U35470 ( .A(n4690), .ZN(n4696) );
  NAND2_X1 U35480 ( .A1(n3153), .A2(n3127), .ZN(n3898) );
  NAND2_X1 U35490 ( .A1(n2808), .A2(n3901), .ZN(n4354) );
  NAND2_X1 U35500 ( .A1(n4354), .A2(n4356), .ZN(n2810) );
  NAND2_X1 U35510 ( .A1(n2810), .A2(n3902), .ZN(n3134) );
  NAND2_X1 U35520 ( .A1(n2947), .A2(n3231), .ZN(n3907) );
  INV_X1 U35530 ( .A(n3231), .ZN(n2949) );
  NAND2_X1 U35540 ( .A1(n4363), .A2(n2949), .ZN(n3904) );
  AND2_X1 U35550 ( .A1(n3907), .A2(n3904), .ZN(n3857) );
  NAND2_X1 U35560 ( .A1(n3134), .A2(n3857), .ZN(n2811) );
  NAND2_X1 U35570 ( .A1(n2811), .A2(n3907), .ZN(n3181) );
  INV_X1 U35580 ( .A(n3908), .ZN(n2812) );
  AND2_X1 U35590 ( .A1(n3998), .A2(n3249), .ZN(n3245) );
  INV_X1 U35600 ( .A(n3998), .ZN(n3275) );
  NAND2_X1 U35610 ( .A1(n3275), .A2(n3303), .ZN(n3923) );
  INV_X1 U35620 ( .A(n3272), .ZN(n3319) );
  NAND2_X1 U35630 ( .A1(n3997), .A2(n3319), .ZN(n3921) );
  INV_X1 U35640 ( .A(n3997), .ZN(n3288) );
  NAND2_X1 U35650 ( .A1(n3288), .A2(n3272), .ZN(n3913) );
  NAND2_X1 U35660 ( .A1(n2813), .A2(n3913), .ZN(n3283) );
  INV_X1 U35670 ( .A(n2814), .ZN(n2815) );
  OR2_X1 U35680 ( .A1(n3283), .A2(n2815), .ZN(n2816) );
  NAND2_X1 U35690 ( .A1(n3353), .A2(n3332), .ZN(n3918) );
  NAND2_X1 U35700 ( .A1(n3994), .A2(n3369), .ZN(n3915) );
  AND2_X1 U35710 ( .A1(n3993), .A2(n3379), .ZN(n3930) );
  NAND2_X1 U35720 ( .A1(n3447), .A2(n3347), .ZN(n3917) );
  NAND2_X1 U35730 ( .A1(n2817), .A2(n3917), .ZN(n3445) );
  NAND2_X1 U35740 ( .A1(n3992), .A2(n3446), .ZN(n3933) );
  NAND2_X1 U35750 ( .A1(n3445), .A2(n3933), .ZN(n2818) );
  NAND2_X1 U35760 ( .A1(n3390), .A2(n2890), .ZN(n3931) );
  NAND2_X1 U35770 ( .A1(n2818), .A2(n3931), .ZN(n3402) );
  NAND2_X1 U35780 ( .A1(n3990), .A2(n3537), .ZN(n3479) );
  NAND2_X1 U35790 ( .A1(n3989), .A2(n3560), .ZN(n2819) );
  NAND2_X1 U35800 ( .A1(n3479), .A2(n2819), .ZN(n2822) );
  INV_X1 U35810 ( .A(n3401), .ZN(n2820) );
  NOR2_X1 U3582 ( .A1(n2822), .A2(n2820), .ZN(n3934) );
  NAND2_X1 U3583 ( .A1(n3402), .A2(n3934), .ZN(n2826) );
  NAND2_X1 U3584 ( .A1(n2821), .A2(n3525), .ZN(n3481) );
  NAND2_X1 U3585 ( .A1(n3399), .A2(n3481), .ZN(n2825) );
  INV_X1 U3586 ( .A(n2822), .ZN(n2824) );
  NOR2_X1 U3587 ( .A1(n3989), .A2(n3560), .ZN(n2823) );
  AOI21_X1 U3588 ( .B1(n2825), .B2(n2824), .A(n2823), .ZN(n3936) );
  NAND2_X1 U3589 ( .A1(n2826), .A2(n3936), .ZN(n3820) );
  INV_X1 U3590 ( .A(n3428), .ZN(n3886) );
  NAND2_X1 U3591 ( .A1(n3820), .A2(n3886), .ZN(n3430) );
  NAND2_X1 U3592 ( .A1(n3430), .A2(n3816), .ZN(n3459) );
  INV_X1 U3593 ( .A(n3987), .ZN(n4529) );
  NAND2_X1 U3594 ( .A1(n4529), .A2(n3584), .ZN(n3819) );
  INV_X1 U3595 ( .A(n3584), .ZN(n3808) );
  NAND2_X1 U3596 ( .A1(n3987), .A2(n3808), .ZN(n3818) );
  NAND2_X1 U3597 ( .A1(n3819), .A2(n3818), .ZN(n3883) );
  OR2_X1 U3598 ( .A1(n3459), .A2(n3883), .ZN(n2827) );
  NAND2_X1 U3599 ( .A1(n2827), .A2(n3818), .ZN(n3495) );
  INV_X1 U3600 ( .A(n3502), .ZN(n3887) );
  NAND2_X1 U3601 ( .A1(n3495), .A2(n3887), .ZN(n2828) );
  NAND2_X1 U3602 ( .A1(n2828), .A2(n3821), .ZN(n4231) );
  NAND2_X1 U3603 ( .A1(n4533), .A2(n3598), .ZN(n4312) );
  NAND2_X1 U3604 ( .A1(n4317), .A2(n4312), .ZN(n2831) );
  NAND2_X1 U3605 ( .A1(n4339), .A2(n4327), .ZN(n2829) );
  AND2_X1 U3606 ( .A1(n4315), .A2(n2829), .ZN(n4232) );
  NOR2_X1 U3607 ( .A1(n4339), .A2(n4327), .ZN(n2830) );
  AOI21_X1 U3608 ( .B1(n2831), .B2(n4232), .A(n2830), .ZN(n4286) );
  INV_X1 U3609 ( .A(n4290), .ZN(n4301) );
  OR2_X1 U3610 ( .A1(n4322), .A2(n4301), .ZN(n2832) );
  NAND2_X1 U3611 ( .A1(n4231), .A2(n4234), .ZN(n2833) );
  NAND2_X1 U3612 ( .A1(n4557), .A2(n4434), .ZN(n4229) );
  NAND2_X1 U3613 ( .A1(n4232), .A2(n4229), .ZN(n3944) );
  AND2_X1 U3614 ( .A1(n4322), .A2(n4301), .ZN(n4233) );
  AOI21_X1 U3615 ( .B1(n4234), .B2(n3944), .A(n4233), .ZN(n3823) );
  OR2_X1 U3616 ( .A1(n4258), .A2(n4415), .ZN(n4235) );
  NAND2_X1 U3617 ( .A1(n4236), .A2(n4235), .ZN(n3950) );
  INV_X1 U3618 ( .A(n3950), .ZN(n2834) );
  NAND2_X1 U3619 ( .A1(n3984), .A2(n4225), .ZN(n2836) );
  NAND2_X1 U3620 ( .A1(n2836), .A2(n2835), .ZN(n3953) );
  AND2_X1 U3621 ( .A1(n4258), .A2(n4415), .ZN(n3948) );
  AND2_X1 U3622 ( .A1(n4236), .A2(n3948), .ZN(n2837) );
  NOR2_X1 U3623 ( .A1(n3953), .A2(n2837), .ZN(n3827) );
  NAND2_X1 U3624 ( .A1(n4243), .A2(n4218), .ZN(n3881) );
  OR2_X1 U3625 ( .A1(n3984), .A2(n4225), .ZN(n4206) );
  AND2_X1 U3626 ( .A1(n3881), .A2(n4206), .ZN(n3952) );
  NAND2_X1 U3627 ( .A1(n3983), .A2(n4399), .ZN(n3880) );
  NAND2_X1 U3628 ( .A1(n2838), .A2(n3880), .ZN(n4191) );
  AND2_X1 U3629 ( .A1(n4178), .A2(n4197), .ZN(n3892) );
  OR2_X1 U3630 ( .A1(n4191), .A2(n3892), .ZN(n4173) );
  NAND2_X1 U3631 ( .A1(n4385), .A2(n4176), .ZN(n3853) );
  OR2_X1 U3632 ( .A1(n4178), .A2(n4197), .ZN(n4172) );
  AND2_X1 U3633 ( .A1(n3853), .A2(n4172), .ZN(n3961) );
  AND2_X1 U3634 ( .A1(n4194), .A2(n4183), .ZN(n3852) );
  AND2_X1 U3635 ( .A1(n4177), .A2(n4384), .ZN(n3959) );
  INV_X1 U3636 ( .A(n3959), .ZN(n2839) );
  OR2_X1 U3637 ( .A1(n4177), .A2(n4384), .ZN(n2840) );
  INV_X1 U3638 ( .A(n2840), .ZN(n3838) );
  INV_X1 U3639 ( .A(n3895), .ZN(n2841) );
  XNOR2_X1 U3640 ( .A(n2899), .B(n2841), .ZN(n2854) );
  NAND2_X1 U3641 ( .A1(n3976), .A2(n4519), .ZN(n2842) );
  INV_X1 U3642 ( .A(n3963), .ZN(n3850) );
  NAND2_X1 U3643 ( .A1(n4518), .A2(n3850), .ZN(n3845) );
  OR2_X1 U3644 ( .A1(n4134), .A2(n2843), .ZN(n2848) );
  INV_X1 U3645 ( .A(REG2_REG_29__SCAN_IN), .ZN(n4130) );
  NAND2_X1 U3646 ( .A1(n2538), .A2(REG0_REG_29__SCAN_IN), .ZN(n2845) );
  NAND2_X1 U3647 ( .A1(n2537), .A2(REG1_REG_29__SCAN_IN), .ZN(n2844) );
  OAI211_X1 U3648 ( .C1(n4130), .C2(n2562), .A(n2845), .B(n2844), .ZN(n2846)
         );
  INV_X1 U3649 ( .A(n2846), .ZN(n2847) );
  NAND2_X1 U3650 ( .A1(n2848), .A2(n2847), .ZN(n3981) );
  NAND2_X1 U3651 ( .A1(n2271), .A2(IR_REG_31__SCAN_IN), .ZN(n2849) );
  MUX2_X1 U3652 ( .A(n2849), .B(IR_REG_31__SCAN_IN), .S(n2508), .Z(n2852) );
  INV_X1 U3653 ( .A(n2850), .ZN(n2851) );
  AND2_X1 U3654 ( .A1(n3981), .A2(n4362), .ZN(n2853) );
  AOI21_X1 U3655 ( .B1(n2854), .B2(n4342), .A(n2853), .ZN(n4147) );
  AOI22_X1 U3656 ( .A1(n4177), .A2(n4291), .B1(n4380), .B2(n4143), .ZN(n2855)
         );
  OAI211_X1 U3657 ( .C1(n4152), .C2(n4441), .A(n4147), .B(n2855), .ZN(n2894)
         );
  NOR2_X1 U3658 ( .A1(n2856), .A2(n2863), .ZN(n2857) );
  MUX2_X1 U3659 ( .A(n2863), .B(n2857), .S(IR_REG_25__SCAN_IN), .Z(n2859) );
  NAND2_X1 U3660 ( .A1(n3015), .A2(B_REG_SCAN_IN), .ZN(n2862) );
  MUX2_X1 U3661 ( .A(n2862), .B(B_REG_SCAN_IN), .S(n2868), .Z(n2865) );
  NAND2_X1 U3662 ( .A1(n2866), .A2(n3015), .ZN(n3036) );
  NAND2_X1 U3663 ( .A1(n2984), .A2(n3036), .ZN(n2886) );
  NAND2_X1 U3664 ( .A1(n4690), .A2(n3866), .ZN(n3002) );
  NAND2_X1 U3665 ( .A1(n3963), .A2(n4116), .ZN(n2986) );
  NAND2_X1 U3666 ( .A1(n3042), .A2(n2986), .ZN(n3120) );
  NAND2_X1 U3667 ( .A1(n3002), .A2(n3120), .ZN(n2873) );
  NOR2_X1 U3668 ( .A1(n3118), .A2(n2873), .ZN(n2885) );
  NOR4_X1 U3669 ( .A1(D_REG_30__SCAN_IN), .A2(D_REG_13__SCAN_IN), .A3(
        D_REG_31__SCAN_IN), .A4(D_REG_12__SCAN_IN), .ZN(n2877) );
  NOR4_X1 U3670 ( .A1(D_REG_8__SCAN_IN), .A2(D_REG_4__SCAN_IN), .A3(
        D_REG_15__SCAN_IN), .A4(D_REG_26__SCAN_IN), .ZN(n2876) );
  NOR4_X1 U3671 ( .A1(D_REG_25__SCAN_IN), .A2(D_REG_19__SCAN_IN), .A3(
        D_REG_10__SCAN_IN), .A4(D_REG_6__SCAN_IN), .ZN(n2875) );
  NOR4_X1 U3672 ( .A1(D_REG_11__SCAN_IN), .A2(D_REG_20__SCAN_IN), .A3(
        D_REG_7__SCAN_IN), .A4(D_REG_18__SCAN_IN), .ZN(n2874) );
  NAND4_X1 U3673 ( .A1(n2877), .A2(n2876), .A3(n2875), .A4(n2874), .ZN(n2883)
         );
  NOR2_X1 U3674 ( .A1(D_REG_29__SCAN_IN), .A2(D_REG_27__SCAN_IN), .ZN(n2881)
         );
  NOR4_X1 U3675 ( .A1(D_REG_28__SCAN_IN), .A2(D_REG_5__SCAN_IN), .A3(
        D_REG_23__SCAN_IN), .A4(D_REG_22__SCAN_IN), .ZN(n2880) );
  NOR4_X1 U3676 ( .A1(D_REG_9__SCAN_IN), .A2(D_REG_14__SCAN_IN), .A3(
        D_REG_3__SCAN_IN), .A4(D_REG_24__SCAN_IN), .ZN(n2879) );
  NOR4_X1 U3677 ( .A1(D_REG_21__SCAN_IN), .A2(D_REG_17__SCAN_IN), .A3(
        D_REG_16__SCAN_IN), .A4(D_REG_2__SCAN_IN), .ZN(n2878) );
  NAND4_X1 U3678 ( .A1(n2881), .A2(n2880), .A3(n2879), .A4(n2878), .ZN(n2882)
         );
  NOR2_X1 U3679 ( .A1(n2883), .A2(n2882), .ZN(n2884) );
  INV_X1 U3680 ( .A(n2868), .ZN(n2887) );
  NAND2_X1 U3681 ( .A1(n2887), .A2(n2866), .ZN(n3038) );
  MUX2_X1 U3682 ( .A(REG1_REG_28__SCAN_IN), .B(n2894), .S(n4716), .Z(n2889) );
  INV_X1 U3683 ( .A(n2889), .ZN(n2892) );
  NAND2_X1 U3684 ( .A1(n3250), .A2(n3249), .ZN(n3263) );
  NAND2_X1 U3685 ( .A1(n3489), .A2(n3560), .ZN(n3488) );
  NAND2_X1 U3686 ( .A1(n4299), .A2(n4415), .ZN(n4278) );
  INV_X1 U3687 ( .A(n2914), .ZN(n2891) );
  OAI21_X1 U3688 ( .B1(n4160), .B2(n3686), .A(n2891), .ZN(n4141) );
  NAND2_X1 U3689 ( .A1(n2892), .A2(n2489), .ZN(U3546) );
  MUX2_X1 U3690 ( .A(REG0_REG_28__SCAN_IN), .B(n2894), .S(n4704), .Z(n2895) );
  INV_X1 U3691 ( .A(n2895), .ZN(n2896) );
  NAND2_X1 U3692 ( .A1(n2896), .A2(n2486), .ZN(U3514) );
  OAI21_X1 U3693 ( .B1(n2897), .B2(n3895), .A(n2490), .ZN(n2898) );
  XNOR2_X1 U3694 ( .A(n3981), .B(n4133), .ZN(n3896) );
  XNOR2_X1 U3695 ( .A(n2898), .B(n3896), .ZN(n4129) );
  NAND2_X1 U3696 ( .A1(n4129), .A2(n4694), .ZN(n2909) );
  INV_X1 U3697 ( .A(n3896), .ZN(n2900) );
  INV_X1 U3698 ( .A(REG2_REG_30__SCAN_IN), .ZN(n2903) );
  NAND2_X1 U3699 ( .A1(n2537), .A2(REG1_REG_30__SCAN_IN), .ZN(n2902) );
  NAND2_X1 U3700 ( .A1(n2538), .A2(REG0_REG_30__SCAN_IN), .ZN(n2901) );
  OAI211_X1 U3701 ( .C1(n2562), .C2(n2903), .A(n2902), .B(n2901), .ZN(n3980)
         );
  INV_X1 U3702 ( .A(n3980), .ZN(n2906) );
  INV_X1 U3703 ( .A(B_REG_SCAN_IN), .ZN(n2905) );
  XNOR2_X1 U3704 ( .A(n2904), .B(n2482), .ZN(n4001) );
  OAI21_X1 U3705 ( .B1(n2905), .B2(n4001), .A(n4362), .ZN(n4122) );
  OAI22_X1 U3706 ( .A1(n2907), .A2(n4366), .B1(n2906), .B2(n4122), .ZN(n4137)
         );
  OAI22_X1 U3707 ( .A1(n4131), .A2(n4435), .B1(n2913), .B2(n4433), .ZN(n2908)
         );
  NAND2_X1 U3708 ( .A1(n2912), .A2(n2911), .ZN(n2915) );
  NAND2_X1 U3709 ( .A1(n2914), .A2(n2913), .ZN(n4377) );
  OAI21_X1 U3710 ( .B1(n2914), .B2(n2913), .A(n4377), .ZN(n4135) );
  NAND2_X1 U3711 ( .A1(n2915), .A2(n2485), .ZN(U3515) );
  INV_X1 U3712 ( .A(REG1_REG_29__SCAN_IN), .ZN(n2917) );
  NAND2_X1 U3713 ( .A1(n4713), .A2(n2917), .ZN(n2918) );
  NAND2_X1 U3714 ( .A1(n2919), .A2(n2491), .ZN(U3547) );
  INV_X2 U3715 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  NAND2_X2 U3716 ( .A1(n2921), .A2(n3124), .ZN(n3618) );
  NAND2_X2 U3717 ( .A1(n2921), .A2(n2923), .ZN(n2934) );
  BUF_X4 U3718 ( .A(n2934), .Z(n3677) );
  OAI22_X1 U3719 ( .A1(n3390), .A2(n3678), .B1(n3677), .B2(n3446), .ZN(n2925)
         );
  NOR2_X1 U3720 ( .A1(n2922), .A2(n4519), .ZN(n2996) );
  INV_X1 U3721 ( .A(n2996), .ZN(n2924) );
  XNOR2_X1 U3722 ( .A(n2925), .B(n3675), .ZN(n3416) );
  INV_X2 U3723 ( .A(n2934), .ZN(n2926) );
  NAND2_X4 U3724 ( .A1(n2926), .A2(n4678), .ZN(n3674) );
  OAI22_X1 U3725 ( .A1(n3390), .A2(n3674), .B1(n3663), .B2(n3446), .ZN(n3415)
         );
  XNOR2_X1 U3726 ( .A(n3416), .B(n3415), .ZN(n2991) );
  XNOR2_X1 U3727 ( .A(n2927), .B(n3675), .ZN(n2939) );
  INV_X1 U3728 ( .A(n3674), .ZN(n2929) );
  NAND2_X1 U3729 ( .A1(n2929), .A2(n2933), .ZN(n2932) );
  INV_X1 U3730 ( .A(n3618), .ZN(n3585) );
  INV_X1 U3731 ( .A(n2921), .ZN(n2930) );
  AOI22_X1 U3732 ( .A1(n3585), .A2(n3127), .B1(n2930), .B2(IR_REG_0__SCAN_IN), 
        .ZN(n2931) );
  NAND2_X1 U3733 ( .A1(n2932), .A2(n2931), .ZN(n3080) );
  NAND2_X1 U3734 ( .A1(n2933), .A2(n3636), .ZN(n2936) );
  NAND2_X1 U3735 ( .A1(n2926), .A2(n3127), .ZN(n2937) );
  INV_X1 U3736 ( .A(REG1_REG_0__SCAN_IN), .ZN(n2935) );
  NAND2_X1 U3737 ( .A1(n3080), .A2(n3079), .ZN(n3078) );
  NAND2_X1 U3738 ( .A1(n2937), .A2(n3661), .ZN(n2938) );
  AND2_X1 U3739 ( .A1(n3078), .A2(n2938), .ZN(n3151) );
  NOR2_X1 U3740 ( .A1(n3150), .A2(n2941), .ZN(n3142) );
  XNOR2_X1 U3741 ( .A(n2942), .B(n3675), .ZN(n2945) );
  XNOR2_X1 U3742 ( .A(n2945), .B(n2943), .ZN(n3143) );
  NAND2_X1 U3743 ( .A1(n3142), .A2(n3143), .ZN(n3141) );
  OR2_X1 U3744 ( .A1(n2945), .A2(n2944), .ZN(n2946) );
  NAND2_X1 U3745 ( .A1(n3141), .A2(n2946), .ZN(n3172) );
  XNOR2_X1 U3746 ( .A(n2948), .B(n3675), .ZN(n2951) );
  NOR2_X1 U3747 ( .A1(n3663), .A2(n2949), .ZN(n2950) );
  AOI21_X1 U3748 ( .B1(n3665), .B2(n4363), .A(n2950), .ZN(n2952) );
  XNOR2_X1 U3749 ( .A(n2951), .B(n2952), .ZN(n3171) );
  INV_X1 U3750 ( .A(n2951), .ZN(n2953) );
  AOI21_X1 U3751 ( .B1(n3172), .B2(n3171), .A(n2483), .ZN(n3214) );
  OAI22_X1 U3752 ( .A1(n3305), .A2(n3674), .B1(n3663), .B2(n3215), .ZN(n2956)
         );
  OAI22_X1 U3753 ( .A1(n3305), .A2(n3663), .B1(n3677), .B2(n3215), .ZN(n2954)
         );
  XNOR2_X1 U3754 ( .A(n2954), .B(n2232), .ZN(n2955) );
  XOR2_X1 U3755 ( .A(n2956), .B(n2955), .Z(n3213) );
  NAND2_X1 U3756 ( .A1(n3214), .A2(n3213), .ZN(n3212) );
  NAND2_X1 U3757 ( .A1(n3212), .A2(n2957), .ZN(n3237) );
  OAI22_X1 U3758 ( .A1(n3275), .A2(n3674), .B1(n3663), .B2(n3249), .ZN(n2962)
         );
  NAND2_X1 U3759 ( .A1(n3998), .A2(n3636), .ZN(n2959) );
  NAND2_X1 U3760 ( .A1(n2926), .A2(n3303), .ZN(n2958) );
  NAND2_X1 U3761 ( .A1(n2959), .A2(n2958), .ZN(n2960) );
  XNOR2_X1 U3762 ( .A(n2960), .B(n2232), .ZN(n2961) );
  XOR2_X1 U3763 ( .A(n2962), .B(n2961), .Z(n3236) );
  OAI22_X1 U3764 ( .A1(n3288), .A2(n3674), .B1(n3663), .B2(n3319), .ZN(n2965)
         );
  INV_X1 U3765 ( .A(n2965), .ZN(n3313) );
  OAI22_X1 U3766 ( .A1(n3288), .A2(n3678), .B1(n3677), .B2(n3319), .ZN(n2964)
         );
  XNOR2_X1 U3767 ( .A(n2964), .B(n3675), .ZN(n3314) );
  OAI22_X1 U3768 ( .A1(n3368), .A2(n3674), .B1(n3663), .B2(n3570), .ZN(n2967)
         );
  OAI22_X1 U3769 ( .A1(n3368), .A2(n3678), .B1(n3677), .B2(n3570), .ZN(n2966)
         );
  XNOR2_X1 U3770 ( .A(n2966), .B(n2232), .ZN(n2968) );
  XOR2_X1 U3771 ( .A(n2967), .B(n2968), .Z(n3565) );
  NAND2_X1 U3772 ( .A1(n3994), .A2(n3585), .ZN(n2970) );
  NAND2_X1 U3773 ( .A1(n2926), .A2(n3332), .ZN(n2969) );
  NAND2_X1 U3774 ( .A1(n2970), .A2(n2969), .ZN(n2971) );
  XNOR2_X1 U3775 ( .A(n2971), .B(n3661), .ZN(n2976) );
  INV_X1 U3776 ( .A(n2976), .ZN(n2974) );
  NOR2_X1 U3777 ( .A1(n3663), .A2(n3369), .ZN(n2972) );
  AOI21_X1 U3778 ( .B1(n3665), .B2(n3994), .A(n2972), .ZN(n2975) );
  INV_X1 U3779 ( .A(n2975), .ZN(n2973) );
  AND2_X1 U3780 ( .A1(n2976), .A2(n2975), .ZN(n3365) );
  NOR2_X1 U3781 ( .A1(n3663), .A2(n3379), .ZN(n2977) );
  AOI21_X1 U3782 ( .B1(n3665), .B2(n3993), .A(n2977), .ZN(n2979) );
  OAI22_X1 U3783 ( .A1(n3447), .A2(n3678), .B1(n3677), .B2(n3379), .ZN(n2978)
         );
  XNOR2_X1 U3784 ( .A(n2978), .B(n2232), .ZN(n2981) );
  XOR2_X1 U3785 ( .A(n2979), .B(n2981), .Z(n3376) );
  INV_X1 U3786 ( .A(n2979), .ZN(n2980) );
  OR2_X1 U3787 ( .A1(n2981), .A2(n2980), .ZN(n2982) );
  INV_X1 U3788 ( .A(n3042), .ZN(n2988) );
  NAND2_X1 U3789 ( .A1(n3126), .A2(n2986), .ZN(n2987) );
  NAND2_X1 U3790 ( .A1(n2988), .A2(n2987), .ZN(n2992) );
  OR2_X1 U3791 ( .A1(n3118), .A2(n2992), .ZN(n2989) );
  AOI211_X1 U3792 ( .C1(n2991), .C2(n2990), .A(n3813), .B(n2270), .ZN(n3009)
         );
  NAND2_X1 U3793 ( .A1(n2992), .A2(n4433), .ZN(n2993) );
  NAND2_X1 U3794 ( .A1(n3005), .A2(n2993), .ZN(n2994) );
  NAND2_X1 U3795 ( .A1(n2994), .A2(n3120), .ZN(n3112) );
  NAND2_X1 U3796 ( .A1(n2921), .A2(n3041), .ZN(n2995) );
  OAI21_X1 U3797 ( .B1(n3112), .B2(n2995), .A(STATE_REG_SCAN_IN), .ZN(n2998)
         );
  NAND2_X1 U3798 ( .A1(n4666), .A2(n2996), .ZN(n2997) );
  NAND2_X1 U3799 ( .A1(n3005), .A2(n3974), .ZN(n3111) );
  NOR2_X1 U3800 ( .A1(n4563), .A2(n2999), .ZN(n3008) );
  NAND2_X1 U3801 ( .A1(n3974), .A2(n3083), .ZN(n3000) );
  NAND2_X1 U3802 ( .A1(REG3_REG_10__SCAN_IN), .A2(U3149), .ZN(n4582) );
  OAI21_X1 U3803 ( .B1(n4528), .B2(n3447), .A(n4582), .ZN(n3007) );
  OR2_X1 U3804 ( .A1(n3118), .A2(n4433), .ZN(n3001) );
  OR2_X1 U3805 ( .A1(n3005), .A2(n3001), .ZN(n3003) );
  NAND2_X1 U3806 ( .A1(n3974), .A2(n3046), .ZN(n3004) );
  OAI22_X1 U3807 ( .A1(n4531), .A2(n3446), .B1(n3538), .B2(n4546), .ZN(n3006)
         );
  OR4_X1 U3808 ( .A1(n3009), .A2(n3008), .A3(n3007), .A4(n3006), .ZN(U3214) );
  INV_X1 U3809 ( .A(n4022), .ZN(n4031) );
  INV_X1 U3810 ( .A(DATAI_2_), .ZN(n3010) );
  MUX2_X1 U3811 ( .A(n4031), .B(n3010), .S(U3149), .Z(n3011) );
  INV_X1 U3812 ( .A(n3011), .ZN(U3350) );
  INV_X1 U3813 ( .A(DATAI_8_), .ZN(n3012) );
  INV_X1 U3814 ( .A(n3161), .ZN(n4046) );
  MUX2_X1 U3815 ( .A(n3012), .B(n4046), .S(STATE_REG_SCAN_IN), .Z(n3013) );
  INV_X1 U3816 ( .A(n3013), .ZN(U3344) );
  NAND2_X1 U3817 ( .A1(U3149), .A2(DATAI_25_), .ZN(n3014) );
  OAI21_X1 U3818 ( .B1(n3015), .B2(U3149), .A(n3014), .ZN(U3327) );
  INV_X1 U3819 ( .A(DATAI_26_), .ZN(n4967) );
  NAND2_X1 U3820 ( .A1(n3016), .A2(STATE_REG_SCAN_IN), .ZN(n3017) );
  OAI21_X1 U3821 ( .B1(STATE_REG_SCAN_IN), .B2(n4967), .A(n3017), .ZN(U3326)
         );
  INV_X1 U3822 ( .A(DATAI_27_), .ZN(n4968) );
  INV_X1 U3823 ( .A(n4001), .ZN(n3018) );
  NAND2_X1 U3824 ( .A1(n3018), .A2(STATE_REG_SCAN_IN), .ZN(n3019) );
  OAI21_X1 U3825 ( .B1(STATE_REG_SCAN_IN), .B2(n4968), .A(n3019), .ZN(U3325)
         );
  INV_X1 U3826 ( .A(DATAI_20_), .ZN(n4970) );
  NAND2_X1 U3827 ( .A1(n3850), .A2(STATE_REG_SCAN_IN), .ZN(n3020) );
  OAI21_X1 U3828 ( .B1(STATE_REG_SCAN_IN), .B2(n4970), .A(n3020), .ZN(U3332)
         );
  INV_X1 U3829 ( .A(DATAI_31_), .ZN(n5068) );
  INV_X1 U3830 ( .A(IR_REG_30__SCAN_IN), .ZN(n3021) );
  NAND4_X1 U3831 ( .A1(n3022), .A2(IR_REG_31__SCAN_IN), .A3(STATE_REG_SCAN_IN), 
        .A4(n3021), .ZN(n3023) );
  OAI21_X1 U3832 ( .B1(STATE_REG_SCAN_IN), .B2(n5068), .A(n3023), .ZN(U3321)
         );
  INV_X1 U3833 ( .A(DATAI_12_), .ZN(n3024) );
  MUX2_X1 U3834 ( .A(n3024), .B(n4043), .S(STATE_REG_SCAN_IN), .Z(n3025) );
  INV_X1 U3835 ( .A(n3025), .ZN(U3340) );
  INV_X1 U3836 ( .A(DATAI_22_), .ZN(n4791) );
  NAND2_X1 U3837 ( .A1(n3976), .A2(STATE_REG_SCAN_IN), .ZN(n3026) );
  OAI21_X1 U3838 ( .B1(STATE_REG_SCAN_IN), .B2(n4791), .A(n3026), .ZN(U3330)
         );
  INV_X1 U3839 ( .A(DATAI_28_), .ZN(n3028) );
  NAND2_X1 U3840 ( .A1(n3083), .A2(STATE_REG_SCAN_IN), .ZN(n3027) );
  OAI21_X1 U3841 ( .B1(STATE_REG_SCAN_IN), .B2(n3028), .A(n3027), .ZN(U3324)
         );
  INV_X1 U3842 ( .A(DATAI_24_), .ZN(n3030) );
  NAND2_X1 U3843 ( .A1(n2868), .A2(STATE_REG_SCAN_IN), .ZN(n3029) );
  OAI21_X1 U3844 ( .B1(STATE_REG_SCAN_IN), .B2(n3030), .A(n3029), .ZN(U3328)
         );
  INV_X1 U3845 ( .A(DATAI_30_), .ZN(n3033) );
  NAND2_X1 U3846 ( .A1(n3031), .A2(STATE_REG_SCAN_IN), .ZN(n3032) );
  OAI21_X1 U3847 ( .B1(STATE_REG_SCAN_IN), .B2(n3033), .A(n3032), .ZN(U3322)
         );
  INV_X1 U3848 ( .A(D_REG_1__SCAN_IN), .ZN(n5058) );
  INV_X1 U3849 ( .A(n3036), .ZN(n3037) );
  AOI22_X1 U3850 ( .A1(n4664), .A2(n5058), .B1(n3037), .B2(n4666), .ZN(U3459)
         );
  INV_X1 U3851 ( .A(D_REG_0__SCAN_IN), .ZN(n3040) );
  INV_X1 U3852 ( .A(n3038), .ZN(n3039) );
  AOI22_X1 U3853 ( .A1(n4664), .A2(n3040), .B1(n3039), .B2(n4666), .ZN(U3458)
         );
  OR2_X1 U3854 ( .A1(n3041), .A2(U3149), .ZN(n3978) );
  NAND2_X1 U3855 ( .A1(n3118), .A2(n3978), .ZN(n3045) );
  AOI21_X1 U3856 ( .B1(n3042), .B2(n3041), .A(n2741), .ZN(n3044) );
  INV_X1 U3857 ( .A(n3044), .ZN(n3043) );
  NOR2_X1 U3858 ( .A1(n4636), .A2(U4043), .ZN(U3148) );
  NOR2_X1 U3859 ( .A1(n3046), .A2(n4001), .ZN(n3973) );
  INV_X1 U3860 ( .A(REG2_REG_2__SCAN_IN), .ZN(n4023) );
  MUX2_X1 U3861 ( .A(REG2_REG_2__SCAN_IN), .B(n4023), .S(n4022), .Z(n3049) );
  INV_X1 U3862 ( .A(REG2_REG_1__SCAN_IN), .ZN(n3047) );
  AND2_X1 U3863 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n4011)
         );
  NAND2_X1 U3864 ( .A1(n4010), .A2(n4011), .ZN(n4025) );
  NAND2_X1 U3865 ( .A1(n4025), .A2(n4024), .ZN(n3048) );
  NAND2_X1 U3866 ( .A1(n3049), .A2(n3048), .ZN(n4028) );
  OAI21_X1 U3867 ( .B1(n4023), .B2(n4031), .A(n4028), .ZN(n3057) );
  XOR2_X1 U3868 ( .A(n4527), .B(n3057), .Z(n3058) );
  INV_X1 U3869 ( .A(REG2_REG_3__SCAN_IN), .ZN(n3227) );
  XNOR2_X1 U3870 ( .A(n3058), .B(n3227), .ZN(n3054) );
  INV_X1 U3871 ( .A(REG1_REG_2__SCAN_IN), .ZN(n4707) );
  MUX2_X1 U3872 ( .A(REG1_REG_2__SCAN_IN), .B(n4707), .S(n4022), .Z(n4021) );
  INV_X1 U3873 ( .A(REG1_REG_1__SCAN_IN), .ZN(n3050) );
  NAND2_X1 U3874 ( .A1(n4014), .A2(n4013), .ZN(n4012) );
  NAND2_X1 U3875 ( .A1(n4012), .A2(n3051), .ZN(n4020) );
  INV_X1 U3876 ( .A(n4637), .ZN(n3169) );
  AOI211_X1 U3877 ( .C1(n3207), .C2(n3052), .A(n3063), .B(n3169), .ZN(n3053)
         );
  AOI21_X1 U3878 ( .B1(n4593), .B2(n3054), .A(n3053), .ZN(n3056) );
  AOI22_X1 U3879 ( .A1(n4636), .A2(ADDR_REG_3__SCAN_IN), .B1(
        REG3_REG_3__SCAN_IN), .B2(U3149), .ZN(n3055) );
  OAI211_X1 U3880 ( .C1(n2441), .C2(n4642), .A(n3056), .B(n3055), .ZN(U3243)
         );
  AOI22_X1 U3881 ( .A1(n3058), .A2(REG2_REG_3__SCAN_IN), .B1(n4527), .B2(n3057), .ZN(n3059) );
  INV_X1 U3882 ( .A(REG2_REG_5__SCAN_IN), .ZN(n3301) );
  MUX2_X1 U3883 ( .A(n3301), .B(REG2_REG_5__SCAN_IN), .S(n4525), .Z(n3091) );
  XNOR2_X1 U3884 ( .A(n3101), .B(n4524), .ZN(n3103) );
  XNOR2_X1 U3885 ( .A(n3103), .B(REG2_REG_6__SCAN_IN), .ZN(n3069) );
  INV_X1 U3886 ( .A(n4642), .ZN(n4045) );
  NOR2_X1 U3887 ( .A1(STATE_REG_SCAN_IN), .A2(n3060), .ZN(n3316) );
  AOI21_X1 U3888 ( .B1(n4636), .B2(ADDR_REG_6__SCAN_IN), .A(n3316), .ZN(n3061)
         );
  INV_X1 U3889 ( .A(n3061), .ZN(n3067) );
  INV_X1 U3890 ( .A(REG1_REG_4__SCAN_IN), .ZN(n4709) );
  XNOR2_X1 U3891 ( .A(n4525), .B(REG1_REG_5__SCAN_IN), .ZN(n3088) );
  INV_X1 U3892 ( .A(REG1_REG_6__SCAN_IN), .ZN(n3267) );
  NOR2_X1 U3893 ( .A1(n3065), .A2(n3267), .ZN(n3099) );
  AOI211_X1 U3894 ( .C1(n3065), .C2(n3267), .A(n3169), .B(n3099), .ZN(n3066)
         );
  AOI211_X1 U3895 ( .C1(n4045), .C2(n4524), .A(n3067), .B(n3066), .ZN(n3068)
         );
  OAI21_X1 U3896 ( .B1(n3069), .B2(n4630), .A(n3068), .ZN(U3246) );
  XOR2_X1 U3897 ( .A(REG2_REG_4__SCAN_IN), .B(n3070), .Z(n3077) );
  NAND2_X1 U3898 ( .A1(U3149), .A2(REG3_REG_4__SCAN_IN), .ZN(n3216) );
  INV_X1 U3899 ( .A(n3216), .ZN(n3071) );
  AOI21_X1 U3900 ( .B1(n4636), .B2(ADDR_REG_4__SCAN_IN), .A(n3071), .ZN(n3072)
         );
  OAI21_X1 U3901 ( .B1(n4642), .B2(n2371), .A(n3072), .ZN(n3076) );
  AOI211_X1 U3902 ( .C1(n4709), .C2(n3074), .A(n3073), .B(n3169), .ZN(n3075)
         );
  AOI211_X1 U3903 ( .C1(n4593), .C2(n3077), .A(n3076), .B(n3075), .ZN(n3086)
         );
  NOR2_X1 U3904 ( .A1(n3080), .A2(n3079), .ZN(n3081) );
  OR2_X1 U3905 ( .A1(n3082), .A2(n3081), .ZN(n3114) );
  NAND3_X1 U3906 ( .A1(n3114), .A2(n3083), .A3(n4001), .ZN(n3085) );
  INV_X1 U3907 ( .A(IR_REG_0__SCAN_IN), .ZN(n4002) );
  OAI21_X1 U3908 ( .B1(REG2_REG_0__SCAN_IN), .B2(n4001), .A(n3083), .ZN(n4004)
         );
  AOI22_X1 U3909 ( .A1(n4002), .A2(n4004), .B1(n3973), .B2(n4011), .ZN(n3084)
         );
  NAND3_X1 U3910 ( .A1(n3085), .A2(U4043), .A3(n3084), .ZN(n4035) );
  NAND2_X1 U3911 ( .A1(n3086), .A2(n4035), .ZN(U3244) );
  AOI211_X1 U3912 ( .C1(n3089), .C2(n3088), .A(n3169), .B(n3087), .ZN(n3097)
         );
  AOI211_X1 U3913 ( .C1(n3092), .C2(n3091), .A(n3090), .B(n4630), .ZN(n3096)
         );
  INV_X1 U3914 ( .A(n4525), .ZN(n3094) );
  INV_X1 U3915 ( .A(REG3_REG_5__SCAN_IN), .ZN(n4998) );
  NOR2_X1 U3916 ( .A1(STATE_REG_SCAN_IN), .A2(n4998), .ZN(n3238) );
  AOI21_X1 U3917 ( .B1(n4636), .B2(ADDR_REG_5__SCAN_IN), .A(n3238), .ZN(n3093)
         );
  OAI21_X1 U3918 ( .B1(n4642), .B2(n3094), .A(n3093), .ZN(n3095) );
  OR3_X1 U3919 ( .A1(n3097), .A2(n3096), .A3(n3095), .ZN(U3245) );
  INV_X1 U3920 ( .A(REG1_REG_7__SCAN_IN), .ZN(n4711) );
  MUX2_X1 U3921 ( .A(REG1_REG_7__SCAN_IN), .B(n4711), .S(n4523), .Z(n3100) );
  XNOR2_X1 U3922 ( .A(n3159), .B(n3100), .ZN(n3109) );
  INV_X1 U3923 ( .A(n3101), .ZN(n3102) );
  AOI22_X1 U3924 ( .A1(n3103), .A2(REG2_REG_6__SCAN_IN), .B1(n4524), .B2(n3102), .ZN(n3105) );
  INV_X1 U3925 ( .A(REG2_REG_7__SCAN_IN), .ZN(n3293) );
  MUX2_X1 U3926 ( .A(n3293), .B(REG2_REG_7__SCAN_IN), .S(n4523), .Z(n3104) );
  AOI211_X1 U3927 ( .C1(n3105), .C2(n3104), .A(n4630), .B(n3163), .ZN(n3108)
         );
  INV_X1 U3928 ( .A(n4523), .ZN(n3160) );
  AND2_X1 U3929 ( .A1(U3149), .A2(REG3_REG_7__SCAN_IN), .ZN(n3567) );
  AOI21_X1 U3930 ( .B1(n4636), .B2(ADDR_REG_7__SCAN_IN), .A(n3567), .ZN(n3106)
         );
  OAI21_X1 U3931 ( .B1(n4642), .B2(n3160), .A(n3106), .ZN(n3107) );
  AOI211_X1 U3932 ( .C1(n3109), .C2(n4637), .A(n3108), .B(n3107), .ZN(n3110)
         );
  INV_X1 U3933 ( .A(n3110), .ZN(U3247) );
  INV_X1 U3934 ( .A(n3111), .ZN(n3113) );
  NOR3_X1 U3935 ( .A1(n3113), .A2(n3112), .A3(n3118), .ZN(n3158) );
  INV_X1 U3936 ( .A(REG3_REG_0__SCAN_IN), .ZN(n3117) );
  AOI21_X1 U3937 ( .B1(n3127), .B2(n4559), .A(n3115), .ZN(n3116) );
  OAI21_X1 U3938 ( .B1(n3158), .B2(n3117), .A(n3116), .ZN(U3229) );
  NAND2_X1 U3939 ( .A1(n2933), .A2(n3192), .ZN(n3900) );
  AND2_X1 U3940 ( .A1(n3898), .A2(n3900), .ZN(n4675) );
  OAI21_X1 U3941 ( .B1(n5058), .B2(n3118), .A(n4664), .ZN(n3119) );
  NAND4_X1 U3942 ( .A1(n3122), .A2(n3121), .A3(n3120), .A4(n3119), .ZN(n3123)
         );
  NAND2_X1 U3943 ( .A1(n3124), .A2(n4519), .ZN(n3222) );
  INV_X1 U3944 ( .A(n3222), .ZN(n3125) );
  NAND2_X1 U3945 ( .A1(n4654), .A2(n3125), .ZN(n4309) );
  NAND2_X1 U3946 ( .A1(n3127), .A2(n3126), .ZN(n4673) );
  AOI21_X1 U3947 ( .B1(n4366), .B2(n4298), .A(n4675), .ZN(n3128) );
  AOI21_X1 U3948 ( .B1(n4362), .B2(n2543), .A(n3128), .ZN(n4674) );
  OAI21_X1 U3949 ( .B1(n3129), .B2(n4673), .A(n4674), .ZN(n3130) );
  AOI22_X1 U3950 ( .A1(n3130), .A2(n4654), .B1(REG3_REG_0__SCAN_IN), .B2(n4643), .ZN(n3132) );
  NAND2_X1 U3951 ( .A1(n4663), .A2(REG2_REG_0__SCAN_IN), .ZN(n3131) );
  OAI211_X1 U3952 ( .C1(n4675), .C2(n4309), .A(n3132), .B(n3131), .ZN(U3290)
         );
  XNOR2_X1 U3953 ( .A(n3133), .B(n3857), .ZN(n3224) );
  XNOR2_X1 U3954 ( .A(n3134), .B(n3857), .ZN(n3135) );
  AOI22_X1 U3955 ( .A1(n3135), .A2(n4342), .B1(n4362), .B2(n3999), .ZN(n3225)
         );
  AOI22_X1 U3956 ( .A1(n4000), .A2(n4291), .B1(n4380), .B2(n3231), .ZN(n3136)
         );
  OAI211_X1 U3957 ( .C1(n4441), .C2(n3224), .A(n3225), .B(n3136), .ZN(n3209)
         );
  AND2_X1 U3958 ( .A1(n4683), .A2(n3231), .ZN(n3137) );
  OR2_X1 U3959 ( .A1(n3137), .A2(n3178), .ZN(n3234) );
  INV_X1 U3960 ( .A(REG0_REG_3__SCAN_IN), .ZN(n3138) );
  OAI22_X1 U3961 ( .A1(n4515), .A2(n3234), .B1(n4704), .B2(n3138), .ZN(n3139)
         );
  AOI21_X1 U3962 ( .B1(n3209), .B2(n4704), .A(n3139), .ZN(n3140) );
  INV_X1 U3963 ( .A(n3140), .ZN(U3473) );
  INV_X1 U3964 ( .A(REG3_REG_2__SCAN_IN), .ZN(n3148) );
  OAI21_X1 U3965 ( .B1(n3143), .B2(n3142), .A(n3141), .ZN(n3144) );
  NAND2_X1 U3966 ( .A1(n3144), .A2(n4554), .ZN(n3147) );
  AOI21_X1 U3967 ( .B1(n4369), .B2(n4559), .A(n3145), .ZN(n3146) );
  OAI211_X1 U3968 ( .C1(n3158), .C2(n3148), .A(n3147), .B(n3146), .ZN(U3234)
         );
  INV_X1 U3969 ( .A(REG3_REG_1__SCAN_IN), .ZN(n3157) );
  AOI211_X1 U3970 ( .C1(n3151), .C2(n3149), .A(n3813), .B(n3150), .ZN(n3152)
         );
  INV_X1 U3971 ( .A(n3152), .ZN(n3156) );
  OAI22_X1 U3972 ( .A1(n3153), .A2(n4528), .B1(n4546), .B2(n3228), .ZN(n3154)
         );
  AOI21_X1 U3973 ( .B1(n3197), .B2(n4559), .A(n3154), .ZN(n3155) );
  OAI211_X1 U3974 ( .C1(n3158), .C2(n3157), .A(n3156), .B(n3155), .ZN(U3219)
         );
  XNOR2_X1 U3975 ( .A(n3162), .B(n3161), .ZN(n4037) );
  XOR2_X1 U3976 ( .A(REG1_REG_8__SCAN_IN), .B(n4037), .Z(n3170) );
  XNOR2_X1 U3977 ( .A(REG2_REG_8__SCAN_IN), .B(n4047), .ZN(n3164) );
  NAND2_X1 U3978 ( .A1(n4593), .A2(n3164), .ZN(n3165) );
  NAND2_X1 U3979 ( .A1(REG3_REG_8__SCAN_IN), .A2(U3149), .ZN(n3370) );
  NAND2_X1 U3980 ( .A1(n3165), .A2(n3370), .ZN(n3167) );
  NOR2_X1 U3981 ( .A1(n4642), .A2(n4046), .ZN(n3166) );
  AOI211_X1 U3982 ( .C1(n4636), .C2(ADDR_REG_8__SCAN_IN), .A(n3167), .B(n3166), 
        .ZN(n3168) );
  OAI21_X1 U3983 ( .B1(n3170), .B2(n3169), .A(n3168), .ZN(U3248) );
  XOR2_X1 U3984 ( .A(n3172), .B(n3171), .Z(n3176) );
  OAI22_X1 U3985 ( .A1(n3228), .A2(n4528), .B1(n4546), .B2(n3305), .ZN(n3174)
         );
  MUX2_X1 U3986 ( .A(U3149), .B(n3811), .S(n4828), .Z(n3173) );
  AOI211_X1 U3987 ( .C1(n3231), .C2(n4559), .A(n3174), .B(n3173), .ZN(n3175)
         );
  OAI21_X1 U3988 ( .B1(n3176), .B2(n3813), .A(n3175), .ZN(U3215) );
  INV_X1 U3989 ( .A(n3250), .ZN(n3177) );
  OAI211_X1 U3990 ( .C1(n3178), .C2(n3215), .A(n3177), .B(n4701), .ZN(n4687)
         );
  NOR2_X1 U3991 ( .A1(n4687), .A2(n4519), .ZN(n3187) );
  XNOR2_X1 U3992 ( .A(n3179), .B(n3180), .ZN(n3188) );
  INV_X1 U3993 ( .A(n3180), .ZN(n3858) );
  XNOR2_X1 U3994 ( .A(n3181), .B(n3858), .ZN(n3185) );
  AOI22_X1 U3995 ( .A1(n3998), .A2(n4362), .B1(n3182), .B2(n4380), .ZN(n3183)
         );
  OAI21_X1 U3996 ( .B1(n2947), .B2(n4435), .A(n3183), .ZN(n3184) );
  AOI21_X1 U3997 ( .B1(n3185), .B2(n4342), .A(n3184), .ZN(n3186) );
  OAI21_X1 U3998 ( .B1(n3188), .B2(n4298), .A(n3186), .ZN(n4688) );
  AOI211_X1 U3999 ( .C1(n4643), .C2(n3211), .A(n3187), .B(n4688), .ZN(n3190)
         );
  INV_X1 U4000 ( .A(n3188), .ZN(n4691) );
  INV_X1 U4001 ( .A(n4309), .ZN(n4658) );
  AOI22_X1 U4002 ( .A1(n4691), .A2(n4658), .B1(REG2_REG_4__SCAN_IN), .B2(n4663), .ZN(n3189) );
  OAI21_X1 U4003 ( .B1(n3190), .B2(n4663), .A(n3189), .ZN(U3286) );
  INV_X2 U4004 ( .A(n4663), .ZN(n4654) );
  NAND2_X1 U4005 ( .A1(n4654), .A2(n4116), .ZN(n4347) );
  OAI21_X1 U4006 ( .B1(n3192), .B2(n3191), .A(n4370), .ZN(n4677) );
  AND2_X1 U4007 ( .A1(n3195), .A2(n3194), .ZN(n3196) );
  AOI22_X1 U4008 ( .A1(n4658), .A2(n3196), .B1(REG3_REG_1__SCAN_IN), .B2(n4643), .ZN(n3206) );
  INV_X1 U4009 ( .A(n3196), .ZN(n4679) );
  NAND2_X1 U4010 ( .A1(n4380), .A2(n3197), .ZN(n3199) );
  NAND2_X1 U4011 ( .A1(n2933), .A2(n4291), .ZN(n3198) );
  OAI211_X1 U4012 ( .C1(n3228), .C2(n4293), .A(n3199), .B(n3198), .ZN(n3200)
         );
  INV_X1 U4013 ( .A(n3200), .ZN(n3203) );
  NAND2_X1 U4014 ( .A1(n3201), .A2(n4342), .ZN(n3202) );
  OAI211_X1 U4015 ( .C1(n4679), .C2(n4298), .A(n3203), .B(n3202), .ZN(n4680)
         );
  MUX2_X1 U4016 ( .A(REG2_REG_1__SCAN_IN), .B(n4680), .S(n4654), .Z(n3204) );
  INV_X1 U4017 ( .A(n3204), .ZN(n3205) );
  OAI211_X1 U4018 ( .C1(n4328), .C2(n4677), .A(n3206), .B(n3205), .ZN(U3289)
         );
  INV_X1 U4019 ( .A(REG1_REG_3__SCAN_IN), .ZN(n3207) );
  OAI22_X1 U4020 ( .A1(n4458), .A2(n3234), .B1(n4716), .B2(n3207), .ZN(n3208)
         );
  AOI21_X1 U4021 ( .B1(n3209), .B2(n4716), .A(n3208), .ZN(n3210) );
  INV_X1 U4022 ( .A(n3210), .ZN(U3521) );
  INV_X1 U4023 ( .A(n3211), .ZN(n3221) );
  OAI211_X1 U4024 ( .C1(n3214), .C2(n3213), .A(n3212), .B(n4554), .ZN(n3220)
         );
  OAI22_X1 U4025 ( .A1(n4531), .A2(n3215), .B1(n2947), .B2(n4528), .ZN(n3218)
         );
  OAI21_X1 U4026 ( .B1(n4546), .B2(n3275), .A(n3216), .ZN(n3217) );
  NOR2_X1 U4027 ( .A1(n3218), .A2(n3217), .ZN(n3219) );
  OAI211_X1 U4028 ( .C1(n4563), .C2(n3221), .A(n3220), .B(n3219), .ZN(U3227)
         );
  NAND2_X1 U4029 ( .A1(n4298), .A2(n3222), .ZN(n3223) );
  OAI22_X1 U4030 ( .A1(n3225), .A2(n4663), .B1(n3224), .B2(n4353), .ZN(n3226)
         );
  INV_X1 U4031 ( .A(n3226), .ZN(n3233) );
  OAI22_X1 U4032 ( .A1(n4654), .A2(n3227), .B1(REG3_REG_3__SCAN_IN), .B2(n4651), .ZN(n3230) );
  NAND2_X1 U4033 ( .A1(n4654), .A2(n4291), .ZN(n4277) );
  NOR2_X1 U4034 ( .A1(n4277), .A2(n3228), .ZN(n3229) );
  AOI211_X1 U4035 ( .C1(n4282), .C2(n3231), .A(n3230), .B(n3229), .ZN(n3232)
         );
  OAI211_X1 U4036 ( .C1(n4328), .C2(n3234), .A(n3233), .B(n3232), .ZN(U3287)
         );
  OAI211_X1 U4037 ( .C1(n3237), .C2(n3236), .A(n3235), .B(n4554), .ZN(n3243)
         );
  OAI22_X1 U4038 ( .A1(n4531), .A2(n3249), .B1(n3288), .B2(n4546), .ZN(n3241)
         );
  INV_X1 U4039 ( .A(n3238), .ZN(n3239) );
  OAI21_X1 U4040 ( .B1(n4528), .B2(n3305), .A(n3239), .ZN(n3240) );
  NOR2_X1 U4041 ( .A1(n3241), .A2(n3240), .ZN(n3242) );
  OAI211_X1 U4042 ( .C1(n4563), .C2(n3300), .A(n3243), .B(n3242), .ZN(U3224)
         );
  INV_X1 U40430 ( .A(n3245), .ZN(n3910) );
  AND2_X1 U4044 ( .A1(n3910), .A2(n3923), .ZN(n3871) );
  XOR2_X1 U4045 ( .A(n3244), .B(n3871), .Z(n3306) );
  XOR2_X1 U4046 ( .A(n3246), .B(n3871), .Z(n3247) );
  AOI22_X1 U4047 ( .A1(n3247), .A2(n4342), .B1(n4362), .B2(n3997), .ZN(n3311)
         );
  AOI22_X1 U4048 ( .A1(n3999), .A2(n4291), .B1(n4380), .B2(n3303), .ZN(n3248)
         );
  OAI211_X1 U4049 ( .C1(n4441), .C2(n3306), .A(n3311), .B(n3248), .ZN(n3257)
         );
  OR2_X1 U4050 ( .A1(n3250), .A2(n3249), .ZN(n3251) );
  NAND2_X1 U4051 ( .A1(n3263), .A2(n3251), .ZN(n3299) );
  INV_X1 U4052 ( .A(REG0_REG_5__SCAN_IN), .ZN(n3252) );
  OAI22_X1 U4053 ( .A1(n4515), .A2(n3299), .B1(n4704), .B2(n3252), .ZN(n3253)
         );
  AOI21_X1 U4054 ( .B1(n3257), .B2(n4704), .A(n3253), .ZN(n3254) );
  INV_X1 U4055 ( .A(n3254), .ZN(U3477) );
  INV_X1 U4056 ( .A(REG1_REG_5__SCAN_IN), .ZN(n3255) );
  OAI22_X1 U4057 ( .A1(n4458), .A2(n3299), .B1(n4716), .B2(n3255), .ZN(n3256)
         );
  AOI21_X1 U4058 ( .B1(n3257), .B2(n4716), .A(n3256), .ZN(n3258) );
  INV_X1 U4059 ( .A(n3258), .ZN(U3523) );
  AND2_X1 U4060 ( .A1(n3913), .A2(n3921), .ZN(n3884) );
  XNOR2_X1 U4061 ( .A(n3259), .B(n3884), .ZN(n3276) );
  XNOR2_X1 U4062 ( .A(n3260), .B(n3884), .ZN(n3261) );
  AOI22_X1 U4063 ( .A1(n3261), .A2(n4342), .B1(n4362), .B2(n3995), .ZN(n3281)
         );
  AOI22_X1 U4064 ( .A1(n3998), .A2(n4291), .B1(n3272), .B2(n4380), .ZN(n3262)
         );
  OAI211_X1 U4065 ( .C1(n3276), .C2(n4441), .A(n3281), .B(n3262), .ZN(n3269)
         );
  NAND2_X1 U4066 ( .A1(n3263), .A2(n3272), .ZN(n3264) );
  NAND2_X1 U4067 ( .A1(n3290), .A2(n3264), .ZN(n3271) );
  INV_X1 U4068 ( .A(REG0_REG_6__SCAN_IN), .ZN(n4993) );
  OAI22_X1 U4069 ( .A1(n4515), .A2(n3271), .B1(n4704), .B2(n4993), .ZN(n3265)
         );
  AOI21_X1 U4070 ( .B1(n3269), .B2(n4704), .A(n3265), .ZN(n3266) );
  INV_X1 U4071 ( .A(n3266), .ZN(U3479) );
  OAI22_X1 U4072 ( .A1(n4458), .A2(n3271), .B1(n4716), .B2(n3267), .ZN(n3268)
         );
  AOI21_X1 U4073 ( .B1(n3269), .B2(n4716), .A(n3268), .ZN(n3270) );
  INV_X1 U4074 ( .A(n3270), .ZN(U3524) );
  INV_X1 U4075 ( .A(n3271), .ZN(n3279) );
  AOI22_X1 U4076 ( .A1(n4663), .A2(REG2_REG_6__SCAN_IN), .B1(n3321), .B2(n4643), .ZN(n3274) );
  NAND2_X1 U4077 ( .A1(n4282), .A2(n3272), .ZN(n3273) );
  OAI211_X1 U4078 ( .C1(n3275), .C2(n4277), .A(n3274), .B(n3273), .ZN(n3278)
         );
  NOR2_X1 U4079 ( .A1(n3276), .A2(n4353), .ZN(n3277) );
  AOI211_X1 U4080 ( .C1(n3279), .C2(n4657), .A(n3278), .B(n3277), .ZN(n3280)
         );
  OAI21_X1 U4081 ( .B1(n4663), .B2(n3281), .A(n3280), .ZN(U3284) );
  XNOR2_X1 U4082 ( .A(n3282), .B(n2261), .ZN(n4695) );
  INV_X1 U4083 ( .A(n4695), .ZN(n3298) );
  XNOR2_X1 U4084 ( .A(n3283), .B(n2261), .ZN(n3284) );
  NAND2_X1 U4085 ( .A1(n3284), .A2(n4342), .ZN(n3287) );
  NOR2_X1 U4086 ( .A1(n3570), .A2(n4433), .ZN(n3285) );
  AOI21_X1 U4087 ( .B1(n3994), .B2(n4362), .A(n3285), .ZN(n3286) );
  OAI211_X1 U4088 ( .C1(n3288), .C2(n4435), .A(n3287), .B(n3286), .ZN(n4692)
         );
  NAND2_X1 U4089 ( .A1(n4692), .A2(n4654), .ZN(n3297) );
  INV_X1 U4090 ( .A(n3331), .ZN(n3289) );
  AOI211_X1 U4091 ( .C1(n3291), .C2(n3290), .A(n4678), .B(n3289), .ZN(n4693)
         );
  INV_X1 U4092 ( .A(n4347), .ZN(n3295) );
  INV_X1 U4093 ( .A(n3572), .ZN(n3292) );
  OAI22_X1 U4094 ( .A1(n4654), .A2(n3293), .B1(n3292), .B2(n4651), .ZN(n3294)
         );
  AOI21_X1 U4095 ( .B1(n4693), .B2(n3295), .A(n3294), .ZN(n3296) );
  OAI211_X1 U4096 ( .C1(n3298), .C2(n4353), .A(n3297), .B(n3296), .ZN(U3283)
         );
  INV_X1 U4097 ( .A(n3299), .ZN(n3309) );
  OAI22_X1 U4098 ( .A1(n4654), .A2(n3301), .B1(n3300), .B2(n4651), .ZN(n3302)
         );
  AOI21_X1 U4099 ( .B1(n3303), .B2(n4282), .A(n3302), .ZN(n3304) );
  OAI21_X1 U4100 ( .B1(n3305), .B2(n4277), .A(n3304), .ZN(n3308) );
  NOR2_X1 U4101 ( .A1(n3306), .A2(n4353), .ZN(n3307) );
  AOI211_X1 U4102 ( .C1(n3309), .C2(n4657), .A(n3308), .B(n3307), .ZN(n3310)
         );
  OAI21_X1 U4103 ( .B1(n4663), .B2(n3311), .A(n3310), .ZN(U3285) );
  XNOR2_X1 U4104 ( .A(n3314), .B(n3313), .ZN(n3315) );
  XNOR2_X1 U4105 ( .A(n3312), .B(n3315), .ZN(n3323) );
  AOI21_X1 U4106 ( .B1(n3805), .B2(n3995), .A(n3316), .ZN(n3318) );
  NAND2_X1 U4107 ( .A1(n4556), .A2(n3998), .ZN(n3317) );
  OAI211_X1 U4108 ( .C1(n4531), .C2(n3319), .A(n3318), .B(n3317), .ZN(n3320)
         );
  AOI21_X1 U4109 ( .B1(n3811), .B2(n3321), .A(n3320), .ZN(n3322) );
  OAI21_X1 U4110 ( .B1(n3323), .B2(n3813), .A(n3322), .ZN(U3236) );
  AND2_X1 U4111 ( .A1(n3918), .A2(n3915), .ZN(n3869) );
  XNOR2_X1 U4112 ( .A(n3324), .B(n3869), .ZN(n4659) );
  INV_X1 U4113 ( .A(n4659), .ZN(n3330) );
  INV_X1 U4114 ( .A(n4298), .ZN(n4359) );
  XNOR2_X1 U4115 ( .A(n3325), .B(n3869), .ZN(n3328) );
  OAI22_X1 U4116 ( .A1(n3368), .A2(n4435), .B1(n3369), .B2(n4433), .ZN(n3326)
         );
  AOI21_X1 U4117 ( .B1(n4362), .B2(n3993), .A(n3326), .ZN(n3327) );
  OAI21_X1 U4118 ( .B1(n3328), .B2(n4366), .A(n3327), .ZN(n3329) );
  AOI21_X1 U4119 ( .B1(n4359), .B2(n4659), .A(n3329), .ZN(n4662) );
  OAI21_X1 U4120 ( .B1(n4696), .B2(n3330), .A(n4662), .ZN(n3335) );
  INV_X1 U4121 ( .A(n3335), .ZN(n3334) );
  AOI21_X1 U4122 ( .B1(n3332), .B2(n3331), .A(n3342), .ZN(n4656) );
  INV_X1 U4123 ( .A(n4515), .ZN(n3357) );
  AOI22_X1 U4124 ( .A1(n4656), .A2(n3357), .B1(n4702), .B2(REG0_REG_8__SCAN_IN), .ZN(n3333) );
  OAI21_X1 U4125 ( .B1(n3334), .B2(n4702), .A(n3333), .ZN(U3483) );
  INV_X1 U4126 ( .A(REG1_REG_8__SCAN_IN), .ZN(n3338) );
  NAND2_X1 U4127 ( .A1(n3335), .A2(n4716), .ZN(n3337) );
  INV_X1 U4128 ( .A(n4458), .ZN(n3359) );
  NAND2_X1 U4129 ( .A1(n4656), .A2(n3359), .ZN(n3336) );
  OAI211_X1 U4130 ( .C1(n4716), .C2(n3338), .A(n3337), .B(n3336), .ZN(U3526)
         );
  AND2_X1 U4131 ( .A1(n2296), .A2(n3917), .ZN(n3872) );
  XNOR2_X1 U4132 ( .A(n3339), .B(n3872), .ZN(n3340) );
  OAI22_X1 U4133 ( .A1(n3340), .A2(n4366), .B1(n3390), .B2(n4293), .ZN(n3354)
         );
  INV_X1 U4134 ( .A(n3354), .ZN(n3352) );
  XOR2_X1 U4135 ( .A(n3872), .B(n3341), .Z(n3356) );
  OR2_X1 U4136 ( .A1(n3342), .A2(n3379), .ZN(n3343) );
  AND2_X1 U4137 ( .A1(n3343), .A2(n3441), .ZN(n3360) );
  NAND2_X1 U4138 ( .A1(n3360), .A2(n4657), .ZN(n3349) );
  INV_X1 U4139 ( .A(REG2_REG_9__SCAN_IN), .ZN(n3344) );
  OAI22_X1 U4140 ( .A1(n3345), .A2(n4651), .B1(n3344), .B2(n4654), .ZN(n3346)
         );
  AOI21_X1 U4141 ( .B1(n4282), .B2(n3347), .A(n3346), .ZN(n3348) );
  OAI211_X1 U4142 ( .C1(n3353), .C2(n4277), .A(n3349), .B(n3348), .ZN(n3350)
         );
  AOI21_X1 U4143 ( .B1(n3356), .B2(n4273), .A(n3350), .ZN(n3351) );
  OAI21_X1 U4144 ( .B1(n4663), .B2(n3352), .A(n3351), .ZN(U3281) );
  OAI22_X1 U4145 ( .A1(n3353), .A2(n4435), .B1(n4433), .B2(n3379), .ZN(n3355)
         );
  AOI211_X1 U4146 ( .C1(n4694), .C2(n3356), .A(n3355), .B(n3354), .ZN(n3362)
         );
  AOI22_X1 U4147 ( .A1(n3360), .A2(n3357), .B1(REG0_REG_9__SCAN_IN), .B2(n4702), .ZN(n3358) );
  OAI21_X1 U4148 ( .B1(n3362), .B2(n4702), .A(n3358), .ZN(U3485) );
  AOI22_X1 U4149 ( .A1(n3360), .A2(n3359), .B1(REG1_REG_9__SCAN_IN), .B2(n4713), .ZN(n3361) );
  OAI21_X1 U4150 ( .B1(n3362), .B2(n4713), .A(n3361), .ZN(U3527) );
  INV_X1 U4151 ( .A(n3363), .ZN(n4652) );
  NOR2_X1 U4152 ( .A1(n2272), .A2(n3365), .ZN(n3366) );
  XNOR2_X1 U4153 ( .A(n3364), .B(n3366), .ZN(n3367) );
  NAND2_X1 U4154 ( .A1(n3367), .A2(n4554), .ZN(n3374) );
  OAI22_X1 U4155 ( .A1(n4531), .A2(n3369), .B1(n3368), .B2(n4528), .ZN(n3372)
         );
  OAI21_X1 U4156 ( .B1(n4546), .B2(n3447), .A(n3370), .ZN(n3371) );
  NOR2_X1 U4157 ( .A1(n3372), .A2(n3371), .ZN(n3373) );
  OAI211_X1 U4158 ( .C1(n4563), .C2(n4652), .A(n3374), .B(n3373), .ZN(U3218)
         );
  XOR2_X1 U4159 ( .A(n3376), .B(n3375), .Z(n3383) );
  NOR2_X1 U4160 ( .A1(STATE_REG_SCAN_IN), .A2(n2613), .ZN(n4578) );
  AOI21_X1 U4161 ( .B1(n3805), .B2(n3992), .A(n4578), .ZN(n3378) );
  NAND2_X1 U4162 ( .A1(n4556), .A2(n3994), .ZN(n3377) );
  OAI211_X1 U4163 ( .C1(n4531), .C2(n3379), .A(n3378), .B(n3377), .ZN(n3380)
         );
  AOI21_X1 U4164 ( .B1(n3811), .B2(n3381), .A(n3380), .ZN(n3382) );
  OAI21_X1 U4165 ( .B1(n3383), .B2(n3813), .A(n3382), .ZN(U3228) );
  OR2_X1 U4166 ( .A1(n3444), .A2(n3384), .ZN(n3386) );
  NAND2_X1 U4167 ( .A1(n3386), .A2(n3385), .ZN(n3388) );
  INV_X1 U4168 ( .A(n3387), .ZN(n3854) );
  XNOR2_X1 U4169 ( .A(n3388), .B(n3854), .ZN(n4697) );
  XNOR2_X1 U4170 ( .A(n3402), .B(n3854), .ZN(n3392) );
  AOI22_X1 U4171 ( .A1(n3990), .A2(n4362), .B1(n4380), .B2(n3417), .ZN(n3389)
         );
  OAI21_X1 U4172 ( .B1(n3390), .B2(n4435), .A(n3389), .ZN(n3391) );
  AOI21_X1 U4173 ( .B1(n3392), .B2(n4342), .A(n3391), .ZN(n3393) );
  OAI21_X1 U4174 ( .B1(n4697), .B2(n4298), .A(n3393), .ZN(n4698) );
  NAND2_X1 U4175 ( .A1(n4698), .A2(n4654), .ZN(n3398) );
  AOI21_X1 U4176 ( .B1(n3417), .B2(n3442), .A(n3405), .ZN(n4700) );
  INV_X1 U4177 ( .A(REG2_REG_11__SCAN_IN), .ZN(n3395) );
  INV_X1 U4178 ( .A(n3424), .ZN(n3394) );
  OAI22_X1 U4179 ( .A1(n4654), .A2(n3395), .B1(n3394), .B2(n4651), .ZN(n3396)
         );
  AOI21_X1 U4180 ( .B1(n4700), .B2(n4657), .A(n3396), .ZN(n3397) );
  OAI211_X1 U4181 ( .C1(n4697), .C2(n4309), .A(n3398), .B(n3397), .ZN(U3279)
         );
  INV_X1 U4182 ( .A(n3399), .ZN(n3400) );
  AOI21_X1 U4183 ( .B1(n3402), .B2(n3401), .A(n3400), .ZN(n3482) );
  AND2_X1 U4184 ( .A1(n3481), .A2(n3479), .ZN(n3870) );
  XNOR2_X1 U4185 ( .A(n3482), .B(n3870), .ZN(n3403) );
  OAI22_X1 U4186 ( .A1(n3403), .A2(n4366), .B1(n3704), .B2(n4293), .ZN(n3469)
         );
  INV_X1 U4187 ( .A(n3469), .ZN(n3414) );
  XOR2_X1 U4188 ( .A(n3870), .B(n3404), .Z(n3471) );
  NOR2_X1 U4189 ( .A1(n3405), .A2(n3537), .ZN(n3406) );
  OR2_X1 U4190 ( .A1(n3489), .A2(n3406), .ZN(n3477) );
  INV_X1 U4191 ( .A(REG2_REG_12__SCAN_IN), .ZN(n3408) );
  INV_X1 U4192 ( .A(n3407), .ZN(n3543) );
  OAI22_X1 U4193 ( .A1(n4654), .A2(n3408), .B1(n3543), .B2(n4651), .ZN(n3410)
         );
  NOR2_X1 U4194 ( .A1(n4277), .A2(n3538), .ZN(n3409) );
  AOI211_X1 U4195 ( .C1(n4282), .C2(n3525), .A(n3410), .B(n3409), .ZN(n3411)
         );
  OAI21_X1 U4196 ( .B1(n3477), .B2(n4328), .A(n3411), .ZN(n3412) );
  AOI21_X1 U4197 ( .B1(n3471), .B2(n4273), .A(n3412), .ZN(n3413) );
  OAI21_X1 U4198 ( .B1(n4663), .B2(n3414), .A(n3413), .ZN(U3278) );
  INV_X1 U4199 ( .A(n3618), .ZN(n3628) );
  AOI22_X1 U4200 ( .A1(n3991), .A2(n3665), .B1(n3628), .B2(n3417), .ZN(n3520)
         );
  OAI22_X1 U4201 ( .A1(n3538), .A2(n3678), .B1(n3677), .B2(n3422), .ZN(n3418)
         );
  XNOR2_X1 U4202 ( .A(n2455), .B(n3523), .ZN(n3419) );
  XNOR2_X1 U4203 ( .A(n3521), .B(n3419), .ZN(n3426) );
  AND2_X1 U4204 ( .A1(U3149), .A2(REG3_REG_11__SCAN_IN), .ZN(n4600) );
  AOI21_X1 U4205 ( .B1(n4556), .B2(n3992), .A(n4600), .ZN(n3421) );
  NAND2_X1 U4206 ( .A1(n3805), .A2(n3990), .ZN(n3420) );
  OAI211_X1 U4207 ( .C1(n4531), .C2(n3422), .A(n3421), .B(n3420), .ZN(n3423)
         );
  AOI21_X1 U4208 ( .B1(n3811), .B2(n3424), .A(n3423), .ZN(n3425) );
  OAI21_X1 U4209 ( .B1(n3426), .B2(n3813), .A(n3425), .ZN(U3233) );
  OAI21_X1 U4210 ( .B1(n3429), .B2(n3428), .A(n3427), .ZN(n4447) );
  OAI21_X1 U4211 ( .B1(n3886), .B2(n3820), .A(n3430), .ZN(n3431) );
  NAND2_X1 U4212 ( .A1(n3431), .A2(n4342), .ZN(n3433) );
  AOI22_X1 U4213 ( .A1(n3987), .A2(n4362), .B1(n4380), .B2(n3435), .ZN(n3432)
         );
  OAI211_X1 U4214 ( .C1(n3704), .C2(n4435), .A(n3433), .B(n3432), .ZN(n3434)
         );
  AOI21_X1 U4215 ( .B1(n4447), .B2(n4359), .A(n3434), .ZN(n4451) );
  NAND2_X1 U4216 ( .A1(n3488), .A2(n3435), .ZN(n4448) );
  AND3_X1 U4217 ( .A1(n4449), .A2(n4657), .A3(n4448), .ZN(n3439) );
  INV_X1 U4218 ( .A(REG2_REG_14__SCAN_IN), .ZN(n3437) );
  INV_X1 U4219 ( .A(n3436), .ZN(n3710) );
  OAI22_X1 U4220 ( .A1(n4654), .A2(n3437), .B1(n3710), .B2(n4651), .ZN(n3438)
         );
  AOI211_X1 U4221 ( .C1(n4447), .C2(n4658), .A(n3439), .B(n3438), .ZN(n3440)
         );
  OAI21_X1 U4222 ( .B1(n4451), .B2(n4663), .A(n3440), .ZN(U3276) );
  INV_X1 U4223 ( .A(n3441), .ZN(n3443) );
  OAI21_X1 U4224 ( .B1(n3443), .B2(n3446), .A(n3442), .ZN(n4645) );
  INV_X1 U4225 ( .A(REG0_REG_10__SCAN_IN), .ZN(n3453) );
  XNOR2_X1 U4226 ( .A(n3444), .B(n3856), .ZN(n4647) );
  XOR2_X1 U4227 ( .A(n3445), .B(n3856), .Z(n3450) );
  OAI22_X1 U4228 ( .A1(n3447), .A2(n4435), .B1(n3446), .B2(n4433), .ZN(n3448)
         );
  AOI21_X1 U4229 ( .B1(n4362), .B2(n3991), .A(n3448), .ZN(n3449) );
  OAI21_X1 U4230 ( .B1(n3450), .B2(n4366), .A(n3449), .ZN(n3451) );
  AOI21_X1 U4231 ( .B1(n4359), .B2(n4647), .A(n3451), .ZN(n4650) );
  INV_X1 U4232 ( .A(n4650), .ZN(n3452) );
  AOI21_X1 U4233 ( .B1(n4690), .B2(n4647), .A(n3452), .ZN(n3455) );
  MUX2_X1 U4234 ( .A(n3453), .B(n3455), .S(n4704), .Z(n3454) );
  OAI21_X1 U4235 ( .B1(n4645), .B2(n4515), .A(n3454), .ZN(U3487) );
  INV_X1 U4236 ( .A(REG1_REG_10__SCAN_IN), .ZN(n3456) );
  MUX2_X1 U4237 ( .A(n3456), .B(n3455), .S(n4716), .Z(n3457) );
  OAI21_X1 U4238 ( .B1(n4645), .B2(n4458), .A(n3457), .ZN(U3528) );
  XNOR2_X1 U4239 ( .A(n3458), .B(n3883), .ZN(n3513) );
  INV_X1 U4240 ( .A(n3513), .ZN(n3468) );
  XNOR2_X1 U4241 ( .A(n3459), .B(n3883), .ZN(n3460) );
  OAI22_X1 U4242 ( .A1(n3460), .A2(n4366), .B1(n4436), .B2(n4293), .ZN(n3512)
         );
  INV_X1 U4243 ( .A(n4449), .ZN(n3462) );
  INV_X1 U4244 ( .A(n3504), .ZN(n3461) );
  OAI21_X1 U4245 ( .B1(n3462), .B2(n3808), .A(n3461), .ZN(n3519) );
  AOI22_X1 U4246 ( .A1(n4663), .A2(REG2_REG_15__SCAN_IN), .B1(n3810), .B2(
        n4643), .ZN(n3463) );
  OAI21_X1 U4247 ( .B1(n3579), .B2(n4277), .A(n3463), .ZN(n3464) );
  AOI21_X1 U4248 ( .B1(n3584), .B2(n4282), .A(n3464), .ZN(n3465) );
  OAI21_X1 U4249 ( .B1(n3519), .B2(n4328), .A(n3465), .ZN(n3466) );
  AOI21_X1 U4250 ( .B1(n3512), .B2(n4654), .A(n3466), .ZN(n3467) );
  OAI21_X1 U4251 ( .B1(n3468), .B2(n4353), .A(n3467), .ZN(U3275) );
  INV_X1 U4252 ( .A(REG0_REG_12__SCAN_IN), .ZN(n3472) );
  OAI22_X1 U4253 ( .A1(n3538), .A2(n4435), .B1(n3537), .B2(n4433), .ZN(n3470)
         );
  AOI211_X1 U4254 ( .C1(n4694), .C2(n3471), .A(n3470), .B(n3469), .ZN(n3474)
         );
  MUX2_X1 U4255 ( .A(n3472), .B(n3474), .S(n4704), .Z(n3473) );
  OAI21_X1 U4256 ( .B1(n3477), .B2(n4515), .A(n3473), .ZN(U3491) );
  INV_X1 U4257 ( .A(REG1_REG_12__SCAN_IN), .ZN(n3475) );
  MUX2_X1 U4258 ( .A(n3475), .B(n3474), .S(n4716), .Z(n3476) );
  OAI21_X1 U4259 ( .B1(n3477), .B2(n4458), .A(n3476), .ZN(U3530) );
  OAI22_X1 U4260 ( .A1(n3579), .A2(n4293), .B1(n4433), .B2(n3560), .ZN(n3486)
         );
  XNOR2_X1 U4261 ( .A(n3989), .B(n3478), .ZN(n3876) );
  INV_X1 U4262 ( .A(n3479), .ZN(n3480) );
  AOI21_X1 U4263 ( .B1(n3482), .B2(n3481), .A(n3480), .ZN(n3483) );
  XOR2_X1 U4264 ( .A(n3876), .B(n3483), .Z(n3484) );
  NOR2_X1 U4265 ( .A1(n3484), .A2(n4366), .ZN(n3485) );
  AOI211_X1 U4266 ( .C1(n4291), .C2(n3990), .A(n3486), .B(n3485), .ZN(n4453)
         );
  XNOR2_X1 U4267 ( .A(n3487), .B(n3876), .ZN(n4455) );
  OAI21_X1 U4268 ( .B1(n3489), .B2(n3560), .A(n3488), .ZN(n4516) );
  NOR2_X1 U4269 ( .A1(n3490), .A2(n4651), .ZN(n3491) );
  AOI21_X1 U4270 ( .B1(n4663), .B2(REG2_REG_13__SCAN_IN), .A(n3491), .ZN(n3492) );
  OAI21_X1 U4271 ( .B1(n4516), .B2(n4328), .A(n3492), .ZN(n3493) );
  AOI21_X1 U4272 ( .B1(n4455), .B2(n4273), .A(n3493), .ZN(n3494) );
  OAI21_X1 U4273 ( .B1(n4453), .B2(n4663), .A(n3494), .ZN(U3277) );
  XNOR2_X1 U4274 ( .A(n3495), .B(n3502), .ZN(n3500) );
  NAND2_X1 U4275 ( .A1(n4380), .A2(n3496), .ZN(n3498) );
  NAND2_X1 U4276 ( .A1(n3987), .A2(n4291), .ZN(n3497) );
  OAI211_X1 U4277 ( .C1(n4533), .C2(n4293), .A(n3498), .B(n3497), .ZN(n3499)
         );
  AOI21_X1 U4278 ( .B1(n3500), .B2(n4342), .A(n3499), .ZN(n4443) );
  OAI21_X1 U4279 ( .B1(n3503), .B2(n3502), .A(n3501), .ZN(n4442) );
  OR2_X1 U4280 ( .A1(n4442), .A2(n4353), .ZN(n3510) );
  NOR2_X1 U4281 ( .A1(n3504), .A2(n4530), .ZN(n3505) );
  OR2_X1 U4282 ( .A1(n3546), .A2(n3505), .ZN(n4508) );
  INV_X1 U4283 ( .A(n4508), .ZN(n3508) );
  INV_X1 U4284 ( .A(REG2_REG_16__SCAN_IN), .ZN(n3506) );
  OAI22_X1 U4285 ( .A1(n4654), .A2(n3506), .B1(n4543), .B2(n4651), .ZN(n3507)
         );
  AOI21_X1 U4286 ( .B1(n3508), .B2(n4657), .A(n3507), .ZN(n3509) );
  OAI211_X1 U4287 ( .C1(n4663), .C2(n4443), .A(n3510), .B(n3509), .ZN(U3274)
         );
  INV_X1 U4288 ( .A(REG0_REG_15__SCAN_IN), .ZN(n3514) );
  OAI22_X1 U4289 ( .A1(n3579), .A2(n4435), .B1(n3808), .B2(n4433), .ZN(n3511)
         );
  AOI211_X1 U4290 ( .C1(n3513), .C2(n4694), .A(n3512), .B(n3511), .ZN(n3516)
         );
  MUX2_X1 U4291 ( .A(n3514), .B(n3516), .S(n4704), .Z(n3515) );
  OAI21_X1 U4292 ( .B1(n3519), .B2(n4515), .A(n3515), .ZN(U3497) );
  INV_X1 U4293 ( .A(REG1_REG_15__SCAN_IN), .ZN(n3517) );
  MUX2_X1 U4294 ( .A(n3517), .B(n3516), .S(n4716), .Z(n3518) );
  OAI21_X1 U4295 ( .B1(n4458), .B2(n3519), .A(n3518), .ZN(U3533) );
  NAND2_X1 U4296 ( .A1(n3521), .A2(n3520), .ZN(n3524) );
  NAND2_X1 U4297 ( .A1(n3990), .A2(n3636), .ZN(n3527) );
  NAND2_X1 U4298 ( .A1(n2926), .A2(n3525), .ZN(n3526) );
  NAND2_X1 U4299 ( .A1(n3527), .A2(n3526), .ZN(n3528) );
  XNOR2_X1 U4300 ( .A(n3528), .B(n3661), .ZN(n3533) );
  INV_X1 U4301 ( .A(n3533), .ZN(n3531) );
  NOR2_X1 U4302 ( .A1(n3663), .A2(n3537), .ZN(n3529) );
  AOI21_X1 U4303 ( .B1(n3665), .B2(n3990), .A(n3529), .ZN(n3532) );
  INV_X1 U4304 ( .A(n3532), .ZN(n3530) );
  NAND2_X1 U4305 ( .A1(n3531), .A2(n3530), .ZN(n3554) );
  INV_X1 U4306 ( .A(n3554), .ZN(n3534) );
  AND2_X1 U4307 ( .A1(n3533), .A2(n3532), .ZN(n3553) );
  NOR2_X1 U4308 ( .A1(n3534), .A2(n3553), .ZN(n3535) );
  XNOR2_X1 U4309 ( .A(n3555), .B(n3535), .ZN(n3536) );
  NAND2_X1 U4310 ( .A1(n3536), .A2(n4554), .ZN(n3542) );
  OAI22_X1 U4311 ( .A1(n4531), .A2(n3537), .B1(n3704), .B2(n4546), .ZN(n3540)
         );
  NAND2_X1 U4312 ( .A1(REG3_REG_12__SCAN_IN), .A2(U3149), .ZN(n4053) );
  OAI21_X1 U4313 ( .B1(n4528), .B2(n3538), .A(n4053), .ZN(n3539) );
  NOR2_X1 U4314 ( .A1(n3540), .A2(n3539), .ZN(n3541) );
  OAI211_X1 U4315 ( .C1(n4563), .C2(n3543), .A(n3542), .B(n3541), .ZN(U3221)
         );
  XNOR2_X1 U4316 ( .A(n3544), .B(n3867), .ZN(n4439) );
  INV_X1 U4317 ( .A(n4439), .ZN(n3552) );
  XNOR2_X1 U4318 ( .A(n4231), .B(n3867), .ZN(n3545) );
  OAI22_X1 U4319 ( .A1(n3545), .A2(n4366), .B1(n4325), .B2(n4293), .ZN(n4438)
         );
  OAI21_X1 U4320 ( .B1(n3546), .B2(n4434), .A(n4344), .ZN(n4506) );
  AOI22_X1 U4321 ( .A1(n4663), .A2(REG2_REG_17__SCAN_IN), .B1(n3762), .B2(
        n4643), .ZN(n3547) );
  OAI21_X1 U4322 ( .B1(n4436), .B2(n4277), .A(n3547), .ZN(n3548) );
  AOI21_X1 U4323 ( .B1(n3598), .B2(n4282), .A(n3548), .ZN(n3549) );
  OAI21_X1 U4324 ( .B1(n4506), .B2(n4328), .A(n3549), .ZN(n3550) );
  AOI21_X1 U4325 ( .B1(n4438), .B2(n4654), .A(n3550), .ZN(n3551) );
  OAI21_X1 U4326 ( .B1(n3552), .B2(n4353), .A(n3551), .ZN(U3273) );
  OAI22_X1 U4327 ( .A1(n3704), .A2(n3618), .B1(n3677), .B2(n3560), .ZN(n3556)
         );
  OAI22_X1 U4328 ( .A1(n3704), .A2(n3674), .B1(n3663), .B2(n3560), .ZN(n3577)
         );
  XNOR2_X1 U4329 ( .A(n3575), .B(n3577), .ZN(n3557) );
  XNOR2_X1 U4330 ( .A(n3576), .B(n3557), .ZN(n3564) );
  NOR2_X1 U4331 ( .A1(STATE_REG_SCAN_IN), .A2(n2659), .ZN(n4070) );
  AOI21_X1 U4332 ( .B1(n4556), .B2(n3990), .A(n4070), .ZN(n3559) );
  NAND2_X1 U4333 ( .A1(n3805), .A2(n3988), .ZN(n3558) );
  OAI211_X1 U4334 ( .C1(n4531), .C2(n3560), .A(n3559), .B(n3558), .ZN(n3561)
         );
  AOI21_X1 U4335 ( .B1(n3811), .B2(n3562), .A(n3561), .ZN(n3563) );
  OAI21_X1 U4336 ( .B1(n3564), .B2(n3813), .A(n3563), .ZN(U3231) );
  XNOR2_X1 U4337 ( .A(n3566), .B(n3565), .ZN(n3574) );
  AOI21_X1 U4338 ( .B1(n3805), .B2(n3994), .A(n3567), .ZN(n3569) );
  NAND2_X1 U4339 ( .A1(n4556), .A2(n3997), .ZN(n3568) );
  OAI211_X1 U4340 ( .C1(n4531), .C2(n3570), .A(n3569), .B(n3568), .ZN(n3571)
         );
  AOI21_X1 U4341 ( .B1(n3811), .B2(n3572), .A(n3571), .ZN(n3573) );
  OAI21_X1 U4342 ( .B1(n3574), .B2(n3813), .A(n3573), .ZN(U3210) );
  OAI22_X1 U4343 ( .A1(n3579), .A2(n3678), .B1(n3677), .B2(n3705), .ZN(n3578)
         );
  XNOR2_X1 U4344 ( .A(n3578), .B(n2232), .ZN(n3581) );
  OAI22_X1 U4345 ( .A1(n3579), .A2(n3674), .B1(n3663), .B2(n3705), .ZN(n3580)
         );
  NAND2_X1 U4346 ( .A1(n3581), .A2(n3580), .ZN(n3699) );
  OR2_X1 U4347 ( .A1(n3581), .A2(n3580), .ZN(n3700) );
  NAND2_X1 U4348 ( .A1(n3582), .A2(n3700), .ZN(n3588) );
  OAI22_X1 U4349 ( .A1(n4529), .A2(n3663), .B1(n3677), .B2(n3808), .ZN(n3583)
         );
  XOR2_X1 U4350 ( .A(n3675), .B(n3583), .Z(n3589) );
  NAND2_X1 U4351 ( .A1(n3588), .A2(n3589), .ZN(n3803) );
  NAND2_X1 U4352 ( .A1(n3665), .A2(n3987), .ZN(n3587) );
  NAND2_X1 U4353 ( .A1(n3585), .A2(n3584), .ZN(n3586) );
  NAND2_X1 U4354 ( .A1(n3587), .A2(n3586), .ZN(n4536) );
  INV_X1 U4355 ( .A(n3588), .ZN(n3591) );
  NAND2_X1 U4356 ( .A1(n3591), .A2(n3590), .ZN(n3802) );
  OAI22_X1 U4357 ( .A1(n4436), .A2(n3678), .B1(n3677), .B2(n4530), .ZN(n3592)
         );
  XNOR2_X1 U4358 ( .A(n3592), .B(n3675), .ZN(n3594) );
  OAI22_X1 U4359 ( .A1(n4436), .A2(n3674), .B1(n3663), .B2(n4530), .ZN(n3593)
         );
  NOR2_X1 U4360 ( .A1(n3594), .A2(n3593), .ZN(n3595) );
  INV_X1 U4361 ( .A(n3595), .ZN(n3596) );
  OAI22_X1 U4362 ( .A1(n4533), .A2(n3678), .B1(n3677), .B2(n4434), .ZN(n3597)
         );
  XNOR2_X1 U4363 ( .A(n3597), .B(n3675), .ZN(n3601) );
  OR2_X1 U4364 ( .A1(n3674), .A2(n4533), .ZN(n3600) );
  NAND2_X1 U4365 ( .A1(n3636), .A2(n3598), .ZN(n3599) );
  NAND2_X1 U4366 ( .A1(n3600), .A2(n3599), .ZN(n3602) );
  NAND2_X1 U4367 ( .A1(n3601), .A2(n3602), .ZN(n3757) );
  INV_X1 U4368 ( .A(n3601), .ZN(n3604) );
  INV_X1 U4369 ( .A(n3602), .ZN(n3603) );
  NAND2_X1 U4370 ( .A1(n3604), .A2(n3603), .ZN(n3756) );
  OAI22_X1 U4371 ( .A1(n4325), .A2(n3663), .B1(n3677), .B2(n4346), .ZN(n3605)
         );
  XNOR2_X1 U4372 ( .A(n3605), .B(n2232), .ZN(n3608) );
  OR2_X1 U4373 ( .A1(n3674), .A2(n4325), .ZN(n3607) );
  NAND2_X1 U4374 ( .A1(n3636), .A2(n4558), .ZN(n3606) );
  NAND2_X1 U4375 ( .A1(n3607), .A2(n3606), .ZN(n3609) );
  NAND2_X1 U4376 ( .A1(n3608), .A2(n3609), .ZN(n4548) );
  INV_X1 U4377 ( .A(n3608), .ZN(n3611) );
  INV_X1 U4378 ( .A(n3609), .ZN(n3610) );
  NAND2_X1 U4379 ( .A1(n3611), .A2(n3610), .ZN(n4549) );
  OAI22_X1 U4380 ( .A1(n4545), .A2(n3674), .B1(n3663), .B2(n4327), .ZN(n3614)
         );
  OAI22_X1 U4381 ( .A1(n4545), .A2(n3663), .B1(n3677), .B2(n4327), .ZN(n3612)
         );
  XNOR2_X1 U4382 ( .A(n3612), .B(n3675), .ZN(n3613) );
  XOR2_X1 U4383 ( .A(n3614), .B(n3613), .Z(n3724) );
  NAND2_X1 U4384 ( .A1(n3723), .A2(n3724), .ZN(n3722) );
  INV_X1 U4385 ( .A(n3613), .ZN(n3616) );
  INV_X1 U4386 ( .A(n3614), .ZN(n3615) );
  NAND2_X1 U4387 ( .A1(n3616), .A2(n3615), .ZN(n3617) );
  NAND2_X1 U4388 ( .A1(n3722), .A2(n3617), .ZN(n3730) );
  NAND2_X1 U4389 ( .A1(n4322), .A2(n3636), .ZN(n3620) );
  NAND2_X1 U4390 ( .A1(n2926), .A2(n4290), .ZN(n3619) );
  NAND2_X1 U4391 ( .A1(n3620), .A2(n3619), .ZN(n3621) );
  XNOR2_X1 U4392 ( .A(n3621), .B(n3661), .ZN(n3632) );
  INV_X1 U4393 ( .A(n3632), .ZN(n3624) );
  NOR2_X1 U4394 ( .A1(n3663), .A2(n4301), .ZN(n3622) );
  AOI21_X1 U4395 ( .B1(n3665), .B2(n4322), .A(n3622), .ZN(n3631) );
  INV_X1 U4396 ( .A(n3631), .ZN(n3623) );
  NAND2_X1 U4397 ( .A1(n3624), .A2(n3623), .ZN(n3775) );
  NAND2_X1 U4398 ( .A1(n4258), .A2(n3636), .ZN(n3626) );
  NAND2_X1 U4399 ( .A1(n2926), .A2(n4281), .ZN(n3625) );
  NAND2_X1 U4400 ( .A1(n3626), .A2(n3625), .ZN(n3627) );
  XNOR2_X1 U4401 ( .A(n3627), .B(n2232), .ZN(n3733) );
  NAND2_X1 U4402 ( .A1(n4258), .A2(n3665), .ZN(n3630) );
  NAND2_X1 U4403 ( .A1(n3628), .A2(n4281), .ZN(n3629) );
  NAND2_X1 U4404 ( .A1(n3630), .A2(n3629), .ZN(n3732) );
  NAND2_X1 U4405 ( .A1(n3632), .A2(n3631), .ZN(n3774) );
  OAI21_X1 U4406 ( .B1(n3733), .B2(n3732), .A(n3774), .ZN(n3633) );
  INV_X1 U4407 ( .A(n3733), .ZN(n3635) );
  INV_X1 U4408 ( .A(n3732), .ZN(n3634) );
  NOR2_X1 U4409 ( .A1(n3635), .A2(n3634), .ZN(n3782) );
  AOI22_X1 U4410 ( .A1(n4268), .A2(n3636), .B1(n2926), .B2(n4257), .ZN(n3637)
         );
  XNOR2_X1 U4411 ( .A(n3637), .B(n3675), .ZN(n3639) );
  AOI22_X1 U4412 ( .A1(n4268), .A2(n3665), .B1(n3636), .B2(n4257), .ZN(n3640)
         );
  XNOR2_X1 U4413 ( .A(n3639), .B(n3640), .ZN(n3785) );
  OR2_X1 U4414 ( .A1(n3782), .A2(n3785), .ZN(n3638) );
  INV_X1 U4415 ( .A(n3639), .ZN(n3642) );
  INV_X1 U4416 ( .A(n3640), .ZN(n3641) );
  NOR2_X1 U4417 ( .A1(n3642), .A2(n3641), .ZN(n3713) );
  NAND2_X1 U4418 ( .A1(n3984), .A2(n3636), .ZN(n3644) );
  NAND2_X1 U4419 ( .A1(n2926), .A2(n4240), .ZN(n3643) );
  NAND2_X1 U4420 ( .A1(n3644), .A2(n3643), .ZN(n3645) );
  XNOR2_X1 U4421 ( .A(n3645), .B(n3661), .ZN(n3648) );
  NOR2_X1 U4422 ( .A1(n3663), .A2(n4225), .ZN(n3646) );
  AOI21_X1 U4423 ( .B1(n3984), .B2(n3665), .A(n3646), .ZN(n3647) );
  XNOR2_X1 U4424 ( .A(n3648), .B(n3647), .ZN(n3712) );
  NOR2_X1 U4425 ( .A1(n3648), .A2(n3647), .ZN(n3650) );
  OAI22_X1 U4426 ( .A1(n4243), .A2(n3674), .B1(n3663), .B2(n4399), .ZN(n3651)
         );
  OAI22_X1 U4427 ( .A1(n4243), .A2(n3618), .B1(n3677), .B2(n4399), .ZN(n3649)
         );
  XNOR2_X1 U4428 ( .A(n3649), .B(n2232), .ZN(n3767) );
  NAND2_X1 U4429 ( .A1(n3765), .A2(n3767), .ZN(n3652) );
  NAND2_X1 U4430 ( .A1(n3652), .A2(n3766), .ZN(n3743) );
  NAND2_X1 U4431 ( .A1(n4178), .A2(n3636), .ZN(n3654) );
  NAND2_X1 U4432 ( .A1(n2926), .A2(n2284), .ZN(n3653) );
  NAND2_X1 U4433 ( .A1(n3654), .A2(n3653), .ZN(n3655) );
  XNOR2_X1 U4434 ( .A(n3655), .B(n3661), .ZN(n3658) );
  NOR2_X1 U4435 ( .A1(n3663), .A2(n4197), .ZN(n3656) );
  AOI21_X1 U4436 ( .B1(n4178), .B2(n3665), .A(n3656), .ZN(n3657) );
  NAND2_X1 U4437 ( .A1(n3658), .A2(n3657), .ZN(n3744) );
  OR2_X1 U4438 ( .A1(n3658), .A2(n3657), .ZN(n3745) );
  NAND2_X1 U4439 ( .A1(n4194), .A2(n3636), .ZN(n3660) );
  NAND2_X1 U4440 ( .A1(n2926), .A2(n4176), .ZN(n3659) );
  NAND2_X1 U4441 ( .A1(n3660), .A2(n3659), .ZN(n3662) );
  XNOR2_X1 U4442 ( .A(n3662), .B(n3661), .ZN(n3667) );
  NOR2_X1 U4443 ( .A1(n3663), .A2(n4183), .ZN(n3664) );
  AOI21_X1 U4444 ( .B1(n4194), .B2(n3665), .A(n3664), .ZN(n3666) );
  NAND2_X1 U4445 ( .A1(n3667), .A2(n3666), .ZN(n3793) );
  OAI22_X1 U4446 ( .A1(n4146), .A2(n3618), .B1(n3677), .B2(n4384), .ZN(n3669)
         );
  XNOR2_X1 U4447 ( .A(n3669), .B(n3675), .ZN(n3671) );
  OAI22_X1 U4448 ( .A1(n4146), .A2(n3674), .B1(n3663), .B2(n4384), .ZN(n3670)
         );
  INV_X1 U4449 ( .A(n3670), .ZN(n3673) );
  INV_X1 U4450 ( .A(n3671), .ZN(n3672) );
  OAI22_X1 U4451 ( .A1(n4131), .A2(n3674), .B1(n3663), .B2(n3686), .ZN(n3676)
         );
  XNOR2_X1 U4452 ( .A(n3676), .B(n2232), .ZN(n3680) );
  OAI22_X1 U4453 ( .A1(n4131), .A2(n3678), .B1(n3677), .B2(n3686), .ZN(n3679)
         );
  XNOR2_X1 U4454 ( .A(n3680), .B(n3679), .ZN(n3681) );
  XNOR2_X1 U4455 ( .A(n3682), .B(n3681), .ZN(n3683) );
  NAND2_X1 U4456 ( .A1(n3683), .A2(n4554), .ZN(n3690) );
  INV_X1 U4457 ( .A(n3684), .ZN(n4142) );
  INV_X1 U4458 ( .A(n3981), .ZN(n3837) );
  OAI22_X1 U4459 ( .A1(n3837), .A2(n4546), .B1(STATE_REG_SCAN_IN), .B2(n3685), 
        .ZN(n3688) );
  OAI22_X1 U4460 ( .A1(n4146), .A2(n4528), .B1(n4531), .B2(n3686), .ZN(n3687)
         );
  AOI211_X1 U4461 ( .C1(n4142), .C2(n3811), .A(n3688), .B(n3687), .ZN(n3689)
         );
  NAND2_X1 U4462 ( .A1(n3690), .A2(n3689), .ZN(U3217) );
  XNOR2_X1 U4463 ( .A(n3691), .B(n3692), .ZN(n3698) );
  INV_X1 U4464 ( .A(n3693), .ZN(n4163) );
  OAI22_X1 U4465 ( .A1(n4385), .A2(n4528), .B1(n4531), .B2(n4384), .ZN(n3696)
         );
  OAI22_X1 U4466 ( .A1(n4131), .A2(n4546), .B1(STATE_REG_SCAN_IN), .B2(n3694), 
        .ZN(n3695) );
  AOI211_X1 U4467 ( .C1(n4163), .C2(n3811), .A(n3696), .B(n3695), .ZN(n3697)
         );
  OAI21_X1 U4468 ( .B1(n3698), .B2(n3813), .A(n3697), .ZN(U3211) );
  NAND2_X1 U4469 ( .A1(n3700), .A2(n3699), .ZN(n3702) );
  XOR2_X1 U4470 ( .A(n3702), .B(n3701), .Z(n3703) );
  NAND2_X1 U4471 ( .A1(n3703), .A2(n4554), .ZN(n3709) );
  OAI22_X1 U4472 ( .A1(n4531), .A2(n3705), .B1(n3704), .B2(n4528), .ZN(n3707)
         );
  NAND2_X1 U4473 ( .A1(REG3_REG_14__SCAN_IN), .A2(U3149), .ZN(n4602) );
  OAI21_X1 U4474 ( .B1(n4546), .B2(n4529), .A(n4602), .ZN(n3706) );
  NOR2_X1 U4475 ( .A1(n3707), .A2(n3706), .ZN(n3708) );
  OAI211_X1 U4476 ( .C1(n4563), .C2(n3710), .A(n3709), .B(n3708), .ZN(U3212)
         );
  INV_X1 U4477 ( .A(n3711), .ZN(n4244) );
  OAI21_X1 U4478 ( .B1(n2242), .B2(n3713), .A(n3712), .ZN(n3716) );
  INV_X1 U4479 ( .A(n3714), .ZN(n3715) );
  NAND3_X1 U4480 ( .A1(n3716), .A2(n3715), .A3(n4554), .ZN(n3720) );
  OAI22_X1 U4481 ( .A1(n4531), .A2(n4225), .B1(n4243), .B2(n4546), .ZN(n3718)
         );
  INV_X1 U4482 ( .A(n4268), .ZN(n3738) );
  INV_X1 U4483 ( .A(REG3_REG_23__SCAN_IN), .ZN(n5070) );
  OAI22_X1 U4484 ( .A1(n4528), .A2(n3738), .B1(STATE_REG_SCAN_IN), .B2(n5070), 
        .ZN(n3717) );
  NOR2_X1 U4485 ( .A1(n3718), .A2(n3717), .ZN(n3719) );
  OAI211_X1 U4486 ( .C1(n4563), .C2(n4244), .A(n3720), .B(n3719), .ZN(U3213)
         );
  INV_X1 U4487 ( .A(n3721), .ZN(n4329) );
  OAI21_X1 U4488 ( .B1(n3724), .B2(n3723), .A(n3722), .ZN(n3725) );
  NAND2_X1 U4489 ( .A1(n3725), .A2(n4554), .ZN(n3729) );
  INV_X1 U4490 ( .A(n4322), .ZN(n4416) );
  OAI22_X1 U4491 ( .A1(n4531), .A2(n4327), .B1(n4416), .B2(n4546), .ZN(n3727)
         );
  NAND2_X1 U4492 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n4115) );
  OAI21_X1 U4493 ( .B1(n4528), .B2(n4325), .A(n4115), .ZN(n3726) );
  NOR2_X1 U4494 ( .A1(n3727), .A2(n3726), .ZN(n3728) );
  OAI211_X1 U4495 ( .C1(n4563), .C2(n4329), .A(n3729), .B(n3728), .ZN(U3216)
         );
  INV_X1 U4496 ( .A(n3774), .ZN(n3731) );
  OAI21_X1 U4497 ( .B1(n3730), .B2(n3731), .A(n3775), .ZN(n3735) );
  XNOR2_X1 U4498 ( .A(n3733), .B(n3732), .ZN(n3734) );
  XNOR2_X1 U4499 ( .A(n3735), .B(n3734), .ZN(n3736) );
  NAND2_X1 U4500 ( .A1(n3736), .A2(n4554), .ZN(n3742) );
  OAI22_X1 U4501 ( .A1(n4531), .A2(n4415), .B1(n4416), .B2(n4528), .ZN(n3740)
         );
  OAI22_X1 U4502 ( .A1(n4546), .A2(n3738), .B1(STATE_REG_SCAN_IN), .B2(n3737), 
        .ZN(n3739) );
  NOR2_X1 U4503 ( .A1(n3740), .A2(n3739), .ZN(n3741) );
  OAI211_X1 U4504 ( .C1(n4563), .C2(n4274), .A(n3742), .B(n3741), .ZN(U3220)
         );
  NAND2_X1 U4505 ( .A1(n3745), .A2(n3744), .ZN(n3746) );
  XNOR2_X1 U4506 ( .A(n3743), .B(n3746), .ZN(n3753) );
  INV_X1 U4507 ( .A(n4200), .ZN(n3751) );
  AOI22_X1 U4508 ( .A1(n2284), .A2(n4559), .B1(n4194), .B2(n3805), .ZN(n3750)
         );
  OAI22_X1 U4509 ( .A1(n4243), .A2(n4528), .B1(STATE_REG_SCAN_IN), .B2(n3747), 
        .ZN(n3748) );
  INV_X1 U4510 ( .A(n3748), .ZN(n3749) );
  OAI211_X1 U4511 ( .C1(n4563), .C2(n3751), .A(n3750), .B(n3749), .ZN(n3752)
         );
  AOI21_X1 U4512 ( .B1(n3753), .B2(n4554), .A(n3752), .ZN(n3754) );
  INV_X1 U4513 ( .A(n3754), .ZN(U3222) );
  NAND2_X1 U4514 ( .A1(n3757), .A2(n3756), .ZN(n3758) );
  XNOR2_X1 U4515 ( .A(n3755), .B(n3758), .ZN(n3764) );
  NOR2_X1 U4516 ( .A1(STATE_REG_SCAN_IN), .A2(n2708), .ZN(n4635) );
  AOI21_X1 U4517 ( .B1(n4556), .B2(n3986), .A(n4635), .ZN(n3760) );
  NAND2_X1 U4518 ( .A1(n3805), .A2(n3985), .ZN(n3759) );
  OAI211_X1 U4519 ( .C1(n4531), .C2(n4434), .A(n3760), .B(n3759), .ZN(n3761)
         );
  AOI21_X1 U4520 ( .B1(n3811), .B2(n3762), .A(n3761), .ZN(n3763) );
  OAI21_X1 U4521 ( .B1(n3764), .B2(n3813), .A(n3763), .ZN(U3225) );
  NAND2_X1 U4522 ( .A1(n3766), .A2(n3765), .ZN(n3768) );
  XNOR2_X1 U4523 ( .A(n3768), .B(n3767), .ZN(n3772) );
  AOI22_X1 U4524 ( .A1(n4556), .A2(n3984), .B1(REG3_REG_24__SCAN_IN), .B2(
        U3149), .ZN(n3770) );
  AOI22_X1 U4525 ( .A1(n4559), .A2(n4218), .B1(n4178), .B2(n3805), .ZN(n3769)
         );
  OAI211_X1 U4526 ( .C1(n4563), .C2(n4214), .A(n3770), .B(n3769), .ZN(n3771)
         );
  AOI21_X1 U4527 ( .B1(n3772), .B2(n4554), .A(n3771), .ZN(n3773) );
  INV_X1 U4528 ( .A(n3773), .ZN(U3226) );
  NAND2_X1 U4529 ( .A1(n3775), .A2(n3774), .ZN(n3776) );
  XOR2_X1 U4530 ( .A(n3776), .B(n3730), .Z(n3777) );
  NAND2_X1 U4531 ( .A1(n3777), .A2(n4554), .ZN(n3781) );
  OAI22_X1 U4532 ( .A1(n4531), .A2(n4301), .B1(n4294), .B2(n4546), .ZN(n3779)
         );
  OAI22_X1 U4533 ( .A1(n4528), .A2(n4545), .B1(STATE_REG_SCAN_IN), .B2(n4815), 
        .ZN(n3778) );
  NOR2_X1 U4534 ( .A1(n3779), .A2(n3778), .ZN(n3780) );
  OAI211_X1 U4535 ( .C1(n4563), .C2(n4303), .A(n3781), .B(n3780), .ZN(U3230)
         );
  OR2_X1 U4536 ( .A1(n3783), .A2(n3782), .ZN(n3784) );
  AOI21_X1 U4537 ( .B1(n3785), .B2(n3784), .A(n2242), .ZN(n3792) );
  INV_X1 U4538 ( .A(n4261), .ZN(n3790) );
  INV_X1 U4539 ( .A(REG3_REG_22__SCAN_IN), .ZN(n3786) );
  OAI22_X1 U4540 ( .A1(n4528), .A2(n4294), .B1(STATE_REG_SCAN_IN), .B2(n3786), 
        .ZN(n3789) );
  OAI22_X1 U4541 ( .A1(n4531), .A2(n3787), .B1(n4400), .B2(n4546), .ZN(n3788)
         );
  AOI211_X1 U4542 ( .C1(n3811), .C2(n3790), .A(n3789), .B(n3788), .ZN(n3791)
         );
  OAI21_X1 U4543 ( .B1(n3792), .B2(n3813), .A(n3791), .ZN(U3232) );
  NAND2_X1 U4544 ( .A1(n2264), .A2(n3793), .ZN(n3794) );
  INV_X1 U4545 ( .A(n4185), .ZN(n3795) );
  NOR2_X1 U4546 ( .A1(n4563), .A2(n3795), .ZN(n3799) );
  NAND2_X1 U4547 ( .A1(n4177), .A2(n3805), .ZN(n3797) );
  AOI22_X1 U4548 ( .A1(n4178), .A2(n4556), .B1(REG3_REG_26__SCAN_IN), .B2(
        U3149), .ZN(n3796) );
  OAI211_X1 U4549 ( .C1(n4531), .C2(n4183), .A(n3797), .B(n3796), .ZN(n3798)
         );
  INV_X1 U4550 ( .A(n3801), .ZN(U3237) );
  NAND2_X1 U4551 ( .A1(n3802), .A2(n3803), .ZN(n3804) );
  XOR2_X1 U4552 ( .A(n4536), .B(n3804), .Z(n3814) );
  AND2_X1 U4553 ( .A1(U3149), .A2(REG3_REG_15__SCAN_IN), .ZN(n4615) );
  AOI21_X1 U4554 ( .B1(n3805), .B2(n3986), .A(n4615), .ZN(n3807) );
  NAND2_X1 U4555 ( .A1(n4556), .A2(n3988), .ZN(n3806) );
  OAI211_X1 U4556 ( .C1(n4531), .C2(n3808), .A(n3807), .B(n3806), .ZN(n3809)
         );
  AOI21_X1 U4557 ( .B1(n3811), .B2(n3810), .A(n3809), .ZN(n3812) );
  OAI21_X1 U4558 ( .B1(n3814), .B2(n3813), .A(n3812), .ZN(U3238) );
  INV_X1 U4559 ( .A(n3880), .ZN(n3815) );
  NOR2_X1 U4560 ( .A1(n3892), .A2(n3815), .ZN(n3956) );
  INV_X1 U4561 ( .A(n3956), .ZN(n3830) );
  NAND2_X1 U4562 ( .A1(n3816), .A2(n3819), .ZN(n3938) );
  NAND2_X1 U4563 ( .A1(n3818), .A2(n3817), .ZN(n3928) );
  NAND2_X1 U4564 ( .A1(n3928), .A2(n3819), .ZN(n3937) );
  OAI21_X1 U4565 ( .B1(n3820), .B2(n3938), .A(n3937), .ZN(n3822) );
  INV_X1 U4566 ( .A(n3821), .ZN(n3940) );
  AOI21_X1 U4567 ( .B1(n3822), .B2(n3943), .A(n3940), .ZN(n3825) );
  INV_X1 U4568 ( .A(n4234), .ZN(n3824) );
  OAI21_X1 U4569 ( .B1(n3825), .B2(n3824), .A(n3823), .ZN(n3826) );
  INV_X1 U4570 ( .A(n3826), .ZN(n3828) );
  OAI21_X1 U4571 ( .B1(n3828), .B2(n3950), .A(n3827), .ZN(n3829) );
  OAI221_X1 U4572 ( .B1(n3830), .B2(n3952), .C1(n3830), .C2(n3829), .A(n3961), 
        .ZN(n3834) );
  NAND2_X1 U4573 ( .A1(n2235), .A2(DATAI_30_), .ZN(n4121) );
  INV_X1 U4574 ( .A(REG2_REG_31__SCAN_IN), .ZN(n4126) );
  NAND2_X1 U4575 ( .A1(n2537), .A2(REG1_REG_31__SCAN_IN), .ZN(n3832) );
  NAND2_X1 U4576 ( .A1(n2538), .A2(REG0_REG_31__SCAN_IN), .ZN(n3831) );
  OAI211_X1 U4577 ( .C1(n2562), .C2(n4126), .A(n3832), .B(n3831), .ZN(n4124)
         );
  NAND2_X1 U4578 ( .A1(n2235), .A2(DATAI_31_), .ZN(n4125) );
  NAND2_X1 U4579 ( .A1(n4124), .A2(n4125), .ZN(n3851) );
  OAI21_X1 U4580 ( .B1(n3980), .B2(n4121), .A(n3851), .ZN(n3865) );
  AOI21_X1 U4581 ( .B1(n3837), .B2(n4133), .A(n3865), .ZN(n3840) );
  INV_X1 U4582 ( .A(n3840), .ZN(n3833) );
  NOR4_X1 U4583 ( .A1(n3834), .A2(n3839), .A3(n3838), .A4(n3833), .ZN(n3844)
         );
  INV_X1 U4584 ( .A(n3835), .ZN(n3836) );
  OAI21_X1 U4585 ( .B1(n3837), .B2(n4133), .A(n3836), .ZN(n3841) );
  NOR2_X1 U4586 ( .A1(n3852), .A2(n3841), .ZN(n3957) );
  NOR2_X1 U4587 ( .A1(n3839), .A2(n3838), .ZN(n3842) );
  OAI21_X1 U4588 ( .B1(n3842), .B2(n3841), .A(n3840), .ZN(n3848) );
  AOI21_X1 U4589 ( .B1(n4154), .B2(n3957), .A(n3848), .ZN(n3843) );
  OAI22_X1 U4590 ( .A1(n3844), .A2(n3843), .B1(n4124), .B2(n4121), .ZN(n3971)
         );
  NAND2_X1 U4591 ( .A1(n3980), .A2(n4121), .ZN(n3847) );
  AOI21_X1 U4592 ( .B1(n3847), .B2(n4124), .A(n4125), .ZN(n3846) );
  NOR2_X1 U4593 ( .A1(n3846), .A2(n3845), .ZN(n3970) );
  OAI21_X1 U4594 ( .B1(n4124), .B2(n4125), .A(n3847), .ZN(n3966) );
  INV_X1 U4595 ( .A(n3848), .ZN(n3849) );
  AOI211_X1 U4596 ( .C1(n3851), .C2(n3966), .A(n3850), .B(n3849), .ZN(n3969)
         );
  XNOR2_X1 U4597 ( .A(n3984), .B(n4225), .ZN(n4227) );
  INV_X1 U4598 ( .A(n4227), .ZN(n4238) );
  NAND2_X1 U4599 ( .A1(n2319), .A2(n3853), .ZN(n4174) );
  INV_X1 U4600 ( .A(n4337), .ZN(n3855) );
  NAND4_X1 U4601 ( .A1(n3855), .A2(n3854), .A3(n2261), .A4(n4356), .ZN(n3861)
         );
  NAND4_X1 U4602 ( .A1(n3859), .A2(n3858), .A3(n3857), .A4(n3856), .ZN(n3860)
         );
  NOR2_X1 U4603 ( .A1(n3861), .A2(n3860), .ZN(n3878) );
  INV_X1 U4604 ( .A(n3862), .ZN(n3863) );
  OR2_X1 U4605 ( .A1(n3864), .A2(n3863), .ZN(n4288) );
  INV_X1 U4606 ( .A(n3865), .ZN(n3868) );
  NAND4_X1 U4607 ( .A1(n4288), .A2(n3868), .A3(n3867), .A4(n3866), .ZN(n3874)
         );
  NAND4_X1 U4608 ( .A1(n3872), .A2(n3871), .A3(n3870), .A4(n3869), .ZN(n3873)
         );
  NOR2_X1 U4609 ( .A1(n3874), .A2(n3873), .ZN(n3877) );
  XNOR2_X1 U4610 ( .A(n4545), .B(n3875), .ZN(n4310) );
  INV_X1 U4611 ( .A(n4310), .ZN(n4318) );
  NAND4_X1 U4612 ( .A1(n3878), .A2(n3877), .A3(n4318), .A4(n3876), .ZN(n3879)
         );
  NOR2_X1 U4613 ( .A1(n4174), .A2(n3879), .ZN(n3891) );
  NAND2_X1 U4614 ( .A1(n3881), .A2(n3880), .ZN(n4208) );
  INV_X1 U4615 ( .A(n3948), .ZN(n3882) );
  INV_X1 U4616 ( .A(n3883), .ZN(n3885) );
  AND4_X1 U4617 ( .A1(n3887), .A2(n3886), .A3(n3885), .A4(n3884), .ZN(n3888)
         );
  NAND4_X1 U4618 ( .A1(n4255), .A2(n4270), .A3(n3888), .A4(n4675), .ZN(n3889)
         );
  NOR2_X1 U4619 ( .A1(n4208), .A2(n3889), .ZN(n3890) );
  AND4_X1 U4620 ( .A1(n4154), .A2(n4238), .A3(n3891), .A4(n3890), .ZN(n3897)
         );
  INV_X1 U4621 ( .A(n3892), .ZN(n3893) );
  NAND2_X1 U4622 ( .A1(n3893), .A2(n4172), .ZN(n4192) );
  INV_X1 U4623 ( .A(n4192), .ZN(n3894) );
  NAND4_X1 U4624 ( .A1(n3897), .A2(n3896), .A3(n3895), .A4(n3894), .ZN(n3965)
         );
  OAI211_X1 U4625 ( .C1(n2286), .C2(n4518), .A(n3900), .B(n3899), .ZN(n3903)
         );
  NAND3_X1 U4626 ( .A1(n3903), .A2(n3902), .A3(n3901), .ZN(n3906) );
  NAND3_X1 U4627 ( .A1(n3906), .A2(n3905), .A3(n3904), .ZN(n3909) );
  NAND3_X1 U4628 ( .A1(n3909), .A2(n3908), .A3(n3907), .ZN(n3912) );
  NAND4_X1 U4629 ( .A1(n3912), .A2(n3911), .A3(n3910), .A4(n3921), .ZN(n3914)
         );
  NAND3_X1 U4630 ( .A1(n3914), .A2(n2261), .A3(n3913), .ZN(n3920) );
  AND2_X1 U4631 ( .A1(n3916), .A2(n3915), .ZN(n3922) );
  INV_X1 U4632 ( .A(n3917), .ZN(n3919) );
  AOI211_X1 U4633 ( .C1(n3920), .C2(n3922), .A(n3919), .B(n2301), .ZN(n3929)
         );
  INV_X1 U4634 ( .A(n3922), .ZN(n3924) );
  NOR3_X1 U4635 ( .A1(n2303), .A2(n3924), .A3(n3923), .ZN(n3926) );
  INV_X1 U4636 ( .A(n3931), .ZN(n3925) );
  OAI21_X1 U4637 ( .B1(n3926), .B2(n3925), .A(n3937), .ZN(n3927) );
  OAI21_X1 U4638 ( .B1(n3929), .B2(n3928), .A(n3927), .ZN(n3935) );
  NAND2_X1 U4639 ( .A1(n3931), .A2(n3930), .ZN(n3932) );
  NAND4_X1 U4640 ( .A1(n3935), .A2(n3934), .A3(n3933), .A4(n3932), .ZN(n3942)
         );
  INV_X1 U4641 ( .A(n3936), .ZN(n3939) );
  OAI21_X1 U4642 ( .B1(n3939), .B2(n3938), .A(n3937), .ZN(n3941) );
  AOI21_X1 U4643 ( .B1(n3942), .B2(n3941), .A(n3940), .ZN(n3947) );
  INV_X1 U4644 ( .A(n3943), .ZN(n3946) );
  INV_X1 U4645 ( .A(n3944), .ZN(n3945) );
  OAI21_X1 U4646 ( .B1(n3947), .B2(n3946), .A(n3945), .ZN(n3949) );
  AOI211_X1 U4647 ( .C1(n3949), .C2(n4234), .A(n3948), .B(n4233), .ZN(n3951)
         );
  NOR2_X1 U4648 ( .A1(n3951), .A2(n3950), .ZN(n3954) );
  OAI21_X1 U4649 ( .B1(n3954), .B2(n3953), .A(n3952), .ZN(n3955) );
  NAND2_X1 U4650 ( .A1(n3956), .A2(n3955), .ZN(n3960) );
  INV_X1 U4651 ( .A(n3957), .ZN(n3958) );
  AOI211_X1 U4652 ( .C1(n3961), .C2(n3960), .A(n3959), .B(n3958), .ZN(n3962)
         );
  INV_X1 U4653 ( .A(n3962), .ZN(n3964) );
  MUX2_X1 U4654 ( .A(n3965), .B(n3964), .S(n3963), .Z(n3967) );
  NOR2_X1 U4655 ( .A1(n3967), .A2(n3966), .ZN(n3968) );
  AOI211_X1 U4656 ( .C1(n3971), .C2(n3970), .A(n3969), .B(n3968), .ZN(n3972)
         );
  XNOR2_X1 U4657 ( .A(n3972), .B(n4116), .ZN(n3979) );
  NAND2_X1 U4658 ( .A1(n3974), .A2(n3973), .ZN(n3975) );
  OAI211_X1 U4659 ( .C1(n3976), .C2(n3978), .A(n3975), .B(B_REG_SCAN_IN), .ZN(
        n3977) );
  OAI21_X1 U4660 ( .B1(n3979), .B2(n3978), .A(n3977), .ZN(U3239) );
  MUX2_X1 U4661 ( .A(DATAO_REG_31__SCAN_IN), .B(n4124), .S(U4043), .Z(U3581)
         );
  MUX2_X1 U4662 ( .A(DATAO_REG_30__SCAN_IN), .B(n3980), .S(U4043), .Z(U3580)
         );
  MUX2_X1 U4663 ( .A(DATAO_REG_29__SCAN_IN), .B(n3981), .S(U4043), .Z(U3579)
         );
  MUX2_X1 U4664 ( .A(DATAO_REG_28__SCAN_IN), .B(n4157), .S(U4043), .Z(U3578)
         );
  MUX2_X1 U4665 ( .A(DATAO_REG_27__SCAN_IN), .B(n4177), .S(U4043), .Z(U3577)
         );
  MUX2_X1 U4666 ( .A(DATAO_REG_26__SCAN_IN), .B(n4194), .S(U4043), .Z(U3576)
         );
  MUX2_X1 U4667 ( .A(DATAO_REG_25__SCAN_IN), .B(n4178), .S(U4043), .Z(U3575)
         );
  MUX2_X1 U4668 ( .A(DATAO_REG_24__SCAN_IN), .B(n3983), .S(n3996), .Z(U3574)
         );
  MUX2_X1 U4669 ( .A(DATAO_REG_23__SCAN_IN), .B(n3984), .S(U4043), .Z(U3573)
         );
  MUX2_X1 U4670 ( .A(DATAO_REG_22__SCAN_IN), .B(n4268), .S(n3996), .Z(U3572)
         );
  MUX2_X1 U4671 ( .A(DATAO_REG_21__SCAN_IN), .B(n4258), .S(U4043), .Z(U3571)
         );
  MUX2_X1 U4672 ( .A(DATAO_REG_20__SCAN_IN), .B(n4322), .S(n3996), .Z(U3570)
         );
  MUX2_X1 U4673 ( .A(DATAO_REG_19__SCAN_IN), .B(n4339), .S(n3996), .Z(U3569)
         );
  MUX2_X1 U4674 ( .A(DATAO_REG_18__SCAN_IN), .B(n3985), .S(n3996), .Z(U3568)
         );
  MUX2_X1 U4675 ( .A(DATAO_REG_17__SCAN_IN), .B(n4557), .S(n3996), .Z(U3567)
         );
  MUX2_X1 U4676 ( .A(DATAO_REG_16__SCAN_IN), .B(n3986), .S(n3996), .Z(U3566)
         );
  MUX2_X1 U4677 ( .A(DATAO_REG_15__SCAN_IN), .B(n3987), .S(n3996), .Z(U3565)
         );
  MUX2_X1 U4678 ( .A(DATAO_REG_14__SCAN_IN), .B(n3988), .S(n3996), .Z(U3564)
         );
  MUX2_X1 U4679 ( .A(DATAO_REG_13__SCAN_IN), .B(n3989), .S(n3996), .Z(U3563)
         );
  MUX2_X1 U4680 ( .A(DATAO_REG_12__SCAN_IN), .B(n3990), .S(n3996), .Z(U3562)
         );
  MUX2_X1 U4681 ( .A(DATAO_REG_11__SCAN_IN), .B(n3991), .S(n3996), .Z(U3561)
         );
  MUX2_X1 U4682 ( .A(DATAO_REG_10__SCAN_IN), .B(n3992), .S(n3996), .Z(U3560)
         );
  MUX2_X1 U4683 ( .A(DATAO_REG_9__SCAN_IN), .B(n3993), .S(n3996), .Z(U3559) );
  MUX2_X1 U4684 ( .A(DATAO_REG_8__SCAN_IN), .B(n3994), .S(n3996), .Z(U3558) );
  MUX2_X1 U4685 ( .A(DATAO_REG_7__SCAN_IN), .B(n3995), .S(n3996), .Z(U3557) );
  MUX2_X1 U4686 ( .A(DATAO_REG_6__SCAN_IN), .B(n3997), .S(n3996), .Z(U3556) );
  MUX2_X1 U4687 ( .A(DATAO_REG_5__SCAN_IN), .B(n3998), .S(U4043), .Z(U3555) );
  MUX2_X1 U4688 ( .A(DATAO_REG_4__SCAN_IN), .B(n3999), .S(U4043), .Z(U3554) );
  MUX2_X1 U4689 ( .A(DATAO_REG_3__SCAN_IN), .B(n4363), .S(U4043), .Z(U3553) );
  MUX2_X1 U4690 ( .A(DATAO_REG_2__SCAN_IN), .B(n4000), .S(U4043), .Z(U3552) );
  MUX2_X1 U4691 ( .A(DATAO_REG_1__SCAN_IN), .B(n2543), .S(U4043), .Z(U3551) );
  MUX2_X1 U4692 ( .A(DATAO_REG_0__SCAN_IN), .B(n2933), .S(U4043), .Z(U3550) );
  NAND3_X1 U4693 ( .A1(n4637), .A2(IR_REG_0__SCAN_IN), .A3(n2935), .ZN(n4009)
         );
  AOI21_X1 U4694 ( .B1(n2935), .B2(n4001), .A(n4004), .ZN(n4003) );
  MUX2_X1 U4695 ( .A(n4004), .B(n4003), .S(n4002), .Z(n4005) );
  AOI22_X1 U4696 ( .A1(n4006), .A2(n4005), .B1(REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n4008) );
  NAND2_X1 U4697 ( .A1(n4636), .A2(ADDR_REG_0__SCAN_IN), .ZN(n4007) );
  NAND3_X1 U4698 ( .A1(n4009), .A2(n4008), .A3(n4007), .ZN(U3240) );
  OAI211_X1 U4699 ( .C1(n4011), .C2(n4010), .A(n4593), .B(n4025), .ZN(n4017)
         );
  OAI211_X1 U4700 ( .C1(n4014), .C2(n4013), .A(n4637), .B(n4012), .ZN(n4016)
         );
  AOI22_X1 U4701 ( .A1(n4636), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n4015) );
  NAND4_X1 U4702 ( .A1(n4018), .A2(n4017), .A3(n4016), .A4(n4015), .ZN(U3241)
         );
  AOI22_X1 U4703 ( .A1(n4636), .A2(ADDR_REG_2__SCAN_IN), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n4034) );
  OAI211_X1 U4704 ( .C1(n4021), .C2(n4020), .A(n4637), .B(n4019), .ZN(n4030)
         );
  MUX2_X1 U4705 ( .A(n4023), .B(REG2_REG_2__SCAN_IN), .S(n4022), .Z(n4026) );
  NAND3_X1 U4706 ( .A1(n4026), .A2(n4025), .A3(n4024), .ZN(n4027) );
  NAND3_X1 U4707 ( .A1(n4593), .A2(n4028), .A3(n4027), .ZN(n4029) );
  AND2_X1 U4708 ( .A1(n4030), .A2(n4029), .ZN(n4033) );
  OR2_X1 U4709 ( .A1(n4642), .A2(n4031), .ZN(n4032) );
  NAND4_X1 U4710 ( .A1(n4035), .A2(n4034), .A3(n4033), .A4(n4032), .ZN(U3242)
         );
  INV_X1 U4711 ( .A(REG1_REG_11__SCAN_IN), .ZN(n4714) );
  INV_X1 U4712 ( .A(n4522), .ZN(n4598) );
  NAND2_X1 U4713 ( .A1(n4567), .A2(REG1_REG_9__SCAN_IN), .ZN(n4040) );
  INV_X1 U4714 ( .A(REG1_REG_9__SCAN_IN), .ZN(n4038) );
  MUX2_X1 U4715 ( .A(n4038), .B(REG1_REG_9__SCAN_IN), .S(n4567), .Z(n4039) );
  INV_X1 U4716 ( .A(n4039), .ZN(n4569) );
  NAND2_X1 U4717 ( .A1(n4570), .A2(n4569), .ZN(n4568) );
  NAND2_X1 U4718 ( .A1(n4040), .A2(n4568), .ZN(n4041) );
  NAND2_X1 U4719 ( .A1(n4049), .A2(n4041), .ZN(n4042) );
  INV_X1 U4720 ( .A(n4049), .ZN(n4672) );
  XNOR2_X1 U4721 ( .A(n4041), .B(n4672), .ZN(n4586) );
  NAND2_X1 U4722 ( .A1(REG1_REG_10__SCAN_IN), .A2(n4586), .ZN(n4585) );
  NAND2_X1 U4723 ( .A1(n4042), .A2(n4585), .ZN(n4591) );
  MUX2_X1 U4724 ( .A(REG1_REG_11__SCAN_IN), .B(n4714), .S(n4522), .Z(n4590) );
  NAND2_X1 U4725 ( .A1(n4591), .A2(n4590), .ZN(n4589) );
  OAI211_X1 U4726 ( .C1(n4044), .C2(REG1_REG_12__SCAN_IN), .A(n4637), .B(n4065), .ZN(n4057) );
  AOI22_X1 U4727 ( .A1(n4045), .A2(n4064), .B1(n4636), .B2(
        ADDR_REG_12__SCAN_IN), .ZN(n4056) );
  MUX2_X1 U4728 ( .A(REG2_REG_11__SCAN_IN), .B(n3395), .S(n4522), .Z(n4594) );
  NAND2_X1 U4729 ( .A1(n4567), .A2(REG2_REG_9__SCAN_IN), .ZN(n4048) );
  MUX2_X1 U4730 ( .A(REG2_REG_9__SCAN_IN), .B(n3344), .S(n4567), .Z(n4572) );
  INV_X1 U4731 ( .A(REG2_REG_8__SCAN_IN), .ZN(n4653) );
  NAND2_X1 U4732 ( .A1(n4572), .A2(n4573), .ZN(n4571) );
  NAND2_X1 U4733 ( .A1(n4048), .A2(n4571), .ZN(n4050) );
  NAND2_X1 U4734 ( .A1(n4049), .A2(n4050), .ZN(n4051) );
  XNOR2_X1 U4735 ( .A(n4050), .B(n4672), .ZN(n4581) );
  NAND2_X1 U4736 ( .A1(REG2_REG_10__SCAN_IN), .A2(n4581), .ZN(n4580) );
  NAND2_X1 U4737 ( .A1(n4051), .A2(n4580), .ZN(n4595) );
  NAND2_X1 U4738 ( .A1(n4594), .A2(n4595), .ZN(n4592) );
  OAI211_X1 U4739 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4052), .A(n4593), .B(n4059), .ZN(n4054) );
  AND2_X1 U4740 ( .A1(n4054), .A2(n4053), .ZN(n4055) );
  NAND3_X1 U4741 ( .A1(n4057), .A2(n4056), .A3(n4055), .ZN(U3252) );
  INV_X1 U4742 ( .A(REG2_REG_13__SCAN_IN), .ZN(n4058) );
  NOR2_X1 U4743 ( .A1(n4073), .A2(n4058), .ZN(n4090) );
  AOI21_X1 U4744 ( .B1(n4058), .B2(n4073), .A(n4090), .ZN(n4062) );
  OAI21_X1 U4745 ( .B1(n4043), .B2(n4060), .A(n4059), .ZN(n4091) );
  OAI21_X1 U4746 ( .B1(n4062), .B2(n4091), .A(n4593), .ZN(n4061) );
  AOI21_X1 U4747 ( .B1(n4062), .B2(n4091), .A(n4061), .ZN(n4075) );
  NAND2_X1 U4748 ( .A1(n4064), .A2(n4063), .ZN(n4066) );
  NAND2_X1 U4749 ( .A1(n4521), .A2(REG1_REG_13__SCAN_IN), .ZN(n4077) );
  INV_X1 U4750 ( .A(n4077), .ZN(n4067) );
  AOI21_X1 U4751 ( .B1(n4456), .B2(n4073), .A(n4067), .ZN(n4068) );
  NAND2_X1 U4752 ( .A1(n4068), .A2(n4069), .ZN(n4076) );
  OAI211_X1 U4753 ( .C1(n4069), .C2(n4068), .A(n4637), .B(n4076), .ZN(n4072)
         );
  AOI21_X1 U4754 ( .B1(n4636), .B2(ADDR_REG_13__SCAN_IN), .A(n4070), .ZN(n4071) );
  OAI211_X1 U4755 ( .C1(n4642), .C2(n4073), .A(n4072), .B(n4071), .ZN(n4074)
         );
  OR2_X1 U4756 ( .A1(n4075), .A2(n4074), .ZN(U3253) );
  XOR2_X1 U4757 ( .A(REG1_REG_18__SCAN_IN), .B(n4520), .Z(n4110) );
  NOR2_X1 U4758 ( .A1(n4099), .A2(REG1_REG_17__SCAN_IN), .ZN(n4084) );
  NAND2_X1 U4759 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4096), .ZN(n4080) );
  INV_X1 U4760 ( .A(n4096), .ZN(n4670) );
  AOI22_X1 U4761 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4096), .B1(n4670), .B2(
        n3517), .ZN(n4618) );
  NAND2_X1 U4762 ( .A1(n4077), .A2(n4076), .ZN(n4078) );
  NAND2_X1 U4763 ( .A1(n4093), .A2(n4078), .ZN(n4079) );
  INV_X1 U4764 ( .A(n4093), .ZN(n4671) );
  XNOR2_X1 U4765 ( .A(n4078), .B(n4671), .ZN(n4608) );
  NAND2_X1 U4766 ( .A1(REG1_REG_14__SCAN_IN), .A2(n4608), .ZN(n4607) );
  NAND2_X1 U4767 ( .A1(n4079), .A2(n4607), .ZN(n4617) );
  NAND2_X1 U4768 ( .A1(n4618), .A2(n4617), .ZN(n4616) );
  NOR2_X1 U4769 ( .A1(n4668), .A2(n4081), .ZN(n4082) );
  INV_X1 U4770 ( .A(n4668), .ZN(n4629) );
  INV_X1 U4771 ( .A(REG1_REG_17__SCAN_IN), .ZN(n4083) );
  AOI22_X1 U4772 ( .A1(n4099), .A2(n4083), .B1(REG1_REG_17__SCAN_IN), .B2(
        n4667), .ZN(n4638) );
  XOR2_X1 U4773 ( .A(n4110), .B(n4111), .Z(n4104) );
  INV_X1 U4774 ( .A(n4520), .ZN(n4087) );
  INV_X1 U4775 ( .A(REG3_REG_18__SCAN_IN), .ZN(n4544) );
  NOR2_X1 U4776 ( .A1(STATE_REG_SCAN_IN), .A2(n4544), .ZN(n4085) );
  AOI21_X1 U4777 ( .B1(n4636), .B2(ADDR_REG_18__SCAN_IN), .A(n4085), .ZN(n4086) );
  OAI21_X1 U4778 ( .B1(n4642), .B2(n4087), .A(n4086), .ZN(n4103) );
  NOR2_X1 U4779 ( .A1(n4520), .A2(n4348), .ZN(n4088) );
  AOI21_X1 U4780 ( .B1(n4520), .B2(n4348), .A(n4088), .ZN(n4101) );
  NOR2_X1 U4781 ( .A1(n4099), .A2(REG2_REG_17__SCAN_IN), .ZN(n4089) );
  AOI21_X1 U4782 ( .B1(REG2_REG_17__SCAN_IN), .B2(n4099), .A(n4089), .ZN(n4633) );
  NOR2_X1 U4783 ( .A1(n4671), .A2(n4092), .ZN(n4094) );
  XOR2_X1 U4784 ( .A(n4093), .B(n4092), .Z(n4604) );
  NAND2_X1 U4785 ( .A1(REG2_REG_15__SCAN_IN), .A2(n4096), .ZN(n4095) );
  OAI21_X1 U4786 ( .B1(REG2_REG_15__SCAN_IN), .B2(n4096), .A(n4095), .ZN(n4612) );
  NAND2_X1 U4787 ( .A1(n4097), .A2(n4629), .ZN(n4098) );
  XNOR2_X1 U4788 ( .A(n4097), .B(n4668), .ZN(n4622) );
  NAND2_X1 U4789 ( .A1(n4622), .A2(n3506), .ZN(n4621) );
  NAND2_X1 U4790 ( .A1(n4098), .A2(n4621), .ZN(n4631) );
  AOI211_X1 U4791 ( .C1(n4104), .C2(n4637), .A(n4103), .B(n4102), .ZN(n4105)
         );
  INV_X1 U4792 ( .A(n4105), .ZN(U3258) );
  INV_X1 U4793 ( .A(REG2_REG_19__SCAN_IN), .ZN(n4106) );
  MUX2_X1 U4794 ( .A(REG2_REG_19__SCAN_IN), .B(n4106), .S(n4519), .Z(n4108) );
  XOR2_X1 U4795 ( .A(n4108), .B(n4107), .Z(n4120) );
  INV_X1 U4796 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4109) );
  MUX2_X1 U4797 ( .A(n4109), .B(REG1_REG_19__SCAN_IN), .S(n4519), .Z(n4113) );
  AOI22_X1 U4798 ( .A1(n4111), .A2(n4110), .B1(REG1_REG_18__SCAN_IN), .B2(
        n4520), .ZN(n4112) );
  XOR2_X1 U4799 ( .A(n4113), .B(n4112), .Z(n4118) );
  NAND2_X1 U4800 ( .A1(n4636), .A2(ADDR_REG_19__SCAN_IN), .ZN(n4114) );
  OAI211_X1 U4801 ( .C1(n4642), .C2(n4116), .A(n4115), .B(n4114), .ZN(n4117)
         );
  AOI21_X1 U4802 ( .B1(n4118), .B2(n4637), .A(n4117), .ZN(n4119) );
  OAI21_X1 U4803 ( .B1(n4120), .B2(n4630), .A(n4119), .ZN(U3259) );
  XNOR2_X1 U4804 ( .A(n4376), .B(n4125), .ZN(n4462) );
  INV_X1 U4805 ( .A(n4122), .ZN(n4123) );
  NAND2_X1 U4806 ( .A1(n4124), .A2(n4123), .ZN(n4378) );
  OAI21_X1 U4807 ( .B1(n4125), .B2(n4433), .A(n4378), .ZN(n4459) );
  NOR2_X1 U4808 ( .A1(n4654), .A2(n4126), .ZN(n4127) );
  AOI21_X1 U4809 ( .B1(n4654), .B2(n4459), .A(n4127), .ZN(n4128) );
  OAI21_X1 U4810 ( .B1(n4462), .B2(n4328), .A(n4128), .ZN(U3260) );
  INV_X1 U4811 ( .A(n4129), .ZN(n4140) );
  OAI22_X1 U4812 ( .A1(n4131), .A2(n4277), .B1(n4654), .B2(n4130), .ZN(n4132)
         );
  AOI21_X1 U4813 ( .B1(n4133), .B2(n4282), .A(n4132), .ZN(n4139) );
  OAI22_X1 U4814 ( .A1(n4135), .A2(n4328), .B1(n4134), .B2(n4651), .ZN(n4136)
         );
  OAI21_X1 U4815 ( .B1(n4137), .B2(n4136), .A(n4654), .ZN(n4138) );
  OAI211_X1 U4816 ( .C1(n4140), .C2(n4353), .A(n4139), .B(n4138), .ZN(U3354)
         );
  INV_X1 U4817 ( .A(n4141), .ZN(n4150) );
  AOI22_X1 U4818 ( .A1(n4142), .A2(n4643), .B1(REG2_REG_28__SCAN_IN), .B2(
        n4663), .ZN(n4145) );
  NAND2_X1 U4819 ( .A1(n4282), .A2(n4143), .ZN(n4144) );
  OAI211_X1 U4820 ( .C1(n4146), .C2(n4277), .A(n4145), .B(n4144), .ZN(n4149)
         );
  NOR2_X1 U4821 ( .A1(n4147), .A2(n4663), .ZN(n4148) );
  AOI211_X1 U4822 ( .C1(n4657), .C2(n4150), .A(n4149), .B(n4148), .ZN(n4151)
         );
  OAI21_X1 U4823 ( .B1(n4152), .B2(n4353), .A(n4151), .ZN(U3262) );
  XNOR2_X1 U4824 ( .A(n4153), .B(n4154), .ZN(n4388) );
  INV_X1 U4825 ( .A(n4388), .ZN(n4170) );
  XNOR2_X1 U4826 ( .A(n4155), .B(n4154), .ZN(n4156) );
  NAND2_X1 U4827 ( .A1(n4156), .A2(n4342), .ZN(n4159) );
  NAND2_X1 U4828 ( .A1(n4157), .A2(n4362), .ZN(n4158) );
  NAND2_X1 U4829 ( .A1(n4159), .A2(n4158), .ZN(n4387) );
  INV_X1 U4830 ( .A(n4182), .ZN(n4162) );
  INV_X1 U4831 ( .A(n4160), .ZN(n4161) );
  OAI21_X1 U4832 ( .B1(n4162), .B2(n4384), .A(n4161), .ZN(n4469) );
  AOI22_X1 U4833 ( .A1(n4163), .A2(n4643), .B1(REG2_REG_27__SCAN_IN), .B2(
        n4663), .ZN(n4164) );
  OAI21_X1 U4834 ( .B1(n4385), .B2(n4277), .A(n4164), .ZN(n4165) );
  AOI21_X1 U4835 ( .B1(n4166), .B2(n4282), .A(n4165), .ZN(n4167) );
  OAI21_X1 U4836 ( .B1(n4469), .B2(n4328), .A(n4167), .ZN(n4168) );
  AOI21_X1 U4837 ( .B1(n4387), .B2(n4654), .A(n4168), .ZN(n4169) );
  OAI21_X1 U4838 ( .B1(n4170), .B2(n4353), .A(n4169), .ZN(U3263) );
  XNOR2_X1 U4839 ( .A(n4171), .B(n4174), .ZN(n4392) );
  INV_X1 U4840 ( .A(n4392), .ZN(n4189) );
  NAND2_X1 U4841 ( .A1(n4173), .A2(n4172), .ZN(n4175) );
  XNOR2_X1 U4842 ( .A(n4175), .B(n4174), .ZN(n4181) );
  AOI22_X1 U4843 ( .A1(n4177), .A2(n4362), .B1(n4380), .B2(n4176), .ZN(n4180)
         );
  NAND2_X1 U4844 ( .A1(n4178), .A2(n4291), .ZN(n4179) );
  OAI211_X1 U4845 ( .C1(n4181), .C2(n4366), .A(n4180), .B(n4179), .ZN(n4391)
         );
  INV_X1 U4846 ( .A(n4199), .ZN(n4184) );
  OAI21_X1 U4847 ( .B1(n4184), .B2(n4183), .A(n4182), .ZN(n4473) );
  AOI22_X1 U4848 ( .A1(n4663), .A2(REG2_REG_26__SCAN_IN), .B1(n4185), .B2(
        n4643), .ZN(n4186) );
  OAI21_X1 U4849 ( .B1(n4473), .B2(n4328), .A(n4186), .ZN(n4187) );
  AOI21_X1 U4850 ( .B1(n4391), .B2(n4654), .A(n4187), .ZN(n4188) );
  OAI21_X1 U4851 ( .B1(n4189), .B2(n4353), .A(n4188), .ZN(U3264) );
  XOR2_X1 U4852 ( .A(n4192), .B(n4190), .Z(n4396) );
  INV_X1 U4853 ( .A(n4396), .ZN(n4204) );
  XOR2_X1 U4854 ( .A(n4192), .B(n4191), .Z(n4196) );
  OAI22_X1 U4855 ( .A1(n4243), .A2(n4435), .B1(n4197), .B2(n4433), .ZN(n4193)
         );
  AOI21_X1 U4856 ( .B1(n4362), .B2(n4194), .A(n4193), .ZN(n4195) );
  OAI21_X1 U4857 ( .B1(n4196), .B2(n4366), .A(n4195), .ZN(n4395) );
  OR2_X1 U4858 ( .A1(n4212), .A2(n4197), .ZN(n4198) );
  NAND2_X1 U4859 ( .A1(n4199), .A2(n4198), .ZN(n4477) );
  AOI22_X1 U4860 ( .A1(n4663), .A2(REG2_REG_25__SCAN_IN), .B1(n4200), .B2(
        n4643), .ZN(n4201) );
  OAI21_X1 U4861 ( .B1(n4477), .B2(n4328), .A(n4201), .ZN(n4202) );
  AOI21_X1 U4862 ( .B1(n4395), .B2(n4654), .A(n4202), .ZN(n4203) );
  OAI21_X1 U4863 ( .B1(n4204), .B2(n4353), .A(n4203), .ZN(U3265) );
  XOR2_X1 U4864 ( .A(n4208), .B(n4205), .Z(n4403) );
  INV_X1 U4865 ( .A(n4403), .ZN(n4222) );
  NAND2_X1 U4866 ( .A1(n4207), .A2(n4206), .ZN(n4209) );
  XNOR2_X1 U4867 ( .A(n4209), .B(n4208), .ZN(n4211) );
  OAI22_X1 U4868 ( .A1(n4211), .A2(n4366), .B1(n4210), .B2(n4293), .ZN(n4402)
         );
  INV_X1 U4869 ( .A(n4212), .ZN(n4213) );
  OAI21_X1 U4870 ( .B1(n4223), .B2(n4399), .A(n4213), .ZN(n4481) );
  OAI22_X1 U4871 ( .A1(n4654), .A2(n4215), .B1(n4214), .B2(n4651), .ZN(n4217)
         );
  NOR2_X1 U4872 ( .A1(n4277), .A2(n4400), .ZN(n4216) );
  AOI211_X1 U4873 ( .C1(n4282), .C2(n4218), .A(n4217), .B(n4216), .ZN(n4219)
         );
  OAI21_X1 U4874 ( .B1(n4481), .B2(n4328), .A(n4219), .ZN(n4220) );
  AOI21_X1 U4875 ( .B1(n4402), .B2(n4654), .A(n4220), .ZN(n4221) );
  OAI21_X1 U4876 ( .B1(n4222), .B2(n4353), .A(n4221), .ZN(U3266) );
  INV_X1 U4877 ( .A(n4250), .ZN(n4226) );
  INV_X1 U4878 ( .A(n4223), .ZN(n4224) );
  OAI21_X1 U4879 ( .B1(n4226), .B2(n4225), .A(n4224), .ZN(n4485) );
  XNOR2_X1 U4880 ( .A(n4228), .B(n4227), .ZN(n4407) );
  NAND2_X1 U4881 ( .A1(n4407), .A2(n4273), .ZN(n4248) );
  INV_X1 U4882 ( .A(n4229), .ZN(n4230) );
  NOR2_X1 U4883 ( .A1(n4231), .A2(n4230), .ZN(n4314) );
  NAND2_X1 U4884 ( .A1(n4314), .A2(n4232), .ZN(n4287) );
  AOI21_X1 U4885 ( .B1(n4287), .B2(n4234), .A(n4233), .ZN(n4267) );
  NAND2_X1 U4886 ( .A1(n4267), .A2(n4270), .ZN(n4266) );
  NAND2_X1 U4887 ( .A1(n4235), .A2(n4266), .ZN(n4254) );
  NAND2_X1 U4888 ( .A1(n4255), .A2(n4254), .ZN(n4253) );
  NAND2_X1 U4889 ( .A1(n4236), .A2(n4253), .ZN(n4237) );
  XNOR2_X1 U4890 ( .A(n4238), .B(n4237), .ZN(n4239) );
  NAND2_X1 U4891 ( .A1(n4239), .A2(n4342), .ZN(n4242) );
  AOI22_X1 U4892 ( .A1(n4268), .A2(n4291), .B1(n4380), .B2(n4240), .ZN(n4241)
         );
  OAI211_X1 U4893 ( .C1(n4243), .C2(n4293), .A(n4242), .B(n4241), .ZN(n4406)
         );
  OAI22_X1 U4894 ( .A1(n4654), .A2(n4245), .B1(n4244), .B2(n4651), .ZN(n4246)
         );
  AOI21_X1 U4895 ( .B1(n4406), .B2(n4654), .A(n4246), .ZN(n4247) );
  OAI211_X1 U4896 ( .C1(n4485), .C2(n4328), .A(n4248), .B(n4247), .ZN(U3267)
         );
  NAND2_X1 U4897 ( .A1(n4278), .A2(n4257), .ZN(n4249) );
  NAND2_X1 U4898 ( .A1(n4250), .A2(n4249), .ZN(n4489) );
  AOI21_X1 U4899 ( .B1(n4255), .B2(n4252), .A(n4251), .ZN(n4411) );
  NAND2_X1 U4900 ( .A1(n4411), .A2(n4273), .ZN(n4265) );
  OAI21_X1 U4901 ( .B1(n4255), .B2(n4254), .A(n4253), .ZN(n4256) );
  NAND2_X1 U4902 ( .A1(n4256), .A2(n4342), .ZN(n4260) );
  AOI22_X1 U4903 ( .A1(n4258), .A2(n4291), .B1(n4257), .B2(n4380), .ZN(n4259)
         );
  OAI211_X1 U4904 ( .C1(n4400), .C2(n4293), .A(n4260), .B(n4259), .ZN(n4410)
         );
  INV_X1 U4905 ( .A(n4410), .ZN(n4262) );
  OAI22_X1 U4906 ( .A1(n4262), .A2(n4663), .B1(n4261), .B2(n4651), .ZN(n4263)
         );
  AOI21_X1 U4907 ( .B1(REG2_REG_22__SCAN_IN), .B2(n4663), .A(n4263), .ZN(n4264) );
  OAI211_X1 U4908 ( .C1(n4489), .C2(n4328), .A(n4265), .B(n4264), .ZN(U3268)
         );
  OAI21_X1 U4909 ( .B1(n4270), .B2(n4267), .A(n4266), .ZN(n4269) );
  AOI22_X1 U4910 ( .A1(n4269), .A2(n4342), .B1(n4362), .B2(n4268), .ZN(n4414)
         );
  INV_X1 U4911 ( .A(n4270), .ZN(n4272) );
  XOR2_X1 U4912 ( .A(n4272), .B(n4271), .Z(n4419) );
  NAND2_X1 U4913 ( .A1(n4419), .A2(n4273), .ZN(n4284) );
  INV_X1 U4914 ( .A(n4274), .ZN(n4275) );
  AOI22_X1 U4915 ( .A1(n4663), .A2(REG2_REG_21__SCAN_IN), .B1(n4275), .B2(
        n4643), .ZN(n4276) );
  OAI21_X1 U4916 ( .B1(n4416), .B2(n4277), .A(n4276), .ZN(n4280) );
  OAI21_X1 U4917 ( .B1(n4299), .B2(n4415), .A(n4278), .ZN(n4493) );
  NOR2_X1 U4918 ( .A1(n4493), .A2(n4328), .ZN(n4279) );
  AOI211_X1 U4919 ( .C1(n4282), .C2(n4281), .A(n4280), .B(n4279), .ZN(n4283)
         );
  OAI211_X1 U4920 ( .C1(n4663), .C2(n4414), .A(n4284), .B(n4283), .ZN(U3269)
         );
  XNOR2_X1 U4921 ( .A(n4285), .B(n4288), .ZN(n4422) );
  NAND2_X1 U4922 ( .A1(n4287), .A2(n4286), .ZN(n4289) );
  XNOR2_X1 U4923 ( .A(n4289), .B(n4288), .ZN(n4296) );
  AOI22_X1 U4924 ( .A1(n4339), .A2(n4291), .B1(n4380), .B2(n4290), .ZN(n4292)
         );
  OAI21_X1 U4925 ( .B1(n4294), .B2(n4293), .A(n4292), .ZN(n4295) );
  AOI21_X1 U4926 ( .B1(n4296), .B2(n4342), .A(n4295), .ZN(n4297) );
  OAI21_X1 U4927 ( .B1(n4422), .B2(n4298), .A(n4297), .ZN(n4423) );
  NAND2_X1 U4928 ( .A1(n4423), .A2(n4654), .ZN(n4308) );
  INV_X1 U4929 ( .A(n4326), .ZN(n4302) );
  INV_X1 U4930 ( .A(n4299), .ZN(n4300) );
  OAI21_X1 U4931 ( .B1(n4302), .B2(n4301), .A(n4300), .ZN(n4497) );
  INV_X1 U4932 ( .A(n4497), .ZN(n4306) );
  INV_X1 U4933 ( .A(REG2_REG_20__SCAN_IN), .ZN(n4304) );
  OAI22_X1 U4934 ( .A1(n4654), .A2(n4304), .B1(n4303), .B2(n4651), .ZN(n4305)
         );
  AOI21_X1 U4935 ( .B1(n4306), .B2(n4657), .A(n4305), .ZN(n4307) );
  OAI211_X1 U4936 ( .C1(n4422), .C2(n4309), .A(n4308), .B(n4307), .ZN(U3270)
         );
  XNOR2_X1 U4937 ( .A(n4311), .B(n4310), .ZN(n4428) );
  INV_X1 U4938 ( .A(n4428), .ZN(n4333) );
  INV_X1 U4939 ( .A(n4312), .ZN(n4313) );
  NOR2_X1 U4940 ( .A1(n4314), .A2(n4313), .ZN(n4338) );
  INV_X1 U4941 ( .A(n4315), .ZN(n4316) );
  AOI21_X1 U4942 ( .B1(n4338), .B2(n4317), .A(n4316), .ZN(n4319) );
  XNOR2_X1 U4943 ( .A(n4319), .B(n4318), .ZN(n4320) );
  NAND2_X1 U4944 ( .A1(n4320), .A2(n4342), .ZN(n4324) );
  NOR2_X1 U4945 ( .A1(n4433), .A2(n4327), .ZN(n4321) );
  AOI21_X1 U4946 ( .B1(n4322), .B2(n4362), .A(n4321), .ZN(n4323) );
  OAI211_X1 U4947 ( .C1(n4325), .C2(n4435), .A(n4324), .B(n4323), .ZN(n4427)
         );
  OAI21_X1 U4948 ( .B1(n2280), .B2(n4327), .A(n4326), .ZN(n4501) );
  NOR2_X1 U4949 ( .A1(n4501), .A2(n4328), .ZN(n4331) );
  OAI22_X1 U4950 ( .A1(n4654), .A2(n4106), .B1(n4329), .B2(n4651), .ZN(n4330)
         );
  AOI211_X1 U4951 ( .C1(n4427), .C2(n4654), .A(n4331), .B(n4330), .ZN(n4332)
         );
  OAI21_X1 U4952 ( .B1(n4333), .B2(n4353), .A(n4332), .ZN(U3271) );
  OAI21_X1 U4953 ( .B1(n4335), .B2(n4337), .A(n4334), .ZN(n4336) );
  INV_X1 U4954 ( .A(n4336), .ZN(n4432) );
  XNOR2_X1 U4955 ( .A(n4338), .B(n4337), .ZN(n4343) );
  AOI22_X1 U4956 ( .A1(n4339), .A2(n4362), .B1(n4380), .B2(n4558), .ZN(n4340)
         );
  OAI21_X1 U4957 ( .B1(n4533), .B2(n4435), .A(n4340), .ZN(n4341) );
  AOI21_X1 U4958 ( .B1(n4343), .B2(n4342), .A(n4341), .ZN(n4431) );
  INV_X1 U4959 ( .A(n4431), .ZN(n4351) );
  OAI211_X1 U4960 ( .C1(n2278), .C2(n4346), .A(n4701), .B(n4345), .ZN(n4430)
         );
  NOR2_X1 U4961 ( .A1(n4430), .A2(n4347), .ZN(n4350) );
  OAI22_X1 U4962 ( .A1(n4654), .A2(n4348), .B1(n4562), .B2(n4651), .ZN(n4349)
         );
  AOI211_X1 U4963 ( .C1(n4351), .C2(n4654), .A(n4350), .B(n4349), .ZN(n4352)
         );
  OAI21_X1 U4964 ( .B1(n4432), .B2(n4353), .A(n4352), .ZN(U3272) );
  XNOR2_X1 U4965 ( .A(n4354), .B(n2809), .ZN(n4367) );
  NAND2_X1 U4966 ( .A1(n4357), .A2(n4356), .ZN(n4358) );
  NAND2_X1 U4967 ( .A1(n4355), .A2(n4358), .ZN(n4686) );
  NAND2_X1 U4968 ( .A1(n4686), .A2(n4359), .ZN(n4365) );
  NOR2_X1 U4969 ( .A1(n4360), .A2(n4433), .ZN(n4361) );
  AOI21_X1 U4970 ( .B1(n4363), .B2(n4362), .A(n4361), .ZN(n4364) );
  OAI211_X1 U4971 ( .C1(n4367), .C2(n4366), .A(n4365), .B(n2273), .ZN(n4684)
         );
  MUX2_X1 U4972 ( .A(n4684), .B(REG2_REG_2__SCAN_IN), .S(n4663), .Z(n4368) );
  INV_X1 U4973 ( .A(n4368), .ZN(n4373) );
  AOI22_X1 U4974 ( .A1(n4658), .A2(n4686), .B1(REG3_REG_2__SCAN_IN), .B2(n4643), .ZN(n4372) );
  NAND2_X1 U4975 ( .A1(n4370), .A2(n4369), .ZN(n4682) );
  NAND3_X1 U4976 ( .A1(n4657), .A2(n4683), .A3(n4682), .ZN(n4371) );
  NAND3_X1 U4977 ( .A1(n4373), .A2(n4372), .A3(n4371), .ZN(U3288) );
  NAND2_X1 U4978 ( .A1(n4716), .A2(n4459), .ZN(n4375) );
  NAND2_X1 U4979 ( .A1(n4713), .A2(REG1_REG_31__SCAN_IN), .ZN(n4374) );
  OAI211_X1 U4980 ( .C1(n4462), .C2(n4458), .A(n4375), .B(n4374), .ZN(U3549)
         );
  AOI21_X1 U4981 ( .B1(n4381), .B2(n4377), .A(n4376), .ZN(n4564) );
  INV_X1 U4982 ( .A(n4564), .ZN(n4465) );
  INV_X1 U4983 ( .A(REG1_REG_30__SCAN_IN), .ZN(n4382) );
  INV_X1 U4984 ( .A(n4378), .ZN(n4379) );
  AOI21_X1 U4985 ( .B1(n4381), .B2(n4380), .A(n4379), .ZN(n4566) );
  MUX2_X1 U4986 ( .A(n4382), .B(n4566), .S(n4716), .Z(n4383) );
  OAI21_X1 U4987 ( .B1(n4465), .B2(n4458), .A(n4383), .ZN(U3548) );
  INV_X1 U4988 ( .A(REG1_REG_27__SCAN_IN), .ZN(n4389) );
  OAI22_X1 U4989 ( .A1(n4385), .A2(n4435), .B1(n4384), .B2(n4433), .ZN(n4386)
         );
  AOI211_X1 U4990 ( .C1(n4388), .C2(n4694), .A(n4387), .B(n4386), .ZN(n4466)
         );
  MUX2_X1 U4991 ( .A(n4389), .B(n4466), .S(n4716), .Z(n4390) );
  OAI21_X1 U4992 ( .B1(n4458), .B2(n4469), .A(n4390), .ZN(U3545) );
  INV_X1 U4993 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4393) );
  AOI21_X1 U4994 ( .B1(n4392), .B2(n4694), .A(n4391), .ZN(n4470) );
  MUX2_X1 U4995 ( .A(n4393), .B(n4470), .S(n4716), .Z(n4394) );
  OAI21_X1 U4996 ( .B1(n4458), .B2(n4473), .A(n4394), .ZN(U3544) );
  INV_X1 U4997 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4397) );
  AOI21_X1 U4998 ( .B1(n4396), .B2(n4694), .A(n4395), .ZN(n4474) );
  MUX2_X1 U4999 ( .A(n4397), .B(n4474), .S(n4716), .Z(n4398) );
  OAI21_X1 U5000 ( .B1(n4458), .B2(n4477), .A(n4398), .ZN(U3543) );
  INV_X1 U5001 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4404) );
  OAI22_X1 U5002 ( .A1(n4400), .A2(n4435), .B1(n4433), .B2(n4399), .ZN(n4401)
         );
  AOI211_X1 U5003 ( .C1(n4403), .C2(n4694), .A(n4402), .B(n4401), .ZN(n4478)
         );
  MUX2_X1 U5004 ( .A(n4404), .B(n4478), .S(n4716), .Z(n4405) );
  OAI21_X1 U5005 ( .B1(n4458), .B2(n4481), .A(n4405), .ZN(U3542) );
  INV_X1 U5006 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4408) );
  AOI21_X1 U5007 ( .B1(n4407), .B2(n4694), .A(n4406), .ZN(n4482) );
  MUX2_X1 U5008 ( .A(n4408), .B(n4482), .S(n4716), .Z(n4409) );
  OAI21_X1 U5009 ( .B1(n4458), .B2(n4485), .A(n4409), .ZN(U3541) );
  INV_X1 U5010 ( .A(REG1_REG_22__SCAN_IN), .ZN(n4412) );
  AOI21_X1 U5011 ( .B1(n4411), .B2(n4694), .A(n4410), .ZN(n4486) );
  MUX2_X1 U5012 ( .A(n4412), .B(n4486), .S(n4716), .Z(n4413) );
  OAI21_X1 U5013 ( .B1(n4458), .B2(n4489), .A(n4413), .ZN(U3540) );
  INV_X1 U5014 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4420) );
  INV_X1 U5015 ( .A(n4414), .ZN(n4418) );
  OAI22_X1 U5016 ( .A1(n4416), .A2(n4435), .B1(n4433), .B2(n4415), .ZN(n4417)
         );
  AOI211_X1 U5017 ( .C1(n4419), .C2(n4694), .A(n4418), .B(n4417), .ZN(n4490)
         );
  MUX2_X1 U5018 ( .A(n4420), .B(n4490), .S(n4716), .Z(n4421) );
  OAI21_X1 U5019 ( .B1(n4458), .B2(n4493), .A(n4421), .ZN(U3539) );
  INV_X1 U5020 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4425) );
  INV_X1 U5021 ( .A(n4422), .ZN(n4424) );
  AOI21_X1 U5022 ( .B1(n4690), .B2(n4424), .A(n4423), .ZN(n4494) );
  MUX2_X1 U5023 ( .A(n4425), .B(n4494), .S(n4716), .Z(n4426) );
  OAI21_X1 U5024 ( .B1(n4458), .B2(n4497), .A(n4426), .ZN(U3538) );
  AOI21_X1 U5025 ( .B1(n4428), .B2(n4694), .A(n4427), .ZN(n4498) );
  MUX2_X1 U5026 ( .A(n4109), .B(n4498), .S(n4716), .Z(n4429) );
  OAI21_X1 U5027 ( .B1(n4458), .B2(n4501), .A(n4429), .ZN(U3537) );
  OAI211_X1 U5028 ( .C1(n4432), .C2(n4441), .A(n4431), .B(n4430), .ZN(n4502)
         );
  MUX2_X1 U5029 ( .A(REG1_REG_18__SCAN_IN), .B(n4502), .S(n4716), .Z(U3536) );
  OAI22_X1 U5030 ( .A1(n4436), .A2(n4435), .B1(n4434), .B2(n4433), .ZN(n4437)
         );
  AOI211_X1 U5031 ( .C1(n4439), .C2(n4694), .A(n4438), .B(n4437), .ZN(n4503)
         );
  MUX2_X1 U5032 ( .A(n4083), .B(n4503), .S(n4716), .Z(n4440) );
  OAI21_X1 U5033 ( .B1(n4458), .B2(n4506), .A(n4440), .ZN(U3535) );
  OR2_X1 U5034 ( .A1(n4442), .A2(n4441), .ZN(n4444) );
  NAND2_X1 U5035 ( .A1(n4444), .A2(n4443), .ZN(n4507) );
  MUX2_X1 U5036 ( .A(REG1_REG_16__SCAN_IN), .B(n4507), .S(n4716), .Z(n4445) );
  INV_X1 U5037 ( .A(n4445), .ZN(n4446) );
  OAI21_X1 U5038 ( .B1(n4458), .B2(n4508), .A(n4446), .ZN(U3534) );
  INV_X1 U5039 ( .A(n4447), .ZN(n4452) );
  NAND3_X1 U5040 ( .A1(n4449), .A2(n4701), .A3(n4448), .ZN(n4450) );
  OAI211_X1 U5041 ( .C1(n4452), .C2(n4696), .A(n4451), .B(n4450), .ZN(n4511)
         );
  MUX2_X1 U5042 ( .A(REG1_REG_14__SCAN_IN), .B(n4511), .S(n4716), .Z(U3532) );
  INV_X1 U5043 ( .A(REG1_REG_13__SCAN_IN), .ZN(n4456) );
  INV_X1 U5044 ( .A(n4453), .ZN(n4454) );
  AOI21_X1 U5045 ( .B1(n4455), .B2(n4694), .A(n4454), .ZN(n4512) );
  MUX2_X1 U5046 ( .A(n4456), .B(n4512), .S(n4716), .Z(n4457) );
  OAI21_X1 U5047 ( .B1(n4458), .B2(n4516), .A(n4457), .ZN(U3531) );
  NAND2_X1 U5048 ( .A1(n4704), .A2(n4459), .ZN(n4461) );
  NAND2_X1 U5049 ( .A1(n4702), .A2(REG0_REG_31__SCAN_IN), .ZN(n4460) );
  OAI211_X1 U5050 ( .C1(n4462), .C2(n4515), .A(n4461), .B(n4460), .ZN(U3517)
         );
  INV_X1 U5051 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4463) );
  MUX2_X1 U5052 ( .A(n4463), .B(n4566), .S(n4704), .Z(n4464) );
  OAI21_X1 U5053 ( .B1(n4465), .B2(n4515), .A(n4464), .ZN(U3516) );
  INV_X1 U5054 ( .A(REG0_REG_27__SCAN_IN), .ZN(n4467) );
  MUX2_X1 U5055 ( .A(n4467), .B(n4466), .S(n4704), .Z(n4468) );
  OAI21_X1 U5056 ( .B1(n4469), .B2(n4515), .A(n4468), .ZN(U3513) );
  INV_X1 U5057 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4471) );
  MUX2_X1 U5058 ( .A(n4471), .B(n4470), .S(n4704), .Z(n4472) );
  OAI21_X1 U5059 ( .B1(n4473), .B2(n4515), .A(n4472), .ZN(U3512) );
  INV_X1 U5060 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4475) );
  MUX2_X1 U5061 ( .A(n4475), .B(n4474), .S(n4704), .Z(n4476) );
  OAI21_X1 U5062 ( .B1(n4477), .B2(n4515), .A(n4476), .ZN(U3511) );
  INV_X1 U5063 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4479) );
  MUX2_X1 U5064 ( .A(n4479), .B(n4478), .S(n4704), .Z(n4480) );
  OAI21_X1 U5065 ( .B1(n4481), .B2(n4515), .A(n4480), .ZN(U3510) );
  INV_X1 U5066 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4483) );
  MUX2_X1 U5067 ( .A(n4483), .B(n4482), .S(n4704), .Z(n4484) );
  OAI21_X1 U5068 ( .B1(n4485), .B2(n4515), .A(n4484), .ZN(U3509) );
  INV_X1 U5069 ( .A(REG0_REG_22__SCAN_IN), .ZN(n4487) );
  MUX2_X1 U5070 ( .A(n4487), .B(n4486), .S(n4704), .Z(n4488) );
  OAI21_X1 U5071 ( .B1(n4489), .B2(n4515), .A(n4488), .ZN(U3508) );
  INV_X1 U5072 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4491) );
  MUX2_X1 U5073 ( .A(n4491), .B(n4490), .S(n4704), .Z(n4492) );
  OAI21_X1 U5074 ( .B1(n4493), .B2(n4515), .A(n4492), .ZN(U3507) );
  INV_X1 U5075 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4495) );
  MUX2_X1 U5076 ( .A(n4495), .B(n4494), .S(n4704), .Z(n4496) );
  OAI21_X1 U5077 ( .B1(n4497), .B2(n4515), .A(n4496), .ZN(U3506) );
  INV_X1 U5078 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4499) );
  MUX2_X1 U5079 ( .A(n4499), .B(n4498), .S(n4704), .Z(n4500) );
  OAI21_X1 U5080 ( .B1(n4501), .B2(n4515), .A(n4500), .ZN(U3505) );
  MUX2_X1 U5081 ( .A(REG0_REG_18__SCAN_IN), .B(n4502), .S(n4704), .Z(U3503) );
  INV_X1 U5082 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4504) );
  MUX2_X1 U5083 ( .A(n4504), .B(n4503), .S(n4704), .Z(n4505) );
  OAI21_X1 U5084 ( .B1(n4506), .B2(n4515), .A(n4505), .ZN(U3501) );
  MUX2_X1 U5085 ( .A(REG0_REG_16__SCAN_IN), .B(n4507), .S(n4704), .Z(n4510) );
  NOR2_X1 U5086 ( .A1(n4508), .A2(n4515), .ZN(n4509) );
  MUX2_X1 U5087 ( .A(REG0_REG_14__SCAN_IN), .B(n4511), .S(n4704), .Z(U3495) );
  INV_X1 U5088 ( .A(REG0_REG_13__SCAN_IN), .ZN(n4513) );
  MUX2_X1 U5089 ( .A(n4513), .B(n4512), .S(n4704), .Z(n4514) );
  OAI21_X1 U5090 ( .B1(n4516), .B2(n4515), .A(n4514), .ZN(U3493) );
  MUX2_X1 U5091 ( .A(n4517), .B(DATAI_29_), .S(U3149), .Z(U3323) );
  MUX2_X1 U5092 ( .A(n4518), .B(DATAI_21_), .S(U3149), .Z(U3331) );
  MUX2_X1 U5093 ( .A(DATAI_19_), .B(n4519), .S(STATE_REG_SCAN_IN), .Z(U3333)
         );
  MUX2_X1 U5094 ( .A(n4520), .B(DATAI_18_), .S(U3149), .Z(U3334) );
  MUX2_X1 U5095 ( .A(n4521), .B(DATAI_13_), .S(U3149), .Z(U3339) );
  MUX2_X1 U5096 ( .A(n4522), .B(DATAI_11_), .S(U3149), .Z(U3341) );
  MUX2_X1 U5097 ( .A(n4567), .B(DATAI_9_), .S(U3149), .Z(U3343) );
  MUX2_X1 U5098 ( .A(n4523), .B(DATAI_7_), .S(U3149), .Z(U3345) );
  MUX2_X1 U5099 ( .A(n4524), .B(DATAI_6_), .S(U3149), .Z(U3346) );
  MUX2_X1 U5100 ( .A(n4525), .B(DATAI_5_), .S(U3149), .Z(U3347) );
  MUX2_X1 U5101 ( .A(DATAI_4_), .B(n4526), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U5102 ( .A(n4527), .B(DATAI_3_), .S(U3149), .Z(U3349) );
  OAI22_X1 U5103 ( .A1(n4531), .A2(n4530), .B1(n4529), .B2(n4528), .ZN(n4535)
         );
  NOR2_X1 U5104 ( .A1(STATE_REG_SCAN_IN), .A2(n5067), .ZN(n4624) );
  INV_X1 U5105 ( .A(n4624), .ZN(n4532) );
  OAI21_X1 U5106 ( .B1(n4546), .B2(n4533), .A(n4532), .ZN(n4534) );
  NOR2_X1 U5107 ( .A1(n4535), .A2(n4534), .ZN(n4542) );
  INV_X1 U5108 ( .A(n3802), .ZN(n4537) );
  OAI21_X1 U5109 ( .B1(n4537), .B2(n4536), .A(n3803), .ZN(n4539) );
  XNOR2_X1 U5110 ( .A(n4539), .B(n4538), .ZN(n4540) );
  NAND2_X1 U5111 ( .A1(n4540), .A2(n4554), .ZN(n4541) );
  OAI211_X1 U5112 ( .C1(n4563), .C2(n4543), .A(n4542), .B(n4541), .ZN(U3223)
         );
  OAI22_X1 U5113 ( .A1(n4546), .A2(n4545), .B1(STATE_REG_SCAN_IN), .B2(n4544), 
        .ZN(n4547) );
  INV_X1 U5114 ( .A(n4547), .ZN(n4561) );
  INV_X1 U5115 ( .A(n4549), .ZN(n4552) );
  AND2_X1 U5116 ( .A1(n4549), .A2(n4548), .ZN(n4551) );
  OAI22_X1 U5117 ( .A1(n4553), .A2(n4552), .B1(n4551), .B2(n4550), .ZN(n4555)
         );
  AOI222_X1 U5118 ( .A1(n4559), .A2(n4558), .B1(n4557), .B2(n4556), .C1(n4555), 
        .C2(n4554), .ZN(n4560) );
  OAI211_X1 U5119 ( .C1(n4563), .C2(n4562), .A(n4561), .B(n4560), .ZN(U3235)
         );
  AOI22_X1 U5120 ( .A1(n4564), .A2(n4657), .B1(REG2_REG_30__SCAN_IN), .B2(
        n4663), .ZN(n4565) );
  OAI21_X1 U5121 ( .B1(n4663), .B2(n4566), .A(n4565), .ZN(U3261) );
  INV_X1 U5122 ( .A(n4567), .ZN(n4576) );
  OAI211_X1 U5123 ( .C1(n4570), .C2(n4569), .A(n4637), .B(n4568), .ZN(n4575)
         );
  OAI211_X1 U5124 ( .C1(n4573), .C2(n4572), .A(n4593), .B(n4571), .ZN(n4574)
         );
  OAI211_X1 U5125 ( .C1(n4642), .C2(n4576), .A(n4575), .B(n4574), .ZN(n4577)
         );
  AOI211_X1 U5126 ( .C1(n4636), .C2(ADDR_REG_9__SCAN_IN), .A(n4578), .B(n4577), 
        .ZN(n4579) );
  INV_X1 U5127 ( .A(n4579), .ZN(U3249) );
  OAI211_X1 U5128 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4581), .A(n4593), .B(n4580), .ZN(n4583) );
  NAND2_X1 U5129 ( .A1(n4583), .A2(n4582), .ZN(n4584) );
  AOI21_X1 U5130 ( .B1(n4636), .B2(ADDR_REG_10__SCAN_IN), .A(n4584), .ZN(n4588) );
  OAI211_X1 U5131 ( .C1(REG1_REG_10__SCAN_IN), .C2(n4586), .A(n4637), .B(n4585), .ZN(n4587) );
  OAI211_X1 U5132 ( .C1(n4642), .C2(n4672), .A(n4588), .B(n4587), .ZN(U3250)
         );
  OAI211_X1 U5133 ( .C1(n4591), .C2(n4590), .A(n4589), .B(n4637), .ZN(n4597)
         );
  OAI211_X1 U5134 ( .C1(n4595), .C2(n4594), .A(n4593), .B(n4592), .ZN(n4596)
         );
  OAI211_X1 U5135 ( .C1(n4642), .C2(n4598), .A(n4597), .B(n4596), .ZN(n4599)
         );
  AOI211_X1 U5136 ( .C1(n4636), .C2(ADDR_REG_11__SCAN_IN), .A(n4600), .B(n4599), .ZN(n4601) );
  INV_X1 U5137 ( .A(n4601), .ZN(U3251) );
  INV_X1 U5138 ( .A(n4602), .ZN(n4606) );
  AOI211_X1 U5139 ( .C1(n3437), .C2(n4604), .A(n4603), .B(n4630), .ZN(n4605)
         );
  AOI211_X1 U5140 ( .C1(n4636), .C2(ADDR_REG_14__SCAN_IN), .A(n4606), .B(n4605), .ZN(n4610) );
  OAI211_X1 U5141 ( .C1(REG1_REG_14__SCAN_IN), .C2(n4608), .A(n4637), .B(n4607), .ZN(n4609) );
  OAI211_X1 U5142 ( .C1(n4642), .C2(n4671), .A(n4610), .B(n4609), .ZN(U3254)
         );
  AOI211_X1 U5143 ( .C1(n4613), .C2(n4612), .A(n4611), .B(n4630), .ZN(n4614)
         );
  AOI211_X1 U5144 ( .C1(n4636), .C2(ADDR_REG_15__SCAN_IN), .A(n4615), .B(n4614), .ZN(n4620) );
  OAI211_X1 U5145 ( .C1(n4618), .C2(n4617), .A(n4637), .B(n4616), .ZN(n4619)
         );
  OAI211_X1 U5146 ( .C1(n4642), .C2(n4670), .A(n4620), .B(n4619), .ZN(U3255)
         );
  AOI221_X1 U5147 ( .B1(n4622), .B2(n4621), .C1(n3506), .C2(n4621), .A(n4630), 
        .ZN(n4623) );
  AOI211_X1 U5148 ( .C1(n4636), .C2(ADDR_REG_16__SCAN_IN), .A(n4624), .B(n4623), .ZN(n4628) );
  OAI221_X1 U5149 ( .B1(n4626), .B2(REG1_REG_16__SCAN_IN), .C1(n4626), .C2(
        n4625), .A(n4637), .ZN(n4627) );
  OAI211_X1 U5150 ( .C1(n4642), .C2(n4629), .A(n4628), .B(n4627), .ZN(U3256)
         );
  AOI221_X1 U5151 ( .B1(n4633), .B2(n4632), .C1(n4631), .C2(n4632), .A(n4630), 
        .ZN(n4634) );
  AOI211_X1 U5152 ( .C1(n4636), .C2(ADDR_REG_17__SCAN_IN), .A(n4635), .B(n4634), .ZN(n4641) );
  OAI221_X1 U5153 ( .B1(n4639), .B2(n2259), .C1(n4639), .C2(n4638), .A(n4637), 
        .ZN(n4640) );
  OAI211_X1 U5154 ( .C1(n4642), .C2(n4667), .A(n4641), .B(n4640), .ZN(U3257)
         );
  AOI22_X1 U5155 ( .A1(n4644), .A2(n4643), .B1(REG2_REG_10__SCAN_IN), .B2(
        n4663), .ZN(n4649) );
  INV_X1 U5156 ( .A(n4645), .ZN(n4646) );
  AOI22_X1 U5157 ( .A1(n4647), .A2(n4658), .B1(n4657), .B2(n4646), .ZN(n4648)
         );
  OAI211_X1 U5158 ( .C1(n4663), .C2(n4650), .A(n4649), .B(n4648), .ZN(U3280)
         );
  OAI22_X1 U5159 ( .A1(n4654), .A2(n4653), .B1(n4652), .B2(n4651), .ZN(n4655)
         );
  INV_X1 U5160 ( .A(n4655), .ZN(n4661) );
  AOI22_X1 U5161 ( .A1(n4659), .A2(n4658), .B1(n4657), .B2(n4656), .ZN(n4660)
         );
  OAI211_X1 U5162 ( .C1(n4663), .C2(n4662), .A(n4661), .B(n4660), .ZN(U3282)
         );
  INV_X1 U5163 ( .A(D_REG_31__SCAN_IN), .ZN(n5032) );
  NOR2_X1 U5164 ( .A1(n4665), .A2(n5032), .ZN(U3291) );
  INV_X1 U5165 ( .A(D_REG_30__SCAN_IN), .ZN(n5029) );
  NOR2_X1 U5166 ( .A1(n4665), .A2(n5029), .ZN(U3292) );
  AND2_X1 U5167 ( .A1(n4664), .A2(D_REG_29__SCAN_IN), .ZN(U3293) );
  INV_X1 U5168 ( .A(D_REG_28__SCAN_IN), .ZN(n5054) );
  NOR2_X1 U5169 ( .A1(n4665), .A2(n5054), .ZN(U3294) );
  AND2_X1 U5170 ( .A1(n4664), .A2(D_REG_27__SCAN_IN), .ZN(U3295) );
  INV_X1 U5171 ( .A(D_REG_26__SCAN_IN), .ZN(n5025) );
  NOR2_X1 U5172 ( .A1(n4665), .A2(n5025), .ZN(U3296) );
  INV_X1 U5173 ( .A(D_REG_25__SCAN_IN), .ZN(n5045) );
  NOR2_X1 U5174 ( .A1(n4665), .A2(n5045), .ZN(U3297) );
  INV_X1 U5175 ( .A(D_REG_24__SCAN_IN), .ZN(n4743) );
  NOR2_X1 U5176 ( .A1(n4665), .A2(n4743), .ZN(U3298) );
  AND2_X1 U5177 ( .A1(n4664), .A2(D_REG_23__SCAN_IN), .ZN(U3299) );
  AND2_X1 U5178 ( .A1(n4664), .A2(D_REG_22__SCAN_IN), .ZN(U3300) );
  AND2_X1 U5179 ( .A1(n4664), .A2(D_REG_21__SCAN_IN), .ZN(U3301) );
  INV_X1 U5180 ( .A(D_REG_20__SCAN_IN), .ZN(n5038) );
  NOR2_X1 U5181 ( .A1(n4665), .A2(n5038), .ZN(U3302) );
  INV_X1 U5182 ( .A(D_REG_19__SCAN_IN), .ZN(n5044) );
  NOR2_X1 U5183 ( .A1(n4665), .A2(n5044), .ZN(U3303) );
  INV_X1 U5184 ( .A(D_REG_18__SCAN_IN), .ZN(n5041) );
  NOR2_X1 U5185 ( .A1(n4665), .A2(n5041), .ZN(U3304) );
  AND2_X1 U5186 ( .A1(n4664), .A2(D_REG_17__SCAN_IN), .ZN(U3305) );
  AND2_X1 U5187 ( .A1(n4664), .A2(D_REG_16__SCAN_IN), .ZN(U3306) );
  INV_X1 U5188 ( .A(D_REG_15__SCAN_IN), .ZN(n5026) );
  NOR2_X1 U5189 ( .A1(n4665), .A2(n5026), .ZN(U3307) );
  INV_X1 U5190 ( .A(D_REG_14__SCAN_IN), .ZN(n4827) );
  NOR2_X1 U5191 ( .A1(n4665), .A2(n4827), .ZN(U3308) );
  INV_X1 U5192 ( .A(D_REG_13__SCAN_IN), .ZN(n5028) );
  NOR2_X1 U5193 ( .A1(n4665), .A2(n5028), .ZN(U3309) );
  INV_X1 U5194 ( .A(D_REG_12__SCAN_IN), .ZN(n5031) );
  NOR2_X1 U5195 ( .A1(n4665), .A2(n5031), .ZN(U3310) );
  INV_X1 U5196 ( .A(D_REG_11__SCAN_IN), .ZN(n5039) );
  NOR2_X1 U5197 ( .A1(n4665), .A2(n5039), .ZN(U3311) );
  INV_X1 U5198 ( .A(D_REG_10__SCAN_IN), .ZN(n5048) );
  NOR2_X1 U5199 ( .A1(n4665), .A2(n5048), .ZN(U3312) );
  INV_X1 U5200 ( .A(D_REG_9__SCAN_IN), .ZN(n4792) );
  NOR2_X1 U5201 ( .A1(n4665), .A2(n4792), .ZN(U3313) );
  INV_X1 U5202 ( .A(D_REG_8__SCAN_IN), .ZN(n4877) );
  NOR2_X1 U5203 ( .A1(n4665), .A2(n4877), .ZN(U3314) );
  INV_X1 U5204 ( .A(D_REG_7__SCAN_IN), .ZN(n5042) );
  NOR2_X1 U5205 ( .A1(n4665), .A2(n5042), .ZN(U3315) );
  INV_X1 U5206 ( .A(D_REG_6__SCAN_IN), .ZN(n5047) );
  NOR2_X1 U5207 ( .A1(n4665), .A2(n5047), .ZN(U3316) );
  INV_X1 U5208 ( .A(D_REG_5__SCAN_IN), .ZN(n5092) );
  NOR2_X1 U5209 ( .A1(n4665), .A2(n5092), .ZN(U3317) );
  INV_X1 U5210 ( .A(D_REG_4__SCAN_IN), .ZN(n5022) );
  NOR2_X1 U5211 ( .A1(n4665), .A2(n5022), .ZN(U3318) );
  INV_X1 U5212 ( .A(D_REG_3__SCAN_IN), .ZN(n4834) );
  NOR2_X1 U5213 ( .A1(n4665), .A2(n4834), .ZN(U3319) );
  INV_X1 U5214 ( .A(D_REG_2__SCAN_IN), .ZN(n4845) );
  NOR2_X1 U5215 ( .A1(n4665), .A2(n4845), .ZN(U3320) );
  INV_X1 U5216 ( .A(DATAI_23_), .ZN(n4971) );
  AOI21_X1 U5217 ( .B1(U3149), .B2(n4971), .A(n4666), .ZN(U3329) );
  AOI22_X1 U5218 ( .A1(STATE_REG_SCAN_IN), .A2(n4667), .B1(n4794), .B2(U3149), 
        .ZN(U3335) );
  OAI22_X1 U5219 ( .A1(U3149), .A2(n4668), .B1(DATAI_16_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4669) );
  INV_X1 U5220 ( .A(n4669), .ZN(U3336) );
  INV_X1 U5221 ( .A(DATAI_15_), .ZN(n4742) );
  AOI22_X1 U5222 ( .A1(STATE_REG_SCAN_IN), .A2(n4670), .B1(n4742), .B2(U3149), 
        .ZN(U3337) );
  INV_X1 U5223 ( .A(DATAI_14_), .ZN(n4981) );
  AOI22_X1 U5224 ( .A1(STATE_REG_SCAN_IN), .A2(n4671), .B1(n4981), .B2(U3149), 
        .ZN(U3338) );
  INV_X1 U5225 ( .A(DATAI_10_), .ZN(n4817) );
  AOI22_X1 U5226 ( .A1(STATE_REG_SCAN_IN), .A2(n4672), .B1(n4817), .B2(U3149), 
        .ZN(U3342) );
  OAI211_X1 U5227 ( .C1(n4675), .C2(n4696), .A(n4674), .B(n4673), .ZN(n4676)
         );
  INV_X1 U5228 ( .A(n4676), .ZN(n4705) );
  INV_X1 U5229 ( .A(REG0_REG_0__SCAN_IN), .ZN(n5006) );
  AOI22_X1 U5230 ( .A1(n4704), .A2(n4705), .B1(n5006), .B2(n4702), .ZN(U3467)
         );
  OAI22_X1 U5231 ( .A1(n4679), .A2(n4696), .B1(n4678), .B2(n4677), .ZN(n4681)
         );
  NOR2_X1 U5232 ( .A1(n4681), .A2(n4680), .ZN(n4706) );
  INV_X1 U5233 ( .A(REG0_REG_1__SCAN_IN), .ZN(n4864) );
  AOI22_X1 U5234 ( .A1(n4704), .A2(n4706), .B1(n4864), .B2(n4702), .ZN(U3469)
         );
  AND3_X1 U5235 ( .A1(n4683), .A2(n4701), .A3(n4682), .ZN(n4685) );
  AOI211_X1 U5236 ( .C1(n4690), .C2(n4686), .A(n4685), .B(n4684), .ZN(n4708)
         );
  INV_X1 U5237 ( .A(REG0_REG_2__SCAN_IN), .ZN(n5072) );
  AOI22_X1 U5238 ( .A1(n4704), .A2(n4708), .B1(n5072), .B2(n4702), .ZN(U3471)
         );
  INV_X1 U5239 ( .A(n4687), .ZN(n4689) );
  AOI211_X1 U5240 ( .C1(n4691), .C2(n4690), .A(n4689), .B(n4688), .ZN(n4710)
         );
  INV_X1 U5241 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4804) );
  AOI22_X1 U5242 ( .A1(n4704), .A2(n4710), .B1(n4804), .B2(n4702), .ZN(U3475)
         );
  AOI211_X1 U5243 ( .C1(n4695), .C2(n4694), .A(n4693), .B(n4692), .ZN(n4712)
         );
  INV_X1 U5244 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4996) );
  AOI22_X1 U5245 ( .A1(n4704), .A2(n4712), .B1(n4996), .B2(n4702), .ZN(U3481)
         );
  NOR2_X1 U5246 ( .A1(n4697), .A2(n4696), .ZN(n4699) );
  AOI211_X1 U5247 ( .C1(n4701), .C2(n4700), .A(n4699), .B(n4698), .ZN(n4715)
         );
  INV_X1 U5248 ( .A(REG0_REG_11__SCAN_IN), .ZN(n4703) );
  AOI22_X1 U5249 ( .A1(n4704), .A2(n4715), .B1(n4703), .B2(n4702), .ZN(U3489)
         );
  AOI22_X1 U5250 ( .A1(n4716), .A2(n4705), .B1(n2935), .B2(n4713), .ZN(U3518)
         );
  AOI22_X1 U5251 ( .A1(n4716), .A2(n4706), .B1(n3050), .B2(n4713), .ZN(U3519)
         );
  AOI22_X1 U5252 ( .A1(n4716), .A2(n4708), .B1(n4707), .B2(n4713), .ZN(U3520)
         );
  AOI22_X1 U5253 ( .A1(n4716), .A2(n4710), .B1(n4709), .B2(n4713), .ZN(U3522)
         );
  AOI22_X1 U5254 ( .A1(n4716), .A2(n4712), .B1(n4711), .B2(n4713), .ZN(U3525)
         );
  AOI22_X1 U5255 ( .A1(n4716), .A2(n4715), .B1(n4714), .B2(n4713), .ZN(U3529)
         );
  OAI22_X1 U5256 ( .A1(D_REG_13__SCAN_IN), .A2(keyinput_g100), .B1(
        keyinput_g40), .B2(REG3_REG_28__SCAN_IN), .ZN(n4717) );
  AOI221_X1 U5257 ( .B1(D_REG_13__SCAN_IN), .B2(keyinput_g100), .C1(
        REG3_REG_28__SCAN_IN), .C2(keyinput_g40), .A(n4717), .ZN(n4724) );
  OAI22_X1 U5258 ( .A1(REG3_REG_14__SCAN_IN), .A2(keyinput_g35), .B1(
        REG0_REG_2__SCAN_IN), .B2(keyinput_g121), .ZN(n4718) );
  AOI221_X1 U5259 ( .B1(REG3_REG_14__SCAN_IN), .B2(keyinput_g35), .C1(
        keyinput_g121), .C2(REG0_REG_2__SCAN_IN), .A(n4718), .ZN(n4723) );
  OAI22_X1 U5260 ( .A1(IR_REG_3__SCAN_IN), .A2(keyinput_g58), .B1(
        keyinput_g103), .B2(D_REG_16__SCAN_IN), .ZN(n4719) );
  AOI221_X1 U5261 ( .B1(IR_REG_3__SCAN_IN), .B2(keyinput_g58), .C1(
        D_REG_16__SCAN_IN), .C2(keyinput_g103), .A(n4719), .ZN(n4722) );
  OAI22_X1 U5262 ( .A1(IR_REG_5__SCAN_IN), .A2(keyinput_g60), .B1(
        REG3_REG_12__SCAN_IN), .B2(keyinput_g44), .ZN(n4720) );
  AOI221_X1 U5263 ( .B1(IR_REG_5__SCAN_IN), .B2(keyinput_g60), .C1(
        keyinput_g44), .C2(REG3_REG_12__SCAN_IN), .A(n4720), .ZN(n4721) );
  NAND4_X1 U5264 ( .A1(n4724), .A2(n4723), .A3(n4722), .A4(n4721), .ZN(n4755)
         );
  OAI22_X1 U5265 ( .A1(D_REG_29__SCAN_IN), .A2(keyinput_g116), .B1(DATAI_29_), 
        .B2(keyinput_g2), .ZN(n4725) );
  AOI221_X1 U5266 ( .B1(D_REG_29__SCAN_IN), .B2(keyinput_g116), .C1(
        keyinput_g2), .C2(DATAI_29_), .A(n4725), .ZN(n4732) );
  OAI22_X1 U5267 ( .A1(IR_REG_0__SCAN_IN), .A2(keyinput_g55), .B1(
        D_REG_23__SCAN_IN), .B2(keyinput_g110), .ZN(n4726) );
  AOI221_X1 U5268 ( .B1(IR_REG_0__SCAN_IN), .B2(keyinput_g55), .C1(
        keyinput_g110), .C2(D_REG_23__SCAN_IN), .A(n4726), .ZN(n4731) );
  OAI22_X1 U5269 ( .A1(IR_REG_20__SCAN_IN), .A2(keyinput_g75), .B1(
        keyinput_g11), .B2(DATAI_20_), .ZN(n4727) );
  AOI221_X1 U5270 ( .B1(IR_REG_20__SCAN_IN), .B2(keyinput_g75), .C1(DATAI_20_), 
        .C2(keyinput_g11), .A(n4727), .ZN(n4730) );
  OAI22_X1 U5271 ( .A1(DATAI_21_), .A2(keyinput_g10), .B1(REG0_REG_7__SCAN_IN), 
        .B2(keyinput_g126), .ZN(n4728) );
  AOI221_X1 U5272 ( .B1(DATAI_21_), .B2(keyinput_g10), .C1(keyinput_g126), 
        .C2(REG0_REG_7__SCAN_IN), .A(n4728), .ZN(n4729) );
  NAND4_X1 U5273 ( .A1(n4732), .A2(n4731), .A3(n4730), .A4(n4729), .ZN(n4754)
         );
  OAI22_X1 U5274 ( .A1(REG3_REG_25__SCAN_IN), .A2(keyinput_g45), .B1(DATAI_16_), .B2(keyinput_g15), .ZN(n4733) );
  AOI221_X1 U5275 ( .B1(REG3_REG_25__SCAN_IN), .B2(keyinput_g45), .C1(
        keyinput_g15), .C2(DATAI_16_), .A(n4733), .ZN(n4740) );
  OAI22_X1 U5276 ( .A1(IR_REG_30__SCAN_IN), .A2(keyinput_g85), .B1(
        keyinput_g49), .B2(REG3_REG_24__SCAN_IN), .ZN(n4734) );
  AOI221_X1 U5277 ( .B1(IR_REG_30__SCAN_IN), .B2(keyinput_g85), .C1(
        REG3_REG_24__SCAN_IN), .C2(keyinput_g49), .A(n4734), .ZN(n4739) );
  OAI22_X1 U5278 ( .A1(IR_REG_14__SCAN_IN), .A2(keyinput_g69), .B1(
        D_REG_12__SCAN_IN), .B2(keyinput_g99), .ZN(n4735) );
  AOI221_X1 U5279 ( .B1(IR_REG_14__SCAN_IN), .B2(keyinput_g69), .C1(
        keyinput_g99), .C2(D_REG_12__SCAN_IN), .A(n4735), .ZN(n4738) );
  OAI22_X1 U5280 ( .A1(REG3_REG_7__SCAN_IN), .A2(keyinput_g33), .B1(
        keyinput_g7), .B2(DATAI_24_), .ZN(n4736) );
  AOI221_X1 U5281 ( .B1(REG3_REG_7__SCAN_IN), .B2(keyinput_g33), .C1(DATAI_24_), .C2(keyinput_g7), .A(n4736), .ZN(n4737) );
  NAND4_X1 U5282 ( .A1(n4740), .A2(n4739), .A3(n4738), .A4(n4737), .ZN(n4753)
         );
  AOI22_X1 U5283 ( .A1(n4743), .A2(keyinput_g111), .B1(keyinput_g16), .B2(
        n4742), .ZN(n4741) );
  OAI221_X1 U5284 ( .B1(n4743), .B2(keyinput_g111), .C1(n4742), .C2(
        keyinput_g16), .A(n4741), .ZN(n4751) );
  AOI22_X1 U5285 ( .A1(REG3_REG_19__SCAN_IN), .A2(keyinput_g39), .B1(
        D_REG_27__SCAN_IN), .B2(keyinput_g114), .ZN(n4744) );
  OAI221_X1 U5286 ( .B1(REG3_REG_19__SCAN_IN), .B2(keyinput_g39), .C1(
        D_REG_27__SCAN_IN), .C2(keyinput_g114), .A(n4744), .ZN(n4750) );
  AOI22_X1 U5287 ( .A1(IR_REG_25__SCAN_IN), .A2(keyinput_g80), .B1(n2453), 
        .B2(keyinput_g65), .ZN(n4745) );
  OAI221_X1 U5288 ( .B1(IR_REG_25__SCAN_IN), .B2(keyinput_g80), .C1(n2453), 
        .C2(keyinput_g65), .A(n4745), .ZN(n4749) );
  XNOR2_X1 U5289 ( .A(IR_REG_31__SCAN_IN), .B(keyinput_g86), .ZN(n4747) );
  XNOR2_X1 U5290 ( .A(IR_REG_18__SCAN_IN), .B(keyinput_g73), .ZN(n4746) );
  NAND2_X1 U5291 ( .A1(n4747), .A2(n4746), .ZN(n4748) );
  OR4_X1 U5292 ( .A1(n4751), .A2(n4750), .A3(n4749), .A4(n4748), .ZN(n4752) );
  NOR4_X1 U5293 ( .A1(n4755), .A2(n4754), .A3(n4753), .A4(n4752), .ZN(n5095)
         );
  OAI22_X1 U5294 ( .A1(D_REG_22__SCAN_IN), .A2(keyinput_g109), .B1(
        keyinput_g42), .B2(REG3_REG_1__SCAN_IN), .ZN(n4756) );
  AOI221_X1 U5295 ( .B1(D_REG_22__SCAN_IN), .B2(keyinput_g109), .C1(
        REG3_REG_1__SCAN_IN), .C2(keyinput_g42), .A(n4756), .ZN(n4763) );
  OAI22_X1 U5296 ( .A1(D_REG_21__SCAN_IN), .A2(keyinput_g108), .B1(
        D_REG_17__SCAN_IN), .B2(keyinput_g104), .ZN(n4757) );
  AOI221_X1 U5297 ( .B1(D_REG_21__SCAN_IN), .B2(keyinput_g108), .C1(
        keyinput_g104), .C2(D_REG_17__SCAN_IN), .A(n4757), .ZN(n4762) );
  OAI22_X1 U5298 ( .A1(IR_REG_16__SCAN_IN), .A2(keyinput_g71), .B1(DATAI_12_), 
        .B2(keyinput_g19), .ZN(n4758) );
  AOI221_X1 U5299 ( .B1(IR_REG_16__SCAN_IN), .B2(keyinput_g71), .C1(
        keyinput_g19), .C2(DATAI_12_), .A(n4758), .ZN(n4761) );
  OAI22_X1 U5300 ( .A1(DATAI_8_), .A2(keyinput_g23), .B1(DATAI_5_), .B2(
        keyinput_g26), .ZN(n4759) );
  AOI221_X1 U5301 ( .B1(DATAI_8_), .B2(keyinput_g23), .C1(keyinput_g26), .C2(
        DATAI_5_), .A(n4759), .ZN(n4760) );
  NAND4_X1 U5302 ( .A1(n4763), .A2(n4762), .A3(n4761), .A4(n4760), .ZN(n4893)
         );
  AOI22_X1 U5303 ( .A1(REG0_REG_3__SCAN_IN), .A2(keyinput_g122), .B1(
        IR_REG_28__SCAN_IN), .B2(keyinput_g83), .ZN(n4764) );
  OAI221_X1 U5304 ( .B1(REG0_REG_3__SCAN_IN), .B2(keyinput_g122), .C1(
        IR_REG_28__SCAN_IN), .C2(keyinput_g83), .A(n4764), .ZN(n4771) );
  AOI22_X1 U5305 ( .A1(DATAI_14_), .A2(keyinput_g17), .B1(IR_REG_13__SCAN_IN), 
        .B2(keyinput_g68), .ZN(n4765) );
  OAI221_X1 U5306 ( .B1(DATAI_14_), .B2(keyinput_g17), .C1(IR_REG_13__SCAN_IN), 
        .C2(keyinput_g68), .A(n4765), .ZN(n4770) );
  AOI22_X1 U5307 ( .A1(REG0_REG_6__SCAN_IN), .A2(keyinput_g125), .B1(
        IR_REG_4__SCAN_IN), .B2(keyinput_g59), .ZN(n4766) );
  OAI221_X1 U5308 ( .B1(REG0_REG_6__SCAN_IN), .B2(keyinput_g125), .C1(
        IR_REG_4__SCAN_IN), .C2(keyinput_g59), .A(n4766), .ZN(n4769) );
  AOI22_X1 U5309 ( .A1(DATAI_3_), .A2(keyinput_g28), .B1(REG3_REG_4__SCAN_IN), 
        .B2(keyinput_g50), .ZN(n4767) );
  OAI221_X1 U5310 ( .B1(DATAI_3_), .B2(keyinput_g28), .C1(REG3_REG_4__SCAN_IN), 
        .C2(keyinput_g50), .A(n4767), .ZN(n4768) );
  NOR4_X1 U5311 ( .A1(n4771), .A2(n4770), .A3(n4769), .A4(n4768), .ZN(n4789)
         );
  AOI22_X1 U5312 ( .A1(REG0_REG_8__SCAN_IN), .A2(keyinput_g127), .B1(
        IR_REG_19__SCAN_IN), .B2(keyinput_g74), .ZN(n4772) );
  OAI221_X1 U5313 ( .B1(REG0_REG_8__SCAN_IN), .B2(keyinput_g127), .C1(
        IR_REG_19__SCAN_IN), .C2(keyinput_g74), .A(n4772), .ZN(n4779) );
  AOI22_X1 U5314 ( .A1(D_REG_18__SCAN_IN), .A2(keyinput_g105), .B1(
        D_REG_7__SCAN_IN), .B2(keyinput_g94), .ZN(n4773) );
  OAI221_X1 U5315 ( .B1(D_REG_18__SCAN_IN), .B2(keyinput_g105), .C1(
        D_REG_7__SCAN_IN), .C2(keyinput_g94), .A(n4773), .ZN(n4778) );
  AOI22_X1 U5316 ( .A1(D_REG_25__SCAN_IN), .A2(keyinput_g112), .B1(
        D_REG_28__SCAN_IN), .B2(keyinput_g115), .ZN(n4774) );
  OAI221_X1 U5317 ( .B1(D_REG_25__SCAN_IN), .B2(keyinput_g112), .C1(
        D_REG_28__SCAN_IN), .C2(keyinput_g115), .A(n4774), .ZN(n4777) );
  AOI22_X1 U5318 ( .A1(DATAI_9_), .A2(keyinput_g22), .B1(D_REG_0__SCAN_IN), 
        .B2(keyinput_g87), .ZN(n4775) );
  OAI221_X1 U5319 ( .B1(DATAI_9_), .B2(keyinput_g22), .C1(D_REG_0__SCAN_IN), 
        .C2(keyinput_g87), .A(n4775), .ZN(n4776) );
  NOR4_X1 U5320 ( .A1(n4779), .A2(n4778), .A3(n4777), .A4(n4776), .ZN(n4788)
         );
  OAI22_X1 U5321 ( .A1(DATAI_18_), .A2(keyinput_g13), .B1(keyinput_g1), .B2(
        DATAI_30_), .ZN(n4780) );
  AOI221_X1 U5322 ( .B1(DATAI_18_), .B2(keyinput_g13), .C1(DATAI_30_), .C2(
        keyinput_g1), .A(n4780), .ZN(n4786) );
  OAI22_X1 U5323 ( .A1(DATAI_25_), .A2(keyinput_g6), .B1(keyinput_g29), .B2(
        DATAI_2_), .ZN(n4781) );
  AOI221_X1 U5324 ( .B1(DATAI_25_), .B2(keyinput_g6), .C1(DATAI_2_), .C2(
        keyinput_g29), .A(n4781), .ZN(n4785) );
  OAI22_X1 U5325 ( .A1(REG3_REG_21__SCAN_IN), .A2(keyinput_g43), .B1(
        keyinput_g3), .B2(DATAI_28_), .ZN(n4782) );
  AOI221_X1 U5326 ( .B1(REG3_REG_21__SCAN_IN), .B2(keyinput_g43), .C1(
        DATAI_28_), .C2(keyinput_g3), .A(n4782), .ZN(n4784) );
  XNOR2_X1 U5327 ( .A(IR_REG_8__SCAN_IN), .B(keyinput_g63), .ZN(n4783) );
  AND4_X1 U5328 ( .A1(n4786), .A2(n4785), .A3(n4784), .A4(n4783), .ZN(n4787)
         );
  NAND3_X1 U5329 ( .A1(n4789), .A2(n4788), .A3(n4787), .ZN(n4892) );
  AOI22_X1 U5330 ( .A1(n4792), .A2(keyinput_g96), .B1(keyinput_g9), .B2(n4791), 
        .ZN(n4790) );
  OAI221_X1 U5331 ( .B1(n4792), .B2(keyinput_g96), .C1(n4791), .C2(keyinput_g9), .A(n4790), .ZN(n4802) );
  INV_X1 U5332 ( .A(DATAI_4_), .ZN(n4795) );
  AOI22_X1 U5333 ( .A1(n4795), .A2(keyinput_g27), .B1(n4794), .B2(keyinput_g14), .ZN(n4793) );
  OAI221_X1 U5334 ( .B1(n4795), .B2(keyinput_g27), .C1(n4794), .C2(
        keyinput_g14), .A(n4793), .ZN(n4801) );
  AOI22_X1 U5335 ( .A1(n5067), .A2(keyinput_g46), .B1(n2480), .B2(keyinput_g70), .ZN(n4796) );
  OAI221_X1 U5336 ( .B1(n5067), .B2(keyinput_g46), .C1(n2480), .C2(
        keyinput_g70), .A(n4796), .ZN(n4800) );
  XOR2_X1 U5337 ( .A(n3117), .B(keyinput_g52), .Z(n4798) );
  XNOR2_X1 U5338 ( .A(IR_REG_23__SCAN_IN), .B(keyinput_g78), .ZN(n4797) );
  NAND2_X1 U5339 ( .A1(n4798), .A2(n4797), .ZN(n4799) );
  NOR4_X1 U5340 ( .A1(n4802), .A2(n4801), .A3(n4800), .A4(n4799), .ZN(n4841)
         );
  AOI22_X1 U5341 ( .A1(n5047), .A2(keyinput_g93), .B1(keyinput_g123), .B2(
        n4804), .ZN(n4803) );
  OAI221_X1 U5342 ( .B1(n5047), .B2(keyinput_g93), .C1(n4804), .C2(
        keyinput_g123), .A(n4803), .ZN(n4813) );
  AOI22_X1 U5343 ( .A1(n4806), .A2(keyinput_g81), .B1(keyinput_g97), .B2(n5048), .ZN(n4805) );
  OAI221_X1 U5344 ( .B1(n4806), .B2(keyinput_g81), .C1(n5048), .C2(
        keyinput_g97), .A(n4805), .ZN(n4812) );
  AOI22_X1 U5345 ( .A1(n5068), .A2(keyinput_g0), .B1(n4967), .B2(keyinput_g5), 
        .ZN(n4807) );
  OAI221_X1 U5346 ( .B1(n5068), .B2(keyinput_g0), .C1(n4967), .C2(keyinput_g5), 
        .A(n4807), .ZN(n4811) );
  XNOR2_X1 U5347 ( .A(IR_REG_9__SCAN_IN), .B(keyinput_g64), .ZN(n4809) );
  XNOR2_X1 U5348 ( .A(DATAI_0_), .B(keyinput_g31), .ZN(n4808) );
  NAND2_X1 U5349 ( .A1(n4809), .A2(n4808), .ZN(n4810) );
  NOR4_X1 U5350 ( .A1(n4813), .A2(n4812), .A3(n4811), .A4(n4810), .ZN(n4840)
         );
  AOI22_X1 U5351 ( .A1(n4815), .A2(keyinput_g53), .B1(keyinput_g4), .B2(n4968), 
        .ZN(n4814) );
  OAI221_X1 U5352 ( .B1(n4815), .B2(keyinput_g53), .C1(n4968), .C2(keyinput_g4), .A(n4814), .ZN(n4824) );
  AOI22_X1 U5353 ( .A1(n4817), .A2(keyinput_g21), .B1(U3149), .B2(keyinput_g32), .ZN(n4816) );
  OAI221_X1 U5354 ( .B1(n4817), .B2(keyinput_g21), .C1(U3149), .C2(
        keyinput_g32), .A(n4816), .ZN(n4823) );
  XNOR2_X1 U5355 ( .A(n5044), .B(keyinput_g106), .ZN(n4822) );
  XNOR2_X1 U5356 ( .A(IR_REG_27__SCAN_IN), .B(keyinput_g82), .ZN(n4820) );
  XNOR2_X1 U5357 ( .A(IR_REG_2__SCAN_IN), .B(keyinput_g57), .ZN(n4819) );
  XNOR2_X1 U5358 ( .A(IR_REG_22__SCAN_IN), .B(keyinput_g77), .ZN(n4818) );
  NAND3_X1 U5359 ( .A1(n4820), .A2(n4819), .A3(n4818), .ZN(n4821) );
  NOR4_X1 U5360 ( .A1(n4824), .A2(n4823), .A3(n4822), .A4(n4821), .ZN(n4839)
         );
  AOI22_X1 U5361 ( .A1(n5029), .A2(keyinput_g117), .B1(n4826), .B2(
        keyinput_g61), .ZN(n4825) );
  OAI221_X1 U5362 ( .B1(n5029), .B2(keyinput_g117), .C1(n4826), .C2(
        keyinput_g61), .A(n4825), .ZN(n4831) );
  XNOR2_X1 U5363 ( .A(n4827), .B(keyinput_g101), .ZN(n4830) );
  XNOR2_X1 U5364 ( .A(n4828), .B(keyinput_g38), .ZN(n4829) );
  OR3_X1 U5365 ( .A1(n4831), .A2(n4830), .A3(n4829), .ZN(n4837) );
  INV_X1 U5366 ( .A(DATAI_6_), .ZN(n4994) );
  AOI22_X1 U5367 ( .A1(n5032), .A2(keyinput_g118), .B1(keyinput_g25), .B2(
        n4994), .ZN(n4832) );
  OAI221_X1 U5368 ( .B1(n5032), .B2(keyinput_g118), .C1(n4994), .C2(
        keyinput_g25), .A(n4832), .ZN(n4836) );
  AOI22_X1 U5369 ( .A1(n4834), .A2(keyinput_g90), .B1(keyinput_g124), .B2(
        n3252), .ZN(n4833) );
  OAI221_X1 U5370 ( .B1(n4834), .B2(keyinput_g90), .C1(n3252), .C2(
        keyinput_g124), .A(n4833), .ZN(n4835) );
  NOR3_X1 U5371 ( .A1(n4837), .A2(n4836), .A3(n4835), .ZN(n4838) );
  NAND4_X1 U5372 ( .A1(n4841), .A2(n4840), .A3(n4839), .A4(n4838), .ZN(n4891)
         );
  AOI22_X1 U5373 ( .A1(n5025), .A2(keyinput_g113), .B1(n5022), .B2(
        keyinput_g91), .ZN(n4842) );
  OAI221_X1 U5374 ( .B1(n5025), .B2(keyinput_g113), .C1(n5022), .C2(
        keyinput_g91), .A(n4842), .ZN(n4852) );
  AOI22_X1 U5375 ( .A1(n4845), .A2(keyinput_g89), .B1(n4844), .B2(keyinput_g72), .ZN(n4843) );
  OAI221_X1 U5376 ( .B1(n4845), .B2(keyinput_g89), .C1(n4844), .C2(
        keyinput_g72), .A(n4843), .ZN(n4851) );
  XNOR2_X1 U5377 ( .A(n5026), .B(keyinput_g102), .ZN(n4850) );
  XNOR2_X1 U5378 ( .A(IR_REG_21__SCAN_IN), .B(keyinput_g76), .ZN(n4848) );
  XNOR2_X1 U5379 ( .A(IR_REG_1__SCAN_IN), .B(keyinput_g56), .ZN(n4847) );
  XNOR2_X1 U5380 ( .A(IR_REG_12__SCAN_IN), .B(keyinput_g67), .ZN(n4846) );
  NAND3_X1 U5381 ( .A1(n4848), .A2(n4847), .A3(n4846), .ZN(n4849) );
  NOR4_X1 U5382 ( .A1(n4852), .A2(n4851), .A3(n4850), .A4(n4849), .ZN(n4889)
         );
  AOI22_X1 U5383 ( .A1(n5058), .A2(keyinput_g88), .B1(keyinput_g12), .B2(n4854), .ZN(n4853) );
  OAI221_X1 U5384 ( .B1(n5058), .B2(keyinput_g88), .C1(n4854), .C2(
        keyinput_g12), .A(n4853), .ZN(n4862) );
  AOI22_X1 U5385 ( .A1(n5070), .A2(keyinput_g36), .B1(keyinput_g119), .B2(
        n5006), .ZN(n4855) );
  OAI221_X1 U5386 ( .B1(n5070), .B2(keyinput_g36), .C1(n5006), .C2(
        keyinput_g119), .A(n4855), .ZN(n4861) );
  INV_X1 U5387 ( .A(REG3_REG_10__SCAN_IN), .ZN(n5071) );
  AOI22_X1 U5388 ( .A1(n5039), .A2(keyinput_g98), .B1(keyinput_g37), .B2(n5071), .ZN(n4856) );
  OAI221_X1 U5389 ( .B1(n5039), .B2(keyinput_g98), .C1(n5071), .C2(
        keyinput_g37), .A(n4856), .ZN(n4860) );
  XOR2_X1 U5390 ( .A(n4998), .B(keyinput_g47), .Z(n4858) );
  XNOR2_X1 U5391 ( .A(IR_REG_7__SCAN_IN), .B(keyinput_g62), .ZN(n4857) );
  NAND2_X1 U5392 ( .A1(n4858), .A2(n4857), .ZN(n4859) );
  NOR4_X1 U5393 ( .A1(n4862), .A2(n4861), .A3(n4860), .A4(n4859), .ZN(n4888)
         );
  INV_X1 U5394 ( .A(DATAI_13_), .ZN(n4865) );
  AOI22_X1 U5395 ( .A1(n4865), .A2(keyinput_g18), .B1(keyinput_g120), .B2(
        n4864), .ZN(n4863) );
  OAI221_X1 U5396 ( .B1(n4865), .B2(keyinput_g18), .C1(n4864), .C2(
        keyinput_g120), .A(n4863), .ZN(n4874) );
  XNOR2_X1 U5397 ( .A(n4866), .B(keyinput_g66), .ZN(n4873) );
  XNOR2_X1 U5398 ( .A(keyinput_g8), .B(n4971), .ZN(n4872) );
  XNOR2_X1 U5399 ( .A(REG3_REG_27__SCAN_IN), .B(keyinput_g34), .ZN(n4870) );
  XNOR2_X1 U5400 ( .A(IR_REG_29__SCAN_IN), .B(keyinput_g84), .ZN(n4869) );
  XNOR2_X1 U5401 ( .A(DATAI_7_), .B(keyinput_g24), .ZN(n4868) );
  XNOR2_X1 U5402 ( .A(IR_REG_24__SCAN_IN), .B(keyinput_g79), .ZN(n4867) );
  NAND4_X1 U5403 ( .A1(n4870), .A2(n4869), .A3(n4868), .A4(n4867), .ZN(n4871)
         );
  NOR4_X1 U5404 ( .A1(n4874), .A2(n4873), .A3(n4872), .A4(n4871), .ZN(n4887)
         );
  AOI22_X1 U5405 ( .A1(n5057), .A2(keyinput_g41), .B1(n2659), .B2(keyinput_g54), .ZN(n4875) );
  OAI221_X1 U5406 ( .B1(n5057), .B2(keyinput_g41), .C1(n2659), .C2(
        keyinput_g54), .A(n4875), .ZN(n4885) );
  AOI22_X1 U5407 ( .A1(n5038), .A2(keyinput_g107), .B1(n4877), .B2(
        keyinput_g95), .ZN(n4876) );
  OAI221_X1 U5408 ( .B1(n5038), .B2(keyinput_g107), .C1(n4877), .C2(
        keyinput_g95), .A(n4876), .ZN(n4884) );
  INV_X1 U5409 ( .A(DATAI_11_), .ZN(n4879) );
  AOI22_X1 U5410 ( .A1(n2708), .A2(keyinput_g48), .B1(keyinput_g20), .B2(n4879), .ZN(n4878) );
  OAI221_X1 U5411 ( .B1(n2708), .B2(keyinput_g48), .C1(n4879), .C2(
        keyinput_g20), .A(n4878), .ZN(n4883) );
  XOR2_X1 U5412 ( .A(n2613), .B(keyinput_g51), .Z(n4881) );
  XNOR2_X1 U5413 ( .A(DATAI_1_), .B(keyinput_g30), .ZN(n4880) );
  NAND2_X1 U5414 ( .A1(n4881), .A2(n4880), .ZN(n4882) );
  NOR4_X1 U5415 ( .A1(n4885), .A2(n4884), .A3(n4883), .A4(n4882), .ZN(n4886)
         );
  NAND4_X1 U5416 ( .A1(n4889), .A2(n4888), .A3(n4887), .A4(n4886), .ZN(n4890)
         );
  NOR4_X1 U5417 ( .A1(n4893), .A2(n4892), .A3(n4891), .A4(n4890), .ZN(n5094)
         );
  XOR2_X1 U5418 ( .A(DATAI_9_), .B(keyinput_f22), .Z(n4900) );
  AOI22_X1 U5419 ( .A1(REG3_REG_25__SCAN_IN), .A2(keyinput_f45), .B1(
        STATE_REG_SCAN_IN), .B2(keyinput_f32), .ZN(n4894) );
  OAI221_X1 U5420 ( .B1(REG3_REG_25__SCAN_IN), .B2(keyinput_f45), .C1(
        STATE_REG_SCAN_IN), .C2(keyinput_f32), .A(n4894), .ZN(n4899) );
  AOI22_X1 U5421 ( .A1(DATAI_2_), .A2(keyinput_f29), .B1(DATAI_28_), .B2(
        keyinput_f3), .ZN(n4895) );
  OAI221_X1 U5422 ( .B1(DATAI_2_), .B2(keyinput_f29), .C1(DATAI_28_), .C2(
        keyinput_f3), .A(n4895), .ZN(n4898) );
  AOI22_X1 U5423 ( .A1(DATAI_24_), .A2(keyinput_f7), .B1(REG3_REG_0__SCAN_IN), 
        .B2(keyinput_f52), .ZN(n4896) );
  OAI221_X1 U5424 ( .B1(DATAI_24_), .B2(keyinput_f7), .C1(REG3_REG_0__SCAN_IN), 
        .C2(keyinput_f52), .A(n4896), .ZN(n4897) );
  NOR4_X1 U5425 ( .A1(n4900), .A2(n4899), .A3(n4898), .A4(n4897), .ZN(n4928)
         );
  AOI22_X1 U5426 ( .A1(REG3_REG_19__SCAN_IN), .A2(keyinput_f39), .B1(
        REG3_REG_27__SCAN_IN), .B2(keyinput_f34), .ZN(n4901) );
  OAI221_X1 U5427 ( .B1(REG3_REG_19__SCAN_IN), .B2(keyinput_f39), .C1(
        REG3_REG_27__SCAN_IN), .C2(keyinput_f34), .A(n4901), .ZN(n4908) );
  AOI22_X1 U5428 ( .A1(REG3_REG_20__SCAN_IN), .A2(keyinput_f53), .B1(
        REG3_REG_21__SCAN_IN), .B2(keyinput_f43), .ZN(n4902) );
  OAI221_X1 U5429 ( .B1(REG3_REG_20__SCAN_IN), .B2(keyinput_f53), .C1(
        REG3_REG_21__SCAN_IN), .C2(keyinput_f43), .A(n4902), .ZN(n4907) );
  AOI22_X1 U5430 ( .A1(DATAI_30_), .A2(keyinput_f1), .B1(DATAI_22_), .B2(
        keyinput_f9), .ZN(n4903) );
  OAI221_X1 U5431 ( .B1(DATAI_30_), .B2(keyinput_f1), .C1(DATAI_22_), .C2(
        keyinput_f9), .A(n4903), .ZN(n4906) );
  AOI22_X1 U5432 ( .A1(DATAI_19_), .A2(keyinput_f12), .B1(DATAI_21_), .B2(
        keyinput_f10), .ZN(n4904) );
  OAI221_X1 U5433 ( .B1(DATAI_19_), .B2(keyinput_f12), .C1(DATAI_21_), .C2(
        keyinput_f10), .A(n4904), .ZN(n4905) );
  NOR4_X1 U5434 ( .A1(n4908), .A2(n4907), .A3(n4906), .A4(n4905), .ZN(n4927)
         );
  AOI22_X1 U5435 ( .A1(DATAI_18_), .A2(keyinput_f13), .B1(REG3_REG_7__SCAN_IN), 
        .B2(keyinput_f33), .ZN(n4909) );
  OAI221_X1 U5436 ( .B1(DATAI_18_), .B2(keyinput_f13), .C1(REG3_REG_7__SCAN_IN), .C2(keyinput_f33), .A(n4909), .ZN(n4916) );
  AOI22_X1 U5437 ( .A1(REG3_REG_13__SCAN_IN), .A2(keyinput_f54), .B1(
        REG3_REG_14__SCAN_IN), .B2(keyinput_f35), .ZN(n4910) );
  OAI221_X1 U5438 ( .B1(REG3_REG_13__SCAN_IN), .B2(keyinput_f54), .C1(
        REG3_REG_14__SCAN_IN), .C2(keyinput_f35), .A(n4910), .ZN(n4915) );
  AOI22_X1 U5439 ( .A1(DATAI_15_), .A2(keyinput_f16), .B1(D_REG_29__SCAN_IN), 
        .B2(keyinput_f116), .ZN(n4911) );
  OAI221_X1 U5440 ( .B1(DATAI_15_), .B2(keyinput_f16), .C1(D_REG_29__SCAN_IN), 
        .C2(keyinput_f116), .A(n4911), .ZN(n4914) );
  AOI22_X1 U5441 ( .A1(D_REG_23__SCAN_IN), .A2(keyinput_f110), .B1(
        D_REG_27__SCAN_IN), .B2(keyinput_f114), .ZN(n4912) );
  OAI221_X1 U5442 ( .B1(D_REG_23__SCAN_IN), .B2(keyinput_f110), .C1(
        D_REG_27__SCAN_IN), .C2(keyinput_f114), .A(n4912), .ZN(n4913) );
  NOR4_X1 U5443 ( .A1(n4916), .A2(n4915), .A3(n4914), .A4(n4913), .ZN(n4926)
         );
  AOI22_X1 U5444 ( .A1(D_REG_21__SCAN_IN), .A2(keyinput_f108), .B1(
        D_REG_22__SCAN_IN), .B2(keyinput_f109), .ZN(n4917) );
  OAI221_X1 U5445 ( .B1(D_REG_21__SCAN_IN), .B2(keyinput_f108), .C1(
        D_REG_22__SCAN_IN), .C2(keyinput_f109), .A(n4917), .ZN(n4924) );
  AOI22_X1 U5446 ( .A1(D_REG_16__SCAN_IN), .A2(keyinput_f103), .B1(
        D_REG_17__SCAN_IN), .B2(keyinput_f104), .ZN(n4918) );
  OAI221_X1 U5447 ( .B1(D_REG_16__SCAN_IN), .B2(keyinput_f103), .C1(
        D_REG_17__SCAN_IN), .C2(keyinput_f104), .A(n4918), .ZN(n4923) );
  AOI22_X1 U5448 ( .A1(IR_REG_30__SCAN_IN), .A2(keyinput_f85), .B1(
        IR_REG_16__SCAN_IN), .B2(keyinput_f71), .ZN(n4919) );
  OAI221_X1 U5449 ( .B1(IR_REG_30__SCAN_IN), .B2(keyinput_f85), .C1(
        IR_REG_16__SCAN_IN), .C2(keyinput_f71), .A(n4919), .ZN(n4922) );
  AOI22_X1 U5450 ( .A1(DATAI_16_), .A2(keyinput_f15), .B1(IR_REG_15__SCAN_IN), 
        .B2(keyinput_f70), .ZN(n4920) );
  OAI221_X1 U5451 ( .B1(DATAI_16_), .B2(keyinput_f15), .C1(IR_REG_15__SCAN_IN), 
        .C2(keyinput_f70), .A(n4920), .ZN(n4921) );
  NOR4_X1 U5452 ( .A1(n4924), .A2(n4923), .A3(n4922), .A4(n4921), .ZN(n4925)
         );
  NAND4_X1 U5453 ( .A1(n4928), .A2(n4927), .A3(n4926), .A4(n4925), .ZN(n5087)
         );
  AOI22_X1 U5454 ( .A1(DATAI_8_), .A2(keyinput_f23), .B1(DATAI_12_), .B2(
        keyinput_f19), .ZN(n4929) );
  OAI221_X1 U5455 ( .B1(DATAI_8_), .B2(keyinput_f23), .C1(DATAI_12_), .C2(
        keyinput_f19), .A(n4929), .ZN(n4936) );
  AOI22_X1 U5456 ( .A1(REG0_REG_3__SCAN_IN), .A2(keyinput_f122), .B1(DATAI_5_), 
        .B2(keyinput_f26), .ZN(n4930) );
  OAI221_X1 U5457 ( .B1(REG0_REG_3__SCAN_IN), .B2(keyinput_f122), .C1(DATAI_5_), .C2(keyinput_f26), .A(n4930), .ZN(n4935) );
  AOI22_X1 U5458 ( .A1(IR_REG_28__SCAN_IN), .A2(keyinput_f83), .B1(
        IR_REG_12__SCAN_IN), .B2(keyinput_f67), .ZN(n4931) );
  OAI221_X1 U5459 ( .B1(IR_REG_28__SCAN_IN), .B2(keyinput_f83), .C1(
        IR_REG_12__SCAN_IN), .C2(keyinput_f67), .A(n4931), .ZN(n4934) );
  AOI22_X1 U5460 ( .A1(DATAI_10_), .A2(keyinput_f21), .B1(IR_REG_10__SCAN_IN), 
        .B2(keyinput_f65), .ZN(n4932) );
  OAI221_X1 U5461 ( .B1(DATAI_10_), .B2(keyinput_f21), .C1(IR_REG_10__SCAN_IN), 
        .C2(keyinput_f65), .A(n4932), .ZN(n4933) );
  NOR4_X1 U5462 ( .A1(n4936), .A2(n4935), .A3(n4934), .A4(n4933), .ZN(n4965)
         );
  AOI22_X1 U5463 ( .A1(IR_REG_6__SCAN_IN), .A2(keyinput_f61), .B1(
        IR_REG_7__SCAN_IN), .B2(keyinput_f62), .ZN(n4937) );
  OAI221_X1 U5464 ( .B1(IR_REG_6__SCAN_IN), .B2(keyinput_f61), .C1(
        IR_REG_7__SCAN_IN), .C2(keyinput_f62), .A(n4937), .ZN(n4944) );
  AOI22_X1 U5465 ( .A1(DATAI_4_), .A2(keyinput_f27), .B1(REG0_REG_5__SCAN_IN), 
        .B2(keyinput_f124), .ZN(n4938) );
  OAI221_X1 U5466 ( .B1(DATAI_4_), .B2(keyinput_f27), .C1(REG0_REG_5__SCAN_IN), 
        .C2(keyinput_f124), .A(n4938), .ZN(n4943) );
  AOI22_X1 U5467 ( .A1(IR_REG_3__SCAN_IN), .A2(keyinput_f58), .B1(
        IR_REG_4__SCAN_IN), .B2(keyinput_f59), .ZN(n4939) );
  OAI221_X1 U5468 ( .B1(IR_REG_3__SCAN_IN), .B2(keyinput_f58), .C1(
        IR_REG_4__SCAN_IN), .C2(keyinput_f59), .A(n4939), .ZN(n4942) );
  AOI22_X1 U5469 ( .A1(REG0_REG_4__SCAN_IN), .A2(keyinput_f123), .B1(
        REG0_REG_1__SCAN_IN), .B2(keyinput_f120), .ZN(n4940) );
  OAI221_X1 U5470 ( .B1(REG0_REG_4__SCAN_IN), .B2(keyinput_f123), .C1(
        REG0_REG_1__SCAN_IN), .C2(keyinput_f120), .A(n4940), .ZN(n4941) );
  NOR4_X1 U5471 ( .A1(n4944), .A2(n4943), .A3(n4942), .A4(n4941), .ZN(n4964)
         );
  AOI22_X1 U5472 ( .A1(DATAI_1_), .A2(keyinput_f30), .B1(IR_REG_1__SCAN_IN), 
        .B2(keyinput_f56), .ZN(n4945) );
  OAI221_X1 U5473 ( .B1(DATAI_1_), .B2(keyinput_f30), .C1(IR_REG_1__SCAN_IN), 
        .C2(keyinput_f56), .A(n4945), .ZN(n4952) );
  AOI22_X1 U5474 ( .A1(REG3_REG_9__SCAN_IN), .A2(keyinput_f51), .B1(
        IR_REG_9__SCAN_IN), .B2(keyinput_f64), .ZN(n4946) );
  OAI221_X1 U5475 ( .B1(REG3_REG_9__SCAN_IN), .B2(keyinput_f51), .C1(
        IR_REG_9__SCAN_IN), .C2(keyinput_f64), .A(n4946), .ZN(n4951) );
  AOI22_X1 U5476 ( .A1(DATAI_11_), .A2(keyinput_f20), .B1(IR_REG_19__SCAN_IN), 
        .B2(keyinput_f74), .ZN(n4947) );
  OAI221_X1 U5477 ( .B1(DATAI_11_), .B2(keyinput_f20), .C1(IR_REG_19__SCAN_IN), 
        .C2(keyinput_f74), .A(n4947), .ZN(n4950) );
  AOI22_X1 U5478 ( .A1(D_REG_2__SCAN_IN), .A2(keyinput_f89), .B1(
        IR_REG_20__SCAN_IN), .B2(keyinput_f75), .ZN(n4948) );
  OAI221_X1 U5479 ( .B1(D_REG_2__SCAN_IN), .B2(keyinput_f89), .C1(
        IR_REG_20__SCAN_IN), .C2(keyinput_f75), .A(n4948), .ZN(n4949) );
  NOR4_X1 U5480 ( .A1(n4952), .A2(n4951), .A3(n4950), .A4(n4949), .ZN(n4963)
         );
  AOI22_X1 U5481 ( .A1(D_REG_14__SCAN_IN), .A2(keyinput_f101), .B1(
        D_REG_9__SCAN_IN), .B2(keyinput_f96), .ZN(n4953) );
  OAI221_X1 U5482 ( .B1(D_REG_14__SCAN_IN), .B2(keyinput_f101), .C1(
        D_REG_9__SCAN_IN), .C2(keyinput_f96), .A(n4953), .ZN(n4961) );
  AOI22_X1 U5483 ( .A1(D_REG_24__SCAN_IN), .A2(keyinput_f111), .B1(
        D_REG_3__SCAN_IN), .B2(keyinput_f90), .ZN(n4954) );
  OAI221_X1 U5484 ( .B1(D_REG_24__SCAN_IN), .B2(keyinput_f111), .C1(
        D_REG_3__SCAN_IN), .C2(keyinput_f90), .A(n4954), .ZN(n4960) );
  AOI22_X1 U5485 ( .A1(D_REG_8__SCAN_IN), .A2(keyinput_f95), .B1(
        IR_REG_26__SCAN_IN), .B2(keyinput_f81), .ZN(n4955) );
  OAI221_X1 U5486 ( .B1(D_REG_8__SCAN_IN), .B2(keyinput_f95), .C1(
        IR_REG_26__SCAN_IN), .C2(keyinput_f81), .A(n4955), .ZN(n4959) );
  INV_X1 U5487 ( .A(DATAI_25_), .ZN(n4957) );
  AOI22_X1 U5488 ( .A1(DATAI_13_), .A2(keyinput_f18), .B1(n4957), .B2(
        keyinput_f6), .ZN(n4956) );
  OAI221_X1 U5489 ( .B1(DATAI_13_), .B2(keyinput_f18), .C1(n4957), .C2(
        keyinput_f6), .A(n4956), .ZN(n4958) );
  NOR4_X1 U5490 ( .A1(n4961), .A2(n4960), .A3(n4959), .A4(n4958), .ZN(n4962)
         );
  NAND4_X1 U5491 ( .A1(n4965), .A2(n4964), .A3(n4963), .A4(n4962), .ZN(n5086)
         );
  AOI22_X1 U5492 ( .A1(n4968), .A2(keyinput_f4), .B1(keyinput_f5), .B2(n4967), 
        .ZN(n4966) );
  OAI221_X1 U5493 ( .B1(n4968), .B2(keyinput_f4), .C1(n4967), .C2(keyinput_f5), 
        .A(n4966), .ZN(n4979) );
  AOI22_X1 U5494 ( .A1(n4971), .A2(keyinput_f8), .B1(keyinput_f11), .B2(n4970), 
        .ZN(n4969) );
  OAI221_X1 U5495 ( .B1(n4971), .B2(keyinput_f8), .C1(n4970), .C2(keyinput_f11), .A(n4969), .ZN(n4978) );
  AOI22_X1 U5496 ( .A1(n3685), .A2(keyinput_f40), .B1(keyinput_f49), .B2(n4973), .ZN(n4972) );
  OAI221_X1 U5497 ( .B1(n3685), .B2(keyinput_f40), .C1(n4973), .C2(
        keyinput_f49), .A(n4972), .ZN(n4977) );
  XNOR2_X1 U5498 ( .A(REG3_REG_3__SCAN_IN), .B(keyinput_f38), .ZN(n4975) );
  XNOR2_X1 U5499 ( .A(DATAI_17_), .B(keyinput_f14), .ZN(n4974) );
  NAND2_X1 U5500 ( .A1(n4975), .A2(n4974), .ZN(n4976) );
  NOR4_X1 U5501 ( .A1(n4979), .A2(n4978), .A3(n4977), .A4(n4976), .ZN(n5020)
         );
  AOI22_X1 U5502 ( .A1(n4982), .A2(keyinput_f69), .B1(keyinput_f17), .B2(n4981), .ZN(n4980) );
  OAI221_X1 U5503 ( .B1(n4982), .B2(keyinput_f69), .C1(n4981), .C2(
        keyinput_f17), .A(n4980), .ZN(n4991) );
  XNOR2_X1 U5504 ( .A(n4983), .B(keyinput_f73), .ZN(n4990) );
  XNOR2_X1 U5505 ( .A(keyinput_f42), .B(n3157), .ZN(n4989) );
  XNOR2_X1 U5506 ( .A(IR_REG_27__SCAN_IN), .B(keyinput_f82), .ZN(n4987) );
  XNOR2_X1 U5507 ( .A(IR_REG_0__SCAN_IN), .B(keyinput_f55), .ZN(n4986) );
  XNOR2_X1 U5508 ( .A(IR_REG_17__SCAN_IN), .B(keyinput_f72), .ZN(n4985) );
  XNOR2_X1 U5509 ( .A(IR_REG_31__SCAN_IN), .B(keyinput_f86), .ZN(n4984) );
  NAND4_X1 U5510 ( .A1(n4987), .A2(n4986), .A3(n4985), .A4(n4984), .ZN(n4988)
         );
  NOR4_X1 U5511 ( .A1(n4991), .A2(n4990), .A3(n4989), .A4(n4988), .ZN(n5019)
         );
  AOI22_X1 U5512 ( .A1(n4994), .A2(keyinput_f25), .B1(keyinput_f125), .B2(
        n4993), .ZN(n4992) );
  OAI221_X1 U5513 ( .B1(n4994), .B2(keyinput_f25), .C1(n4993), .C2(
        keyinput_f125), .A(n4992), .ZN(n5005) );
  INV_X1 U5514 ( .A(DATAI_7_), .ZN(n4997) );
  AOI22_X1 U5515 ( .A1(n4997), .A2(keyinput_f24), .B1(n4996), .B2(
        keyinput_f126), .ZN(n4995) );
  OAI221_X1 U5516 ( .B1(n4997), .B2(keyinput_f24), .C1(n4996), .C2(
        keyinput_f126), .A(n4995), .ZN(n5004) );
  XOR2_X1 U5517 ( .A(n4998), .B(keyinput_f47), .Z(n5002) );
  XNOR2_X1 U5518 ( .A(IR_REG_11__SCAN_IN), .B(keyinput_f66), .ZN(n5001) );
  XNOR2_X1 U5519 ( .A(IR_REG_13__SCAN_IN), .B(keyinput_f68), .ZN(n5000) );
  XNOR2_X1 U5520 ( .A(IR_REG_5__SCAN_IN), .B(keyinput_f60), .ZN(n4999) );
  NAND4_X1 U5521 ( .A1(n5002), .A2(n5001), .A3(n5000), .A4(n4999), .ZN(n5003)
         );
  NOR3_X1 U5522 ( .A1(n5005), .A2(n5004), .A3(n5003), .ZN(n5018) );
  XOR2_X1 U5523 ( .A(n5006), .B(keyinput_f119), .Z(n5010) );
  XNOR2_X1 U5524 ( .A(keyinput_f127), .B(REG0_REG_8__SCAN_IN), .ZN(n5009) );
  XNOR2_X1 U5525 ( .A(IR_REG_21__SCAN_IN), .B(keyinput_f76), .ZN(n5008) );
  XNOR2_X1 U5526 ( .A(IR_REG_8__SCAN_IN), .B(keyinput_f63), .ZN(n5007) );
  NAND4_X1 U5527 ( .A1(n5010), .A2(n5009), .A3(n5008), .A4(n5007), .ZN(n5016)
         );
  XNOR2_X1 U5528 ( .A(REG3_REG_4__SCAN_IN), .B(keyinput_f50), .ZN(n5014) );
  XNOR2_X1 U5529 ( .A(DATAI_0_), .B(keyinput_f31), .ZN(n5013) );
  XNOR2_X1 U5530 ( .A(DATAI_3_), .B(keyinput_f28), .ZN(n5012) );
  XNOR2_X1 U5531 ( .A(IR_REG_2__SCAN_IN), .B(keyinput_f57), .ZN(n5011) );
  NAND4_X1 U5532 ( .A1(n5014), .A2(n5013), .A3(n5012), .A4(n5011), .ZN(n5015)
         );
  NOR2_X1 U5533 ( .A1(n5016), .A2(n5015), .ZN(n5017) );
  NAND4_X1 U5534 ( .A1(n5020), .A2(n5019), .A3(n5018), .A4(n5017), .ZN(n5085)
         );
  AOI22_X1 U5535 ( .A1(n5023), .A2(keyinput_f77), .B1(keyinput_f91), .B2(n5022), .ZN(n5021) );
  OAI221_X1 U5536 ( .B1(n5023), .B2(keyinput_f77), .C1(n5022), .C2(
        keyinput_f91), .A(n5021), .ZN(n5036) );
  AOI22_X1 U5537 ( .A1(n5026), .A2(keyinput_f102), .B1(keyinput_f113), .B2(
        n5025), .ZN(n5024) );
  OAI221_X1 U5538 ( .B1(n5026), .B2(keyinput_f102), .C1(n5025), .C2(
        keyinput_f113), .A(n5024), .ZN(n5035) );
  AOI22_X1 U5539 ( .A1(n5029), .A2(keyinput_f117), .B1(keyinput_f100), .B2(
        n5028), .ZN(n5027) );
  OAI221_X1 U5540 ( .B1(n5029), .B2(keyinput_f117), .C1(n5028), .C2(
        keyinput_f100), .A(n5027), .ZN(n5034) );
  AOI22_X1 U5541 ( .A1(n5032), .A2(keyinput_f118), .B1(keyinput_f99), .B2(
        n5031), .ZN(n5030) );
  OAI221_X1 U5542 ( .B1(n5032), .B2(keyinput_f118), .C1(n5031), .C2(
        keyinput_f99), .A(n5030), .ZN(n5033) );
  NOR4_X1 U5543 ( .A1(n5036), .A2(n5035), .A3(n5034), .A4(n5033), .ZN(n5083)
         );
  AOI22_X1 U5544 ( .A1(n5039), .A2(keyinput_f98), .B1(keyinput_f107), .B2(
        n5038), .ZN(n5037) );
  OAI221_X1 U5545 ( .B1(n5039), .B2(keyinput_f98), .C1(n5038), .C2(
        keyinput_f107), .A(n5037), .ZN(n5052) );
  AOI22_X1 U5546 ( .A1(n5042), .A2(keyinput_f94), .B1(keyinput_f105), .B2(
        n5041), .ZN(n5040) );
  OAI221_X1 U5547 ( .B1(n5042), .B2(keyinput_f94), .C1(n5041), .C2(
        keyinput_f105), .A(n5040), .ZN(n5051) );
  AOI22_X1 U5548 ( .A1(n5045), .A2(keyinput_f112), .B1(keyinput_f106), .B2(
        n5044), .ZN(n5043) );
  OAI221_X1 U5549 ( .B1(n5045), .B2(keyinput_f112), .C1(n5044), .C2(
        keyinput_f106), .A(n5043), .ZN(n5050) );
  AOI22_X1 U5550 ( .A1(n5048), .A2(keyinput_f97), .B1(keyinput_f93), .B2(n5047), .ZN(n5046) );
  OAI221_X1 U5551 ( .B1(n5048), .B2(keyinput_f97), .C1(n5047), .C2(
        keyinput_f93), .A(n5046), .ZN(n5049) );
  NOR4_X1 U5552 ( .A1(n5052), .A2(n5051), .A3(n5050), .A4(n5049), .ZN(n5082)
         );
  AOI22_X1 U5553 ( .A1(n5054), .A2(keyinput_f115), .B1(keyinput_f48), .B2(
        n2708), .ZN(n5053) );
  OAI221_X1 U5554 ( .B1(n5054), .B2(keyinput_f115), .C1(n2708), .C2(
        keyinput_f48), .A(n5053), .ZN(n5065) );
  INV_X1 U5555 ( .A(DATAI_29_), .ZN(n5056) );
  AOI22_X1 U5556 ( .A1(n5057), .A2(keyinput_f41), .B1(keyinput_f2), .B2(n5056), 
        .ZN(n5055) );
  OAI221_X1 U5557 ( .B1(n5057), .B2(keyinput_f41), .C1(n5056), .C2(keyinput_f2), .A(n5055), .ZN(n5064) );
  XNOR2_X1 U5558 ( .A(n5058), .B(keyinput_f88), .ZN(n5063) );
  XNOR2_X1 U5559 ( .A(IR_REG_24__SCAN_IN), .B(keyinput_f79), .ZN(n5061) );
  XNOR2_X1 U5560 ( .A(REG3_REG_12__SCAN_IN), .B(keyinput_f44), .ZN(n5060) );
  XNOR2_X1 U5561 ( .A(IR_REG_29__SCAN_IN), .B(keyinput_f84), .ZN(n5059) );
  NAND3_X1 U5562 ( .A1(n5061), .A2(n5060), .A3(n5059), .ZN(n5062) );
  NOR4_X1 U5563 ( .A1(n5065), .A2(n5064), .A3(n5063), .A4(n5062), .ZN(n5081)
         );
  AOI22_X1 U5564 ( .A1(n5068), .A2(keyinput_f0), .B1(n5067), .B2(keyinput_f46), 
        .ZN(n5066) );
  OAI221_X1 U5565 ( .B1(n5068), .B2(keyinput_f0), .C1(n5067), .C2(keyinput_f46), .A(n5066), .ZN(n5079) );
  AOI22_X1 U5566 ( .A1(n5071), .A2(keyinput_f37), .B1(n5070), .B2(keyinput_f36), .ZN(n5069) );
  OAI221_X1 U5567 ( .B1(n5071), .B2(keyinput_f37), .C1(n5070), .C2(
        keyinput_f36), .A(n5069), .ZN(n5078) );
  XOR2_X1 U5568 ( .A(n5072), .B(keyinput_f121), .Z(n5076) );
  XNOR2_X1 U5569 ( .A(IR_REG_25__SCAN_IN), .B(keyinput_f80), .ZN(n5075) );
  XNOR2_X1 U5570 ( .A(IR_REG_23__SCAN_IN), .B(keyinput_f78), .ZN(n5074) );
  XNOR2_X1 U5571 ( .A(D_REG_0__SCAN_IN), .B(keyinput_f87), .ZN(n5073) );
  NAND4_X1 U5572 ( .A1(n5076), .A2(n5075), .A3(n5074), .A4(n5073), .ZN(n5077)
         );
  NOR3_X1 U5573 ( .A1(n5079), .A2(n5078), .A3(n5077), .ZN(n5080) );
  NAND4_X1 U5574 ( .A1(n5083), .A2(n5082), .A3(n5081), .A4(n5080), .ZN(n5084)
         );
  OR4_X1 U5575 ( .A1(n5087), .A2(n5086), .A3(n5085), .A4(n5084), .ZN(n5089) );
  AOI21_X1 U5576 ( .B1(keyinput_f92), .B2(n5089), .A(keyinput_g92), .ZN(n5091)
         );
  INV_X1 U5577 ( .A(keyinput_f92), .ZN(n5088) );
  AOI21_X1 U5578 ( .B1(n5089), .B2(n5088), .A(n5092), .ZN(n5090) );
  AOI22_X1 U5579 ( .A1(n5092), .A2(n5091), .B1(keyinput_g92), .B2(n5090), .ZN(
        n5093) );
  AOI21_X1 U5580 ( .B1(n5095), .B2(n5094), .A(n5093), .ZN(n5097) );
  AOI22_X1 U5581 ( .A1(STATE_REG_SCAN_IN), .A2(IR_REG_0__SCAN_IN), .B1(
        DATAI_0_), .B2(U3149), .ZN(n5096) );
  XNOR2_X1 U5582 ( .A(n5097), .B(n5096), .ZN(U3352) );
  CLKBUF_X1 U2475 ( .A(n3675), .Z(n2232) );
endmodule

