

module b21_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, 
        ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, 
        ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, 
        ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, 
        ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, 
        P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, 
        P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, 
        P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, 
        P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, 
        P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, 
        P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, 
        P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, 
        P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, 
        P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, 
        P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, 
        P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, 
        P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, 
        P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, 
        P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, 
        P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, 
        P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, 
        P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, 
        P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, 
        P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, 
        P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, 
        P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, 
        P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, 
        P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, 
        P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, 
        P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, 
        P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, 
        P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, 
        P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, 
        P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, 
        P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, 
        P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, 
        P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, 
        P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, 
        P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, 
        P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, 
        P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, 
        P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, 
        P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, 
        P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, 
        P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, 
        P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, 
        P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, 
        P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, 
        P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3152, P2_U3151, P2_U3966, keyinput127, keyinput126, 
        keyinput125, keyinput124, keyinput123, keyinput122, keyinput121, 
        keyinput120, keyinput119, keyinput118, keyinput117, keyinput116, 
        keyinput115, keyinput114, keyinput113, keyinput112, keyinput111, 
        keyinput110, keyinput109, keyinput108, keyinput107, keyinput106, 
        keyinput105, keyinput104, keyinput103, keyinput102, keyinput101, 
        keyinput100, keyinput99, keyinput98, keyinput97, keyinput96, 
        keyinput95, keyinput94, keyinput93, keyinput92, keyinput91, keyinput90, 
        keyinput89, keyinput88, keyinput87, keyinput86, keyinput85, keyinput84, 
        keyinput83, keyinput82, keyinput81, keyinput80, keyinput79, keyinput78, 
        keyinput77, keyinput76, keyinput75, keyinput74, keyinput73, keyinput72, 
        keyinput71, keyinput70, keyinput69, keyinput68, keyinput67, keyinput66, 
        keyinput65, keyinput64, keyinput63, keyinput62, keyinput61, keyinput60, 
        keyinput59, keyinput58, keyinput57, keyinput56, keyinput55, keyinput54, 
        keyinput53, keyinput52, keyinput51, keyinput50, keyinput49, keyinput48, 
        keyinput47, keyinput46, keyinput45, keyinput44, keyinput43, keyinput42, 
        keyinput41, keyinput40, keyinput39, keyinput38, keyinput37, keyinput36, 
        keyinput35, keyinput34, keyinput33, keyinput32, keyinput31, keyinput30, 
        keyinput29, keyinput28, keyinput27, keyinput26, keyinput25, keyinput24, 
        keyinput23, keyinput22, keyinput21, keyinput20, keyinput19, keyinput18, 
        keyinput17, keyinput16, keyinput15, keyinput14, keyinput13, keyinput12, 
        keyinput11, keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, 
        keyinput5, keyinput4, keyinput3, keyinput2, keyinput1, keyinput0 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput127, keyinput126, keyinput125,
         keyinput124, keyinput123, keyinput122, keyinput121, keyinput120,
         keyinput119, keyinput118, keyinput117, keyinput116, keyinput115,
         keyinput114, keyinput113, keyinput112, keyinput111, keyinput110,
         keyinput109, keyinput108, keyinput107, keyinput106, keyinput105,
         keyinput104, keyinput103, keyinput102, keyinput101, keyinput100,
         keyinput99, keyinput98, keyinput97, keyinput96, keyinput95,
         keyinput94, keyinput93, keyinput92, keyinput91, keyinput90,
         keyinput89, keyinput88, keyinput87, keyinput86, keyinput85,
         keyinput84, keyinput83, keyinput82, keyinput81, keyinput80,
         keyinput79, keyinput78, keyinput77, keyinput76, keyinput75,
         keyinput74, keyinput73, keyinput72, keyinput71, keyinput70,
         keyinput69, keyinput68, keyinput67, keyinput66, keyinput65,
         keyinput64, keyinput63, keyinput62, keyinput61, keyinput60,
         keyinput59, keyinput58, keyinput57, keyinput56, keyinput55,
         keyinput54, keyinput53, keyinput52, keyinput51, keyinput50,
         keyinput49, keyinput48, keyinput47, keyinput46, keyinput45,
         keyinput44, keyinput43, keyinput42, keyinput41, keyinput40,
         keyinput39, keyinput38, keyinput37, keyinput36, keyinput35,
         keyinput34, keyinput33, keyinput32, keyinput31, keyinput30,
         keyinput29, keyinput28, keyinput27, keyinput26, keyinput25,
         keyinput24, keyinput23, keyinput22, keyinput21, keyinput20,
         keyinput19, keyinput18, keyinput17, keyinput16, keyinput15,
         keyinput14, keyinput13, keyinput12, keyinput11, keyinput10, keyinput9,
         keyinput8, keyinput7, keyinput6, keyinput5, keyinput4, keyinput3,
         keyinput2, keyinput1, keyinput0;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4366, n4367, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377,
         n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387,
         n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397,
         n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407,
         n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417,
         n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427,
         n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437,
         n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447,
         n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457,
         n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467,
         n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477,
         n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487,
         n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497,
         n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507,
         n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517,
         n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527,
         n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537,
         n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547,
         n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557,
         n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567,
         n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577,
         n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587,
         n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597,
         n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607,
         n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617,
         n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627,
         n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637,
         n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647,
         n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657,
         n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667,
         n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677,
         n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687,
         n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697,
         n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707,
         n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717,
         n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727,
         n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737,
         n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747,
         n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757,
         n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767,
         n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777,
         n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787,
         n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797,
         n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807,
         n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817,
         n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827,
         n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837,
         n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847,
         n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857,
         n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867,
         n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877,
         n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887,
         n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897,
         n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907,
         n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917,
         n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927,
         n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937,
         n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947,
         n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957,
         n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967,
         n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977,
         n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987,
         n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997,
         n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007,
         n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017,
         n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027,
         n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037,
         n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047,
         n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057,
         n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067,
         n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077,
         n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087,
         n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097,
         n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107,
         n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117,
         n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127,
         n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137,
         n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147,
         n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157,
         n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167,
         n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177,
         n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187,
         n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197,
         n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207,
         n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217,
         n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227,
         n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237,
         n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247,
         n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257,
         n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267,
         n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277,
         n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287,
         n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297,
         n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307,
         n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317,
         n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327,
         n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337,
         n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347,
         n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357,
         n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367,
         n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377,
         n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387,
         n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397,
         n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407,
         n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417,
         n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427,
         n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437,
         n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447,
         n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457,
         n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467,
         n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477,
         n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487,
         n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497,
         n5498, n5499, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508,
         n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518,
         n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528,
         n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538,
         n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548,
         n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558,
         n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568,
         n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578,
         n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588,
         n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598,
         n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608,
         n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618,
         n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628,
         n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638,
         n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648,
         n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658,
         n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668,
         n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678,
         n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688,
         n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698,
         n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708,
         n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718,
         n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728,
         n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738,
         n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748,
         n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758,
         n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768,
         n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778,
         n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788,
         n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798,
         n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808,
         n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818,
         n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828,
         n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838,
         n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848,
         n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858,
         n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868,
         n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878,
         n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888,
         n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898,
         n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908,
         n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918,
         n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928,
         n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938,
         n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948,
         n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958,
         n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968,
         n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978,
         n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988,
         n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998,
         n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008,
         n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018,
         n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028,
         n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038,
         n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048,
         n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058,
         n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068,
         n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078,
         n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088,
         n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098,
         n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108,
         n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118,
         n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128,
         n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138,
         n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148,
         n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158,
         n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168,
         n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178,
         n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188,
         n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198,
         n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208,
         n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218,
         n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228,
         n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238,
         n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248,
         n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258,
         n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268,
         n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278,
         n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288,
         n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298,
         n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308,
         n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318,
         n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328,
         n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338,
         n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348,
         n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358,
         n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368,
         n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378,
         n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388,
         n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398,
         n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408,
         n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418,
         n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428,
         n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438,
         n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448,
         n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458,
         n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468,
         n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478,
         n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488,
         n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498,
         n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508,
         n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518,
         n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528,
         n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538,
         n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548,
         n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558,
         n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568,
         n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578,
         n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588,
         n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598,
         n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608,
         n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618,
         n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628,
         n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638,
         n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648,
         n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658,
         n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668,
         n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678,
         n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688,
         n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698,
         n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708,
         n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718,
         n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728,
         n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738,
         n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748,
         n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758,
         n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768,
         n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778,
         n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788,
         n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798,
         n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808,
         n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818,
         n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828,
         n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838,
         n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848,
         n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858,
         n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868,
         n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878,
         n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888,
         n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898,
         n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908,
         n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918,
         n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928,
         n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938,
         n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948,
         n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958,
         n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968,
         n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978,
         n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988,
         n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998,
         n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008,
         n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018,
         n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028,
         n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038,
         n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048,
         n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058,
         n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068,
         n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078,
         n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088,
         n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098,
         n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108,
         n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118,
         n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128,
         n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138,
         n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148,
         n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158,
         n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168,
         n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178,
         n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188,
         n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198,
         n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208,
         n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218,
         n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228,
         n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238,
         n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248,
         n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258,
         n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268,
         n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278,
         n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288,
         n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298,
         n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308,
         n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318,
         n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328,
         n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338,
         n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348,
         n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358,
         n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368,
         n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378,
         n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388,
         n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398,
         n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408,
         n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418,
         n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428,
         n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438,
         n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448,
         n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458,
         n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468,
         n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478,
         n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488,
         n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498,
         n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508,
         n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518,
         n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528,
         n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538,
         n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548,
         n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558,
         n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568,
         n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578,
         n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588,
         n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598,
         n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608,
         n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618,
         n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628,
         n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638,
         n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648,
         n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658,
         n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668,
         n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678,
         n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688,
         n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698,
         n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708,
         n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718,
         n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728,
         n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738,
         n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748,
         n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758,
         n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768,
         n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778,
         n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788,
         n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798,
         n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808,
         n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818,
         n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828,
         n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838,
         n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848,
         n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858,
         n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868,
         n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878,
         n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888,
         n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898,
         n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908,
         n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918,
         n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928,
         n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938,
         n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948,
         n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958,
         n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968,
         n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978,
         n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988,
         n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998,
         n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008,
         n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018,
         n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028,
         n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038,
         n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048,
         n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058,
         n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068,
         n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078,
         n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088,
         n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098,
         n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108,
         n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118,
         n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128,
         n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138,
         n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148,
         n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158,
         n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168,
         n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178,
         n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188,
         n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198,
         n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208,
         n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218,
         n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228,
         n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238,
         n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248,
         n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258,
         n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268,
         n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278,
         n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288,
         n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298,
         n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308,
         n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318,
         n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328,
         n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338,
         n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348,
         n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358,
         n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368,
         n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378,
         n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388,
         n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398,
         n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408,
         n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418,
         n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428,
         n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438,
         n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448,
         n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458,
         n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468,
         n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478,
         n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488,
         n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498,
         n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508,
         n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518,
         n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528,
         n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538,
         n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548,
         n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558,
         n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568,
         n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578,
         n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588,
         n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598,
         n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608,
         n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618,
         n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628,
         n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638,
         n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648,
         n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658,
         n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668,
         n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678,
         n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688,
         n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698,
         n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708,
         n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718,
         n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728,
         n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738,
         n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748,
         n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758,
         n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768,
         n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778,
         n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788,
         n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798,
         n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808,
         n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818,
         n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828,
         n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838,
         n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848,
         n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858,
         n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868,
         n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878,
         n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888,
         n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898,
         n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908,
         n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918,
         n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928,
         n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938,
         n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948,
         n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958,
         n8959, n8960, n8961, n8962, n8963, n8964, n8966, n8967, n8968, n8969,
         n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979,
         n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989,
         n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999,
         n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009,
         n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019,
         n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029,
         n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039,
         n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049,
         n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059,
         n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069,
         n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079,
         n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089,
         n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099,
         n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109,
         n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119,
         n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129,
         n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139,
         n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149,
         n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159,
         n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169,
         n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179,
         n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189,
         n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199,
         n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209,
         n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219,
         n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229,
         n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239,
         n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249,
         n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259,
         n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269,
         n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279,
         n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289,
         n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299,
         n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309,
         n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319,
         n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329,
         n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339,
         n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349,
         n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359,
         n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369,
         n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379,
         n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389,
         n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399,
         n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409,
         n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419,
         n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429,
         n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439,
         n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449,
         n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459,
         n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469,
         n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479,
         n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489,
         n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499,
         n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509,
         n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519,
         n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529,
         n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539,
         n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549,
         n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559,
         n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569,
         n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579,
         n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589,
         n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599,
         n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609,
         n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619,
         n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629,
         n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639,
         n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649,
         n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659,
         n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669,
         n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679,
         n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689,
         n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699,
         n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709,
         n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719,
         n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729,
         n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739,
         n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749,
         n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759,
         n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769,
         n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779,
         n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789,
         n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799,
         n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809,
         n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9819, n9820,
         n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830,
         n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840,
         n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850,
         n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860,
         n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870,
         n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880,
         n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890,
         n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900,
         n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910,
         n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920,
         n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930,
         n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940,
         n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950,
         n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960,
         n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970,
         n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980,
         n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990,
         n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273;

  NAND2_X1 U4871 ( .A1(n4901), .A2(n4900), .ZN(n8722) );
  OAI21_X1 U4872 ( .B1(n7872), .B2(P2_REG2_REG_14__SCAN_IN), .A(n7869), .ZN(
        n8086) );
  OR2_X1 U4873 ( .A1(n6917), .A2(n4647), .ZN(n4646) );
  AND2_X1 U4874 ( .A1(n4649), .A2(n4648), .ZN(n6917) );
  OAI21_X1 U4875 ( .B1(n5600), .B2(n5599), .A(n5598), .ZN(n5607) );
  AOI21_X1 U4876 ( .B1(P2_REG2_REG_4__SCAN_IN), .B2(n6559), .A(n6573), .ZN(
        n6549) );
  AOI21_X1 U4877 ( .B1(P2_REG2_REG_2__SCAN_IN), .B2(n6556), .A(n9477), .ZN(
        n6785) );
  AOI21_X1 U4878 ( .B1(P2_REG2_REG_1__SCAN_IN), .B2(n6554), .A(n9462), .ZN(
        n9478) );
  INV_X1 U4879 ( .A(n5239), .ZN(n5447) );
  NOR2_X1 U4880 ( .A1(n5147), .A2(n5146), .ZN(n4920) );
  AND2_X1 U4881 ( .A1(n4642), .A2(n4644), .ZN(n8234) );
  INV_X1 U4882 ( .A(n4392), .ZN(n6169) );
  AND3_X1 U4883 ( .A1(n4366), .A2(n4916), .A3(n5785), .ZN(n5789) );
  NAND2_X1 U4884 ( .A1(n5833), .A2(n5777), .ZN(n5883) );
  NAND2_X1 U4885 ( .A1(n5131), .A2(n5130), .ZN(n7328) );
  AOI21_X1 U4886 ( .B1(n8787), .B2(n8795), .A(n6445), .ZN(n8783) );
  INV_X1 U4887 ( .A(n9022), .ZN(n9767) );
  INV_X1 U4888 ( .A(n8209), .ZN(n9762) );
  NAND2_X1 U4889 ( .A1(n5244), .A2(n4924), .ZN(n5264) );
  XNOR2_X1 U4890 ( .A(n5142), .B(SI_6_), .ZN(n5145) );
  INV_X1 U4891 ( .A(n6152), .ZN(n5848) );
  NAND2_X1 U4892 ( .A1(n5654), .A2(n5653), .ZN(n9395) );
  AND2_X1 U4893 ( .A1(n8453), .A2(n9229), .ZN(n9239) );
  INV_X1 U4894 ( .A(n5447), .ZN(n6607) );
  INV_X1 U4895 ( .A(n8734), .ZN(n9827) );
  AND4_X2 U4896 ( .A1(n4400), .A2(n5776), .A3(n5775), .A4(n5779), .ZN(n4366)
         );
  INV_X2 U4897 ( .A(n5875), .ZN(n5937) );
  CLKBUF_X2 U4898 ( .A(n9716), .Z(n4367) );
  INV_X1 U4899 ( .A(n5505), .ZN(n4989) );
  AOI22_X2 U4900 ( .A1(n8722), .A2(n6446), .B1(n6476), .B2(n8714), .ZN(n8709)
         );
  XNOR2_X2 U4901 ( .A(n4985), .B(n4984), .ZN(n5743) );
  NAND2_X4 U4904 ( .A1(n4502), .A2(n4501), .ZN(n4973) );
  OR2_X1 U4907 ( .A1(n6509), .A2(n6508), .ZN(n6510) );
  NOR2_X1 U4908 ( .A1(n5720), .A2(n5721), .ZN(n6509) );
  OAI21_X1 U4909 ( .B1(n8977), .B2(n4696), .A(n4479), .ZN(n5720) );
  AND3_X1 U4910 ( .A1(n8977), .A2(n4483), .A3(n4482), .ZN(n9009) );
  NAND2_X1 U4911 ( .A1(n4671), .A2(n9040), .ZN(n8977) );
  AND2_X1 U4912 ( .A1(n9043), .A2(n5627), .ZN(n4671) );
  AND2_X1 U4913 ( .A1(n4545), .A2(n4426), .ZN(n4543) );
  AOI21_X1 U4914 ( .B1(n8235), .B2(n4665), .A(n9827), .ZN(n4664) );
  XNOR2_X1 U4915 ( .A(n6205), .B(n6204), .ZN(n8964) );
  NAND2_X1 U4916 ( .A1(n4913), .A2(n4912), .ZN(n8854) );
  NAND2_X2 U4917 ( .A1(n5631), .A2(n5630), .ZN(n9402) );
  NAND2_X1 U4918 ( .A1(n5611), .A2(n5610), .ZN(n9407) );
  OR2_X1 U4919 ( .A1(n7547), .A2(n7552), .ZN(n7549) );
  OAI21_X2 U4920 ( .B1(n7612), .B2(n6432), .A(n6270), .ZN(n7624) );
  AOI21_X1 U4921 ( .B1(n4787), .B2(n4425), .A(n4788), .ZN(n7372) );
  OAI21_X1 U4922 ( .B1(n4791), .B2(n4789), .A(n4420), .ZN(n4788) );
  NAND2_X1 U4923 ( .A1(n5966), .A2(n5965), .ZN(n7670) );
  NAND2_X1 U4924 ( .A1(n5936), .A2(n5935), .ZN(n7646) );
  OAI21_X1 U4925 ( .B1(n5415), .B2(n5414), .A(n5413), .ZN(n5444) );
  NAND2_X1 U4926 ( .A1(n5956), .A2(n5955), .ZN(n9891) );
  OAI21_X1 U4927 ( .B1(n5348), .B2(n5326), .A(n5327), .ZN(n5329) );
  NAND2_X1 U4928 ( .A1(n9087), .A2(n9767), .ZN(n8426) );
  NAND2_X2 U4929 ( .A1(n6523), .A2(n6521), .ZN(n6522) );
  OAI211_X1 U4930 ( .C1(n5042), .C2(n6617), .A(n5107), .B(n5106), .ZN(n7251)
         );
  NAND2_X1 U4931 ( .A1(n5869), .A2(n4469), .ZN(n7510) );
  NAND2_X1 U4932 ( .A1(n5844), .A2(n5843), .ZN(n6419) );
  NAND4_X1 U4933 ( .A1(n5121), .A2(n5120), .A3(n5119), .A4(n5118), .ZN(n9085)
         );
  OR2_X2 U4934 ( .A1(n6936), .A2(n7088), .ZN(n8274) );
  INV_X2 U4935 ( .A(n5709), .ZN(n8288) );
  AND2_X2 U4936 ( .A1(n6906), .A2(n6513), .ZN(n5096) );
  NAND2_X1 U4937 ( .A1(n5937), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5831) );
  AOI21_X1 U4938 ( .B1(n5105), .B2(n5104), .A(n4929), .ZN(n5125) );
  NAND4_X1 U4939 ( .A1(n5867), .A2(n5866), .A3(n5865), .A4(n5864), .ZN(n8654)
         );
  AND2_X1 U4940 ( .A1(n5858), .A2(n4556), .ZN(n6951) );
  BUF_X2 U4941 ( .A(n5114), .Z(n8287) );
  NAND2_X1 U4942 ( .A1(n4930), .A2(n4525), .ZN(n6901) );
  CLKBUF_X1 U4943 ( .A(n5739), .Z(n8514) );
  NOR3_X1 U4944 ( .A1(n4920), .A2(n4708), .A3(n5176), .ZN(n4492) );
  NAND2_X1 U4945 ( .A1(n5808), .A2(n5807), .ZN(n7941) );
  NAND2_X1 U4946 ( .A1(n4959), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4982) );
  NAND2_X1 U4947 ( .A1(n8967), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5787) );
  NAND2_X1 U4948 ( .A1(n9457), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4944) );
  INV_X1 U4949 ( .A(n6898), .ZN(n8543) );
  XNOR2_X1 U4950 ( .A(n5047), .B(SI_2_), .ZN(n5045) );
  NAND2_X2 U4951 ( .A1(n6607), .A2(P1_U3084), .ZN(n8557) );
  XNOR2_X1 U4952 ( .A(n4977), .B(n10084), .ZN(n9104) );
  NAND2_X2 U4953 ( .A1(n6607), .A2(P2_U3152), .ZN(n8973) );
  NAND2_X1 U4954 ( .A1(n4957), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4960) );
  INV_X2 U4955 ( .A(n7974), .ZN(n4370) );
  NOR2_X1 U4956 ( .A1(n5784), .A2(n5783), .ZN(n5785) );
  AND2_X1 U4957 ( .A1(n5122), .A2(n5740), .ZN(n4603) );
  AND2_X1 U4958 ( .A1(n5122), .A2(n4953), .ZN(n5150) );
  NOR2_X1 U4959 ( .A1(n4703), .A2(n4955), .ZN(n4701) );
  NAND2_X1 U4960 ( .A1(n5857), .A2(n5856), .ZN(n9473) );
  INV_X1 U4961 ( .A(n5883), .ZN(n5779) );
  NAND2_X1 U4962 ( .A1(n5793), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5905) );
  AND4_X1 U4963 ( .A1(n5772), .A2(n5818), .A3(n5813), .A4(n5812), .ZN(n5776)
         );
  AND2_X1 U4964 ( .A1(n5044), .A2(n5017), .ZN(n4834) );
  AND2_X1 U4965 ( .A1(n4582), .A2(n4581), .ZN(n4935) );
  AND2_X1 U4966 ( .A1(n4669), .A2(n4931), .ZN(n4444) );
  INV_X1 U4967 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n6405) );
  INV_X1 U4968 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n4943) );
  INV_X4 U4969 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  NOR2_X1 U4970 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n5777) );
  NOR2_X1 U4971 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n4581) );
  NOR2_X1 U4972 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n4582) );
  INV_X1 U4973 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n4958) );
  INV_X1 U4974 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n4931) );
  INV_X1 U4975 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5949) );
  INV_X1 U4976 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n6035) );
  INV_X1 U4977 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n4670) );
  INV_X4 U4978 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  INV_X1 U4979 ( .A(n5096), .ZN(n4371) );
  AND2_X2 U4980 ( .A1(n6906), .A2(n6513), .ZN(n4398) );
  AND2_X1 U4981 ( .A1(n8295), .A2(n9370), .ZN(n8400) );
  NAND2_X1 U4982 ( .A1(n5210), .A2(n10029), .ZN(n5237) );
  NOR2_X1 U4983 ( .A1(n9129), .A2(n4600), .ZN(n4599) );
  INV_X1 U4984 ( .A(n9231), .ZN(n4600) );
  INV_X1 U4985 ( .A(n5888), .ZN(n6192) );
  OR2_X1 U4986 ( .A1(n8184), .A2(n8829), .ZN(n4922) );
  OR2_X1 U4987 ( .A1(n8920), .A2(n8841), .ZN(n6441) );
  AND2_X1 U4988 ( .A1(n9107), .A2(n8394), .ZN(n8500) );
  NAND2_X1 U4989 ( .A1(n4454), .A2(n4459), .ZN(n4453) );
  AOI21_X1 U4990 ( .B1(n4463), .B2(n6325), .A(n8743), .ZN(n6330) );
  NOR2_X1 U4991 ( .A1(n8681), .A2(n7171), .ZN(n4748) );
  AND2_X1 U4992 ( .A1(n6352), .A2(n6350), .ZN(n6360) );
  AND2_X1 U4993 ( .A1(n9173), .A2(n8382), .ZN(n4711) );
  NAND2_X1 U4994 ( .A1(n8384), .A2(n8383), .ZN(n4580) );
  NAND2_X1 U4995 ( .A1(n5298), .A2(n5297), .ZN(n5350) );
  INV_X1 U4996 ( .A(n5290), .ZN(n5295) );
  NAND2_X1 U4997 ( .A1(n7696), .A2(n7697), .ZN(n4820) );
  OR2_X1 U4998 ( .A1(n8860), .A2(n6209), .ZN(n6352) );
  OR2_X1 U4999 ( .A1(n8891), .A2(n8774), .ZN(n6327) );
  OR2_X1 U5000 ( .A1(n8896), .A2(n8613), .ZN(n6326) );
  AOI21_X1 U5001 ( .B1(n7209), .B2(n4731), .A(n4730), .ZN(n7551) );
  INV_X1 U5002 ( .A(n6260), .ZN(n4730) );
  AND2_X1 U5003 ( .A1(n6429), .A2(n6259), .ZN(n4731) );
  NAND2_X1 U5004 ( .A1(n8653), .A2(n9869), .ZN(n7093) );
  NAND2_X1 U5005 ( .A1(n6036), .A2(n6035), .ZN(n6187) );
  NAND2_X1 U5006 ( .A1(n9395), .A2(n9245), .ZN(n8466) );
  OAI21_X1 U5007 ( .B1(n4622), .B2(n4620), .A(n4417), .ZN(n4619) );
  INV_X1 U5008 ( .A(n9125), .ZN(n4620) );
  OR2_X1 U5009 ( .A1(n7930), .A2(n8018), .ZN(n8335) );
  OR2_X1 U5010 ( .A1(n5193), .A2(n6750), .ZN(n5218) );
  NAND2_X1 U5011 ( .A1(n6166), .A2(n6165), .ZN(n6181) );
  NAND2_X1 U5012 ( .A1(n5553), .A2(n5552), .ZN(n5578) );
  NAND2_X1 U5013 ( .A1(n5551), .A2(n5550), .ZN(n5553) );
  NAND2_X1 U5014 ( .A1(n5446), .A2(n5445), .ZN(n5476) );
  NAND2_X1 U5015 ( .A1(n5238), .A2(n5237), .ZN(n5244) );
  OAI21_X1 U5016 ( .B1(n5149), .B2(n4490), .A(n4416), .ZN(n5238) );
  INV_X1 U5017 ( .A(n4492), .ZN(n4490) );
  INV_X1 U5018 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n4704) );
  NAND2_X1 U5019 ( .A1(n4491), .A2(n4494), .ZN(n5180) );
  NOR2_X1 U5020 ( .A1(n4920), .A2(n5176), .ZN(n4491) );
  NAND2_X1 U5021 ( .A1(n8256), .A2(n8255), .ZN(n8568) );
  XNOR2_X1 U5022 ( .A(n6951), .B(n6957), .ZN(n6952) );
  INV_X1 U5023 ( .A(n6064), .ZN(n6063) );
  AND2_X1 U5024 ( .A1(n6921), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n4647) );
  AOI21_X1 U5025 ( .B1(n4902), .B2(n4904), .A(n4414), .ZN(n4900) );
  NAND2_X1 U5026 ( .A1(n8761), .A2(n8774), .ZN(n4907) );
  AND2_X1 U5027 ( .A1(n8913), .A2(n8804), .ZN(n6443) );
  AOI22_X1 U5028 ( .A1(n8854), .A2(n6440), .B1(n8179), .B2(n8852), .ZN(n8150)
         );
  NAND2_X1 U5029 ( .A1(n6017), .A2(n6016), .ZN(n8111) );
  AND4_X1 U5030 ( .A1(n6012), .A2(n6011), .A3(n6010), .A4(n6009), .ZN(n8120)
         );
  OR2_X1 U5031 ( .A1(n9528), .A2(n7843), .ZN(n4759) );
  OR3_X1 U5033 ( .A1(n8404), .A2(n8500), .A3(n4570), .ZN(n4569) );
  AND2_X1 U5034 ( .A1(n8405), .A2(n8406), .ZN(n4570) );
  MUX2_X1 U5035 ( .A(n8403), .B(n8402), .S(n8406), .Z(n8404) );
  NAND2_X1 U5036 ( .A1(n4568), .A2(n5505), .ZN(n4567) );
  OAI21_X1 U5037 ( .B1(n4569), .B2(n8508), .A(n8507), .ZN(n4568) );
  AND2_X1 U5038 ( .A1(n4947), .A2(n4948), .ZN(n5114) );
  OR2_X1 U5039 ( .A1(n9395), .A2(n9245), .ZN(n9211) );
  AOI21_X1 U5040 ( .B1(n4599), .B2(n4597), .A(n4412), .ZN(n4596) );
  INV_X1 U5041 ( .A(n9130), .ZN(n4597) );
  INV_X1 U5042 ( .A(n4599), .ZN(n4598) );
  AOI21_X1 U5043 ( .B1(n9253), .B2(n9127), .A(n9126), .ZN(n9237) );
  AOI21_X1 U5044 ( .B1(n4633), .B2(n4631), .A(n4630), .ZN(n4629) );
  NOR2_X1 U5045 ( .A1(n9358), .A2(n9345), .ZN(n4630) );
  INV_X1 U5046 ( .A(n4614), .ZN(n8046) );
  AOI21_X1 U5047 ( .B1(n4609), .B2(n4607), .A(n4422), .ZN(n4606) );
  NAND2_X1 U5048 ( .A1(n4609), .A2(n7960), .ZN(n4608) );
  INV_X2 U5049 ( .A(n5129), .ZN(n8389) );
  NAND2_X1 U5050 ( .A1(n5042), .A2(n5447), .ZN(n5129) );
  XNOR2_X1 U5051 ( .A(n4946), .B(P1_IR_REG_29__SCAN_IN), .ZN(n4948) );
  OR2_X1 U5052 ( .A1(n4945), .A2(n9456), .ZN(n4946) );
  XNOR2_X1 U5053 ( .A(n5673), .B(n5672), .ZN(n7812) );
  NAND2_X1 U5054 ( .A1(n4723), .A2(n5646), .ZN(n5673) );
  INV_X1 U5055 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n4669) );
  INV_X1 U5056 ( .A(n9216), .ZN(n9245) );
  AND2_X1 U5057 ( .A1(n7567), .A2(n6270), .ZN(n4458) );
  NAND2_X1 U5058 ( .A1(n6265), .A2(n6266), .ZN(n4459) );
  AOI21_X1 U5059 ( .B1(n4460), .B2(n4456), .A(n4455), .ZN(n4454) );
  NAND2_X1 U5060 ( .A1(n6262), .A2(n7552), .ZN(n4460) );
  INV_X1 U5061 ( .A(n4459), .ZN(n4456) );
  INV_X1 U5062 ( .A(n6269), .ZN(n4455) );
  AOI21_X1 U5063 ( .B1(n4576), .B2(n4574), .A(n4419), .ZN(n4573) );
  NOR2_X1 U5064 ( .A1(n8406), .A2(n4575), .ZN(n4574) );
  OAI21_X1 U5065 ( .B1(n8328), .B2(n8327), .A(n8416), .ZN(n4576) );
  OAI21_X1 U5066 ( .B1(n4447), .B2(n4446), .A(n4445), .ZN(n6306) );
  NAND2_X1 U5067 ( .A1(n6312), .A2(n6318), .ZN(n4446) );
  AND2_X1 U5068 ( .A1(n6309), .A2(n6342), .ZN(n4466) );
  NAND2_X1 U5069 ( .A1(n8652), .A2(n9823), .ZN(n6252) );
  INV_X1 U5070 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5818) );
  INV_X1 U5071 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5816) );
  INV_X1 U5072 ( .A(n4925), .ZN(n4477) );
  NOR2_X1 U5073 ( .A1(n5185), .A2(n4710), .ZN(n4709) );
  INV_X1 U5074 ( .A(n5179), .ZN(n4710) );
  INV_X1 U5075 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4505) );
  INV_X1 U5076 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4503) );
  AOI21_X1 U5077 ( .B1(n4823), .B2(n4829), .A(n4413), .ZN(n4822) );
  NAND2_X1 U5078 ( .A1(n8036), .A2(n4800), .ZN(n4799) );
  INV_X1 U5079 ( .A(n7830), .ZN(n4800) );
  NAND2_X1 U5080 ( .A1(n6217), .A2(n4747), .ZN(n4746) );
  INV_X1 U5081 ( .A(n4748), .ZN(n4747) );
  NAND2_X1 U5082 ( .A1(n8688), .A2(n4748), .ZN(n4745) );
  INV_X1 U5083 ( .A(n6357), .ZN(n4462) );
  INV_X1 U5084 ( .A(n9473), .ZN(n6554) );
  INV_X1 U5085 ( .A(n4766), .ZN(n4763) );
  INV_X1 U5086 ( .A(n4765), .ZN(n4764) );
  OR2_X1 U5087 ( .A1(n8876), .A2(n8702), .ZN(n6339) );
  NOR2_X1 U5088 ( .A1(n8876), .A2(n8883), .ZN(n4550) );
  NAND2_X1 U5089 ( .A1(n4767), .A2(n8723), .ZN(n4766) );
  NOR2_X1 U5090 ( .A1(n8765), .A2(n4906), .ZN(n4905) );
  INV_X1 U5091 ( .A(n4921), .ZN(n4906) );
  NAND2_X1 U5092 ( .A1(n8798), .A2(n4770), .ZN(n4769) );
  NOR2_X1 U5093 ( .A1(n8782), .A2(n4771), .ZN(n4770) );
  INV_X1 U5094 ( .A(n6322), .ZN(n4771) );
  INV_X1 U5095 ( .A(n4741), .ZN(n4735) );
  NOR2_X1 U5096 ( .A1(n8149), .A2(n4742), .ZN(n4741) );
  INV_X1 U5097 ( .A(n6363), .ZN(n4742) );
  OAI21_X1 U5098 ( .B1(n8149), .B2(n4740), .A(n6312), .ZN(n4739) );
  NAND2_X1 U5099 ( .A1(n6297), .A2(n6363), .ZN(n4740) );
  NOR2_X1 U5100 ( .A1(n4739), .A2(n8827), .ZN(n4737) );
  AND2_X1 U5101 ( .A1(n6034), .A2(n6298), .ZN(n6296) );
  NAND2_X1 U5102 ( .A1(n7551), .A2(n5947), .ZN(n7476) );
  NAND2_X1 U5103 ( .A1(n4564), .A2(n7563), .ZN(n4563) );
  NOR2_X1 U5104 ( .A1(n7129), .A2(n7221), .ZN(n4564) );
  NAND2_X1 U5105 ( .A1(n5794), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5918) );
  INV_X1 U5106 ( .A(n5905), .ZN(n5794) );
  NAND2_X1 U5107 ( .A1(n6252), .A2(n6235), .ZN(n7094) );
  INV_X1 U5108 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5778) );
  NAND2_X1 U5109 ( .A1(n5786), .A2(n4918), .ZN(n4917) );
  INV_X1 U5110 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5786) );
  INV_X1 U5111 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n4918) );
  INV_X1 U5112 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5820) );
  INV_X1 U5113 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5812) );
  AND2_X1 U5114 ( .A1(n7857), .A2(n5371), .ZN(n5377) );
  NOR2_X1 U5115 ( .A1(n4693), .A2(n4689), .ZN(n4688) );
  INV_X1 U5116 ( .A(n5235), .ZN(n4689) );
  INV_X1 U5117 ( .A(n4694), .ZN(n4693) );
  AND2_X1 U5118 ( .A1(n5377), .A2(n4691), .ZN(n4690) );
  NAND2_X1 U5119 ( .A1(n4694), .A2(n4692), .ZN(n4691) );
  INV_X1 U5120 ( .A(n7713), .ZN(n4692) );
  AND2_X1 U5121 ( .A1(n4473), .A2(n8008), .ZN(n5378) );
  NAND2_X1 U5122 ( .A1(n5371), .A2(n5370), .ZN(n4473) );
  NAND2_X1 U5123 ( .A1(n4433), .A2(n4700), .ZN(n4699) );
  NAND2_X1 U5124 ( .A1(n4377), .A2(n9003), .ZN(n4698) );
  INV_X1 U5125 ( .A(n9064), .ZN(n4700) );
  INV_X1 U5126 ( .A(n4926), .ZN(n4697) );
  NAND2_X1 U5127 ( .A1(n5332), .A2(n5129), .ZN(n4499) );
  NAND2_X1 U5128 ( .A1(n4395), .A2(n4500), .ZN(n4497) );
  INV_X1 U5129 ( .A(n5332), .ZN(n4500) );
  AND3_X1 U5130 ( .A1(n4932), .A2(n4933), .A3(n4934), .ZN(n4524) );
  OR2_X1 U5131 ( .A1(n5246), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n5310) );
  INV_X1 U5132 ( .A(n9196), .ZN(n4849) );
  INV_X1 U5133 ( .A(n9151), .ZN(n4847) );
  OR2_X1 U5134 ( .A1(n9179), .A2(n9157), .ZN(n8458) );
  OR2_X1 U5135 ( .A1(n9385), .A2(n9176), .ZN(n9151) );
  AND2_X1 U5136 ( .A1(n8466), .A2(n9229), .ZN(n9149) );
  OR2_X1 U5137 ( .A1(n9391), .A2(n9131), .ZN(n8467) );
  OR2_X1 U5138 ( .A1(n9410), .A2(n9291), .ZN(n9146) );
  OR2_X1 U5139 ( .A1(n9417), .A2(n9124), .ZN(n8469) );
  NOR2_X1 U5140 ( .A1(n8049), .A2(n7905), .ZN(n4864) );
  NOR2_X1 U5141 ( .A1(n7930), .A2(n7959), .ZN(n4533) );
  INV_X1 U5142 ( .A(n7536), .ZN(n4589) );
  OR2_X1 U5143 ( .A1(n7534), .A2(n8327), .ZN(n4862) );
  NOR2_X1 U5144 ( .A1(n4537), .A2(n7595), .ZN(n4535) );
  NAND2_X1 U5145 ( .A1(n4584), .A2(n4374), .ZN(n4586) );
  OR2_X1 U5146 ( .A1(n7581), .A2(n7328), .ZN(n4537) );
  NAND2_X1 U5147 ( .A1(n5155), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5193) );
  NAND2_X1 U5148 ( .A1(n9773), .A2(n9085), .ZN(n8434) );
  NAND2_X1 U5149 ( .A1(n5115), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5157) );
  INV_X1 U5150 ( .A(n5116), .ZN(n5115) );
  XNOR2_X1 U5151 ( .A(n6200), .B(n6199), .ZN(n6197) );
  OAI21_X1 U5152 ( .B1(n5629), .B2(n4726), .A(n4724), .ZN(n5680) );
  INV_X1 U5153 ( .A(n4725), .ZN(n4724) );
  OAI21_X1 U5154 ( .B1(n4728), .B2(n4726), .A(n5674), .ZN(n4725) );
  NAND2_X1 U5155 ( .A1(n5646), .A2(n4727), .ZN(n4726) );
  AOI21_X1 U5156 ( .B1(n5495), .B2(n4716), .A(n4714), .ZN(n4713) );
  INV_X1 U5157 ( .A(n4716), .ZN(n4715) );
  INV_X1 U5158 ( .A(n5523), .ZN(n4714) );
  OR2_X1 U5159 ( .A1(n5351), .A2(P1_IR_REG_13__SCAN_IN), .ZN(n5423) );
  NOR2_X1 U5160 ( .A1(n5347), .A2(n4722), .ZN(n4721) );
  INV_X1 U5161 ( .A(n5263), .ZN(n4722) );
  OR2_X1 U5162 ( .A1(n5303), .A2(n5302), .ZN(n5349) );
  XNOR2_X1 U5163 ( .A(n5291), .B(SI_11_), .ZN(n5285) );
  NAND2_X1 U5164 ( .A1(n5264), .A2(n5263), .ZN(n5348) );
  AND2_X1 U5165 ( .A1(n5263), .A2(n5243), .ZN(n4924) );
  NAND2_X1 U5166 ( .A1(n5182), .A2(n5181), .ZN(n5207) );
  AND2_X1 U5167 ( .A1(n5237), .A2(n5212), .ZN(n4923) );
  NAND2_X1 U5168 ( .A1(n5180), .A2(n4709), .ZN(n5208) );
  INV_X1 U5169 ( .A(n5145), .ZN(n5146) );
  NAND2_X1 U5170 ( .A1(n5149), .A2(n5148), .ZN(n4494) );
  NAND2_X1 U5171 ( .A1(n5125), .A2(n5124), .ZN(n5149) );
  NOR2_X1 U5172 ( .A1(n7833), .A2(n4802), .ZN(n4801) );
  INV_X1 U5173 ( .A(n4804), .ZN(n4802) );
  AND2_X1 U5174 ( .A1(n8560), .A2(n4783), .ZN(n4782) );
  NAND2_X1 U5175 ( .A1(n4784), .A2(n8270), .ZN(n4783) );
  INV_X1 U5176 ( .A(n8622), .ZN(n4784) );
  NAND2_X1 U5177 ( .A1(n8656), .A2(n8274), .ZN(n6953) );
  NAND2_X1 U5178 ( .A1(n4830), .A2(n4390), .ZN(n4827) );
  NAND2_X1 U5179 ( .A1(n8600), .A2(n4831), .ZN(n4830) );
  INV_X1 U5180 ( .A(n8243), .ZN(n4831) );
  AOI21_X1 U5181 ( .B1(n8172), .B2(n8171), .A(n8170), .ZN(n8176) );
  AND2_X1 U5182 ( .A1(n8169), .A2(n8168), .ZN(n8170) );
  NAND2_X1 U5183 ( .A1(n6019), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6028) );
  NAND2_X1 U5184 ( .A1(n7433), .A2(n7171), .ZN(n7088) );
  NAND2_X1 U5185 ( .A1(n4812), .A2(n4811), .ZN(n7758) );
  INV_X1 U5186 ( .A(n7703), .ZN(n4813) );
  NAND2_X1 U5187 ( .A1(n5797), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5968) );
  INV_X1 U5188 ( .A(n5957), .ZN(n5797) );
  OR2_X1 U5189 ( .A1(n6028), .A2(n8071), .ZN(n6041) );
  INV_X2 U5190 ( .A(n8274), .ZN(n8271) );
  INV_X1 U5191 ( .A(n6393), .ZN(n6392) );
  AND4_X1 U5192 ( .A1(n5946), .A2(n5945), .A3(n5944), .A4(n5943), .ZN(n7553)
         );
  OR2_X1 U5193 ( .A1(n5890), .A2(n5862), .ZN(n5866) );
  OR2_X1 U5194 ( .A1(n9473), .A2(n4661), .ZN(n4660) );
  NAND2_X1 U5195 ( .A1(n9473), .A2(n4661), .ZN(n4659) );
  NOR2_X1 U5196 ( .A1(n6585), .A2(n6584), .ZN(n6806) );
  OR2_X1 U5197 ( .A1(n6810), .A2(n6809), .ZN(n4652) );
  AND2_X1 U5198 ( .A1(n8750), .A2(n4386), .ZN(n8686) );
  NAND2_X1 U5199 ( .A1(n8750), .A2(n4548), .ZN(n8694) );
  AND2_X1 U5200 ( .A1(n6339), .A2(n6338), .ZN(n6447) );
  NAND2_X1 U5201 ( .A1(n6447), .A2(n6135), .ZN(n4765) );
  INV_X1 U5202 ( .A(n6447), .ZN(n8713) );
  NOR2_X1 U5203 ( .A1(n8745), .A2(n4766), .ZN(n8726) );
  NAND2_X1 U5204 ( .A1(n8723), .A2(n6222), .ZN(n8739) );
  INV_X1 U5205 ( .A(n8891), .ZN(n8761) );
  OR2_X1 U5206 ( .A1(n8780), .A2(n8613), .ZN(n4921) );
  NAND2_X1 U5207 ( .A1(n8898), .A2(n4905), .ZN(n4908) );
  AND2_X1 U5208 ( .A1(n6327), .A2(n6325), .ZN(n8765) );
  NOR2_X1 U5209 ( .A1(n8903), .A2(n6444), .ZN(n6445) );
  AND2_X1 U5210 ( .A1(n6114), .A2(n6113), .ZN(n8774) );
  OR2_X1 U5211 ( .A1(n8903), .A2(n8775), .ZN(n6322) );
  INV_X1 U5212 ( .A(n4769), .ZN(n8771) );
  NAND2_X1 U5213 ( .A1(n6326), .A2(n6311), .ZN(n8782) );
  NOR2_X1 U5214 ( .A1(n8818), .A2(n8908), .ZN(n4553) );
  NAND2_X1 U5215 ( .A1(n4553), .A2(n4552), .ZN(n8788) );
  AND2_X1 U5216 ( .A1(n6322), .A2(n6308), .ZN(n8786) );
  AND2_X1 U5217 ( .A1(n6060), .A2(n6059), .ZN(n8829) );
  NAND2_X1 U5218 ( .A1(n8837), .A2(n4741), .ZN(n4738) );
  INV_X1 U5219 ( .A(n4739), .ZN(n4736) );
  NOR2_X1 U5220 ( .A1(n8920), .A2(n8844), .ZN(n8817) );
  NAND2_X1 U5221 ( .A1(n6048), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6212) );
  AOI21_X1 U5222 ( .B1(n4753), .B2(n4750), .A(n4752), .ZN(n4749) );
  INV_X1 U5223 ( .A(n6296), .ZN(n8030) );
  NAND2_X1 U5224 ( .A1(n8111), .A2(n8640), .ZN(n4914) );
  OR2_X1 U5225 ( .A1(n7948), .A2(n7949), .ZN(n4915) );
  NOR2_X1 U5226 ( .A1(n6226), .A2(n4758), .ZN(n4757) );
  INV_X1 U5227 ( .A(n4759), .ZN(n4758) );
  AOI21_X1 U5228 ( .B1(n4757), .B2(n4755), .A(n4754), .ZN(n4753) );
  AND2_X1 U5229 ( .A1(n6228), .A2(n6227), .ZN(n7841) );
  NAND2_X1 U5230 ( .A1(n7741), .A2(n6438), .ZN(n7796) );
  AOI21_X1 U5231 ( .B1(n7743), .B2(n7742), .A(n6285), .ZN(n7803) );
  NAND2_X1 U5232 ( .A1(n7803), .A2(n7804), .ZN(n7807) );
  OR2_X1 U5233 ( .A1(n5991), .A2(n5990), .ZN(n5993) );
  NAND2_X1 U5234 ( .A1(n4894), .A2(n4893), .ZN(n4892) );
  NOR2_X1 U5235 ( .A1(n7572), .A2(n6431), .ZN(n4893) );
  OR2_X1 U5236 ( .A1(n7700), .A2(n8645), .ZN(n4899) );
  OR2_X1 U5237 ( .A1(n7618), .A2(n9891), .ZN(n7635) );
  AND4_X1 U5238 ( .A1(n5933), .A2(n5932), .A3(n5931), .A4(n5930), .ZN(n7474)
         );
  NAND2_X1 U5239 ( .A1(n7085), .A2(n7094), .ZN(n4911) );
  AND4_X1 U5240 ( .A1(n5879), .A2(n5878), .A3(n5877), .A4(n5876), .ZN(n7211)
         );
  AND4_X1 U5241 ( .A1(n5924), .A2(n5923), .A3(n5922), .A4(n5921), .ZN(n7554)
         );
  AND2_X1 U5242 ( .A1(n7207), .A2(n7222), .ZN(n5911) );
  XNOR2_X1 U5243 ( .A(n7221), .B(n8651), .ZN(n7222) );
  NAND2_X1 U5244 ( .A1(n7510), .A2(n4451), .ZN(n7359) );
  INV_X1 U5245 ( .A(n8654), .ZN(n4451) );
  NOR2_X1 U5246 ( .A1(n7505), .A2(n7510), .ZN(n7504) );
  XNOR2_X1 U5247 ( .A(n8654), .B(n5870), .ZN(n7493) );
  NAND2_X1 U5248 ( .A1(n6050), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n4471) );
  NAND2_X1 U5249 ( .A1(n8867), .A2(n9882), .ZN(n4544) );
  OR2_X1 U5250 ( .A1(n8870), .A2(n9532), .ZN(n4545) );
  AND2_X1 U5251 ( .A1(n5886), .A2(n5885), .ZN(n9869) );
  NAND2_X1 U5252 ( .A1(n6565), .A2(n4554), .ZN(n4556) );
  NAND2_X1 U5253 ( .A1(n4555), .A2(n4410), .ZN(n4554) );
  NAND2_X1 U5254 ( .A1(n4467), .A2(n4366), .ZN(n5808) );
  AND2_X1 U5255 ( .A1(n5785), .A2(n4468), .ZN(n4467) );
  INV_X1 U5256 ( .A(n4917), .ZN(n4468) );
  NOR2_X1 U5257 ( .A1(n6188), .A2(P2_IR_REG_18__SCAN_IN), .ZN(n6189) );
  INV_X1 U5258 ( .A(n6187), .ZN(n6190) );
  NAND2_X1 U5259 ( .A1(n4472), .A2(n5368), .ZN(n7979) );
  INV_X1 U5260 ( .A(n5378), .ZN(n4472) );
  NAND2_X1 U5261 ( .A1(n5354), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n5398) );
  INV_X1 U5262 ( .A(n5356), .ZN(n5354) );
  INV_X1 U5263 ( .A(n9053), .ZN(n4680) );
  AND2_X1 U5264 ( .A1(n5494), .A2(n4680), .ZN(n4679) );
  INV_X1 U5265 ( .A(n5470), .ZN(n4676) );
  NOR2_X1 U5266 ( .A1(n6615), .A2(n6607), .ZN(n4526) );
  NAND2_X1 U5267 ( .A1(n8142), .A2(n8137), .ZN(n8160) );
  AND2_X1 U5268 ( .A1(n5572), .A2(n5592), .ZN(n4672) );
  AND2_X1 U5269 ( .A1(n9370), .A2(n9106), .ZN(n8540) );
  OR2_X1 U5270 ( .A1(n9111), .A2(n9158), .ZN(n8539) );
  NAND2_X1 U5271 ( .A1(n4919), .A2(n4874), .ZN(n4873) );
  AND3_X1 U5272 ( .A1(n4524), .A2(n4935), .A3(n5740), .ZN(n4522) );
  INV_X1 U5273 ( .A(n4939), .ZN(n4521) );
  NAND2_X1 U5274 ( .A1(n8509), .A2(n4989), .ZN(n4566) );
  AND2_X1 U5275 ( .A1(n4947), .A2(n8109), .ZN(n6642) );
  AND2_X1 U5276 ( .A1(n9626), .A2(n6699), .ZN(n9642) );
  NAND2_X1 U5277 ( .A1(n9656), .A2(n9655), .ZN(n4511) );
  NAND2_X1 U5278 ( .A1(n4511), .A2(n4510), .ZN(n4509) );
  NAND2_X1 U5279 ( .A1(n9667), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n4510) );
  NAND2_X1 U5280 ( .A1(n4509), .A2(n4508), .ZN(n4507) );
  INV_X1 U5281 ( .A(n6704), .ZN(n4508) );
  NOR2_X1 U5282 ( .A1(n7402), .A2(n4512), .ZN(n7767) );
  AND2_X1 U5283 ( .A1(n7403), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4512) );
  NOR2_X1 U5284 ( .A1(n9189), .A2(n9179), .ZN(n9178) );
  AND2_X1 U5285 ( .A1(n8465), .A2(n8535), .ZN(n9153) );
  NAND2_X1 U5286 ( .A1(n9134), .A2(n8497), .ZN(n9172) );
  AND2_X1 U5287 ( .A1(n8458), .A2(n8444), .ZN(n9173) );
  AOI21_X1 U5288 ( .B1(n4853), .B2(n4852), .A(n8441), .ZN(n4851) );
  INV_X1 U5289 ( .A(n9149), .ZN(n4852) );
  NAND2_X1 U5290 ( .A1(n9238), .A2(n9149), .ZN(n9212) );
  NAND2_X1 U5291 ( .A1(n4595), .A2(n4594), .ZN(n9202) );
  AOI21_X1 U5292 ( .B1(n4596), .B2(n4598), .A(n9214), .ZN(n4594) );
  NAND2_X1 U5293 ( .A1(n9211), .A2(n8466), .ZN(n9231) );
  OR2_X1 U5294 ( .A1(n5632), .A2(n10069), .ZN(n5657) );
  NAND2_X1 U5295 ( .A1(n9254), .A2(n9148), .ZN(n9238) );
  AND2_X1 U5296 ( .A1(n9239), .A2(n9240), .ZN(n9148) );
  NAND2_X1 U5297 ( .A1(n9257), .A2(n9147), .ZN(n9254) );
  AND2_X1 U5298 ( .A1(n9255), .A2(n9256), .ZN(n9147) );
  INV_X1 U5299 ( .A(n4617), .ZN(n9253) );
  NAND2_X1 U5300 ( .A1(n4624), .A2(n9125), .ZN(n4621) );
  INV_X1 U5301 ( .A(n4619), .ZN(n4618) );
  NOR2_X1 U5302 ( .A1(n9292), .A2(n9410), .ZN(n9274) );
  AOI21_X1 U5303 ( .B1(n4624), .B2(n4623), .A(n4421), .ZN(n4622) );
  INV_X1 U5304 ( .A(n9122), .ZN(n4623) );
  OAI21_X1 U5305 ( .B1(n9308), .B2(n9144), .A(n9143), .ZN(n9287) );
  NAND2_X1 U5306 ( .A1(n8469), .A2(n9145), .ZN(n9288) );
  NAND2_X1 U5307 ( .A1(n9420), .A2(n9327), .ZN(n9122) );
  NOR2_X1 U5308 ( .A1(n4636), .A2(n9119), .ZN(n4635) );
  INV_X1 U5309 ( .A(n4384), .ZN(n4636) );
  NAND2_X1 U5310 ( .A1(n4634), .A2(n4640), .ZN(n4633) );
  INV_X1 U5311 ( .A(n4637), .ZN(n4634) );
  AND2_X1 U5312 ( .A1(n8422), .A2(n9139), .ZN(n9546) );
  NOR2_X1 U5313 ( .A1(n9546), .A2(n4638), .ZN(n4637) );
  INV_X1 U5314 ( .A(n4641), .ZN(n4638) );
  OR2_X1 U5315 ( .A1(n9117), .A2(n9538), .ZN(n4641) );
  NOR2_X1 U5316 ( .A1(n7904), .A2(n4612), .ZN(n4611) );
  INV_X1 U5317 ( .A(n7779), .ZN(n4612) );
  NAND2_X1 U5318 ( .A1(n4610), .A2(n4616), .ZN(n4609) );
  NAND2_X1 U5319 ( .A1(n7905), .A2(n4613), .ZN(n4610) );
  NAND2_X1 U5320 ( .A1(n4391), .A2(n7779), .ZN(n4613) );
  NOR2_X1 U5321 ( .A1(n9505), .A2(n9504), .ZN(n9506) );
  INV_X1 U5322 ( .A(n8391), .ZN(n5506) );
  INV_X1 U5323 ( .A(n8479), .ZN(n4592) );
  INV_X1 U5324 ( .A(n7421), .ZN(n4583) );
  NAND2_X1 U5325 ( .A1(n8434), .A2(n8310), .ZN(n8307) );
  NAND2_X1 U5326 ( .A1(n8307), .A2(n7173), .ZN(n7296) );
  NAND2_X1 U5327 ( .A1(n9714), .A2(n6903), .ZN(n8521) );
  NAND2_X1 U5328 ( .A1(n4367), .A2(n9715), .ZN(n9714) );
  INV_X1 U5329 ( .A(n9348), .ZN(n9711) );
  NAND2_X1 U5330 ( .A1(n8393), .A2(n8392), .ZN(n9376) );
  NAND2_X1 U5331 ( .A1(n5483), .A2(n5482), .ZN(n9432) );
  INV_X1 U5332 ( .A(n6901), .ZN(n9757) );
  NOR2_X1 U5333 ( .A1(n4967), .A2(n4871), .ZN(n4945) );
  NAND2_X1 U5334 ( .A1(n4872), .A2(n4975), .ZN(n4871) );
  NAND2_X1 U5335 ( .A1(n4705), .A2(n6144), .ZN(n6161) );
  NAND2_X1 U5336 ( .A1(n6142), .A2(n6143), .ZN(n4705) );
  NAND2_X1 U5337 ( .A1(n5701), .A2(n5700), .ZN(n6142) );
  NAND2_X1 U5338 ( .A1(n4983), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4985) );
  XNOR2_X1 U5339 ( .A(n4960), .B(P1_IR_REG_20__SCAN_IN), .ZN(n6898) );
  NAND2_X1 U5340 ( .A1(n4718), .A2(n5499), .ZN(n5522) );
  NAND2_X1 U5341 ( .A1(n5497), .A2(n5496), .ZN(n4718) );
  XNOR2_X1 U5342 ( .A(n5075), .B(SI_3_), .ZN(n5073) );
  NAND2_X1 U5343 ( .A1(n5824), .A2(n5823), .ZN(n9528) );
  NAND2_X1 U5344 ( .A1(n6094), .A2(n6093), .ZN(n8896) );
  AND2_X1 U5345 ( .A1(n6071), .A2(n6070), .ZN(n8579) );
  AND3_X1 U5346 ( .A1(n6045), .A2(n6044), .A3(n6043), .ZN(n8179) );
  NAND2_X1 U5347 ( .A1(n7011), .A2(n4794), .ZN(n4793) );
  INV_X1 U5348 ( .A(n7071), .ZN(n4794) );
  INV_X1 U5349 ( .A(n4792), .ZN(n4791) );
  OAI21_X1 U5350 ( .B1(n7061), .B2(n4793), .A(n4795), .ZN(n4792) );
  NAND2_X1 U5351 ( .A1(n7069), .A2(n7070), .ZN(n4795) );
  OR2_X1 U5352 ( .A1(n8261), .A2(n8260), .ZN(n8262) );
  OR2_X1 U5353 ( .A1(n4809), .A2(n7002), .ZN(n4807) );
  AND2_X1 U5354 ( .A1(n7003), .A2(n7144), .ZN(n4808) );
  NAND2_X1 U5355 ( .A1(n8116), .A2(n8069), .ZN(n8131) );
  NAND2_X1 U5356 ( .A1(n6027), .A2(n6026), .ZN(n8930) );
  XNOR2_X1 U5357 ( .A(n8258), .B(n8259), .ZN(n8591) );
  NAND2_X1 U5358 ( .A1(n6038), .A2(n6037), .ZN(n8923) );
  NAND2_X1 U5359 ( .A1(n7060), .A2(n7061), .ZN(n7059) );
  AND2_X1 U5360 ( .A1(n6937), .A2(n9882), .ZN(n8629) );
  AND2_X1 U5361 ( .A1(n6134), .A2(n6133), .ZN(n8714) );
  INV_X1 U5362 ( .A(n8263), .ZN(n8767) );
  INV_X1 U5363 ( .A(n6866), .ZN(n4648) );
  INV_X1 U5364 ( .A(n4666), .ZN(n4665) );
  OAI21_X1 U5365 ( .B1(n8236), .B2(n9811), .A(n9809), .ZN(n4666) );
  OAI22_X1 U5366 ( .A1(n8238), .A2(n8657), .B1(n9811), .B2(n8237), .ZN(n4668)
         );
  AOI21_X1 U5367 ( .B1(n6475), .B2(n8843), .A(n6474), .ZN(n8869) );
  NAND2_X1 U5368 ( .A1(n6473), .A2(n6472), .ZN(n6474) );
  XNOR2_X1 U5369 ( .A(n6466), .B(n6448), .ZN(n6475) );
  OAI21_X1 U5370 ( .B1(n8709), .B2(n4881), .A(n4876), .ZN(n8870) );
  NAND2_X1 U5371 ( .A1(n6467), .A2(n4882), .ZN(n4881) );
  AOI21_X1 U5372 ( .B1(n8709), .B2(n4880), .A(n4877), .ZN(n4876) );
  AND2_X1 U5373 ( .A1(n4883), .A2(n6448), .ZN(n4880) );
  XNOR2_X1 U5374 ( .A(n6212), .B(P2_IR_REG_19__SCAN_IN), .ZN(n8734) );
  NAND2_X1 U5375 ( .A1(n7812), .A2(n8389), .ZN(n5654) );
  OR2_X1 U5376 ( .A1(n9207), .A2(n6500), .ZN(n5692) );
  NAND2_X1 U5377 ( .A1(n5664), .A2(n5663), .ZN(n9216) );
  OR2_X1 U5378 ( .A1(n9225), .A2(n6500), .ZN(n5664) );
  NAND4_X1 U5379 ( .A1(n5198), .A2(n5197), .A3(n5196), .A4(n5195), .ZN(n9083)
         );
  NAND2_X1 U5380 ( .A1(n5095), .A2(n4388), .ZN(n9086) );
  INV_X1 U5381 ( .A(n5042), .ZN(n9601) );
  AND2_X1 U5382 ( .A1(n9642), .A2(n9643), .ZN(n9645) );
  OAI21_X1 U5383 ( .B1(n9097), .B2(n9659), .A(n4520), .ZN(n4519) );
  OR2_X1 U5384 ( .A1(n9098), .A2(n9636), .ZN(n4520) );
  OAI21_X1 U5385 ( .B1(n9101), .B2(n9100), .A(n9099), .ZN(n4516) );
  NAND2_X1 U5386 ( .A1(n9160), .A2(n4540), .ZN(n9374) );
  OR2_X1 U5387 ( .A1(n9178), .A2(n9161), .ZN(n4540) );
  NAND2_X1 U5388 ( .A1(n4393), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4986) );
  OAI21_X1 U5389 ( .B1(n6254), .B2(n4411), .A(n4449), .ZN(n6236) );
  NOR2_X1 U5390 ( .A1(n4450), .A2(n5898), .ZN(n4449) );
  INV_X1 U5391 ( .A(n6259), .ZN(n4450) );
  INV_X1 U5392 ( .A(n8410), .ZN(n4575) );
  AND2_X1 U5393 ( .A1(n6271), .A2(n4458), .ZN(n4457) );
  NAND2_X1 U5394 ( .A1(n4578), .A2(n8406), .ZN(n4577) );
  INV_X1 U5395 ( .A(n8332), .ZN(n4578) );
  AOI21_X1 U5396 ( .B1(n6314), .B2(n6362), .A(n4448), .ZN(n4447) );
  NAND2_X1 U5397 ( .A1(n6315), .A2(n6363), .ZN(n4448) );
  AND2_X1 U5398 ( .A1(n6321), .A2(n6316), .ZN(n4445) );
  OAI21_X1 U5399 ( .B1(n4465), .B2(n4464), .A(n6324), .ZN(n4463) );
  NOR2_X1 U5400 ( .A1(n6311), .A2(n6342), .ZN(n4464) );
  AOI211_X1 U5401 ( .C1(n6310), .C2(n6353), .A(n8782), .B(n4466), .ZN(n4465)
         );
  INV_X1 U5402 ( .A(n5207), .ZN(n4708) );
  INV_X1 U5403 ( .A(n8576), .ZN(n4825) );
  AND2_X1 U5404 ( .A1(n6218), .A2(n6351), .ZN(n6361) );
  OR2_X1 U5405 ( .A1(n8883), .A2(n8714), .ZN(n6334) );
  AND2_X1 U5406 ( .A1(n8006), .A2(n5344), .ZN(n5371) );
  INV_X1 U5407 ( .A(n8387), .ZN(n8399) );
  OAI21_X1 U5408 ( .B1(n6181), .B2(n6180), .A(n6179), .ZN(n6200) );
  INV_X1 U5409 ( .A(n5672), .ZN(n4727) );
  AND2_X1 U5410 ( .A1(n5499), .A2(n4717), .ZN(n4716) );
  INV_X1 U5411 ( .A(n5521), .ZN(n4717) );
  OR2_X1 U5412 ( .A1(n5326), .A2(n5295), .ZN(n5346) );
  NAND2_X1 U5413 ( .A1(n4492), .A2(n4489), .ZN(n4488) );
  INV_X1 U5414 ( .A(n5148), .ZN(n4489) );
  INV_X1 U5415 ( .A(n4707), .ZN(n4706) );
  OAI21_X1 U5416 ( .B1(n4709), .B2(n4708), .A(n4923), .ZN(n4707) );
  NAND2_X1 U5417 ( .A1(n5241), .A2(n5240), .ZN(n5263) );
  AOI21_X1 U5418 ( .B1(n4376), .B2(n4799), .A(n4407), .ZN(n4798) );
  INV_X1 U5419 ( .A(n7345), .ZN(n4789) );
  INV_X1 U5420 ( .A(n4793), .ZN(n4790) );
  NOR2_X1 U5421 ( .A1(n8658), .A2(n4443), .ZN(n8231) );
  NAND2_X1 U5422 ( .A1(n8699), .A2(n4886), .ZN(n4885) );
  NAND2_X1 U5423 ( .A1(n6447), .A2(n4888), .ZN(n4886) );
  NOR2_X1 U5424 ( .A1(n8871), .A2(n4549), .ZN(n4548) );
  INV_X1 U5425 ( .A(n4550), .ZN(n4549) );
  NOR2_X1 U5426 ( .A1(n4903), .A2(n8744), .ZN(n4902) );
  NOR2_X1 U5427 ( .A1(n4905), .A2(n4904), .ZN(n4903) );
  INV_X1 U5428 ( .A(n4907), .ZN(n4904) );
  NOR2_X1 U5429 ( .A1(n7700), .A2(n7763), .ZN(n4559) );
  INV_X1 U5430 ( .A(n7478), .ZN(n7472) );
  INV_X1 U5431 ( .A(n6426), .ZN(n4910) );
  NOR2_X1 U5432 ( .A1(n7094), .A2(n5897), .ZN(n7092) );
  NOR2_X1 U5433 ( .A1(n7356), .A2(n6233), .ZN(n7091) );
  INV_X1 U5434 ( .A(n7359), .ZN(n6233) );
  INV_X1 U5435 ( .A(n7493), .ZN(n7496) );
  INV_X1 U5436 ( .A(n8656), .ZN(n5860) );
  NAND2_X1 U5437 ( .A1(n8656), .A2(n6951), .ZN(n6367) );
  NAND2_X1 U5438 ( .A1(n8777), .A2(n8761), .ZN(n8751) );
  INV_X1 U5439 ( .A(n7307), .ZN(n7310) );
  AND2_X1 U5440 ( .A1(n6237), .A2(n6367), .ZN(n7309) );
  NAND2_X1 U5441 ( .A1(n5854), .A2(n6607), .ZN(n4555) );
  OR2_X1 U5442 ( .A1(n5925), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n5934) );
  AND2_X1 U5443 ( .A1(n8995), .A2(n4476), .ZN(n4475) );
  NAND2_X1 U5444 ( .A1(n9032), .A2(n4477), .ZN(n4476) );
  AND2_X1 U5445 ( .A1(n7819), .A2(n4438), .ZN(n4694) );
  NAND2_X1 U5446 ( .A1(n8387), .A2(n4579), .ZN(n8401) );
  NOR2_X1 U5447 ( .A1(n9152), .A2(n9078), .ZN(n4579) );
  OR2_X1 U5448 ( .A1(n9376), .A2(n9177), .ZN(n8465) );
  INV_X1 U5449 ( .A(n9232), .ZN(n9131) );
  NOR2_X1 U5450 ( .A1(n9402), .A2(n9407), .ZN(n4530) );
  NOR2_X1 U5451 ( .A1(n4529), .A2(n9395), .ZN(n4528) );
  INV_X1 U5452 ( .A(n4530), .ZN(n4529) );
  AND2_X1 U5453 ( .A1(n9420), .A2(n9290), .ZN(n9144) );
  OR2_X1 U5454 ( .A1(n9420), .A2(n9290), .ZN(n9143) );
  OR2_X1 U5455 ( .A1(n9360), .A2(n9140), .ZN(n4844) );
  OR2_X1 U5456 ( .A1(n9432), .A2(n8991), .ZN(n8472) );
  INV_X1 U5457 ( .A(n9120), .ZN(n4632) );
  NOR2_X1 U5458 ( .A1(n4635), .A2(n9120), .ZN(n4631) );
  NOR2_X1 U5459 ( .A1(n4611), .A2(n4615), .ZN(n4607) );
  AOI21_X1 U5460 ( .B1(n4860), .B2(n8327), .A(n4859), .ZN(n4858) );
  INV_X1 U5461 ( .A(n8330), .ZN(n4859) );
  OR2_X1 U5462 ( .A1(n7409), .A2(n7595), .ZN(n8317) );
  NAND2_X1 U5463 ( .A1(n5088), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5116) );
  INV_X1 U5464 ( .A(n4367), .ZN(n9702) );
  NAND2_X1 U5465 ( .A1(n5738), .A2(n4989), .ZN(n6907) );
  NAND2_X1 U5466 ( .A1(n9274), .A2(n9270), .ZN(n9263) );
  NAND2_X1 U5467 ( .A1(n5680), .A2(n5679), .ZN(n5701) );
  NOR2_X1 U5468 ( .A1(n5647), .A2(n4729), .ZN(n4728) );
  INV_X1 U5469 ( .A(n5628), .ZN(n4729) );
  XNOR2_X1 U5470 ( .A(n4982), .B(P1_IR_REG_21__SCAN_IN), .ZN(n5739) );
  INV_X1 U5471 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n4956) );
  NAND2_X1 U5472 ( .A1(n4720), .A2(n4719), .ZN(n5415) );
  AOI21_X1 U5473 ( .B1(n4372), .B2(n5382), .A(n4418), .ZN(n4719) );
  NAND2_X1 U5474 ( .A1(n5264), .A2(n4401), .ZN(n4720) );
  NOR2_X1 U5475 ( .A1(n5295), .A2(n5294), .ZN(n5302) );
  AND2_X1 U5476 ( .A1(n5293), .A2(n5327), .ZN(n5294) );
  NAND2_X1 U5477 ( .A1(n4995), .A2(n4994), .ZN(n5021) );
  NAND3_X1 U5478 ( .A1(n4712), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n4501) );
  INV_X1 U5479 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4712) );
  NAND2_X1 U5480 ( .A1(n7828), .A2(n7829), .ZN(n4804) );
  OR2_X1 U5481 ( .A1(n7831), .A2(n7830), .ZN(n4803) );
  AOI21_X1 U5482 ( .B1(n4782), .B2(n4785), .A(n4423), .ZN(n4780) );
  INV_X1 U5483 ( .A(n8270), .ZN(n4785) );
  NAND2_X1 U5484 ( .A1(n4818), .A2(n4820), .ZN(n4814) );
  OR2_X1 U5485 ( .A1(n4816), .A2(n4821), .ZN(n4815) );
  INV_X1 U5486 ( .A(n4820), .ZN(n4816) );
  INV_X1 U5487 ( .A(n5891), .ZN(n5793) );
  NAND2_X1 U5488 ( .A1(n8257), .A2(n8568), .ZN(n8258) );
  AND2_X1 U5489 ( .A1(n7137), .A2(n4385), .ZN(n4809) );
  NOR2_X1 U5490 ( .A1(n8173), .A2(n8174), .ZN(n8243) );
  NAND2_X1 U5491 ( .A1(n6084), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6096) );
  INV_X1 U5492 ( .A(n6085), .ZN(n6084) );
  NOR2_X1 U5493 ( .A1(n7440), .A2(n7349), .ZN(n4819) );
  NAND2_X1 U5494 ( .A1(n6039), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6053) );
  INV_X1 U5495 ( .A(n6006), .ZN(n6004) );
  OR2_X1 U5496 ( .A1(n7831), .A2(n4799), .ZN(n4797) );
  AND2_X1 U5497 ( .A1(n7088), .A2(n6387), .ZN(n6947) );
  NAND2_X1 U5498 ( .A1(n4424), .A2(n6218), .ZN(n4744) );
  OAI21_X1 U5499 ( .B1(n4461), .B2(n6356), .A(n6388), .ZN(n6393) );
  AOI21_X1 U5500 ( .B1(n6349), .B2(n4399), .A(n4462), .ZN(n4461) );
  NAND2_X1 U5501 ( .A1(n6388), .A2(n9827), .ZN(n6936) );
  AND4_X1 U5502 ( .A1(n5985), .A2(n5984), .A3(n5983), .A4(n5982), .ZN(n7760)
         );
  NOR2_X1 U5503 ( .A1(n9464), .A2(n4658), .ZN(n9462) );
  NAND2_X1 U5504 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n4658) );
  AOI21_X1 U5505 ( .B1(P2_REG2_REG_3__SCAN_IN), .B2(n6557), .A(n6784), .ZN(
        n6575) );
  OR2_X1 U5506 ( .A1(n6800), .A2(n6799), .ZN(n6801) );
  OR2_X1 U5507 ( .A1(n6863), .A2(n4650), .ZN(n4649) );
  AND2_X1 U5508 ( .A1(n6864), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n4650) );
  NOR2_X1 U5509 ( .A1(n7451), .A2(n7450), .ZN(n7517) );
  NOR2_X1 U5510 ( .A1(n8091), .A2(n8090), .ZN(n8226) );
  OR2_X1 U5511 ( .A1(n8226), .A2(n4655), .ZN(n4654) );
  AND2_X1 U5512 ( .A1(n8227), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n4655) );
  NAND2_X1 U5513 ( .A1(n6158), .A2(n8634), .ZN(n6159) );
  NAND2_X1 U5514 ( .A1(n8634), .A2(n8838), .ZN(n6473) );
  INV_X1 U5515 ( .A(n4885), .ZN(n4882) );
  INV_X1 U5516 ( .A(n4884), .ZN(n4883) );
  OAI21_X1 U5517 ( .B1(n4885), .B2(n4888), .A(n4887), .ZN(n4884) );
  NAND2_X1 U5518 ( .A1(n6158), .A2(n8715), .ZN(n4887) );
  INV_X1 U5519 ( .A(n4878), .ZN(n4877) );
  OAI21_X1 U5520 ( .B1(n6467), .B2(n4883), .A(n4879), .ZN(n4878) );
  OAI21_X1 U5521 ( .B1(n6467), .B2(n4882), .A(n4883), .ZN(n4879) );
  INV_X1 U5522 ( .A(n4762), .ZN(n4761) );
  OAI21_X1 U5523 ( .B1(n4765), .B2(n4763), .A(n6339), .ZN(n4762) );
  XNOR2_X1 U5524 ( .A(n8871), .B(n8634), .ZN(n8692) );
  NAND2_X1 U5525 ( .A1(n4889), .A2(n8702), .ZN(n4888) );
  AND2_X1 U5526 ( .A1(n8765), .A2(n6311), .ZN(n4768) );
  OR2_X1 U5527 ( .A1(n6117), .A2(n8586), .ZN(n6127) );
  OR2_X1 U5528 ( .A1(n6096), .A2(n6095), .ZN(n6107) );
  NAND2_X1 U5529 ( .A1(n6106), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6117) );
  INV_X1 U5530 ( .A(n6107), .ZN(n6106) );
  NOR2_X1 U5531 ( .A1(n8788), .A2(n8896), .ZN(n8777) );
  INV_X1 U5532 ( .A(n8786), .ZN(n8795) );
  NAND2_X1 U5533 ( .A1(n4891), .A2(n4890), .ZN(n8787) );
  NAND2_X1 U5534 ( .A1(n8811), .A2(n8831), .ZN(n4890) );
  NAND2_X1 U5535 ( .A1(n8807), .A2(n4402), .ZN(n4891) );
  OAI21_X1 U5536 ( .B1(n4737), .B2(n4734), .A(n4732), .ZN(n8803) );
  NOR2_X1 U5537 ( .A1(n4735), .A2(n4734), .ZN(n4733) );
  INV_X1 U5538 ( .A(n6316), .ZN(n4734) );
  AOI21_X1 U5539 ( .B1(n4375), .B2(n7949), .A(n4406), .ZN(n4912) );
  NAND2_X1 U5540 ( .A1(n7948), .A2(n4375), .ZN(n4913) );
  OR2_X1 U5541 ( .A1(n8846), .A2(n8923), .ZN(n8844) );
  AND2_X1 U5542 ( .A1(n6363), .A2(n6362), .ZN(n8853) );
  NOR2_X1 U5543 ( .A1(n8111), .A2(n7950), .ZN(n8023) );
  NAND2_X1 U5544 ( .A1(n7637), .A2(n4557), .ZN(n7950) );
  AND2_X1 U5545 ( .A1(n4378), .A2(n4558), .ZN(n4557) );
  OAI22_X1 U5546 ( .A1(n7796), .A2(n7804), .B1(n9528), .B2(n8642), .ZN(n7848)
         );
  NAND2_X1 U5547 ( .A1(n7637), .A2(n4378), .ZN(n7849) );
  AND2_X1 U5548 ( .A1(n7637), .A2(n4559), .ZN(n7797) );
  NAND2_X1 U5549 ( .A1(n5798), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5991) );
  INV_X1 U5550 ( .A(n5980), .ZN(n5798) );
  AND2_X1 U5551 ( .A1(n7637), .A2(n9900), .ZN(n7749) );
  AND4_X1 U5552 ( .A1(n5973), .A2(n5972), .A3(n5971), .A4(n5970), .ZN(n7707)
         );
  AND4_X1 U5553 ( .A1(n5998), .A2(n5997), .A3(n5996), .A4(n5995), .ZN(n8643)
         );
  NOR2_X1 U5554 ( .A1(n7635), .A2(n7670), .ZN(n7637) );
  NAND2_X1 U5555 ( .A1(n7476), .A2(n5948), .ZN(n7612) );
  NOR2_X1 U5556 ( .A1(n4563), .A2(n7646), .ZN(n4561) );
  AND4_X1 U5557 ( .A1(n5962), .A2(n5961), .A3(n5960), .A4(n5959), .ZN(n7473)
         );
  NAND2_X1 U5558 ( .A1(n6267), .A2(n6266), .ZN(n7478) );
  AND2_X1 U5559 ( .A1(n6264), .A2(n7477), .ZN(n7552) );
  NAND2_X1 U5560 ( .A1(n5795), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5941) );
  NOR2_X1 U5561 ( .A1(n7216), .A2(n4562), .ZN(n7560) );
  INV_X1 U5562 ( .A(n4564), .ZN(n4562) );
  NOR2_X1 U5563 ( .A1(n7216), .A2(n7221), .ZN(n7217) );
  OR2_X1 U5564 ( .A1(n9852), .A2(n7312), .ZN(n7505) );
  OR2_X1 U5565 ( .A1(n6419), .A2(n7197), .ZN(n6938) );
  AND2_X1 U5566 ( .A1(n9848), .A2(n6936), .ZN(n9882) );
  AND2_X1 U5567 ( .A1(n9842), .A2(n6450), .ZN(n9837) );
  AND2_X1 U5568 ( .A1(n6189), .A2(n6216), .ZN(n4833) );
  NOR2_X1 U5569 ( .A1(n4917), .A2(P2_IR_REG_28__SCAN_IN), .ZN(n4916) );
  INV_X1 U5570 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5790) );
  NAND2_X1 U5571 ( .A1(n6408), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6397) );
  NAND2_X1 U5572 ( .A1(n6187), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6047) );
  AND2_X1 U5573 ( .A1(n5775), .A2(n6014), .ZN(n4832) );
  OR2_X1 U5574 ( .A1(n5913), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n5925) );
  AND2_X1 U5575 ( .A1(n5113), .A2(n9020), .ZN(n4682) );
  AND2_X1 U5576 ( .A1(n4684), .A2(n5137), .ZN(n4683) );
  INV_X1 U5577 ( .A(n5087), .ZN(n4686) );
  NAND2_X1 U5578 ( .A1(n5381), .A2(n5380), .ZN(n7983) );
  AND2_X1 U5579 ( .A1(n5379), .A2(n5378), .ZN(n5380) );
  AND2_X1 U5580 ( .A1(n5062), .A2(n5060), .ZN(n6875) );
  OR2_X1 U5581 ( .A1(n5059), .A2(n5058), .ZN(n5060) );
  AOI21_X1 U5582 ( .B1(n4487), .B2(n4481), .A(n4480), .ZN(n4479) );
  NOR2_X1 U5583 ( .A1(n4696), .A2(n8978), .ZN(n4481) );
  OAI21_X1 U5584 ( .B1(n4696), .B2(n4482), .A(n4415), .ZN(n4480) );
  AND2_X1 U5585 ( .A1(n5340), .A2(n4497), .ZN(n4496) );
  NAND2_X1 U5586 ( .A1(n9018), .A2(n5087), .ZN(n7228) );
  INV_X1 U5587 ( .A(n9011), .ZN(n4482) );
  NAND2_X1 U5588 ( .A1(n4487), .A2(n4486), .ZN(n4483) );
  NAND2_X1 U5589 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5090) );
  NAND2_X1 U5590 ( .A1(n9019), .A2(n9020), .ZN(n9018) );
  INV_X1 U5591 ( .A(n9031), .ZN(n4478) );
  AND2_X1 U5592 ( .A1(n5372), .A2(n5373), .ZN(n8010) );
  OR2_X1 U5593 ( .A1(n5335), .A2(n5315), .ZN(n5356) );
  NAND2_X1 U5594 ( .A1(n5270), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5333) );
  INV_X1 U5595 ( .A(n6777), .ZN(n5014) );
  NAND2_X1 U5596 ( .A1(n8159), .A2(n5470), .ZN(n4681) );
  NAND2_X1 U5597 ( .A1(n4681), .A2(n5494), .ZN(n9054) );
  OR2_X1 U5599 ( .A1(n9607), .A2(n9608), .ZN(n9609) );
  NAND2_X1 U5600 ( .A1(n6849), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4506) );
  NOR2_X1 U5601 ( .A1(n7768), .A2(n7769), .ZN(n7883) );
  NAND2_X1 U5602 ( .A1(n8286), .A2(n8285), .ZN(n9111) );
  AND2_X1 U5603 ( .A1(n9163), .A2(n5754), .ZN(n9180) );
  AOI21_X1 U5604 ( .B1(n4848), .B2(n4854), .A(n4847), .ZN(n4846) );
  AND2_X1 U5605 ( .A1(n9274), .A2(n4527), .ZN(n9206) );
  AND2_X1 U5606 ( .A1(n4528), .A2(n9210), .ZN(n4527) );
  NAND2_X1 U5607 ( .A1(n9274), .A2(n4528), .ZN(n9223) );
  NAND2_X1 U5608 ( .A1(n5613), .A2(n5612), .ZN(n5632) );
  INV_X1 U5609 ( .A(n5616), .ZN(n5613) );
  OR2_X1 U5610 ( .A1(n9407), .A2(n9244), .ZN(n9240) );
  AND2_X1 U5611 ( .A1(n9240), .A2(n8468), .ZN(n9255) );
  OAI21_X1 U5612 ( .B1(n9287), .B2(n9288), .A(n9145), .ZN(n9278) );
  INV_X1 U5613 ( .A(n5531), .ZN(n5533) );
  OR2_X1 U5614 ( .A1(n5557), .A2(n5556), .ZN(n5616) );
  NAND2_X1 U5615 ( .A1(n4837), .A2(n4835), .ZN(n9308) );
  AOI21_X1 U5616 ( .B1(n4838), .B2(n4840), .A(n4836), .ZN(n4835) );
  INV_X1 U5617 ( .A(n9142), .ZN(n4836) );
  NOR2_X1 U5618 ( .A1(n9316), .A2(n9420), .ZN(n9302) );
  INV_X1 U5619 ( .A(n4841), .ZN(n4840) );
  AOI21_X1 U5620 ( .B1(n4843), .B2(n9140), .A(n4842), .ZN(n4841) );
  INV_X1 U5621 ( .A(n9323), .ZN(n4842) );
  INV_X1 U5622 ( .A(n4839), .ZN(n4838) );
  OAI21_X1 U5623 ( .B1(n4840), .B2(n4843), .A(n9322), .ZN(n4839) );
  AND2_X1 U5624 ( .A1(n8471), .A2(n9142), .ZN(n9322) );
  NAND2_X1 U5625 ( .A1(n5456), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n5485) );
  INV_X1 U5626 ( .A(n5458), .ZN(n5456) );
  NOR2_X1 U5627 ( .A1(n9353), .A2(n9432), .ZN(n9333) );
  OAI21_X1 U5628 ( .B1(n9138), .B2(n9137), .A(n9546), .ZN(n9536) );
  INV_X1 U5629 ( .A(n5398), .ZN(n5396) );
  OR2_X1 U5630 ( .A1(n5427), .A2(n7896), .ZN(n5458) );
  AND2_X1 U5631 ( .A1(n4373), .A2(n9565), .ZN(n4532) );
  NAND2_X1 U5632 ( .A1(n4863), .A2(n4865), .ZN(n8050) );
  AOI21_X1 U5633 ( .B1(n4867), .B2(n4869), .A(n4866), .ZN(n4865) );
  AND2_X1 U5634 ( .A1(n8419), .A2(n8341), .ZN(n8487) );
  NAND2_X1 U5635 ( .A1(n7788), .A2(n4533), .ZN(n7966) );
  NAND2_X1 U5636 ( .A1(n7788), .A2(n7793), .ZN(n7916) );
  AND2_X1 U5637 ( .A1(n9506), .A2(n9582), .ZN(n7788) );
  NAND2_X1 U5638 ( .A1(n4856), .A2(n4855), .ZN(n7781) );
  AOI21_X1 U5639 ( .B1(n4858), .B2(n4861), .A(n8331), .ZN(n4855) );
  OR2_X1 U5640 ( .A1(n7534), .A2(n4857), .ZN(n4856) );
  INV_X1 U5641 ( .A(n4858), .ZN(n4857) );
  NAND2_X1 U5642 ( .A1(n4862), .A2(n4860), .ZN(n9493) );
  NAND2_X1 U5643 ( .A1(n5216), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n5249) );
  OR2_X1 U5644 ( .A1(n5249), .A2(n6692), .ZN(n5272) );
  NAND2_X1 U5645 ( .A1(n4585), .A2(n7724), .ZN(n9491) );
  OR2_X1 U5646 ( .A1(n9786), .A2(n9497), .ZN(n7724) );
  NOR2_X1 U5647 ( .A1(n7725), .A2(n4589), .ZN(n4588) );
  NAND2_X1 U5648 ( .A1(n4536), .A2(n4382), .ZN(n9505) );
  NAND2_X1 U5649 ( .A1(n4862), .A2(n8317), .ZN(n7730) );
  NAND2_X1 U5650 ( .A1(n4536), .A2(n4535), .ZN(n7540) );
  AND2_X1 U5651 ( .A1(n8317), .A2(n8436), .ZN(n8479) );
  OR2_X1 U5652 ( .A1(n7415), .A2(n7417), .ZN(n7419) );
  INV_X1 U5653 ( .A(n4591), .ZN(n4590) );
  NOR2_X1 U5654 ( .A1(n7185), .A2(n4537), .ZN(n7423) );
  NAND2_X1 U5655 ( .A1(n7296), .A2(n7295), .ZN(n7297) );
  INV_X1 U5656 ( .A(n7294), .ZN(n7295) );
  AOI22_X1 U5657 ( .A1(n5506), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n9601), .B2(
        n9652), .ZN(n5131) );
  NOR2_X1 U5658 ( .A1(n7185), .A2(n7328), .ZN(n7284) );
  INV_X1 U5659 ( .A(n9086), .ZN(n7180) );
  INV_X1 U5660 ( .A(n9084), .ZN(n7413) );
  NAND2_X1 U5661 ( .A1(n7380), .A2(n6894), .ZN(n6895) );
  NAND2_X1 U5662 ( .A1(n8294), .A2(n8293), .ZN(n9370) );
  NAND2_X1 U5663 ( .A1(n5584), .A2(n5583), .ZN(n9410) );
  NAND2_X1 U5664 ( .A1(n5453), .A2(n5452), .ZN(n9435) );
  OR2_X1 U5665 ( .A1(n7044), .A2(n7043), .ZN(n9787) );
  XNOR2_X1 U5666 ( .A(n6197), .B(SI_30_), .ZN(n8554) );
  XNOR2_X1 U5667 ( .A(n6181), .B(n6168), .ZN(n8390) );
  OAI21_X1 U5668 ( .B1(n5680), .B2(n5679), .A(n5701), .ZN(n7922) );
  AOI21_X1 U5669 ( .B1(n5264), .B2(n4721), .A(n4372), .ZN(n5385) );
  INV_X1 U5670 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5311) );
  NAND2_X1 U5671 ( .A1(n5150), .A2(n4702), .ZN(n5246) );
  NAND2_X1 U5672 ( .A1(n5208), .A2(n5207), .ZN(n5236) );
  NAND2_X1 U5673 ( .A1(n5180), .A2(n5179), .ZN(n5186) );
  INV_X1 U5674 ( .A(n4920), .ZN(n4493) );
  XNOR2_X1 U5675 ( .A(n5098), .B(SI_4_), .ZN(n5102) );
  NAND2_X1 U5676 ( .A1(n5074), .A2(n5073), .ZN(n5105) );
  NAND2_X1 U5677 ( .A1(n4514), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5018) );
  INV_X1 U5678 ( .A(n5016), .ZN(n4514) );
  NAND2_X1 U5679 ( .A1(n5018), .A2(n5017), .ZN(n5043) );
  NAND2_X1 U5680 ( .A1(n4781), .A2(n8270), .ZN(n8561) );
  NAND2_X1 U5681 ( .A1(n7940), .A2(n6169), .ZN(n6138) );
  NAND2_X1 U5682 ( .A1(n4803), .A2(n4804), .ZN(n7832) );
  NOR2_X1 U5683 ( .A1(n6996), .A2(n6995), .ZN(n7145) );
  OR2_X1 U5684 ( .A1(n8627), .A2(n8828), .ZN(n8602) );
  AND2_X1 U5685 ( .A1(n8176), .A2(n8175), .ZN(n8244) );
  AND2_X1 U5686 ( .A1(n4782), .A2(n4786), .ZN(n4775) );
  OAI22_X1 U5687 ( .A1(n4778), .A2(n4777), .B1(n4786), .B2(n4780), .ZN(n4776)
         );
  NOR2_X1 U5688 ( .A1(n4782), .A2(n4786), .ZN(n4778) );
  INV_X1 U5689 ( .A(n4780), .ZN(n4777) );
  NAND2_X1 U5690 ( .A1(n4780), .A2(n8278), .ZN(n4779) );
  NAND2_X1 U5691 ( .A1(n4773), .A2(n6954), .ZN(n4772) );
  OAI22_X1 U5692 ( .A1(n6950), .A2(n8271), .B1(n9847), .B2(n6957), .ZN(n6981)
         );
  NAND2_X1 U5693 ( .A1(n4826), .A2(n4827), .ZN(n8577) );
  NAND2_X1 U5694 ( .A1(n8176), .A2(n4828), .ZN(n4826) );
  NAND2_X1 U5695 ( .A1(n7136), .A2(n7003), .ZN(n7027) );
  NAND2_X1 U5696 ( .A1(n6105), .A2(n6104), .ZN(n8891) );
  NOR2_X1 U5697 ( .A1(n8244), .A2(n8243), .ZN(n8601) );
  NAND2_X1 U5698 ( .A1(n6062), .A2(n6061), .ZN(n8913) );
  INV_X1 U5699 ( .A(n4817), .ZN(n7699) );
  AOI21_X1 U5700 ( .B1(n7370), .B2(n4819), .A(n4821), .ZN(n4817) );
  NOR2_X1 U5701 ( .A1(n6961), .A2(n6960), .ZN(n6996) );
  OAI22_X1 U5702 ( .A1(n8131), .A2(n8130), .B1(n8129), .B2(n8128), .ZN(n8172)
         );
  INV_X1 U5703 ( .A(n8625), .ZN(n8615) );
  OR2_X1 U5704 ( .A1(n6544), .A2(n7013), .ZN(n8638) );
  NAND4_X1 U5705 ( .A1(n5896), .A2(n5895), .A3(n5894), .A4(n5893), .ZN(n8653)
         );
  OR2_X1 U5706 ( .A1(n5888), .A2(n5887), .ZN(n5896) );
  OR2_X1 U5707 ( .A1(n5875), .A2(n5861), .ZN(n5867) );
  NOR2_X1 U5708 ( .A1(n6806), .A2(n4432), .ZN(n6810) );
  INV_X1 U5709 ( .A(n4652), .ZN(n6820) );
  AND2_X1 U5710 ( .A1(n4652), .A2(n4651), .ZN(n6824) );
  NAND2_X1 U5711 ( .A1(n6821), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n4651) );
  INV_X1 U5712 ( .A(n4649), .ZN(n6867) );
  INV_X1 U5713 ( .A(n6918), .ZN(n4645) );
  INV_X1 U5714 ( .A(n4646), .ZN(n6919) );
  AOI21_X1 U5715 ( .B1(P2_REG2_REG_10__SCAN_IN), .B2(n7113), .A(n4396), .ZN(
        n7110) );
  NOR2_X1 U5716 ( .A1(n7517), .A2(n4657), .ZN(n7520) );
  AND2_X1 U5717 ( .A1(n7518), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n4657) );
  NAND2_X1 U5718 ( .A1(n7520), .A2(n7519), .ZN(n7679) );
  NAND2_X1 U5719 ( .A1(n7679), .A2(n4656), .ZN(n7680) );
  OR2_X1 U5720 ( .A1(n7684), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n4656) );
  AND2_X1 U5721 ( .A1(n4654), .A2(n4653), .ZN(n8658) );
  INV_X1 U5722 ( .A(n8659), .ZN(n4653) );
  INV_X1 U5723 ( .A(n4654), .ZN(n8660) );
  NAND2_X1 U5724 ( .A1(n6208), .A2(n6207), .ZN(n8860) );
  OR2_X1 U5725 ( .A1(n8726), .A2(n4765), .ZN(n8717) );
  NAND2_X1 U5726 ( .A1(n6116), .A2(n6115), .ZN(n8887) );
  NAND2_X1 U5727 ( .A1(n7812), .A2(n6169), .ZN(n6116) );
  AND2_X1 U5728 ( .A1(n4908), .A2(n4907), .ZN(n8740) );
  NAND2_X1 U5729 ( .A1(n8898), .A2(n4921), .ZN(n8758) );
  NOR2_X1 U5730 ( .A1(n8771), .A2(n6103), .ZN(n8764) );
  NAND2_X1 U5731 ( .A1(n8798), .A2(n6322), .ZN(n8772) );
  INV_X1 U5732 ( .A(n4553), .ZN(n8790) );
  NAND2_X1 U5733 ( .A1(n4738), .A2(n4736), .ZN(n8826) );
  NAND2_X1 U5734 ( .A1(n6052), .A2(n6051), .ZN(n8920) );
  OAI21_X1 U5735 ( .B1(n8837), .B2(n6297), .A(n6363), .ZN(n8152) );
  NAND2_X1 U5736 ( .A1(n4915), .A2(n4375), .ZN(n8029) );
  AND2_X1 U5737 ( .A1(n4915), .A2(n4914), .ZN(n8031) );
  OAI21_X1 U5738 ( .B1(n7803), .B2(n4756), .A(n4753), .ZN(n7945) );
  INV_X1 U5739 ( .A(n4757), .ZN(n4756) );
  NAND2_X1 U5740 ( .A1(n7807), .A2(n4759), .ZN(n7842) );
  NAND2_X1 U5741 ( .A1(n4895), .A2(n4896), .ZN(n7739) );
  AND2_X1 U5742 ( .A1(n4892), .A2(n4899), .ZN(n4895) );
  NOR2_X1 U5743 ( .A1(n7471), .A2(n6431), .ZN(n4897) );
  AND2_X1 U5744 ( .A1(n7209), .A2(n6259), .ZN(n7126) );
  NAND2_X1 U5745 ( .A1(n4911), .A2(n6426), .ZN(n7224) );
  INV_X1 U5746 ( .A(n4470), .ZN(n4469) );
  OAI21_X1 U5747 ( .B1(n4392), .B2(n6622), .A(n4471), .ZN(n4470) );
  INV_X1 U5748 ( .A(n8851), .ZN(n8755) );
  NAND2_X1 U5749 ( .A1(n4546), .A2(n4543), .ZN(n8949) );
  NAND2_X1 U5750 ( .A1(n8868), .A2(n9883), .ZN(n4546) );
  XNOR2_X1 U5751 ( .A(n5810), .B(n5809), .ZN(n8240) );
  NAND2_X1 U5752 ( .A1(n5808), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5810) );
  OAI21_X1 U5753 ( .B1(n6410), .B2(P2_IR_REG_26__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5806) );
  XNOR2_X1 U5754 ( .A(n6397), .B(n6405), .ZN(n7433) );
  XNOR2_X1 U5755 ( .A(n6191), .B(n6216), .ZN(n7171) );
  INV_X1 U5756 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n10082) );
  INV_X1 U5757 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n10073) );
  INV_X1 U5758 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6609) );
  MUX2_X1 U5759 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5855), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n5857) );
  INV_X1 U5760 ( .A(n9083), .ZN(n7409) );
  AND2_X1 U5761 ( .A1(n5720), .A2(n5721), .ZN(n5748) );
  NAND2_X1 U5762 ( .A1(n5706), .A2(n5705), .ZN(n9385) );
  INV_X1 U5763 ( .A(n9080), .ZN(n7988) );
  AND2_X1 U5764 ( .A1(n7981), .A2(n7979), .ZN(n5376) );
  NAND2_X1 U5765 ( .A1(n7655), .A2(n5235), .ZN(n7715) );
  OR2_X1 U5766 ( .A1(n5494), .A2(n4680), .ZN(n4678) );
  NAND2_X1 U5767 ( .A1(n8159), .A2(n4675), .ZN(n4674) );
  NOR2_X1 U5768 ( .A1(n4679), .A2(n4676), .ZN(n4675) );
  NAND2_X1 U5769 ( .A1(n5508), .A2(n5507), .ZN(n9425) );
  NAND2_X1 U5770 ( .A1(n6486), .A2(n6485), .ZN(n9179) );
  NAND2_X1 U5771 ( .A1(n6484), .A2(n8389), .ZN(n6486) );
  OAI21_X1 U5772 ( .B1(n4526), .B2(n4380), .A(n5042), .ZN(n4525) );
  NAND2_X1 U5773 ( .A1(n9028), .A2(n9032), .ZN(n8996) );
  NAND2_X1 U5774 ( .A1(n5555), .A2(n5554), .ZN(n9417) );
  CLKBUF_X1 U5775 ( .A(n7817), .Z(n7818) );
  CLKBUF_X1 U5776 ( .A(n9073), .Z(n9037) );
  NAND2_X1 U5777 ( .A1(n9054), .A2(n9053), .ZN(n9052) );
  INV_X1 U5778 ( .A(n9079), .ZN(n8052) );
  NAND2_X1 U5779 ( .A1(n4565), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4976) );
  NAND2_X1 U5780 ( .A1(n4523), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4977) );
  INV_X1 U5781 ( .A(n4873), .ZN(n4604) );
  NAND2_X1 U5782 ( .A1(n4567), .A2(n4566), .ZN(n8510) );
  INV_X1 U5783 ( .A(n4569), .ZN(n8506) );
  NAND4_X1 U5784 ( .A1(n5041), .A2(n5040), .A3(n5039), .A4(n5038), .ZN(n9088)
         );
  NAND4_X1 U5785 ( .A1(n6891), .A2(n6890), .A3(n6889), .A4(n6888), .ZN(n9712)
         );
  NAND2_X1 U5786 ( .A1(n5114), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5002) );
  CLKBUF_X1 U5787 ( .A(P1_IR_REG_0__SCAN_IN), .Z(n9949) );
  NAND2_X1 U5788 ( .A1(n9627), .A2(n9628), .ZN(n9626) );
  NOR2_X1 U5789 ( .A1(n9645), .A2(n4394), .ZN(n6734) );
  INV_X1 U5790 ( .A(n4511), .ZN(n9658) );
  INV_X1 U5791 ( .A(n4509), .ZN(n6705) );
  INV_X1 U5792 ( .A(n4507), .ZN(n6848) );
  XNOR2_X1 U5793 ( .A(n7767), .B(n7766), .ZN(n7405) );
  NOR2_X1 U5794 ( .A1(n7405), .A2(n7404), .ZN(n7768) );
  INV_X1 U5795 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5477) );
  INV_X1 U5796 ( .A(n9370), .ZN(n9107) );
  AND2_X1 U5797 ( .A1(n9172), .A2(n9171), .ZN(n9378) );
  NAND2_X1 U5798 ( .A1(n4850), .A2(n4851), .ZN(n9195) );
  OR2_X1 U5799 ( .A1(n9238), .A2(n4854), .ZN(n4850) );
  NAND2_X1 U5800 ( .A1(n9212), .A2(n4853), .ZN(n9213) );
  OAI21_X1 U5801 ( .B1(n9237), .B2(n4598), .A(n4596), .ZN(n9204) );
  AND2_X1 U5802 ( .A1(n4601), .A2(n4602), .ZN(n9222) );
  NAND2_X1 U5803 ( .A1(n9237), .A2(n9130), .ZN(n4601) );
  OAI21_X1 U5804 ( .B1(n9123), .B2(n4625), .A(n4622), .ZN(n9273) );
  NAND2_X1 U5805 ( .A1(n4626), .A2(n4624), .ZN(n9285) );
  AND2_X1 U5806 ( .A1(n4626), .A2(n4379), .ZN(n9286) );
  NAND2_X1 U5807 ( .A1(n9123), .A2(n9122), .ZN(n4626) );
  NAND2_X1 U5808 ( .A1(n4628), .A2(n4633), .ZN(n9351) );
  NAND2_X1 U5809 ( .A1(n9115), .A2(n4635), .ZN(n4628) );
  NAND2_X1 U5810 ( .A1(n5426), .A2(n5425), .ZN(n9544) );
  NAND2_X1 U5811 ( .A1(n4639), .A2(n4641), .ZN(n9545) );
  NAND2_X1 U5812 ( .A1(n9115), .A2(n4384), .ZN(n4639) );
  NAND2_X1 U5813 ( .A1(n5314), .A2(n5313), .ZN(n7959) );
  NAND2_X1 U5814 ( .A1(n4605), .A2(n4609), .ZN(n7958) );
  NAND2_X1 U5815 ( .A1(n7780), .A2(n4611), .ZN(n4605) );
  OAI21_X1 U5816 ( .B1(n7780), .B2(n4391), .A(n7779), .ZN(n7906) );
  NAND2_X1 U5817 ( .A1(n5269), .A2(n5268), .ZN(n7782) );
  NAND2_X1 U5818 ( .A1(n5248), .A2(n5247), .ZN(n9504) );
  OR2_X1 U5819 ( .A1(n4587), .A2(n4593), .ZN(n7726) );
  NAND2_X1 U5820 ( .A1(n4591), .A2(n7536), .ZN(n4587) );
  INV_X1 U5821 ( .A(n7296), .ZN(n7293) );
  INV_X1 U5822 ( .A(n9806), .ZN(n9803) );
  OAI211_X1 U5823 ( .C1(n9788), .C2(n9374), .A(n9377), .B(n4408), .ZN(n9443)
         );
  AND2_X1 U5824 ( .A1(n9376), .A2(n9436), .ZN(n4539) );
  INV_X1 U5825 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n4942) );
  XNOR2_X1 U5826 ( .A(n6161), .B(n6160), .ZN(n6484) );
  XNOR2_X1 U5827 ( .A(n6142), .B(n6143), .ZN(n7940) );
  INV_X1 U5828 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n10148) );
  INV_X1 U5829 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6618) );
  NAND2_X1 U5830 ( .A1(n4834), .A2(n5016), .ZN(n5069) );
  XNOR2_X1 U5831 ( .A(n4513), .B(n5044), .ZN(n6710) );
  NAND2_X1 U5832 ( .A1(n5043), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4513) );
  INV_X1 U5833 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6606) );
  NAND2_X1 U5834 ( .A1(n7059), .A2(n7011), .ZN(n7072) );
  OAI21_X1 U5835 ( .B1(n7060), .B2(n4793), .A(n4791), .ZN(n7346) );
  AOI21_X1 U5836 ( .B1(n9813), .B2(P2_ADDR_REG_19__SCAN_IN), .A(n8239), .ZN(
        n4662) );
  NAND2_X1 U5837 ( .A1(n4668), .A2(n9827), .ZN(n4667) );
  INV_X1 U5838 ( .A(n4664), .ZN(n4663) );
  NAND2_X1 U5839 ( .A1(n4542), .A2(n4541), .ZN(P2_U3517) );
  NAND2_X1 U5840 ( .A1(n9907), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n4541) );
  NAND2_X1 U5841 ( .A1(n8949), .A2(n9909), .ZN(n4542) );
  AOI21_X1 U5842 ( .B1(n9668), .B2(P1_ADDR_REG_19__SCAN_IN), .A(n9102), .ZN(
        n4517) );
  NAND2_X1 U5843 ( .A1(n4516), .A2(n5505), .ZN(n4515) );
  NAND2_X1 U5844 ( .A1(n4519), .A2(n4989), .ZN(n4518) );
  NAND2_X1 U5845 ( .A1(n4377), .A2(n4697), .ZN(n4696) );
  AND2_X1 U5846 ( .A1(n5350), .A2(n5349), .ZN(n4372) );
  AND2_X1 U5847 ( .A1(n4533), .A2(n9572), .ZN(n4373) );
  NOR2_X1 U5848 ( .A1(n7419), .A2(n8479), .ZN(n4374) );
  INV_X2 U5849 ( .A(n5055), .ZN(n6490) );
  AND2_X1 U5850 ( .A1(n8030), .A2(n4914), .ZN(n4375) );
  INV_X1 U5851 ( .A(n5239), .ZN(n5601) );
  OR2_X1 U5852 ( .A1(n4801), .A2(n8037), .ZN(n4376) );
  AND2_X1 U5853 ( .A1(n4433), .A2(n5671), .ZN(n4377) );
  NAND2_X1 U5854 ( .A1(n6334), .A2(n6135), .ZN(n6446) );
  AND2_X1 U5855 ( .A1(n4559), .A2(n7802), .ZN(n4378) );
  OR2_X1 U5856 ( .A1(n9420), .A2(n9327), .ZN(n4379) );
  INV_X1 U5857 ( .A(n6957), .ZN(n8247) );
  AOI21_X1 U5858 ( .B1(n8711), .B2(n5848), .A(n6141), .ZN(n8702) );
  AND2_X1 U5859 ( .A1(n6607), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4380) );
  OR2_X1 U5860 ( .A1(n8233), .A2(n4644), .ZN(n4381) );
  NAND2_X1 U5861 ( .A1(n5977), .A2(n5976), .ZN(n7700) );
  AND2_X1 U5862 ( .A1(n4535), .A2(n4538), .ZN(n4382) );
  AND2_X1 U5863 ( .A1(n8860), .A2(n6209), .ZN(n6355) );
  AND2_X1 U5864 ( .A1(n4844), .A2(n4843), .ZN(n4383) );
  INV_X1 U5865 ( .A(n4861), .ZN(n4860) );
  NAND2_X1 U5866 ( .A1(n8316), .A2(n8317), .ZN(n4861) );
  INV_X1 U5867 ( .A(n4869), .ZN(n4868) );
  INV_X1 U5868 ( .A(n4829), .ZN(n4828) );
  NAND2_X1 U5869 ( .A1(n4390), .A2(n8175), .ZN(n4829) );
  OR2_X1 U5870 ( .A1(n9565), .A2(n9116), .ZN(n4384) );
  NAND2_X1 U5871 ( .A1(n6999), .A2(n6998), .ZN(n4385) );
  AND2_X1 U5872 ( .A1(n4548), .A2(n4547), .ZN(n4386) );
  AND2_X1 U5873 ( .A1(n4898), .A2(n4899), .ZN(n4387) );
  NAND2_X1 U5874 ( .A1(n4379), .A2(n9288), .ZN(n4625) );
  NAND2_X1 U5875 ( .A1(n5353), .A2(n5352), .ZN(n8048) );
  INV_X1 U5876 ( .A(n6227), .ZN(n4754) );
  NAND2_X1 U5877 ( .A1(n4810), .A2(n4809), .ZN(n7136) );
  INV_X1 U5878 ( .A(n7087), .ZN(n6388) );
  AND2_X1 U5879 ( .A1(n6347), .A2(n6346), .ZN(n6467) );
  AND3_X1 U5880 ( .A1(n5094), .A2(n5093), .A3(n5092), .ZN(n4388) );
  NAND2_X1 U5881 ( .A1(n4485), .A2(n4484), .ZN(n4487) );
  NAND2_X1 U5882 ( .A1(n5779), .A2(n5778), .ZN(n5811) );
  NAND2_X1 U5883 ( .A1(n6157), .A2(n6156), .ZN(n8634) );
  NOR2_X1 U5884 ( .A1(n7221), .A2(n8651), .ZN(n4389) );
  OR2_X1 U5885 ( .A1(n8913), .A2(n8579), .ZN(n6316) );
  NAND2_X1 U5886 ( .A1(n8246), .A2(n8245), .ZN(n4390) );
  INV_X1 U5887 ( .A(n7433), .ZN(n6219) );
  NOR2_X1 U5888 ( .A1(n7782), .A2(n9496), .ZN(n4391) );
  NAND2_X1 U5889 ( .A1(n6565), .A2(n6607), .ZN(n4392) );
  NAND2_X1 U5890 ( .A1(n5150), .A2(n4701), .ZN(n4393) );
  AND2_X1 U5891 ( .A1(n9652), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n4394) );
  OAI21_X1 U5892 ( .B1(n8591), .B2(n8592), .A(n8262), .ZN(n8584) );
  XNOR2_X1 U5893 ( .A(n5791), .B(n5790), .ZN(n5792) );
  AND2_X1 U5894 ( .A1(n6492), .A2(n4499), .ZN(n4395) );
  AND2_X1 U5895 ( .A1(n4646), .A2(n4645), .ZN(n4396) );
  NAND2_X1 U5896 ( .A1(n5739), .A2(n8543), .ZN(n4987) );
  OR3_X1 U5897 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .A3(
        P2_IR_REG_0__SCAN_IN), .ZN(n4397) );
  NAND2_X1 U5898 ( .A1(n5150), .A2(n4954), .ZN(n5188) );
  AND3_X1 U5899 ( .A1(n6351), .A2(n6348), .A3(n6350), .ZN(n4399) );
  XNOR2_X1 U5900 ( .A(n5178), .B(SI_7_), .ZN(n5176) );
  AND3_X1 U5901 ( .A1(n5774), .A2(n5773), .A3(n5778), .ZN(n4400) );
  INV_X1 U5902 ( .A(n8278), .ZN(n4786) );
  NAND2_X1 U5903 ( .A1(n5529), .A2(n5528), .ZN(n9420) );
  NAND2_X1 U5904 ( .A1(n4498), .A2(n5332), .ZN(n7930) );
  AND2_X1 U5905 ( .A1(n4721), .A2(n5382), .ZN(n4401) );
  OR2_X1 U5906 ( .A1(n8811), .A2(n8831), .ZN(n4402) );
  AND2_X1 U5907 ( .A1(n4507), .A2(n4506), .ZN(n4403) );
  OR2_X1 U5908 ( .A1(n8726), .A2(n6136), .ZN(n4404) );
  NAND2_X1 U5909 ( .A1(n4478), .A2(n4925), .ZN(n9028) );
  NOR2_X1 U5910 ( .A1(n8233), .A2(n4643), .ZN(n4405) );
  NAND2_X1 U5911 ( .A1(n8750), .A2(n4550), .ZN(n4551) );
  NAND2_X1 U5912 ( .A1(n5989), .A2(n5988), .ZN(n7763) );
  INV_X1 U5913 ( .A(n8871), .ZN(n6158) );
  NAND2_X1 U5914 ( .A1(n6146), .A2(n6145), .ZN(n8871) );
  AND2_X1 U5915 ( .A1(n6439), .A2(n8132), .ZN(n4406) );
  OR2_X1 U5916 ( .A1(n8887), .A2(n8263), .ZN(n8723) );
  NAND2_X1 U5917 ( .A1(n9391), .A2(n9131), .ZN(n9150) );
  INV_X1 U5918 ( .A(n8049), .ZN(n4867) );
  NOR2_X1 U5919 ( .A1(n8060), .A2(n8062), .ZN(n4407) );
  NOR2_X1 U5920 ( .A1(n9375), .A2(n4539), .ZN(n4408) );
  INV_X1 U5921 ( .A(n7960), .ZN(n4615) );
  NAND2_X1 U5922 ( .A1(n9576), .A2(n7988), .ZN(n7960) );
  INV_X1 U5923 ( .A(n7904), .ZN(n4616) );
  INV_X1 U5924 ( .A(n8883), .ZN(n6476) );
  NAND2_X1 U5925 ( .A1(n6125), .A2(n6124), .ZN(n8883) );
  OR2_X1 U5926 ( .A1(n4967), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n4409) );
  INV_X1 U5927 ( .A(n4703), .ZN(n4702) );
  NAND2_X1 U5928 ( .A1(n4954), .A2(n4704), .ZN(n4703) );
  NAND2_X1 U5929 ( .A1(n5601), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n4410) );
  AND2_X1 U5930 ( .A1(n7359), .A2(n6234), .ZN(n4411) );
  NOR2_X1 U5931 ( .A1(n9395), .A2(n9216), .ZN(n4412) );
  NOR2_X1 U5932 ( .A1(n8249), .A2(n8248), .ZN(n4413) );
  NAND2_X1 U5933 ( .A1(n8467), .A2(n9150), .ZN(n9203) );
  INV_X1 U5934 ( .A(n9203), .ZN(n9214) );
  INV_X1 U5935 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n10084) );
  INV_X1 U5936 ( .A(n9119), .ZN(n4640) );
  AND2_X1 U5937 ( .A1(n9544), .A2(n9361), .ZN(n9119) );
  NOR2_X1 U5938 ( .A1(n8887), .A2(n8767), .ZN(n4414) );
  AND2_X1 U5939 ( .A1(n4698), .A2(n4699), .ZN(n4415) );
  AND2_X1 U5940 ( .A1(n4488), .A2(n4706), .ZN(n4416) );
  NAND2_X1 U5941 ( .A1(n9410), .A2(n9258), .ZN(n4417) );
  AND2_X1 U5942 ( .A1(n5384), .A2(SI_14_), .ZN(n4418) );
  NAND2_X1 U5943 ( .A1(n8335), .A2(n8484), .ZN(n4419) );
  NAND2_X1 U5944 ( .A1(n7343), .A2(n7344), .ZN(n4420) );
  NAND2_X1 U5945 ( .A1(n6183), .A2(n6182), .ZN(n8688) );
  NOR2_X1 U5946 ( .A1(n9298), .A2(n9124), .ZN(n4421) );
  AND2_X1 U5947 ( .A1(n7959), .A2(n9080), .ZN(n4422) );
  OAI21_X1 U5948 ( .B1(n4821), .B2(n4819), .A(n7698), .ZN(n4818) );
  AND2_X1 U5949 ( .A1(n8273), .A2(n8272), .ZN(n4423) );
  INV_X1 U5950 ( .A(n4625), .ZN(n4624) );
  NAND2_X1 U5951 ( .A1(n6360), .A2(n4745), .ZN(n4424) );
  OR2_X1 U5952 ( .A1(n9504), .A2(n7821), .ZN(n8329) );
  AND2_X1 U5953 ( .A1(n4790), .A2(n7345), .ZN(n4425) );
  AND2_X1 U5954 ( .A1(n8869), .A2(n4544), .ZN(n4426) );
  AND2_X1 U5955 ( .A1(n8522), .A2(n8518), .ZN(n4427) );
  NAND2_X1 U5956 ( .A1(n5395), .A2(n5394), .ZN(n9117) );
  AND2_X1 U5957 ( .A1(n4633), .A2(n4632), .ZN(n4428) );
  NOR2_X1 U5958 ( .A1(n4873), .A2(P1_IR_REG_27__SCAN_IN), .ZN(n4872) );
  INV_X1 U5959 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n6216) );
  INV_X1 U5960 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n6014) );
  AND2_X1 U5961 ( .A1(n4457), .A2(n4453), .ZN(n4429) );
  AND2_X1 U5962 ( .A1(n4851), .A2(n4849), .ZN(n4848) );
  INV_X1 U5963 ( .A(n4824), .ZN(n4823) );
  NAND2_X1 U5964 ( .A1(n4827), .A2(n4825), .ZN(n4824) );
  AND2_X2 U5965 ( .A1(n5792), .A2(n8971), .ZN(n6030) );
  INV_X1 U5966 ( .A(n4586), .ZN(n4593) );
  NAND2_X1 U5967 ( .A1(n7783), .A2(n8486), .ZN(n7910) );
  NOR2_X1 U5968 ( .A1(n8050), .A2(n8489), .ZN(n9138) );
  INV_X1 U5969 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5813) );
  AND2_X1 U5970 ( .A1(n4797), .A2(n4376), .ZN(n4430) );
  AND2_X1 U5971 ( .A1(n7910), .A2(n4868), .ZN(n4431) );
  NAND2_X1 U5972 ( .A1(n4674), .A2(n4678), .ZN(n8985) );
  AND2_X1 U5973 ( .A1(n6807), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n4432) );
  INV_X1 U5974 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n4874) );
  AND4_X1 U5975 ( .A1(n4832), .A2(n4400), .A3(n5776), .A4(n5779), .ZN(n6036)
         );
  OR2_X1 U5976 ( .A1(n5699), .A2(n5698), .ZN(n4433) );
  NAND2_X1 U5977 ( .A1(n6073), .A2(n6072), .ZN(n8908) );
  AND2_X1 U5978 ( .A1(n6283), .A2(n5999), .ZN(n7742) );
  INV_X1 U5979 ( .A(n7742), .ZN(n4898) );
  NAND2_X1 U5980 ( .A1(n6171), .A2(n6170), .ZN(n8867) );
  INV_X1 U5981 ( .A(n8867), .ZN(n4547) );
  NAND2_X1 U5982 ( .A1(n6138), .A2(n6137), .ZN(n8876) );
  INV_X1 U5983 ( .A(n6293), .ZN(n4752) );
  AND2_X1 U5984 ( .A1(n4738), .A2(n4737), .ZN(n4434) );
  NAND2_X1 U5985 ( .A1(n9274), .A2(n4530), .ZN(n4531) );
  INV_X1 U5986 ( .A(n4677), .ZN(n9055) );
  NOR2_X1 U5987 ( .A1(n4681), .A2(n5494), .ZN(n4677) );
  AND2_X1 U5988 ( .A1(n4803), .A2(n4801), .ZN(n4435) );
  AND2_X1 U5989 ( .A1(n4639), .A2(n4637), .ZN(n4436) );
  NAND2_X1 U5990 ( .A1(n5682), .A2(n5681), .ZN(n9391) );
  INV_X1 U5991 ( .A(n9129), .ZN(n4602) );
  INV_X1 U5992 ( .A(n7804), .ZN(n4755) );
  NAND2_X1 U5993 ( .A1(n4583), .A2(n4592), .ZN(n4591) );
  NAND2_X1 U5994 ( .A1(n6904), .A2(n8518), .ZN(n7163) );
  NAND2_X1 U5995 ( .A1(n6083), .A2(n6082), .ZN(n8903) );
  INV_X1 U5996 ( .A(n8903), .ZN(n4552) );
  NAND2_X1 U5997 ( .A1(n4940), .A2(n5122), .ZN(n4437) );
  OR2_X1 U5998 ( .A1(n8048), .A2(n8052), .ZN(n8419) );
  INV_X1 U5999 ( .A(n8419), .ZN(n4866) );
  INV_X1 U6000 ( .A(n7420), .ZN(n4584) );
  NAND2_X1 U6001 ( .A1(n5262), .A2(n5261), .ZN(n4438) );
  OR2_X1 U6002 ( .A1(n4590), .A2(n4593), .ZN(n4439) );
  OR2_X1 U6003 ( .A1(n7216), .A2(n4563), .ZN(n4440) );
  NAND2_X1 U6004 ( .A1(n7788), .A2(n4373), .ZN(n4534) );
  AND2_X1 U6005 ( .A1(n4810), .A2(n4385), .ZN(n4441) );
  AND2_X1 U6006 ( .A1(n4695), .A2(n4438), .ZN(n4442) );
  NAND2_X1 U6007 ( .A1(n6219), .A2(n8734), .ZN(n6387) );
  XNOR2_X1 U6008 ( .A(n4976), .B(n4975), .ZN(n5759) );
  AND2_X1 U6009 ( .A1(n8229), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n4443) );
  NAND2_X1 U6010 ( .A1(n5215), .A2(n5214), .ZN(n9786) );
  INV_X1 U6011 ( .A(n9786), .ZN(n4538) );
  NAND2_X1 U6012 ( .A1(n6003), .A2(n6002), .ZN(n9521) );
  INV_X1 U6013 ( .A(n9521), .ZN(n4558) );
  OR2_X1 U6014 ( .A1(n8198), .A2(n7251), .ZN(n7185) );
  INV_X1 U6015 ( .A(n7185), .ZN(n4536) );
  INV_X1 U6016 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6406) );
  INV_X1 U6017 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5421) );
  XNOR2_X1 U6018 ( .A(n6214), .B(P2_IR_REG_20__SCAN_IN), .ZN(n7087) );
  INV_X1 U6019 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4504) );
  INV_X1 U6020 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n4661) );
  NOR2_X2 U6021 ( .A1(n9100), .A2(n6764), .ZN(n9686) );
  OR2_X2 U6022 ( .A1(n6525), .A2(P1_U3084), .ZN(n9089) );
  AND3_X2 U6023 ( .A1(n5016), .A2(n4834), .A3(n4444), .ZN(n5122) );
  NAND2_X1 U6024 ( .A1(n4695), .A2(n4694), .ZN(n7817) );
  NAND2_X1 U6025 ( .A1(n4673), .A2(n4672), .ZN(n9044) );
  OAI21_X1 U6026 ( .B1(n9002), .B2(n9003), .A(n5671), .ZN(n9066) );
  NAND2_X1 U6027 ( .A1(n6263), .A2(n4454), .ZN(n4452) );
  NAND2_X1 U6028 ( .A1(n4429), .A2(n4452), .ZN(n6274) );
  OAI21_X1 U6029 ( .B1(n6263), .B2(n4459), .A(n4454), .ZN(n6276) );
  NAND2_X1 U6030 ( .A1(n4366), .A2(n5785), .ZN(n6410) );
  AND2_X2 U6031 ( .A1(n6565), .A2(n5447), .ZN(n6050) );
  NAND2_X2 U6032 ( .A1(n8240), .A2(n7941), .ZN(n6565) );
  NAND2_X1 U6033 ( .A1(n9029), .A2(n9032), .ZN(n4474) );
  NAND2_X1 U6034 ( .A1(n4474), .A2(n4475), .ZN(n4673) );
  NAND2_X1 U6035 ( .A1(n4483), .A2(n8977), .ZN(n9010) );
  INV_X1 U6036 ( .A(n5627), .ZN(n4484) );
  NAND2_X1 U6037 ( .A1(n9040), .A2(n9043), .ZN(n4485) );
  INV_X1 U6038 ( .A(n8978), .ZN(n4486) );
  AND2_X1 U6039 ( .A1(n4494), .A2(n4493), .ZN(n5177) );
  NAND2_X1 U6040 ( .A1(n6688), .A2(n4395), .ZN(n4495) );
  NAND2_X1 U6041 ( .A1(n4495), .A2(n4496), .ZN(n5341) );
  NAND2_X1 U6042 ( .A1(n6688), .A2(n8389), .ZN(n4498) );
  NAND3_X1 U6043 ( .A1(n4504), .A2(n4505), .A3(n4503), .ZN(n4502) );
  NAND3_X1 U6044 ( .A1(n4518), .A2(n4517), .A3(n4515), .ZN(P1_U3260) );
  NAND2_X1 U6045 ( .A1(n4524), .A2(n4935), .ZN(n4955) );
  NAND4_X1 U6047 ( .A1(n5122), .A2(n4522), .A3(n4604), .A4(n4521), .ZN(n4523)
         );
  NAND2_X2 U6048 ( .A1(n5759), .A2(n9104), .ZN(n5042) );
  NAND2_X2 U6049 ( .A1(n5042), .A2(n6607), .ZN(n8391) );
  INV_X1 U6050 ( .A(n4531), .ZN(n9246) );
  NAND2_X1 U6051 ( .A1(n7788), .A2(n4532), .ZN(n9547) );
  INV_X1 U6052 ( .A(n4534), .ZN(n8053) );
  NOR2_X2 U6053 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5833) );
  NAND2_X1 U6054 ( .A1(n8750), .A2(n6476), .ZN(n8729) );
  INV_X1 U6055 ( .A(n4551), .ZN(n8710) );
  INV_X1 U6056 ( .A(n7216), .ZN(n4560) );
  NAND2_X1 U6057 ( .A1(n4560), .A2(n4561), .ZN(n7618) );
  XNOR2_X1 U6058 ( .A(n5011), .B(n6901), .ZN(n9716) );
  NAND2_X1 U6059 ( .A1(n4603), .A2(n4940), .ZN(n4967) );
  NAND3_X1 U6060 ( .A1(n4603), .A2(n4872), .A3(n4940), .ZN(n4565) );
  OAI22_X1 U6061 ( .A1(n8381), .A2(n9391), .B1(n8385), .B2(n8466), .ZN(n8371)
         );
  OAI21_X1 U6062 ( .B1(n4572), .B2(n4571), .A(n8370), .ZN(n8381) );
  OAI21_X1 U6063 ( .B1(n8367), .B2(n8385), .A(n8369), .ZN(n4571) );
  NOR2_X1 U6064 ( .A1(n8368), .A2(n8406), .ZN(n4572) );
  AOI21_X1 U6065 ( .B1(n4577), .B2(n4573), .A(n8338), .ZN(n8348) );
  NAND2_X2 U6066 ( .A1(n4580), .A2(n4711), .ZN(n8387) );
  NAND3_X1 U6067 ( .A1(n4586), .A2(n4591), .A3(n4588), .ZN(n4585) );
  NAND2_X1 U6068 ( .A1(n9237), .A2(n4596), .ZN(n4595) );
  OAI21_X1 U6069 ( .B1(n7780), .B2(n4608), .A(n4606), .ZN(n4614) );
  OAI21_X1 U6070 ( .B1(n9123), .B2(n4621), .A(n4618), .ZN(n4617) );
  NAND2_X1 U6071 ( .A1(n9118), .A2(n4428), .ZN(n4627) );
  NAND2_X1 U6072 ( .A1(n4627), .A2(n4629), .ZN(n9332) );
  INV_X1 U6073 ( .A(n8233), .ZN(n4642) );
  INV_X1 U6074 ( .A(n8232), .ZN(n4643) );
  NAND2_X1 U6075 ( .A1(n8232), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n4644) );
  NAND2_X1 U6076 ( .A1(n4660), .A2(n4659), .ZN(n9464) );
  NAND3_X1 U6077 ( .A1(n4667), .A2(n4663), .A3(n4662), .ZN(P2_U3264) );
  NAND3_X1 U6078 ( .A1(n5016), .A2(n4834), .A3(n4931), .ZN(n5071) );
  AND2_X2 U6079 ( .A1(n4998), .A2(n4670), .ZN(n5016) );
  NAND3_X1 U6080 ( .A1(n5412), .A2(n5438), .A3(n7994), .ZN(n8142) );
  NAND2_X1 U6081 ( .A1(n5412), .A2(n7994), .ZN(n8138) );
  NAND2_X1 U6082 ( .A1(n4673), .A2(n5572), .ZN(n5597) );
  NAND2_X1 U6083 ( .A1(n5113), .A2(n4686), .ZN(n4684) );
  NAND2_X1 U6084 ( .A1(n9019), .A2(n4682), .ZN(n4685) );
  NAND2_X1 U6085 ( .A1(n4685), .A2(n4683), .ZN(n5141) );
  NAND2_X1 U6086 ( .A1(n7656), .A2(n4688), .ZN(n4687) );
  NAND2_X1 U6087 ( .A1(n4687), .A2(n4690), .ZN(n5381) );
  NAND2_X1 U6088 ( .A1(n7715), .A2(n7713), .ZN(n4695) );
  NOR2_X1 U6089 ( .A1(n9009), .A2(n4926), .ZN(n9002) );
  NAND3_X1 U6090 ( .A1(n5150), .A2(n4701), .A3(n4956), .ZN(n4957) );
  AOI21_X1 U6091 ( .B1(P2_REG2_REG_5__SCAN_IN), .B2(n6586), .A(n6583), .ZN(
        n6585) );
  OAI21_X1 U6092 ( .B1(n5497), .B2(n4715), .A(n4713), .ZN(n5551) );
  NAND2_X1 U6093 ( .A1(n5629), .A2(n4728), .ZN(n4723) );
  NAND2_X1 U6094 ( .A1(n5629), .A2(n5628), .ZN(n5648) );
  NAND2_X1 U6095 ( .A1(n8837), .A2(n4733), .ZN(n4732) );
  NAND3_X1 U6096 ( .A1(n6195), .A2(n6218), .A3(n4746), .ZN(n4743) );
  NAND2_X1 U6097 ( .A1(n4743), .A2(n4744), .ZN(n6210) );
  NAND2_X1 U6098 ( .A1(n4751), .A2(n4749), .ZN(n8026) );
  NOR2_X1 U6099 ( .A1(n6224), .A2(n4757), .ZN(n4750) );
  NAND3_X1 U6100 ( .A1(n7803), .A2(n4753), .A3(n6299), .ZN(n4751) );
  NAND2_X1 U6101 ( .A1(n4760), .A2(n4761), .ZN(n8698) );
  NAND2_X1 U6102 ( .A1(n8745), .A2(n4764), .ZN(n4760) );
  INV_X1 U6103 ( .A(n6446), .ZN(n4767) );
  NAND2_X1 U6104 ( .A1(n4769), .A2(n4768), .ZN(n8746) );
  NOR2_X1 U6105 ( .A1(n6982), .A2(n6981), .ZN(n6980) );
  NAND2_X1 U6106 ( .A1(n4772), .A2(n6955), .ZN(n6982) );
  INV_X1 U6107 ( .A(n6952), .ZN(n4773) );
  NAND2_X1 U6108 ( .A1(n8621), .A2(n4775), .ZN(n4774) );
  OAI211_X1 U6109 ( .C1(n8621), .C2(n4779), .A(n4776), .B(n4774), .ZN(n8284)
         );
  NAND2_X1 U6110 ( .A1(n8621), .A2(n8622), .ZN(n4781) );
  INV_X1 U6111 ( .A(n7060), .ZN(n4787) );
  NAND2_X1 U6112 ( .A1(n4796), .A2(n4798), .ZN(n8065) );
  NAND2_X1 U6113 ( .A1(n7831), .A2(n4376), .ZN(n4796) );
  NAND2_X1 U6114 ( .A1(n4807), .A2(n4805), .ZN(n7026) );
  AOI21_X1 U6115 ( .B1(n4808), .B2(n7145), .A(n4806), .ZN(n4805) );
  INV_X1 U6116 ( .A(n7028), .ZN(n4806) );
  NAND2_X1 U6117 ( .A1(n7145), .A2(n7144), .ZN(n4810) );
  NAND2_X1 U6118 ( .A1(n7370), .A2(n4814), .ZN(n4811) );
  AOI21_X1 U6119 ( .B1(n4814), .B2(n4815), .A(n4813), .ZN(n4812) );
  OAI21_X1 U6120 ( .B1(n7370), .B2(n4815), .A(n4814), .ZN(n7704) );
  NAND2_X1 U6121 ( .A1(n7370), .A2(n7350), .ZN(n7441) );
  NOR2_X1 U6122 ( .A1(n7439), .A2(n7438), .ZN(n4821) );
  OAI21_X1 U6123 ( .B1(n8176), .B2(n4824), .A(n4822), .ZN(n8250) );
  NAND2_X1 U6124 ( .A1(n6190), .A2(n6189), .ZN(n6215) );
  NAND2_X1 U6125 ( .A1(n6190), .A2(n4833), .ZN(n6408) );
  NAND2_X1 U6126 ( .A1(n6904), .A2(n4427), .ZN(n8186) );
  NAND2_X1 U6127 ( .A1(n8186), .A2(n8431), .ZN(n7164) );
  OAI21_X1 U6128 ( .B1(n9360), .B2(n4840), .A(n4838), .ZN(n9325) );
  NAND2_X1 U6129 ( .A1(n9360), .A2(n4838), .ZN(n4837) );
  INV_X1 U6130 ( .A(n4844), .ZN(n9341) );
  INV_X1 U6131 ( .A(n9141), .ZN(n4843) );
  NAND2_X1 U6132 ( .A1(n9238), .A2(n4848), .ZN(n4845) );
  NAND2_X1 U6133 ( .A1(n4845), .A2(n4846), .ZN(n9174) );
  INV_X1 U6134 ( .A(n4854), .ZN(n4853) );
  NAND2_X1 U6135 ( .A1(n9214), .A2(n9211), .ZN(n4854) );
  NAND2_X1 U6136 ( .A1(n7783), .A2(n4864), .ZN(n4863) );
  NAND2_X1 U6137 ( .A1(n7910), .A2(n8333), .ZN(n7911) );
  NAND2_X1 U6138 ( .A1(n8333), .A2(n4870), .ZN(n4869) );
  INV_X1 U6139 ( .A(n8483), .ZN(n4870) );
  NAND3_X2 U6140 ( .A1(n4875), .A2(n5852), .A3(n5853), .ZN(n8656) );
  AND2_X1 U6141 ( .A1(n5851), .A2(n5850), .ZN(n4875) );
  OAI21_X1 U6142 ( .B1(n8709), .B2(n6447), .A(n4888), .ZN(n8693) );
  INV_X1 U6143 ( .A(n8876), .ZN(n4889) );
  AOI21_X2 U6144 ( .B1(n8816), .B2(n8827), .A(n6443), .ZN(n8807) );
  INV_X1 U6145 ( .A(n7471), .ZN(n4894) );
  NAND2_X1 U6146 ( .A1(n6436), .A2(n6437), .ZN(n4896) );
  NAND3_X1 U6147 ( .A1(n4896), .A2(n4387), .A3(n4892), .ZN(n7741) );
  NOR2_X1 U6148 ( .A1(n6436), .A2(n4897), .ZN(n7571) );
  NAND2_X1 U6149 ( .A1(n8898), .A2(n4902), .ZN(n4901) );
  INV_X1 U6150 ( .A(n4908), .ZN(n8757) );
  NAND2_X1 U6151 ( .A1(n4911), .A2(n4909), .ZN(n6428) );
  NOR2_X1 U6152 ( .A1(n4389), .A2(n4910), .ZN(n4909) );
  INV_X1 U6153 ( .A(n4915), .ZN(n7947) );
  INV_X1 U6154 ( .A(n8971), .ZN(n5801) );
  NAND2_X4 U6155 ( .A1(n8078), .A2(n8971), .ZN(n6152) );
  XNOR2_X2 U6156 ( .A(n5787), .B(P2_IR_REG_30__SCAN_IN), .ZN(n8971) );
  NAND2_X1 U6157 ( .A1(n6030), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5850) );
  NAND2_X2 U6158 ( .A1(n5801), .A2(n5792), .ZN(n5888) );
  CLKBUF_X1 U6159 ( .A(n6775), .Z(n8207) );
  CLKBUF_X1 U6160 ( .A(n9029), .Z(n9031) );
  OR2_X1 U6161 ( .A1(n5890), .A2(n5826), .ZN(n5829) );
  NAND2_X1 U6162 ( .A1(n5597), .A2(n5596), .ZN(n9043) );
  AOI22_X1 U6163 ( .A1(n6359), .A2(n6358), .B1(n6947), .B2(n6392), .ZN(n6396)
         );
  INV_X1 U6164 ( .A(n5202), .ZN(n5205) );
  NAND2_X1 U6165 ( .A1(n5004), .A2(n5003), .ZN(n5005) );
  AOI22_X1 U6166 ( .A1(n4398), .A2(n8214), .B1(n4990), .B2(n9949), .ZN(n4991)
         );
  NAND2_X1 U6167 ( .A1(n7279), .A2(n7178), .ZN(n8308) );
  CLKBUF_X1 U6168 ( .A(n7471), .Z(n7627) );
  OR2_X1 U6169 ( .A1(n5789), .A2(n5788), .ZN(n5791) );
  INV_X1 U6170 ( .A(n5792), .ZN(n8078) );
  OR2_X1 U6171 ( .A1(n6565), .A2(n9473), .ZN(n5858) );
  INV_X2 U6172 ( .A(n6565), .ZN(n6049) );
  INV_X1 U6173 ( .A(n6642), .ZN(n5063) );
  NAND2_X1 U6174 ( .A1(n8150), .A2(n6441), .ZN(n6442) );
  INV_X1 U6175 ( .A(n9301), .ZN(n9123) );
  AOI21_X1 U6176 ( .B1(n8746), .B2(n6327), .A(n8739), .ZN(n8745) );
  AND2_X1 U6177 ( .A1(n4961), .A2(n4941), .ZN(n4919) );
  OAI22_X1 U6178 ( .A1(n7203), .A2(n7202), .B1(n5859), .B2(n8656), .ZN(n7306)
         );
  INV_X1 U6179 ( .A(n8930), .ZN(n6439) );
  NAND2_X1 U6180 ( .A1(n5050), .A2(n5049), .ZN(n5074) );
  INV_X1 U6181 ( .A(n6467), .ZN(n6448) );
  NAND2_X1 U6182 ( .A1(n5023), .A2(n5022), .ZN(n5046) );
  AND2_X1 U6183 ( .A1(n6092), .A2(n6091), .ZN(n8775) );
  NAND2_X1 U6184 ( .A1(n5546), .A2(n5547), .ZN(n4925) );
  INV_X1 U6185 ( .A(n9075), .ZN(n5747) );
  AND2_X1 U6186 ( .A1(n5642), .A2(n5641), .ZN(n4926) );
  AND3_X1 U6187 ( .A1(n6033), .A2(n6032), .A3(n6031), .ZN(n8132) );
  OR2_X1 U6188 ( .A1(n8870), .A2(n8855), .ZN(n4927) );
  XOR2_X1 U6189 ( .A(n8903), .B(n8276), .Z(n4928) );
  NOR2_X1 U6190 ( .A1(n5103), .A2(n5102), .ZN(n4929) );
  NAND2_X1 U6191 ( .A1(n7286), .A2(n9708), .ZN(n9725) );
  OR2_X1 U6192 ( .A1(n5042), .A2(n6603), .ZN(n4930) );
  OR2_X1 U6193 ( .A1(n7227), .A2(n7232), .ZN(n5113) );
  INV_X1 U6194 ( .A(n7093), .ZN(n5897) );
  AND2_X1 U6195 ( .A1(n7475), .A2(n6266), .ZN(n5948) );
  AND3_X1 U6196 ( .A1(n5949), .A2(n5816), .A3(n5820), .ZN(n5775) );
  INV_X1 U6197 ( .A(n5090), .ZN(n5088) );
  NAND2_X1 U6198 ( .A1(n8251), .A2(n4928), .ZN(n8252) );
  INV_X1 U6199 ( .A(n6041), .ZN(n6039) );
  INV_X1 U6200 ( .A(n6020), .ZN(n6019) );
  NAND2_X1 U6201 ( .A1(n8633), .A2(n8682), .ZN(n6472) );
  INV_X1 U6202 ( .A(n8775), .ZN(n6444) );
  INV_X1 U6203 ( .A(n5918), .ZN(n5795) );
  INV_X1 U6204 ( .A(n7763), .ZN(n8940) );
  OR2_X1 U6205 ( .A1(n7089), .A2(n7101), .ZN(n7216) );
  CLKBUF_X3 U6206 ( .A(n5026), .Z(n6492) );
  INV_X1 U6207 ( .A(n5657), .ZN(n5655) );
  INV_X1 U6208 ( .A(n5157), .ZN(n5155) );
  INV_X1 U6209 ( .A(n5218), .ZN(n5216) );
  INV_X1 U6210 ( .A(n8474), .ZN(n6892) );
  OR2_X1 U6211 ( .A1(n5346), .A2(n5345), .ZN(n5347) );
  INV_X1 U6212 ( .A(n5285), .ZN(n5326) );
  AND2_X1 U6213 ( .A1(n8113), .A2(n8063), .ZN(n8064) );
  NAND2_X1 U6214 ( .A1(n6063), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6074) );
  OR2_X1 U6215 ( .A1(n5968), .A2(n5967), .ZN(n5980) );
  NAND2_X1 U6216 ( .A1(n6004), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6020) );
  OR2_X1 U6217 ( .A1(n6127), .A2(n6126), .ZN(n6150) );
  OR2_X1 U6218 ( .A1(n6074), .A2(n10062), .ZN(n6085) );
  OR2_X1 U6219 ( .A1(n5993), .A2(n10059), .ZN(n6006) );
  NAND2_X1 U6220 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5891) );
  NAND2_X1 U6221 ( .A1(n8231), .A2(n8680), .ZN(n8232) );
  OR2_X1 U6222 ( .A1(n5941), .A2(n5796), .ZN(n5957) );
  AND2_X1 U6223 ( .A1(n6260), .A2(n6261), .ZN(n6429) );
  INV_X1 U6224 ( .A(n7510), .ZN(n5870) );
  INV_X1 U6225 ( .A(n7094), .ZN(n7086) );
  INV_X1 U6226 ( .A(n7243), .ZN(n5173) );
  NAND2_X1 U6227 ( .A1(n5205), .A2(n5204), .ZN(n7591) );
  INV_X1 U6228 ( .A(n5272), .ZN(n5270) );
  NAND2_X1 U6229 ( .A1(n5655), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n5684) );
  NAND2_X1 U6230 ( .A1(n5533), .A2(n5532), .ZN(n5557) );
  OR2_X1 U6231 ( .A1(n5333), .A2(n6842), .ZN(n5335) );
  NAND2_X1 U6232 ( .A1(n6642), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n4999) );
  AOI21_X1 U6233 ( .B1(n9174), .B2(n9173), .A(n9152), .ZN(n9155) );
  NAND2_X1 U6234 ( .A1(n5396), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5427) );
  INV_X1 U6235 ( .A(n9376), .ZN(n9161) );
  OR2_X1 U6236 ( .A1(n9703), .A2(n8209), .ZN(n7388) );
  INV_X1 U6237 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5740) );
  NAND2_X1 U6238 ( .A1(n6161), .A2(n6160), .ZN(n6166) );
  NAND2_X1 U6239 ( .A1(n5444), .A2(n5443), .ZN(n5446) );
  NAND2_X1 U6240 ( .A1(n5287), .A2(n5286), .ZN(n5290) );
  NAND2_X1 U6241 ( .A1(n5207), .A2(n5184), .ZN(n5185) );
  INV_X1 U6242 ( .A(n8634), .ZN(n8715) );
  OR2_X1 U6243 ( .A1(n6053), .A2(n8178), .ZN(n6064) );
  OR2_X1 U6244 ( .A1(n8068), .A2(n8067), .ZN(n8069) );
  OR2_X1 U6245 ( .A1(n8627), .A2(n8830), .ZN(n8603) );
  AND2_X1 U6246 ( .A1(n6150), .A2(n6128), .ZN(n8732) );
  AND2_X1 U6247 ( .A1(n6102), .A2(n6101), .ZN(n8613) );
  OR2_X1 U6248 ( .A1(n5888), .A2(n5871), .ZN(n5879) );
  INV_X1 U6249 ( .A(n8739), .ZN(n8744) );
  INV_X1 U6250 ( .A(n7944), .ZN(n7949) );
  INV_X1 U6251 ( .A(n7841), .ZN(n7847) );
  INV_X1 U6252 ( .A(n6437), .ZN(n7572) );
  XNOR2_X1 U6253 ( .A(n5201), .B(n7160), .ZN(n7592) );
  AND2_X1 U6254 ( .A1(n5112), .A2(n5111), .ZN(n7232) );
  OR2_X1 U6255 ( .A1(n5670), .A2(n5669), .ZN(n5671) );
  AND2_X1 U6256 ( .A1(n8543), .A2(n4989), .ZN(n7043) );
  OR2_X1 U6257 ( .A1(n5684), .A2(n5683), .ZN(n5753) );
  OR2_X1 U6258 ( .A1(n5485), .A2(n5484), .ZN(n5531) );
  INV_X1 U6259 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6750) );
  INV_X1 U6260 ( .A(n9217), .ZN(n9176) );
  NAND2_X1 U6261 ( .A1(n9151), .A2(n8443), .ZN(n9196) );
  AND2_X1 U6262 ( .A1(n9402), .A2(n9259), .ZN(n9129) );
  INV_X1 U6263 ( .A(n9117), .ZN(n9565) );
  AND2_X1 U6264 ( .A1(n6900), .A2(n6899), .ZN(n9499) );
  INV_X1 U6265 ( .A(n4947), .ZN(n8555) );
  AND2_X1 U6266 ( .A1(n5445), .A2(n5419), .ZN(n5443) );
  INV_X1 U6267 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9456) );
  AND2_X1 U6268 ( .A1(n7018), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8625) );
  INV_X1 U6269 ( .A(n7514), .ZN(n6399) );
  AND2_X1 U6270 ( .A1(n6123), .A2(n6122), .ZN(n8263) );
  OR2_X1 U6271 ( .A1(n5888), .A2(n5903), .ZN(n5910) );
  NAND2_X1 U6272 ( .A1(n6316), .A2(n6318), .ZN(n8827) );
  OR2_X1 U6273 ( .A1(n9838), .A2(n7080), .ZN(n9825) );
  INV_X1 U6274 ( .A(n8685), .ZN(n8858) );
  OR2_X1 U6275 ( .A1(n9840), .A2(n6451), .ZN(n7104) );
  INV_X1 U6276 ( .A(n9014), .ZN(n9067) );
  OR2_X1 U6277 ( .A1(n5753), .A2(n5750), .ZN(n9163) );
  INV_X1 U6278 ( .A(n5758), .ZN(n6500) );
  NAND2_X1 U6279 ( .A1(n8335), .A2(n8412), .ZN(n7905) );
  INV_X1 U6280 ( .A(n9346), .ZN(n9713) );
  OR2_X1 U6281 ( .A1(n6886), .A2(n5749), .ZN(n9708) );
  AND2_X1 U6282 ( .A1(n9725), .A2(n7041), .ZN(n9543) );
  OR2_X1 U6283 ( .A1(n9793), .A2(n9502), .ZN(n9783) );
  INV_X1 U6284 ( .A(n8514), .ZN(n5744) );
  XNOR2_X1 U6285 ( .A(n5126), .B(SI_5_), .ZN(n5124) );
  OR2_X1 U6286 ( .A1(n6416), .A2(n6415), .ZN(n6417) );
  OR3_X1 U6287 ( .A1(n6024), .A2(n6023), .A3(n6022), .ZN(n8640) );
  INV_X1 U6288 ( .A(n6482), .ZN(n6483) );
  NAND2_X1 U6289 ( .A1(n6477), .A2(n9825), .ZN(n9834) );
  INV_X1 U6290 ( .A(n9909), .ZN(n9907) );
  INV_X1 U6291 ( .A(n9839), .ZN(n9843) );
  INV_X1 U6292 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n10216) );
  INV_X1 U6293 ( .A(n6556), .ZN(n9487) );
  NAND2_X1 U6294 ( .A1(n5692), .A2(n5691), .ZN(n9232) );
  INV_X1 U6295 ( .A(n9543), .ZN(n9357) );
  INV_X1 U6296 ( .A(n9795), .ZN(n9794) );
  INV_X1 U6297 ( .A(n4948), .ZN(n8109) );
  INV_X1 U6298 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n10150) );
  INV_X1 U6299 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n10181) );
  NAND2_X1 U6300 ( .A1(n4927), .A2(n6483), .ZN(P2_U3267) );
  NOR2_X1 U6301 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n4934) );
  NOR2_X1 U6302 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n4933) );
  NOR2_X1 U6303 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n4932) );
  NOR2_X1 U6304 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n4938) );
  NOR2_X1 U6305 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n4937) );
  NOR2_X1 U6306 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n4936) );
  NAND4_X1 U6307 ( .A1(n4938), .A2(n4937), .A3(n4936), .A4(n4958), .ZN(n4939)
         );
  INV_X1 U6308 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n4961) );
  INV_X1 U6309 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n4941) );
  NAND2_X1 U6310 ( .A1(n4945), .A2(n4942), .ZN(n9457) );
  XNOR2_X2 U6311 ( .A(n4944), .B(n4943), .ZN(n4947) );
  NAND2_X1 U6312 ( .A1(n6642), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n4952) );
  AND2_X2 U6313 ( .A1(n8555), .A2(n8109), .ZN(n5154) );
  NAND2_X1 U6314 ( .A1(n5154), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n4951) );
  NAND2_X1 U6315 ( .A1(n5114), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n4950) );
  AND2_X2 U6316 ( .A1(n8555), .A2(n4948), .ZN(n5037) );
  NAND2_X1 U6317 ( .A1(n5037), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n4949) );
  NAND4_X1 U6318 ( .A1(n4952), .A2(n4951), .A3(n4950), .A4(n4949), .ZN(n6638)
         );
  INV_X1 U6319 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n4953) );
  INV_X1 U6320 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n4954) );
  NAND2_X1 U6321 ( .A1(n4960), .A2(n4958), .ZN(n4959) );
  INV_X1 U6322 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n4981) );
  INV_X1 U6323 ( .A(n4987), .ZN(n6906) );
  NAND2_X1 U6324 ( .A1(n4409), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4963) );
  NAND2_X1 U6325 ( .A1(n4963), .A2(n4961), .ZN(n4965) );
  NAND2_X1 U6326 ( .A1(n4965), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4962) );
  XNOR2_X1 U6327 ( .A(n4962), .B(P1_IR_REG_26__SCAN_IN), .ZN(n5725) );
  INV_X1 U6328 ( .A(n4963), .ZN(n4964) );
  NAND2_X1 U6329 ( .A1(n4964), .A2(P1_IR_REG_25__SCAN_IN), .ZN(n4966) );
  NAND2_X1 U6330 ( .A1(n4966), .A2(n4965), .ZN(n7814) );
  NAND2_X1 U6331 ( .A1(n4967), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4968) );
  XNOR2_X1 U6332 ( .A(n4968), .B(n4874), .ZN(n7644) );
  NOR2_X1 U6333 ( .A1(n7814), .A2(n7644), .ZN(n4969) );
  NAND2_X2 U6334 ( .A1(n5725), .A2(n4969), .ZN(n6513) );
  NAND2_X1 U6335 ( .A1(n6638), .A2(n4398), .ZN(n4980) );
  INV_X1 U6336 ( .A(SI_0_), .ZN(n4971) );
  INV_X1 U6337 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n4970) );
  OAI21_X1 U6338 ( .B1(n6607), .B2(n4971), .A(n4970), .ZN(n4974) );
  AND2_X1 U6339 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n4972) );
  NAND2_X1 U6340 ( .A1(n4973), .A2(n4972), .ZN(n4995) );
  AND2_X1 U6341 ( .A1(n4974), .A2(n4995), .ZN(n6600) );
  INV_X1 U6342 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n4975) );
  MUX2_X1 U6343 ( .A(n9949), .B(n6600), .S(n5042), .Z(n8214) );
  AND2_X2 U6344 ( .A1(n4987), .A2(n6513), .ZN(n5026) );
  INV_X1 U6345 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n10055) );
  NOR2_X1 U6346 ( .A1(n6513), .A2(n10055), .ZN(n4978) );
  AOI21_X1 U6347 ( .B1(n8214), .B2(n5026), .A(n4978), .ZN(n4979) );
  NAND2_X1 U6348 ( .A1(n4980), .A2(n4979), .ZN(n6521) );
  INV_X1 U6349 ( .A(n6521), .ZN(n4988) );
  NAND2_X1 U6350 ( .A1(n4982), .A2(n4981), .ZN(n4983) );
  INV_X1 U6351 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n4984) );
  INV_X1 U6352 ( .A(n5743), .ZN(n5738) );
  XNOR2_X2 U6353 ( .A(n4986), .B(P1_IR_REG_19__SCAN_IN), .ZN(n5505) );
  NAND2_X1 U6354 ( .A1(n6907), .A2(n4987), .ZN(n5055) );
  NAND2_X1 U6355 ( .A1(n4988), .A2(n5055), .ZN(n4993) );
  NAND2_X1 U6356 ( .A1(n5743), .A2(n7043), .ZN(n6908) );
  AND2_X4 U6357 ( .A1(n5026), .A2(n6908), .ZN(n5640) );
  NAND2_X1 U6358 ( .A1(n6638), .A2(n5640), .ZN(n4992) );
  INV_X1 U6359 ( .A(n6513), .ZN(n4990) );
  AND2_X1 U6360 ( .A1(n4992), .A2(n4991), .ZN(n6523) );
  NAND2_X1 U6361 ( .A1(n4993), .A2(n6522), .ZN(n5009) );
  INV_X1 U6362 ( .A(n5009), .ZN(n5007) );
  INV_X1 U6363 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6604) );
  NAND3_X1 U6364 ( .A1(n5239), .A2(SI_0_), .A3(P1_DATAO_REG_0__SCAN_IN), .ZN(
        n4994) );
  INV_X1 U6365 ( .A(SI_1_), .ZN(n4996) );
  XNOR2_X1 U6366 ( .A(n5021), .B(n4996), .ZN(n5020) );
  MUX2_X1 U6367 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n4973), .Z(n5019) );
  XNOR2_X1 U6368 ( .A(n5020), .B(n5019), .ZN(n6615) );
  INV_X1 U6369 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n4998) );
  NAND2_X1 U6370 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n9949), .ZN(n4997) );
  XNOR2_X1 U6371 ( .A(n4998), .B(n4997), .ZN(n6603) );
  NAND2_X1 U6372 ( .A1(n6901), .A2(n5026), .ZN(n5004) );
  NAND2_X1 U6373 ( .A1(n5154), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5001) );
  NAND2_X1 U6374 ( .A1(n5037), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5000) );
  NAND4_X2 U6375 ( .A1(n5002), .A2(n5001), .A3(n5000), .A4(n4999), .ZN(n5011)
         );
  NAND2_X1 U6376 ( .A1(n5011), .A2(n4398), .ZN(n5003) );
  XNOR2_X1 U6377 ( .A(n5005), .B(n6490), .ZN(n5008) );
  INV_X1 U6378 ( .A(n5008), .ZN(n5006) );
  NAND2_X1 U6379 ( .A1(n5007), .A2(n5006), .ZN(n5010) );
  NAND2_X1 U6380 ( .A1(n5009), .A2(n5008), .ZN(n8203) );
  NAND2_X1 U6381 ( .A1(n5010), .A2(n8203), .ZN(n6774) );
  INV_X1 U6382 ( .A(n6774), .ZN(n5015) );
  NAND2_X1 U6383 ( .A1(n5011), .A2(n5640), .ZN(n5013) );
  NAND2_X1 U6384 ( .A1(n5096), .A2(n6901), .ZN(n5012) );
  NAND2_X1 U6385 ( .A1(n5013), .A2(n5012), .ZN(n6777) );
  NAND2_X1 U6386 ( .A1(n5015), .A2(n5014), .ZN(n6775) );
  NAND2_X1 U6387 ( .A1(n6775), .A2(n8203), .ZN(n5036) );
  NAND2_X1 U6388 ( .A1(n5114), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6891) );
  NAND2_X1 U6389 ( .A1(n6642), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n6890) );
  NAND2_X1 U6390 ( .A1(n5154), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6889) );
  NAND2_X1 U6391 ( .A1(n5037), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n6888) );
  NAND2_X1 U6392 ( .A1(n9712), .A2(n5096), .ZN(n5028) );
  INV_X1 U6393 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5017) );
  OAI21_X1 U6394 ( .B1(n5018), .B2(n5017), .A(n5043), .ZN(n6605) );
  OR2_X1 U6395 ( .A1(n8391), .A2(n6606), .ZN(n5025) );
  NAND2_X1 U6396 ( .A1(n5020), .A2(n5019), .ZN(n5023) );
  NAND2_X1 U6397 ( .A1(n5021), .A2(SI_1_), .ZN(n5022) );
  MUX2_X1 U6398 ( .A(n6609), .B(n6606), .S(n4973), .Z(n5047) );
  XNOR2_X1 U6399 ( .A(n5046), .B(n5045), .ZN(n6608) );
  OR2_X1 U6400 ( .A1(n5129), .A2(n6608), .ZN(n5024) );
  OAI211_X1 U6401 ( .C1(n5042), .C2(n6605), .A(n5025), .B(n5024), .ZN(n8209)
         );
  NAND2_X1 U6402 ( .A1(n8209), .A2(n6492), .ZN(n5027) );
  NAND2_X1 U6403 ( .A1(n5028), .A2(n5027), .ZN(n5029) );
  XNOR2_X1 U6404 ( .A(n5029), .B(n6490), .ZN(n5031) );
  AND2_X1 U6405 ( .A1(n5096), .A2(n8209), .ZN(n5030) );
  AOI21_X1 U6406 ( .B1(n9712), .B2(n5640), .A(n5030), .ZN(n5032) );
  NAND2_X1 U6407 ( .A1(n5031), .A2(n5032), .ZN(n6877) );
  INV_X1 U6408 ( .A(n5031), .ZN(n5034) );
  INV_X1 U6409 ( .A(n5032), .ZN(n5033) );
  NAND2_X1 U6410 ( .A1(n5034), .A2(n5033), .ZN(n5035) );
  AND2_X1 U6411 ( .A1(n6877), .A2(n5035), .ZN(n8205) );
  NAND2_X1 U6412 ( .A1(n5036), .A2(n8205), .ZN(n6874) );
  NAND2_X1 U6413 ( .A1(n6874), .A2(n6877), .ZN(n5061) );
  INV_X1 U6414 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n6681) );
  NAND2_X1 U6415 ( .A1(n5037), .A2(n6681), .ZN(n5041) );
  NAND2_X1 U6416 ( .A1(n5114), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5040) );
  NAND2_X1 U6417 ( .A1(n5154), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5039) );
  NAND2_X1 U6418 ( .A1(n6642), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5038) );
  NAND2_X1 U6419 ( .A1(n9088), .A2(n5096), .ZN(n5054) );
  INV_X1 U6420 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5044) );
  INV_X1 U6421 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n9978) );
  OR2_X1 U6422 ( .A1(n8391), .A2(n9978), .ZN(n5052) );
  NAND2_X1 U6423 ( .A1(n5046), .A2(n5045), .ZN(n5050) );
  INV_X1 U6424 ( .A(n5047), .ZN(n5048) );
  NAND2_X1 U6425 ( .A1(n5048), .A2(SI_2_), .ZN(n5049) );
  INV_X1 U6426 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6610) );
  MUX2_X1 U6427 ( .A(n6610), .B(n9978), .S(n4973), .Z(n5075) );
  XNOR2_X1 U6428 ( .A(n5074), .B(n5073), .ZN(n6622) );
  OR2_X1 U6429 ( .A1(n5129), .A2(n6622), .ZN(n5051) );
  OAI211_X1 U6430 ( .C1(n5042), .C2(n6710), .A(n5052), .B(n5051), .ZN(n7049)
         );
  NAND2_X1 U6431 ( .A1(n7049), .A2(n6492), .ZN(n5053) );
  NAND2_X1 U6432 ( .A1(n5054), .A2(n5053), .ZN(n5056) );
  XNOR2_X1 U6433 ( .A(n5056), .B(n6490), .ZN(n5059) );
  AND2_X1 U6434 ( .A1(n5096), .A2(n7049), .ZN(n5057) );
  AOI21_X1 U6435 ( .B1(n9088), .B2(n5640), .A(n5057), .ZN(n5058) );
  NAND2_X1 U6436 ( .A1(n5059), .A2(n5058), .ZN(n5062) );
  NAND2_X1 U6437 ( .A1(n5061), .A2(n6875), .ZN(n6879) );
  NAND2_X1 U6438 ( .A1(n6879), .A2(n5062), .ZN(n9019) );
  NAND2_X1 U6439 ( .A1(n8287), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5068) );
  INV_X4 U6440 ( .A(n5063), .ZN(n8289) );
  NAND2_X1 U6441 ( .A1(n8289), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5067) );
  INV_X1 U6442 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n10215) );
  NAND2_X1 U6443 ( .A1(n6681), .A2(n10215), .ZN(n5064) );
  AND2_X1 U6444 ( .A1(n5064), .A2(n5090), .ZN(n9023) );
  NAND2_X1 U6445 ( .A1(n5037), .A2(n9023), .ZN(n5066) );
  NAND2_X1 U6446 ( .A1(n5154), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5065) );
  NAND4_X1 U6447 ( .A1(n5068), .A2(n5067), .A3(n5066), .A4(n5065), .ZN(n9087)
         );
  NAND2_X1 U6448 ( .A1(n9087), .A2(n5096), .ZN(n5081) );
  NAND2_X1 U6449 ( .A1(n5069), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5070) );
  MUX2_X1 U6450 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5070), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n5072) );
  NAND2_X1 U6451 ( .A1(n5072), .A2(n5071), .ZN(n9612) );
  INV_X1 U6452 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6611) );
  OR2_X1 U6453 ( .A1(n8391), .A2(n6611), .ZN(n5079) );
  INV_X1 U6454 ( .A(n5075), .ZN(n5076) );
  NAND2_X1 U6455 ( .A1(n5076), .A2(SI_3_), .ZN(n5100) );
  NAND2_X1 U6456 ( .A1(n5105), .A2(n5100), .ZN(n5077) );
  INV_X1 U6457 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6614) );
  MUX2_X1 U6458 ( .A(n6614), .B(n6611), .S(n4973), .Z(n5098) );
  XNOR2_X1 U6459 ( .A(n5077), .B(n5102), .ZN(n6613) );
  OR2_X1 U6460 ( .A1(n5129), .A2(n6613), .ZN(n5078) );
  OAI211_X1 U6461 ( .C1(n5042), .C2(n9612), .A(n5079), .B(n5078), .ZN(n9022)
         );
  NAND2_X1 U6462 ( .A1(n9022), .A2(n6492), .ZN(n5080) );
  NAND2_X1 U6463 ( .A1(n5081), .A2(n5080), .ZN(n5082) );
  INV_X1 U6464 ( .A(n6490), .ZN(n7160) );
  XNOR2_X1 U6465 ( .A(n5082), .B(n7160), .ZN(n5084) );
  AND2_X1 U6466 ( .A1(n5096), .A2(n9022), .ZN(n5083) );
  AOI21_X1 U6467 ( .B1(n9087), .B2(n5640), .A(n5083), .ZN(n5085) );
  XNOR2_X1 U6468 ( .A(n5084), .B(n5085), .ZN(n9020) );
  INV_X1 U6469 ( .A(n5084), .ZN(n5086) );
  NAND2_X1 U6470 ( .A1(n5086), .A2(n5085), .ZN(n5087) );
  NAND2_X1 U6471 ( .A1(n8287), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5095) );
  INV_X1 U6472 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5089) );
  NAND2_X1 U6473 ( .A1(n5090), .A2(n5089), .ZN(n5091) );
  AND2_X1 U6474 ( .A1(n5116), .A2(n5091), .ZN(n7233) );
  NAND2_X1 U6475 ( .A1(n5037), .A2(n7233), .ZN(n5094) );
  NAND2_X1 U6476 ( .A1(n5154), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5093) );
  NAND2_X1 U6477 ( .A1(n8289), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5092) );
  NAND2_X1 U6478 ( .A1(n9086), .A2(n5096), .ZN(n5109) );
  NAND2_X1 U6479 ( .A1(n5071), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5097) );
  XNOR2_X1 U6480 ( .A(n5097), .B(P1_IR_REG_5__SCAN_IN), .ZN(n9639) );
  INV_X1 U6481 ( .A(n9639), .ZN(n6617) );
  INV_X1 U6482 ( .A(n5098), .ZN(n5099) );
  NAND2_X1 U6483 ( .A1(n5099), .A2(SI_4_), .ZN(n5101) );
  AND2_X1 U6484 ( .A1(n5100), .A2(n5101), .ZN(n5104) );
  INV_X1 U6485 ( .A(n5101), .ZN(n5103) );
  INV_X1 U6486 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6621) );
  MUX2_X1 U6487 ( .A(n6621), .B(n6618), .S(n5601), .Z(n5126) );
  XNOR2_X1 U6488 ( .A(n5125), .B(n5124), .ZN(n6620) );
  OR2_X1 U6489 ( .A1(n5129), .A2(n6620), .ZN(n5107) );
  OR2_X1 U6490 ( .A1(n8391), .A2(n6618), .ZN(n5106) );
  NAND2_X1 U6491 ( .A1(n7251), .A2(n6492), .ZN(n5108) );
  NAND2_X1 U6492 ( .A1(n5109), .A2(n5108), .ZN(n5110) );
  XNOR2_X1 U6493 ( .A(n5110), .B(n6490), .ZN(n7227) );
  NAND2_X1 U6494 ( .A1(n9086), .A2(n5640), .ZN(n5112) );
  NAND2_X1 U6495 ( .A1(n5096), .A2(n7251), .ZN(n5111) );
  NAND2_X1 U6496 ( .A1(n8289), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5121) );
  NAND2_X1 U6497 ( .A1(n5114), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5120) );
  INV_X1 U6498 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n7327) );
  NAND2_X1 U6499 ( .A1(n5116), .A2(n7327), .ZN(n5117) );
  AND2_X1 U6500 ( .A1(n5157), .A2(n5117), .ZN(n7329) );
  NAND2_X1 U6501 ( .A1(n5037), .A2(n7329), .ZN(n5119) );
  NAND2_X1 U6502 ( .A1(n5154), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5118) );
  NAND2_X1 U6503 ( .A1(n9085), .A2(n5096), .ZN(n5133) );
  OR2_X1 U6504 ( .A1(n5122), .A2(n9456), .ZN(n5123) );
  XNOR2_X1 U6505 ( .A(n5123), .B(P1_IR_REG_6__SCAN_IN), .ZN(n9652) );
  INV_X1 U6506 ( .A(n5126), .ZN(n5127) );
  NAND2_X1 U6507 ( .A1(n5127), .A2(SI_5_), .ZN(n5143) );
  NAND2_X1 U6508 ( .A1(n5149), .A2(n5143), .ZN(n5128) );
  MUX2_X1 U6509 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n4973), .Z(n5142) );
  XNOR2_X1 U6510 ( .A(n5128), .B(n5145), .ZN(n6625) );
  NAND2_X1 U6511 ( .A1(n6625), .A2(n8389), .ZN(n5130) );
  NAND2_X1 U6512 ( .A1(n7328), .A2(n6492), .ZN(n5132) );
  NAND2_X1 U6513 ( .A1(n5133), .A2(n5132), .ZN(n5134) );
  XNOR2_X1 U6514 ( .A(n5134), .B(n6490), .ZN(n7324) );
  NAND2_X1 U6515 ( .A1(n9085), .A2(n5640), .ZN(n5136) );
  NAND2_X1 U6516 ( .A1(n7328), .A2(n5096), .ZN(n5135) );
  AND2_X1 U6517 ( .A1(n5136), .A2(n5135), .ZN(n5138) );
  AOI22_X1 U6518 ( .A1(n7232), .A2(n7227), .B1(n7324), .B2(n5138), .ZN(n5137)
         );
  INV_X1 U6519 ( .A(n7324), .ZN(n5139) );
  INV_X1 U6520 ( .A(n5138), .ZN(n7323) );
  NAND2_X1 U6521 ( .A1(n5139), .A2(n7323), .ZN(n5140) );
  NAND2_X1 U6522 ( .A1(n5141), .A2(n5140), .ZN(n7240) );
  INV_X1 U6523 ( .A(n7240), .ZN(n5174) );
  NAND2_X1 U6524 ( .A1(n5142), .A2(SI_6_), .ZN(n5144) );
  AND2_X1 U6525 ( .A1(n5143), .A2(n5144), .ZN(n5148) );
  INV_X1 U6526 ( .A(n5144), .ZN(n5147) );
  MUX2_X1 U6527 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n4973), .Z(n5178) );
  XNOR2_X1 U6528 ( .A(n5177), .B(n5176), .ZN(n6629) );
  NAND2_X1 U6529 ( .A1(n6629), .A2(n8389), .ZN(n5153) );
  OR2_X1 U6530 ( .A1(n5150), .A2(n9456), .ZN(n5151) );
  XNOR2_X1 U6531 ( .A(n5151), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6719) );
  AOI22_X1 U6532 ( .A1(n5506), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n9601), .B2(
        n6719), .ZN(n5152) );
  NAND2_X1 U6533 ( .A1(n5153), .A2(n5152), .ZN(n7581) );
  NAND2_X1 U6534 ( .A1(n7581), .A2(n6492), .ZN(n5164) );
  NAND2_X1 U6535 ( .A1(n8287), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5162) );
  NAND2_X1 U6536 ( .A1(n5154), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5161) );
  INV_X1 U6537 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5156) );
  NAND2_X1 U6538 ( .A1(n5157), .A2(n5156), .ZN(n5158) );
  AND2_X1 U6539 ( .A1(n5193), .A2(n5158), .ZN(n7287) );
  NAND2_X1 U6540 ( .A1(n5037), .A2(n7287), .ZN(n5160) );
  NAND2_X1 U6541 ( .A1(n8289), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5159) );
  NAND4_X1 U6542 ( .A1(n5162), .A2(n5161), .A3(n5160), .A4(n5159), .ZN(n9084)
         );
  NAND2_X1 U6543 ( .A1(n9084), .A2(n5096), .ZN(n5163) );
  NAND2_X1 U6544 ( .A1(n5164), .A2(n5163), .ZN(n5165) );
  XNOR2_X1 U6545 ( .A(n5165), .B(n6490), .ZN(n5168) );
  NAND2_X1 U6546 ( .A1(n7581), .A2(n5096), .ZN(n5167) );
  NAND2_X1 U6547 ( .A1(n9084), .A2(n5640), .ZN(n5166) );
  AND2_X1 U6548 ( .A1(n5167), .A2(n5166), .ZN(n5169) );
  NAND2_X1 U6549 ( .A1(n5168), .A2(n5169), .ZN(n5175) );
  INV_X1 U6550 ( .A(n5168), .ZN(n5171) );
  INV_X1 U6551 ( .A(n5169), .ZN(n5170) );
  NAND2_X1 U6552 ( .A1(n5171), .A2(n5170), .ZN(n5172) );
  NAND2_X1 U6553 ( .A1(n5175), .A2(n5172), .ZN(n7243) );
  NAND2_X1 U6554 ( .A1(n5174), .A2(n5173), .ZN(n7241) );
  NAND2_X1 U6555 ( .A1(n7241), .A2(n5175), .ZN(n5202) );
  NAND2_X1 U6556 ( .A1(n5178), .A2(SI_7_), .ZN(n5179) );
  MUX2_X1 U6557 ( .A(n10073), .B(n10181), .S(n4973), .Z(n5182) );
  INV_X1 U6558 ( .A(SI_8_), .ZN(n5181) );
  INV_X1 U6559 ( .A(n5182), .ZN(n5183) );
  NAND2_X1 U6560 ( .A1(n5183), .A2(SI_8_), .ZN(n5184) );
  NAND2_X1 U6561 ( .A1(n5186), .A2(n5185), .ZN(n5187) );
  NAND2_X1 U6562 ( .A1(n5208), .A2(n5187), .ZN(n6633) );
  NAND2_X1 U6563 ( .A1(n6633), .A2(n8389), .ZN(n5192) );
  NAND2_X1 U6564 ( .A1(n5188), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5189) );
  MUX2_X1 U6565 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5189), .S(
        P1_IR_REG_8__SCAN_IN), .Z(n5190) );
  AND2_X1 U6566 ( .A1(n5190), .A2(n5246), .ZN(n6708) );
  AOI22_X1 U6567 ( .A1(n5506), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n9601), .B2(
        n6708), .ZN(n5191) );
  NAND2_X1 U6568 ( .A1(n5192), .A2(n5191), .ZN(n7595) );
  NAND2_X1 U6569 ( .A1(n8289), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5198) );
  NAND2_X1 U6570 ( .A1(n8287), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5197) );
  NAND2_X1 U6571 ( .A1(n5193), .A2(n6750), .ZN(n5194) );
  AND2_X1 U6572 ( .A1(n5218), .A2(n5194), .ZN(n7596) );
  NAND2_X1 U6573 ( .A1(n5037), .A2(n7596), .ZN(n5196) );
  INV_X1 U6574 ( .A(n5154), .ZN(n5709) );
  NAND2_X1 U6575 ( .A1(n8288), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5195) );
  AOI22_X1 U6576 ( .A1(n7595), .A2(n5096), .B1(n5640), .B2(n9083), .ZN(n5203)
         );
  NAND2_X1 U6577 ( .A1(n5202), .A2(n5203), .ZN(n7590) );
  NAND2_X1 U6578 ( .A1(n7595), .A2(n6492), .ZN(n5200) );
  NAND2_X1 U6579 ( .A1(n9083), .A2(n4398), .ZN(n5199) );
  NAND2_X1 U6580 ( .A1(n5200), .A2(n5199), .ZN(n5201) );
  NAND2_X1 U6581 ( .A1(n7590), .A2(n7592), .ZN(n5206) );
  INV_X1 U6582 ( .A(n5203), .ZN(n5204) );
  NAND2_X1 U6583 ( .A1(n5206), .A2(n7591), .ZN(n7657) );
  INV_X1 U6584 ( .A(n7657), .ZN(n5234) );
  INV_X1 U6585 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n5209) );
  MUX2_X1 U6586 ( .A(n10082), .B(n5209), .S(n4973), .Z(n5210) );
  INV_X1 U6587 ( .A(SI_9_), .ZN(n10029) );
  INV_X1 U6588 ( .A(n5210), .ZN(n5211) );
  NAND2_X1 U6589 ( .A1(n5211), .A2(SI_9_), .ZN(n5212) );
  XNOR2_X1 U6590 ( .A(n5236), .B(n4923), .ZN(n6636) );
  NAND2_X1 U6591 ( .A1(n6636), .A2(n8389), .ZN(n5215) );
  NAND2_X1 U6592 ( .A1(n5246), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5213) );
  XNOR2_X1 U6593 ( .A(n5213), .B(P1_IR_REG_9__SCAN_IN), .ZN(n9667) );
  AOI22_X1 U6594 ( .A1(n5506), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n9601), .B2(
        n9667), .ZN(n5214) );
  NAND2_X1 U6595 ( .A1(n9786), .A2(n6492), .ZN(n5225) );
  INV_X1 U6596 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5217) );
  NAND2_X1 U6597 ( .A1(n5218), .A2(n5217), .ZN(n5219) );
  AND2_X1 U6598 ( .A1(n5249), .A2(n5219), .ZN(n7660) );
  NAND2_X1 U6599 ( .A1(n5758), .A2(n7660), .ZN(n5223) );
  NAND2_X1 U6600 ( .A1(n8287), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5222) );
  NAND2_X1 U6601 ( .A1(n8288), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5221) );
  NAND2_X1 U6602 ( .A1(n8289), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5220) );
  NAND4_X1 U6603 ( .A1(n5223), .A2(n5222), .A3(n5221), .A4(n5220), .ZN(n9497)
         );
  NAND2_X1 U6604 ( .A1(n9497), .A2(n4398), .ZN(n5224) );
  NAND2_X1 U6605 ( .A1(n5225), .A2(n5224), .ZN(n5226) );
  XNOR2_X1 U6606 ( .A(n5226), .B(n6490), .ZN(n5228) );
  AND2_X1 U6607 ( .A1(n9497), .A2(n5640), .ZN(n5227) );
  AOI21_X1 U6608 ( .B1(n9786), .B2(n4398), .A(n5227), .ZN(n5229) );
  NAND2_X1 U6609 ( .A1(n5228), .A2(n5229), .ZN(n5235) );
  INV_X1 U6610 ( .A(n5228), .ZN(n5231) );
  INV_X1 U6611 ( .A(n5229), .ZN(n5230) );
  NAND2_X1 U6612 ( .A1(n5231), .A2(n5230), .ZN(n5232) );
  NAND2_X1 U6613 ( .A1(n5235), .A2(n5232), .ZN(n7658) );
  INV_X1 U6614 ( .A(n7658), .ZN(n5233) );
  NAND2_X1 U6615 ( .A1(n5234), .A2(n5233), .ZN(n7655) );
  INV_X1 U6616 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6650) );
  MUX2_X1 U6617 ( .A(n6650), .B(n10148), .S(n5601), .Z(n5241) );
  INV_X1 U6618 ( .A(SI_10_), .ZN(n5240) );
  INV_X1 U6619 ( .A(n5241), .ZN(n5242) );
  NAND2_X1 U6620 ( .A1(n5242), .A2(SI_10_), .ZN(n5243) );
  OR2_X1 U6621 ( .A1(n5244), .A2(n4924), .ZN(n5245) );
  NAND2_X1 U6622 ( .A1(n5264), .A2(n5245), .ZN(n6648) );
  NAND2_X1 U6623 ( .A1(n6648), .A2(n8389), .ZN(n5248) );
  NAND2_X1 U6624 ( .A1(n5310), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5265) );
  XNOR2_X1 U6625 ( .A(n5265), .B(P1_IR_REG_10__SCAN_IN), .ZN(n6849) );
  AOI22_X1 U6626 ( .A1(n5506), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n9601), .B2(
        n6849), .ZN(n5247) );
  NAND2_X1 U6627 ( .A1(n9504), .A2(n6492), .ZN(n5256) );
  NAND2_X1 U6628 ( .A1(n8287), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5254) );
  NAND2_X1 U6629 ( .A1(n8288), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5253) );
  INV_X1 U6630 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n6692) );
  NAND2_X1 U6631 ( .A1(n5249), .A2(n6692), .ZN(n5250) );
  AND2_X1 U6632 ( .A1(n5272), .A2(n5250), .ZN(n9503) );
  NAND2_X1 U6633 ( .A1(n5758), .A2(n9503), .ZN(n5252) );
  NAND2_X1 U6634 ( .A1(n8289), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5251) );
  NAND4_X1 U6635 ( .A1(n5254), .A2(n5253), .A3(n5252), .A4(n5251), .ZN(n9082)
         );
  NAND2_X1 U6636 ( .A1(n9082), .A2(n4398), .ZN(n5255) );
  NAND2_X1 U6637 ( .A1(n5256), .A2(n5255), .ZN(n5257) );
  XNOR2_X1 U6638 ( .A(n5257), .B(n6490), .ZN(n5262) );
  INV_X1 U6639 ( .A(n5262), .ZN(n5260) );
  AND2_X1 U6640 ( .A1(n9082), .A2(n5640), .ZN(n5258) );
  AOI21_X1 U6641 ( .B1(n9504), .B2(n4398), .A(n5258), .ZN(n5261) );
  INV_X1 U6642 ( .A(n5261), .ZN(n5259) );
  NAND2_X1 U6643 ( .A1(n5260), .A2(n5259), .ZN(n7713) );
  INV_X1 U6644 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n10222) );
  MUX2_X1 U6645 ( .A(n10222), .B(n10150), .S(n4973), .Z(n5291) );
  XNOR2_X1 U6646 ( .A(n5348), .B(n5285), .ZN(n6651) );
  NAND2_X1 U6647 ( .A1(n6651), .A2(n8389), .ZN(n5269) );
  INV_X1 U6648 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5308) );
  NAND2_X1 U6649 ( .A1(n5265), .A2(n5308), .ZN(n5266) );
  NAND2_X1 U6650 ( .A1(n5266), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5267) );
  XNOR2_X1 U6651 ( .A(n5267), .B(P1_IR_REG_11__SCAN_IN), .ZN(n9672) );
  AOI22_X1 U6652 ( .A1(n5506), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n9601), .B2(
        n9672), .ZN(n5268) );
  NAND2_X1 U6653 ( .A1(n7782), .A2(n6492), .ZN(n5279) );
  NAND2_X1 U6654 ( .A1(n8289), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5277) );
  NAND2_X1 U6655 ( .A1(n8287), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5276) );
  INV_X1 U6656 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5271) );
  NAND2_X1 U6657 ( .A1(n5272), .A2(n5271), .ZN(n5273) );
  AND2_X1 U6658 ( .A1(n5333), .A2(n5273), .ZN(n7823) );
  NAND2_X1 U6659 ( .A1(n5758), .A2(n7823), .ZN(n5275) );
  NAND2_X1 U6660 ( .A1(n8288), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5274) );
  NAND4_X1 U6661 ( .A1(n5277), .A2(n5276), .A3(n5275), .A4(n5274), .ZN(n9496)
         );
  NAND2_X1 U6662 ( .A1(n9496), .A2(n5096), .ZN(n5278) );
  NAND2_X1 U6663 ( .A1(n5279), .A2(n5278), .ZN(n5280) );
  XNOR2_X1 U6664 ( .A(n5280), .B(n7160), .ZN(n5284) );
  AND2_X1 U6665 ( .A1(n9496), .A2(n5640), .ZN(n5281) );
  AOI21_X1 U6666 ( .B1(n7782), .B2(n5096), .A(n5281), .ZN(n5282) );
  XNOR2_X1 U6667 ( .A(n5284), .B(n5282), .ZN(n7819) );
  INV_X1 U6668 ( .A(n5282), .ZN(n5283) );
  NAND2_X1 U6669 ( .A1(n5284), .A2(n5283), .ZN(n7857) );
  INV_X1 U6670 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6689) );
  INV_X1 U6671 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6691) );
  MUX2_X1 U6672 ( .A(n6689), .B(n6691), .S(n4973), .Z(n5287) );
  INV_X1 U6673 ( .A(SI_12_), .ZN(n5286) );
  NOR2_X1 U6674 ( .A1(n5348), .A2(n5346), .ZN(n5304) );
  INV_X1 U6675 ( .A(n5287), .ZN(n5288) );
  NAND2_X1 U6676 ( .A1(n5288), .A2(SI_12_), .ZN(n5289) );
  NAND2_X1 U6677 ( .A1(n5290), .A2(n5289), .ZN(n5328) );
  INV_X1 U6678 ( .A(n5328), .ZN(n5293) );
  INV_X1 U6679 ( .A(n5291), .ZN(n5292) );
  NAND2_X1 U6680 ( .A1(n5292), .A2(SI_11_), .ZN(n5327) );
  OR2_X1 U6681 ( .A1(n5304), .A2(n5302), .ZN(n5301) );
  INV_X1 U6682 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n5296) );
  MUX2_X1 U6683 ( .A(n10216), .B(n5296), .S(n5601), .Z(n5298) );
  INV_X1 U6684 ( .A(SI_13_), .ZN(n5297) );
  INV_X1 U6685 ( .A(n5298), .ZN(n5299) );
  NAND2_X1 U6686 ( .A1(n5299), .A2(SI_13_), .ZN(n5300) );
  NAND2_X1 U6687 ( .A1(n5350), .A2(n5300), .ZN(n5303) );
  NAND2_X1 U6688 ( .A1(n5301), .A2(n5303), .ZN(n5306) );
  OR2_X1 U6689 ( .A1(n5304), .A2(n5349), .ZN(n5305) );
  NAND2_X1 U6690 ( .A1(n5306), .A2(n5305), .ZN(n6653) );
  NAND2_X1 U6691 ( .A1(n6653), .A2(n8389), .ZN(n5314) );
  INV_X1 U6692 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n5307) );
  NAND2_X1 U6693 ( .A1(n5308), .A2(n5307), .ZN(n5309) );
  NOR2_X1 U6694 ( .A1(n5310), .A2(n5309), .ZN(n5330) );
  NAND2_X1 U6695 ( .A1(n5330), .A2(n5311), .ZN(n5351) );
  NAND2_X1 U6696 ( .A1(n5351), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5312) );
  XNOR2_X1 U6697 ( .A(n5312), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7403) );
  AOI22_X1 U6698 ( .A1(n5506), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n9601), .B2(
        n7403), .ZN(n5313) );
  NAND2_X1 U6699 ( .A1(n7959), .A2(n6492), .ZN(n5322) );
  NAND2_X1 U6700 ( .A1(n8287), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5320) );
  NAND2_X1 U6701 ( .A1(n8288), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5319) );
  INV_X1 U6702 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n6842) );
  INV_X1 U6703 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5315) );
  NAND2_X1 U6704 ( .A1(n5335), .A2(n5315), .ZN(n5316) );
  AND2_X1 U6705 ( .A1(n5356), .A2(n5316), .ZN(n8020) );
  NAND2_X1 U6706 ( .A1(n5758), .A2(n8020), .ZN(n5318) );
  NAND2_X1 U6707 ( .A1(n8289), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5317) );
  NAND4_X1 U6708 ( .A1(n5320), .A2(n5319), .A3(n5318), .A4(n5317), .ZN(n9080)
         );
  NAND2_X1 U6709 ( .A1(n9080), .A2(n4398), .ZN(n5321) );
  NAND2_X1 U6710 ( .A1(n5322), .A2(n5321), .ZN(n5323) );
  XNOR2_X1 U6711 ( .A(n5323), .B(n7160), .ZN(n5372) );
  NAND2_X1 U6712 ( .A1(n7959), .A2(n5096), .ZN(n5325) );
  NAND2_X1 U6713 ( .A1(n9080), .A2(n5640), .ZN(n5324) );
  NAND2_X1 U6714 ( .A1(n5325), .A2(n5324), .ZN(n5373) );
  INV_X1 U6715 ( .A(n8010), .ZN(n5344) );
  XNOR2_X1 U6716 ( .A(n5329), .B(n5328), .ZN(n6688) );
  OR2_X1 U6717 ( .A1(n5330), .A2(n9456), .ZN(n5331) );
  XNOR2_X1 U6718 ( .A(n5331), .B(P1_IR_REG_12__SCAN_IN), .ZN(n6974) );
  AOI22_X1 U6719 ( .A1(n5506), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n9601), .B2(
        n6974), .ZN(n5332) );
  NAND2_X1 U6720 ( .A1(n8287), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5339) );
  NAND2_X1 U6721 ( .A1(n8288), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5338) );
  NAND2_X1 U6722 ( .A1(n5333), .A2(n6842), .ZN(n5334) );
  AND2_X1 U6723 ( .A1(n5335), .A2(n5334), .ZN(n7862) );
  NAND2_X1 U6724 ( .A1(n5758), .A2(n7862), .ZN(n5337) );
  NAND2_X1 U6725 ( .A1(n8289), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5336) );
  NAND4_X1 U6726 ( .A1(n5339), .A2(n5338), .A3(n5337), .A4(n5336), .ZN(n9081)
         );
  NAND2_X1 U6727 ( .A1(n9081), .A2(n5096), .ZN(n5340) );
  XNOR2_X1 U6728 ( .A(n5341), .B(n6490), .ZN(n7859) );
  INV_X1 U6729 ( .A(n7859), .ZN(n5343) );
  AND2_X1 U6730 ( .A1(n9081), .A2(n5640), .ZN(n5342) );
  AOI21_X1 U6731 ( .B1(n7930), .B2(n4398), .A(n5342), .ZN(n5369) );
  INV_X1 U6732 ( .A(n5369), .ZN(n7858) );
  NAND2_X1 U6733 ( .A1(n5343), .A2(n7858), .ZN(n8006) );
  INV_X1 U6734 ( .A(n5350), .ZN(n5345) );
  INV_X1 U6735 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6659) );
  INV_X1 U6736 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6657) );
  MUX2_X1 U6737 ( .A(n6659), .B(n6657), .S(n5447), .Z(n5383) );
  XNOR2_X1 U6738 ( .A(n5383), .B(SI_14_), .ZN(n5382) );
  XNOR2_X1 U6739 ( .A(n5385), .B(n5382), .ZN(n6656) );
  NAND2_X1 U6740 ( .A1(n6656), .A2(n8389), .ZN(n5353) );
  NAND2_X1 U6741 ( .A1(n5423), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5390) );
  XNOR2_X1 U6742 ( .A(n5390), .B(P1_IR_REG_14__SCAN_IN), .ZN(n7773) );
  AOI22_X1 U6743 ( .A1(n9601), .A2(n7773), .B1(n5506), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n5352) );
  NAND2_X1 U6744 ( .A1(n8048), .A2(n6492), .ZN(n5363) );
  NAND2_X1 U6745 ( .A1(n8289), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5361) );
  NAND2_X1 U6746 ( .A1(n8287), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5360) );
  INV_X1 U6747 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5355) );
  NAND2_X1 U6748 ( .A1(n5356), .A2(n5355), .ZN(n5357) );
  AND2_X1 U6749 ( .A1(n5398), .A2(n5357), .ZN(n7990) );
  NAND2_X1 U6750 ( .A1(n5758), .A2(n7990), .ZN(n5359) );
  NAND2_X1 U6751 ( .A1(n8288), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5358) );
  NAND4_X1 U6752 ( .A1(n5361), .A2(n5360), .A3(n5359), .A4(n5358), .ZN(n9079)
         );
  NAND2_X1 U6753 ( .A1(n9079), .A2(n4398), .ZN(n5362) );
  NAND2_X1 U6754 ( .A1(n5363), .A2(n5362), .ZN(n5364) );
  XNOR2_X1 U6755 ( .A(n5364), .B(n6490), .ZN(n5368) );
  AND2_X1 U6756 ( .A1(n5377), .A2(n5368), .ZN(n5365) );
  NAND2_X1 U6757 ( .A1(n7817), .A2(n5365), .ZN(n7980) );
  NAND2_X1 U6758 ( .A1(n8048), .A2(n5096), .ZN(n5367) );
  NAND2_X1 U6759 ( .A1(n9079), .A2(n5640), .ZN(n5366) );
  NAND2_X1 U6760 ( .A1(n5367), .A2(n5366), .ZN(n7981) );
  INV_X1 U6761 ( .A(n5368), .ZN(n5379) );
  NAND2_X1 U6762 ( .A1(n7859), .A2(n5369), .ZN(n8004) );
  INV_X1 U6763 ( .A(n8004), .ZN(n5370) );
  INV_X1 U6764 ( .A(n5372), .ZN(n5375) );
  INV_X1 U6765 ( .A(n5373), .ZN(n5374) );
  NAND2_X1 U6766 ( .A1(n5375), .A2(n5374), .ZN(n8008) );
  NAND2_X1 U6767 ( .A1(n7980), .A2(n5376), .ZN(n7978) );
  INV_X1 U6768 ( .A(n5383), .ZN(n5384) );
  INV_X1 U6769 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6758) );
  INV_X1 U6770 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6760) );
  MUX2_X1 U6771 ( .A(n6758), .B(n6760), .S(n5447), .Z(n5387) );
  INV_X1 U6772 ( .A(SI_15_), .ZN(n5386) );
  NAND2_X1 U6773 ( .A1(n5387), .A2(n5386), .ZN(n5413) );
  INV_X1 U6774 ( .A(n5387), .ZN(n5388) );
  NAND2_X1 U6775 ( .A1(n5388), .A2(SI_15_), .ZN(n5389) );
  NAND2_X1 U6776 ( .A1(n5413), .A2(n5389), .ZN(n5414) );
  XNOR2_X1 U6777 ( .A(n5415), .B(n5414), .ZN(n6757) );
  NAND2_X1 U6778 ( .A1(n6757), .A2(n8389), .ZN(n5395) );
  INV_X1 U6779 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5420) );
  NAND2_X1 U6780 ( .A1(n5390), .A2(n5420), .ZN(n5391) );
  NAND2_X1 U6781 ( .A1(n5391), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5392) );
  XNOR2_X1 U6782 ( .A(n5392), .B(n5421), .ZN(n7890) );
  OAI22_X1 U6783 ( .A1(n7890), .A2(n5042), .B1(n8391), .B2(n6760), .ZN(n5393)
         );
  INV_X1 U6784 ( .A(n5393), .ZN(n5394) );
  NAND2_X1 U6785 ( .A1(n9117), .A2(n6492), .ZN(n5405) );
  NAND2_X1 U6786 ( .A1(n8289), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5403) );
  NAND2_X1 U6787 ( .A1(n8287), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5402) );
  INV_X1 U6788 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n5397) );
  NAND2_X1 U6789 ( .A1(n5398), .A2(n5397), .ZN(n5399) );
  AND2_X1 U6790 ( .A1(n5427), .A2(n5399), .ZN(n8054) );
  NAND2_X1 U6791 ( .A1(n5758), .A2(n8054), .ZN(n5401) );
  NAND2_X1 U6792 ( .A1(n5154), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5400) );
  NAND4_X1 U6793 ( .A1(n5403), .A2(n5402), .A3(n5401), .A4(n5400), .ZN(n9538)
         );
  NAND2_X1 U6794 ( .A1(n9538), .A2(n4398), .ZN(n5404) );
  NAND2_X1 U6795 ( .A1(n5405), .A2(n5404), .ZN(n5406) );
  XNOR2_X1 U6796 ( .A(n5406), .B(n6490), .ZN(n5409) );
  NAND3_X1 U6797 ( .A1(n7978), .A2(n7983), .A3(n5409), .ZN(n7993) );
  NAND2_X1 U6798 ( .A1(n9117), .A2(n5096), .ZN(n5408) );
  NAND2_X1 U6799 ( .A1(n9538), .A2(n5640), .ZN(n5407) );
  NAND2_X1 U6800 ( .A1(n5408), .A2(n5407), .ZN(n7996) );
  NAND2_X1 U6801 ( .A1(n7993), .A2(n7996), .ZN(n5412) );
  NAND2_X1 U6802 ( .A1(n7978), .A2(n7983), .ZN(n5411) );
  INV_X1 U6803 ( .A(n5409), .ZN(n5410) );
  NAND2_X1 U6804 ( .A1(n5411), .A2(n5410), .ZN(n7994) );
  INV_X1 U6805 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n6773) );
  INV_X1 U6806 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n6762) );
  MUX2_X1 U6807 ( .A(n6773), .B(n6762), .S(n5601), .Z(n5417) );
  INV_X1 U6808 ( .A(SI_16_), .ZN(n5416) );
  NAND2_X1 U6809 ( .A1(n5417), .A2(n5416), .ZN(n5445) );
  INV_X1 U6810 ( .A(n5417), .ZN(n5418) );
  NAND2_X1 U6811 ( .A1(n5418), .A2(SI_16_), .ZN(n5419) );
  XNOR2_X1 U6812 ( .A(n5444), .B(n5443), .ZN(n6761) );
  NAND2_X1 U6813 ( .A1(n6761), .A2(n8389), .ZN(n5426) );
  NAND2_X1 U6814 ( .A1(n5421), .A2(n5420), .ZN(n5422) );
  NOR2_X1 U6815 ( .A1(n5423), .A2(n5422), .ZN(n5450) );
  OR2_X1 U6816 ( .A1(n5450), .A2(n9456), .ZN(n5424) );
  XNOR2_X1 U6817 ( .A(n5424), .B(P1_IR_REG_16__SCAN_IN), .ZN(n8103) );
  AOI22_X1 U6818 ( .A1(n8103), .A2(n9601), .B1(n5506), .B2(
        P2_DATAO_REG_16__SCAN_IN), .ZN(n5425) );
  NAND2_X1 U6819 ( .A1(n9544), .A2(n6492), .ZN(n5434) );
  NAND2_X1 U6820 ( .A1(n8287), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n5432) );
  NAND2_X1 U6821 ( .A1(n8289), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5431) );
  INV_X1 U6822 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n7896) );
  NAND2_X1 U6823 ( .A1(n5427), .A2(n7896), .ZN(n5428) );
  AND2_X1 U6824 ( .A1(n5458), .A2(n5428), .ZN(n9542) );
  NAND2_X1 U6825 ( .A1(n5758), .A2(n9542), .ZN(n5430) );
  NAND2_X1 U6826 ( .A1(n8288), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5429) );
  NAND4_X1 U6827 ( .A1(n5432), .A2(n5431), .A3(n5430), .A4(n5429), .ZN(n9361)
         );
  NAND2_X1 U6828 ( .A1(n9361), .A2(n4398), .ZN(n5433) );
  NAND2_X1 U6829 ( .A1(n5434), .A2(n5433), .ZN(n5435) );
  XNOR2_X1 U6830 ( .A(n5435), .B(n7160), .ZN(n5439) );
  NAND2_X1 U6831 ( .A1(n9544), .A2(n5096), .ZN(n5437) );
  NAND2_X1 U6832 ( .A1(n9361), .A2(n5640), .ZN(n5436) );
  NAND2_X1 U6833 ( .A1(n5437), .A2(n5436), .ZN(n5440) );
  AND2_X1 U6834 ( .A1(n5439), .A2(n5440), .ZN(n8139) );
  INV_X1 U6835 ( .A(n8139), .ZN(n5438) );
  INV_X1 U6836 ( .A(n5439), .ZN(n5442) );
  INV_X1 U6837 ( .A(n5440), .ZN(n5441) );
  NAND2_X1 U6838 ( .A1(n5442), .A2(n5441), .ZN(n8137) );
  INV_X1 U6839 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n10113) );
  INV_X1 U6840 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n5448) );
  MUX2_X1 U6841 ( .A(n10113), .B(n5448), .S(n5601), .Z(n5472) );
  XNOR2_X1 U6842 ( .A(n5472), .B(SI_17_), .ZN(n5471) );
  XNOR2_X1 U6843 ( .A(n5476), .B(n5471), .ZN(n6797) );
  NAND2_X1 U6844 ( .A1(n6797), .A2(n8389), .ZN(n5453) );
  INV_X1 U6845 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5449) );
  NAND2_X1 U6846 ( .A1(n5450), .A2(n5449), .ZN(n5451) );
  NAND2_X1 U6847 ( .A1(n5451), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5478) );
  XNOR2_X1 U6848 ( .A(n5478), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9095) );
  AOI22_X1 U6849 ( .A1(n9095), .A2(n9601), .B1(n5506), .B2(
        P2_DATAO_REG_17__SCAN_IN), .ZN(n5452) );
  NAND2_X1 U6850 ( .A1(n9435), .A2(n6492), .ZN(n5464) );
  INV_X1 U6851 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n5462) );
  NAND2_X1 U6852 ( .A1(n8287), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n5455) );
  NAND2_X1 U6853 ( .A1(n8289), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5454) );
  AND2_X1 U6854 ( .A1(n5455), .A2(n5454), .ZN(n5461) );
  INV_X1 U6855 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n5457) );
  NAND2_X1 U6856 ( .A1(n5458), .A2(n5457), .ZN(n5459) );
  NAND2_X1 U6857 ( .A1(n5485), .A2(n5459), .ZN(n8163) );
  OR2_X1 U6858 ( .A1(n8163), .A2(n6500), .ZN(n5460) );
  OAI211_X1 U6859 ( .C1(n5709), .C2(n5462), .A(n5461), .B(n5460), .ZN(n9539)
         );
  NAND2_X1 U6860 ( .A1(n9539), .A2(n5096), .ZN(n5463) );
  NAND2_X1 U6861 ( .A1(n5464), .A2(n5463), .ZN(n5465) );
  XNOR2_X1 U6862 ( .A(n5465), .B(n7160), .ZN(n5467) );
  AND2_X1 U6863 ( .A1(n9539), .A2(n5640), .ZN(n5466) );
  AOI21_X1 U6864 ( .B1(n9435), .B2(n4398), .A(n5466), .ZN(n5468) );
  XNOR2_X1 U6865 ( .A(n5467), .B(n5468), .ZN(n8161) );
  NAND2_X1 U6866 ( .A1(n8160), .A2(n8161), .ZN(n8159) );
  INV_X1 U6867 ( .A(n5467), .ZN(n5469) );
  NAND2_X1 U6868 ( .A1(n5469), .A2(n5468), .ZN(n5470) );
  INV_X1 U6869 ( .A(n5471), .ZN(n5475) );
  INV_X1 U6870 ( .A(n5472), .ZN(n5473) );
  NAND2_X1 U6871 ( .A1(n5473), .A2(SI_17_), .ZN(n5474) );
  OAI21_X2 U6872 ( .B1(n5476), .B2(n5475), .A(n5474), .ZN(n5497) );
  MUX2_X1 U6873 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n5447), .Z(n5498) );
  XNOR2_X1 U6874 ( .A(n5498), .B(SI_18_), .ZN(n5495) );
  XNOR2_X1 U6875 ( .A(n5497), .B(n5495), .ZN(n6872) );
  NAND2_X1 U6876 ( .A1(n6872), .A2(n8389), .ZN(n5483) );
  NAND2_X1 U6877 ( .A1(n5478), .A2(n5477), .ZN(n5479) );
  NAND2_X1 U6878 ( .A1(n5479), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5480) );
  XNOR2_X1 U6879 ( .A(n5480), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9685) );
  INV_X1 U6880 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n10186) );
  NOR2_X1 U6881 ( .A1(n8391), .A2(n10186), .ZN(n5481) );
  AOI21_X1 U6882 ( .B1(n9685), .B2(n9601), .A(n5481), .ZN(n5482) );
  NAND2_X1 U6883 ( .A1(n9432), .A2(n6492), .ZN(n5490) );
  INV_X1 U6884 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n5484) );
  NAND2_X1 U6885 ( .A1(n5485), .A2(n5484), .ZN(n5486) );
  NAND2_X1 U6886 ( .A1(n5531), .A2(n5486), .ZN(n9335) );
  AOI22_X1 U6887 ( .A1(n8287), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n5154), .B2(
        P1_REG2_REG_18__SCAN_IN), .ZN(n5488) );
  NAND2_X1 U6888 ( .A1(n8289), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n5487) );
  OAI211_X1 U6889 ( .C1(n9335), .C2(n6500), .A(n5488), .B(n5487), .ZN(n9362)
         );
  NAND2_X1 U6890 ( .A1(n9362), .A2(n4398), .ZN(n5489) );
  NAND2_X1 U6891 ( .A1(n5490), .A2(n5489), .ZN(n5491) );
  XNOR2_X1 U6892 ( .A(n5491), .B(n6490), .ZN(n5494) );
  NAND2_X1 U6893 ( .A1(n9432), .A2(n5096), .ZN(n5493) );
  NAND2_X1 U6894 ( .A1(n9362), .A2(n5640), .ZN(n5492) );
  NAND2_X1 U6895 ( .A1(n5493), .A2(n5492), .ZN(n9053) );
  INV_X1 U6896 ( .A(n5495), .ZN(n5496) );
  NAND2_X1 U6897 ( .A1(n5498), .A2(SI_18_), .ZN(n5499) );
  INV_X1 U6898 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n6990) );
  INV_X1 U6899 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n6988) );
  MUX2_X1 U6900 ( .A(n6990), .B(n6988), .S(n5447), .Z(n5502) );
  INV_X1 U6901 ( .A(SI_19_), .ZN(n5501) );
  NAND2_X1 U6902 ( .A1(n5502), .A2(n5501), .ZN(n5523) );
  INV_X1 U6903 ( .A(n5502), .ZN(n5503) );
  NAND2_X1 U6904 ( .A1(n5503), .A2(SI_19_), .ZN(n5504) );
  NAND2_X1 U6905 ( .A1(n5523), .A2(n5504), .ZN(n5521) );
  XNOR2_X1 U6906 ( .A(n5522), .B(n5521), .ZN(n6987) );
  NAND2_X1 U6907 ( .A1(n6987), .A2(n8389), .ZN(n5508) );
  AOI22_X1 U6908 ( .A1(n5506), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n5505), .B2(
        n9601), .ZN(n5507) );
  NAND2_X1 U6909 ( .A1(n9425), .A2(n6492), .ZN(n5515) );
  XNOR2_X1 U6910 ( .A(n5531), .B(P1_REG3_REG_19__SCAN_IN), .ZN(n9319) );
  NAND2_X1 U6911 ( .A1(n9319), .A2(n5758), .ZN(n5513) );
  INV_X1 U6912 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n10226) );
  NAND2_X1 U6913 ( .A1(n8287), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n5510) );
  NAND2_X1 U6914 ( .A1(n8288), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n5509) );
  OAI211_X1 U6915 ( .C1(n5063), .C2(n10226), .A(n5510), .B(n5509), .ZN(n5511)
         );
  INV_X1 U6916 ( .A(n5511), .ZN(n5512) );
  NAND2_X1 U6917 ( .A1(n5513), .A2(n5512), .ZN(n9309) );
  NAND2_X1 U6918 ( .A1(n9309), .A2(n5096), .ZN(n5514) );
  NAND2_X1 U6919 ( .A1(n5515), .A2(n5514), .ZN(n5516) );
  XNOR2_X1 U6920 ( .A(n5516), .B(n7160), .ZN(n8986) );
  NAND2_X1 U6921 ( .A1(n9425), .A2(n4398), .ZN(n5518) );
  NAND2_X1 U6922 ( .A1(n9309), .A2(n5640), .ZN(n5517) );
  NAND2_X1 U6923 ( .A1(n5518), .A2(n5517), .ZN(n8987) );
  OAI21_X1 U6924 ( .B1(n8985), .B2(n8986), .A(n8987), .ZN(n5520) );
  NAND2_X1 U6925 ( .A1(n8985), .A2(n8986), .ZN(n5519) );
  NAND2_X1 U6926 ( .A1(n5520), .A2(n5519), .ZN(n9029) );
  INV_X1 U6927 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n10057) );
  INV_X1 U6928 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n9998) );
  MUX2_X1 U6929 ( .A(n10057), .B(n9998), .S(n5601), .Z(n5525) );
  INV_X1 U6930 ( .A(SI_20_), .ZN(n5524) );
  NAND2_X1 U6931 ( .A1(n5525), .A2(n5524), .ZN(n5552) );
  INV_X1 U6932 ( .A(n5525), .ZN(n5526) );
  NAND2_X1 U6933 ( .A1(n5526), .A2(SI_20_), .ZN(n5527) );
  AND2_X1 U6934 ( .A1(n5552), .A2(n5527), .ZN(n5550) );
  XNOR2_X1 U6935 ( .A(n5551), .B(n5550), .ZN(n7123) );
  NAND2_X1 U6936 ( .A1(n7123), .A2(n8389), .ZN(n5529) );
  OR2_X1 U6937 ( .A1(n8391), .A2(n9998), .ZN(n5528) );
  NAND2_X1 U6938 ( .A1(n9420), .A2(n6492), .ZN(n5542) );
  INV_X1 U6939 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n10119) );
  INV_X1 U6940 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n5530) );
  OAI21_X1 U6941 ( .B1(n5531), .B2(n10119), .A(n5530), .ZN(n5534) );
  AND2_X1 U6942 ( .A1(P1_REG3_REG_19__SCAN_IN), .A2(P1_REG3_REG_20__SCAN_IN), 
        .ZN(n5532) );
  NAND2_X1 U6943 ( .A1(n5534), .A2(n5557), .ZN(n9303) );
  OR2_X1 U6944 ( .A1(n9303), .A2(n6500), .ZN(n5540) );
  INV_X1 U6945 ( .A(n8287), .ZN(n5689) );
  INV_X1 U6946 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n5537) );
  NAND2_X1 U6947 ( .A1(n8289), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n5536) );
  NAND2_X1 U6948 ( .A1(n8288), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n5535) );
  OAI211_X1 U6949 ( .C1(n5689), .C2(n5537), .A(n5536), .B(n5535), .ZN(n5538)
         );
  INV_X1 U6950 ( .A(n5538), .ZN(n5539) );
  NAND2_X1 U6951 ( .A1(n5540), .A2(n5539), .ZN(n9327) );
  NAND2_X1 U6952 ( .A1(n9327), .A2(n5096), .ZN(n5541) );
  NAND2_X1 U6953 ( .A1(n5542), .A2(n5541), .ZN(n5543) );
  XNOR2_X1 U6954 ( .A(n5543), .B(n7160), .ZN(n5546) );
  NAND2_X1 U6955 ( .A1(n9420), .A2(n5096), .ZN(n5545) );
  NAND2_X1 U6956 ( .A1(n9327), .A2(n5640), .ZN(n5544) );
  NAND2_X1 U6957 ( .A1(n5545), .A2(n5544), .ZN(n5547) );
  INV_X1 U6958 ( .A(n5546), .ZN(n5549) );
  INV_X1 U6959 ( .A(n5547), .ZN(n5548) );
  NAND2_X1 U6960 ( .A1(n5549), .A2(n5548), .ZN(n9032) );
  INV_X1 U6961 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7172) );
  INV_X1 U6962 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n8558) );
  MUX2_X1 U6963 ( .A(n7172), .B(n8558), .S(n5447), .Z(n5574) );
  XNOR2_X1 U6964 ( .A(n5574), .B(SI_21_), .ZN(n5573) );
  XNOR2_X1 U6965 ( .A(n5578), .B(n5573), .ZN(n7170) );
  NAND2_X1 U6966 ( .A1(n7170), .A2(n8389), .ZN(n5555) );
  OR2_X1 U6967 ( .A1(n8391), .A2(n8558), .ZN(n5554) );
  NAND2_X1 U6968 ( .A1(n9417), .A2(n6492), .ZN(n5566) );
  INV_X1 U6969 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n5556) );
  NAND2_X1 U6970 ( .A1(n5557), .A2(n5556), .ZN(n5558) );
  AND2_X1 U6971 ( .A1(n5616), .A2(n5558), .ZN(n9295) );
  NAND2_X1 U6972 ( .A1(n9295), .A2(n5758), .ZN(n5564) );
  INV_X1 U6973 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n5561) );
  NAND2_X1 U6974 ( .A1(n8289), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5560) );
  NAND2_X1 U6975 ( .A1(n8288), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n5559) );
  OAI211_X1 U6976 ( .C1(n5689), .C2(n5561), .A(n5560), .B(n5559), .ZN(n5562)
         );
  INV_X1 U6977 ( .A(n5562), .ZN(n5563) );
  NAND2_X1 U6978 ( .A1(n5564), .A2(n5563), .ZN(n9310) );
  NAND2_X1 U6979 ( .A1(n9310), .A2(n4398), .ZN(n5565) );
  NAND2_X1 U6980 ( .A1(n5566), .A2(n5565), .ZN(n5567) );
  XNOR2_X1 U6981 ( .A(n5567), .B(n7160), .ZN(n5569) );
  AND2_X1 U6982 ( .A1(n9310), .A2(n5640), .ZN(n5568) );
  AOI21_X1 U6983 ( .B1(n9417), .B2(n5096), .A(n5568), .ZN(n5570) );
  XNOR2_X1 U6984 ( .A(n5569), .B(n5570), .ZN(n8995) );
  INV_X1 U6985 ( .A(n5569), .ZN(n5571) );
  NAND2_X1 U6986 ( .A1(n5571), .A2(n5570), .ZN(n5572) );
  INV_X1 U6987 ( .A(n5573), .ZN(n5577) );
  INV_X1 U6988 ( .A(n5574), .ZN(n5575) );
  NAND2_X1 U6989 ( .A1(n5575), .A2(SI_21_), .ZN(n5576) );
  OAI21_X2 U6990 ( .B1(n5578), .B2(n5577), .A(n5576), .ZN(n5600) );
  INV_X1 U6991 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7434) );
  INV_X1 U6992 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n10098) );
  MUX2_X1 U6993 ( .A(n7434), .B(n10098), .S(n5601), .Z(n5580) );
  INV_X1 U6994 ( .A(SI_22_), .ZN(n5579) );
  NAND2_X1 U6995 ( .A1(n5580), .A2(n5579), .ZN(n5598) );
  INV_X1 U6996 ( .A(n5580), .ZN(n5581) );
  NAND2_X1 U6997 ( .A1(n5581), .A2(SI_22_), .ZN(n5582) );
  NAND2_X1 U6998 ( .A1(n5598), .A2(n5582), .ZN(n5599) );
  XNOR2_X1 U6999 ( .A(n5600), .B(n5599), .ZN(n7432) );
  NAND2_X1 U7000 ( .A1(n7432), .A2(n8389), .ZN(n5584) );
  OR2_X1 U7001 ( .A1(n8391), .A2(n10098), .ZN(n5583) );
  XNOR2_X1 U7002 ( .A(n5616), .B(P1_REG3_REG_22__SCAN_IN), .ZN(n9275) );
  NAND2_X1 U7003 ( .A1(n9275), .A2(n5758), .ZN(n5590) );
  INV_X1 U7004 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n5587) );
  NAND2_X1 U7005 ( .A1(n8289), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5586) );
  NAND2_X1 U7006 ( .A1(n8288), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n5585) );
  OAI211_X1 U7007 ( .C1(n5689), .C2(n5587), .A(n5586), .B(n5585), .ZN(n5588)
         );
  INV_X1 U7008 ( .A(n5588), .ZN(n5589) );
  NAND2_X1 U7009 ( .A1(n5590), .A2(n5589), .ZN(n9258) );
  AND2_X1 U7010 ( .A1(n9258), .A2(n5640), .ZN(n5591) );
  AOI21_X1 U7011 ( .B1(n9410), .B2(n5096), .A(n5591), .ZN(n5596) );
  INV_X1 U7012 ( .A(n5596), .ZN(n5592) );
  NAND2_X1 U7013 ( .A1(n9410), .A2(n6492), .ZN(n5594) );
  NAND2_X1 U7014 ( .A1(n9258), .A2(n5096), .ZN(n5593) );
  NAND2_X1 U7015 ( .A1(n5594), .A2(n5593), .ZN(n5595) );
  XNOR2_X1 U7016 ( .A(n5595), .B(n6490), .ZN(n9042) );
  NAND2_X1 U7017 ( .A1(n9044), .A2(n9042), .ZN(n9040) );
  INV_X1 U7018 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n5602) );
  INV_X1 U7019 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n5609) );
  MUX2_X1 U7020 ( .A(n5602), .B(n5609), .S(n5447), .Z(n5603) );
  INV_X1 U7021 ( .A(SI_23_), .ZN(n10063) );
  NAND2_X1 U7022 ( .A1(n5603), .A2(n10063), .ZN(n5628) );
  INV_X1 U7023 ( .A(n5603), .ZN(n5604) );
  NAND2_X1 U7024 ( .A1(n5604), .A2(SI_23_), .ZN(n5605) );
  AND2_X1 U7025 ( .A1(n5628), .A2(n5605), .ZN(n5606) );
  OR2_X1 U7027 ( .A1(n5607), .A2(n5606), .ZN(n5608) );
  NAND2_X1 U7028 ( .A1(n5629), .A2(n5608), .ZN(n7446) );
  NAND2_X1 U7029 ( .A1(n7446), .A2(n8389), .ZN(n5611) );
  OR2_X1 U7030 ( .A1(n8391), .A2(n5609), .ZN(n5610) );
  NAND2_X1 U7031 ( .A1(n9407), .A2(n6492), .ZN(n5625) );
  AND2_X1 U7032 ( .A1(P1_REG3_REG_22__SCAN_IN), .A2(P1_REG3_REG_23__SCAN_IN), 
        .ZN(n5612) );
  INV_X1 U7033 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n5615) );
  INV_X1 U7034 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n5614) );
  OAI21_X1 U7035 ( .B1(n5616), .B2(n5615), .A(n5614), .ZN(n5617) );
  NAND2_X1 U7036 ( .A1(n5632), .A2(n5617), .ZN(n9266) );
  OR2_X1 U7037 ( .A1(n9266), .A2(n6500), .ZN(n5623) );
  INV_X1 U7038 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n5620) );
  NAND2_X1 U7039 ( .A1(n8289), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5619) );
  NAND2_X1 U7040 ( .A1(n5154), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n5618) );
  OAI211_X1 U7041 ( .C1(n5689), .C2(n5620), .A(n5619), .B(n5618), .ZN(n5621)
         );
  INV_X1 U7042 ( .A(n5621), .ZN(n5622) );
  NAND2_X1 U7043 ( .A1(n5623), .A2(n5622), .ZN(n9280) );
  NAND2_X1 U7044 ( .A1(n9280), .A2(n4398), .ZN(n5624) );
  NAND2_X1 U7045 ( .A1(n5625), .A2(n5624), .ZN(n5626) );
  XNOR2_X1 U7046 ( .A(n5626), .B(n7160), .ZN(n5627) );
  AOI22_X1 U7047 ( .A1(n9407), .A2(n5096), .B1(n5640), .B2(n9280), .ZN(n8978)
         );
  INV_X1 U7048 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7667) );
  INV_X1 U7049 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7643) );
  MUX2_X1 U7050 ( .A(n7667), .B(n7643), .S(n5447), .Z(n5644) );
  XNOR2_X1 U7051 ( .A(n5644), .B(SI_24_), .ZN(n5643) );
  XNOR2_X1 U7052 ( .A(n5648), .B(n5643), .ZN(n7642) );
  NAND2_X1 U7053 ( .A1(n7642), .A2(n8389), .ZN(n5631) );
  OR2_X1 U7054 ( .A1(n8391), .A2(n7643), .ZN(n5630) );
  INV_X1 U7055 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n10069) );
  NAND2_X1 U7056 ( .A1(n5632), .A2(n10069), .ZN(n5633) );
  AND2_X1 U7057 ( .A1(n5657), .A2(n5633), .ZN(n9247) );
  NAND2_X1 U7058 ( .A1(n9247), .A2(n5758), .ZN(n5638) );
  INV_X1 U7059 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n10151) );
  NAND2_X1 U7060 ( .A1(n8289), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5635) );
  NAND2_X1 U7061 ( .A1(n8288), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5634) );
  OAI211_X1 U7062 ( .C1(n5689), .C2(n10151), .A(n5635), .B(n5634), .ZN(n5636)
         );
  INV_X1 U7063 ( .A(n5636), .ZN(n5637) );
  NAND2_X1 U7064 ( .A1(n5638), .A2(n5637), .ZN(n9259) );
  AOI22_X1 U7065 ( .A1(n9402), .A2(n6492), .B1(n5096), .B2(n9259), .ZN(n5639)
         );
  XNOR2_X1 U7066 ( .A(n5639), .B(n7160), .ZN(n5642) );
  AOI22_X1 U7067 ( .A1(n9402), .A2(n5096), .B1(n5640), .B2(n9259), .ZN(n5641)
         );
  XNOR2_X1 U7068 ( .A(n5642), .B(n5641), .ZN(n9011) );
  INV_X1 U7069 ( .A(n5643), .ZN(n5647) );
  INV_X1 U7070 ( .A(n5644), .ZN(n5645) );
  NAND2_X1 U7071 ( .A1(n5645), .A2(SI_24_), .ZN(n5646) );
  INV_X1 U7072 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n10075) );
  INV_X1 U7073 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7816) );
  MUX2_X1 U7074 ( .A(n10075), .B(n7816), .S(n5601), .Z(n5650) );
  INV_X1 U7075 ( .A(SI_25_), .ZN(n5649) );
  NAND2_X1 U7076 ( .A1(n5650), .A2(n5649), .ZN(n5674) );
  INV_X1 U7077 ( .A(n5650), .ZN(n5651) );
  NAND2_X1 U7078 ( .A1(n5651), .A2(SI_25_), .ZN(n5652) );
  NAND2_X1 U7079 ( .A1(n5674), .A2(n5652), .ZN(n5672) );
  OR2_X1 U7080 ( .A1(n8391), .A2(n7816), .ZN(n5653) );
  INV_X1 U7081 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n5656) );
  NAND2_X1 U7082 ( .A1(n5657), .A2(n5656), .ZN(n5658) );
  NAND2_X1 U7083 ( .A1(n5684), .A2(n5658), .ZN(n9225) );
  INV_X1 U7084 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n5661) );
  NAND2_X1 U7085 ( .A1(n8288), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5660) );
  NAND2_X1 U7086 ( .A1(n8289), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5659) );
  OAI211_X1 U7087 ( .C1(n5689), .C2(n5661), .A(n5660), .B(n5659), .ZN(n5662)
         );
  INV_X1 U7088 ( .A(n5662), .ZN(n5663) );
  AOI22_X1 U7089 ( .A1(n9395), .A2(n4398), .B1(n5640), .B2(n9216), .ZN(n5668)
         );
  NAND2_X1 U7090 ( .A1(n9395), .A2(n6492), .ZN(n5666) );
  NAND2_X1 U7091 ( .A1(n9216), .A2(n5096), .ZN(n5665) );
  NAND2_X1 U7092 ( .A1(n5666), .A2(n5665), .ZN(n5667) );
  XNOR2_X1 U7093 ( .A(n5667), .B(n7160), .ZN(n5670) );
  XOR2_X1 U7094 ( .A(n5668), .B(n5670), .Z(n9003) );
  INV_X1 U7095 ( .A(n5668), .ZN(n5669) );
  INV_X1 U7096 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7924) );
  INV_X1 U7097 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7927) );
  MUX2_X1 U7098 ( .A(n7924), .B(n7927), .S(n5447), .Z(n5676) );
  INV_X1 U7099 ( .A(SI_26_), .ZN(n5675) );
  NAND2_X1 U7100 ( .A1(n5676), .A2(n5675), .ZN(n5700) );
  INV_X1 U7101 ( .A(n5676), .ZN(n5677) );
  NAND2_X1 U7102 ( .A1(n5677), .A2(SI_26_), .ZN(n5678) );
  AND2_X1 U7103 ( .A1(n5700), .A2(n5678), .ZN(n5679) );
  NAND2_X1 U7104 ( .A1(n7922), .A2(n8389), .ZN(n5682) );
  OR2_X1 U7105 ( .A1(n8391), .A2(n7927), .ZN(n5681) );
  NAND2_X1 U7106 ( .A1(n9391), .A2(n6492), .ZN(n5694) );
  INV_X1 U7107 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n5683) );
  NAND2_X1 U7108 ( .A1(n5684), .A2(n5683), .ZN(n5685) );
  NAND2_X1 U7109 ( .A1(n5753), .A2(n5685), .ZN(n9207) );
  INV_X1 U7110 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n5688) );
  NAND2_X1 U7111 ( .A1(n8289), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5687) );
  NAND2_X1 U7112 ( .A1(n5154), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n5686) );
  OAI211_X1 U7113 ( .C1(n5689), .C2(n5688), .A(n5687), .B(n5686), .ZN(n5690)
         );
  INV_X1 U7114 ( .A(n5690), .ZN(n5691) );
  NAND2_X1 U7115 ( .A1(n9232), .A2(n5096), .ZN(n5693) );
  NAND2_X1 U7116 ( .A1(n5694), .A2(n5693), .ZN(n5695) );
  XNOR2_X1 U7117 ( .A(n5695), .B(n7160), .ZN(n5699) );
  NAND2_X1 U7118 ( .A1(n9391), .A2(n4398), .ZN(n5697) );
  NAND2_X1 U7119 ( .A1(n9232), .A2(n5640), .ZN(n5696) );
  NAND2_X1 U7120 ( .A1(n5697), .A2(n5696), .ZN(n5698) );
  NAND2_X1 U7121 ( .A1(n5699), .A2(n5698), .ZN(n9064) );
  INV_X1 U7122 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n7943) );
  INV_X1 U7123 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n7939) );
  MUX2_X1 U7124 ( .A(n7943), .B(n7939), .S(n5601), .Z(n5702) );
  INV_X1 U7125 ( .A(SI_27_), .ZN(n10041) );
  NAND2_X1 U7126 ( .A1(n5702), .A2(n10041), .ZN(n6144) );
  INV_X1 U7127 ( .A(n5702), .ZN(n5703) );
  NAND2_X1 U7128 ( .A1(n5703), .A2(SI_27_), .ZN(n5704) );
  AND2_X1 U7129 ( .A1(n6144), .A2(n5704), .ZN(n6143) );
  NAND2_X1 U7130 ( .A1(n7940), .A2(n8389), .ZN(n5706) );
  OR2_X1 U7131 ( .A1(n8391), .A2(n7939), .ZN(n5705) );
  NAND2_X1 U7132 ( .A1(n9385), .A2(n6492), .ZN(n5715) );
  XNOR2_X1 U7133 ( .A(n5753), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n9192) );
  NAND2_X1 U7134 ( .A1(n9192), .A2(n5758), .ZN(n5713) );
  INV_X1 U7135 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n5710) );
  NAND2_X1 U7136 ( .A1(n8287), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n5708) );
  NAND2_X1 U7137 ( .A1(n8289), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5707) );
  OAI211_X1 U7138 ( .C1(n5710), .C2(n5709), .A(n5708), .B(n5707), .ZN(n5711)
         );
  INV_X1 U7139 ( .A(n5711), .ZN(n5712) );
  NAND2_X1 U7140 ( .A1(n5713), .A2(n5712), .ZN(n9217) );
  NAND2_X1 U7141 ( .A1(n9217), .A2(n4398), .ZN(n5714) );
  NAND2_X1 U7142 ( .A1(n5715), .A2(n5714), .ZN(n5716) );
  XNOR2_X1 U7143 ( .A(n5716), .B(n6490), .ZN(n5719) );
  AND2_X1 U7144 ( .A1(n9217), .A2(n5640), .ZN(n5717) );
  AOI21_X1 U7145 ( .B1(n9385), .B2(n4398), .A(n5717), .ZN(n5718) );
  NAND2_X1 U7146 ( .A1(n5719), .A2(n5718), .ZN(n6506) );
  OAI21_X1 U7147 ( .B1(n5719), .B2(n5718), .A(n6506), .ZN(n5721) );
  NAND2_X1 U7148 ( .A1(n7814), .A2(P1_B_REG_SCAN_IN), .ZN(n5723) );
  INV_X1 U7149 ( .A(n7644), .ZN(n5722) );
  MUX2_X1 U7150 ( .A(n5723), .B(P1_B_REG_SCAN_IN), .S(n5722), .Z(n5724) );
  AND2_X1 U7151 ( .A1(n5724), .A2(n5725), .ZN(n9729) );
  INV_X1 U7152 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n6624) );
  INV_X1 U7153 ( .A(n5725), .ZN(n7925) );
  AND2_X1 U7154 ( .A1(n7925), .A2(n7644), .ZN(n5726) );
  AOI21_X1 U7155 ( .B1(n9729), .B2(n6624), .A(n5726), .ZN(n6829) );
  NOR4_X1 U7156 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_17__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_23__SCAN_IN), .ZN(n5730) );
  NOR4_X1 U7157 ( .A1(P1_D_REG_13__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_11__SCAN_IN), .A4(P1_D_REG_14__SCAN_IN), .ZN(n5729) );
  INV_X1 U7158 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n10158) );
  INV_X1 U7159 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n10196) );
  INV_X1 U7160 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n10040) );
  INV_X1 U7161 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n10092) );
  NAND4_X1 U7162 ( .A1(n10158), .A2(n10196), .A3(n10040), .A4(n10092), .ZN(
        n5727) );
  NOR2_X1 U7163 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n5727), .ZN(n9959) );
  NOR4_X1 U7164 ( .A1(P1_D_REG_27__SCAN_IN), .A2(P1_D_REG_24__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n5728) );
  NAND4_X1 U7165 ( .A1(n5730), .A2(n5729), .A3(n9959), .A4(n5728), .ZN(n5735)
         );
  NOR4_X1 U7166 ( .A1(P1_D_REG_28__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_3__SCAN_IN), .A4(P1_D_REG_19__SCAN_IN), .ZN(n5733) );
  NOR4_X1 U7167 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_8__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n5732) );
  NOR4_X1 U7168 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_25__SCAN_IN), .A3(
        P1_D_REG_6__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5731) );
  INV_X1 U7169 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n9734) );
  NAND4_X1 U7170 ( .A1(n5733), .A2(n5732), .A3(n5731), .A4(n9734), .ZN(n5734)
         );
  OAI21_X1 U7171 ( .B1(n5735), .B2(n5734), .A(n9729), .ZN(n6830) );
  NAND2_X1 U7172 ( .A1(n6829), .A2(n6830), .ZN(n6769) );
  INV_X1 U7173 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n9754) );
  NAND2_X1 U7174 ( .A1(n9729), .A2(n9754), .ZN(n5737) );
  NAND2_X1 U7175 ( .A1(n7925), .A2(n7814), .ZN(n5736) );
  NAND2_X1 U7176 ( .A1(n5737), .A2(n5736), .ZN(n7038) );
  OR2_X1 U7177 ( .A1(n6769), .A2(n7038), .ZN(n5764) );
  INV_X1 U7178 ( .A(n5764), .ZN(n5746) );
  NAND2_X1 U7179 ( .A1(n5738), .A2(n8514), .ZN(n8508) );
  NAND2_X1 U7180 ( .A1(n4437), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5741) );
  XNOR2_X1 U7181 ( .A(n5741), .B(n5740), .ZN(n7447) );
  AND2_X1 U7182 ( .A1(n7447), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5742) );
  AND2_X1 U7183 ( .A1(n6513), .A2(n5742), .ZN(n9755) );
  AND2_X1 U7184 ( .A1(n8508), .A2(n9755), .ZN(n5745) );
  NAND2_X1 U7185 ( .A1(n5743), .A2(n5744), .ZN(n7044) );
  NAND3_X1 U7186 ( .A1(n5746), .A2(n5745), .A3(n9787), .ZN(n9075) );
  OAI21_X1 U7187 ( .B1(n6509), .B2(n5748), .A(n5747), .ZN(n5771) );
  OR2_X1 U7188 ( .A1(n7044), .A2(n8543), .ZN(n9706) );
  INV_X1 U7189 ( .A(n9755), .ZN(n9730) );
  OR2_X1 U7190 ( .A1(n9706), .A2(n9730), .ZN(n5763) );
  NAND2_X1 U7191 ( .A1(n5743), .A2(n5505), .ZN(n8406) );
  OR2_X1 U7192 ( .A1(n8406), .A2(n6898), .ZN(n6886) );
  NAND2_X1 U7193 ( .A1(n9755), .A2(n5744), .ZN(n5749) );
  OAI21_X1 U7194 ( .B1(n5763), .B2(n5764), .A(n9708), .ZN(n9073) );
  NAND2_X1 U7195 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n5750) );
  INV_X1 U7196 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n5752) );
  INV_X1 U7197 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n5751) );
  OAI21_X1 U7198 ( .B1(n5753), .B2(n5752), .A(n5751), .ZN(n5754) );
  INV_X1 U7199 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n10038) );
  NAND2_X1 U7200 ( .A1(n8288), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n5756) );
  NAND2_X1 U7201 ( .A1(n8287), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n5755) );
  OAI211_X1 U7202 ( .C1(n5063), .C2(n10038), .A(n5756), .B(n5755), .ZN(n5757)
         );
  AOI21_X1 U7203 ( .B1(n9180), .B2(n5758), .A(n5757), .ZN(n9157) );
  OR2_X1 U7204 ( .A1(n6907), .A2(n4987), .ZN(n7161) );
  OR2_X1 U7205 ( .A1(n7161), .A2(n9730), .ZN(n8548) );
  NOR2_X1 U7206 ( .A1(n8548), .A2(n5764), .ZN(n5760) );
  NAND2_X1 U7207 ( .A1(n5760), .A2(n5759), .ZN(n9014) );
  INV_X1 U7208 ( .A(n5759), .ZN(n6764) );
  AND2_X1 U7209 ( .A1(n5760), .A2(n6764), .ZN(n9068) );
  AOI22_X1 U7210 ( .A1(n9232), .A2(n9068), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3084), .ZN(n5768) );
  OR2_X1 U7211 ( .A1(n8508), .A2(n7043), .ZN(n6768) );
  AND3_X1 U7212 ( .A1(n6768), .A2(n6513), .A3(n7447), .ZN(n5761) );
  NAND2_X1 U7213 ( .A1(n5764), .A2(n9787), .ZN(n6778) );
  NAND2_X1 U7214 ( .A1(n5761), .A2(n6778), .ZN(n5762) );
  NAND2_X1 U7215 ( .A1(n5762), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5766) );
  INV_X1 U7216 ( .A(n5763), .ZN(n5765) );
  NAND2_X1 U7217 ( .A1(n5765), .A2(n5764), .ZN(n6780) );
  NAND2_X1 U7218 ( .A1(n5766), .A2(n6780), .ZN(n9049) );
  NAND2_X1 U7219 ( .A1(n9192), .A2(n9049), .ZN(n5767) );
  OAI211_X1 U7220 ( .C1(n9157), .C2(n9014), .A(n5768), .B(n5767), .ZN(n5769)
         );
  AOI21_X1 U7221 ( .B1(n9385), .B2(n9073), .A(n5769), .ZN(n5770) );
  NAND2_X1 U7222 ( .A1(n5771), .A2(n5770), .ZN(P1_U3212) );
  INV_X1 U7223 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5772) );
  NOR2_X1 U7224 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n5774) );
  NOR2_X1 U7225 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n5773) );
  INV_X1 U7226 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n6211) );
  INV_X1 U7227 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5780) );
  NAND2_X1 U7228 ( .A1(n6211), .A2(n5780), .ZN(n6188) );
  INV_X1 U7229 ( .A(n6188), .ZN(n5782) );
  NOR2_X1 U7230 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .ZN(
        n5781) );
  NAND4_X1 U7231 ( .A1(n5782), .A2(n5781), .A3(n6405), .A4(n6216), .ZN(n5784)
         );
  INV_X1 U7232 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n6046) );
  NAND4_X1 U7233 ( .A1(n6046), .A2(n6406), .A3(n6035), .A4(n6014), .ZN(n5783)
         );
  NAND2_X1 U7234 ( .A1(n5789), .A2(n5790), .ZN(n8967) );
  INV_X1 U7235 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5788) );
  NAND2_X1 U7236 ( .A1(n6192), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5805) );
  NAND2_X1 U7237 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_REG3_REG_9__SCAN_IN), 
        .ZN(n5796) );
  INV_X1 U7238 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n5967) );
  INV_X1 U7239 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5990) );
  INV_X1 U7240 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n10059) );
  NAND2_X1 U7241 ( .A1(n5993), .A2(n10059), .ZN(n5799) );
  NAND2_X1 U7242 ( .A1(n6006), .A2(n5799), .ZN(n7837) );
  OR2_X1 U7243 ( .A1(n6152), .A2(n7837), .ZN(n5804) );
  INV_X2 U7244 ( .A(n6030), .ZN(n5890) );
  INV_X1 U7245 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n5800) );
  OR2_X1 U7246 ( .A1(n5890), .A2(n5800), .ZN(n5803) );
  NAND2_X2 U7247 ( .A1(n5801), .A2(n8078), .ZN(n5875) );
  INV_X1 U7248 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n7683) );
  OR2_X1 U7249 ( .A1(n5875), .A2(n7683), .ZN(n5802) );
  NAND4_X1 U7250 ( .A1(n5805), .A2(n5804), .A3(n5803), .A4(n5802), .ZN(n8642)
         );
  INV_X1 U7251 ( .A(n8642), .ZN(n7843) );
  MUX2_X1 U7252 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5806), .S(
        P2_IR_REG_27__SCAN_IN), .Z(n5807) );
  INV_X1 U7253 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5809) );
  NAND2_X1 U7254 ( .A1(n6656), .A2(n6169), .ZN(n5824) );
  NOR2_X1 U7255 ( .A1(n5811), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n5899) );
  NAND2_X1 U7256 ( .A1(n5899), .A2(n5812), .ZN(n5913) );
  INV_X1 U7257 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5814) );
  NAND3_X1 U7258 ( .A1(n5949), .A2(n5813), .A3(n5814), .ZN(n5815) );
  NOR2_X1 U7259 ( .A1(n5934), .A2(n5815), .ZN(n5974) );
  NAND2_X1 U7260 ( .A1(n5974), .A2(n5816), .ZN(n5817) );
  NAND2_X1 U7261 ( .A1(n5817), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5987) );
  NAND2_X1 U7262 ( .A1(n5987), .A2(n5818), .ZN(n5819) );
  NAND2_X1 U7263 ( .A1(n5819), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5821) );
  NAND2_X1 U7264 ( .A1(n5821), .A2(n5820), .ZN(n6000) );
  OR2_X1 U7265 ( .A1(n5821), .A2(n5820), .ZN(n5822) );
  AND2_X1 U7266 ( .A1(n6000), .A2(n5822), .ZN(n7872) );
  AOI22_X1 U7267 ( .A1(n7872), .A2(n6049), .B1(n6206), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n5823) );
  INV_X1 U7268 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n5825) );
  OR2_X1 U7269 ( .A1(n6152), .A2(n5825), .ZN(n5830) );
  INV_X1 U7270 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n5826) );
  INV_X1 U7271 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n5827) );
  OR2_X1 U7272 ( .A1(n5888), .A2(n5827), .ZN(n5828) );
  NAND4_X2 U7273 ( .A1(n5831), .A2(n5830), .A3(n5829), .A4(n5828), .ZN(n8655)
         );
  INV_X1 U7274 ( .A(n4392), .ZN(n5912) );
  INV_X1 U7275 ( .A(n6608), .ZN(n5832) );
  NAND2_X1 U7276 ( .A1(n5912), .A2(n5832), .ZN(n5837) );
  NAND2_X1 U7277 ( .A1(n6050), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n5836) );
  OR2_X1 U7278 ( .A1(n5833), .A2(n5788), .ZN(n5834) );
  XNOR2_X2 U7279 ( .A(n5834), .B(P2_IR_REG_2__SCAN_IN), .ZN(n6556) );
  NAND2_X1 U7280 ( .A1(n6049), .A2(n6556), .ZN(n5835) );
  AND3_X2 U7281 ( .A1(n5837), .A2(n5836), .A3(n5835), .ZN(n9858) );
  OR2_X1 U7282 ( .A1(n8655), .A2(n9858), .ZN(n6244) );
  NAND2_X1 U7283 ( .A1(n8655), .A2(n9858), .ZN(n6246) );
  NAND2_X1 U7284 ( .A1(n6244), .A2(n6246), .ZN(n7307) );
  INV_X1 U7285 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n7337) );
  OR2_X1 U7286 ( .A1(n6152), .A2(n7337), .ZN(n5844) );
  INV_X1 U7287 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n5838) );
  OR2_X1 U7288 ( .A1(n5888), .A2(n5838), .ZN(n5842) );
  INV_X1 U7289 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n5839) );
  OR2_X1 U7290 ( .A1(n5875), .A2(n5839), .ZN(n5841) );
  NAND2_X1 U7291 ( .A1(n6030), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5840) );
  AND3_X1 U7292 ( .A1(n5842), .A2(n5841), .A3(n5840), .ZN(n5843) );
  INV_X1 U7293 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n9816) );
  NAND2_X1 U7294 ( .A1(n6607), .A2(SI_0_), .ZN(n5846) );
  INV_X1 U7295 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5845) );
  XNOR2_X1 U7296 ( .A(n5846), .B(n5845), .ZN(n8975) );
  MUX2_X1 U7297 ( .A(n9816), .B(n8975), .S(n6565), .Z(n7197) );
  INV_X1 U7298 ( .A(n5875), .ZN(n5847) );
  NAND2_X1 U7299 ( .A1(n5847), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5853) );
  NAND2_X1 U7300 ( .A1(n5848), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n5852) );
  INV_X1 U7301 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n5849) );
  OR2_X1 U7302 ( .A1(n5888), .A2(n5849), .ZN(n5851) );
  INV_X1 U7303 ( .A(n6615), .ZN(n5854) );
  NAND2_X1 U7304 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5855) );
  INV_X1 U7305 ( .A(n5833), .ZN(n5856) );
  INV_X1 U7306 ( .A(n6951), .ZN(n5859) );
  NAND2_X1 U7307 ( .A1(n5860), .A2(n5859), .ZN(n6368) );
  NAND2_X1 U7308 ( .A1(n6938), .A2(n6368), .ZN(n6237) );
  NAND2_X1 U7309 ( .A1(n7310), .A2(n7309), .ZN(n7308) );
  NAND2_X1 U7310 ( .A1(n7308), .A2(n6244), .ZN(n7497) );
  INV_X1 U7311 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n5861) );
  INV_X1 U7312 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n5862) );
  INV_X1 U7313 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n5863) );
  OR2_X1 U7314 ( .A1(n5888), .A2(n5863), .ZN(n5865) );
  OR2_X1 U7315 ( .A1(n6152), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5864) );
  NAND2_X1 U7316 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n4397), .ZN(n5868) );
  XNOR2_X1 U7317 ( .A(n5868), .B(P2_IR_REG_3__SCAN_IN), .ZN(n6557) );
  NAND2_X1 U7318 ( .A1(n6049), .A2(n6557), .ZN(n5869) );
  NAND2_X1 U7319 ( .A1(n7497), .A2(n7496), .ZN(n7495) );
  INV_X1 U7320 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n5871) );
  INV_X1 U7321 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n5872) );
  OR2_X1 U7322 ( .A1(n5890), .A2(n5872), .ZN(n5878) );
  INV_X1 U7323 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5873) );
  NAND2_X1 U7324 ( .A1(n5891), .A2(n5873), .ZN(n5874) );
  NAND2_X1 U7325 ( .A1(n5905), .A2(n5874), .ZN(n9824) );
  OR2_X1 U7326 ( .A1(n6152), .A2(n9824), .ZN(n5877) );
  INV_X1 U7327 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6560) );
  OR2_X1 U7328 ( .A1(n5875), .A2(n6560), .ZN(n5876) );
  OR2_X1 U7329 ( .A1(n6620), .A2(n4392), .ZN(n5882) );
  NAND2_X1 U7330 ( .A1(n5811), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5880) );
  XNOR2_X1 U7331 ( .A(n5880), .B(P2_IR_REG_5__SCAN_IN), .ZN(n6586) );
  AOI22_X1 U7332 ( .A1(n6050), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n6049), .B2(
        n6586), .ZN(n5881) );
  NAND2_X1 U7333 ( .A1(n5882), .A2(n5881), .ZN(n7101) );
  NAND2_X1 U7334 ( .A1(n7211), .A2(n7101), .ZN(n6235) );
  NAND2_X1 U7335 ( .A1(n5883), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5884) );
  XNOR2_X1 U7336 ( .A(n5884), .B(P2_IR_REG_4__SCAN_IN), .ZN(n6559) );
  AOI22_X1 U7337 ( .A1(n6050), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n6049), .B2(
        n6559), .ZN(n5886) );
  OR2_X1 U7338 ( .A1(n6613), .A2(n4392), .ZN(n5885) );
  INV_X1 U7339 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n5887) );
  INV_X1 U7340 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n5889) );
  OR2_X1 U7341 ( .A1(n5890), .A2(n5889), .ZN(n5895) );
  OAI21_X1 U7342 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(P2_REG3_REG_4__SCAN_IN), 
        .A(n5891), .ZN(n7363) );
  OR2_X1 U7343 ( .A1(n6152), .A2(n7363), .ZN(n5894) );
  INV_X1 U7344 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n5892) );
  OR2_X1 U7345 ( .A1(n5875), .A2(n5892), .ZN(n5893) );
  OR2_X1 U7346 ( .A1(n9869), .A2(n8653), .ZN(n6234) );
  NAND2_X1 U7347 ( .A1(n6234), .A2(n7093), .ZN(n7356) );
  NAND3_X1 U7348 ( .A1(n7495), .A2(n6235), .A3(n7091), .ZN(n7208) );
  INV_X1 U7349 ( .A(n6235), .ZN(n5898) );
  INV_X1 U7350 ( .A(n7211), .ZN(n8652) );
  INV_X1 U7351 ( .A(n7101), .ZN(n9823) );
  OR2_X1 U7352 ( .A1(n5898), .A2(n7092), .ZN(n7207) );
  NAND2_X1 U7353 ( .A1(n6625), .A2(n5912), .ZN(n5902) );
  OR2_X1 U7354 ( .A1(n5899), .A2(n5788), .ZN(n5900) );
  XNOR2_X1 U7355 ( .A(n5900), .B(P2_IR_REG_6__SCAN_IN), .ZN(n6807) );
  AOI22_X1 U7356 ( .A1(n6050), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n6049), .B2(
        n6807), .ZN(n5901) );
  NAND2_X1 U7357 ( .A1(n5902), .A2(n5901), .ZN(n7221) );
  INV_X1 U7358 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n5903) );
  INV_X1 U7359 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7215) );
  OR2_X1 U7360 ( .A1(n5890), .A2(n7215), .ZN(n5909) );
  INV_X1 U7361 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n5904) );
  NAND2_X1 U7362 ( .A1(n5905), .A2(n5904), .ZN(n5906) );
  NAND2_X1 U7363 ( .A1(n5918), .A2(n5906), .ZN(n7214) );
  OR2_X1 U7364 ( .A1(n6152), .A2(n7214), .ZN(n5908) );
  INV_X1 U7365 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6590) );
  OR2_X1 U7366 ( .A1(n5875), .A2(n6590), .ZN(n5907) );
  NAND4_X1 U7367 ( .A1(n5910), .A2(n5909), .A3(n5908), .A4(n5907), .ZN(n8651)
         );
  NAND2_X1 U7368 ( .A1(n7208), .A2(n5911), .ZN(n7209) );
  INV_X1 U7369 ( .A(n8651), .ZN(n7029) );
  NAND2_X1 U7370 ( .A1(n7221), .A2(n7029), .ZN(n6259) );
  NAND2_X1 U7371 ( .A1(n6629), .A2(n5912), .ZN(n5916) );
  NAND2_X1 U7372 ( .A1(n5913), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5914) );
  XNOR2_X1 U7373 ( .A(n5914), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6821) );
  AOI22_X1 U7374 ( .A1(n6050), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6049), .B2(
        n6821), .ZN(n5915) );
  NAND2_X1 U7375 ( .A1(n5916), .A2(n5915), .ZN(n7129) );
  NAND2_X1 U7376 ( .A1(n6192), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5924) );
  INV_X1 U7377 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n5917) );
  OR2_X1 U7378 ( .A1(n5890), .A2(n5917), .ZN(n5923) );
  INV_X1 U7379 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n7019) );
  NAND2_X1 U7380 ( .A1(n5918), .A2(n7019), .ZN(n5919) );
  NAND2_X1 U7381 ( .A1(n5941), .A2(n5919), .ZN(n7461) );
  OR2_X1 U7382 ( .A1(n6152), .A2(n7461), .ZN(n5922) );
  INV_X1 U7383 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n5920) );
  OR2_X1 U7384 ( .A1(n5875), .A2(n5920), .ZN(n5921) );
  OR2_X1 U7385 ( .A1(n7129), .A2(n7554), .ZN(n6260) );
  NAND2_X1 U7386 ( .A1(n7129), .A2(n7554), .ZN(n6261) );
  NAND2_X1 U7387 ( .A1(n6633), .A2(n6169), .ZN(n5928) );
  NAND2_X1 U7388 ( .A1(n5925), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5926) );
  XNOR2_X1 U7389 ( .A(n5926), .B(P2_IR_REG_8__SCAN_IN), .ZN(n6864) );
  AOI22_X1 U7390 ( .A1(n6050), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6049), .B2(
        n6864), .ZN(n5927) );
  NAND2_X1 U7391 ( .A1(n5928), .A2(n5927), .ZN(n9881) );
  NAND2_X1 U7392 ( .A1(n6192), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5933) );
  INV_X1 U7393 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n6822) );
  OR2_X1 U7394 ( .A1(n5890), .A2(n6822), .ZN(n5932) );
  INV_X1 U7395 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n5940) );
  XNOR2_X1 U7396 ( .A(n5941), .B(n5940), .ZN(n7562) );
  OR2_X1 U7397 ( .A1(n6152), .A2(n7562), .ZN(n5931) );
  INV_X1 U7398 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n5929) );
  OR2_X1 U7399 ( .A1(n5875), .A2(n5929), .ZN(n5930) );
  OR2_X1 U7400 ( .A1(n9881), .A2(n7474), .ZN(n6264) );
  NAND2_X1 U7401 ( .A1(n9881), .A2(n7474), .ZN(n7477) );
  NAND2_X1 U7402 ( .A1(n6636), .A2(n6169), .ZN(n5936) );
  NAND2_X1 U7403 ( .A1(n5934), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5950) );
  XNOR2_X1 U7404 ( .A(n5950), .B(P2_IR_REG_9__SCAN_IN), .ZN(n6921) );
  AOI22_X1 U7405 ( .A1(n6050), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6049), .B2(
        n6921), .ZN(n5935) );
  NAND2_X1 U7406 ( .A1(n5937), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5946) );
  INV_X1 U7407 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n5938) );
  OR2_X1 U7408 ( .A1(n5888), .A2(n5938), .ZN(n5945) );
  INV_X1 U7409 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7486) );
  OR2_X1 U7410 ( .A1(n5890), .A2(n7486), .ZN(n5944) );
  INV_X1 U7411 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5939) );
  OAI21_X1 U7412 ( .B1(n5941), .B2(n5940), .A(n5939), .ZN(n5942) );
  NAND2_X1 U7413 ( .A1(n5942), .A2(n5957), .ZN(n7485) );
  OR2_X1 U7414 ( .A1(n6152), .A2(n7485), .ZN(n5943) );
  OR2_X1 U7415 ( .A1(n7646), .A2(n7553), .ZN(n6267) );
  NAND2_X1 U7416 ( .A1(n7646), .A2(n7553), .ZN(n6266) );
  AND2_X1 U7417 ( .A1(n7552), .A2(n7472), .ZN(n5947) );
  OR2_X1 U7418 ( .A1(n7478), .A2(n7477), .ZN(n7475) );
  NAND2_X1 U7419 ( .A1(n6648), .A2(n6169), .ZN(n5956) );
  NAND2_X1 U7420 ( .A1(n5950), .A2(n5949), .ZN(n5951) );
  NAND2_X1 U7421 ( .A1(n5951), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5953) );
  INV_X1 U7422 ( .A(n5953), .ZN(n5952) );
  NAND2_X1 U7423 ( .A1(n5952), .A2(P2_IR_REG_10__SCAN_IN), .ZN(n5954) );
  NAND2_X1 U7424 ( .A1(n5953), .A2(n5813), .ZN(n5963) );
  AND2_X1 U7425 ( .A1(n5954), .A2(n5963), .ZN(n7113) );
  AOI22_X1 U7426 ( .A1(n6050), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n7113), .B2(
        n6049), .ZN(n5955) );
  NAND2_X1 U7427 ( .A1(n6192), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5962) );
  INV_X1 U7428 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7617) );
  OR2_X1 U7429 ( .A1(n5890), .A2(n7617), .ZN(n5961) );
  INV_X1 U7430 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n10223) );
  NAND2_X1 U7431 ( .A1(n5957), .A2(n10223), .ZN(n5958) );
  NAND2_X1 U7432 ( .A1(n5968), .A2(n5958), .ZN(n7616) );
  OR2_X1 U7433 ( .A1(n6152), .A2(n7616), .ZN(n5960) );
  INV_X1 U7434 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n6924) );
  OR2_X1 U7435 ( .A1(n5875), .A2(n6924), .ZN(n5959) );
  OR2_X1 U7436 ( .A1(n9891), .A2(n7473), .ZN(n6270) );
  NAND2_X1 U7437 ( .A1(n9891), .A2(n7473), .ZN(n6275) );
  NAND2_X1 U7438 ( .A1(n6270), .A2(n6275), .ZN(n6432) );
  NAND2_X1 U7439 ( .A1(n6651), .A2(n6169), .ZN(n5966) );
  NAND2_X1 U7440 ( .A1(n5963), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5964) );
  XNOR2_X1 U7441 ( .A(n5964), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7454) );
  AOI22_X1 U7442 ( .A1(n7454), .A2(n6049), .B1(n6206), .B2(
        P1_DATAO_REG_11__SCAN_IN), .ZN(n5965) );
  NAND2_X1 U7443 ( .A1(n6192), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5973) );
  INV_X1 U7444 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7633) );
  OR2_X1 U7445 ( .A1(n5890), .A2(n7633), .ZN(n5972) );
  NAND2_X1 U7446 ( .A1(n5968), .A2(n5967), .ZN(n5969) );
  NAND2_X1 U7447 ( .A1(n5980), .A2(n5969), .ZN(n7632) );
  OR2_X1 U7448 ( .A1(n6152), .A2(n7632), .ZN(n5971) );
  INV_X1 U7449 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n7111) );
  OR2_X1 U7450 ( .A1(n5875), .A2(n7111), .ZN(n5970) );
  NAND2_X1 U7451 ( .A1(n7670), .A2(n7707), .ZN(n6366) );
  NAND2_X1 U7452 ( .A1(n7624), .A2(n6366), .ZN(n7568) );
  NAND2_X1 U7453 ( .A1(n6688), .A2(n6169), .ZN(n5977) );
  OR2_X1 U7454 ( .A1(n5974), .A2(n5788), .ZN(n5975) );
  XNOR2_X1 U7455 ( .A(n5975), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7518) );
  AOI22_X1 U7456 ( .A1(n6050), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n7518), .B2(
        n6049), .ZN(n5976) );
  NAND2_X1 U7457 ( .A1(n6192), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5985) );
  INV_X1 U7458 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n5978) );
  OR2_X1 U7459 ( .A1(n5890), .A2(n5978), .ZN(n5984) );
  INV_X1 U7460 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n5979) );
  NAND2_X1 U7461 ( .A1(n5980), .A2(n5979), .ZN(n5981) );
  NAND2_X1 U7462 ( .A1(n5991), .A2(n5981), .ZN(n7574) );
  OR2_X1 U7463 ( .A1(n6152), .A2(n7574), .ZN(n5983) );
  INV_X1 U7464 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7521) );
  OR2_X1 U7465 ( .A1(n5875), .A2(n7521), .ZN(n5982) );
  OR2_X1 U7466 ( .A1(n7700), .A2(n7760), .ZN(n6365) );
  OR2_X1 U7467 ( .A1(n7670), .A2(n7707), .ZN(n7567) );
  AND2_X1 U7468 ( .A1(n6365), .A2(n7567), .ZN(n6278) );
  NAND2_X1 U7469 ( .A1(n7568), .A2(n6278), .ZN(n5986) );
  NAND2_X1 U7470 ( .A1(n7700), .A2(n7760), .ZN(n6364) );
  NAND2_X1 U7471 ( .A1(n5986), .A2(n6364), .ZN(n7743) );
  NAND2_X1 U7472 ( .A1(n6653), .A2(n6169), .ZN(n5989) );
  XNOR2_X1 U7473 ( .A(n5987), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7684) );
  AOI22_X1 U7474 ( .A1(n7684), .A2(n6049), .B1(n6206), .B2(
        P1_DATAO_REG_13__SCAN_IN), .ZN(n5988) );
  NAND2_X1 U7475 ( .A1(n6192), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5998) );
  INV_X1 U7476 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n7748) );
  OR2_X1 U7477 ( .A1(n5890), .A2(n7748), .ZN(n5997) );
  NAND2_X1 U7478 ( .A1(n5991), .A2(n5990), .ZN(n5992) );
  NAND2_X1 U7479 ( .A1(n5993), .A2(n5992), .ZN(n7759) );
  OR2_X1 U7480 ( .A1(n6152), .A2(n7759), .ZN(n5996) );
  INV_X1 U7481 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n5994) );
  OR2_X1 U7482 ( .A1(n5875), .A2(n5994), .ZN(n5995) );
  OR2_X1 U7483 ( .A1(n7763), .A2(n8643), .ZN(n6283) );
  NAND2_X1 U7484 ( .A1(n7763), .A2(n8643), .ZN(n5999) );
  INV_X1 U7485 ( .A(n5999), .ZN(n6285) );
  XNOR2_X1 U7486 ( .A(n9528), .B(n8642), .ZN(n7804) );
  NAND2_X1 U7487 ( .A1(n6757), .A2(n6169), .ZN(n6003) );
  NAND2_X1 U7488 ( .A1(n6000), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6001) );
  XNOR2_X1 U7489 ( .A(n6001), .B(P2_IR_REG_15__SCAN_IN), .ZN(n7874) );
  AOI22_X1 U7490 ( .A1(n7874), .A2(n6049), .B1(n6206), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n6002) );
  NAND2_X1 U7491 ( .A1(n6192), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n6012) );
  INV_X1 U7492 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n7851) );
  OR2_X1 U7493 ( .A1(n5890), .A2(n7851), .ZN(n6011) );
  INV_X1 U7494 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n6005) );
  NAND2_X1 U7495 ( .A1(n6006), .A2(n6005), .ZN(n6007) );
  NAND2_X1 U7496 ( .A1(n6020), .A2(n6007), .ZN(n8042) );
  OR2_X1 U7497 ( .A1(n6152), .A2(n8042), .ZN(n6010) );
  INV_X1 U7498 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n6008) );
  OR2_X1 U7499 ( .A1(n5875), .A2(n6008), .ZN(n6009) );
  NOR2_X1 U7500 ( .A1(n9521), .A2(n8120), .ZN(n6226) );
  NAND2_X1 U7501 ( .A1(n9521), .A2(n8120), .ZN(n6227) );
  NAND2_X1 U7502 ( .A1(n6761), .A2(n6169), .ZN(n6017) );
  NOR2_X1 U7503 ( .A1(n4366), .A2(n5788), .ZN(n6013) );
  MUX2_X1 U7504 ( .A(n5788), .B(n6013), .S(P2_IR_REG_16__SCAN_IN), .Z(n6015)
         );
  OR2_X1 U7505 ( .A1(n6015), .A2(n6036), .ZN(n8221) );
  INV_X1 U7506 ( .A(n8221), .ZN(n8227) );
  AOI22_X1 U7507 ( .A1(n6050), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6049), .B2(
        n8227), .ZN(n6016) );
  INV_X1 U7508 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n7952) );
  NAND2_X1 U7509 ( .A1(n6192), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n6018) );
  OAI21_X1 U7510 ( .B1(n5890), .B2(n7952), .A(n6018), .ZN(n6024) );
  INV_X1 U7511 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n10197) );
  NAND2_X1 U7512 ( .A1(n6020), .A2(n10197), .ZN(n6021) );
  NAND2_X1 U7513 ( .A1(n6028), .A2(n6021), .ZN(n8119) );
  NOR2_X1 U7514 ( .A1(n8119), .A2(n6152), .ZN(n6023) );
  INV_X1 U7515 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n10210) );
  NOR2_X1 U7516 ( .A1(n5875), .A2(n10210), .ZN(n6022) );
  INV_X1 U7517 ( .A(n8640), .ZN(n8073) );
  AND2_X1 U7518 ( .A1(n8111), .A2(n8073), .ZN(n6224) );
  OR2_X1 U7519 ( .A1(n8111), .A2(n8073), .ZN(n6293) );
  NAND2_X1 U7520 ( .A1(n6797), .A2(n6169), .ZN(n6027) );
  OR2_X1 U7521 ( .A1(n6036), .A2(n5788), .ZN(n6025) );
  XNOR2_X1 U7522 ( .A(n6025), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8229) );
  AOI22_X1 U7523 ( .A1(n6050), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6049), .B2(
        n8229), .ZN(n6026) );
  INV_X1 U7524 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8071) );
  NAND2_X1 U7525 ( .A1(n6028), .A2(n8071), .ZN(n6029) );
  AND2_X1 U7526 ( .A1(n6041), .A2(n6029), .ZN(n8070) );
  NAND2_X1 U7527 ( .A1(n8070), .A2(n5848), .ZN(n6033) );
  AOI22_X1 U7528 ( .A1(n6192), .A2(P2_REG0_REG_17__SCAN_IN), .B1(n6030), .B2(
        P2_REG2_REG_17__SCAN_IN), .ZN(n6032) );
  NAND2_X1 U7529 ( .A1(n5937), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n6031) );
  OR2_X1 U7530 ( .A1(n8930), .A2(n8132), .ZN(n6034) );
  NAND2_X1 U7531 ( .A1(n8930), .A2(n8132), .ZN(n6298) );
  INV_X1 U7532 ( .A(n6034), .ZN(n6301) );
  AOI21_X1 U7533 ( .B1(n8026), .B2(n6296), .A(n6301), .ZN(n8837) );
  NAND2_X1 U7534 ( .A1(n6872), .A2(n6169), .ZN(n6038) );
  XNOR2_X1 U7535 ( .A(n6047), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8230) );
  AOI22_X1 U7536 ( .A1(n6050), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6049), .B2(
        n8230), .ZN(n6037) );
  INV_X1 U7537 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n6040) );
  NAND2_X1 U7538 ( .A1(n6041), .A2(n6040), .ZN(n6042) );
  NAND2_X1 U7539 ( .A1(n6053), .A2(n6042), .ZN(n8847) );
  OR2_X1 U7540 ( .A1(n8847), .A2(n6152), .ZN(n6045) );
  AOI22_X1 U7541 ( .A1(n6192), .A2(P2_REG0_REG_18__SCAN_IN), .B1(n6030), .B2(
        P2_REG2_REG_18__SCAN_IN), .ZN(n6044) );
  INV_X1 U7542 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8220) );
  OR2_X1 U7543 ( .A1(n5875), .A2(n8220), .ZN(n6043) );
  AND2_X1 U7544 ( .A1(n8923), .A2(n8179), .ZN(n6297) );
  OR2_X1 U7545 ( .A1(n8923), .A2(n8179), .ZN(n6363) );
  NAND2_X1 U7546 ( .A1(n6987), .A2(n6169), .ZN(n6052) );
  NAND2_X1 U7547 ( .A1(n6047), .A2(n6046), .ZN(n6048) );
  AOI22_X1 U7548 ( .A1(n6050), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n6049), .B2(
        n8734), .ZN(n6051) );
  INV_X1 U7549 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n8178) );
  NAND2_X1 U7550 ( .A1(n6053), .A2(n8178), .ZN(n6054) );
  AND2_X1 U7551 ( .A1(n6064), .A2(n6054), .ZN(n8181) );
  NAND2_X1 U7552 ( .A1(n8181), .A2(n5848), .ZN(n6060) );
  INV_X1 U7553 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n6057) );
  NAND2_X1 U7554 ( .A1(n5937), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n6056) );
  NAND2_X1 U7555 ( .A1(n6192), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n6055) );
  OAI211_X1 U7556 ( .C1(n5890), .C2(n6057), .A(n6056), .B(n6055), .ZN(n6058)
         );
  INV_X1 U7557 ( .A(n6058), .ZN(n6059) );
  OR2_X1 U7558 ( .A1(n8920), .A2(n8829), .ZN(n6315) );
  NAND2_X1 U7559 ( .A1(n8920), .A2(n8829), .ZN(n6312) );
  NAND2_X1 U7560 ( .A1(n6315), .A2(n6312), .ZN(n8149) );
  NAND2_X1 U7561 ( .A1(n7123), .A2(n6169), .ZN(n6062) );
  NAND2_X1 U7562 ( .A1(n6206), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n6061) );
  INV_X1 U7563 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n10090) );
  NAND2_X1 U7564 ( .A1(n6064), .A2(n10090), .ZN(n6065) );
  NAND2_X1 U7565 ( .A1(n6074), .A2(n6065), .ZN(n8821) );
  OR2_X1 U7566 ( .A1(n8821), .A2(n6152), .ZN(n6071) );
  INV_X1 U7567 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n6068) );
  NAND2_X1 U7568 ( .A1(n6192), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n6067) );
  NAND2_X1 U7569 ( .A1(n5937), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n6066) );
  OAI211_X1 U7570 ( .C1(n5890), .C2(n6068), .A(n6067), .B(n6066), .ZN(n6069)
         );
  INV_X1 U7571 ( .A(n6069), .ZN(n6070) );
  NAND2_X1 U7572 ( .A1(n8913), .A2(n8579), .ZN(n6318) );
  NAND2_X1 U7573 ( .A1(n7170), .A2(n6169), .ZN(n6073) );
  NAND2_X1 U7574 ( .A1(n6206), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n6072) );
  INV_X1 U7575 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n10062) );
  NAND2_X1 U7576 ( .A1(n6074), .A2(n10062), .ZN(n6075) );
  AND2_X1 U7577 ( .A1(n6085), .A2(n6075), .ZN(n8808) );
  NAND2_X1 U7578 ( .A1(n8808), .A2(n5848), .ZN(n6081) );
  INV_X1 U7579 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n6078) );
  NAND2_X1 U7580 ( .A1(n6192), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n6077) );
  NAND2_X1 U7581 ( .A1(n5937), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n6076) );
  OAI211_X1 U7582 ( .C1(n5890), .C2(n6078), .A(n6077), .B(n6076), .ZN(n6079)
         );
  INV_X1 U7583 ( .A(n6079), .ZN(n6080) );
  NAND2_X1 U7584 ( .A1(n6081), .A2(n6080), .ZN(n8637) );
  XNOR2_X1 U7585 ( .A(n8908), .B(n8637), .ZN(n8806) );
  INV_X1 U7586 ( .A(n8637), .ZN(n8831) );
  AND2_X1 U7587 ( .A1(n8908), .A2(n8831), .ZN(n6305) );
  AOI21_X1 U7588 ( .B1(n8803), .B2(n8806), .A(n6305), .ZN(n8794) );
  NAND2_X1 U7589 ( .A1(n7432), .A2(n6169), .ZN(n6083) );
  NAND2_X1 U7590 ( .A1(n6206), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n6082) );
  INV_X1 U7591 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n8614) );
  NAND2_X1 U7592 ( .A1(n6085), .A2(n8614), .ZN(n6086) );
  NAND2_X1 U7593 ( .A1(n6096), .A2(n6086), .ZN(n8791) );
  OR2_X1 U7594 ( .A1(n8791), .A2(n6152), .ZN(n6092) );
  INV_X1 U7595 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n6089) );
  NAND2_X1 U7596 ( .A1(n6030), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n6088) );
  NAND2_X1 U7597 ( .A1(n5937), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n6087) );
  OAI211_X1 U7598 ( .C1(n5888), .C2(n6089), .A(n6088), .B(n6087), .ZN(n6090)
         );
  INV_X1 U7599 ( .A(n6090), .ZN(n6091) );
  NAND2_X1 U7600 ( .A1(n8903), .A2(n8775), .ZN(n6308) );
  NAND2_X1 U7601 ( .A1(n8794), .A2(n8786), .ZN(n8798) );
  NAND2_X1 U7602 ( .A1(n7446), .A2(n6169), .ZN(n6094) );
  NAND2_X1 U7603 ( .A1(n6206), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n6093) );
  INV_X1 U7604 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n6095) );
  NAND2_X1 U7605 ( .A1(n6096), .A2(n6095), .ZN(n6097) );
  AND2_X1 U7606 ( .A1(n6107), .A2(n6097), .ZN(n8778) );
  NAND2_X1 U7607 ( .A1(n8778), .A2(n5848), .ZN(n6102) );
  INV_X1 U7608 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n10001) );
  NAND2_X1 U7609 ( .A1(n6030), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n6099) );
  NAND2_X1 U7610 ( .A1(n5937), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n6098) );
  OAI211_X1 U7611 ( .C1(n10001), .C2(n5888), .A(n6099), .B(n6098), .ZN(n6100)
         );
  INV_X1 U7612 ( .A(n6100), .ZN(n6101) );
  NAND2_X1 U7613 ( .A1(n8896), .A2(n8613), .ZN(n6311) );
  INV_X1 U7614 ( .A(n6311), .ZN(n6103) );
  NAND2_X1 U7615 ( .A1(n7642), .A2(n6169), .ZN(n6105) );
  NAND2_X1 U7616 ( .A1(n6206), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n6104) );
  INV_X1 U7617 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n8593) );
  NAND2_X1 U7618 ( .A1(n6107), .A2(n8593), .ZN(n6108) );
  NAND2_X1 U7619 ( .A1(n6117), .A2(n6108), .ZN(n8760) );
  OR2_X1 U7620 ( .A1(n8760), .A2(n6152), .ZN(n6114) );
  INV_X1 U7621 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n6111) );
  NAND2_X1 U7622 ( .A1(n5937), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n6110) );
  NAND2_X1 U7623 ( .A1(n6030), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n6109) );
  OAI211_X1 U7624 ( .C1(n5888), .C2(n6111), .A(n6110), .B(n6109), .ZN(n6112)
         );
  INV_X1 U7625 ( .A(n6112), .ZN(n6113) );
  NAND2_X1 U7626 ( .A1(n8891), .A2(n8774), .ZN(n6325) );
  NAND2_X1 U7627 ( .A1(n6206), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n6115) );
  INV_X1 U7628 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8586) );
  NAND2_X1 U7629 ( .A1(n6117), .A2(n8586), .ZN(n6118) );
  NAND2_X1 U7630 ( .A1(n6127), .A2(n6118), .ZN(n8742) );
  OR2_X1 U7631 ( .A1(n8742), .A2(n6152), .ZN(n6123) );
  INV_X1 U7632 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n10003) );
  NAND2_X1 U7633 ( .A1(n6030), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n6120) );
  INV_X1 U7634 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n10120) );
  OR2_X1 U7635 ( .A1(n5875), .A2(n10120), .ZN(n6119) );
  OAI211_X1 U7636 ( .C1(n5888), .C2(n10003), .A(n6120), .B(n6119), .ZN(n6121)
         );
  INV_X1 U7637 ( .A(n6121), .ZN(n6122) );
  NAND2_X1 U7638 ( .A1(n8887), .A2(n8263), .ZN(n6222) );
  NAND2_X1 U7639 ( .A1(n7922), .A2(n6169), .ZN(n6125) );
  NAND2_X1 U7640 ( .A1(n6206), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n6124) );
  INV_X1 U7641 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n6126) );
  NAND2_X1 U7642 ( .A1(n6127), .A2(n6126), .ZN(n6128) );
  NAND2_X1 U7643 ( .A1(n8732), .A2(n5848), .ZN(n6134) );
  INV_X1 U7644 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n6131) );
  NAND2_X1 U7645 ( .A1(n5937), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n6130) );
  NAND2_X1 U7646 ( .A1(n6030), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n6129) );
  OAI211_X1 U7647 ( .C1(n5888), .C2(n6131), .A(n6130), .B(n6129), .ZN(n6132)
         );
  INV_X1 U7648 ( .A(n6132), .ZN(n6133) );
  NAND2_X1 U7649 ( .A1(n8883), .A2(n8714), .ZN(n6135) );
  INV_X1 U7650 ( .A(n6135), .ZN(n6136) );
  NAND2_X1 U7651 ( .A1(n6206), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n6137) );
  XNOR2_X1 U7652 ( .A(n6150), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n8711) );
  INV_X1 U7653 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n10097) );
  NAND2_X1 U7654 ( .A1(n6030), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n6140) );
  NAND2_X1 U7655 ( .A1(n5937), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n6139) );
  OAI211_X1 U7656 ( .C1(n10097), .C2(n5888), .A(n6140), .B(n6139), .ZN(n6141)
         );
  NAND2_X1 U7657 ( .A1(n8876), .A2(n8702), .ZN(n6338) );
  MUX2_X1 U7658 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(P1_DATAO_REG_28__SCAN_IN), 
        .S(n6607), .Z(n6162) );
  INV_X1 U7659 ( .A(SI_28_), .ZN(n6163) );
  XNOR2_X1 U7660 ( .A(n6162), .B(n6163), .ZN(n6160) );
  NAND2_X1 U7661 ( .A1(n6484), .A2(n6169), .ZN(n6146) );
  NAND2_X1 U7662 ( .A1(n6206), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n6145) );
  INV_X1 U7663 ( .A(n6150), .ZN(n6148) );
  AND2_X1 U7664 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .ZN(n6147) );
  NAND2_X1 U7665 ( .A1(n6148), .A2(n6147), .ZN(n6172) );
  INV_X1 U7666 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n10178) );
  INV_X1 U7667 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n6149) );
  OAI21_X1 U7668 ( .B1(n6150), .B2(n10178), .A(n6149), .ZN(n6151) );
  NAND2_X1 U7669 ( .A1(n6172), .A2(n6151), .ZN(n8279) );
  OR2_X1 U7670 ( .A1(n8279), .A2(n6152), .ZN(n6157) );
  INV_X1 U7671 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n10076) );
  NAND2_X1 U7672 ( .A1(n5847), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6154) );
  NAND2_X1 U7673 ( .A1(n6030), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n6153) );
  OAI211_X1 U7674 ( .C1(n5888), .C2(n10076), .A(n6154), .B(n6153), .ZN(n6155)
         );
  INV_X1 U7675 ( .A(n6155), .ZN(n6156) );
  NAND2_X1 U7676 ( .A1(n8698), .A2(n8692), .ZN(n8704) );
  NAND2_X1 U7677 ( .A1(n8704), .A2(n6159), .ZN(n6466) );
  INV_X1 U7678 ( .A(n6162), .ZN(n6164) );
  NAND2_X1 U7679 ( .A1(n6164), .A2(n6163), .ZN(n6165) );
  INV_X1 U7680 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n10023) );
  INV_X1 U7681 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n6167) );
  MUX2_X1 U7682 ( .A(n10023), .B(n6167), .S(n6607), .Z(n6177) );
  XNOR2_X1 U7683 ( .A(n6177), .B(SI_29_), .ZN(n6168) );
  NAND2_X1 U7684 ( .A1(n8390), .A2(n6169), .ZN(n6171) );
  NAND2_X1 U7685 ( .A1(n6206), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n6170) );
  INV_X1 U7686 ( .A(n6172), .ZN(n6478) );
  INV_X1 U7687 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n6175) );
  NAND2_X1 U7688 ( .A1(n6192), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6174) );
  INV_X1 U7689 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n10133) );
  OR2_X1 U7690 ( .A1(n5875), .A2(n10133), .ZN(n6173) );
  OAI211_X1 U7691 ( .C1(n5890), .C2(n6175), .A(n6174), .B(n6173), .ZN(n6176)
         );
  AOI21_X1 U7692 ( .B1(n6478), .B2(n5848), .A(n6176), .ZN(n8701) );
  NOR2_X1 U7693 ( .A1(n8867), .A2(n8701), .ZN(n6221) );
  NAND2_X1 U7694 ( .A1(n8867), .A2(n8701), .ZN(n6346) );
  OAI21_X1 U7695 ( .B1(n6466), .B2(n6221), .A(n6346), .ZN(n6195) );
  INV_X1 U7696 ( .A(n6177), .ZN(n6178) );
  NOR2_X1 U7697 ( .A1(n6178), .A2(SI_29_), .ZN(n6180) );
  NAND2_X1 U7698 ( .A1(n6178), .A2(SI_29_), .ZN(n6179) );
  MUX2_X1 U7699 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n6607), .Z(n6199) );
  NAND2_X1 U7700 ( .A1(n8554), .A2(n6169), .ZN(n6183) );
  NAND2_X1 U7701 ( .A1(n6206), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n6182) );
  NAND2_X1 U7702 ( .A1(n6192), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n6186) );
  NAND2_X1 U7703 ( .A1(n6030), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n6185) );
  NAND2_X1 U7704 ( .A1(n5937), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n6184) );
  AND3_X1 U7705 ( .A1(n6186), .A2(n6185), .A3(n6184), .ZN(n6469) );
  NOR2_X1 U7706 ( .A1(n8688), .A2(n6469), .ZN(n6217) );
  NAND2_X1 U7707 ( .A1(n6215), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6191) );
  INV_X1 U7708 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n10208) );
  NAND2_X1 U7709 ( .A1(n6030), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n6194) );
  NAND2_X1 U7710 ( .A1(n6192), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n6193) );
  OAI211_X1 U7711 ( .C1(n5875), .C2(n10208), .A(n6194), .B(n6193), .ZN(n8681)
         );
  INV_X1 U7712 ( .A(n8688), .ZN(n6196) );
  INV_X1 U7713 ( .A(n6197), .ZN(n6198) );
  NAND2_X1 U7714 ( .A1(n6198), .A2(SI_30_), .ZN(n6202) );
  NAND2_X1 U7715 ( .A1(n6200), .A2(n6199), .ZN(n6201) );
  NAND2_X1 U7716 ( .A1(n6202), .A2(n6201), .ZN(n6205) );
  MUX2_X1 U7717 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n6607), .Z(n6203) );
  XNOR2_X1 U7718 ( .A(n6203), .B(SI_31_), .ZN(n6204) );
  NAND2_X1 U7719 ( .A1(n8964), .A2(n6169), .ZN(n6208) );
  NAND2_X1 U7720 ( .A1(n6206), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n6207) );
  INV_X1 U7721 ( .A(n8681), .ZN(n6209) );
  NAND2_X1 U7722 ( .A1(n8688), .A2(n6469), .ZN(n6350) );
  XNOR2_X1 U7723 ( .A(n6210), .B(n9827), .ZN(n6359) );
  NAND2_X1 U7724 ( .A1(n6212), .A2(n6211), .ZN(n6213) );
  NAND2_X1 U7725 ( .A1(n6213), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6214) );
  INV_X1 U7726 ( .A(n7171), .ZN(n6414) );
  NAND2_X1 U7727 ( .A1(n7087), .A2(n6414), .ZN(n6468) );
  NAND2_X1 U7728 ( .A1(n8274), .A2(n6468), .ZN(n6358) );
  INV_X1 U7729 ( .A(n6355), .ZN(n6218) );
  INV_X1 U7730 ( .A(n6217), .ZN(n6351) );
  NAND2_X1 U7731 ( .A1(n8734), .A2(n6414), .ZN(n6220) );
  OR2_X1 U7732 ( .A1(n6219), .A2(n6220), .ZN(n6353) );
  MUX2_X1 U7733 ( .A(n6360), .B(n6361), .S(n6353), .Z(n6357) );
  INV_X1 U7734 ( .A(n6221), .ZN(n6347) );
  INV_X1 U7735 ( .A(n6353), .ZN(n6342) );
  OR3_X1 U7736 ( .A1(n8871), .A2(n8715), .A3(n6342), .ZN(n6345) );
  INV_X1 U7737 ( .A(n6222), .ZN(n6223) );
  OAI21_X1 U7738 ( .B1(n6446), .B2(n6223), .A(n6353), .ZN(n6333) );
  INV_X1 U7739 ( .A(n6224), .ZN(n6299) );
  NAND2_X1 U7740 ( .A1(n6293), .A2(n6299), .ZN(n7944) );
  MUX2_X1 U7741 ( .A(n4754), .B(n6226), .S(n6342), .Z(n6225) );
  NOR2_X1 U7742 ( .A1(n7944), .A2(n6225), .ZN(n6295) );
  INV_X1 U7743 ( .A(n6226), .ZN(n6228) );
  AND2_X1 U7744 ( .A1(n6275), .A2(n6266), .ZN(n6229) );
  MUX2_X1 U7745 ( .A(n6267), .B(n6229), .S(n6353), .Z(n6230) );
  AND2_X1 U7746 ( .A1(n6230), .A2(n6270), .ZN(n6269) );
  NAND2_X1 U7747 ( .A1(n6235), .A2(n6234), .ZN(n6232) );
  NAND2_X1 U7748 ( .A1(n6252), .A2(n7093), .ZN(n6231) );
  MUX2_X1 U7749 ( .A(n6232), .B(n6231), .S(n6353), .Z(n6254) );
  NAND2_X1 U7750 ( .A1(n6236), .A2(n6353), .ZN(n6243) );
  INV_X1 U7751 ( .A(n6254), .ZN(n6241) );
  NAND2_X1 U7752 ( .A1(n6419), .A2(n7197), .ZN(n6939) );
  AND2_X1 U7753 ( .A1(n6939), .A2(n6414), .ZN(n6238) );
  OAI211_X1 U7754 ( .C1(n6238), .C2(n6237), .A(n6246), .B(n6367), .ZN(n6239)
         );
  NAND3_X1 U7755 ( .A1(n6239), .A2(n6244), .A3(n6353), .ZN(n6240) );
  NAND3_X1 U7756 ( .A1(n6241), .A2(n7496), .A3(n6240), .ZN(n6242) );
  NAND2_X1 U7757 ( .A1(n6243), .A2(n6242), .ZN(n6249) );
  OR2_X1 U7758 ( .A1(n7221), .A2(n7029), .ZN(n6251) );
  NAND2_X1 U7759 ( .A1(n6939), .A2(n6367), .ZN(n6245) );
  NAND3_X1 U7760 ( .A1(n6245), .A2(n6244), .A3(n6368), .ZN(n6247) );
  NAND3_X1 U7761 ( .A1(n6247), .A2(n6342), .A3(n6246), .ZN(n6248) );
  NAND3_X1 U7762 ( .A1(n6249), .A2(n6251), .A3(n6248), .ZN(n6257) );
  NAND2_X1 U7763 ( .A1(n8654), .A2(n5870), .ZN(n6250) );
  AND2_X1 U7764 ( .A1(n7093), .A2(n6250), .ZN(n6253) );
  OAI211_X1 U7765 ( .C1(n6254), .C2(n6253), .A(n6252), .B(n6251), .ZN(n6255)
         );
  NAND2_X1 U7766 ( .A1(n6255), .A2(n6342), .ZN(n6256) );
  NAND2_X1 U7767 ( .A1(n6257), .A2(n6256), .ZN(n6258) );
  OAI211_X1 U7768 ( .C1(n6353), .C2(n6259), .A(n6258), .B(n6429), .ZN(n6263)
         );
  MUX2_X1 U7769 ( .A(n6261), .B(n6260), .S(n6342), .Z(n6262) );
  MUX2_X1 U7770 ( .A(n6264), .B(n7477), .S(n6342), .Z(n6265) );
  INV_X1 U7771 ( .A(n6267), .ZN(n6268) );
  NAND2_X1 U7772 ( .A1(n6269), .A2(n6268), .ZN(n6271) );
  AND2_X1 U7773 ( .A1(n6364), .A2(n6366), .ZN(n6273) );
  INV_X1 U7774 ( .A(n6365), .ZN(n6272) );
  AOI21_X1 U7775 ( .B1(n6274), .B2(n6273), .A(n6272), .ZN(n6281) );
  NAND3_X1 U7776 ( .A1(n6276), .A2(n6366), .A3(n6275), .ZN(n6279) );
  INV_X1 U7777 ( .A(n6364), .ZN(n6277) );
  AOI21_X1 U7778 ( .B1(n6279), .B2(n6278), .A(n6277), .ZN(n6280) );
  MUX2_X1 U7779 ( .A(n6281), .B(n6280), .S(n6342), .Z(n6282) );
  NAND2_X1 U7780 ( .A1(n6282), .A2(n7742), .ZN(n6288) );
  INV_X1 U7781 ( .A(n6283), .ZN(n6284) );
  MUX2_X1 U7782 ( .A(n6285), .B(n6284), .S(n6342), .Z(n6286) );
  INV_X1 U7783 ( .A(n6286), .ZN(n6287) );
  NAND3_X1 U7784 ( .A1(n6288), .A2(n7804), .A3(n6287), .ZN(n6292) );
  NAND2_X1 U7785 ( .A1(n8642), .A2(n6353), .ZN(n6290) );
  NAND2_X1 U7786 ( .A1(n7843), .A2(n6342), .ZN(n6289) );
  MUX2_X1 U7787 ( .A(n6290), .B(n6289), .S(n9528), .Z(n6291) );
  NAND3_X1 U7788 ( .A1(n7841), .A2(n6292), .A3(n6291), .ZN(n6294) );
  AOI22_X1 U7789 ( .A1(n6295), .A2(n6294), .B1(n4752), .B2(n6353), .ZN(n6304)
         );
  INV_X1 U7790 ( .A(n6297), .ZN(n6362) );
  OAI211_X1 U7791 ( .C1(n8030), .C2(n6299), .A(n6362), .B(n6298), .ZN(n6300)
         );
  MUX2_X1 U7792 ( .A(n6301), .B(n6300), .S(n6342), .Z(n6302) );
  INV_X1 U7793 ( .A(n6302), .ZN(n6303) );
  OAI21_X1 U7794 ( .B1(n6304), .B2(n8030), .A(n6303), .ZN(n6314) );
  OR2_X1 U7795 ( .A1(n8908), .A2(n8831), .ZN(n6321) );
  INV_X1 U7796 ( .A(n6305), .ZN(n6317) );
  NAND3_X1 U7797 ( .A1(n6306), .A2(n6308), .A3(n6317), .ZN(n6307) );
  NAND2_X1 U7798 ( .A1(n6307), .A2(n6322), .ZN(n6310) );
  INV_X1 U7799 ( .A(n6308), .ZN(n6309) );
  INV_X1 U7800 ( .A(n6312), .ZN(n6313) );
  AOI21_X1 U7801 ( .B1(n6314), .B2(n6363), .A(n6313), .ZN(n6320) );
  NAND2_X1 U7802 ( .A1(n6316), .A2(n6315), .ZN(n6319) );
  OAI211_X1 U7803 ( .C1(n6320), .C2(n6319), .A(n6318), .B(n6317), .ZN(n6323)
         );
  NAND4_X1 U7804 ( .A1(n6323), .A2(n6322), .A3(n6342), .A4(n6321), .ZN(n6324)
         );
  INV_X1 U7805 ( .A(n6327), .ZN(n8743) );
  AOI21_X1 U7806 ( .B1(n6327), .B2(n6326), .A(n6353), .ZN(n6329) );
  NAND3_X1 U7807 ( .A1(n8891), .A2(n8774), .A3(n6342), .ZN(n6328) );
  OAI211_X1 U7808 ( .C1(n6330), .C2(n6329), .A(n8744), .B(n6328), .ZN(n6332)
         );
  INV_X1 U7809 ( .A(n6334), .ZN(n6331) );
  AOI21_X1 U7810 ( .B1(n6333), .B2(n6332), .A(n6331), .ZN(n6337) );
  AOI21_X1 U7811 ( .B1(n6334), .B2(n8723), .A(n6353), .ZN(n6336) );
  NAND3_X1 U7812 ( .A1(n8883), .A2(n8714), .A3(n6342), .ZN(n6335) );
  OAI211_X1 U7813 ( .C1(n6337), .C2(n6336), .A(n6447), .B(n6335), .ZN(n6341)
         );
  MUX2_X1 U7814 ( .A(n6339), .B(n6338), .S(n6353), .Z(n6340) );
  NAND3_X1 U7815 ( .A1(n6341), .A2(n8692), .A3(n6340), .ZN(n6344) );
  NAND3_X1 U7816 ( .A1(n8871), .A2(n8715), .A3(n6342), .ZN(n6343) );
  NAND4_X1 U7817 ( .A1(n6467), .A2(n6345), .A3(n6344), .A4(n6343), .ZN(n6349)
         );
  MUX2_X1 U7818 ( .A(n6347), .B(n6346), .S(n6353), .Z(n6348) );
  INV_X1 U7819 ( .A(n6352), .ZN(n6354) );
  MUX2_X1 U7820 ( .A(n6355), .B(n6354), .S(n6353), .Z(n6356) );
  INV_X1 U7821 ( .A(n6360), .ZN(n6385) );
  INV_X1 U7822 ( .A(n6361), .ZN(n6384) );
  INV_X1 U7823 ( .A(n8806), .ZN(n6379) );
  INV_X1 U7824 ( .A(n8827), .ZN(n6377) );
  INV_X1 U7825 ( .A(n8149), .ZN(n8151) );
  NAND2_X1 U7826 ( .A1(n6365), .A2(n6364), .ZN(n6437) );
  NAND2_X1 U7827 ( .A1(n7567), .A2(n6366), .ZN(n7630) );
  INV_X1 U7828 ( .A(n6432), .ZN(n7611) );
  INV_X1 U7829 ( .A(n7552), .ZN(n6371) );
  AND2_X1 U7830 ( .A1(n6938), .A2(n6939), .ZN(n7341) );
  AND2_X2 U7831 ( .A1(n6368), .A2(n6367), .ZN(n7203) );
  AND4_X1 U7832 ( .A1(n7341), .A2(n7203), .A3(n7087), .A4(n7310), .ZN(n6369)
         );
  INV_X1 U7833 ( .A(n7356), .ZN(n7358) );
  NAND4_X1 U7834 ( .A1(n6369), .A2(n7086), .A3(n7358), .A4(n7496), .ZN(n6370)
         );
  INV_X1 U7835 ( .A(n6429), .ZN(n7125) );
  NOR3_X1 U7836 ( .A1(n6371), .A2(n6370), .A3(n7125), .ZN(n6372) );
  NAND4_X1 U7837 ( .A1(n7611), .A2(n7472), .A3(n6372), .A4(n7222), .ZN(n6373)
         );
  NOR4_X1 U7838 ( .A1(n4898), .A2(n6437), .A3(n7630), .A4(n6373), .ZN(n6374)
         );
  NAND4_X1 U7839 ( .A1(n7949), .A2(n7841), .A3(n6374), .A4(n7804), .ZN(n6375)
         );
  NOR2_X1 U7840 ( .A1(n6375), .A2(n8030), .ZN(n6376) );
  NAND4_X1 U7841 ( .A1(n6377), .A2(n8151), .A3(n8853), .A4(n6376), .ZN(n6378)
         );
  NOR4_X1 U7842 ( .A1(n8782), .A2(n8795), .A3(n6379), .A4(n6378), .ZN(n6380)
         );
  NAND4_X1 U7843 ( .A1(n4767), .A2(n8744), .A3(n8765), .A4(n6380), .ZN(n6381)
         );
  NOR2_X1 U7844 ( .A1(n8713), .A2(n6381), .ZN(n6382) );
  NAND3_X1 U7845 ( .A1(n6467), .A2(n6382), .A3(n8692), .ZN(n6383) );
  NOR3_X1 U7846 ( .A1(n6385), .A2(n6384), .A3(n6383), .ZN(n6386) );
  XNOR2_X1 U7847 ( .A(n6386), .B(n9827), .ZN(n6390) );
  INV_X1 U7848 ( .A(n6387), .ZN(n6389) );
  AOI22_X1 U7849 ( .A1(n6390), .A2(n7171), .B1(n6389), .B2(n6388), .ZN(n6391)
         );
  INV_X1 U7850 ( .A(n6391), .ZN(n6394) );
  NAND2_X1 U7851 ( .A1(n6394), .A2(n6393), .ZN(n6395) );
  NAND2_X1 U7852 ( .A1(n6396), .A2(n6395), .ZN(n6400) );
  NAND2_X1 U7853 ( .A1(n6397), .A2(n6405), .ZN(n6398) );
  NAND2_X1 U7854 ( .A1(n6398), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6401) );
  XNOR2_X1 U7855 ( .A(n6401), .B(P2_IR_REG_23__SCAN_IN), .ZN(n7013) );
  NAND2_X1 U7856 ( .A1(n7013), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7514) );
  NAND2_X1 U7857 ( .A1(n6400), .A2(n6399), .ZN(n6418) );
  NAND2_X1 U7858 ( .A1(n6401), .A2(n6406), .ZN(n6402) );
  NAND2_X1 U7859 ( .A1(n6402), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6403) );
  XNOR2_X1 U7860 ( .A(n6403), .B(P2_IR_REG_24__SCAN_IN), .ZN(n6449) );
  INV_X1 U7861 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6404) );
  NAND3_X1 U7862 ( .A1(n6406), .A2(n6405), .A3(n6404), .ZN(n6407) );
  OAI21_X1 U7863 ( .B1(n6408), .B2(n6407), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n6409) );
  MUX2_X1 U7864 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6409), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n6411) );
  AND2_X1 U7865 ( .A1(n6411), .A2(n6410), .ZN(n9841) );
  NAND2_X1 U7866 ( .A1(n6410), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6412) );
  XNOR2_X1 U7867 ( .A(n6412), .B(P2_IR_REG_26__SCAN_IN), .ZN(n9842) );
  AND2_X1 U7868 ( .A1(n9841), .A2(n9842), .ZN(n6413) );
  NAND2_X1 U7869 ( .A1(n6449), .A2(n6413), .ZN(n7015) );
  NOR2_X1 U7870 ( .A1(n7013), .A2(P2_U3152), .ZN(n9845) );
  NAND2_X1 U7871 ( .A1(n7015), .A2(n9845), .ZN(n9838) );
  NAND2_X1 U7872 ( .A1(n6219), .A2(n6414), .ZN(n6941) );
  OR2_X1 U7873 ( .A1(n6941), .A2(n8240), .ZN(n8828) );
  NOR4_X1 U7874 ( .A1(n9838), .A2(n7941), .A3(n6936), .A4(n8828), .ZN(n6416)
         );
  OAI21_X1 U7875 ( .B1(n7514), .B2(n6219), .A(P2_B_REG_SCAN_IN), .ZN(n6415) );
  NAND2_X1 U7876 ( .A1(n6418), .A2(n6417), .ZN(P2_U3244) );
  INV_X1 U7877 ( .A(n8908), .ZN(n8811) );
  INV_X1 U7878 ( .A(n8120), .ZN(n8641) );
  INV_X1 U7879 ( .A(n7197), .ZN(n9847) );
  NAND2_X1 U7880 ( .A1(n6419), .A2(n9847), .ZN(n6950) );
  INV_X1 U7881 ( .A(n6950), .ZN(n7202) );
  NAND2_X1 U7882 ( .A1(n7306), .A2(n7307), .ZN(n6421) );
  INV_X1 U7883 ( .A(n9858), .ZN(n7312) );
  OR2_X1 U7884 ( .A1(n8655), .A2(n7312), .ZN(n6420) );
  NAND2_X1 U7885 ( .A1(n6421), .A2(n6420), .ZN(n7492) );
  NAND2_X1 U7886 ( .A1(n7492), .A2(n7493), .ZN(n6423) );
  OR2_X1 U7887 ( .A1(n8654), .A2(n7510), .ZN(n6422) );
  NAND2_X1 U7888 ( .A1(n6423), .A2(n6422), .ZN(n7355) );
  NAND2_X1 U7889 ( .A1(n7355), .A2(n7356), .ZN(n6425) );
  INV_X1 U7890 ( .A(n8653), .ZN(n7147) );
  NAND2_X1 U7891 ( .A1(n7147), .A2(n9869), .ZN(n6424) );
  NAND2_X1 U7892 ( .A1(n6425), .A2(n6424), .ZN(n7085) );
  NAND2_X1 U7893 ( .A1(n7211), .A2(n9823), .ZN(n6426) );
  NAND2_X1 U7894 ( .A1(n7221), .A2(n8651), .ZN(n6427) );
  NAND2_X1 U7895 ( .A1(n6428), .A2(n6427), .ZN(n7124) );
  INV_X1 U7896 ( .A(n7554), .ZN(n8650) );
  OAI22_X1 U7897 ( .A1(n7124), .A2(n6429), .B1(n7129), .B2(n8650), .ZN(n7547)
         );
  INV_X1 U7898 ( .A(n7474), .ZN(n8649) );
  NAND2_X1 U7899 ( .A1(n9881), .A2(n8649), .ZN(n6430) );
  NAND2_X1 U7900 ( .A1(n7549), .A2(n6430), .ZN(n7471) );
  INV_X1 U7901 ( .A(n7473), .ZN(n8647) );
  AND2_X1 U7902 ( .A1(n9891), .A2(n8647), .ZN(n6433) );
  OR2_X1 U7903 ( .A1(n7472), .A2(n6433), .ZN(n7626) );
  INV_X1 U7904 ( .A(n7707), .ZN(n8646) );
  AND2_X1 U7905 ( .A1(n7670), .A2(n8646), .ZN(n6435) );
  OR2_X1 U7906 ( .A1(n7626), .A2(n6435), .ZN(n6431) );
  INV_X1 U7907 ( .A(n7553), .ZN(n8648) );
  OR2_X1 U7908 ( .A1(n7646), .A2(n8648), .ZN(n7606) );
  AND2_X1 U7909 ( .A1(n6432), .A2(n7606), .ZN(n7605) );
  OR2_X1 U7910 ( .A1(n6433), .A2(n7605), .ZN(n7628) );
  AND2_X1 U7911 ( .A1(n7630), .A2(n7628), .ZN(n6434) );
  NOR2_X1 U7912 ( .A1(n6435), .A2(n6434), .ZN(n6436) );
  INV_X1 U7913 ( .A(n7760), .ZN(n8645) );
  NAND2_X1 U7914 ( .A1(n7763), .A2(n8644), .ZN(n6438) );
  NAND2_X1 U7915 ( .A1(n7848), .A2(n7847), .ZN(n7846) );
  OAI21_X1 U7916 ( .B1(n9521), .B2(n8641), .A(n7846), .ZN(n7948) );
  INV_X1 U7917 ( .A(n8132), .ZN(n8839) );
  INV_X1 U7918 ( .A(n8179), .ZN(n8639) );
  NAND2_X1 U7919 ( .A1(n8923), .A2(n8639), .ZN(n6440) );
  INV_X1 U7920 ( .A(n8923), .ZN(n8852) );
  INV_X1 U7921 ( .A(n8829), .ZN(n8841) );
  INV_X1 U7922 ( .A(n8920), .ZN(n8184) );
  NAND2_X1 U7923 ( .A1(n6442), .A2(n4922), .ZN(n8816) );
  INV_X1 U7924 ( .A(n8579), .ZN(n8804) );
  NAND2_X1 U7925 ( .A1(n8783), .A2(n8782), .ZN(n8898) );
  INV_X1 U7926 ( .A(n8896), .ZN(n8780) );
  INV_X1 U7927 ( .A(n8702), .ZN(n8635) );
  INV_X1 U7928 ( .A(n8692), .ZN(n8699) );
  NOR2_X1 U7929 ( .A1(n6449), .A2(n9842), .ZN(n9840) );
  INV_X1 U7930 ( .A(P2_B_REG_SCAN_IN), .ZN(n10015) );
  INV_X1 U7931 ( .A(n6449), .ZN(n7669) );
  INV_X1 U7932 ( .A(n9841), .ZN(n7813) );
  OAI221_X1 U7933 ( .B1(P2_B_REG_SCAN_IN), .B2(n6449), .C1(n10015), .C2(n7669), 
        .A(n7813), .ZN(n6450) );
  INV_X1 U7934 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n10025) );
  AND2_X1 U7935 ( .A1(n9837), .A2(n10025), .ZN(n6451) );
  INV_X1 U7936 ( .A(n9838), .ZN(n6464) );
  INV_X1 U7937 ( .A(n6941), .ZN(n6545) );
  NAND2_X1 U7938 ( .A1(n6545), .A2(n6936), .ZN(n7079) );
  INV_X1 U7939 ( .A(n9842), .ZN(n7923) );
  INV_X1 U7940 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n9844) );
  AND2_X1 U7941 ( .A1(n9837), .A2(n9844), .ZN(n6452) );
  AOI21_X1 U7942 ( .B1(n7813), .B2(n7923), .A(n6452), .ZN(n7078) );
  NOR4_X1 U7943 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_17__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n6456) );
  NOR4_X1 U7944 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_16__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n6455) );
  NOR4_X1 U7945 ( .A1(P2_D_REG_25__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n6454) );
  NOR4_X1 U7946 ( .A1(P2_D_REG_20__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_22__SCAN_IN), .ZN(n6453) );
  NAND4_X1 U7947 ( .A1(n6456), .A2(n6455), .A3(n6454), .A4(n6453), .ZN(n6461)
         );
  NOR2_X1 U7948 ( .A1(P2_D_REG_24__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .ZN(
        n9976) );
  NOR4_X1 U7949 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_31__SCAN_IN), .A3(
        P2_D_REG_14__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n6459) );
  NOR4_X1 U7950 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_5__SCAN_IN), .A3(
        P2_D_REG_6__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n6458) );
  NOR4_X1 U7951 ( .A1(P2_D_REG_12__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_2__SCAN_IN), .A4(P2_D_REG_3__SCAN_IN), .ZN(n6457) );
  NAND4_X1 U7952 ( .A1(n9976), .A2(n6459), .A3(n6458), .A4(n6457), .ZN(n6460)
         );
  OAI21_X1 U7953 ( .B1(n6461), .B2(n6460), .A(n9837), .ZN(n7084) );
  NAND2_X1 U7954 ( .A1(n7078), .A2(n7084), .ZN(n6933) );
  INV_X1 U7955 ( .A(n6933), .ZN(n6462) );
  AND2_X1 U7956 ( .A1(n7079), .A2(n6462), .ZN(n6463) );
  NAND3_X1 U7957 ( .A1(n7104), .A2(n6464), .A3(n6463), .ZN(n6477) );
  OR3_X1 U7958 ( .A1(n6219), .A2(n7087), .A3(n9827), .ZN(n9886) );
  INV_X1 U7959 ( .A(n9886), .ZN(n9897) );
  NAND2_X1 U7960 ( .A1(n9897), .A2(n7171), .ZN(n7080) );
  OR2_X1 U7961 ( .A1(n7087), .A2(n7171), .ZN(n6948) );
  XNOR2_X1 U7962 ( .A(n6948), .B(n6219), .ZN(n6465) );
  NAND2_X1 U7963 ( .A1(n6465), .A2(n9827), .ZN(n7747) );
  OR2_X1 U7964 ( .A1(n6948), .A2(n9827), .ZN(n7489) );
  NAND2_X1 U7965 ( .A1(n7747), .A2(n7489), .ZN(n9819) );
  NAND2_X1 U7966 ( .A1(n9834), .A2(n9819), .ZN(n8855) );
  NAND2_X1 U7967 ( .A1(n6468), .A2(n6387), .ZN(n8843) );
  INV_X1 U7968 ( .A(n8828), .ZN(n8838) );
  INV_X1 U7969 ( .A(n6469), .ZN(n8633) );
  INV_X1 U7970 ( .A(n7941), .ZN(n6471) );
  INV_X1 U7971 ( .A(n8240), .ZN(n6470) );
  OR2_X1 U7972 ( .A1(n6941), .A2(n6470), .ZN(n8830) );
  AOI21_X1 U7973 ( .B1(n6471), .B2(P2_B_REG_SCAN_IN), .A(n8830), .ZN(n8682) );
  INV_X2 U7974 ( .A(n9834), .ZN(n9836) );
  INV_X1 U7975 ( .A(n8913), .ZN(n8824) );
  NAND2_X1 U7976 ( .A1(n6951), .A2(n7197), .ZN(n9852) );
  NAND2_X1 U7977 ( .A1(n7504), .A2(n9869), .ZN(n7089) );
  INV_X1 U7978 ( .A(n7129), .ZN(n7464) );
  INV_X1 U7979 ( .A(n9881), .ZN(n7563) );
  INV_X1 U7980 ( .A(n7700), .ZN(n9900) );
  INV_X1 U7981 ( .A(n9528), .ZN(n7802) );
  NAND2_X1 U7982 ( .A1(n6439), .A2(n8023), .ZN(n8846) );
  NAND2_X1 U7983 ( .A1(n8824), .A2(n8817), .ZN(n8818) );
  NOR2_X2 U7984 ( .A1(n8751), .A2(n8887), .ZN(n8750) );
  AOI21_X1 U7985 ( .B1(n8867), .B2(n8694), .A(n8686), .ZN(n8868) );
  OR2_X1 U7986 ( .A1(n6477), .A2(n8274), .ZN(n8685) );
  NOR2_X1 U7987 ( .A1(n6388), .A2(n7088), .ZN(n9821) );
  NAND2_X1 U7988 ( .A1(n9834), .A2(n9821), .ZN(n8851) );
  INV_X1 U7989 ( .A(n9825), .ZN(n8848) );
  AOI22_X1 U7990 ( .A1(n6478), .A2(n8848), .B1(P2_REG2_REG_29__SCAN_IN), .B2(
        n9836), .ZN(n6479) );
  OAI21_X1 U7991 ( .B1(n4547), .B2(n8851), .A(n6479), .ZN(n6480) );
  AOI21_X1 U7992 ( .B1(n8868), .B2(n8858), .A(n6480), .ZN(n6481) );
  OAI21_X1 U7993 ( .B1(n8869), .B2(n9836), .A(n6481), .ZN(n6482) );
  INV_X1 U7994 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n7977) );
  OR2_X1 U7995 ( .A1(n8391), .A2(n7977), .ZN(n6485) );
  NAND2_X1 U7996 ( .A1(n9179), .A2(n5096), .ZN(n6489) );
  INV_X1 U7997 ( .A(n5640), .ZN(n6487) );
  OR2_X1 U7998 ( .A1(n9157), .A2(n6487), .ZN(n6488) );
  NAND2_X1 U7999 ( .A1(n6489), .A2(n6488), .ZN(n6491) );
  XNOR2_X1 U8000 ( .A(n6491), .B(n6490), .ZN(n6495) );
  NAND2_X1 U8001 ( .A1(n9179), .A2(n6492), .ZN(n6493) );
  OAI21_X1 U8002 ( .B1(n9157), .B2(n4371), .A(n6493), .ZN(n6494) );
  XNOR2_X1 U8003 ( .A(n6495), .B(n6494), .ZN(n6503) );
  NAND3_X1 U8004 ( .A1(n6509), .A2(n5747), .A3(n6503), .ZN(n6512) );
  INV_X1 U8005 ( .A(n9068), .ZN(n9058) );
  AOI22_X1 U8006 ( .A1(n9180), .A2(n9049), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n6502) );
  NAND2_X1 U8007 ( .A1(n8288), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6498) );
  NAND2_X1 U8008 ( .A1(n8289), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6497) );
  NAND2_X1 U8009 ( .A1(n8287), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n6496) );
  AND3_X1 U8010 ( .A1(n6498), .A2(n6497), .A3(n6496), .ZN(n6499) );
  OAI21_X1 U8011 ( .B1(n9163), .B2(n6500), .A(n6499), .ZN(n9078) );
  NAND2_X1 U8012 ( .A1(n9078), .A2(n9067), .ZN(n6501) );
  OAI211_X1 U8013 ( .C1(n9176), .C2(n9058), .A(n6502), .B(n6501), .ZN(n6505)
         );
  INV_X1 U8014 ( .A(n6503), .ZN(n6507) );
  NOR3_X1 U8015 ( .A1(n6507), .A2(n9075), .A3(n6506), .ZN(n6504) );
  AOI211_X1 U8016 ( .C1(n9179), .C2(n9073), .A(n6505), .B(n6504), .ZN(n6511)
         );
  NAND3_X1 U8017 ( .A1(n6507), .A2(n5747), .A3(n6506), .ZN(n6508) );
  NAND3_X1 U8018 ( .A1(n6512), .A2(n6511), .A3(n6510), .ZN(P1_U3218) );
  INV_X1 U8019 ( .A(n7447), .ZN(n6514) );
  OR2_X1 U8020 ( .A1(n6513), .A2(n6514), .ZN(n6525) );
  INV_X1 U8021 ( .A(n9089), .ZN(P1_U4006) );
  OR2_X1 U8022 ( .A1(n7015), .A2(P2_U3152), .ZN(n6544) );
  INV_X2 U8023 ( .A(n8638), .ZN(P2_U3966) );
  OR2_X1 U8024 ( .A1(n8508), .A2(n6514), .ZN(n6515) );
  NAND2_X1 U8025 ( .A1(n6515), .A2(n6525), .ZN(n9602) );
  OR2_X1 U8026 ( .A1(n9602), .A2(n9601), .ZN(n6516) );
  NAND2_X1 U8027 ( .A1(n6516), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  OR2_X1 U8028 ( .A1(n5759), .A2(P1_U3084), .ZN(n7975) );
  INV_X1 U8029 ( .A(n9104), .ZN(n6517) );
  OR2_X1 U8030 ( .A1(n7975), .A2(n6517), .ZN(n6534) );
  INV_X1 U8031 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n10114) );
  AOI21_X1 U8032 ( .B1(n6517), .B2(n10114), .A(n7975), .ZN(n6520) );
  NAND2_X1 U8033 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9949), .ZN(n6601) );
  INV_X1 U8034 ( .A(n6601), .ZN(n6519) );
  AND2_X1 U8035 ( .A1(n9949), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6667) );
  NAND2_X1 U8036 ( .A1(n6764), .A2(n6667), .ZN(n6518) );
  OAI21_X1 U8037 ( .B1(n6520), .B2(n6519), .A(n6518), .ZN(n9603) );
  OAI21_X1 U8038 ( .B1(n6523), .B2(n6521), .A(n6522), .ZN(n8215) );
  NAND2_X1 U8039 ( .A1(n6764), .A2(n9104), .ZN(n9599) );
  NOR2_X1 U8040 ( .A1(n8215), .A2(n9599), .ZN(n6524) );
  AOI211_X1 U8041 ( .C1(n6534), .C2(n9603), .A(n6525), .B(n6524), .ZN(n9620)
         );
  INV_X1 U8042 ( .A(P1_U3083), .ZN(n6526) );
  NAND2_X1 U8043 ( .A1(n6526), .A2(n6525), .ZN(n9699) );
  INV_X1 U8044 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n6527) );
  NOR2_X1 U8045 ( .A1(n9699), .A2(n6527), .ZN(n6542) );
  OR2_X1 U8046 ( .A1(n9104), .A2(P1_U3084), .ZN(n7937) );
  NOR2_X1 U8047 ( .A1(n9602), .A2(n7937), .ZN(n6532) );
  NAND2_X1 U8048 ( .A1(n6532), .A2(n6764), .ZN(n9659) );
  XNOR2_X1 U8049 ( .A(n6605), .B(P1_REG2_REG_2__SCAN_IN), .ZN(n6530) );
  XNOR2_X1 U8050 ( .A(n6603), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n6668) );
  NAND2_X1 U8051 ( .A1(n6668), .A2(n6667), .ZN(n6666) );
  INV_X1 U8052 ( .A(n6603), .ZN(n6665) );
  NAND2_X1 U8053 ( .A1(n6665), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6528) );
  NAND2_X1 U8054 ( .A1(n6666), .A2(n6528), .ZN(n6529) );
  NAND2_X1 U8055 ( .A1(n6530), .A2(n6529), .ZN(n6673) );
  OAI21_X1 U8056 ( .B1(n6530), .B2(n6529), .A(n6673), .ZN(n6531) );
  NOR2_X1 U8057 ( .A1(n9659), .A2(n6531), .ZN(n6541) );
  INV_X1 U8058 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n6539) );
  INV_X1 U8059 ( .A(n6532), .ZN(n9100) );
  INV_X1 U8060 ( .A(n6605), .ZN(n6676) );
  NAND2_X1 U8061 ( .A1(n9686), .A2(n6676), .ZN(n6538) );
  XNOR2_X1 U8062 ( .A(n6605), .B(P1_REG1_REG_2__SCAN_IN), .ZN(n6536) );
  XNOR2_X1 U8063 ( .A(n6603), .B(P1_REG1_REG_1__SCAN_IN), .ZN(n6662) );
  AND2_X1 U8064 ( .A1(n9949), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6661) );
  NAND2_X1 U8065 ( .A1(n6662), .A2(n6661), .ZN(n6660) );
  NAND2_X1 U8066 ( .A1(n6665), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6533) );
  NAND2_X1 U8067 ( .A1(n6660), .A2(n6533), .ZN(n6535) );
  OR2_X1 U8068 ( .A1(n9602), .A2(n6534), .ZN(n9636) );
  INV_X1 U8069 ( .A(n9636), .ZN(n9694) );
  NAND2_X1 U8070 ( .A1(n6536), .A2(n6535), .ZN(n6678) );
  OAI211_X1 U8071 ( .C1(n6536), .C2(n6535), .A(n9694), .B(n6678), .ZN(n6537)
         );
  OAI211_X1 U8072 ( .C1(P1_STATE_REG_SCAN_IN), .C2(n6539), .A(n6538), .B(n6537), .ZN(n6540) );
  OR4_X1 U8073 ( .A1(n9620), .A2(n6542), .A3(n6541), .A4(n6540), .ZN(P1_U3243)
         );
  INV_X1 U8074 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n10230) );
  AOI22_X1 U8075 ( .A1(n6556), .A2(n5826), .B1(P2_REG2_REG_2__SCAN_IN), .B2(
        n9487), .ZN(n9479) );
  NOR2_X1 U8076 ( .A1(n9478), .A2(n9479), .ZN(n9477) );
  INV_X1 U8077 ( .A(n6557), .ZN(n6794) );
  AOI22_X1 U8078 ( .A1(n6557), .A2(n5862), .B1(P2_REG2_REG_3__SCAN_IN), .B2(
        n6794), .ZN(n6786) );
  NOR2_X1 U8079 ( .A1(n6785), .A2(n6786), .ZN(n6784) );
  INV_X1 U8080 ( .A(n6559), .ZN(n6612) );
  AOI22_X1 U8081 ( .A1(n6559), .A2(n5889), .B1(P2_REG2_REG_4__SCAN_IN), .B2(
        n6612), .ZN(n6574) );
  NOR2_X1 U8082 ( .A1(n6575), .A2(n6574), .ZN(n6573) );
  NAND2_X1 U8083 ( .A1(n6586), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6543) );
  OAI21_X1 U8084 ( .B1(n6586), .B2(P2_REG2_REG_5__SCAN_IN), .A(n6543), .ZN(
        n6548) );
  NOR2_X1 U8085 ( .A1(n6549), .A2(n6548), .ZN(n6583) );
  OAI211_X1 U8086 ( .C1(n9838), .C2(n6545), .A(n7514), .B(n6544), .ZN(n6562)
         );
  NAND2_X1 U8087 ( .A1(n6562), .A2(n6565), .ZN(n6546) );
  NAND2_X1 U8088 ( .A1(n6546), .A2(n8638), .ZN(n6550) );
  NOR2_X1 U8089 ( .A1(n8240), .A2(n7941), .ZN(n6547) );
  AND2_X1 U8090 ( .A1(n6550), .A2(n6547), .ZN(n9808) );
  INV_X1 U8091 ( .A(n9808), .ZN(n8657) );
  AOI211_X1 U8092 ( .C1(n6549), .C2(n6548), .A(n6583), .B(n8657), .ZN(n6572)
         );
  NAND2_X1 U8093 ( .A1(n6550), .A2(n8240), .ZN(n9809) );
  INV_X1 U8094 ( .A(n6586), .ZN(n6619) );
  NOR2_X1 U8095 ( .A1(n9809), .A2(n6619), .ZN(n6571) );
  NAND2_X1 U8096 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n9468) );
  INV_X1 U8097 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6551) );
  NAND2_X1 U8098 ( .A1(n9473), .A2(n6551), .ZN(n6553) );
  NAND2_X1 U8099 ( .A1(n6554), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6552) );
  NAND2_X1 U8100 ( .A1(n6553), .A2(n6552), .ZN(n9469) );
  NOR2_X1 U8101 ( .A1(n9468), .A2(n9469), .ZN(n9467) );
  AOI21_X1 U8102 ( .B1(n6554), .B2(P2_REG1_REG_1__SCAN_IN), .A(n9467), .ZN(
        n9482) );
  NAND2_X1 U8103 ( .A1(n6556), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6555) );
  OAI21_X1 U8104 ( .B1(n6556), .B2(P2_REG1_REG_2__SCAN_IN), .A(n6555), .ZN(
        n9483) );
  NOR2_X1 U8105 ( .A1(n9482), .A2(n9483), .ZN(n9481) );
  AOI21_X1 U8106 ( .B1(n6556), .B2(P2_REG1_REG_2__SCAN_IN), .A(n9481), .ZN(
        n6790) );
  MUX2_X1 U8107 ( .A(n5861), .B(P2_REG1_REG_3__SCAN_IN), .S(n6557), .Z(n6789)
         );
  NOR2_X1 U8108 ( .A1(n6790), .A2(n6789), .ZN(n6788) );
  AOI21_X1 U8109 ( .B1(n6557), .B2(P2_REG1_REG_3__SCAN_IN), .A(n6788), .ZN(
        n6578) );
  NAND2_X1 U8110 ( .A1(n6559), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6558) );
  OAI21_X1 U8111 ( .B1(n6559), .B2(P2_REG1_REG_4__SCAN_IN), .A(n6558), .ZN(
        n6577) );
  NOR2_X1 U8112 ( .A1(n6578), .A2(n6577), .ZN(n6576) );
  AOI21_X1 U8113 ( .B1(n6559), .B2(P2_REG1_REG_4__SCAN_IN), .A(n6576), .ZN(
        n6564) );
  MUX2_X1 U8114 ( .A(n6560), .B(P2_REG1_REG_5__SCAN_IN), .S(n6586), .Z(n6563)
         );
  NOR2_X1 U8115 ( .A1(n6564), .A2(n6563), .ZN(n6587) );
  AND2_X1 U8116 ( .A1(n6565), .A2(n7941), .ZN(n6561) );
  NAND2_X1 U8117 ( .A1(n6562), .A2(n6561), .ZN(n9811) );
  AOI211_X1 U8118 ( .C1(n6564), .C2(n6563), .A(n6587), .B(n9811), .ZN(n6570)
         );
  OAI21_X1 U8119 ( .B1(n9838), .B2(n6941), .A(n6565), .ZN(n6567) );
  NAND2_X1 U8120 ( .A1(n9838), .A2(n7514), .ZN(n6566) );
  AND2_X1 U8121 ( .A1(n6567), .A2(n6566), .ZN(n9813) );
  INV_X1 U8122 ( .A(n9813), .ZN(n8675) );
  INV_X1 U8123 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n6568) );
  NAND2_X1 U8124 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3152), .ZN(n7031) );
  OAI21_X1 U8125 ( .B1(n8675), .B2(n6568), .A(n7031), .ZN(n6569) );
  OR4_X1 U8126 ( .A1(n6572), .A2(n6571), .A3(n6570), .A4(n6569), .ZN(P2_U3250)
         );
  AOI211_X1 U8127 ( .C1(n6575), .C2(n6574), .A(n6573), .B(n8657), .ZN(n6582)
         );
  NOR2_X1 U8128 ( .A1(n9809), .A2(n6612), .ZN(n6581) );
  AOI211_X1 U8129 ( .C1(n6578), .C2(n6577), .A(n6576), .B(n9811), .ZN(n6580)
         );
  INV_X1 U8130 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n10160) );
  NAND2_X1 U8131 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3152), .ZN(n7138) );
  OAI21_X1 U8132 ( .B1(n8675), .B2(n10160), .A(n7138), .ZN(n6579) );
  OR4_X1 U8133 ( .A1(n6582), .A2(n6581), .A3(n6580), .A4(n6579), .ZN(P2_U3249)
         );
  XNOR2_X1 U8134 ( .A(n6807), .B(P2_REG2_REG_6__SCAN_IN), .ZN(n6584) );
  AOI211_X1 U8135 ( .C1(n6585), .C2(n6584), .A(n6806), .B(n8657), .ZN(n6599)
         );
  INV_X1 U8136 ( .A(n6807), .ZN(n6627) );
  NOR2_X1 U8137 ( .A1(n9809), .A2(n6627), .ZN(n6598) );
  NAND2_X1 U8138 ( .A1(n6586), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6589) );
  INV_X1 U8139 ( .A(n6587), .ZN(n6588) );
  NAND2_X1 U8140 ( .A1(n6589), .A2(n6588), .ZN(n6591) );
  INV_X1 U8141 ( .A(n6591), .ZN(n6594) );
  XNOR2_X1 U8142 ( .A(n6807), .B(n6590), .ZN(n6592) );
  INV_X1 U8143 ( .A(n6592), .ZN(n6593) );
  AND2_X1 U8144 ( .A1(n6592), .A2(n6591), .ZN(n6800) );
  AOI211_X1 U8145 ( .C1(n6594), .C2(n6593), .A(n6800), .B(n9811), .ZN(n6597)
         );
  INV_X1 U8146 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n6595) );
  NAND2_X1 U8147 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3152), .ZN(n7063) );
  OAI21_X1 U8148 ( .B1(n8675), .B2(n6595), .A(n7063), .ZN(n6596) );
  OR4_X1 U8149 ( .A1(n6599), .A2(n6598), .A3(n6597), .A4(n6596), .ZN(P2_U3251)
         );
  INV_X1 U8150 ( .A(n6600), .ZN(n6602) );
  OAI21_X1 U8151 ( .B1(n6602), .B2(P1_STATE_REG_SCAN_IN), .A(n6601), .ZN(
        P1_U3353) );
  AND2_X1 U8152 ( .A1(n5601), .A2(P1_U3084), .ZN(n7974) );
  OAI222_X1 U8153 ( .A1(n8557), .A2(n6604), .B1(n4370), .B2(n6615), .C1(
        P1_U3084), .C2(n6603), .ZN(P1_U3352) );
  OAI222_X1 U8154 ( .A1(n8557), .A2(n6606), .B1(n4370), .B2(n6608), .C1(
        P1_U3084), .C2(n6605), .ZN(P1_U3351) );
  NOR2_X1 U8155 ( .A1(n6607), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8970) );
  INV_X1 U8156 ( .A(n8970), .ZN(n8242) );
  OAI222_X1 U8157 ( .A1(n8242), .A2(n6609), .B1(n8973), .B2(n6608), .C1(
        P2_U3152), .C2(n9487), .ZN(P2_U3356) );
  OAI222_X1 U8158 ( .A1(n8242), .A2(n6610), .B1(n8973), .B2(n6622), .C1(
        P2_U3152), .C2(n6794), .ZN(P2_U3355) );
  OAI222_X1 U8159 ( .A1(n8557), .A2(n6611), .B1(n4370), .B2(n6613), .C1(
        P1_U3084), .C2(n9612), .ZN(P1_U3349) );
  OAI222_X1 U8160 ( .A1(n8242), .A2(n6614), .B1(n8973), .B2(n6613), .C1(
        P2_U3152), .C2(n6612), .ZN(P2_U3354) );
  INV_X1 U8161 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6616) );
  OAI222_X1 U8162 ( .A1(n8242), .A2(n6616), .B1(n8973), .B2(n6615), .C1(
        P2_U3152), .C2(n9473), .ZN(P2_U3357) );
  OAI222_X1 U8163 ( .A1(n8557), .A2(n6618), .B1(n4370), .B2(n6620), .C1(
        P1_U3084), .C2(n6617), .ZN(P1_U3348) );
  OAI222_X1 U8164 ( .A1(n8242), .A2(n6621), .B1(n8973), .B2(n6620), .C1(
        P2_U3152), .C2(n6619), .ZN(P2_U3353) );
  OAI222_X1 U8165 ( .A1(n8557), .A2(n9978), .B1(n4370), .B2(n6622), .C1(
        P1_U3084), .C2(n6710), .ZN(P1_U3350) );
  NAND2_X1 U8166 ( .A1(n6829), .A2(n9755), .ZN(n6623) );
  OAI21_X1 U8167 ( .B1(n9755), .B2(n6624), .A(n6623), .ZN(P1_U3440) );
  INV_X1 U8168 ( .A(n6625), .ZN(n6628) );
  INV_X1 U8169 ( .A(n8557), .ZN(n9459) );
  AOI22_X1 U8170 ( .A1(n9652), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n9459), .ZN(n6626) );
  OAI21_X1 U8171 ( .B1(n6628), .B2(n4370), .A(n6626), .ZN(P1_U3347) );
  INV_X1 U8172 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n10147) );
  OAI222_X1 U8173 ( .A1(n8242), .A2(n10147), .B1(n8973), .B2(n6628), .C1(
        P2_U3152), .C2(n6627), .ZN(P2_U3352) );
  INV_X1 U8174 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n10122) );
  INV_X1 U8175 ( .A(n6629), .ZN(n6631) );
  INV_X1 U8176 ( .A(n6821), .ZN(n6630) );
  OAI222_X1 U8177 ( .A1(n8242), .A2(n10122), .B1(n8973), .B2(n6631), .C1(
        P2_U3152), .C2(n6630), .ZN(P2_U3351) );
  INV_X1 U8178 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6632) );
  INV_X1 U8179 ( .A(n6719), .ZN(n6740) );
  OAI222_X1 U8180 ( .A1(n8557), .A2(n6632), .B1(n4370), .B2(n6631), .C1(
        P1_U3084), .C2(n6740), .ZN(P1_U3346) );
  INV_X1 U8181 ( .A(n6633), .ZN(n6635) );
  INV_X1 U8182 ( .A(n6864), .ZN(n6634) );
  OAI222_X1 U8183 ( .A1(n8242), .A2(n10073), .B1(n8973), .B2(n6635), .C1(
        P2_U3152), .C2(n6634), .ZN(P2_U3350) );
  INV_X1 U8184 ( .A(n6708), .ZN(n6751) );
  OAI222_X1 U8185 ( .A1(n8557), .A2(n10181), .B1(n4370), .B2(n6635), .C1(
        P1_U3084), .C2(n6751), .ZN(P1_U3345) );
  INV_X1 U8186 ( .A(n6636), .ZN(n6641) );
  AOI22_X1 U8187 ( .A1(n9667), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n9459), .ZN(n6637) );
  OAI21_X1 U8188 ( .B1(n6641), .B2(n4370), .A(n6637), .ZN(P1_U3344) );
  NAND2_X1 U8189 ( .A1(n6638), .A2(P1_U4006), .ZN(n6639) );
  OAI21_X1 U8190 ( .B1(P1_U4006), .B2(n5845), .A(n6639), .ZN(P1_U3555) );
  INV_X1 U8191 ( .A(n6921), .ZN(n6640) );
  OAI222_X1 U8192 ( .A1(n8242), .A2(n10082), .B1(n8973), .B2(n6641), .C1(n6640), .C2(P2_U3152), .ZN(P2_U3349) );
  INV_X1 U8193 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6647) );
  NAND2_X1 U8194 ( .A1(n8287), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6645) );
  NAND2_X1 U8195 ( .A1(n8288), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6644) );
  NAND2_X1 U8196 ( .A1(n6642), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6643) );
  NAND3_X1 U8197 ( .A1(n6645), .A2(n6644), .A3(n6643), .ZN(n8394) );
  NAND2_X1 U8198 ( .A1(n8394), .A2(P1_U4006), .ZN(n6646) );
  OAI21_X1 U8199 ( .B1(P1_U4006), .B2(n6647), .A(n6646), .ZN(P1_U3586) );
  INV_X1 U8200 ( .A(n6648), .ZN(n6649) );
  INV_X1 U8201 ( .A(n6849), .ZN(n6722) );
  OAI222_X1 U8202 ( .A1(n8557), .A2(n10148), .B1(n4370), .B2(n6649), .C1(
        P1_U3084), .C2(n6722), .ZN(P1_U3343) );
  INV_X1 U8203 ( .A(n7113), .ZN(n6930) );
  OAI222_X1 U8204 ( .A1(n8242), .A2(n6650), .B1(n8973), .B2(n6649), .C1(
        P2_U3152), .C2(n6930), .ZN(P2_U3348) );
  INV_X1 U8205 ( .A(n6651), .ZN(n6652) );
  INV_X1 U8206 ( .A(n9672), .ZN(n6847) );
  OAI222_X1 U8207 ( .A1(n4370), .A2(n6652), .B1(n6847), .B2(P1_U3084), .C1(
        n10150), .C2(n8557), .ZN(P1_U3342) );
  INV_X1 U8208 ( .A(n7454), .ZN(n7119) );
  OAI222_X1 U8209 ( .A1(n8242), .A2(n10222), .B1(n8973), .B2(n6652), .C1(n7119), .C2(P2_U3152), .ZN(P2_U3347) );
  INV_X1 U8210 ( .A(n6653), .ZN(n6655) );
  AOI22_X1 U8211 ( .A1(n7403), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n9459), .ZN(n6654) );
  OAI21_X1 U8212 ( .B1(n6655), .B2(n4370), .A(n6654), .ZN(P1_U3340) );
  INV_X1 U8213 ( .A(n7684), .ZN(n7530) );
  OAI222_X1 U8214 ( .A1(n8242), .A2(n10216), .B1(n8973), .B2(n6655), .C1(
        P2_U3152), .C2(n7530), .ZN(P2_U3345) );
  INV_X1 U8215 ( .A(n6656), .ZN(n6658) );
  INV_X1 U8216 ( .A(n7773), .ZN(n7766) );
  OAI222_X1 U8217 ( .A1(n4370), .A2(n6658), .B1(n7766), .B2(P1_U3084), .C1(
        n6657), .C2(n8557), .ZN(P1_U3339) );
  NOR2_X1 U8218 ( .A1(n9813), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U8219 ( .A(n7872), .ZN(n7692) );
  OAI222_X1 U8220 ( .A1(n8242), .A2(n6659), .B1(n8973), .B2(n6658), .C1(n7692), 
        .C2(P2_U3152), .ZN(P2_U3344) );
  INV_X1 U8221 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n6671) );
  OAI21_X1 U8222 ( .B1(n6662), .B2(n6661), .A(n6660), .ZN(n6663) );
  INV_X1 U8223 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n9707) );
  OAI22_X1 U8224 ( .A1(n9636), .A2(n6663), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9707), .ZN(n6664) );
  AOI21_X1 U8225 ( .B1(n9686), .B2(n6665), .A(n6664), .ZN(n6670) );
  INV_X1 U8226 ( .A(n9659), .ZN(n9695) );
  OAI211_X1 U8227 ( .C1(n6668), .C2(n6667), .A(n9695), .B(n6666), .ZN(n6669)
         );
  OAI211_X1 U8228 ( .C1(n6671), .C2(n9699), .A(n6670), .B(n6669), .ZN(P1_U3242) );
  INV_X1 U8229 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n6687) );
  XNOR2_X1 U8230 ( .A(n6710), .B(P1_REG2_REG_3__SCAN_IN), .ZN(n6675) );
  NAND2_X1 U8231 ( .A1(n6676), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6672) );
  NAND2_X1 U8232 ( .A1(n6673), .A2(n6672), .ZN(n6674) );
  NAND2_X1 U8233 ( .A1(n6674), .A2(n6675), .ZN(n6697) );
  OAI211_X1 U8234 ( .C1(n6675), .C2(n6674), .A(n9695), .B(n6697), .ZN(n6686)
         );
  INV_X1 U8235 ( .A(n6710), .ZN(n6695) );
  INV_X1 U8236 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n10089) );
  MUX2_X1 U8237 ( .A(n10089), .B(P1_REG1_REG_3__SCAN_IN), .S(n6710), .Z(n6680)
         );
  NAND2_X1 U8238 ( .A1(n6676), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6677) );
  NAND2_X1 U8239 ( .A1(n6678), .A2(n6677), .ZN(n6679) );
  AND2_X1 U8240 ( .A1(n6680), .A2(n6679), .ZN(n9616) );
  INV_X1 U8241 ( .A(n9616), .ZN(n6713) );
  OAI21_X1 U8242 ( .B1(n6680), .B2(n6679), .A(n6713), .ZN(n6683) );
  NOR2_X1 U8243 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6681), .ZN(n6880) );
  INV_X1 U8244 ( .A(n6880), .ZN(n6682) );
  OAI21_X1 U8245 ( .B1(n9636), .B2(n6683), .A(n6682), .ZN(n6684) );
  AOI21_X1 U8246 ( .B1(n9686), .B2(n6695), .A(n6684), .ZN(n6685) );
  OAI211_X1 U8247 ( .C1(n6687), .C2(n9699), .A(n6686), .B(n6685), .ZN(P1_U3244) );
  INV_X1 U8248 ( .A(n6688), .ZN(n6690) );
  INV_X1 U8249 ( .A(n7518), .ZN(n7522) );
  OAI222_X1 U8250 ( .A1(n8242), .A2(n6689), .B1(n8973), .B2(n6690), .C1(
        P2_U3152), .C2(n7522), .ZN(P2_U3346) );
  INV_X1 U8251 ( .A(n6974), .ZN(n6845) );
  OAI222_X1 U8252 ( .A1(n8557), .A2(n6691), .B1(n4370), .B2(n6690), .C1(
        P1_U3084), .C2(n6845), .ZN(P1_U3341) );
  INV_X1 U8253 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n6728) );
  NOR2_X1 U8254 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6692), .ZN(n7716) );
  INV_X1 U8255 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n7426) );
  XNOR2_X1 U8256 ( .A(n6708), .B(n7426), .ZN(n6745) );
  AOI22_X1 U8257 ( .A1(P1_REG2_REG_7__SCAN_IN), .A2(n6719), .B1(n6740), .B2(
        n7290), .ZN(n6733) );
  INV_X1 U8258 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6693) );
  XNOR2_X1 U8259 ( .A(n9652), .B(n6693), .ZN(n9643) );
  OR2_X1 U8260 ( .A1(n9639), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6699) );
  NOR2_X1 U8261 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n9639), .ZN(n6694) );
  AOI21_X1 U8262 ( .B1(n9639), .B2(P1_REG2_REG_5__SCAN_IN), .A(n6694), .ZN(
        n9628) );
  NAND2_X1 U8263 ( .A1(n6695), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6696) );
  NAND2_X1 U8264 ( .A1(n6697), .A2(n6696), .ZN(n9607) );
  INV_X1 U8265 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n10157) );
  MUX2_X1 U8266 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n10157), .S(n9612), .Z(n9608)
         );
  NAND2_X1 U8267 ( .A1(n9612), .A2(n10157), .ZN(n6698) );
  NAND2_X1 U8268 ( .A1(n9609), .A2(n6698), .ZN(n9627) );
  NAND2_X1 U8269 ( .A1(n6733), .A2(n6734), .ZN(n6732) );
  OAI21_X1 U8270 ( .B1(P1_REG2_REG_7__SCAN_IN), .B2(n6719), .A(n6732), .ZN(
        n6746) );
  NOR2_X1 U8271 ( .A1(n6708), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6700) );
  AOI21_X1 U8272 ( .B1(n6745), .B2(n6746), .A(n6700), .ZN(n9656) );
  OR2_X1 U8273 ( .A1(n9667), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6702) );
  NAND2_X1 U8274 ( .A1(P1_REG2_REG_9__SCAN_IN), .A2(n9667), .ZN(n6701) );
  AND2_X1 U8275 ( .A1(n6702), .A2(n6701), .ZN(n9655) );
  NAND2_X1 U8276 ( .A1(n6849), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6703) );
  OAI21_X1 U8277 ( .B1(n6849), .B2(P1_REG2_REG_10__SCAN_IN), .A(n6703), .ZN(
        n6704) );
  AOI211_X1 U8278 ( .C1(n6705), .C2(n6704), .A(n6848), .B(n9659), .ZN(n6706)
         );
  AOI211_X1 U8279 ( .C1(n9686), .C2(n6849), .A(n7716), .B(n6706), .ZN(n6727)
         );
  NOR2_X1 U8280 ( .A1(P1_REG1_REG_9__SCAN_IN), .A2(n9667), .ZN(n6707) );
  AOI21_X1 U8281 ( .B1(n9667), .B2(P1_REG1_REG_9__SCAN_IN), .A(n6707), .ZN(
        n9662) );
  INV_X1 U8282 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6720) );
  MUX2_X1 U8283 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n6720), .S(n6708), .Z(n6748)
         );
  NOR2_X1 U8284 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(n6719), .ZN(n6709) );
  AOI21_X1 U8285 ( .B1(n6719), .B2(P1_REG1_REG_7__SCAN_IN), .A(n6709), .ZN(
        n6737) );
  XNOR2_X1 U8286 ( .A(n9652), .B(P1_REG1_REG_6__SCAN_IN), .ZN(n9647) );
  XNOR2_X1 U8287 ( .A(n9612), .B(P1_REG1_REG_4__SCAN_IN), .ZN(n9618) );
  NOR2_X1 U8288 ( .A1(n6710), .A2(n10089), .ZN(n9615) );
  INV_X1 U8289 ( .A(n9615), .ZN(n6711) );
  AND2_X1 U8290 ( .A1(n9618), .A2(n6711), .ZN(n6712) );
  NAND2_X1 U8291 ( .A1(n6713), .A2(n6712), .ZN(n9617) );
  INV_X1 U8292 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6714) );
  NAND2_X1 U8293 ( .A1(n9612), .A2(n6714), .ZN(n6715) );
  NAND2_X1 U8294 ( .A1(n9617), .A2(n6715), .ZN(n9630) );
  OR2_X1 U8295 ( .A1(n9639), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6717) );
  NAND2_X1 U8296 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(n9639), .ZN(n6716) );
  NAND2_X1 U8297 ( .A1(n6717), .A2(n6716), .ZN(n9629) );
  NOR2_X1 U8298 ( .A1(n9630), .A2(n9629), .ZN(n9632) );
  AOI21_X1 U8299 ( .B1(n9639), .B2(P1_REG1_REG_5__SCAN_IN), .A(n9632), .ZN(
        n6718) );
  INV_X1 U8300 ( .A(n6718), .ZN(n9646) );
  OAI22_X1 U8301 ( .A1(n9647), .A2(n9646), .B1(n9652), .B2(
        P1_REG1_REG_6__SCAN_IN), .ZN(n6736) );
  NAND2_X1 U8302 ( .A1(n6737), .A2(n6736), .ZN(n6735) );
  OAI21_X1 U8303 ( .B1(P1_REG1_REG_7__SCAN_IN), .B2(n6719), .A(n6735), .ZN(
        n6749) );
  NAND2_X1 U8304 ( .A1(n6748), .A2(n6749), .ZN(n6747) );
  NAND2_X1 U8305 ( .A1(n6751), .A2(n6720), .ZN(n6721) );
  NAND2_X1 U8306 ( .A1(n6747), .A2(n6721), .ZN(n9661) );
  NAND2_X1 U8307 ( .A1(n9662), .A2(n9661), .ZN(n9660) );
  OAI21_X1 U8308 ( .B1(P1_REG1_REG_9__SCAN_IN), .B2(n9667), .A(n9660), .ZN(
        n6724) );
  INV_X1 U8309 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n9519) );
  AOI22_X1 U8310 ( .A1(n6849), .A2(P1_REG1_REG_10__SCAN_IN), .B1(n9519), .B2(
        n6722), .ZN(n6723) );
  NAND2_X1 U8311 ( .A1(n6723), .A2(n6724), .ZN(n6838) );
  OAI21_X1 U8312 ( .B1(n6724), .B2(n6723), .A(n6838), .ZN(n6725) );
  NAND2_X1 U8313 ( .A1(n6725), .A2(n9694), .ZN(n6726) );
  OAI211_X1 U8314 ( .C1(n9699), .C2(n6728), .A(n6727), .B(n6726), .ZN(P1_U3251) );
  INV_X1 U8315 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n6730) );
  NAND2_X1 U8316 ( .A1(P2_U3966), .A2(n8681), .ZN(n6729) );
  OAI21_X1 U8317 ( .B1(P2_U3966), .B2(n6730), .A(n6729), .ZN(P2_U3583) );
  NAND2_X1 U8318 ( .A1(P2_U3966), .A2(n6419), .ZN(n6731) );
  OAI21_X1 U8319 ( .B1(P2_U3966), .B2(n4970), .A(n6731), .ZN(P2_U3552) );
  INV_X1 U8320 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n6744) );
  OAI21_X1 U8321 ( .B1(n6734), .B2(n6733), .A(n6732), .ZN(n6742) );
  INV_X1 U8322 ( .A(n9686), .ZN(n7900) );
  OAI21_X1 U8323 ( .B1(n6737), .B2(n6736), .A(n6735), .ZN(n6738) );
  AND2_X1 U8324 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7244) );
  AOI21_X1 U8325 ( .B1(n9694), .B2(n6738), .A(n7244), .ZN(n6739) );
  OAI21_X1 U8326 ( .B1(n7900), .B2(n6740), .A(n6739), .ZN(n6741) );
  AOI21_X1 U8327 ( .B1(n9695), .B2(n6742), .A(n6741), .ZN(n6743) );
  OAI21_X1 U8328 ( .B1(n9699), .B2(n6744), .A(n6743), .ZN(P1_U3248) );
  XOR2_X1 U8329 ( .A(n6746), .B(n6745), .Z(n6756) );
  OAI21_X1 U8330 ( .B1(n6749), .B2(n6748), .A(n6747), .ZN(n6753) );
  NOR2_X1 U8331 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6750), .ZN(n7594) );
  NOR2_X1 U8332 ( .A1(n7900), .A2(n6751), .ZN(n6752) );
  AOI211_X1 U8333 ( .C1(n9694), .C2(n6753), .A(n7594), .B(n6752), .ZN(n6755)
         );
  INV_X1 U8334 ( .A(n9699), .ZN(n9668) );
  NAND2_X1 U8335 ( .A1(n9668), .A2(P1_ADDR_REG_8__SCAN_IN), .ZN(n6754) );
  OAI211_X1 U8336 ( .C1(n6756), .C2(n9659), .A(n6755), .B(n6754), .ZN(P1_U3249) );
  INV_X1 U8337 ( .A(n6757), .ZN(n6759) );
  INV_X1 U8338 ( .A(n7874), .ZN(n8087) );
  OAI222_X1 U8339 ( .A1(n8242), .A2(n6758), .B1(n8973), .B2(n6759), .C1(
        P2_U3152), .C2(n8087), .ZN(P2_U3343) );
  OAI222_X1 U8340 ( .A1(n8557), .A2(n6760), .B1(n4370), .B2(n6759), .C1(
        P1_U3084), .C2(n7890), .ZN(P1_U3338) );
  INV_X1 U8341 ( .A(n6761), .ZN(n6772) );
  INV_X1 U8342 ( .A(n8103), .ZN(n7899) );
  OAI222_X1 U8343 ( .A1(n4370), .A2(n6772), .B1(n7899), .B2(P1_U3084), .C1(
        n6762), .C2(n8557), .ZN(P1_U3337) );
  INV_X1 U8344 ( .A(n7044), .ZN(n6766) );
  AND2_X1 U8345 ( .A1(n6638), .A2(n8214), .ZN(n9701) );
  INV_X1 U8346 ( .A(n9701), .ZN(n6763) );
  OAI21_X1 U8347 ( .B1(n8214), .B2(n6638), .A(n6763), .ZN(n8473) );
  NAND2_X1 U8348 ( .A1(n7161), .A2(n7044), .ZN(n6765) );
  INV_X1 U8349 ( .A(n5011), .ZN(n6902) );
  OR2_X1 U8350 ( .A1(n8508), .A2(n6764), .ZN(n9348) );
  OAI22_X1 U8351 ( .A1(n8473), .A2(n6765), .B1(n6902), .B2(n9348), .ZN(n7055)
         );
  AOI21_X1 U8352 ( .B1(n8214), .B2(n6766), .A(n7055), .ZN(n6836) );
  OR2_X1 U8353 ( .A1(n6886), .A2(n8514), .ZN(n6767) );
  AND2_X1 U8354 ( .A1(n6767), .A2(n7038), .ZN(n6834) );
  NAND2_X1 U8355 ( .A1(n6768), .A2(n9755), .ZN(n6833) );
  NOR2_X1 U8356 ( .A1(n6833), .A2(n6769), .ZN(n6770) );
  AND2_X2 U8357 ( .A1(n6834), .A2(n6770), .ZN(n9806) );
  NAND2_X1 U8358 ( .A1(n9803), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6771) );
  OAI21_X1 U8359 ( .B1(n6836), .B2(n9803), .A(n6771), .ZN(P1_U3523) );
  OAI222_X1 U8360 ( .A1(n8242), .A2(n6773), .B1(n8973), .B2(n6772), .C1(n8221), 
        .C2(P2_U3152), .ZN(P2_U3342) );
  INV_X1 U8361 ( .A(n8207), .ZN(n6776) );
  AOI21_X1 U8362 ( .B1(n6777), .B2(n6774), .A(n6776), .ZN(n6783) );
  AOI22_X1 U8363 ( .A1(n9068), .A2(n6638), .B1(n6901), .B2(n9073), .ZN(n6782)
         );
  INV_X1 U8364 ( .A(n6833), .ZN(n6779) );
  NAND3_X1 U8365 ( .A1(n6780), .A2(n6779), .A3(n6778), .ZN(n8213) );
  AOI22_X1 U8366 ( .A1(n9067), .A2(n9712), .B1(n8213), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n6781) );
  OAI211_X1 U8367 ( .C1(n6783), .C2(n9075), .A(n6782), .B(n6781), .ZN(P1_U3220) );
  AOI211_X1 U8368 ( .C1(n6786), .C2(n6785), .A(n6784), .B(n8657), .ZN(n6796)
         );
  AND2_X1 U8369 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_U3152), .ZN(n6787) );
  AOI21_X1 U8370 ( .B1(n9813), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n6787), .ZN(
        n6793) );
  INV_X1 U8371 ( .A(n9811), .ZN(n9807) );
  AOI21_X1 U8372 ( .B1(n6790), .B2(n6789), .A(n6788), .ZN(n6791) );
  NAND2_X1 U8373 ( .A1(n9807), .A2(n6791), .ZN(n6792) );
  OAI211_X1 U8374 ( .C1(n9809), .C2(n6794), .A(n6793), .B(n6792), .ZN(n6795)
         );
  OR2_X1 U8375 ( .A1(n6796), .A2(n6795), .ZN(P2_U3248) );
  INV_X1 U8376 ( .A(n6797), .ZN(n6828) );
  AOI22_X1 U8377 ( .A1(n9095), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n9459), .ZN(n6798) );
  OAI21_X1 U8378 ( .B1(n6828), .B2(n4370), .A(n6798), .ZN(P1_U3336) );
  INV_X1 U8379 ( .A(n9809), .ZN(n6870) );
  MUX2_X1 U8380 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n5920), .S(n6821), .Z(n6802)
         );
  AND2_X1 U8381 ( .A1(n6807), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6799) );
  NAND2_X1 U8382 ( .A1(n6801), .A2(n6802), .ZN(n6815) );
  OAI21_X1 U8383 ( .B1(n6802), .B2(n6801), .A(n6815), .ZN(n6805) );
  NAND2_X1 U8384 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_U3152), .ZN(n6804) );
  NAND2_X1 U8385 ( .A1(n9813), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n6803) );
  OAI211_X1 U8386 ( .C1(n9811), .C2(n6805), .A(n6804), .B(n6803), .ZN(n6812)
         );
  NAND2_X1 U8387 ( .A1(n6821), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6808) );
  OAI21_X1 U8388 ( .B1(n6821), .B2(P2_REG2_REG_7__SCAN_IN), .A(n6808), .ZN(
        n6809) );
  AOI211_X1 U8389 ( .C1(n6810), .C2(n6809), .A(n6820), .B(n8657), .ZN(n6811)
         );
  AOI211_X1 U8390 ( .C1(n6870), .C2(n6821), .A(n6812), .B(n6811), .ZN(n6813)
         );
  INV_X1 U8391 ( .A(n6813), .ZN(P2_U3252) );
  INV_X1 U8392 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n6819) );
  MUX2_X1 U8393 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n5929), .S(n6864), .Z(n6817)
         );
  NAND2_X1 U8394 ( .A1(n6821), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6814) );
  NAND2_X1 U8395 ( .A1(n6815), .A2(n6814), .ZN(n6816) );
  NAND2_X1 U8396 ( .A1(n6816), .A2(n6817), .ZN(n6858) );
  OAI211_X1 U8397 ( .C1(n6817), .C2(n6816), .A(n9807), .B(n6858), .ZN(n6818)
         );
  NAND2_X1 U8398 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3152), .ZN(n7073) );
  OAI211_X1 U8399 ( .C1(n6819), .C2(n8675), .A(n6818), .B(n7073), .ZN(n6826)
         );
  MUX2_X1 U8400 ( .A(n6822), .B(P2_REG2_REG_8__SCAN_IN), .S(n6864), .Z(n6823)
         );
  NOR2_X1 U8401 ( .A1(n6823), .A2(n6824), .ZN(n6863) );
  AOI211_X1 U8402 ( .C1(n6824), .C2(n6823), .A(n6863), .B(n8657), .ZN(n6825)
         );
  AOI211_X1 U8403 ( .C1(n6870), .C2(n6864), .A(n6826), .B(n6825), .ZN(n6827)
         );
  INV_X1 U8404 ( .A(n6827), .ZN(P2_U3253) );
  INV_X1 U8405 ( .A(n8229), .ZN(n8668) );
  OAI222_X1 U8406 ( .A1(n8242), .A2(n10113), .B1(n8973), .B2(n6828), .C1(n8668), .C2(P2_U3152), .ZN(P2_U3341) );
  INV_X1 U8407 ( .A(n6829), .ZN(n6831) );
  NAND2_X1 U8408 ( .A1(n6831), .A2(n6830), .ZN(n6832) );
  NOR2_X1 U8409 ( .A1(n6833), .A2(n6832), .ZN(n7039) );
  AND2_X2 U8410 ( .A1(n7039), .A2(n6834), .ZN(n9795) );
  INV_X1 U8411 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n10132) );
  NAND2_X1 U8412 ( .A1(n9794), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n6835) );
  OAI21_X1 U8413 ( .B1(n6836), .B2(n9794), .A(n6835), .ZN(P1_U3454) );
  INV_X1 U8414 ( .A(n8613), .ZN(n8766) );
  NAND2_X1 U8415 ( .A1(n8766), .A2(P2_U3966), .ZN(n6837) );
  OAI21_X1 U8416 ( .B1(P2_U3966), .B2(n5609), .A(n6837), .ZN(P2_U3575) );
  INV_X1 U8417 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n9588) );
  AOI22_X1 U8418 ( .A1(P1_REG1_REG_11__SCAN_IN), .A2(n9672), .B1(n6847), .B2(
        n9588), .ZN(n9677) );
  OAI21_X1 U8419 ( .B1(n6849), .B2(P1_REG1_REG_10__SCAN_IN), .A(n6838), .ZN(
        n9676) );
  NAND2_X1 U8420 ( .A1(n9677), .A2(n9676), .ZN(n9675) );
  OAI21_X1 U8421 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(n9672), .A(n9675), .ZN(
        n6841) );
  INV_X1 U8422 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n6839) );
  MUX2_X1 U8423 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n6839), .S(n6974), .Z(n6840)
         );
  NAND2_X1 U8424 ( .A1(n6840), .A2(n6841), .ZN(n6967) );
  OAI21_X1 U8425 ( .B1(n6841), .B2(n6840), .A(n6967), .ZN(n6855) );
  NAND2_X1 U8426 ( .A1(n9668), .A2(P1_ADDR_REG_12__SCAN_IN), .ZN(n6844) );
  NOR2_X1 U8427 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6842), .ZN(n7861) );
  INV_X1 U8428 ( .A(n7861), .ZN(n6843) );
  OAI211_X1 U8429 ( .C1(n7900), .C2(n6845), .A(n6844), .B(n6843), .ZN(n6854)
         );
  INV_X1 U8430 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n6846) );
  AOI22_X1 U8431 ( .A1(P1_REG2_REG_11__SCAN_IN), .A2(n9672), .B1(n6847), .B2(
        n6846), .ZN(n9674) );
  NAND2_X1 U8432 ( .A1(n9674), .A2(n4403), .ZN(n9673) );
  OAI21_X1 U8433 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n9672), .A(n9673), .ZN(
        n6852) );
  NAND2_X1 U8434 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n6974), .ZN(n6850) );
  OAI21_X1 U8435 ( .B1(n6974), .B2(P1_REG2_REG_12__SCAN_IN), .A(n6850), .ZN(
        n6851) );
  NOR2_X1 U8436 ( .A1(n6851), .A2(n6852), .ZN(n6973) );
  AOI211_X1 U8437 ( .C1(n6852), .C2(n6851), .A(n6973), .B(n9659), .ZN(n6853)
         );
  AOI211_X1 U8438 ( .C1(n9694), .C2(n6855), .A(n6854), .B(n6853), .ZN(n6856)
         );
  INV_X1 U8439 ( .A(n6856), .ZN(P1_U3253) );
  INV_X1 U8440 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n6862) );
  INV_X1 U8441 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n7652) );
  MUX2_X1 U8442 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n7652), .S(n6921), .Z(n6860)
         );
  NAND2_X1 U8443 ( .A1(n6864), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n6857) );
  NAND2_X1 U8444 ( .A1(n6858), .A2(n6857), .ZN(n6859) );
  NAND2_X1 U8445 ( .A1(n6859), .A2(n6860), .ZN(n6923) );
  OAI211_X1 U8446 ( .C1(n6860), .C2(n6859), .A(n9807), .B(n6923), .ZN(n6861)
         );
  NAND2_X1 U8447 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3152), .ZN(n7374) );
  OAI211_X1 U8448 ( .C1(n6862), .C2(n8675), .A(n6861), .B(n7374), .ZN(n6869)
         );
  NAND2_X1 U8449 ( .A1(n6921), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6865) );
  OAI21_X1 U8450 ( .B1(n6921), .B2(P2_REG2_REG_9__SCAN_IN), .A(n6865), .ZN(
        n6866) );
  AOI211_X1 U8451 ( .C1(n6867), .C2(n6866), .A(n6917), .B(n8657), .ZN(n6868)
         );
  AOI211_X1 U8452 ( .C1(n6870), .C2(n6921), .A(n6869), .B(n6868), .ZN(n6871)
         );
  INV_X1 U8453 ( .A(n6871), .ZN(P2_U3254) );
  INV_X1 U8454 ( .A(n6872), .ZN(n6885) );
  AOI22_X1 U8455 ( .A1(n8230), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n8970), .ZN(n6873) );
  OAI21_X1 U8456 ( .B1(n6885), .B2(n8973), .A(n6873), .ZN(P2_U3340) );
  INV_X1 U8457 ( .A(n6875), .ZN(n6876) );
  NAND3_X1 U8458 ( .A1(n6874), .A2(n6877), .A3(n6876), .ZN(n6878) );
  AOI21_X1 U8459 ( .B1(n6879), .B2(n6878), .A(n9075), .ZN(n6884) );
  INV_X1 U8460 ( .A(n9049), .ZN(n9071) );
  AOI22_X1 U8461 ( .A1(n9067), .A2(n9087), .B1(n9068), .B2(n9712), .ZN(n6882)
         );
  AOI21_X1 U8462 ( .B1(n9037), .B2(n7049), .A(n6880), .ZN(n6881) );
  OAI211_X1 U8463 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n9071), .A(n6882), .B(
        n6881), .ZN(n6883) );
  OR2_X1 U8464 ( .A1(n6884), .A2(n6883), .ZN(P1_U3216) );
  INV_X1 U8465 ( .A(n9685), .ZN(n9092) );
  OAI222_X1 U8466 ( .A1(n8557), .A2(n10186), .B1(n4370), .B2(n6885), .C1(
        P1_U3084), .C2(n9092), .ZN(P1_U3335) );
  INV_X1 U8467 ( .A(n6886), .ZN(n9793) );
  NAND2_X1 U8468 ( .A1(n9702), .A2(n9701), .ZN(n9700) );
  NAND2_X1 U8469 ( .A1(n5011), .A2(n6901), .ZN(n6887) );
  NAND2_X1 U8470 ( .A1(n9700), .A2(n6887), .ZN(n7382) );
  INV_X1 U8471 ( .A(n7382), .ZN(n6893) );
  AND4_X1 U8472 ( .A1(n6891), .A2(n6890), .A3(n6889), .A4(n6888), .ZN(n6911)
         );
  NAND2_X1 U8473 ( .A1(n6911), .A2(n8209), .ZN(n8518) );
  NAND2_X1 U8474 ( .A1(n9712), .A2(n9762), .ZN(n8519) );
  AND2_X2 U8475 ( .A1(n8518), .A2(n8519), .ZN(n8474) );
  NAND2_X1 U8476 ( .A1(n6893), .A2(n6892), .ZN(n7380) );
  NAND2_X1 U8477 ( .A1(n6911), .A2(n9762), .ZN(n6894) );
  INV_X1 U8478 ( .A(n9088), .ZN(n7154) );
  NAND2_X1 U8479 ( .A1(n7154), .A2(n7049), .ZN(n8522) );
  INV_X1 U8480 ( .A(n7049), .ZN(n7153) );
  NAND2_X1 U8481 ( .A1(n9088), .A2(n7153), .ZN(n8185) );
  NAND2_X1 U8482 ( .A1(n8522), .A2(n8185), .ZN(n6905) );
  NAND2_X1 U8483 ( .A1(n6895), .A2(n6905), .ZN(n7156) );
  OAI21_X1 U8484 ( .B1(n6895), .B2(n6905), .A(n7156), .ZN(n7037) );
  OR2_X1 U8485 ( .A1(n6901), .A2(n8214), .ZN(n9703) );
  NOR2_X1 U8486 ( .A1(n7388), .A2(n7049), .ZN(n8196) );
  INV_X1 U8487 ( .A(n8196), .ZN(n6897) );
  NAND2_X1 U8488 ( .A1(n7388), .A2(n7049), .ZN(n6896) );
  NAND2_X1 U8489 ( .A1(n6897), .A2(n6896), .ZN(n7046) );
  OR2_X1 U8490 ( .A1(n7044), .A2(n6898), .ZN(n9788) );
  OAI22_X1 U8491 ( .A1(n7046), .A2(n9788), .B1(n7153), .B2(n9787), .ZN(n6915)
         );
  OR2_X1 U8492 ( .A1(n5743), .A2(n4989), .ZN(n6900) );
  OR2_X1 U8493 ( .A1(n5744), .A2(n8543), .ZN(n6899) );
  INV_X1 U8494 ( .A(n8214), .ZN(n9705) );
  NOR2_X1 U8495 ( .A1(n6638), .A2(n9705), .ZN(n9715) );
  NAND2_X1 U8496 ( .A1(n6902), .A2(n6901), .ZN(n6903) );
  NAND2_X1 U8497 ( .A1(n8521), .A2(n8474), .ZN(n6904) );
  XNOR2_X1 U8498 ( .A(n7163), .B(n6905), .ZN(n6914) );
  OR2_X1 U8499 ( .A1(n6907), .A2(n6906), .ZN(n6910) );
  OR2_X1 U8500 ( .A1(n6908), .A2(n5744), .ZN(n6909) );
  NAND2_X1 U8501 ( .A1(n6910), .A2(n6909), .ZN(n9502) );
  OR2_X1 U8502 ( .A1(n8508), .A2(n5759), .ZN(n9346) );
  INV_X1 U8503 ( .A(n9087), .ZN(n7236) );
  OAI22_X1 U8504 ( .A1(n6911), .A2(n9346), .B1(n7236), .B2(n9348), .ZN(n6912)
         );
  AOI21_X1 U8505 ( .B1(n7037), .B2(n9502), .A(n6912), .ZN(n6913) );
  OAI21_X1 U8506 ( .B1(n9499), .B2(n6914), .A(n6913), .ZN(n7040) );
  AOI211_X1 U8507 ( .C1(n9793), .C2(n7037), .A(n6915), .B(n7040), .ZN(n6991)
         );
  NAND2_X1 U8508 ( .A1(n9803), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6916) );
  OAI21_X1 U8509 ( .B1(n6991), .B2(n9803), .A(n6916), .ZN(P1_U3526) );
  AOI22_X1 U8510 ( .A1(n7113), .A2(n7617), .B1(P2_REG2_REG_10__SCAN_IN), .B2(
        n6930), .ZN(n6918) );
  AOI211_X1 U8511 ( .C1(n6919), .C2(n6918), .A(n4396), .B(n8657), .ZN(n6932)
         );
  AND2_X1 U8512 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3152), .ZN(n6920) );
  AOI21_X1 U8513 ( .B1(n9813), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n6920), .ZN(
        n6929) );
  NAND2_X1 U8514 ( .A1(n6921), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n6922) );
  AND2_X1 U8515 ( .A1(n6923), .A2(n6922), .ZN(n6926) );
  MUX2_X1 U8516 ( .A(n6924), .B(P2_REG1_REG_10__SCAN_IN), .S(n7113), .Z(n6925)
         );
  NOR2_X1 U8517 ( .A1(n6926), .A2(n6925), .ZN(n7112) );
  AOI21_X1 U8518 ( .B1(n6926), .B2(n6925), .A(n7112), .ZN(n6927) );
  NAND2_X1 U8519 ( .A1(n9807), .A2(n6927), .ZN(n6928) );
  OAI211_X1 U8520 ( .C1(n9809), .C2(n6930), .A(n6929), .B(n6928), .ZN(n6931)
         );
  OR2_X1 U8521 ( .A1(n6932), .A2(n6931), .ZN(P2_U3255) );
  OR2_X1 U8522 ( .A1(n7104), .A2(n6933), .ZN(n7012) );
  NOR2_X1 U8523 ( .A1(n7012), .A2(n9838), .ZN(n6943) );
  INV_X1 U8524 ( .A(n6943), .ZN(n6934) );
  NAND2_X1 U8525 ( .A1(n6934), .A2(n9825), .ZN(n6937) );
  AND2_X1 U8526 ( .A1(n6937), .A2(n7079), .ZN(n6962) );
  INV_X1 U8527 ( .A(n6936), .ZN(n6935) );
  NAND2_X1 U8528 ( .A1(n6943), .A2(n6935), .ZN(n8627) );
  INV_X1 U8529 ( .A(n8603), .ZN(n8596) );
  INV_X1 U8530 ( .A(n7088), .ZN(n9848) );
  AOI22_X1 U8531 ( .A1(n8596), .A2(n8656), .B1(n8629), .B2(n9847), .ZN(n6946)
         );
  INV_X1 U8532 ( .A(n6938), .ZN(n7193) );
  INV_X1 U8533 ( .A(n6939), .ZN(n6940) );
  MUX2_X1 U8534 ( .A(n9847), .B(n6940), .S(n8274), .Z(n6944) );
  INV_X1 U8535 ( .A(n9882), .ZN(n9899) );
  AND2_X1 U8536 ( .A1(n9899), .A2(n6941), .ZN(n6942) );
  NAND2_X1 U8537 ( .A1(n6943), .A2(n6942), .ZN(n8631) );
  INV_X1 U8538 ( .A(n8631), .ZN(n8611) );
  OAI21_X1 U8539 ( .B1(n7193), .B2(n6944), .A(n8611), .ZN(n6945) );
  OAI211_X1 U8540 ( .C1(n6962), .C2(n7337), .A(n6946), .B(n6945), .ZN(P2_U3234) );
  NAND2_X1 U8541 ( .A1(n6947), .A2(n7171), .ZN(n6949) );
  NAND2_X2 U8542 ( .A1(n6949), .A2(n6948), .ZN(n6957) );
  NAND2_X1 U8543 ( .A1(n6952), .A2(n6953), .ZN(n6955) );
  INV_X1 U8544 ( .A(n6953), .ZN(n6954) );
  INV_X1 U8545 ( .A(n6955), .ZN(n6956) );
  NOR2_X1 U8546 ( .A1(n6980), .A2(n6956), .ZN(n6961) );
  XNOR2_X1 U8547 ( .A(n6957), .B(n9858), .ZN(n6959) );
  NAND2_X1 U8548 ( .A1(n8655), .A2(n8274), .ZN(n6958) );
  NAND2_X1 U8549 ( .A1(n6959), .A2(n6958), .ZN(n6994) );
  OAI21_X1 U8550 ( .B1(n6959), .B2(n6958), .A(n6994), .ZN(n6960) );
  AOI21_X1 U8551 ( .B1(n6961), .B2(n6960), .A(n6996), .ZN(n6965) );
  INV_X1 U8552 ( .A(n6962), .ZN(n6983) );
  AOI22_X1 U8553 ( .A1(n6983), .A2(P2_REG3_REG_2__SCAN_IN), .B1(n8629), .B2(
        n7312), .ZN(n6964) );
  INV_X1 U8554 ( .A(n8602), .ZN(n7150) );
  AOI22_X1 U8555 ( .A1(n7150), .A2(n8656), .B1(n8596), .B2(n8654), .ZN(n6963)
         );
  OAI211_X1 U8556 ( .C1(n6965), .C2(n8631), .A(n6964), .B(n6963), .ZN(P2_U3239) );
  INV_X1 U8557 ( .A(n7403), .ZN(n6972) );
  NAND2_X1 U8558 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n8015) );
  INV_X1 U8559 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n6966) );
  MUX2_X1 U8560 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n6966), .S(n7403), .Z(n6969)
         );
  OAI21_X1 U8561 ( .B1(n6974), .B2(P1_REG1_REG_12__SCAN_IN), .A(n6967), .ZN(
        n6968) );
  NAND2_X1 U8562 ( .A1(n6969), .A2(n6968), .ZN(n7396) );
  OAI21_X1 U8563 ( .B1(n6969), .B2(n6968), .A(n7396), .ZN(n6970) );
  NAND2_X1 U8564 ( .A1(n9694), .A2(n6970), .ZN(n6971) );
  OAI211_X1 U8565 ( .C1(n7900), .C2(n6972), .A(n8015), .B(n6971), .ZN(n6978)
         );
  AOI21_X1 U8566 ( .B1(n6974), .B2(P1_REG2_REG_12__SCAN_IN), .A(n6973), .ZN(
        n6976) );
  XNOR2_X1 U8567 ( .A(n7403), .B(P1_REG2_REG_13__SCAN_IN), .ZN(n6975) );
  NOR2_X1 U8568 ( .A1(n6975), .A2(n6976), .ZN(n7402) );
  AOI211_X1 U8569 ( .C1(n6976), .C2(n6975), .A(n7402), .B(n9659), .ZN(n6977)
         );
  AOI211_X1 U8570 ( .C1(P1_ADDR_REG_13__SCAN_IN), .C2(n9668), .A(n6978), .B(
        n6977), .ZN(n6979) );
  INV_X1 U8571 ( .A(n6979), .ZN(P1_U3254) );
  AOI21_X1 U8572 ( .B1(n6982), .B2(n6981), .A(n6980), .ZN(n6986) );
  AOI22_X1 U8573 ( .A1(n7150), .A2(n6419), .B1(n8596), .B2(n8655), .ZN(n6985)
         );
  AOI22_X1 U8574 ( .A1(n6983), .A2(P2_REG3_REG_1__SCAN_IN), .B1(n8629), .B2(
        n5859), .ZN(n6984) );
  OAI211_X1 U8575 ( .C1(n6986), .C2(n8631), .A(n6985), .B(n6984), .ZN(P2_U3224) );
  INV_X1 U8576 ( .A(n6987), .ZN(n6989) );
  OAI222_X1 U8577 ( .A1(n8557), .A2(n6988), .B1(n4370), .B2(n6989), .C1(
        P1_U3084), .C2(n4989), .ZN(P1_U3334) );
  OAI222_X1 U8578 ( .A1(n8242), .A2(n6990), .B1(n8973), .B2(n6989), .C1(
        P2_U3152), .C2(n9827), .ZN(P2_U3339) );
  INV_X1 U8579 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n6993) );
  OR2_X1 U8580 ( .A1(n6991), .A2(n9794), .ZN(n6992) );
  OAI21_X1 U8581 ( .B1(n9795), .B2(n6993), .A(n6992), .ZN(P1_U3463) );
  INV_X1 U8582 ( .A(n6994), .ZN(n6995) );
  XNOR2_X1 U8583 ( .A(n6957), .B(n7510), .ZN(n6998) );
  NAND2_X1 U8584 ( .A1(n8654), .A2(n8274), .ZN(n6997) );
  XNOR2_X1 U8585 ( .A(n6998), .B(n6997), .ZN(n7144) );
  INV_X1 U8586 ( .A(n6997), .ZN(n6999) );
  AND2_X1 U8587 ( .A1(n8653), .A2(n8274), .ZN(n7001) );
  INV_X1 U8588 ( .A(n9869), .ZN(n7365) );
  XNOR2_X1 U8589 ( .A(n7365), .B(n6957), .ZN(n7000) );
  NOR2_X1 U8590 ( .A1(n7000), .A2(n7001), .ZN(n7002) );
  AOI21_X1 U8591 ( .B1(n7001), .B2(n7000), .A(n7002), .ZN(n7137) );
  INV_X1 U8592 ( .A(n7002), .ZN(n7003) );
  NOR2_X1 U8593 ( .A1(n7211), .A2(n8271), .ZN(n7005) );
  XNOR2_X1 U8594 ( .A(n7101), .B(n6957), .ZN(n7004) );
  NOR2_X1 U8595 ( .A1(n7005), .A2(n7004), .ZN(n7006) );
  AOI21_X1 U8596 ( .B1(n7005), .B2(n7004), .A(n7006), .ZN(n7028) );
  INV_X1 U8597 ( .A(n7006), .ZN(n7007) );
  NAND2_X1 U8598 ( .A1(n7026), .A2(n7007), .ZN(n7060) );
  AND2_X1 U8599 ( .A1(n8651), .A2(n8274), .ZN(n7009) );
  INV_X2 U8600 ( .A(n8247), .ZN(n8276) );
  XNOR2_X1 U8601 ( .A(n7221), .B(n8276), .ZN(n7008) );
  NOR2_X1 U8602 ( .A1(n7008), .A2(n7009), .ZN(n7010) );
  AOI21_X1 U8603 ( .B1(n7009), .B2(n7008), .A(n7010), .ZN(n7061) );
  INV_X1 U8604 ( .A(n7010), .ZN(n7011) );
  XNOR2_X1 U8605 ( .A(n7129), .B(n6957), .ZN(n7069) );
  NOR2_X1 U8606 ( .A1(n7554), .A2(n8271), .ZN(n7070) );
  XNOR2_X1 U8607 ( .A(n7069), .B(n7070), .ZN(n7071) );
  XNOR2_X1 U8608 ( .A(n7072), .B(n7071), .ZN(n7023) );
  NAND2_X1 U8609 ( .A1(n7012), .A2(n7080), .ZN(n7017) );
  INV_X1 U8610 ( .A(n7013), .ZN(n7014) );
  AND3_X1 U8611 ( .A1(n7015), .A2(n7014), .A3(n7079), .ZN(n7016) );
  NAND2_X1 U8612 ( .A1(n7017), .A2(n7016), .ZN(n7018) );
  OAI22_X1 U8613 ( .A1(n8615), .A2(n7461), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7019), .ZN(n7021) );
  OAI22_X1 U8614 ( .A1(n7029), .A2(n8602), .B1(n8603), .B2(n7474), .ZN(n7020)
         );
  AOI211_X1 U8615 ( .C1(n8629), .C2(n7129), .A(n7021), .B(n7020), .ZN(n7022)
         );
  OAI21_X1 U8616 ( .B1(n7023), .B2(n8631), .A(n7022), .ZN(P2_U3215) );
  INV_X1 U8617 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n7025) );
  INV_X1 U8618 ( .A(n9157), .ZN(n9197) );
  NAND2_X1 U8619 ( .A1(n9197), .A2(P1_U4006), .ZN(n7024) );
  OAI21_X1 U8620 ( .B1(P1_U4006), .B2(n7025), .A(n7024), .ZN(P1_U3583) );
  OAI21_X1 U8621 ( .B1(n7028), .B2(n7027), .A(n7026), .ZN(n7034) );
  OAI22_X1 U8622 ( .A1(n7147), .A2(n8602), .B1(n8603), .B2(n7029), .ZN(n7033)
         );
  NAND2_X1 U8623 ( .A1(n8629), .A2(n7101), .ZN(n7030) );
  OAI211_X1 U8624 ( .C1(n8615), .C2(n9824), .A(n7031), .B(n7030), .ZN(n7032)
         );
  AOI211_X1 U8625 ( .C1(n7034), .C2(n8611), .A(n7033), .B(n7032), .ZN(n7035)
         );
  INV_X1 U8626 ( .A(n7035), .ZN(P2_U3229) );
  NAND2_X1 U8627 ( .A1(n8638), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n7036) );
  OAI21_X1 U8628 ( .B1(n8701), .B2(n8638), .A(n7036), .ZN(P2_U3581) );
  INV_X1 U8629 ( .A(n7037), .ZN(n7053) );
  INV_X1 U8630 ( .A(n7038), .ZN(n9752) );
  NAND2_X1 U8631 ( .A1(n7039), .A2(n9752), .ZN(n7286) );
  NOR2_X1 U8632 ( .A1(n4987), .A2(n4989), .ZN(n9724) );
  AND2_X1 U8633 ( .A1(n9725), .A2(n9724), .ZN(n9510) );
  INV_X1 U8634 ( .A(n9510), .ZN(n7052) );
  NAND2_X1 U8635 ( .A1(n7040), .A2(n9725), .ZN(n7051) );
  INV_X1 U8636 ( .A(n9706), .ZN(n7041) );
  INV_X1 U8637 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n7042) );
  OAI22_X1 U8638 ( .A1(n9725), .A2(n7042), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n9708), .ZN(n7048) );
  INV_X1 U8639 ( .A(n7043), .ZN(n8546) );
  NOR2_X1 U8640 ( .A1(n7044), .A2(n8546), .ZN(n7045) );
  NAND2_X1 U8641 ( .A1(n9725), .A2(n7045), .ZN(n9166) );
  NOR2_X1 U8642 ( .A1(n9166), .A2(n7046), .ZN(n7047) );
  AOI211_X1 U8643 ( .C1(n9543), .C2(n7049), .A(n7048), .B(n7047), .ZN(n7050)
         );
  OAI211_X1 U8644 ( .C1(n7053), .C2(n7052), .A(n7051), .B(n7050), .ZN(P1_U3288) );
  INV_X1 U8645 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n8218) );
  NOR2_X1 U8646 ( .A1(n9708), .A2(n8218), .ZN(n7054) );
  OAI21_X1 U8647 ( .B1(n7055), .B2(n7054), .A(n9725), .ZN(n7057) );
  INV_X1 U8648 ( .A(n9166), .ZN(n9366) );
  OAI21_X1 U8649 ( .B1(n9366), .B2(n9543), .A(n8214), .ZN(n7056) );
  OAI211_X1 U8650 ( .C1(n10114), .C2(n9725), .A(n7057), .B(n7056), .ZN(
        P1_U3291) );
  NAND2_X1 U8651 ( .A1(n8638), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n7058) );
  OAI21_X1 U8652 ( .B1(n8714), .B2(n8638), .A(n7058), .ZN(P2_U3578) );
  INV_X1 U8653 ( .A(n7221), .ZN(n9875) );
  INV_X1 U8654 ( .A(n8629), .ZN(n8620) );
  OAI21_X1 U8655 ( .B1(n7061), .B2(n7060), .A(n7059), .ZN(n7062) );
  NAND2_X1 U8656 ( .A1(n7062), .A2(n8611), .ZN(n7068) );
  INV_X1 U8657 ( .A(n7214), .ZN(n7066) );
  INV_X1 U8658 ( .A(n7063), .ZN(n7065) );
  OAI22_X1 U8659 ( .A1(n7211), .A2(n8602), .B1(n8603), .B2(n7554), .ZN(n7064)
         );
  AOI211_X1 U8660 ( .C1(n7066), .C2(n8625), .A(n7065), .B(n7064), .ZN(n7067)
         );
  OAI211_X1 U8661 ( .C1(n9875), .C2(n8620), .A(n7068), .B(n7067), .ZN(P2_U3241) );
  XNOR2_X1 U8662 ( .A(n9881), .B(n8247), .ZN(n7342) );
  NOR2_X1 U8663 ( .A1(n7474), .A2(n8271), .ZN(n7344) );
  XNOR2_X1 U8664 ( .A(n7342), .B(n7344), .ZN(n7345) );
  XNOR2_X1 U8665 ( .A(n7346), .B(n7345), .ZN(n7077) );
  OAI21_X1 U8666 ( .B1(n8615), .B2(n7562), .A(n7073), .ZN(n7075) );
  OAI22_X1 U8667 ( .A1(n7554), .A2(n8602), .B1(n8603), .B2(n7553), .ZN(n7074)
         );
  AOI211_X1 U8668 ( .C1(n8629), .C2(n9881), .A(n7075), .B(n7074), .ZN(n7076)
         );
  OAI21_X1 U8669 ( .B1(n7077), .B2(n8631), .A(n7076), .ZN(P2_U3223) );
  INV_X1 U8670 ( .A(n7078), .ZN(n7081) );
  NAND3_X1 U8671 ( .A1(n7081), .A2(n7080), .A3(n7079), .ZN(n7082) );
  NOR2_X1 U8672 ( .A1(n7082), .A2(n9838), .ZN(n7083) );
  AND2_X1 U8673 ( .A1(n7084), .A2(n7083), .ZN(n7106) );
  AND2_X2 U8674 ( .A1(n7106), .A2(n7104), .ZN(n9909) );
  AND2_X1 U8675 ( .A1(n7747), .A2(n9886), .ZN(n9532) );
  XNOR2_X1 U8676 ( .A(n7085), .B(n7086), .ZN(n9832) );
  OR2_X1 U8677 ( .A1(n7088), .A2(n7087), .ZN(n9901) );
  AOI21_X1 U8678 ( .B1(n7089), .B2(n7101), .A(n9901), .ZN(n7090) );
  AND2_X1 U8679 ( .A1(n7090), .A2(n7216), .ZN(n9828) );
  NAND2_X1 U8680 ( .A1(n7495), .A2(n7091), .ZN(n7357) );
  NAND2_X1 U8681 ( .A1(n7357), .A2(n7092), .ZN(n7097) );
  NAND2_X1 U8682 ( .A1(n7357), .A2(n7093), .ZN(n7095) );
  NAND2_X1 U8683 ( .A1(n7095), .A2(n7094), .ZN(n7096) );
  NAND2_X1 U8684 ( .A1(n7097), .A2(n7096), .ZN(n7098) );
  NAND2_X1 U8685 ( .A1(n7098), .A2(n8843), .ZN(n7100) );
  INV_X1 U8686 ( .A(n8830), .ZN(n8840) );
  AOI22_X1 U8687 ( .A1(n8838), .A2(n8653), .B1(n8651), .B2(n8840), .ZN(n7099)
         );
  NAND2_X1 U8688 ( .A1(n7100), .A2(n7099), .ZN(n9820) );
  AOI211_X1 U8689 ( .C1(n9882), .C2(n7101), .A(n9828), .B(n9820), .ZN(n7102)
         );
  OAI21_X1 U8690 ( .B1(n9532), .B2(n9832), .A(n7102), .ZN(n7107) );
  NAND2_X1 U8691 ( .A1(n7107), .A2(n9909), .ZN(n7103) );
  OAI21_X1 U8692 ( .B1(n9909), .B2(n5871), .A(n7103), .ZN(P2_U3466) );
  INV_X1 U8693 ( .A(n7104), .ZN(n7105) );
  NAND2_X1 U8694 ( .A1(n7106), .A2(n7105), .ZN(n9994) );
  INV_X2 U8695 ( .A(n9994), .ZN(n9996) );
  NAND2_X1 U8696 ( .A1(n7107), .A2(n9996), .ZN(n7108) );
  OAI21_X1 U8697 ( .B1(n9996), .B2(n6560), .A(n7108), .ZN(P2_U3525) );
  AOI22_X1 U8698 ( .A1(n7454), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n7633), .B2(
        n7119), .ZN(n7109) );
  NAND2_X1 U8699 ( .A1(n7110), .A2(n7109), .ZN(n7449) );
  OAI21_X1 U8700 ( .B1(n7110), .B2(n7109), .A(n7449), .ZN(n7121) );
  AOI22_X1 U8701 ( .A1(n9813), .A2(P2_ADDR_REG_11__SCAN_IN), .B1(
        P2_REG3_REG_11__SCAN_IN), .B2(P2_U3152), .ZN(n7118) );
  MUX2_X1 U8702 ( .A(n7111), .B(P2_REG1_REG_11__SCAN_IN), .S(n7454), .Z(n7115)
         );
  AOI21_X1 U8703 ( .B1(n7113), .B2(P2_REG1_REG_10__SCAN_IN), .A(n7112), .ZN(
        n7114) );
  NOR2_X1 U8704 ( .A1(n7114), .A2(n7115), .ZN(n7453) );
  AOI21_X1 U8705 ( .B1(n7115), .B2(n7114), .A(n7453), .ZN(n7116) );
  NAND2_X1 U8706 ( .A1(n9807), .A2(n7116), .ZN(n7117) );
  OAI211_X1 U8707 ( .C1(n9809), .C2(n7119), .A(n7118), .B(n7117), .ZN(n7120)
         );
  AOI21_X1 U8708 ( .B1(n7121), .B2(n9808), .A(n7120), .ZN(n7122) );
  INV_X1 U8709 ( .A(n7122), .ZN(P2_U3256) );
  INV_X1 U8710 ( .A(n7123), .ZN(n7135) );
  OAI222_X1 U8711 ( .A1(n4370), .A2(n7135), .B1(n8543), .B2(P1_U3084), .C1(
        n9998), .C2(n8557), .ZN(P1_U3333) );
  INV_X1 U8712 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n7132) );
  XNOR2_X1 U8713 ( .A(n7124), .B(n7125), .ZN(n7465) );
  XNOR2_X1 U8714 ( .A(n7126), .B(n7125), .ZN(n7127) );
  AOI222_X1 U8715 ( .A1(n8843), .A2(n7127), .B1(n8649), .B2(n8840), .C1(n8651), 
        .C2(n8838), .ZN(n7470) );
  INV_X1 U8716 ( .A(n7217), .ZN(n7128) );
  AOI21_X1 U8717 ( .B1(n7129), .B2(n7128), .A(n7560), .ZN(n7468) );
  INV_X1 U8718 ( .A(n9901), .ZN(n9883) );
  AOI22_X1 U8719 ( .A1(n7468), .A2(n9883), .B1(n9882), .B2(n7129), .ZN(n7130)
         );
  OAI211_X1 U8720 ( .C1(n9532), .C2(n7465), .A(n7470), .B(n7130), .ZN(n7133)
         );
  NAND2_X1 U8721 ( .A1(n7133), .A2(n9909), .ZN(n7131) );
  OAI21_X1 U8722 ( .B1(n9909), .B2(n7132), .A(n7131), .ZN(P2_U3472) );
  NAND2_X1 U8723 ( .A1(n7133), .A2(n9996), .ZN(n7134) );
  OAI21_X1 U8724 ( .B1(n9996), .B2(n5920), .A(n7134), .ZN(P2_U3527) );
  OAI222_X1 U8725 ( .A1(n8242), .A2(n10057), .B1(n8973), .B2(n7135), .C1(n6388), .C2(P2_U3152), .ZN(P2_U3338) );
  OAI21_X1 U8726 ( .B1(n4441), .B2(n7137), .A(n7136), .ZN(n7142) );
  OAI22_X1 U8727 ( .A1(n9869), .A2(n8620), .B1(n8603), .B2(n7211), .ZN(n7141)
         );
  NAND2_X1 U8728 ( .A1(n7150), .A2(n8654), .ZN(n7139) );
  OAI211_X1 U8729 ( .C1(n8615), .C2(n7363), .A(n7139), .B(n7138), .ZN(n7140)
         );
  AOI211_X1 U8730 ( .C1(n7142), .C2(n8611), .A(n7141), .B(n7140), .ZN(n7143)
         );
  INV_X1 U8731 ( .A(n7143), .ZN(P2_U3232) );
  XNOR2_X1 U8732 ( .A(n7145), .B(n7144), .ZN(n7152) );
  INV_X1 U8733 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n7146) );
  OAI22_X1 U8734 ( .A1(n8615), .A2(P2_REG3_REG_3__SCAN_IN), .B1(
        P2_STATE_REG_SCAN_IN), .B2(n7146), .ZN(n7149) );
  OAI22_X1 U8735 ( .A1(n5870), .A2(n8620), .B1(n8603), .B2(n7147), .ZN(n7148)
         );
  AOI211_X1 U8736 ( .C1(n7150), .C2(n8655), .A(n7149), .B(n7148), .ZN(n7151)
         );
  OAI21_X1 U8737 ( .B1(n7152), .B2(n8631), .A(n7151), .ZN(P2_U3220) );
  NAND2_X1 U8738 ( .A1(n7154), .A2(n7153), .ZN(n7155) );
  NAND2_X1 U8739 ( .A1(n7156), .A2(n7155), .ZN(n8190) );
  NAND2_X1 U8740 ( .A1(n7236), .A2(n9022), .ZN(n7280) );
  NAND2_X1 U8741 ( .A1(n7280), .A2(n8426), .ZN(n8189) );
  NAND2_X1 U8742 ( .A1(n8190), .A2(n8189), .ZN(n8191) );
  NAND2_X1 U8743 ( .A1(n7236), .A2(n9767), .ZN(n7157) );
  NAND2_X1 U8744 ( .A1(n8191), .A2(n7157), .ZN(n7420) );
  NAND2_X1 U8745 ( .A1(n7180), .A2(n7251), .ZN(n7279) );
  INV_X1 U8746 ( .A(n7251), .ZN(n7158) );
  NAND2_X1 U8747 ( .A1(n9086), .A2(n7158), .ZN(n8427) );
  AND2_X1 U8748 ( .A1(n7279), .A2(n8427), .ZN(n7292) );
  INV_X1 U8749 ( .A(n7292), .ZN(n7159) );
  OR2_X1 U8750 ( .A1(n7420), .A2(n7292), .ZN(n7174) );
  OAI21_X1 U8751 ( .B1(n4584), .B2(n7159), .A(n7174), .ZN(n7254) );
  AND2_X1 U8752 ( .A1(n7161), .A2(n7160), .ZN(n7162) );
  NAND2_X1 U8753 ( .A1(n9725), .A2(n7162), .ZN(n9368) );
  INV_X1 U8754 ( .A(n9499), .ZN(n9717) );
  INV_X1 U8755 ( .A(n8522), .ZN(n8428) );
  AND2_X1 U8756 ( .A1(n8426), .A2(n8185), .ZN(n8431) );
  NAND2_X1 U8757 ( .A1(n7164), .A2(n7280), .ZN(n7177) );
  XNOR2_X1 U8758 ( .A(n7177), .B(n7292), .ZN(n7165) );
  AOI222_X1 U8759 ( .A1(n9717), .A2(n7165), .B1(n9085), .B2(n9711), .C1(n9087), 
        .C2(n9713), .ZN(n7253) );
  NAND2_X1 U8760 ( .A1(n8196), .A2(n9767), .ZN(n8198) );
  AOI211_X1 U8761 ( .C1(n7251), .C2(n8198), .A(n9788), .B(n4536), .ZN(n7250)
         );
  INV_X1 U8762 ( .A(n9708), .ZN(n9541) );
  AOI22_X1 U8763 ( .A1(n7250), .A2(n4989), .B1(n9541), .B2(n7233), .ZN(n7166)
         );
  INV_X2 U8764 ( .A(n9725), .ZN(n9728) );
  AOI21_X1 U8765 ( .B1(n7253), .B2(n7166), .A(n9728), .ZN(n7167) );
  INV_X1 U8766 ( .A(n7167), .ZN(n7169) );
  AOI22_X1 U8767 ( .A1(n9543), .A2(n7251), .B1(n9728), .B2(
        P1_REG2_REG_5__SCAN_IN), .ZN(n7168) );
  OAI211_X1 U8768 ( .C1(n7254), .C2(n9368), .A(n7169), .B(n7168), .ZN(P1_U3286) );
  INV_X1 U8769 ( .A(n7170), .ZN(n8559) );
  OAI222_X1 U8770 ( .A1(n8242), .A2(n7172), .B1(n8973), .B2(n8559), .C1(n7171), 
        .C2(P2_U3152), .ZN(P2_U3337) );
  NAND2_X1 U8771 ( .A1(n9086), .A2(n7251), .ZN(n7173) );
  AND2_X1 U8772 ( .A1(n7174), .A2(n7173), .ZN(n7176) );
  INV_X1 U8773 ( .A(n9085), .ZN(n7291) );
  NAND2_X1 U8774 ( .A1(n7291), .A2(n7328), .ZN(n8310) );
  INV_X1 U8775 ( .A(n7328), .ZN(n9773) );
  NAND2_X1 U8776 ( .A1(n7174), .A2(n7293), .ZN(n7175) );
  OAI21_X1 U8777 ( .B1(n7176), .B2(n8307), .A(n7175), .ZN(n9777) );
  INV_X1 U8778 ( .A(n9777), .ZN(n7184) );
  INV_X1 U8779 ( .A(n9502), .ZN(n9721) );
  INV_X1 U8780 ( .A(n8307), .ZN(n7179) );
  NAND2_X1 U8781 ( .A1(n7177), .A2(n8427), .ZN(n7178) );
  NAND2_X1 U8782 ( .A1(n8308), .A2(n7179), .ZN(n8311) );
  OAI21_X1 U8783 ( .B1(n7179), .B2(n8308), .A(n8311), .ZN(n7182) );
  OAI22_X1 U8784 ( .A1(n7413), .A2(n9348), .B1(n7180), .B2(n9346), .ZN(n7181)
         );
  AOI21_X1 U8785 ( .B1(n7182), .B2(n9717), .A(n7181), .ZN(n7183) );
  OAI21_X1 U8786 ( .B1(n7184), .B2(n9721), .A(n7183), .ZN(n9775) );
  INV_X1 U8787 ( .A(n9775), .ZN(n7192) );
  INV_X1 U8788 ( .A(n7284), .ZN(n7187) );
  NAND2_X1 U8789 ( .A1(n7185), .A2(n7328), .ZN(n7186) );
  NAND2_X1 U8790 ( .A1(n7187), .A2(n7186), .ZN(n9774) );
  AOI22_X1 U8791 ( .A1(n9728), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n7329), .B2(
        n9541), .ZN(n7189) );
  NAND2_X1 U8792 ( .A1(n9543), .A2(n7328), .ZN(n7188) );
  OAI211_X1 U8793 ( .C1(n9774), .C2(n9166), .A(n7189), .B(n7188), .ZN(n7190)
         );
  AOI21_X1 U8794 ( .B1(n9777), .B2(n9510), .A(n7190), .ZN(n7191) );
  OAI21_X1 U8795 ( .B1(n7192), .B2(n9728), .A(n7191), .ZN(P1_U3285) );
  XNOR2_X1 U8796 ( .A(n7203), .B(n7193), .ZN(n7194) );
  NAND2_X1 U8797 ( .A1(n7194), .A2(n8843), .ZN(n7196) );
  AOI22_X1 U8798 ( .A1(n8838), .A2(n6419), .B1(n8655), .B2(n8840), .ZN(n7195)
         );
  NAND2_X1 U8799 ( .A1(n7196), .A2(n7195), .ZN(n9855) );
  INV_X1 U8800 ( .A(n9855), .ZN(n7206) );
  NOR2_X1 U8801 ( .A1(n9834), .A2(n4661), .ZN(n7201) );
  OR2_X1 U8802 ( .A1(n7197), .A2(n6951), .ZN(n9853) );
  NAND2_X1 U8803 ( .A1(n9853), .A2(n9852), .ZN(n7199) );
  INV_X1 U8804 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7198) );
  OAI22_X1 U8805 ( .A1(n8685), .A2(n7199), .B1(n7198), .B2(n9825), .ZN(n7200)
         );
  AOI211_X1 U8806 ( .C1(n8755), .C2(n5859), .A(n7201), .B(n7200), .ZN(n7205)
         );
  INV_X1 U8807 ( .A(n8855), .ZN(n8813) );
  XNOR2_X1 U8808 ( .A(n7203), .B(n7202), .ZN(n9857) );
  NAND2_X1 U8809 ( .A1(n8813), .A2(n9857), .ZN(n7204) );
  OAI211_X1 U8810 ( .C1(n9836), .C2(n7206), .A(n7205), .B(n7204), .ZN(P2_U3295) );
  AND2_X1 U8811 ( .A1(n7208), .A2(n7207), .ZN(n7210) );
  OAI21_X1 U8812 ( .B1(n7210), .B2(n7222), .A(n7209), .ZN(n7213) );
  OAI22_X1 U8813 ( .A1(n7211), .A2(n8828), .B1(n7554), .B2(n8830), .ZN(n7212)
         );
  AOI21_X1 U8814 ( .B1(n7213), .B2(n8843), .A(n7212), .ZN(n9879) );
  OAI22_X1 U8815 ( .A1(n9834), .A2(n7215), .B1(n7214), .B2(n9825), .ZN(n7220)
         );
  AND2_X1 U8816 ( .A1(n7216), .A2(n7221), .ZN(n7218) );
  OR2_X1 U8817 ( .A1(n7218), .A2(n7217), .ZN(n9876) );
  NOR2_X1 U8818 ( .A1(n9876), .A2(n8685), .ZN(n7219) );
  AOI211_X1 U8819 ( .C1(n8755), .C2(n7221), .A(n7220), .B(n7219), .ZN(n7226)
         );
  INV_X1 U8820 ( .A(n7222), .ZN(n7223) );
  XNOR2_X1 U8821 ( .A(n7224), .B(n7223), .ZN(n9874) );
  NAND2_X1 U8822 ( .A1(n9874), .A2(n8813), .ZN(n7225) );
  OAI211_X1 U8823 ( .C1(n9879), .C2(n9836), .A(n7226), .B(n7225), .ZN(P2_U3290) );
  INV_X1 U8824 ( .A(n7228), .ZN(n7230) );
  INV_X1 U8825 ( .A(n7227), .ZN(n7229) );
  AND2_X1 U8826 ( .A1(n7228), .A2(n7227), .ZN(n7320) );
  AOI21_X1 U8827 ( .B1(n7230), .B2(n7229), .A(n7320), .ZN(n7231) );
  NAND2_X1 U8828 ( .A1(n7231), .A2(n7232), .ZN(n7322) );
  OAI21_X1 U8829 ( .B1(n7232), .B2(n7231), .A(n7322), .ZN(n7238) );
  AND2_X1 U8830 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n9633) );
  AOI21_X1 U8831 ( .B1(n9067), .B2(n9085), .A(n9633), .ZN(n7235) );
  AOI22_X1 U8832 ( .A1(n9049), .A2(n7233), .B1(n7251), .B2(n9037), .ZN(n7234)
         );
  OAI211_X1 U8833 ( .C1(n7236), .C2(n9058), .A(n7235), .B(n7234), .ZN(n7237)
         );
  AOI21_X1 U8834 ( .B1(n7238), .B2(n5747), .A(n7237), .ZN(n7239) );
  INV_X1 U8835 ( .A(n7239), .ZN(P1_U3225) );
  INV_X1 U8836 ( .A(n7241), .ZN(n7242) );
  AOI21_X1 U8837 ( .B1(n7243), .B2(n7240), .A(n7242), .ZN(n7249) );
  AOI21_X1 U8838 ( .B1(n9068), .B2(n9085), .A(n7244), .ZN(n7246) );
  NAND2_X1 U8839 ( .A1(n9049), .A2(n7287), .ZN(n7245) );
  OAI211_X1 U8840 ( .C1(n7409), .C2(n9014), .A(n7246), .B(n7245), .ZN(n7247)
         );
  AOI21_X1 U8841 ( .B1(n7581), .B2(n9073), .A(n7247), .ZN(n7248) );
  OAI21_X1 U8842 ( .B1(n7249), .B2(n9075), .A(n7248), .ZN(P1_U3211) );
  INV_X1 U8843 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n7256) );
  INV_X1 U8844 ( .A(n9783), .ZN(n9440) );
  INV_X1 U8845 ( .A(n9787), .ZN(n9436) );
  AOI21_X1 U8846 ( .B1(n9436), .B2(n7251), .A(n7250), .ZN(n7252) );
  OAI211_X1 U8847 ( .C1(n9440), .C2(n7254), .A(n7253), .B(n7252), .ZN(n7257)
         );
  NAND2_X1 U8848 ( .A1(n7257), .A2(n9806), .ZN(n7255) );
  OAI21_X1 U8849 ( .B1(n9806), .B2(n7256), .A(n7255), .ZN(P1_U3528) );
  INV_X1 U8850 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n7259) );
  NAND2_X1 U8851 ( .A1(n7257), .A2(n9795), .ZN(n7258) );
  OAI21_X1 U8852 ( .B1(n9795), .B2(n7259), .A(n7258), .ZN(P1_U3469) );
  INV_X1 U8853 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10083) );
  INV_X1 U8854 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10060) );
  AOI22_X1 U8855 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(P1_ADDR_REG_18__SCAN_IN), 
        .B1(n10083), .B2(n10060), .ZN(n10261) );
  NOR2_X1 U8856 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(P2_ADDR_REG_17__SCAN_IN), 
        .ZN(n7260) );
  AOI21_X1 U8857 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n7260), .ZN(n9926) );
  INV_X1 U8858 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n7261) );
  INV_X1 U8859 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n10194) );
  AOI22_X1 U8860 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(P2_ADDR_REG_16__SCAN_IN), 
        .B1(n7261), .B2(n10194), .ZN(n9929) );
  NOR2_X1 U8861 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7262) );
  AOI21_X1 U8862 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n7262), .ZN(n9932) );
  NOR2_X1 U8863 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7263) );
  AOI21_X1 U8864 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n7263), .ZN(n9935) );
  NOR2_X1 U8865 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7264) );
  AOI21_X1 U8866 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n7264), .ZN(n9938) );
  NOR2_X1 U8867 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7265) );
  AOI21_X1 U8868 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n7265), .ZN(n9941) );
  NOR2_X1 U8869 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n7266) );
  AOI21_X1 U8870 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n7266), .ZN(n9944) );
  NOR2_X1 U8871 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n7267) );
  AOI21_X1 U8872 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n7267), .ZN(n9947) );
  NOR2_X1 U8873 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n7268) );
  AOI21_X1 U8874 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(P2_ADDR_REG_9__SCAN_IN), 
        .A(n7268), .ZN(n10264) );
  NOR2_X1 U8875 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n7269) );
  AOI21_X1 U8876 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(P2_ADDR_REG_8__SCAN_IN), 
        .A(n7269), .ZN(n10249) );
  NOR2_X1 U8877 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n7270) );
  AOI21_X1 U8878 ( .B1(P1_ADDR_REG_7__SCAN_IN), .B2(P2_ADDR_REG_7__SCAN_IN), 
        .A(n7270), .ZN(n10258) );
  NOR2_X1 U8879 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(P2_ADDR_REG_6__SCAN_IN), 
        .ZN(n7271) );
  AOI21_X1 U8880 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(P1_ADDR_REG_6__SCAN_IN), 
        .A(n7271), .ZN(n10252) );
  NOR2_X1 U8881 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(P2_ADDR_REG_5__SCAN_IN), 
        .ZN(n7272) );
  AOI21_X1 U8882 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(P1_ADDR_REG_5__SCAN_IN), 
        .A(n7272), .ZN(n10255) );
  NAND2_X1 U8883 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n9922) );
  INV_X1 U8884 ( .A(n9922), .ZN(n7273) );
  NAND2_X1 U8885 ( .A1(n9922), .A2(n6671), .ZN(n9920) );
  AOI22_X1 U8886 ( .A1(n7273), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P2_ADDR_REG_1__SCAN_IN), .B2(n9920), .ZN(n10267) );
  NAND2_X1 U8887 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n7274) );
  OAI21_X1 U8888 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(P1_ADDR_REG_2__SCAN_IN), 
        .A(n7274), .ZN(n10266) );
  NOR2_X1 U8889 ( .A1(n10267), .A2(n10266), .ZN(n10265) );
  AOI21_X1 U8890 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(P2_ADDR_REG_2__SCAN_IN), 
        .A(n10265), .ZN(n10270) );
  NAND2_X1 U8891 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7275) );
  OAI21_X1 U8892 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n7275), .ZN(n10269) );
  NOR2_X1 U8893 ( .A1(n10270), .A2(n10269), .ZN(n10268) );
  AOI21_X1 U8894 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(P1_ADDR_REG_3__SCAN_IN), 
        .A(n10268), .ZN(n10273) );
  NOR2_X1 U8895 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(P1_ADDR_REG_4__SCAN_IN), 
        .ZN(n7276) );
  AOI21_X1 U8896 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(P2_ADDR_REG_4__SCAN_IN), 
        .A(n7276), .ZN(n10272) );
  NAND2_X1 U8897 ( .A1(n10273), .A2(n10272), .ZN(n10271) );
  OAI21_X1 U8898 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(P1_ADDR_REG_4__SCAN_IN), 
        .A(n10271), .ZN(n10254) );
  NAND2_X1 U8899 ( .A1(n10255), .A2(n10254), .ZN(n10253) );
  OAI21_X1 U8900 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(P2_ADDR_REG_5__SCAN_IN), 
        .A(n10253), .ZN(n10251) );
  NAND2_X1 U8901 ( .A1(n10252), .A2(n10251), .ZN(n10250) );
  OAI21_X1 U8902 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(P2_ADDR_REG_6__SCAN_IN), 
        .A(n10250), .ZN(n10257) );
  NAND2_X1 U8903 ( .A1(n10258), .A2(n10257), .ZN(n10256) );
  OAI21_X1 U8904 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(P1_ADDR_REG_7__SCAN_IN), 
        .A(n10256), .ZN(n10248) );
  NAND2_X1 U8905 ( .A1(n10249), .A2(n10248), .ZN(n10247) );
  OAI21_X1 U8906 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(P1_ADDR_REG_8__SCAN_IN), 
        .A(n10247), .ZN(n10263) );
  NAND2_X1 U8907 ( .A1(n10264), .A2(n10263), .ZN(n10262) );
  OAI21_X1 U8908 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(P1_ADDR_REG_9__SCAN_IN), 
        .A(n10262), .ZN(n9946) );
  NAND2_X1 U8909 ( .A1(n9947), .A2(n9946), .ZN(n9945) );
  OAI21_X1 U8910 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n9945), .ZN(n9943) );
  NAND2_X1 U8911 ( .A1(n9944), .A2(n9943), .ZN(n9942) );
  OAI21_X1 U8912 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n9942), .ZN(n9940) );
  NAND2_X1 U8913 ( .A1(n9941), .A2(n9940), .ZN(n9939) );
  OAI21_X1 U8914 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n9939), .ZN(n9937) );
  NAND2_X1 U8915 ( .A1(n9938), .A2(n9937), .ZN(n9936) );
  OAI21_X1 U8916 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n9936), .ZN(n9934) );
  NAND2_X1 U8917 ( .A1(n9935), .A2(n9934), .ZN(n9933) );
  OAI21_X1 U8918 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n9933), .ZN(n9931) );
  NAND2_X1 U8919 ( .A1(n9932), .A2(n9931), .ZN(n9930) );
  OAI21_X1 U8920 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n9930), .ZN(n9928) );
  NAND2_X1 U8921 ( .A1(n9929), .A2(n9928), .ZN(n9927) );
  OAI21_X1 U8922 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n9927), .ZN(n9925) );
  NAND2_X1 U8923 ( .A1(n9926), .A2(n9925), .ZN(n9924) );
  OAI21_X1 U8924 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n9924), .ZN(n10260) );
  NAND2_X1 U8925 ( .A1(n10261), .A2(n10260), .ZN(n10259) );
  OAI21_X1 U8926 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(P1_ADDR_REG_18__SCAN_IN), 
        .A(n10259), .ZN(n7278) );
  XNOR2_X1 U8927 ( .A(n4504), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n7277) );
  XNOR2_X1 U8928 ( .A(n7278), .B(n7277), .ZN(ADD_1071_U4) );
  NAND2_X1 U8929 ( .A1(n8310), .A2(n7279), .ZN(n8476) );
  INV_X1 U8930 ( .A(n7280), .ZN(n8429) );
  OR2_X1 U8931 ( .A1(n8476), .A2(n8429), .ZN(n7282) );
  NAND2_X1 U8932 ( .A1(n8434), .A2(n8427), .ZN(n7281) );
  NAND2_X1 U8933 ( .A1(n8310), .A2(n7281), .ZN(n8432) );
  NAND2_X1 U8934 ( .A1(n7282), .A2(n8432), .ZN(n8527) );
  NAND2_X1 U8935 ( .A1(n8311), .A2(n8527), .ZN(n7410) );
  INV_X1 U8936 ( .A(n7581), .ZN(n7414) );
  NAND2_X1 U8937 ( .A1(n7414), .A2(n9084), .ZN(n8425) );
  NAND2_X1 U8938 ( .A1(n7413), .A2(n7581), .ZN(n8435) );
  NAND2_X1 U8939 ( .A1(n8425), .A2(n8435), .ZN(n7300) );
  INV_X1 U8940 ( .A(n7300), .ZN(n8478) );
  XNOR2_X1 U8941 ( .A(n7410), .B(n8478), .ZN(n7283) );
  AOI222_X1 U8942 ( .A1(n9717), .A2(n7283), .B1(n9083), .B2(n9711), .C1(n9085), 
        .C2(n9713), .ZN(n7583) );
  INV_X1 U8943 ( .A(n9788), .ZN(n9704) );
  OAI21_X1 U8944 ( .B1(n7284), .B2(n7414), .A(n9704), .ZN(n7285) );
  NOR2_X1 U8945 ( .A1(n7285), .A2(n7423), .ZN(n7580) );
  NOR2_X1 U8946 ( .A1(n7286), .A2(n5505), .ZN(n9550) );
  INV_X1 U8947 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7290) );
  NAND2_X1 U8948 ( .A1(n9543), .A2(n7581), .ZN(n7289) );
  NAND2_X1 U8949 ( .A1(n9541), .A2(n7287), .ZN(n7288) );
  OAI211_X1 U8950 ( .C1(n9725), .C2(n7290), .A(n7289), .B(n7288), .ZN(n7304)
         );
  AND2_X1 U8951 ( .A1(n9773), .A2(n7291), .ZN(n7294) );
  OR2_X1 U8952 ( .A1(n7292), .A2(n7294), .ZN(n7415) );
  OR2_X1 U8953 ( .A1(n7420), .A2(n7415), .ZN(n7298) );
  AND2_X1 U8954 ( .A1(n7298), .A2(n7297), .ZN(n7301) );
  AND2_X1 U8955 ( .A1(n7297), .A2(n7300), .ZN(n7416) );
  NAND2_X1 U8956 ( .A1(n7298), .A2(n7416), .ZN(n7299) );
  OAI21_X1 U8957 ( .B1(n7301), .B2(n7300), .A(n7299), .ZN(n7302) );
  INV_X1 U8958 ( .A(n7302), .ZN(n7584) );
  NOR2_X1 U8959 ( .A1(n7584), .A2(n9368), .ZN(n7303) );
  AOI211_X1 U8960 ( .C1(n7580), .C2(n9550), .A(n7304), .B(n7303), .ZN(n7305)
         );
  OAI21_X1 U8961 ( .B1(n9728), .B2(n7583), .A(n7305), .ZN(P1_U3284) );
  XNOR2_X1 U8962 ( .A(n7306), .B(n7307), .ZN(n9863) );
  INV_X1 U8963 ( .A(n9863), .ZN(n7319) );
  OAI21_X1 U8964 ( .B1(n7310), .B2(n7309), .A(n7308), .ZN(n7311) );
  AOI222_X1 U8965 ( .A1(n8843), .A2(n7311), .B1(n8654), .B2(n8840), .C1(n8656), 
        .C2(n8838), .ZN(n9860) );
  NOR2_X1 U8966 ( .A1(n9860), .A2(n9836), .ZN(n7317) );
  NOR2_X1 U8967 ( .A1(n8851), .A2(n9858), .ZN(n7316) );
  NOR2_X1 U8968 ( .A1(n9834), .A2(n5826), .ZN(n7315) );
  NAND2_X1 U8969 ( .A1(n9852), .A2(n7312), .ZN(n7313) );
  NAND2_X1 U8970 ( .A1(n7505), .A2(n7313), .ZN(n9859) );
  OAI22_X1 U8971 ( .A1(n8685), .A2(n9859), .B1(n5825), .B2(n9825), .ZN(n7314)
         );
  NOR4_X1 U8972 ( .A1(n7317), .A2(n7316), .A3(n7315), .A4(n7314), .ZN(n7318)
         );
  OAI21_X1 U8973 ( .B1(n7319), .B2(n8855), .A(n7318), .ZN(P2_U3294) );
  INV_X1 U8974 ( .A(n7320), .ZN(n7321) );
  NAND2_X1 U8975 ( .A1(n7322), .A2(n7321), .ZN(n7326) );
  XNOR2_X1 U8976 ( .A(n7324), .B(n7323), .ZN(n7325) );
  XNOR2_X1 U8977 ( .A(n7326), .B(n7325), .ZN(n7335) );
  NOR2_X1 U8978 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7327), .ZN(n9648) );
  AOI21_X1 U8979 ( .B1(n9067), .B2(n9084), .A(n9648), .ZN(n7333) );
  NAND2_X1 U8980 ( .A1(n9073), .A2(n7328), .ZN(n7332) );
  NAND2_X1 U8981 ( .A1(n9049), .A2(n7329), .ZN(n7331) );
  NAND2_X1 U8982 ( .A1(n9068), .A2(n9086), .ZN(n7330) );
  NAND4_X1 U8983 ( .A1(n7333), .A2(n7332), .A3(n7331), .A4(n7330), .ZN(n7334)
         );
  AOI21_X1 U8984 ( .B1(n7335), .B2(n5747), .A(n7334), .ZN(n7336) );
  INV_X1 U8985 ( .A(n7336), .ZN(P1_U3237) );
  INV_X1 U8986 ( .A(n7341), .ZN(n9849) );
  AOI22_X1 U8987 ( .A1(n9849), .A2(n8843), .B1(n8840), .B2(n8656), .ZN(n9851)
         );
  OAI22_X1 U8988 ( .A1(n9851), .A2(n9836), .B1(n7337), .B2(n9825), .ZN(n7338)
         );
  AOI21_X1 U8989 ( .B1(P2_REG2_REG_0__SCAN_IN), .B2(n9836), .A(n7338), .ZN(
        n7340) );
  OAI21_X1 U8990 ( .B1(n8755), .B2(n8858), .A(n9847), .ZN(n7339) );
  OAI211_X1 U8991 ( .C1(n7341), .C2(n8855), .A(n7340), .B(n7339), .ZN(P2_U3296) );
  INV_X1 U8992 ( .A(n7342), .ZN(n7343) );
  NOR2_X1 U8993 ( .A1(n7553), .A2(n8271), .ZN(n7348) );
  XNOR2_X1 U8994 ( .A(n7646), .B(n8276), .ZN(n7347) );
  NOR2_X1 U8995 ( .A1(n7347), .A2(n7348), .ZN(n7349) );
  AOI21_X1 U8996 ( .B1(n7348), .B2(n7347), .A(n7349), .ZN(n7371) );
  NAND2_X1 U8997 ( .A1(n7372), .A2(n7371), .ZN(n7370) );
  INV_X1 U8998 ( .A(n7349), .ZN(n7350) );
  XNOR2_X1 U8999 ( .A(n9891), .B(n6957), .ZN(n7436) );
  NOR2_X1 U9000 ( .A1(n7473), .A2(n8271), .ZN(n7437) );
  XNOR2_X1 U9001 ( .A(n7436), .B(n7437), .ZN(n7440) );
  XNOR2_X1 U9002 ( .A(n7441), .B(n7440), .ZN(n7354) );
  OAI22_X1 U9003 ( .A1(n8615), .A2(n7616), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10223), .ZN(n7352) );
  OAI22_X1 U9004 ( .A1(n7553), .A2(n8602), .B1(n8603), .B2(n7707), .ZN(n7351)
         );
  AOI211_X1 U9005 ( .C1(n8629), .C2(n9891), .A(n7352), .B(n7351), .ZN(n7353)
         );
  OAI21_X1 U9006 ( .B1(n7354), .B2(n8631), .A(n7353), .ZN(P2_U3219) );
  XNOR2_X1 U9007 ( .A(n7355), .B(n7356), .ZN(n9873) );
  INV_X1 U9008 ( .A(n9873), .ZN(n7369) );
  NAND2_X1 U9009 ( .A1(n7357), .A2(n8843), .ZN(n7362) );
  AOI21_X1 U9010 ( .B1(n7495), .B2(n7359), .A(n7358), .ZN(n7361) );
  AOI22_X1 U9011 ( .A1(n8652), .A2(n8840), .B1(n8838), .B2(n8654), .ZN(n7360)
         );
  OAI21_X1 U9012 ( .B1(n7362), .B2(n7361), .A(n7360), .ZN(n9871) );
  XNOR2_X1 U9013 ( .A(n7504), .B(n9869), .ZN(n9870) );
  OAI22_X1 U9014 ( .A1(n9834), .A2(n5889), .B1(n7363), .B2(n9825), .ZN(n7364)
         );
  AOI21_X1 U9015 ( .B1(n8755), .B2(n7365), .A(n7364), .ZN(n7366) );
  OAI21_X1 U9016 ( .B1(n8685), .B2(n9870), .A(n7366), .ZN(n7367) );
  AOI21_X1 U9017 ( .B1(n9871), .B2(n9834), .A(n7367), .ZN(n7368) );
  OAI21_X1 U9018 ( .B1(n7369), .B2(n8855), .A(n7368), .ZN(P2_U3292) );
  INV_X1 U9019 ( .A(n7646), .ZN(n7484) );
  OAI21_X1 U9020 ( .B1(n7372), .B2(n7371), .A(n7370), .ZN(n7373) );
  NAND2_X1 U9021 ( .A1(n7373), .A2(n8611), .ZN(n7379) );
  INV_X1 U9022 ( .A(n7485), .ZN(n7377) );
  INV_X1 U9023 ( .A(n7374), .ZN(n7376) );
  OAI22_X1 U9024 ( .A1(n7474), .A2(n8602), .B1(n8603), .B2(n7473), .ZN(n7375)
         );
  AOI211_X1 U9025 ( .C1(n7377), .C2(n8625), .A(n7376), .B(n7375), .ZN(n7378)
         );
  OAI211_X1 U9026 ( .C1(n7484), .C2(n8620), .A(n7379), .B(n7378), .ZN(P2_U3233) );
  INV_X1 U9027 ( .A(n7380), .ZN(n7381) );
  AOI21_X1 U9028 ( .B1(n8474), .B2(n7382), .A(n7381), .ZN(n7386) );
  AOI22_X1 U9029 ( .A1(n9713), .A2(n5011), .B1(n9088), .B2(n9711), .ZN(n7385)
         );
  XNOR2_X1 U9030 ( .A(n8521), .B(n8474), .ZN(n7383) );
  NAND2_X1 U9031 ( .A1(n7383), .A2(n9717), .ZN(n7384) );
  OAI211_X1 U9032 ( .C1(n7386), .C2(n9721), .A(n7385), .B(n7384), .ZN(n9764)
         );
  INV_X1 U9033 ( .A(n9764), .ZN(n7394) );
  INV_X1 U9034 ( .A(n7386), .ZN(n9766) );
  NAND2_X1 U9035 ( .A1(n9703), .A2(n8209), .ZN(n7387) );
  NAND2_X1 U9036 ( .A1(n7388), .A2(n7387), .ZN(n9763) );
  AND2_X1 U9037 ( .A1(n9541), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n7390) );
  NOR2_X1 U9038 ( .A1(n9357), .A2(n9762), .ZN(n7389) );
  AOI211_X1 U9039 ( .C1(n9728), .C2(P1_REG2_REG_2__SCAN_IN), .A(n7390), .B(
        n7389), .ZN(n7391) );
  OAI21_X1 U9040 ( .B1(n9166), .B2(n9763), .A(n7391), .ZN(n7392) );
  AOI21_X1 U9041 ( .B1(n9510), .B2(n9766), .A(n7392), .ZN(n7393) );
  OAI21_X1 U9042 ( .B1(n9728), .B2(n7394), .A(n7393), .ZN(P1_U3289) );
  NAND2_X1 U9043 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3084), .ZN(n7401) );
  INV_X1 U9044 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n7395) );
  MUX2_X1 U9045 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n7395), .S(n7773), .Z(n7398)
         );
  OAI21_X1 U9046 ( .B1(P1_REG1_REG_13__SCAN_IN), .B2(n7403), .A(n7396), .ZN(
        n7397) );
  NAND2_X1 U9047 ( .A1(n7397), .A2(n7398), .ZN(n7772) );
  OAI21_X1 U9048 ( .B1(n7398), .B2(n7397), .A(n7772), .ZN(n7399) );
  NAND2_X1 U9049 ( .A1(n7399), .A2(n9694), .ZN(n7400) );
  OAI211_X1 U9050 ( .C1(n7900), .C2(n7766), .A(n7401), .B(n7400), .ZN(n7407)
         );
  INV_X1 U9051 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7404) );
  AOI211_X1 U9052 ( .C1(n7405), .C2(n7404), .A(n7768), .B(n9659), .ZN(n7406)
         );
  AOI211_X1 U9053 ( .C1(n9668), .C2(P1_ADDR_REG_14__SCAN_IN), .A(n7407), .B(
        n7406), .ZN(n7408) );
  INV_X1 U9054 ( .A(n7408), .ZN(P1_U3255) );
  INV_X1 U9055 ( .A(n9497), .ZN(n7597) );
  NAND2_X1 U9056 ( .A1(n7595), .A2(n7409), .ZN(n8436) );
  NAND2_X1 U9057 ( .A1(n7410), .A2(n8478), .ZN(n7411) );
  NAND2_X1 U9058 ( .A1(n7411), .A2(n8435), .ZN(n7534) );
  XOR2_X1 U9059 ( .A(n8479), .B(n7534), .Z(n7412) );
  OAI222_X1 U9060 ( .A1(n9348), .A2(n7597), .B1(n9346), .B2(n7413), .C1(n7412), 
        .C2(n9499), .ZN(n9781) );
  INV_X1 U9061 ( .A(n9781), .ZN(n7431) );
  AND2_X1 U9062 ( .A1(n7414), .A2(n7413), .ZN(n7417) );
  OR2_X1 U9063 ( .A1(n7420), .A2(n7419), .ZN(n7418) );
  OR2_X1 U9064 ( .A1(n7417), .A2(n7416), .ZN(n7421) );
  AND2_X1 U9065 ( .A1(n7418), .A2(n7421), .ZN(n7422) );
  AOI21_X1 U9066 ( .B1(n8479), .B2(n7422), .A(n4439), .ZN(n9784) );
  INV_X1 U9067 ( .A(n9368), .ZN(n9552) );
  INV_X1 U9068 ( .A(n7595), .ZN(n9779) );
  OR2_X1 U9069 ( .A1(n7423), .A2(n9779), .ZN(n7424) );
  NAND2_X1 U9070 ( .A1(n7540), .A2(n7424), .ZN(n9780) );
  INV_X1 U9071 ( .A(n7596), .ZN(n7425) );
  OAI22_X1 U9072 ( .A1(n9725), .A2(n7426), .B1(n7425), .B2(n9708), .ZN(n7427)
         );
  AOI21_X1 U9073 ( .B1(n9543), .B2(n7595), .A(n7427), .ZN(n7428) );
  OAI21_X1 U9074 ( .B1(n9780), .B2(n9166), .A(n7428), .ZN(n7429) );
  AOI21_X1 U9075 ( .B1(n9784), .B2(n9552), .A(n7429), .ZN(n7430) );
  OAI21_X1 U9076 ( .B1(n9728), .B2(n7431), .A(n7430), .ZN(P1_U3283) );
  INV_X1 U9077 ( .A(n7432), .ZN(n7435) );
  OAI222_X1 U9078 ( .A1(n8242), .A2(n7434), .B1(n8973), .B2(n7435), .C1(
        P2_U3152), .C2(n7433), .ZN(P2_U3336) );
  OAI222_X1 U9079 ( .A1(n8557), .A2(n10098), .B1(n4370), .B2(n7435), .C1(
        P1_U3084), .C2(n5743), .ZN(P1_U3331) );
  INV_X1 U9080 ( .A(n7436), .ZN(n7439) );
  INV_X1 U9081 ( .A(n7437), .ZN(n7438) );
  NOR2_X1 U9082 ( .A1(n7707), .A2(n8271), .ZN(n7697) );
  XNOR2_X1 U9083 ( .A(n7670), .B(n8276), .ZN(n7696) );
  XOR2_X1 U9084 ( .A(n7697), .B(n7696), .Z(n7698) );
  XNOR2_X1 U9085 ( .A(n7699), .B(n7698), .ZN(n7445) );
  OAI22_X1 U9086 ( .A1(n8615), .A2(n7632), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5967), .ZN(n7443) );
  OAI22_X1 U9087 ( .A1(n7473), .A2(n8602), .B1(n8603), .B2(n7760), .ZN(n7442)
         );
  AOI211_X1 U9088 ( .C1(n8629), .C2(n7670), .A(n7443), .B(n7442), .ZN(n7444)
         );
  OAI21_X1 U9089 ( .B1(n7445), .B2(n8631), .A(n7444), .ZN(P2_U3238) );
  INV_X1 U9090 ( .A(n7446), .ZN(n7516) );
  OR2_X1 U9091 ( .A1(n7447), .A2(P1_U3084), .ZN(n8549) );
  INV_X1 U9092 ( .A(n8549), .ZN(n8544) );
  AOI21_X1 U9093 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(n9459), .A(n8544), .ZN(
        n7448) );
  OAI21_X1 U9094 ( .B1(n7516), .B2(n4370), .A(n7448), .ZN(P1_U3330) );
  OAI21_X1 U9095 ( .B1(n7454), .B2(P2_REG2_REG_11__SCAN_IN), .A(n7449), .ZN(
        n7451) );
  XNOR2_X1 U9096 ( .A(n7518), .B(P2_REG2_REG_12__SCAN_IN), .ZN(n7450) );
  AOI211_X1 U9097 ( .C1(n7451), .C2(n7450), .A(n8657), .B(n7517), .ZN(n7452)
         );
  INV_X1 U9098 ( .A(n7452), .ZN(n7460) );
  AOI21_X1 U9099 ( .B1(n7454), .B2(P2_REG1_REG_11__SCAN_IN), .A(n7453), .ZN(
        n7456) );
  MUX2_X1 U9100 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n7521), .S(n7518), .Z(n7455)
         );
  NAND2_X1 U9101 ( .A1(n7456), .A2(n7455), .ZN(n7524) );
  OAI21_X1 U9102 ( .B1(n7456), .B2(n7455), .A(n7524), .ZN(n7458) );
  INV_X1 U9103 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n10177) );
  NAND2_X1 U9104 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3152), .ZN(n7706) );
  OAI21_X1 U9105 ( .B1(n8675), .B2(n10177), .A(n7706), .ZN(n7457) );
  AOI21_X1 U9106 ( .B1(n9807), .B2(n7458), .A(n7457), .ZN(n7459) );
  OAI211_X1 U9107 ( .C1(n9809), .C2(n7522), .A(n7460), .B(n7459), .ZN(P2_U3257) );
  INV_X1 U9108 ( .A(n7461), .ZN(n7462) );
  AOI22_X1 U9109 ( .A1(n9836), .A2(P2_REG2_REG_7__SCAN_IN), .B1(n7462), .B2(
        n8848), .ZN(n7463) );
  OAI21_X1 U9110 ( .B1(n7464), .B2(n8851), .A(n7463), .ZN(n7467) );
  NOR2_X1 U9111 ( .A1(n7465), .A2(n8855), .ZN(n7466) );
  AOI211_X1 U9112 ( .C1(n7468), .C2(n8858), .A(n7467), .B(n7466), .ZN(n7469)
         );
  OAI21_X1 U9113 ( .B1(n9836), .B2(n7470), .A(n7469), .ZN(P2_U3289) );
  OR2_X1 U9114 ( .A1(n7627), .A2(n7472), .ZN(n7607) );
  OAI21_X1 U9115 ( .B1(n4894), .B2(n7478), .A(n7607), .ZN(n7645) );
  INV_X1 U9116 ( .A(n7747), .ZN(n7494) );
  OAI22_X1 U9117 ( .A1(n7474), .A2(n8828), .B1(n7473), .B2(n8830), .ZN(n7482)
         );
  AND2_X1 U9118 ( .A1(n7476), .A2(n7475), .ZN(n7480) );
  NAND2_X1 U9119 ( .A1(n7551), .A2(n7552), .ZN(n7550) );
  NAND3_X1 U9120 ( .A1(n7550), .A2(n7478), .A3(n7477), .ZN(n7479) );
  INV_X1 U9121 ( .A(n8843), .ZN(n8825) );
  AOI21_X1 U9122 ( .B1(n7480), .B2(n7479), .A(n8825), .ZN(n7481) );
  AOI211_X1 U9123 ( .C1(n7645), .C2(n7494), .A(n7482), .B(n7481), .ZN(n7649)
         );
  INV_X1 U9124 ( .A(n7618), .ZN(n7483) );
  AOI21_X1 U9125 ( .B1(n7646), .B2(n4440), .A(n7483), .ZN(n7647) );
  NOR2_X1 U9126 ( .A1(n7484), .A2(n8851), .ZN(n7488) );
  OAI22_X1 U9127 ( .A1(n9834), .A2(n7486), .B1(n7485), .B2(n9825), .ZN(n7487)
         );
  AOI211_X1 U9128 ( .C1(n7647), .C2(n8858), .A(n7488), .B(n7487), .ZN(n7491)
         );
  OR2_X1 U9129 ( .A1(n9836), .A2(n7489), .ZN(n7755) );
  INV_X1 U9130 ( .A(n7755), .ZN(n7511) );
  NAND2_X1 U9131 ( .A1(n7645), .A2(n7511), .ZN(n7490) );
  OAI211_X1 U9132 ( .C1(n7649), .C2(n9836), .A(n7491), .B(n7490), .ZN(P2_U3287) );
  XNOR2_X1 U9133 ( .A(n7492), .B(n7493), .ZN(n9866) );
  NAND2_X1 U9134 ( .A1(n9866), .A2(n7494), .ZN(n7503) );
  OAI21_X1 U9135 ( .B1(n7497), .B2(n7496), .A(n7495), .ZN(n7501) );
  NAND2_X1 U9136 ( .A1(n8655), .A2(n8838), .ZN(n7499) );
  NAND2_X1 U9137 ( .A1(n8653), .A2(n8840), .ZN(n7498) );
  NAND2_X1 U9138 ( .A1(n7499), .A2(n7498), .ZN(n7500) );
  AOI21_X1 U9139 ( .B1(n7501), .B2(n8843), .A(n7500), .ZN(n7502) );
  AND2_X1 U9140 ( .A1(n7503), .A2(n7502), .ZN(n9868) );
  OAI22_X1 U9141 ( .A1(n9834), .A2(n5862), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n9825), .ZN(n7509) );
  INV_X1 U9142 ( .A(n7504), .ZN(n7507) );
  NAND2_X1 U9143 ( .A1(n7505), .A2(n7510), .ZN(n7506) );
  NAND2_X1 U9144 ( .A1(n7507), .A2(n7506), .ZN(n9864) );
  NOR2_X1 U9145 ( .A1(n9864), .A2(n8685), .ZN(n7508) );
  AOI211_X1 U9146 ( .C1(n8755), .C2(n7510), .A(n7509), .B(n7508), .ZN(n7513)
         );
  NAND2_X1 U9147 ( .A1(n9866), .A2(n7511), .ZN(n7512) );
  OAI211_X1 U9148 ( .C1(n9868), .C2(n9836), .A(n7513), .B(n7512), .ZN(P2_U3293) );
  NAND2_X1 U9149 ( .A1(n8970), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n7515) );
  OAI211_X1 U9150 ( .C1(n7516), .C2(n8973), .A(n7515), .B(n7514), .ZN(P2_U3335) );
  AOI22_X1 U9151 ( .A1(n7684), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n7748), .B2(
        n7530), .ZN(n7519) );
  OAI21_X1 U9152 ( .B1(n7520), .B2(n7519), .A(n7679), .ZN(n7532) );
  AOI22_X1 U9153 ( .A1(n9813), .A2(P2_ADDR_REG_13__SCAN_IN), .B1(
        P2_REG3_REG_13__SCAN_IN), .B2(P2_U3152), .ZN(n7529) );
  NAND2_X1 U9154 ( .A1(n7522), .A2(n7521), .ZN(n7523) );
  NAND2_X1 U9155 ( .A1(n7524), .A2(n7523), .ZN(n7526) );
  AOI22_X1 U9156 ( .A1(n7684), .A2(P2_REG1_REG_13__SCAN_IN), .B1(n5994), .B2(
        n7530), .ZN(n7525) );
  NAND2_X1 U9157 ( .A1(n7525), .A2(n7526), .ZN(n7685) );
  OAI21_X1 U9158 ( .B1(n7526), .B2(n7525), .A(n7685), .ZN(n7527) );
  NAND2_X1 U9159 ( .A1(n9807), .A2(n7527), .ZN(n7528) );
  OAI211_X1 U9160 ( .C1(n9809), .C2(n7530), .A(n7529), .B(n7528), .ZN(n7531)
         );
  AOI21_X1 U9161 ( .B1(n7532), .B2(n9808), .A(n7531), .ZN(n7533) );
  INV_X1 U9162 ( .A(n7533), .ZN(P2_U3258) );
  INV_X1 U9163 ( .A(n8436), .ZN(n8327) );
  NOR2_X1 U9164 ( .A1(n9786), .A2(n7597), .ZN(n8315) );
  NAND2_X1 U9165 ( .A1(n9786), .A2(n7597), .ZN(n9492) );
  INV_X1 U9166 ( .A(n9492), .ZN(n7535) );
  OR2_X1 U9167 ( .A1(n8315), .A2(n7535), .ZN(n8482) );
  XOR2_X1 U9168 ( .A(n7730), .B(n8482), .Z(n7539) );
  NAND2_X1 U9169 ( .A1(n7595), .A2(n9083), .ZN(n7536) );
  XOR2_X1 U9170 ( .A(n8482), .B(n7726), .Z(n9792) );
  NAND2_X1 U9171 ( .A1(n9792), .A2(n9502), .ZN(n7538) );
  AOI22_X1 U9172 ( .A1(n9713), .A2(n9083), .B1(n9082), .B2(n9711), .ZN(n7537)
         );
  OAI211_X1 U9173 ( .C1(n9499), .C2(n7539), .A(n7538), .B(n7537), .ZN(n9790)
         );
  INV_X1 U9174 ( .A(n9790), .ZN(n7546) );
  NAND2_X1 U9175 ( .A1(n7540), .A2(n9786), .ZN(n7541) );
  NAND2_X1 U9176 ( .A1(n9505), .A2(n7541), .ZN(n9789) );
  AOI22_X1 U9177 ( .A1(n9728), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n7660), .B2(
        n9541), .ZN(n7543) );
  NAND2_X1 U9178 ( .A1(n9543), .A2(n9786), .ZN(n7542) );
  OAI211_X1 U9179 ( .C1(n9789), .C2(n9166), .A(n7543), .B(n7542), .ZN(n7544)
         );
  AOI21_X1 U9180 ( .B1(n9792), .B2(n9510), .A(n7544), .ZN(n7545) );
  OAI21_X1 U9181 ( .B1(n7546), .B2(n9728), .A(n7545), .ZN(P1_U3282) );
  NAND2_X1 U9182 ( .A1(n7547), .A2(n7552), .ZN(n7548) );
  NAND2_X1 U9183 ( .A1(n7549), .A2(n7548), .ZN(n9887) );
  OAI21_X1 U9184 ( .B1(n7552), .B2(n7551), .A(n7550), .ZN(n7556) );
  OAI22_X1 U9185 ( .A1(n7554), .A2(n8828), .B1(n7553), .B2(n8830), .ZN(n7555)
         );
  AOI21_X1 U9186 ( .B1(n7556), .B2(n8843), .A(n7555), .ZN(n7558) );
  OR2_X1 U9187 ( .A1(n9887), .A2(n7747), .ZN(n7557) );
  NAND2_X1 U9188 ( .A1(n7558), .A2(n7557), .ZN(n9889) );
  MUX2_X1 U9189 ( .A(n9889), .B(P2_REG2_REG_8__SCAN_IN), .S(n9836), .Z(n7559)
         );
  INV_X1 U9190 ( .A(n7559), .ZN(n7566) );
  OR2_X1 U9191 ( .A1(n7560), .A2(n7563), .ZN(n7561) );
  AND2_X1 U9192 ( .A1(n4440), .A2(n7561), .ZN(n9884) );
  OAI22_X1 U9193 ( .A1(n8851), .A2(n7563), .B1(n9825), .B2(n7562), .ZN(n7564)
         );
  AOI21_X1 U9194 ( .B1(n9884), .B2(n8858), .A(n7564), .ZN(n7565) );
  OAI211_X1 U9195 ( .C1(n9887), .C2(n7755), .A(n7566), .B(n7565), .ZN(P2_U3288) );
  NAND2_X1 U9196 ( .A1(n7568), .A2(n7567), .ZN(n7569) );
  XNOR2_X1 U9197 ( .A(n7569), .B(n7572), .ZN(n7570) );
  OAI222_X1 U9198 ( .A1(n8830), .A2(n8643), .B1(n8828), .B2(n7707), .C1(n8825), 
        .C2(n7570), .ZN(n9903) );
  INV_X1 U9199 ( .A(n9903), .ZN(n7579) );
  XNOR2_X1 U9200 ( .A(n7571), .B(n7572), .ZN(n9906) );
  NOR2_X1 U9201 ( .A1(n7637), .A2(n9900), .ZN(n7573) );
  OR2_X1 U9202 ( .A1(n7749), .A2(n7573), .ZN(n9902) );
  INV_X1 U9203 ( .A(n7574), .ZN(n7710) );
  AOI22_X1 U9204 ( .A1(n9836), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n7710), .B2(
        n8848), .ZN(n7576) );
  NAND2_X1 U9205 ( .A1(n7700), .A2(n8755), .ZN(n7575) );
  OAI211_X1 U9206 ( .C1(n9902), .C2(n8685), .A(n7576), .B(n7575), .ZN(n7577)
         );
  AOI21_X1 U9207 ( .B1(n9906), .B2(n8813), .A(n7577), .ZN(n7578) );
  OAI21_X1 U9208 ( .B1(n7579), .B2(n9836), .A(n7578), .ZN(P2_U3284) );
  INV_X1 U9209 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n7586) );
  AOI21_X1 U9210 ( .B1(n9436), .B2(n7581), .A(n7580), .ZN(n7582) );
  OAI211_X1 U9211 ( .C1(n7584), .C2(n9440), .A(n7583), .B(n7582), .ZN(n7587)
         );
  NAND2_X1 U9212 ( .A1(n7587), .A2(n9806), .ZN(n7585) );
  OAI21_X1 U9213 ( .B1(n9806), .B2(n7586), .A(n7585), .ZN(P1_U3530) );
  INV_X1 U9214 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n7589) );
  NAND2_X1 U9215 ( .A1(n7587), .A2(n9795), .ZN(n7588) );
  OAI21_X1 U9216 ( .B1(n9795), .B2(n7589), .A(n7588), .ZN(P1_U3475) );
  NAND2_X1 U9217 ( .A1(n7591), .A2(n7590), .ZN(n7593) );
  XNOR2_X1 U9218 ( .A(n7593), .B(n7592), .ZN(n7603) );
  AOI21_X1 U9219 ( .B1(n9068), .B2(n9084), .A(n7594), .ZN(n7601) );
  NAND2_X1 U9220 ( .A1(n9073), .A2(n7595), .ZN(n7600) );
  NAND2_X1 U9221 ( .A1(n9049), .A2(n7596), .ZN(n7599) );
  OR2_X1 U9222 ( .A1(n9014), .A2(n7597), .ZN(n7598) );
  NAND4_X1 U9223 ( .A1(n7601), .A2(n7600), .A3(n7599), .A4(n7598), .ZN(n7602)
         );
  AOI21_X1 U9224 ( .B1(n7603), .B2(n5747), .A(n7602), .ZN(n7604) );
  INV_X1 U9225 ( .A(n7604), .ZN(P1_U3219) );
  NAND2_X1 U9226 ( .A1(n7607), .A2(n7605), .ZN(n7610) );
  NAND2_X1 U9227 ( .A1(n7607), .A2(n7606), .ZN(n7608) );
  NAND2_X1 U9228 ( .A1(n7608), .A2(n7611), .ZN(n7609) );
  NAND2_X1 U9229 ( .A1(n7610), .A2(n7609), .ZN(n9890) );
  AOI22_X1 U9230 ( .A1(n8838), .A2(n8648), .B1(n8646), .B2(n8840), .ZN(n7615)
         );
  XNOR2_X1 U9231 ( .A(n7612), .B(n7611), .ZN(n7613) );
  NAND2_X1 U9232 ( .A1(n7613), .A2(n8843), .ZN(n7614) );
  OAI211_X1 U9233 ( .C1(n9890), .C2(n7747), .A(n7615), .B(n7614), .ZN(n9894)
         );
  NAND2_X1 U9234 ( .A1(n9894), .A2(n9834), .ZN(n7623) );
  OAI22_X1 U9235 ( .A1(n9834), .A2(n7617), .B1(n7616), .B2(n9825), .ZN(n7621)
         );
  NAND2_X1 U9236 ( .A1(n7618), .A2(n9891), .ZN(n7619) );
  NAND2_X1 U9237 ( .A1(n7635), .A2(n7619), .ZN(n9893) );
  NOR2_X1 U9238 ( .A1(n9893), .A2(n8685), .ZN(n7620) );
  AOI211_X1 U9239 ( .C1(n8755), .C2(n9891), .A(n7621), .B(n7620), .ZN(n7622)
         );
  OAI211_X1 U9240 ( .C1(n9890), .C2(n7755), .A(n7623), .B(n7622), .ZN(P2_U3286) );
  XNOR2_X1 U9241 ( .A(n7624), .B(n7630), .ZN(n7625) );
  AOI222_X1 U9242 ( .A1(n8843), .A2(n7625), .B1(n8645), .B2(n8840), .C1(n8647), 
        .C2(n8838), .ZN(n7673) );
  OR2_X1 U9243 ( .A1(n7627), .A2(n7626), .ZN(n7629) );
  AND2_X1 U9244 ( .A1(n7629), .A2(n7628), .ZN(n7631) );
  XNOR2_X1 U9245 ( .A(n7631), .B(n7630), .ZN(n7674) );
  OAI22_X1 U9246 ( .A1(n9834), .A2(n7633), .B1(n7632), .B2(n9825), .ZN(n7634)
         );
  AOI21_X1 U9247 ( .B1(n7670), .B2(n8755), .A(n7634), .ZN(n7639) );
  AND2_X1 U9248 ( .A1(n7635), .A2(n7670), .ZN(n7636) );
  NOR2_X1 U9249 ( .A1(n7637), .A2(n7636), .ZN(n7671) );
  NAND2_X1 U9250 ( .A1(n7671), .A2(n8858), .ZN(n7638) );
  OAI211_X1 U9251 ( .C1(n7674), .C2(n8855), .A(n7639), .B(n7638), .ZN(n7640)
         );
  INV_X1 U9252 ( .A(n7640), .ZN(n7641) );
  OAI21_X1 U9253 ( .B1(n7673), .B2(n9836), .A(n7641), .ZN(P2_U3285) );
  INV_X1 U9254 ( .A(n7642), .ZN(n7668) );
  OAI222_X1 U9255 ( .A1(n4370), .A2(n7668), .B1(P1_U3084), .B2(n7644), .C1(
        n7643), .C2(n8557), .ZN(P1_U3329) );
  INV_X1 U9256 ( .A(n7645), .ZN(n7650) );
  AOI22_X1 U9257 ( .A1(n7647), .A2(n9883), .B1(n9882), .B2(n7646), .ZN(n7648)
         );
  OAI211_X1 U9258 ( .C1(n7650), .C2(n9886), .A(n7649), .B(n7648), .ZN(n7653)
         );
  NAND2_X1 U9259 ( .A1(n7653), .A2(n9996), .ZN(n7651) );
  OAI21_X1 U9260 ( .B1(n9996), .B2(n7652), .A(n7651), .ZN(P2_U3529) );
  NAND2_X1 U9261 ( .A1(n7653), .A2(n9909), .ZN(n7654) );
  OAI21_X1 U9262 ( .B1(n9909), .B2(n5938), .A(n7654), .ZN(P2_U3478) );
  NAND2_X1 U9264 ( .A1(n7657), .A2(n7658), .ZN(n7659) );
  AOI21_X1 U9265 ( .B1(n7656), .B2(n7659), .A(n9075), .ZN(n7666) );
  AND2_X1 U9266 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n9663) );
  AOI21_X1 U9267 ( .B1(n9067), .B2(n9082), .A(n9663), .ZN(n7664) );
  NAND2_X1 U9268 ( .A1(n9786), .A2(n9073), .ZN(n7663) );
  NAND2_X1 U9269 ( .A1(n9049), .A2(n7660), .ZN(n7662) );
  NAND2_X1 U9270 ( .A1(n9068), .A2(n9083), .ZN(n7661) );
  NAND4_X1 U9271 ( .A1(n7664), .A2(n7663), .A3(n7662), .A4(n7661), .ZN(n7665)
         );
  OR2_X1 U9272 ( .A1(n7666), .A2(n7665), .ZN(P1_U3229) );
  OAI222_X1 U9273 ( .A1(P2_U3152), .A2(n7669), .B1(n8973), .B2(n7668), .C1(
        n7667), .C2(n8242), .ZN(P2_U3334) );
  INV_X1 U9274 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n7676) );
  AOI22_X1 U9275 ( .A1(n7671), .A2(n9883), .B1(n9882), .B2(n7670), .ZN(n7672)
         );
  OAI211_X1 U9276 ( .C1(n9532), .C2(n7674), .A(n7673), .B(n7672), .ZN(n7677)
         );
  NAND2_X1 U9277 ( .A1(n7677), .A2(n9909), .ZN(n7675) );
  OAI21_X1 U9278 ( .B1(n9909), .B2(n7676), .A(n7675), .ZN(P2_U3484) );
  NAND2_X1 U9279 ( .A1(n7677), .A2(n9996), .ZN(n7678) );
  OAI21_X1 U9280 ( .B1(n9996), .B2(n7111), .A(n7678), .ZN(P2_U3531) );
  AOI22_X1 U9281 ( .A1(n7872), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n5800), .B2(
        n7692), .ZN(n7681) );
  NAND2_X1 U9282 ( .A1(n7681), .A2(n7680), .ZN(n7869) );
  OAI21_X1 U9283 ( .B1(n7681), .B2(n7680), .A(n7869), .ZN(n7694) );
  NAND2_X1 U9284 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3152), .ZN(n7835) );
  INV_X1 U9285 ( .A(n7835), .ZN(n7682) );
  AOI21_X1 U9286 ( .B1(n9813), .B2(P2_ADDR_REG_14__SCAN_IN), .A(n7682), .ZN(
        n7691) );
  MUX2_X1 U9287 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n7683), .S(n7872), .Z(n7688)
         );
  OR2_X1 U9288 ( .A1(n7684), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n7686) );
  NAND2_X1 U9289 ( .A1(n7686), .A2(n7685), .ZN(n7687) );
  NAND2_X1 U9290 ( .A1(n7688), .A2(n7687), .ZN(n7871) );
  OAI21_X1 U9291 ( .B1(n7688), .B2(n7687), .A(n7871), .ZN(n7689) );
  NAND2_X1 U9292 ( .A1(n9807), .A2(n7689), .ZN(n7690) );
  OAI211_X1 U9293 ( .C1(n9809), .C2(n7692), .A(n7691), .B(n7690), .ZN(n7693)
         );
  AOI21_X1 U9294 ( .B1(n9808), .B2(n7694), .A(n7693), .ZN(n7695) );
  INV_X1 U9295 ( .A(n7695), .ZN(P2_U3259) );
  NOR2_X1 U9296 ( .A1(n7760), .A2(n8271), .ZN(n7702) );
  XNOR2_X1 U9297 ( .A(n7700), .B(n6957), .ZN(n7701) );
  NOR2_X1 U9298 ( .A1(n7701), .A2(n7702), .ZN(n7756) );
  AOI21_X1 U9299 ( .B1(n7702), .B2(n7701), .A(n7756), .ZN(n7703) );
  OAI21_X1 U9300 ( .B1(n7704), .B2(n7703), .A(n7758), .ZN(n7705) );
  NAND2_X1 U9301 ( .A1(n7705), .A2(n8611), .ZN(n7712) );
  INV_X1 U9302 ( .A(n7706), .ZN(n7709) );
  OAI22_X1 U9303 ( .A1(n7707), .A2(n8602), .B1(n8603), .B2(n8643), .ZN(n7708)
         );
  AOI211_X1 U9304 ( .C1(n7710), .C2(n8625), .A(n7709), .B(n7708), .ZN(n7711)
         );
  OAI211_X1 U9305 ( .C1(n9900), .C2(n8620), .A(n7712), .B(n7711), .ZN(P2_U3226) );
  NAND2_X1 U9306 ( .A1(n4438), .A2(n7713), .ZN(n7714) );
  XNOR2_X1 U9307 ( .A(n7715), .B(n7714), .ZN(n7723) );
  NAND2_X1 U9308 ( .A1(n9049), .A2(n9503), .ZN(n7720) );
  NAND2_X1 U9309 ( .A1(n9068), .A2(n9497), .ZN(n7719) );
  INV_X1 U9310 ( .A(n9496), .ZN(n7865) );
  OR2_X1 U9311 ( .A1(n9014), .A2(n7865), .ZN(n7718) );
  INV_X1 U9312 ( .A(n7716), .ZN(n7717) );
  NAND4_X1 U9313 ( .A1(n7720), .A2(n7719), .A3(n7718), .A4(n7717), .ZN(n7721)
         );
  AOI21_X1 U9314 ( .B1(n9504), .B2(n9037), .A(n7721), .ZN(n7722) );
  OAI21_X1 U9315 ( .B1(n7723), .B2(n9075), .A(n7722), .ZN(P1_U3215) );
  AND2_X1 U9316 ( .A1(n9786), .A2(n9497), .ZN(n7725) );
  INV_X1 U9317 ( .A(n9082), .ZN(n7821) );
  NAND2_X1 U9318 ( .A1(n9504), .A2(n7821), .ZN(n8320) );
  NAND2_X1 U9319 ( .A1(n8329), .A2(n8320), .ZN(n9494) );
  NAND2_X1 U9320 ( .A1(n9491), .A2(n9494), .ZN(n7728) );
  OR2_X1 U9321 ( .A1(n9504), .A2(n9082), .ZN(n7727) );
  NAND2_X1 U9322 ( .A1(n7728), .A2(n7727), .ZN(n7780) );
  XNOR2_X1 U9323 ( .A(n7782), .B(n9496), .ZN(n8484) );
  INV_X1 U9324 ( .A(n8484), .ZN(n7729) );
  XNOR2_X1 U9325 ( .A(n7780), .B(n7729), .ZN(n9585) );
  AND2_X1 U9326 ( .A1(n8320), .A2(n9492), .ZN(n8330) );
  XNOR2_X1 U9327 ( .A(n7781), .B(n8484), .ZN(n7732) );
  AOI22_X1 U9328 ( .A1(n9713), .A2(n9082), .B1(n9081), .B2(n9711), .ZN(n7731)
         );
  OAI21_X1 U9329 ( .B1(n7732), .B2(n9499), .A(n7731), .ZN(n7733) );
  AOI21_X1 U9330 ( .B1(n9585), .B2(n9502), .A(n7733), .ZN(n9587) );
  INV_X1 U9331 ( .A(n7782), .ZN(n9582) );
  NOR2_X1 U9332 ( .A1(n9506), .A2(n9582), .ZN(n7734) );
  OR2_X1 U9333 ( .A1(n7788), .A2(n7734), .ZN(n9583) );
  AOI22_X1 U9334 ( .A1(n9728), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n7823), .B2(
        n9541), .ZN(n7736) );
  NAND2_X1 U9335 ( .A1(n7782), .A2(n9543), .ZN(n7735) );
  OAI211_X1 U9336 ( .C1(n9583), .C2(n9166), .A(n7736), .B(n7735), .ZN(n7737)
         );
  AOI21_X1 U9337 ( .B1(n9585), .B2(n9510), .A(n7737), .ZN(n7738) );
  OAI21_X1 U9338 ( .B1(n9587), .B2(n9728), .A(n7738), .ZN(P1_U3280) );
  NAND2_X1 U9339 ( .A1(n7739), .A2(n7742), .ZN(n7740) );
  NAND2_X1 U9340 ( .A1(n7741), .A2(n7740), .ZN(n8944) );
  AOI22_X1 U9341 ( .A1(n8645), .A2(n8838), .B1(n8840), .B2(n8642), .ZN(n7746)
         );
  XNOR2_X1 U9342 ( .A(n7743), .B(n7742), .ZN(n7744) );
  NAND2_X1 U9343 ( .A1(n7744), .A2(n8843), .ZN(n7745) );
  OAI211_X1 U9344 ( .C1(n8944), .C2(n7747), .A(n7746), .B(n7745), .ZN(n8946)
         );
  NAND2_X1 U9345 ( .A1(n8946), .A2(n9834), .ZN(n7754) );
  OAI22_X1 U9346 ( .A1(n9834), .A2(n7748), .B1(n7759), .B2(n9825), .ZN(n7752)
         );
  NOR2_X1 U9347 ( .A1(n7749), .A2(n8940), .ZN(n7750) );
  OR2_X1 U9348 ( .A1(n7797), .A2(n7750), .ZN(n8941) );
  NOR2_X1 U9349 ( .A1(n8941), .A2(n8685), .ZN(n7751) );
  AOI211_X1 U9350 ( .C1(n8755), .C2(n7763), .A(n7752), .B(n7751), .ZN(n7753)
         );
  OAI211_X1 U9351 ( .C1(n8944), .C2(n7755), .A(n7754), .B(n7753), .ZN(P2_U3283) );
  INV_X1 U9352 ( .A(n7756), .ZN(n7757) );
  NAND2_X1 U9353 ( .A1(n7758), .A2(n7757), .ZN(n7831) );
  XNOR2_X1 U9354 ( .A(n7763), .B(n8276), .ZN(n7828) );
  NOR2_X1 U9355 ( .A1(n8643), .A2(n8271), .ZN(n7829) );
  XNOR2_X1 U9356 ( .A(n7828), .B(n7829), .ZN(n7830) );
  XNOR2_X1 U9357 ( .A(n7831), .B(n7830), .ZN(n7765) );
  OAI22_X1 U9358 ( .A1(n8615), .A2(n7759), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5990), .ZN(n7762) );
  OAI22_X1 U9359 ( .A1(n7760), .A2(n8602), .B1(n8603), .B2(n7843), .ZN(n7761)
         );
  AOI211_X1 U9360 ( .C1(n7763), .C2(n8629), .A(n7762), .B(n7761), .ZN(n7764)
         );
  OAI21_X1 U9361 ( .B1(n7765), .B2(n8631), .A(n7764), .ZN(P2_U3236) );
  NOR2_X1 U9362 ( .A1(n7767), .A2(n7766), .ZN(n7769) );
  XNOR2_X1 U9363 ( .A(n7883), .B(n7890), .ZN(n7771) );
  INV_X1 U9364 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n7770) );
  NOR2_X1 U9365 ( .A1(n7770), .A2(n7771), .ZN(n7884) );
  AOI211_X1 U9366 ( .C1(n7771), .C2(n7770), .A(n7884), .B(n9659), .ZN(n7778)
         );
  OAI21_X1 U9367 ( .B1(n7773), .B2(P1_REG1_REG_14__SCAN_IN), .A(n7772), .ZN(
        n7889) );
  XNOR2_X1 U9368 ( .A(n7890), .B(n7889), .ZN(n7774) );
  INV_X1 U9369 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9570) );
  NOR2_X1 U9370 ( .A1(n9570), .A2(n7774), .ZN(n7891) );
  AOI211_X1 U9371 ( .C1(n7774), .C2(n9570), .A(n7891), .B(n9636), .ZN(n7777)
         );
  NAND2_X1 U9372 ( .A1(n9668), .A2(P1_ADDR_REG_15__SCAN_IN), .ZN(n7775) );
  NAND2_X1 U9373 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n7997) );
  OAI211_X1 U9374 ( .C1(n7900), .C2(n7890), .A(n7775), .B(n7997), .ZN(n7776)
         );
  OR3_X1 U9375 ( .A1(n7778), .A2(n7777), .A3(n7776), .ZN(P1_U3256) );
  NAND2_X1 U9376 ( .A1(n7782), .A2(n9496), .ZN(n7779) );
  INV_X1 U9377 ( .A(n9081), .ZN(n8018) );
  NAND2_X1 U9378 ( .A1(n7930), .A2(n8018), .ZN(n8412) );
  XNOR2_X1 U9379 ( .A(n7906), .B(n7905), .ZN(n7932) );
  NAND2_X1 U9380 ( .A1(n7782), .A2(n7865), .ZN(n8411) );
  NAND2_X1 U9381 ( .A1(n7781), .A2(n8411), .ZN(n7784) );
  OR2_X1 U9382 ( .A1(n7782), .A2(n7865), .ZN(n7907) );
  NAND2_X1 U9383 ( .A1(n7784), .A2(n7907), .ZN(n7783) );
  INV_X1 U9384 ( .A(n7905), .ZN(n8486) );
  NAND3_X1 U9385 ( .A1(n7784), .A2(n7905), .A3(n7907), .ZN(n7785) );
  NAND3_X1 U9386 ( .A1(n7910), .A2(n9717), .A3(n7785), .ZN(n7787) );
  AOI22_X1 U9387 ( .A1(n9711), .A2(n9080), .B1(n9496), .B2(n9713), .ZN(n7786)
         );
  NAND2_X1 U9388 ( .A1(n7787), .A2(n7786), .ZN(n7928) );
  INV_X1 U9389 ( .A(n7930), .ZN(n7793) );
  INV_X1 U9390 ( .A(n7788), .ZN(n7790) );
  INV_X1 U9391 ( .A(n7916), .ZN(n7789) );
  AOI211_X1 U9392 ( .C1(n7930), .C2(n7790), .A(n9788), .B(n7789), .ZN(n7929)
         );
  NAND2_X1 U9393 ( .A1(n7929), .A2(n9550), .ZN(n7792) );
  AOI22_X1 U9394 ( .A1(n9728), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n7862), .B2(
        n9541), .ZN(n7791) );
  OAI211_X1 U9395 ( .C1(n7793), .C2(n9357), .A(n7792), .B(n7791), .ZN(n7794)
         );
  AOI21_X1 U9396 ( .B1(n7928), .B2(n9725), .A(n7794), .ZN(n7795) );
  OAI21_X1 U9397 ( .B1(n7932), .B2(n9368), .A(n7795), .ZN(P1_U3279) );
  XOR2_X1 U9398 ( .A(n7804), .B(n7796), .Z(n9533) );
  INV_X1 U9399 ( .A(n7797), .ZN(n7799) );
  INV_X1 U9400 ( .A(n7849), .ZN(n7798) );
  AOI21_X1 U9401 ( .B1(n9528), .B2(n7799), .A(n7798), .ZN(n9529) );
  INV_X1 U9402 ( .A(n7837), .ZN(n7800) );
  AOI22_X1 U9403 ( .A1(n9836), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n7800), .B2(
        n8848), .ZN(n7801) );
  OAI21_X1 U9404 ( .B1(n7802), .B2(n8851), .A(n7801), .ZN(n7810) );
  INV_X1 U9405 ( .A(n7803), .ZN(n7805) );
  AOI21_X1 U9406 ( .B1(n7805), .B2(n4755), .A(n8825), .ZN(n7808) );
  OR2_X1 U9407 ( .A1(n8643), .A2(n8828), .ZN(n7806) );
  OAI21_X1 U9408 ( .B1(n8120), .B2(n8830), .A(n7806), .ZN(n7834) );
  AOI21_X1 U9409 ( .B1(n7808), .B2(n7807), .A(n7834), .ZN(n9531) );
  NOR2_X1 U9410 ( .A1(n9531), .A2(n9836), .ZN(n7809) );
  AOI211_X1 U9411 ( .C1(n9529), .C2(n8858), .A(n7810), .B(n7809), .ZN(n7811)
         );
  OAI21_X1 U9412 ( .B1(n9533), .B2(n8855), .A(n7811), .ZN(P2_U3282) );
  INV_X1 U9413 ( .A(n7812), .ZN(n7815) );
  OAI222_X1 U9414 ( .A1(n8242), .A2(n10075), .B1(n8973), .B2(n7815), .C1(
        P2_U3152), .C2(n7813), .ZN(P2_U3333) );
  OAI222_X1 U9415 ( .A1(n8557), .A2(n7816), .B1(n4370), .B2(n7815), .C1(n7814), 
        .C2(P1_U3084), .ZN(P1_U3328) );
  INV_X1 U9416 ( .A(n9073), .ZN(n9063) );
  OAI211_X1 U9417 ( .C1(n4442), .C2(n7819), .A(n7818), .B(n5747), .ZN(n7825)
         );
  AND2_X1 U9418 ( .A1(P1_U3084), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n9671) );
  AOI21_X1 U9419 ( .B1(n9067), .B2(n9081), .A(n9671), .ZN(n7820) );
  OAI21_X1 U9420 ( .B1(n7821), .B2(n9058), .A(n7820), .ZN(n7822) );
  AOI21_X1 U9421 ( .B1(n7823), .B2(n9049), .A(n7822), .ZN(n7824) );
  OAI211_X1 U9422 ( .C1(n9582), .C2(n9063), .A(n7825), .B(n7824), .ZN(P1_U3234) );
  XNOR2_X1 U9423 ( .A(n9528), .B(n8247), .ZN(n7827) );
  NAND2_X1 U9424 ( .A1(n8642), .A2(n8274), .ZN(n7826) );
  NAND2_X1 U9425 ( .A1(n7827), .A2(n7826), .ZN(n8036) );
  OAI21_X1 U9426 ( .B1(n7827), .B2(n7826), .A(n8036), .ZN(n7833) );
  AOI21_X1 U9427 ( .B1(n7833), .B2(n7832), .A(n4435), .ZN(n7840) );
  INV_X1 U9428 ( .A(n8627), .ZN(n8617) );
  NAND2_X1 U9429 ( .A1(n8617), .A2(n7834), .ZN(n7836) );
  OAI211_X1 U9430 ( .C1(n8615), .C2(n7837), .A(n7836), .B(n7835), .ZN(n7838)
         );
  AOI21_X1 U9431 ( .B1(n9528), .B2(n8629), .A(n7838), .ZN(n7839) );
  OAI21_X1 U9432 ( .B1(n7840), .B2(n8631), .A(n7839), .ZN(P2_U3217) );
  XNOR2_X1 U9433 ( .A(n7842), .B(n7841), .ZN(n7845) );
  OAI22_X1 U9434 ( .A1(n8073), .A2(n8830), .B1(n7843), .B2(n8828), .ZN(n8039)
         );
  INV_X1 U9435 ( .A(n8039), .ZN(n7844) );
  OAI21_X1 U9436 ( .B1(n7845), .B2(n8825), .A(n7844), .ZN(n9523) );
  INV_X1 U9437 ( .A(n9523), .ZN(n7856) );
  OAI21_X1 U9438 ( .B1(n7848), .B2(n7847), .A(n7846), .ZN(n9525) );
  NAND2_X1 U9439 ( .A1(n7849), .A2(n9521), .ZN(n7850) );
  NAND2_X1 U9440 ( .A1(n7950), .A2(n7850), .ZN(n9522) );
  OAI22_X1 U9441 ( .A1(n9834), .A2(n7851), .B1(n8042), .B2(n9825), .ZN(n7852)
         );
  AOI21_X1 U9442 ( .B1(n9521), .B2(n8755), .A(n7852), .ZN(n7853) );
  OAI21_X1 U9443 ( .B1(n9522), .B2(n8685), .A(n7853), .ZN(n7854) );
  AOI21_X1 U9444 ( .B1(n9525), .B2(n8813), .A(n7854), .ZN(n7855) );
  OAI21_X1 U9445 ( .B1(n9836), .B2(n7856), .A(n7855), .ZN(P2_U3281) );
  NAND2_X1 U9446 ( .A1(n7818), .A2(n7857), .ZN(n8005) );
  XNOR2_X1 U9447 ( .A(n7859), .B(n7858), .ZN(n7860) );
  XNOR2_X1 U9448 ( .A(n8005), .B(n7860), .ZN(n7868) );
  AOI21_X1 U9449 ( .B1(n9067), .B2(n9080), .A(n7861), .ZN(n7864) );
  NAND2_X1 U9450 ( .A1(n9049), .A2(n7862), .ZN(n7863) );
  OAI211_X1 U9451 ( .C1(n7865), .C2(n9058), .A(n7864), .B(n7863), .ZN(n7866)
         );
  AOI21_X1 U9452 ( .B1(n7930), .B2(n9037), .A(n7866), .ZN(n7867) );
  OAI21_X1 U9453 ( .B1(n7868), .B2(n9075), .A(n7867), .ZN(P1_U3222) );
  XNOR2_X1 U9454 ( .A(n7874), .B(n8086), .ZN(n7870) );
  NAND2_X1 U9455 ( .A1(n7870), .A2(n7851), .ZN(n8088) );
  OAI21_X1 U9456 ( .B1(n7870), .B2(n7851), .A(n8088), .ZN(n7881) );
  NOR2_X1 U9457 ( .A1(n9809), .A2(n8087), .ZN(n7880) );
  INV_X1 U9458 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n10161) );
  OAI21_X1 U9459 ( .B1(n7872), .B2(P2_REG1_REG_14__SCAN_IN), .A(n7871), .ZN(
        n8080) );
  INV_X1 U9460 ( .A(n8080), .ZN(n7873) );
  XNOR2_X1 U9461 ( .A(n7874), .B(n7873), .ZN(n7875) );
  NAND2_X1 U9462 ( .A1(n7875), .A2(n6008), .ZN(n7877) );
  NOR2_X1 U9463 ( .A1(n6008), .A2(n7875), .ZN(n8081) );
  INV_X1 U9464 ( .A(n8081), .ZN(n7876) );
  NAND3_X1 U9465 ( .A1(n9807), .A2(n7877), .A3(n7876), .ZN(n7878) );
  NAND2_X1 U9466 ( .A1(P2_U3152), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8040) );
  OAI211_X1 U9467 ( .C1(n10161), .C2(n8675), .A(n7878), .B(n8040), .ZN(n7879)
         );
  AOI211_X1 U9468 ( .C1(n7881), .C2(n9808), .A(n7880), .B(n7879), .ZN(n7882)
         );
  INV_X1 U9469 ( .A(n7882), .ZN(P2_U3260) );
  NOR2_X1 U9470 ( .A1(n7883), .A2(n7890), .ZN(n7885) );
  NOR2_X1 U9471 ( .A1(n7885), .A2(n7884), .ZN(n7888) );
  NAND2_X1 U9472 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n8103), .ZN(n7886) );
  OAI21_X1 U9473 ( .B1(n8103), .B2(P1_REG2_REG_16__SCAN_IN), .A(n7886), .ZN(
        n7887) );
  NOR2_X1 U9474 ( .A1(n7888), .A2(n7887), .ZN(n8096) );
  AOI211_X1 U9475 ( .C1(n7888), .C2(n7887), .A(n8096), .B(n9659), .ZN(n7903)
         );
  NOR2_X1 U9476 ( .A1(n7890), .A2(n7889), .ZN(n7892) );
  NOR2_X1 U9477 ( .A1(n7892), .A2(n7891), .ZN(n7895) );
  INV_X1 U9478 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n7893) );
  MUX2_X1 U9479 ( .A(n7893), .B(P1_REG1_REG_16__SCAN_IN), .S(n8103), .Z(n7894)
         );
  NOR2_X1 U9480 ( .A1(n7895), .A2(n7894), .ZN(n8102) );
  AOI211_X1 U9481 ( .C1(n7895), .C2(n7894), .A(n8102), .B(n9636), .ZN(n7902)
         );
  NAND2_X1 U9482 ( .A1(n9668), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n7898) );
  NOR2_X1 U9483 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7896), .ZN(n8144) );
  INV_X1 U9484 ( .A(n8144), .ZN(n7897) );
  OAI211_X1 U9485 ( .C1(n7900), .C2(n7899), .A(n7898), .B(n7897), .ZN(n7901)
         );
  OR3_X1 U9486 ( .A1(n7903), .A2(n7902), .A3(n7901), .ZN(P1_U3257) );
  AND2_X1 U9487 ( .A1(n7930), .A2(n9081), .ZN(n7904) );
  OR2_X1 U9488 ( .A1(n7959), .A2(n7988), .ZN(n8340) );
  NAND2_X1 U9489 ( .A1(n7959), .A2(n7988), .ZN(n8334) );
  NAND2_X1 U9490 ( .A1(n8340), .A2(n8334), .ZN(n8483) );
  XNOR2_X1 U9491 ( .A(n7958), .B(n8483), .ZN(n9579) );
  INV_X1 U9492 ( .A(n7907), .ZN(n7908) );
  NAND2_X1 U9493 ( .A1(n8412), .A2(n7908), .ZN(n7909) );
  AND2_X1 U9494 ( .A1(n7909), .A2(n8335), .ZN(n8333) );
  AND2_X1 U9495 ( .A1(n7911), .A2(n8483), .ZN(n7912) );
  OAI21_X1 U9496 ( .B1(n4431), .B2(n7912), .A(n9717), .ZN(n7914) );
  AOI22_X1 U9497 ( .A1(n9713), .A2(n9081), .B1(n9079), .B2(n9711), .ZN(n7913)
         );
  NAND2_X1 U9498 ( .A1(n7914), .A2(n7913), .ZN(n7915) );
  AOI21_X1 U9499 ( .B1(n9579), .B2(n9502), .A(n7915), .ZN(n9581) );
  NAND2_X1 U9500 ( .A1(n7916), .A2(n7959), .ZN(n7917) );
  NAND2_X1 U9501 ( .A1(n7966), .A2(n7917), .ZN(n9577) );
  AOI22_X1 U9502 ( .A1(n9728), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n8020), .B2(
        n9541), .ZN(n7919) );
  NAND2_X1 U9503 ( .A1(n7959), .A2(n9543), .ZN(n7918) );
  OAI211_X1 U9504 ( .C1(n9577), .C2(n9166), .A(n7919), .B(n7918), .ZN(n7920)
         );
  AOI21_X1 U9505 ( .B1(n9579), .B2(n9510), .A(n7920), .ZN(n7921) );
  OAI21_X1 U9506 ( .B1(n9581), .B2(n9728), .A(n7921), .ZN(P1_U3278) );
  INV_X1 U9507 ( .A(n7922), .ZN(n7926) );
  OAI222_X1 U9508 ( .A1(n8242), .A2(n7924), .B1(n8973), .B2(n7926), .C1(
        P2_U3152), .C2(n7923), .ZN(P2_U3332) );
  OAI222_X1 U9509 ( .A1(n8557), .A2(n7927), .B1(n4370), .B2(n7926), .C1(n7925), 
        .C2(P1_U3084), .ZN(P1_U3327) );
  AOI211_X1 U9510 ( .C1(n9436), .C2(n7930), .A(n7929), .B(n7928), .ZN(n7931)
         );
  OAI21_X1 U9511 ( .B1(n7932), .B2(n9440), .A(n7931), .ZN(n7934) );
  NAND2_X1 U9512 ( .A1(n7934), .A2(n9806), .ZN(n7933) );
  OAI21_X1 U9513 ( .B1(n9806), .B2(n6839), .A(n7933), .ZN(P1_U3535) );
  INV_X1 U9514 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n7936) );
  NAND2_X1 U9515 ( .A1(n7934), .A2(n9795), .ZN(n7935) );
  OAI21_X1 U9516 ( .B1(n9795), .B2(n7936), .A(n7935), .ZN(P1_U3490) );
  NAND2_X1 U9517 ( .A1(n7940), .A2(n7974), .ZN(n7938) );
  OAI211_X1 U9518 ( .C1(n8557), .C2(n7939), .A(n7938), .B(n7937), .ZN(P1_U3326) );
  INV_X1 U9519 ( .A(n7940), .ZN(n7942) );
  OAI222_X1 U9520 ( .A1(n8242), .A2(n7943), .B1(n8973), .B2(n7942), .C1(n7941), 
        .C2(P2_U3152), .ZN(P2_U3331) );
  XNOR2_X1 U9521 ( .A(n7945), .B(n7944), .ZN(n7946) );
  OAI222_X1 U9522 ( .A1(n8830), .A2(n8132), .B1(n8828), .B2(n8120), .C1(n7946), 
        .C2(n8825), .ZN(n8936) );
  INV_X1 U9523 ( .A(n8936), .ZN(n7957) );
  AOI21_X1 U9524 ( .B1(n7949), .B2(n7948), .A(n7947), .ZN(n8938) );
  AND2_X1 U9525 ( .A1(n8111), .A2(n7950), .ZN(n7951) );
  OR2_X1 U9526 ( .A1(n7951), .A2(n8023), .ZN(n8935) );
  OAI22_X1 U9527 ( .A1(n9834), .A2(n7952), .B1(n8119), .B2(n9825), .ZN(n7953)
         );
  AOI21_X1 U9528 ( .B1(n8111), .B2(n8755), .A(n7953), .ZN(n7954) );
  OAI21_X1 U9529 ( .B1(n8935), .B2(n8685), .A(n7954), .ZN(n7955) );
  AOI21_X1 U9530 ( .B1(n8938), .B2(n8813), .A(n7955), .ZN(n7956) );
  OAI21_X1 U9531 ( .B1(n9836), .B2(n7957), .A(n7956), .ZN(P2_U3280) );
  INV_X1 U9532 ( .A(n7959), .ZN(n9576) );
  NAND2_X1 U9533 ( .A1(n8048), .A2(n8052), .ZN(n8341) );
  XOR2_X1 U9534 ( .A(n8046), .B(n8487), .Z(n9575) );
  INV_X1 U9535 ( .A(n9575), .ZN(n7973) );
  INV_X1 U9536 ( .A(n8334), .ZN(n7961) );
  OR2_X1 U9537 ( .A1(n4431), .A2(n7961), .ZN(n7962) );
  XNOR2_X1 U9538 ( .A(n7962), .B(n8487), .ZN(n7963) );
  NAND2_X1 U9539 ( .A1(n7963), .A2(n9717), .ZN(n7965) );
  AOI22_X1 U9540 ( .A1(n9713), .A2(n9080), .B1(n9538), .B2(n9711), .ZN(n7964)
         );
  NAND2_X1 U9541 ( .A1(n7965), .A2(n7964), .ZN(n9574) );
  INV_X1 U9542 ( .A(n8048), .ZN(n9572) );
  INV_X1 U9543 ( .A(n7966), .ZN(n7967) );
  OAI211_X1 U9544 ( .C1(n9572), .C2(n7967), .A(n4534), .B(n9704), .ZN(n9571)
         );
  INV_X1 U9545 ( .A(n9550), .ZN(n7970) );
  AOI22_X1 U9546 ( .A1(n9728), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n7990), .B2(
        n9541), .ZN(n7969) );
  NAND2_X1 U9547 ( .A1(n8048), .A2(n9543), .ZN(n7968) );
  OAI211_X1 U9548 ( .C1(n9571), .C2(n7970), .A(n7969), .B(n7968), .ZN(n7971)
         );
  AOI21_X1 U9549 ( .B1(n9574), .B2(n9725), .A(n7971), .ZN(n7972) );
  OAI21_X1 U9550 ( .B1(n7973), .B2(n9368), .A(n7972), .ZN(P1_U3277) );
  NAND2_X1 U9551 ( .A1(n6484), .A2(n7974), .ZN(n7976) );
  OAI211_X1 U9552 ( .C1(n8557), .C2(n7977), .A(n7976), .B(n7975), .ZN(P1_U3325) );
  INV_X1 U9553 ( .A(n7983), .ZN(n7986) );
  AND2_X1 U9554 ( .A1(n7980), .A2(n7979), .ZN(n7982) );
  AOI21_X1 U9555 ( .B1(n7983), .B2(n7982), .A(n7981), .ZN(n7984) );
  NOR2_X1 U9556 ( .A1(n7984), .A2(n9075), .ZN(n7985) );
  OAI21_X1 U9557 ( .B1(n7986), .B2(n7978), .A(n7985), .ZN(n7992) );
  AOI22_X1 U9558 ( .A1(n9067), .A2(n9538), .B1(P1_REG3_REG_14__SCAN_IN), .B2(
        P1_U3084), .ZN(n7987) );
  OAI21_X1 U9559 ( .B1(n7988), .B2(n9058), .A(n7987), .ZN(n7989) );
  AOI21_X1 U9560 ( .B1(n7990), .B2(n9049), .A(n7989), .ZN(n7991) );
  OAI211_X1 U9561 ( .C1(n9572), .C2(n9063), .A(n7992), .B(n7991), .ZN(P1_U3213) );
  NAND2_X1 U9562 ( .A1(n7994), .A2(n7993), .ZN(n7995) );
  XOR2_X1 U9563 ( .A(n7996), .B(n7995), .Z(n8003) );
  INV_X1 U9564 ( .A(n7997), .ZN(n7998) );
  AOI21_X1 U9565 ( .B1(n9067), .B2(n9361), .A(n7998), .ZN(n8000) );
  NAND2_X1 U9566 ( .A1(n9049), .A2(n8054), .ZN(n7999) );
  OAI211_X1 U9567 ( .C1(n8052), .C2(n9058), .A(n8000), .B(n7999), .ZN(n8001)
         );
  AOI21_X1 U9568 ( .B1(n9117), .B2(n9073), .A(n8001), .ZN(n8002) );
  OAI21_X1 U9569 ( .B1(n8003), .B2(n9075), .A(n8002), .ZN(P1_U3239) );
  NAND2_X1 U9570 ( .A1(n8005), .A2(n8004), .ZN(n8007) );
  NAND2_X1 U9571 ( .A1(n8007), .A2(n8006), .ZN(n8009) );
  OR2_X1 U9572 ( .A1(n8009), .A2(n8010), .ZN(n8013) );
  INV_X1 U9573 ( .A(n8008), .ZN(n8012) );
  OAI21_X1 U9574 ( .B1(n8010), .B2(n8012), .A(n8009), .ZN(n8011) );
  OAI21_X1 U9575 ( .B1(n8013), .B2(n8012), .A(n8011), .ZN(n8014) );
  NAND2_X1 U9576 ( .A1(n8014), .A2(n5747), .ZN(n8022) );
  INV_X1 U9577 ( .A(n8015), .ZN(n8016) );
  AOI21_X1 U9578 ( .B1(n9067), .B2(n9079), .A(n8016), .ZN(n8017) );
  OAI21_X1 U9579 ( .B1(n8018), .B2(n9058), .A(n8017), .ZN(n8019) );
  AOI21_X1 U9580 ( .B1(n8020), .B2(n9049), .A(n8019), .ZN(n8021) );
  OAI211_X1 U9581 ( .C1(n9576), .C2(n9063), .A(n8022), .B(n8021), .ZN(P1_U3232) );
  INV_X1 U9582 ( .A(n8023), .ZN(n8025) );
  INV_X1 U9583 ( .A(n8846), .ZN(n8024) );
  AOI211_X1 U9584 ( .C1(n8930), .C2(n8025), .A(n9901), .B(n8024), .ZN(n8929)
         );
  XNOR2_X1 U9585 ( .A(n8026), .B(n8030), .ZN(n8027) );
  AOI222_X1 U9586 ( .A1(n8843), .A2(n8027), .B1(n8639), .B2(n8840), .C1(n8640), 
        .C2(n8838), .ZN(n8932) );
  INV_X1 U9587 ( .A(n8932), .ZN(n8028) );
  AOI21_X1 U9588 ( .B1(n8929), .B2(n9827), .A(n8028), .ZN(n8035) );
  OAI21_X1 U9589 ( .B1(n8031), .B2(n8030), .A(n8029), .ZN(n8928) );
  AOI22_X1 U9590 ( .A1(n9836), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n8070), .B2(
        n8848), .ZN(n8032) );
  OAI21_X1 U9591 ( .B1(n6439), .B2(n8851), .A(n8032), .ZN(n8033) );
  AOI21_X1 U9592 ( .B1(n8928), .B2(n8813), .A(n8033), .ZN(n8034) );
  OAI21_X1 U9593 ( .B1(n8035), .B2(n9836), .A(n8034), .ZN(P2_U3279) );
  NOR2_X1 U9594 ( .A1(n8120), .A2(n8271), .ZN(n8062) );
  INV_X1 U9595 ( .A(n8036), .ZN(n8037) );
  XNOR2_X1 U9596 ( .A(n9521), .B(n8276), .ZN(n8060) );
  INV_X1 U9597 ( .A(n8060), .ZN(n8061) );
  NAND2_X1 U9598 ( .A1(n4430), .A2(n8061), .ZN(n8112) );
  OAI21_X1 U9599 ( .B1(n4430), .B2(n8061), .A(n8112), .ZN(n8038) );
  NOR2_X1 U9600 ( .A1(n8038), .A2(n8062), .ZN(n8115) );
  AOI21_X1 U9601 ( .B1(n8062), .B2(n8038), .A(n8115), .ZN(n8045) );
  NAND2_X1 U9602 ( .A1(n8617), .A2(n8039), .ZN(n8041) );
  OAI211_X1 U9603 ( .C1(n8615), .C2(n8042), .A(n8041), .B(n8040), .ZN(n8043)
         );
  AOI21_X1 U9604 ( .B1(n9521), .B2(n8629), .A(n8043), .ZN(n8044) );
  OAI21_X1 U9605 ( .B1(n8045), .B2(n8631), .A(n8044), .ZN(P2_U3243) );
  OAI21_X1 U9606 ( .B1(n9572), .B2(n8052), .A(n8046), .ZN(n8047) );
  OAI21_X1 U9607 ( .B1(n9079), .B2(n8048), .A(n8047), .ZN(n9115) );
  INV_X1 U9608 ( .A(n9538), .ZN(n9116) );
  OR2_X1 U9609 ( .A1(n9117), .A2(n9116), .ZN(n8421) );
  NAND2_X1 U9610 ( .A1(n9117), .A2(n9116), .ZN(n9534) );
  NAND2_X1 U9611 ( .A1(n8421), .A2(n9534), .ZN(n8489) );
  XNOR2_X1 U9612 ( .A(n9115), .B(n8489), .ZN(n9569) );
  INV_X1 U9613 ( .A(n9569), .ZN(n8059) );
  INV_X1 U9614 ( .A(n9361), .ZN(n8306) );
  NAND2_X1 U9615 ( .A1(n8487), .A2(n8334), .ZN(n8049) );
  AOI21_X1 U9616 ( .B1(n8489), .B2(n8050), .A(n9138), .ZN(n8051) );
  OAI222_X1 U9617 ( .A1(n9348), .A2(n8306), .B1(n9346), .B2(n8052), .C1(n9499), 
        .C2(n8051), .ZN(n9567) );
  OAI21_X1 U9618 ( .B1(n8053), .B2(n9565), .A(n9547), .ZN(n9566) );
  AOI22_X1 U9619 ( .A1(n9728), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n8054), .B2(
        n9541), .ZN(n8056) );
  NAND2_X1 U9620 ( .A1(n9117), .A2(n9543), .ZN(n8055) );
  OAI211_X1 U9621 ( .C1(n9566), .C2(n9166), .A(n8056), .B(n8055), .ZN(n8057)
         );
  AOI21_X1 U9622 ( .B1(n9567), .B2(n9725), .A(n8057), .ZN(n8058) );
  OAI21_X1 U9623 ( .B1(n8059), .B2(n9368), .A(n8058), .ZN(P1_U3276) );
  XNOR2_X1 U9624 ( .A(n8111), .B(n6957), .ZN(n8068) );
  NAND2_X1 U9625 ( .A1(n8640), .A2(n8274), .ZN(n8066) );
  XNOR2_X1 U9626 ( .A(n8068), .B(n8066), .ZN(n8113) );
  NAND2_X1 U9627 ( .A1(n8060), .A2(n8062), .ZN(n8063) );
  NAND2_X1 U9628 ( .A1(n8065), .A2(n8064), .ZN(n8116) );
  INV_X1 U9629 ( .A(n8066), .ZN(n8067) );
  XNOR2_X1 U9630 ( .A(n8930), .B(n8276), .ZN(n8126) );
  NOR2_X1 U9631 ( .A1(n8132), .A2(n8271), .ZN(n8127) );
  XNOR2_X1 U9632 ( .A(n8126), .B(n8127), .ZN(n8130) );
  XNOR2_X1 U9633 ( .A(n8131), .B(n8130), .ZN(n8077) );
  INV_X1 U9634 ( .A(n8070), .ZN(n8072) );
  OAI22_X1 U9635 ( .A1(n8615), .A2(n8072), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8071), .ZN(n8075) );
  OAI22_X1 U9636 ( .A1(n8073), .A2(n8602), .B1(n8603), .B2(n8179), .ZN(n8074)
         );
  AOI211_X1 U9637 ( .C1(n8930), .C2(n8629), .A(n8075), .B(n8074), .ZN(n8076)
         );
  OAI21_X1 U9638 ( .B1(n8077), .B2(n8631), .A(n8076), .ZN(P2_U3230) );
  INV_X1 U9639 ( .A(n8390), .ZN(n8110) );
  AOI22_X1 U9640 ( .A1(n8078), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n8970), .ZN(n8079) );
  OAI21_X1 U9641 ( .B1(n8110), .B2(n8973), .A(n8079), .ZN(P2_U3329) );
  NOR2_X1 U9642 ( .A1(n8087), .A2(n8080), .ZN(n8082) );
  NOR2_X1 U9643 ( .A1(n8082), .A2(n8081), .ZN(n8084) );
  XNOR2_X1 U9644 ( .A(n8221), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n8083) );
  NAND2_X1 U9645 ( .A1(n8083), .A2(n8084), .ZN(n8222) );
  OAI21_X1 U9646 ( .B1(n8084), .B2(n8083), .A(n8222), .ZN(n8094) );
  NOR2_X1 U9647 ( .A1(n10197), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8122) );
  AOI21_X1 U9648 ( .B1(n9813), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n8122), .ZN(
        n8085) );
  OAI21_X1 U9649 ( .B1(n9809), .B2(n8221), .A(n8085), .ZN(n8093) );
  NAND2_X1 U9650 ( .A1(n8087), .A2(n8086), .ZN(n8089) );
  NAND2_X1 U9651 ( .A1(n8089), .A2(n8088), .ZN(n8091) );
  AOI22_X1 U9652 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n8221), .B1(n8227), .B2(
        n7952), .ZN(n8090) );
  AOI211_X1 U9653 ( .C1(n8091), .C2(n8090), .A(n8226), .B(n8657), .ZN(n8092)
         );
  AOI211_X1 U9654 ( .C1(n9807), .C2(n8094), .A(n8093), .B(n8092), .ZN(n8095)
         );
  INV_X1 U9655 ( .A(n8095), .ZN(P2_U3261) );
  AND2_X1 U9656 ( .A1(P1_REG3_REG_17__SCAN_IN), .A2(P1_U3084), .ZN(n8101) );
  AOI21_X1 U9657 ( .B1(n8103), .B2(P1_REG2_REG_16__SCAN_IN), .A(n8096), .ZN(
        n8099) );
  NAND2_X1 U9658 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(n9095), .ZN(n8097) );
  OAI21_X1 U9659 ( .B1(n9095), .B2(P1_REG2_REG_17__SCAN_IN), .A(n8097), .ZN(
        n8098) );
  NOR2_X1 U9660 ( .A1(n8099), .A2(n8098), .ZN(n9090) );
  AOI211_X1 U9661 ( .C1(n8099), .C2(n8098), .A(n9090), .B(n9659), .ZN(n8100)
         );
  AOI211_X1 U9662 ( .C1(n9686), .C2(n9095), .A(n8101), .B(n8100), .ZN(n8108)
         );
  XNOR2_X1 U9663 ( .A(n9095), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n8105) );
  AOI21_X1 U9664 ( .B1(n8103), .B2(P1_REG1_REG_16__SCAN_IN), .A(n8102), .ZN(
        n8104) );
  NOR2_X1 U9665 ( .A1(n8104), .A2(n8105), .ZN(n9094) );
  AOI211_X1 U9666 ( .C1(n8105), .C2(n8104), .A(n9094), .B(n9636), .ZN(n8106)
         );
  AOI21_X1 U9667 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(n9668), .A(n8106), .ZN(
        n8107) );
  NAND2_X1 U9668 ( .A1(n8108), .A2(n8107), .ZN(P1_U3258) );
  OAI222_X1 U9669 ( .A1(n4370), .A2(n8110), .B1(n8109), .B2(P1_U3084), .C1(
        n10023), .C2(n8557), .ZN(P1_U3324) );
  INV_X1 U9670 ( .A(n8111), .ZN(n8934) );
  INV_X1 U9671 ( .A(n8112), .ZN(n8114) );
  NOR3_X1 U9672 ( .A1(n8115), .A2(n8114), .A3(n8113), .ZN(n8118) );
  INV_X1 U9673 ( .A(n8116), .ZN(n8117) );
  OAI21_X1 U9674 ( .B1(n8118), .B2(n8117), .A(n8611), .ZN(n8125) );
  INV_X1 U9675 ( .A(n8119), .ZN(n8123) );
  OAI22_X1 U9676 ( .A1(n8120), .A2(n8602), .B1(n8603), .B2(n8132), .ZN(n8121)
         );
  AOI211_X1 U9677 ( .C1(n8625), .C2(n8123), .A(n8122), .B(n8121), .ZN(n8124)
         );
  OAI211_X1 U9678 ( .C1(n8934), .C2(n8620), .A(n8125), .B(n8124), .ZN(P2_U3228) );
  INV_X1 U9679 ( .A(n8126), .ZN(n8129) );
  INV_X1 U9680 ( .A(n8127), .ZN(n8128) );
  NOR2_X1 U9681 ( .A1(n8179), .A2(n8271), .ZN(n8168) );
  XNOR2_X1 U9682 ( .A(n8923), .B(n8276), .ZN(n8169) );
  XOR2_X1 U9683 ( .A(n8168), .B(n8169), .Z(n8171) );
  XNOR2_X1 U9684 ( .A(n8172), .B(n8171), .ZN(n8136) );
  NAND2_X1 U9685 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8674) );
  OAI21_X1 U9686 ( .B1(n8615), .B2(n8847), .A(n8674), .ZN(n8134) );
  OAI22_X1 U9687 ( .A1(n8132), .A2(n8602), .B1(n8603), .B2(n8829), .ZN(n8133)
         );
  AOI211_X1 U9688 ( .C1(n8923), .C2(n8629), .A(n8134), .B(n8133), .ZN(n8135)
         );
  OAI21_X1 U9689 ( .B1(n8136), .B2(n8631), .A(n8135), .ZN(P2_U3240) );
  INV_X1 U9690 ( .A(n9544), .ZN(n9562) );
  INV_X1 U9691 ( .A(n8137), .ZN(n8141) );
  OAI21_X1 U9692 ( .B1(n8139), .B2(n8141), .A(n8138), .ZN(n8140) );
  OAI21_X1 U9693 ( .B1(n8142), .B2(n8141), .A(n8140), .ZN(n8143) );
  NAND2_X1 U9694 ( .A1(n8143), .A2(n5747), .ZN(n8148) );
  AOI21_X1 U9695 ( .B1(n9067), .B2(n9539), .A(n8144), .ZN(n8145) );
  OAI21_X1 U9696 ( .B1(n9116), .B2(n9058), .A(n8145), .ZN(n8146) );
  AOI21_X1 U9697 ( .B1(n9542), .B2(n9049), .A(n8146), .ZN(n8147) );
  OAI211_X1 U9698 ( .C1(n9562), .C2(n9063), .A(n8148), .B(n8147), .ZN(P1_U3224) );
  XNOR2_X1 U9699 ( .A(n8150), .B(n8149), .ZN(n8922) );
  AOI22_X1 U9700 ( .A1(n8920), .A2(n8755), .B1(n9836), .B2(
        P2_REG2_REG_19__SCAN_IN), .ZN(n8158) );
  XNOR2_X1 U9701 ( .A(n8152), .B(n8151), .ZN(n8153) );
  OAI222_X1 U9702 ( .A1(n8830), .A2(n8579), .B1(n8828), .B2(n8179), .C1(n8825), 
        .C2(n8153), .ZN(n8918) );
  AOI211_X1 U9703 ( .C1(n8920), .C2(n8844), .A(n9901), .B(n8817), .ZN(n8919)
         );
  INV_X1 U9704 ( .A(n8919), .ZN(n8155) );
  INV_X1 U9705 ( .A(n8181), .ZN(n8154) );
  OAI22_X1 U9706 ( .A1(n8155), .A2(n8734), .B1(n9825), .B2(n8154), .ZN(n8156)
         );
  OAI21_X1 U9707 ( .B1(n8918), .B2(n8156), .A(n9834), .ZN(n8157) );
  OAI211_X1 U9708 ( .C1(n8922), .C2(n8855), .A(n8158), .B(n8157), .ZN(P2_U3277) );
  INV_X1 U9709 ( .A(n9435), .ZN(n9358) );
  OAI21_X1 U9710 ( .B1(n8161), .B2(n8160), .A(n8159), .ZN(n8162) );
  NAND2_X1 U9711 ( .A1(n8162), .A2(n5747), .ZN(n8167) );
  INV_X1 U9712 ( .A(n8163), .ZN(n9355) );
  INV_X1 U9713 ( .A(n9362), .ZN(n8991) );
  AOI22_X1 U9714 ( .A1(n9068), .A2(n9361), .B1(P1_REG3_REG_17__SCAN_IN), .B2(
        P1_U3084), .ZN(n8164) );
  OAI21_X1 U9715 ( .B1(n8991), .B2(n9014), .A(n8164), .ZN(n8165) );
  AOI21_X1 U9716 ( .B1(n9355), .B2(n9049), .A(n8165), .ZN(n8166) );
  OAI211_X1 U9717 ( .C1(n9358), .C2(n9063), .A(n8167), .B(n8166), .ZN(P1_U3226) );
  NOR2_X1 U9718 ( .A1(n8829), .A2(n8271), .ZN(n8174) );
  XNOR2_X1 U9719 ( .A(n8920), .B(n8276), .ZN(n8173) );
  AOI21_X1 U9720 ( .B1(n8174), .B2(n8173), .A(n8243), .ZN(n8175) );
  NOR2_X1 U9721 ( .A1(n8176), .A2(n8175), .ZN(n8177) );
  OAI21_X1 U9722 ( .B1(n8177), .B2(n8244), .A(n8611), .ZN(n8183) );
  NOR2_X1 U9723 ( .A1(n8178), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8239) );
  OAI22_X1 U9724 ( .A1(n8179), .A2(n8602), .B1(n8603), .B2(n8579), .ZN(n8180)
         );
  AOI211_X1 U9725 ( .C1(n8625), .C2(n8181), .A(n8239), .B(n8180), .ZN(n8182)
         );
  OAI211_X1 U9726 ( .C1(n8184), .C2(n8620), .A(n8183), .B(n8182), .ZN(P2_U3221) );
  NAND2_X1 U9727 ( .A1(n8186), .A2(n8185), .ZN(n8188) );
  INV_X1 U9728 ( .A(n8189), .ZN(n8187) );
  XNOR2_X1 U9729 ( .A(n8188), .B(n8187), .ZN(n8195) );
  OR2_X1 U9730 ( .A1(n8190), .A2(n8189), .ZN(n8192) );
  NAND2_X1 U9731 ( .A1(n8192), .A2(n8191), .ZN(n9771) );
  NAND2_X1 U9732 ( .A1(n9771), .A2(n9502), .ZN(n8194) );
  AOI22_X1 U9733 ( .A1(n9713), .A2(n9088), .B1(n9086), .B2(n9711), .ZN(n8193)
         );
  OAI211_X1 U9734 ( .C1(n9499), .C2(n8195), .A(n8194), .B(n8193), .ZN(n9769)
         );
  MUX2_X1 U9735 ( .A(n9769), .B(P1_REG2_REG_4__SCAN_IN), .S(n9728), .Z(n8202)
         );
  OR2_X1 U9736 ( .A1(n8196), .A2(n9767), .ZN(n8197) );
  NAND2_X1 U9737 ( .A1(n8198), .A2(n8197), .ZN(n9768) );
  NAND2_X1 U9738 ( .A1(n9771), .A2(n9510), .ZN(n8200) );
  AOI22_X1 U9739 ( .A1(n9543), .A2(n9022), .B1(n9023), .B2(n9541), .ZN(n8199)
         );
  OAI211_X1 U9740 ( .C1(n9166), .C2(n9768), .A(n8200), .B(n8199), .ZN(n8201)
         );
  OR2_X1 U9741 ( .A1(n8202), .A2(n8201), .ZN(P1_U3287) );
  INV_X1 U9742 ( .A(n8203), .ZN(n8204) );
  NOR2_X1 U9743 ( .A1(n8205), .A2(n8204), .ZN(n8208) );
  INV_X1 U9744 ( .A(n6874), .ZN(n8206) );
  AOI21_X1 U9745 ( .B1(n8208), .B2(n8207), .A(n8206), .ZN(n8212) );
  AOI22_X1 U9746 ( .A1(n9068), .A2(n5011), .B1(n8209), .B2(n9037), .ZN(n8211)
         );
  AOI22_X1 U9747 ( .A1(n9067), .A2(n9088), .B1(n8213), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n8210) );
  OAI211_X1 U9748 ( .C1(n8212), .C2(n9075), .A(n8211), .B(n8210), .ZN(P1_U3235) );
  INV_X1 U9749 ( .A(n8213), .ZN(n8219) );
  AOI22_X1 U9750 ( .A1(n9067), .A2(n5011), .B1(n8214), .B2(n9037), .ZN(n8217)
         );
  NAND2_X1 U9751 ( .A1(n8215), .A2(n5747), .ZN(n8216) );
  OAI211_X1 U9752 ( .C1(n8219), .C2(n8218), .A(n8217), .B(n8216), .ZN(P1_U3230) );
  XNOR2_X1 U9753 ( .A(n8230), .B(n8220), .ZN(n8673) );
  XNOR2_X1 U9754 ( .A(n8229), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n8664) );
  NAND2_X1 U9755 ( .A1(n8221), .A2(n10210), .ZN(n8223) );
  NAND2_X1 U9756 ( .A1(n8223), .A2(n8222), .ZN(n8663) );
  NOR2_X1 U9757 ( .A1(n8664), .A2(n8663), .ZN(n8662) );
  AOI21_X1 U9758 ( .B1(n8229), .B2(P2_REG1_REG_17__SCAN_IN), .A(n8662), .ZN(
        n8672) );
  NAND2_X1 U9759 ( .A1(n8673), .A2(n8672), .ZN(n8671) );
  OR2_X1 U9760 ( .A1(n8230), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8224) );
  NAND2_X1 U9761 ( .A1(n8671), .A2(n8224), .ZN(n8225) );
  XNOR2_X1 U9762 ( .A(n8225), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8236) );
  INV_X1 U9763 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n10032) );
  NAND2_X1 U9764 ( .A1(P2_REG2_REG_17__SCAN_IN), .A2(n8229), .ZN(n8228) );
  OAI21_X1 U9765 ( .B1(P2_REG2_REG_17__SCAN_IN), .B2(n8229), .A(n8228), .ZN(
        n8659) );
  INV_X1 U9766 ( .A(n8230), .ZN(n8680) );
  NOR2_X1 U9767 ( .A1(n8231), .A2(n8680), .ZN(n8233) );
  XNOR2_X1 U9768 ( .A(n8234), .B(n6057), .ZN(n8238) );
  NAND2_X1 U9769 ( .A1(n8238), .A2(n9808), .ZN(n8235) );
  INV_X1 U9770 ( .A(n8236), .ZN(n8237) );
  INV_X1 U9771 ( .A(n6484), .ZN(n8241) );
  OAI222_X1 U9772 ( .A1(n8242), .A2(n7025), .B1(n8973), .B2(n8241), .C1(n8240), 
        .C2(P2_U3152), .ZN(P2_U3330) );
  NOR2_X1 U9773 ( .A1(n8579), .A2(n8271), .ZN(n8245) );
  XNOR2_X1 U9774 ( .A(n8913), .B(n8276), .ZN(n8246) );
  XOR2_X1 U9775 ( .A(n8245), .B(n8246), .Z(n8600) );
  XNOR2_X1 U9776 ( .A(n8908), .B(n8247), .ZN(n8249) );
  NAND2_X1 U9777 ( .A1(n8637), .A2(n8274), .ZN(n8248) );
  XNOR2_X1 U9778 ( .A(n8249), .B(n8248), .ZN(n8576) );
  XNOR2_X1 U9779 ( .A(n8250), .B(n4928), .ZN(n8610) );
  NAND2_X1 U9780 ( .A1(n6444), .A2(n8274), .ZN(n8609) );
  NAND2_X1 U9781 ( .A1(n8610), .A2(n8609), .ZN(n8608) );
  INV_X1 U9782 ( .A(n8250), .ZN(n8251) );
  NAND2_X1 U9783 ( .A1(n8608), .A2(n8252), .ZN(n8253) );
  XOR2_X1 U9784 ( .A(n8276), .B(n8896), .Z(n8254) );
  NAND2_X1 U9785 ( .A1(n8253), .A2(n8254), .ZN(n8567) );
  NOR2_X1 U9786 ( .A1(n8613), .A2(n8271), .ZN(n8570) );
  NAND2_X1 U9787 ( .A1(n8567), .A2(n8570), .ZN(n8257) );
  INV_X1 U9788 ( .A(n8253), .ZN(n8256) );
  INV_X1 U9789 ( .A(n8254), .ZN(n8255) );
  XNOR2_X1 U9790 ( .A(n8891), .B(n8276), .ZN(n8259) );
  INV_X1 U9791 ( .A(n8774), .ZN(n8636) );
  NAND2_X1 U9792 ( .A1(n8636), .A2(n8274), .ZN(n8592) );
  INV_X1 U9793 ( .A(n8258), .ZN(n8261) );
  INV_X1 U9794 ( .A(n8259), .ZN(n8260) );
  NOR2_X1 U9795 ( .A1(n8263), .A2(n8271), .ZN(n8264) );
  XNOR2_X1 U9796 ( .A(n8887), .B(n8276), .ZN(n8265) );
  XOR2_X1 U9797 ( .A(n8264), .B(n8265), .Z(n8585) );
  NAND2_X1 U9798 ( .A1(n8584), .A2(n8585), .ZN(n8267) );
  NAND2_X1 U9799 ( .A1(n8265), .A2(n8264), .ZN(n8266) );
  NAND2_X1 U9800 ( .A1(n8267), .A2(n8266), .ZN(n8621) );
  NOR2_X1 U9801 ( .A1(n8714), .A2(n8271), .ZN(n8268) );
  XNOR2_X1 U9802 ( .A(n8883), .B(n8276), .ZN(n8269) );
  XOR2_X1 U9803 ( .A(n8268), .B(n8269), .Z(n8622) );
  NAND2_X1 U9804 ( .A1(n8269), .A2(n8268), .ZN(n8270) );
  NOR2_X1 U9805 ( .A1(n8702), .A2(n8271), .ZN(n8272) );
  XNOR2_X1 U9806 ( .A(n8876), .B(n8276), .ZN(n8273) );
  XOR2_X1 U9807 ( .A(n8272), .B(n8273), .Z(n8560) );
  NAND2_X1 U9808 ( .A1(n8634), .A2(n8274), .ZN(n8275) );
  XOR2_X1 U9809 ( .A(n8276), .B(n8275), .Z(n8277) );
  XNOR2_X1 U9810 ( .A(n8871), .B(n8277), .ZN(n8278) );
  NOR2_X1 U9811 ( .A1(n8702), .A2(n8602), .ZN(n8282) );
  INV_X1 U9812 ( .A(n8279), .ZN(n8696) );
  AOI22_X1 U9813 ( .A1(n8696), .A2(n8625), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3152), .ZN(n8280) );
  OAI21_X1 U9814 ( .B1(n8701), .B2(n8603), .A(n8280), .ZN(n8281) );
  AOI211_X1 U9815 ( .C1(n8871), .C2(n8629), .A(n8282), .B(n8281), .ZN(n8283)
         );
  OAI21_X1 U9816 ( .B1(n8284), .B2(n8631), .A(n8283), .ZN(P2_U3222) );
  NAND2_X1 U9817 ( .A1(n8554), .A2(n8389), .ZN(n8286) );
  INV_X1 U9818 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8556) );
  OR2_X1 U9819 ( .A1(n8391), .A2(n8556), .ZN(n8285) );
  NAND2_X1 U9820 ( .A1(n8287), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n8292) );
  NAND2_X1 U9821 ( .A1(n8288), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n8291) );
  NAND2_X1 U9822 ( .A1(n8289), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n8290) );
  AND3_X1 U9823 ( .A1(n8292), .A2(n8291), .A3(n8290), .ZN(n9158) );
  NAND2_X1 U9824 ( .A1(n8539), .A2(n8394), .ZN(n8295) );
  NAND2_X1 U9825 ( .A1(n8964), .A2(n8389), .ZN(n8294) );
  OR2_X1 U9826 ( .A1(n8391), .A2(n6730), .ZN(n8293) );
  INV_X1 U9827 ( .A(n8400), .ZN(n8464) );
  INV_X1 U9828 ( .A(n9158), .ZN(n9077) );
  NAND2_X1 U9829 ( .A1(n9077), .A2(n8394), .ZN(n8296) );
  NAND2_X1 U9830 ( .A1(n9111), .A2(n8296), .ZN(n8461) );
  INV_X1 U9831 ( .A(n9259), .ZN(n9128) );
  OR2_X1 U9832 ( .A1(n9402), .A2(n9128), .ZN(n8453) );
  NAND2_X1 U9833 ( .A1(n9402), .A2(n9128), .ZN(n9229) );
  INV_X1 U9834 ( .A(n9280), .ZN(n9244) );
  INV_X1 U9835 ( .A(n9407), .ZN(n9270) );
  MUX2_X1 U9836 ( .A(n9244), .B(n9270), .S(n8406), .Z(n8297) );
  NAND2_X1 U9837 ( .A1(n9239), .A2(n8297), .ZN(n8303) );
  OAI21_X1 U9838 ( .B1(n8303), .B2(n9270), .A(n9149), .ZN(n8299) );
  OAI211_X1 U9839 ( .C1(n8303), .C2(n9244), .A(n9211), .B(n8453), .ZN(n8298)
         );
  MUX2_X1 U9840 ( .A(n8299), .B(n8298), .S(n8406), .Z(n8300) );
  INV_X1 U9841 ( .A(n8300), .ZN(n8370) );
  NAND2_X1 U9842 ( .A1(n9407), .A2(n9280), .ZN(n9127) );
  INV_X1 U9843 ( .A(n9127), .ZN(n8301) );
  NAND2_X1 U9844 ( .A1(n9239), .A2(n8301), .ZN(n8302) );
  NAND2_X1 U9845 ( .A1(n8303), .A2(n8302), .ZN(n8369) );
  NAND2_X1 U9846 ( .A1(n9432), .A2(n8991), .ZN(n9323) );
  INV_X1 U9847 ( .A(n9539), .ZN(n9345) );
  AND2_X1 U9848 ( .A1(n9435), .A2(n9345), .ZN(n9140) );
  INV_X1 U9849 ( .A(n9140), .ZN(n8305) );
  NAND2_X1 U9850 ( .A1(n9323), .A2(n8305), .ZN(n8408) );
  OR2_X1 U9851 ( .A1(n9435), .A2(n9345), .ZN(n9339) );
  NAND2_X1 U9852 ( .A1(n8472), .A2(n9339), .ZN(n9141) );
  MUX2_X1 U9853 ( .A(n8408), .B(n9141), .S(n8406), .Z(n8304) );
  INV_X1 U9854 ( .A(n8304), .ZN(n8352) );
  AND2_X1 U9855 ( .A1(n8305), .A2(n9339), .ZN(n9359) );
  OR2_X1 U9856 ( .A1(n9544), .A2(n8306), .ZN(n8422) );
  NAND2_X1 U9857 ( .A1(n9544), .A2(n8306), .ZN(n9139) );
  MUX2_X1 U9858 ( .A(n8422), .B(n9139), .S(n8406), .Z(n8350) );
  OAI211_X1 U9859 ( .C1(n8308), .C2(n8307), .A(n8425), .B(n8434), .ZN(n8309)
         );
  NAND2_X1 U9860 ( .A1(n8309), .A2(n8435), .ZN(n8314) );
  NAND3_X1 U9861 ( .A1(n8311), .A2(n8310), .A3(n8435), .ZN(n8312) );
  NAND2_X1 U9862 ( .A1(n8312), .A2(n8425), .ZN(n8313) );
  MUX2_X1 U9863 ( .A(n8314), .B(n8313), .S(n8406), .Z(n8328) );
  INV_X1 U9864 ( .A(n8328), .ZN(n8326) );
  INV_X1 U9865 ( .A(n8315), .ZN(n8316) );
  NAND2_X1 U9866 ( .A1(n8316), .A2(n8329), .ZN(n8319) );
  INV_X1 U9867 ( .A(n8317), .ZN(n8318) );
  NOR2_X1 U9868 ( .A1(n8319), .A2(n8318), .ZN(n8416) );
  INV_X1 U9869 ( .A(n8319), .ZN(n8323) );
  NAND2_X1 U9870 ( .A1(n9492), .A2(n8436), .ZN(n8322) );
  INV_X1 U9871 ( .A(n8320), .ZN(n8321) );
  AOI21_X1 U9872 ( .B1(n8323), .B2(n8322), .A(n8321), .ZN(n8324) );
  NAND2_X1 U9873 ( .A1(n8412), .A2(n8324), .ZN(n8325) );
  AOI21_X1 U9874 ( .B1(n8326), .B2(n8416), .A(n8325), .ZN(n8332) );
  INV_X1 U9875 ( .A(n8329), .ZN(n8331) );
  OR2_X1 U9876 ( .A1(n8331), .A2(n8330), .ZN(n8410) );
  INV_X1 U9877 ( .A(n8406), .ZN(n8385) );
  AND2_X1 U9878 ( .A1(n8333), .A2(n8340), .ZN(n8415) );
  AND2_X1 U9879 ( .A1(n8419), .A2(n8406), .ZN(n8339) );
  AND2_X1 U9880 ( .A1(n8341), .A2(n8334), .ZN(n8409) );
  NAND2_X1 U9881 ( .A1(n8412), .A2(n8411), .ZN(n8336) );
  AOI21_X1 U9882 ( .B1(n8336), .B2(n8335), .A(n8406), .ZN(n8337) );
  AOI22_X1 U9883 ( .A1(n8415), .A2(n8339), .B1(n8409), .B2(n8337), .ZN(n8338)
         );
  INV_X1 U9884 ( .A(n8339), .ZN(n8345) );
  INV_X1 U9885 ( .A(n8489), .ZN(n8344) );
  NAND2_X1 U9886 ( .A1(n8419), .A2(n8340), .ZN(n8342) );
  NAND3_X1 U9887 ( .A1(n8342), .A2(n8385), .A3(n8341), .ZN(n8343) );
  OAI211_X1 U9888 ( .C1(n8409), .C2(n8345), .A(n8344), .B(n8343), .ZN(n8347)
         );
  MUX2_X1 U9889 ( .A(n8421), .B(n9534), .S(n8385), .Z(n8346) );
  OAI211_X1 U9890 ( .C1(n8348), .C2(n8347), .A(n9546), .B(n8346), .ZN(n8349)
         );
  NAND3_X1 U9891 ( .A1(n9359), .A2(n8350), .A3(n8349), .ZN(n8351) );
  NAND2_X1 U9892 ( .A1(n8352), .A2(n8351), .ZN(n8355) );
  INV_X1 U9893 ( .A(n9309), .ZN(n9347) );
  OR2_X1 U9894 ( .A1(n9425), .A2(n9347), .ZN(n8471) );
  NAND3_X1 U9895 ( .A1(n8355), .A2(n8471), .A3(n8472), .ZN(n8354) );
  INV_X1 U9896 ( .A(n9327), .ZN(n9290) );
  INV_X1 U9897 ( .A(n9144), .ZN(n8353) );
  NAND2_X1 U9898 ( .A1(n9425), .A2(n9347), .ZN(n9142) );
  NAND3_X1 U9899 ( .A1(n8354), .A2(n8353), .A3(n9142), .ZN(n8358) );
  AND2_X1 U9900 ( .A1(n9143), .A2(n8471), .ZN(n8448) );
  AND2_X1 U9901 ( .A1(n9142), .A2(n9323), .ZN(n8447) );
  NAND2_X1 U9902 ( .A1(n8355), .A2(n8447), .ZN(n8356) );
  NAND2_X1 U9903 ( .A1(n8448), .A2(n8356), .ZN(n8357) );
  MUX2_X1 U9904 ( .A(n8358), .B(n8357), .S(n8406), .Z(n8365) );
  INV_X1 U9905 ( .A(n9310), .ZN(n9124) );
  AND2_X1 U9906 ( .A1(n8469), .A2(n9143), .ZN(n8360) );
  NAND2_X1 U9907 ( .A1(n9417), .A2(n9124), .ZN(n9145) );
  INV_X1 U9908 ( .A(n9145), .ZN(n8359) );
  AOI21_X1 U9909 ( .B1(n8365), .B2(n8360), .A(n8359), .ZN(n8361) );
  INV_X1 U9910 ( .A(n9258), .ZN(n9291) );
  INV_X1 U9911 ( .A(n9146), .ZN(n8450) );
  NAND2_X1 U9912 ( .A1(n9410), .A2(n9291), .ZN(n9256) );
  OAI21_X1 U9913 ( .B1(n8361), .B2(n8450), .A(n9256), .ZN(n8368) );
  INV_X1 U9914 ( .A(n8469), .ZN(n8364) );
  NAND2_X1 U9915 ( .A1(n8469), .A2(n9144), .ZN(n8362) );
  AND2_X1 U9916 ( .A1(n8362), .A2(n9145), .ZN(n8363) );
  AND2_X1 U9917 ( .A1(n8363), .A2(n9256), .ZN(n8452) );
  OAI21_X1 U9918 ( .B1(n8365), .B2(n8364), .A(n8452), .ZN(n8366) );
  NAND2_X1 U9919 ( .A1(n8366), .A2(n9146), .ZN(n8367) );
  NAND2_X1 U9920 ( .A1(n8371), .A2(n9131), .ZN(n8375) );
  OAI21_X1 U9921 ( .B1(n9391), .B2(n9211), .A(n9131), .ZN(n8372) );
  MUX2_X1 U9922 ( .A(n9391), .B(n8372), .S(n8385), .Z(n8373) );
  INV_X1 U9923 ( .A(n8373), .ZN(n8374) );
  NAND2_X1 U9924 ( .A1(n8375), .A2(n8374), .ZN(n8384) );
  NAND2_X1 U9925 ( .A1(n9385), .A2(n9176), .ZN(n8443) );
  INV_X1 U9926 ( .A(n9211), .ZN(n8376) );
  INV_X1 U9927 ( .A(n9391), .ZN(n9210) );
  OAI21_X1 U9928 ( .B1(n8376), .B2(n9210), .A(n8443), .ZN(n8379) );
  NAND2_X1 U9929 ( .A1(n8466), .A2(n9232), .ZN(n8377) );
  NAND2_X1 U9930 ( .A1(n9151), .A2(n8377), .ZN(n8378) );
  MUX2_X1 U9931 ( .A(n8379), .B(n8378), .S(n8406), .Z(n8380) );
  OAI21_X1 U9932 ( .B1(n8381), .B2(n9196), .A(n8380), .ZN(n8383) );
  NAND2_X1 U9933 ( .A1(n9179), .A2(n9157), .ZN(n8444) );
  MUX2_X1 U9934 ( .A(n9151), .B(n8443), .S(n8406), .Z(n8382) );
  MUX2_X1 U9935 ( .A(n8458), .B(n8444), .S(n8385), .Z(n8386) );
  AND3_X1 U9936 ( .A1(n8461), .A2(n8387), .A3(n8386), .ZN(n8388) );
  NAND2_X1 U9937 ( .A1(n8464), .A2(n8388), .ZN(n8398) );
  NAND2_X1 U9938 ( .A1(n8390), .A2(n8389), .ZN(n8393) );
  OR2_X1 U9939 ( .A1(n8391), .A2(n10023), .ZN(n8392) );
  INV_X1 U9940 ( .A(n8394), .ZN(n9106) );
  OAI22_X1 U9941 ( .A1(n8398), .A2(n9161), .B1(n8540), .B2(n8461), .ZN(n8405)
         );
  INV_X1 U9942 ( .A(n9078), .ZN(n9177) );
  INV_X1 U9943 ( .A(n8444), .ZN(n8395) );
  OAI21_X1 U9944 ( .B1(n8399), .B2(n8395), .A(n9177), .ZN(n8396) );
  NAND3_X1 U9945 ( .A1(n8396), .A2(n9161), .A3(n8461), .ZN(n8397) );
  OAI211_X1 U9946 ( .C1(n8398), .C2(n9177), .A(n8397), .B(n8464), .ZN(n8403)
         );
  NAND2_X1 U9947 ( .A1(n9376), .A2(n9177), .ZN(n8535) );
  INV_X1 U9948 ( .A(n8458), .ZN(n9152) );
  AOI21_X1 U9949 ( .B1(n8535), .B2(n8401), .A(n8400), .ZN(n8402) );
  NOR4_X1 U9950 ( .A1(n8506), .A2(n8500), .A3(n5738), .A4(n5744), .ZN(n8511)
         );
  INV_X1 U9951 ( .A(n9139), .ZN(n8407) );
  OR2_X1 U9952 ( .A1(n8408), .A2(n8407), .ZN(n8439) );
  INV_X1 U9953 ( .A(n8409), .ZN(n8414) );
  NAND3_X1 U9954 ( .A1(n8412), .A2(n8411), .A3(n8410), .ZN(n8413) );
  NOR2_X1 U9955 ( .A1(n8414), .A2(n8413), .ZN(n8437) );
  INV_X1 U9956 ( .A(n8437), .ZN(n8417) );
  OAI22_X1 U9957 ( .A1(n8417), .A2(n8416), .B1(n8415), .B2(n8414), .ZN(n8418)
         );
  NAND2_X1 U9958 ( .A1(n8418), .A2(n9534), .ZN(n8423) );
  NAND2_X1 U9959 ( .A1(n9534), .A2(n4866), .ZN(n8420) );
  AND4_X1 U9960 ( .A1(n8423), .A2(n8422), .A3(n8421), .A4(n8420), .ZN(n8424)
         );
  OR2_X1 U9961 ( .A1(n8439), .A2(n8424), .ZN(n8529) );
  INV_X1 U9962 ( .A(n8425), .ZN(n8526) );
  OAI211_X1 U9963 ( .C1(n8429), .C2(n8428), .A(n8427), .B(n8426), .ZN(n8475)
         );
  INV_X1 U9964 ( .A(n8476), .ZN(n8430) );
  NAND2_X1 U9965 ( .A1(n8475), .A2(n8430), .ZN(n8433) );
  AND2_X1 U9966 ( .A1(n8432), .A2(n8431), .ZN(n8524) );
  AOI22_X1 U9967 ( .A1(n8434), .A2(n8433), .B1(n7163), .B2(n8524), .ZN(n8440)
         );
  NAND4_X1 U9968 ( .A1(n8437), .A2(n9534), .A3(n8436), .A4(n8435), .ZN(n8438)
         );
  NOR2_X1 U9969 ( .A1(n8439), .A2(n8438), .ZN(n8513) );
  OAI21_X1 U9970 ( .B1(n8526), .B2(n8440), .A(n8513), .ZN(n8446) );
  INV_X1 U9971 ( .A(n9150), .ZN(n8441) );
  NAND2_X1 U9972 ( .A1(n9151), .A2(n8441), .ZN(n8442) );
  NAND3_X1 U9973 ( .A1(n8444), .A2(n8443), .A3(n8442), .ZN(n8460) );
  NAND2_X1 U9974 ( .A1(n9407), .A2(n9244), .ZN(n8468) );
  NAND4_X1 U9975 ( .A1(n9149), .A2(n8452), .A3(n8468), .A4(n9142), .ZN(n8445)
         );
  OR2_X1 U9976 ( .A1(n8460), .A2(n8445), .ZN(n8534) );
  AOI21_X1 U9977 ( .B1(n8529), .B2(n8446), .A(n8534), .ZN(n8462) );
  INV_X1 U9978 ( .A(n8447), .ZN(n8449) );
  OAI211_X1 U9979 ( .C1(n4843), .C2(n8449), .A(n8469), .B(n8448), .ZN(n8451)
         );
  AOI21_X1 U9980 ( .B1(n8452), .B2(n8451), .A(n8450), .ZN(n8455) );
  INV_X1 U9981 ( .A(n8468), .ZN(n8454) );
  OAI211_X1 U9982 ( .C1(n8455), .C2(n8454), .A(n8453), .B(n9240), .ZN(n8456)
         );
  NAND2_X1 U9983 ( .A1(n9149), .A2(n8456), .ZN(n8457) );
  AND4_X1 U9984 ( .A1(n9151), .A2(n9211), .A3(n8467), .A4(n8457), .ZN(n8459)
         );
  OAI211_X1 U9985 ( .C1(n8460), .C2(n8459), .A(n8465), .B(n8458), .ZN(n8536)
         );
  OAI211_X1 U9986 ( .C1(n8462), .C2(n8536), .A(n8461), .B(n8535), .ZN(n8463)
         );
  AOI211_X1 U9987 ( .C1(n8464), .C2(n8463), .A(n5744), .B(n8500), .ZN(n8505)
         );
  INV_X1 U9988 ( .A(n9173), .ZN(n8497) );
  INV_X1 U9989 ( .A(n9255), .ZN(n8494) );
  NAND2_X1 U9990 ( .A1(n9146), .A2(n9256), .ZN(n9279) );
  INV_X1 U9991 ( .A(n9143), .ZN(n8470) );
  NOR2_X1 U9992 ( .A1(n8470), .A2(n9144), .ZN(n9307) );
  NAND2_X1 U9993 ( .A1(n8472), .A2(n9323), .ZN(n9342) );
  INV_X1 U9994 ( .A(n9342), .ZN(n8492) );
  INV_X1 U9995 ( .A(n9359), .ZN(n8490) );
  INV_X1 U9996 ( .A(n9546), .ZN(n9535) );
  NAND4_X1 U9997 ( .A1(n8475), .A2(n8474), .A3(n4367), .A4(n8473), .ZN(n8477)
         );
  NOR2_X1 U9998 ( .A1(n8477), .A2(n8476), .ZN(n8480) );
  NAND4_X1 U9999 ( .A1(n8480), .A2(n8479), .A3(n8478), .A4(n8524), .ZN(n8481)
         );
  NOR4_X1 U10000 ( .A1(n8483), .A2(n8482), .A3(n9494), .A4(n8481), .ZN(n8485)
         );
  NAND4_X1 U10001 ( .A1(n8487), .A2(n8486), .A3(n8485), .A4(n8484), .ZN(n8488)
         );
  NOR4_X1 U10002 ( .A1(n8490), .A2(n9535), .A3(n8489), .A4(n8488), .ZN(n8491)
         );
  NAND4_X1 U10003 ( .A1(n9307), .A2(n9322), .A3(n8492), .A4(n8491), .ZN(n8493)
         );
  NOR4_X1 U10004 ( .A1(n8494), .A2(n9279), .A3(n9288), .A4(n8493), .ZN(n8495)
         );
  NAND3_X1 U10005 ( .A1(n9214), .A2(n9239), .A3(n8495), .ZN(n8496) );
  NOR4_X1 U10006 ( .A1(n8497), .A2(n9196), .A3(n9231), .A4(n8496), .ZN(n8499)
         );
  INV_X1 U10007 ( .A(n8540), .ZN(n8498) );
  NAND4_X1 U10008 ( .A1(n8539), .A2(n9153), .A3(n8499), .A4(n8498), .ZN(n8503)
         );
  INV_X1 U10009 ( .A(n8500), .ZN(n8502) );
  NAND2_X1 U10010 ( .A1(n9111), .A2(n9158), .ZN(n8501) );
  NAND2_X1 U10011 ( .A1(n8502), .A2(n8501), .ZN(n8512) );
  OAI21_X1 U10012 ( .B1(n8503), .B2(n8512), .A(n5744), .ZN(n8507) );
  INV_X1 U10013 ( .A(n8507), .ZN(n8504) );
  NOR2_X1 U10014 ( .A1(n8505), .A2(n8504), .ZN(n8509) );
  NOR3_X1 U10015 ( .A1(n8511), .A2(n8510), .A3(n8543), .ZN(n8553) );
  INV_X1 U10016 ( .A(n8512), .ZN(n8542) );
  INV_X1 U10017 ( .A(n8513), .ZN(n8531) );
  NAND2_X1 U10018 ( .A1(n6638), .A2(n9705), .ZN(n8516) );
  NAND2_X1 U10019 ( .A1(n5011), .A2(n9757), .ZN(n8515) );
  NAND3_X1 U10020 ( .A1(n8516), .A2(n8515), .A3(n8514), .ZN(n8517) );
  NAND2_X1 U10021 ( .A1(n8518), .A2(n8517), .ZN(n8520) );
  OAI21_X1 U10022 ( .B1(n8521), .B2(n8520), .A(n8519), .ZN(n8523) );
  NAND2_X1 U10023 ( .A1(n8523), .A2(n8522), .ZN(n8525) );
  NAND2_X1 U10024 ( .A1(n8525), .A2(n8524), .ZN(n8528) );
  AOI21_X1 U10025 ( .B1(n8528), .B2(n8527), .A(n8526), .ZN(n8530) );
  OAI21_X1 U10026 ( .B1(n8531), .B2(n8530), .A(n8529), .ZN(n8532) );
  INV_X1 U10027 ( .A(n8532), .ZN(n8533) );
  NOR2_X1 U10028 ( .A1(n8534), .A2(n8533), .ZN(n8537) );
  OAI21_X1 U10029 ( .B1(n8537), .B2(n8536), .A(n8535), .ZN(n8538) );
  NAND2_X1 U10030 ( .A1(n8539), .A2(n8538), .ZN(n8541) );
  AOI21_X1 U10031 ( .B1(n8542), .B2(n8541), .A(n8540), .ZN(n8547) );
  NAND3_X1 U10032 ( .A1(n8547), .A2(n5505), .A3(n8543), .ZN(n8545) );
  OAI211_X1 U10033 ( .C1(n8547), .C2(n8546), .A(n8545), .B(n8544), .ZN(n8552)
         );
  NOR3_X1 U10034 ( .A1(n8548), .A2(n5759), .A3(n9104), .ZN(n8551) );
  OAI21_X1 U10035 ( .B1(n5738), .B2(n8549), .A(P1_B_REG_SCAN_IN), .ZN(n8550)
         );
  OAI22_X1 U10036 ( .A1(n8553), .A2(n8552), .B1(n8551), .B2(n8550), .ZN(
        P1_U3240) );
  INV_X1 U10037 ( .A(n8554), .ZN(n8974) );
  OAI222_X1 U10038 ( .A1(n8557), .A2(n8556), .B1(n4370), .B2(n8974), .C1(
        P1_U3084), .C2(n4947), .ZN(P1_U3323) );
  OAI222_X1 U10039 ( .A1(n4370), .A2(n8559), .B1(n5744), .B2(P1_U3084), .C1(
        n8558), .C2(n8557), .ZN(P1_U3332) );
  XNOR2_X1 U10040 ( .A(n8561), .B(n8560), .ZN(n8566) );
  OAI22_X1 U10041 ( .A1(n8714), .A2(n8602), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10178), .ZN(n8562) );
  AOI21_X1 U10042 ( .B1(n8711), .B2(n8625), .A(n8562), .ZN(n8563) );
  OAI21_X1 U10043 ( .B1(n8715), .B2(n8603), .A(n8563), .ZN(n8564) );
  AOI21_X1 U10044 ( .B1(n8876), .B2(n8629), .A(n8564), .ZN(n8565) );
  OAI21_X1 U10045 ( .B1(n8566), .B2(n8631), .A(n8565), .ZN(P2_U3216) );
  NAND2_X1 U10046 ( .A1(n8568), .A2(n8567), .ZN(n8569) );
  XOR2_X1 U10047 ( .A(n8570), .B(n8569), .Z(n8575) );
  NAND2_X1 U10048 ( .A1(n8636), .A2(n8596), .ZN(n8572) );
  AOI22_X1 U10049 ( .A1(n8778), .A2(n8625), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3152), .ZN(n8571) );
  OAI211_X1 U10050 ( .C1(n8775), .C2(n8602), .A(n8572), .B(n8571), .ZN(n8573)
         );
  AOI21_X1 U10051 ( .B1(n8896), .B2(n8629), .A(n8573), .ZN(n8574) );
  OAI21_X1 U10052 ( .B1(n8575), .B2(n8631), .A(n8574), .ZN(P2_U3218) );
  XNOR2_X1 U10053 ( .A(n8577), .B(n8576), .ZN(n8583) );
  INV_X1 U10054 ( .A(n8808), .ZN(n8578) );
  OAI22_X1 U10055 ( .A1(n8615), .A2(n8578), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10062), .ZN(n8581) );
  OAI22_X1 U10056 ( .A1(n8775), .A2(n8603), .B1(n8579), .B2(n8602), .ZN(n8580)
         );
  AOI211_X1 U10057 ( .C1(n8908), .C2(n8629), .A(n8581), .B(n8580), .ZN(n8582)
         );
  OAI21_X1 U10058 ( .B1(n8583), .B2(n8631), .A(n8582), .ZN(P2_U3225) );
  XNOR2_X1 U10059 ( .A(n8584), .B(n8585), .ZN(n8590) );
  OAI22_X1 U10060 ( .A1(n8714), .A2(n8830), .B1(n8774), .B2(n8828), .ZN(n8748)
         );
  OAI22_X1 U10061 ( .A1(n8742), .A2(n8615), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8586), .ZN(n8587) );
  AOI21_X1 U10062 ( .B1(n8748), .B2(n8617), .A(n8587), .ZN(n8589) );
  NAND2_X1 U10063 ( .A1(n8887), .A2(n8629), .ZN(n8588) );
  OAI211_X1 U10064 ( .C1(n8590), .C2(n8631), .A(n8589), .B(n8588), .ZN(
        P2_U3227) );
  XNOR2_X1 U10065 ( .A(n8591), .B(n8592), .ZN(n8599) );
  OAI22_X1 U10066 ( .A1(n8760), .A2(n8615), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8593), .ZN(n8595) );
  NOR2_X1 U10067 ( .A1(n8613), .A2(n8602), .ZN(n8594) );
  AOI211_X1 U10068 ( .C1(n8767), .C2(n8596), .A(n8595), .B(n8594), .ZN(n8598)
         );
  NAND2_X1 U10069 ( .A1(n8891), .A2(n8629), .ZN(n8597) );
  OAI211_X1 U10070 ( .C1(n8599), .C2(n8631), .A(n8598), .B(n8597), .ZN(
        P2_U3231) );
  XNOR2_X1 U10071 ( .A(n8601), .B(n8600), .ZN(n8607) );
  OAI22_X1 U10072 ( .A1(n8615), .A2(n8821), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10090), .ZN(n8605) );
  OAI22_X1 U10073 ( .A1(n8831), .A2(n8603), .B1(n8602), .B2(n8829), .ZN(n8604)
         );
  AOI211_X1 U10074 ( .C1(n8913), .C2(n8629), .A(n8605), .B(n8604), .ZN(n8606)
         );
  OAI21_X1 U10075 ( .B1(n8607), .B2(n8631), .A(n8606), .ZN(P2_U3235) );
  OAI21_X1 U10076 ( .B1(n8610), .B2(n8609), .A(n8608), .ZN(n8612) );
  NAND2_X1 U10077 ( .A1(n8612), .A2(n8611), .ZN(n8619) );
  OAI22_X1 U10078 ( .A1(n8613), .A2(n8830), .B1(n8831), .B2(n8828), .ZN(n8797)
         );
  OAI22_X1 U10079 ( .A1(n8615), .A2(n8791), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8614), .ZN(n8616) );
  AOI21_X1 U10080 ( .B1(n8797), .B2(n8617), .A(n8616), .ZN(n8618) );
  OAI211_X1 U10081 ( .C1(n4552), .C2(n8620), .A(n8619), .B(n8618), .ZN(
        P2_U3237) );
  XNOR2_X1 U10082 ( .A(n8621), .B(n8622), .ZN(n8632) );
  OR2_X1 U10083 ( .A1(n8702), .A2(n8830), .ZN(n8624) );
  NAND2_X1 U10084 ( .A1(n8767), .A2(n8838), .ZN(n8623) );
  AND2_X1 U10085 ( .A1(n8624), .A2(n8623), .ZN(n8727) );
  AOI22_X1 U10086 ( .A1(n8732), .A2(n8625), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3152), .ZN(n8626) );
  OAI21_X1 U10087 ( .B1(n8727), .B2(n8627), .A(n8626), .ZN(n8628) );
  AOI21_X1 U10088 ( .B1(n8883), .B2(n8629), .A(n8628), .ZN(n8630) );
  OAI21_X1 U10089 ( .B1(n8632), .B2(n8631), .A(n8630), .ZN(P2_U3242) );
  MUX2_X1 U10090 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8633), .S(P2_U3966), .Z(
        P2_U3582) );
  MUX2_X1 U10091 ( .A(n8634), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8638), .Z(
        P2_U3580) );
  MUX2_X1 U10092 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8635), .S(P2_U3966), .Z(
        P2_U3579) );
  MUX2_X1 U10093 ( .A(n8767), .B(P2_DATAO_REG_25__SCAN_IN), .S(n8638), .Z(
        P2_U3577) );
  MUX2_X1 U10094 ( .A(n8636), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8638), .Z(
        P2_U3576) );
  MUX2_X1 U10095 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n6444), .S(P2_U3966), .Z(
        P2_U3574) );
  MUX2_X1 U10096 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8637), .S(P2_U3966), .Z(
        P2_U3573) );
  MUX2_X1 U10097 ( .A(n8804), .B(P2_DATAO_REG_20__SCAN_IN), .S(n8638), .Z(
        P2_U3572) );
  MUX2_X1 U10098 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8841), .S(P2_U3966), .Z(
        P2_U3571) );
  MUX2_X1 U10099 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8639), .S(P2_U3966), .Z(
        P2_U3570) );
  MUX2_X1 U10100 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8839), .S(P2_U3966), .Z(
        P2_U3569) );
  MUX2_X1 U10101 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8640), .S(P2_U3966), .Z(
        P2_U3568) );
  MUX2_X1 U10102 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8641), .S(P2_U3966), .Z(
        P2_U3567) );
  MUX2_X1 U10103 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8642), .S(P2_U3966), .Z(
        P2_U3566) );
  INV_X1 U10104 ( .A(n8643), .ZN(n8644) );
  MUX2_X1 U10105 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n8644), .S(P2_U3966), .Z(
        P2_U3565) );
  MUX2_X1 U10106 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n8645), .S(P2_U3966), .Z(
        P2_U3564) );
  MUX2_X1 U10107 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n8646), .S(P2_U3966), .Z(
        P2_U3563) );
  MUX2_X1 U10108 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n8647), .S(P2_U3966), .Z(
        P2_U3562) );
  MUX2_X1 U10109 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n8648), .S(P2_U3966), .Z(
        P2_U3561) );
  MUX2_X1 U10110 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n8649), .S(P2_U3966), .Z(
        P2_U3560) );
  MUX2_X1 U10111 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n8650), .S(P2_U3966), .Z(
        P2_U3559) );
  MUX2_X1 U10112 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n8651), .S(P2_U3966), .Z(
        P2_U3558) );
  MUX2_X1 U10113 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n8652), .S(P2_U3966), .Z(
        P2_U3557) );
  MUX2_X1 U10114 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n8653), .S(P2_U3966), .Z(
        P2_U3556) );
  MUX2_X1 U10115 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n8654), .S(P2_U3966), .Z(
        P2_U3555) );
  MUX2_X1 U10116 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n8655), .S(P2_U3966), .Z(
        P2_U3554) );
  MUX2_X1 U10117 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n8656), .S(P2_U3966), .Z(
        P2_U3553) );
  AOI211_X1 U10118 ( .C1(n8660), .C2(n8659), .A(n8658), .B(n8657), .ZN(n8670)
         );
  AND2_X1 U10119 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(P2_U3152), .ZN(n8661) );
  AOI21_X1 U10120 ( .B1(n9813), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n8661), .ZN(
        n8667) );
  AOI21_X1 U10121 ( .B1(n8664), .B2(n8663), .A(n8662), .ZN(n8665) );
  NAND2_X1 U10122 ( .A1(n9807), .A2(n8665), .ZN(n8666) );
  OAI211_X1 U10123 ( .C1(n9809), .C2(n8668), .A(n8667), .B(n8666), .ZN(n8669)
         );
  OR2_X1 U10124 ( .A1(n8670), .A2(n8669), .ZN(P2_U3262) );
  OAI21_X1 U10125 ( .B1(n8673), .B2(n8672), .A(n8671), .ZN(n8677) );
  OAI21_X1 U10126 ( .B1(n8675), .B2(n10060), .A(n8674), .ZN(n8676) );
  AOI21_X1 U10127 ( .B1(n9807), .B2(n8677), .A(n8676), .ZN(n8679) );
  OAI211_X1 U10128 ( .C1(n4405), .C2(P2_REG2_REG_18__SCAN_IN), .A(n9808), .B(
        n4381), .ZN(n8678) );
  OAI211_X1 U10129 ( .C1(n9809), .C2(n8680), .A(n8679), .B(n8678), .ZN(
        P2_U3263) );
  NAND2_X1 U10130 ( .A1(n6196), .A2(n8686), .ZN(n8864) );
  XNOR2_X1 U10131 ( .A(n8864), .B(n8860), .ZN(n8862) );
  NAND2_X1 U10132 ( .A1(n8682), .A2(n8681), .ZN(n8865) );
  NOR2_X1 U10133 ( .A1(n9836), .A2(n8865), .ZN(n8689) );
  AOI21_X1 U10134 ( .B1(n9836), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8689), .ZN(
        n8684) );
  NAND2_X1 U10135 ( .A1(n8860), .A2(n8755), .ZN(n8683) );
  OAI211_X1 U10136 ( .C1(n8862), .C2(n8685), .A(n8684), .B(n8683), .ZN(
        P2_U3265) );
  INV_X1 U10137 ( .A(n8686), .ZN(n8687) );
  NAND2_X1 U10138 ( .A1(n8688), .A2(n8687), .ZN(n8863) );
  NAND3_X1 U10139 ( .A1(n8864), .A2(n8858), .A3(n8863), .ZN(n8691) );
  AOI21_X1 U10140 ( .B1(n9836), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8689), .ZN(
        n8690) );
  OAI211_X1 U10141 ( .C1(n6196), .C2(n8851), .A(n8691), .B(n8690), .ZN(
        P2_U3266) );
  XNOR2_X1 U10142 ( .A(n8693), .B(n8692), .ZN(n8875) );
  INV_X1 U10143 ( .A(n8694), .ZN(n8695) );
  AOI21_X1 U10144 ( .B1(n8871), .B2(n4551), .A(n8695), .ZN(n8872) );
  AOI22_X1 U10145 ( .A1(n8696), .A2(n8848), .B1(P2_REG2_REG_28__SCAN_IN), .B2(
        n9836), .ZN(n8697) );
  OAI21_X1 U10146 ( .B1(n6158), .B2(n8851), .A(n8697), .ZN(n8707) );
  INV_X1 U10147 ( .A(n8698), .ZN(n8700) );
  AOI21_X1 U10148 ( .B1(n8700), .B2(n8699), .A(n8825), .ZN(n8705) );
  OAI22_X1 U10149 ( .A1(n8702), .A2(n8828), .B1(n8701), .B2(n8830), .ZN(n8703)
         );
  AOI21_X1 U10150 ( .B1(n8705), .B2(n8704), .A(n8703), .ZN(n8874) );
  NOR2_X1 U10151 ( .A1(n8874), .A2(n9836), .ZN(n8706) );
  AOI211_X1 U10152 ( .C1(n8872), .C2(n8858), .A(n8707), .B(n8706), .ZN(n8708)
         );
  OAI21_X1 U10153 ( .B1(n8875), .B2(n8855), .A(n8708), .ZN(P2_U3268) );
  XNOR2_X1 U10154 ( .A(n8709), .B(n8713), .ZN(n8880) );
  AOI21_X1 U10155 ( .B1(n8876), .B2(n8729), .A(n8710), .ZN(n8877) );
  AOI22_X1 U10156 ( .A1(n8711), .A2(n8848), .B1(P2_REG2_REG_27__SCAN_IN), .B2(
        n9836), .ZN(n8712) );
  OAI21_X1 U10157 ( .B1(n4889), .B2(n8851), .A(n8712), .ZN(n8720) );
  AOI21_X1 U10158 ( .B1(n4404), .B2(n8713), .A(n8825), .ZN(n8718) );
  OAI22_X1 U10159 ( .A1(n8715), .A2(n8830), .B1(n8714), .B2(n8828), .ZN(n8716)
         );
  AOI21_X1 U10160 ( .B1(n8718), .B2(n8717), .A(n8716), .ZN(n8879) );
  NOR2_X1 U10161 ( .A1(n8879), .A2(n9836), .ZN(n8719) );
  AOI211_X1 U10162 ( .C1(n8877), .C2(n8858), .A(n8720), .B(n8719), .ZN(n8721)
         );
  OAI21_X1 U10163 ( .B1(n8880), .B2(n8855), .A(n8721), .ZN(P2_U3269) );
  XNOR2_X1 U10164 ( .A(n8722), .B(n4767), .ZN(n8885) );
  AOI22_X1 U10165 ( .A1(n8883), .A2(n8755), .B1(n9836), .B2(
        P2_REG2_REG_26__SCAN_IN), .ZN(n8738) );
  INV_X1 U10166 ( .A(n8745), .ZN(n8724) );
  AOI21_X1 U10167 ( .B1(n8724), .B2(n8723), .A(n4767), .ZN(n8725) );
  OAI21_X1 U10168 ( .B1(n8726), .B2(n8725), .A(n8843), .ZN(n8728) );
  NAND2_X1 U10169 ( .A1(n8728), .A2(n8727), .ZN(n8881) );
  INV_X1 U10170 ( .A(n8750), .ZN(n8731) );
  INV_X1 U10171 ( .A(n8729), .ZN(n8730) );
  AOI211_X1 U10172 ( .C1(n8883), .C2(n8731), .A(n9901), .B(n8730), .ZN(n8882)
         );
  INV_X1 U10173 ( .A(n8882), .ZN(n8735) );
  INV_X1 U10174 ( .A(n8732), .ZN(n8733) );
  OAI22_X1 U10175 ( .A1(n8735), .A2(n8734), .B1(n9825), .B2(n8733), .ZN(n8736)
         );
  OAI21_X1 U10176 ( .B1(n8881), .B2(n8736), .A(n9834), .ZN(n8737) );
  OAI211_X1 U10177 ( .C1(n8885), .C2(n8855), .A(n8738), .B(n8737), .ZN(
        P2_U3270) );
  XNOR2_X1 U10178 ( .A(n8740), .B(n8739), .ZN(n8890) );
  INV_X1 U10179 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n8741) );
  OAI22_X1 U10180 ( .A1(n8742), .A2(n9825), .B1(n8741), .B2(n9834), .ZN(n8754)
         );
  NOR2_X1 U10181 ( .A1(n8744), .A2(n8743), .ZN(n8747) );
  AOI211_X1 U10182 ( .C1(n8747), .C2(n8746), .A(n8825), .B(n8745), .ZN(n8749)
         );
  NOR2_X1 U10183 ( .A1(n8749), .A2(n8748), .ZN(n8889) );
  AOI211_X1 U10184 ( .C1(n8887), .C2(n8751), .A(n9901), .B(n8750), .ZN(n8886)
         );
  NAND2_X1 U10185 ( .A1(n8886), .A2(n9827), .ZN(n8752) );
  AOI21_X1 U10186 ( .B1(n8889), .B2(n8752), .A(n9836), .ZN(n8753) );
  AOI211_X1 U10187 ( .C1(n8755), .C2(n8887), .A(n8754), .B(n8753), .ZN(n8756)
         );
  OAI21_X1 U10188 ( .B1(n8890), .B2(n8855), .A(n8756), .ZN(P2_U3271) );
  AOI21_X1 U10189 ( .B1(n8765), .B2(n8758), .A(n8757), .ZN(n8895) );
  XNOR2_X1 U10190 ( .A(n8891), .B(n8777), .ZN(n8892) );
  INV_X1 U10191 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n8759) );
  OAI22_X1 U10192 ( .A1(n8760), .A2(n9825), .B1(n8759), .B2(n9834), .ZN(n8763)
         );
  NOR2_X1 U10193 ( .A1(n8761), .A2(n8851), .ZN(n8762) );
  AOI211_X1 U10194 ( .C1(n8892), .C2(n8858), .A(n8763), .B(n8762), .ZN(n8770)
         );
  XOR2_X1 U10195 ( .A(n8765), .B(n8764), .Z(n8768) );
  AOI222_X1 U10196 ( .A1(n8843), .A2(n8768), .B1(n8767), .B2(n8840), .C1(n8766), .C2(n8838), .ZN(n8894) );
  OR2_X1 U10197 ( .A1(n8894), .A2(n9836), .ZN(n8769) );
  OAI211_X1 U10198 ( .C1(n8895), .C2(n8855), .A(n8770), .B(n8769), .ZN(
        P2_U3272) );
  AOI21_X1 U10199 ( .B1(n8782), .B2(n8772), .A(n8771), .ZN(n8773) );
  OAI222_X1 U10200 ( .A1(n8828), .A2(n8775), .B1(n8830), .B2(n8774), .C1(n8825), .C2(n8773), .ZN(n8776) );
  INV_X1 U10201 ( .A(n8776), .ZN(n8902) );
  AOI21_X1 U10202 ( .B1(n8896), .B2(n8788), .A(n8777), .ZN(n8897) );
  AOI22_X1 U10203 ( .A1(n8778), .A2(n8848), .B1(P2_REG2_REG_23__SCAN_IN), .B2(
        n9836), .ZN(n8779) );
  OAI21_X1 U10204 ( .B1(n8780), .B2(n8851), .A(n8779), .ZN(n8781) );
  AOI21_X1 U10205 ( .B1(n8897), .B2(n8858), .A(n8781), .ZN(n8785) );
  OR2_X1 U10206 ( .A1(n8783), .A2(n8782), .ZN(n8899) );
  NAND3_X1 U10207 ( .A1(n8899), .A2(n8898), .A3(n8813), .ZN(n8784) );
  OAI211_X1 U10208 ( .C1(n8902), .C2(n9836), .A(n8785), .B(n8784), .ZN(
        P2_U3273) );
  XNOR2_X1 U10209 ( .A(n8787), .B(n8786), .ZN(n8907) );
  INV_X1 U10210 ( .A(n8788), .ZN(n8789) );
  AOI21_X1 U10211 ( .B1(n8903), .B2(n8790), .A(n8789), .ZN(n8904) );
  INV_X1 U10212 ( .A(n8791), .ZN(n8792) );
  AOI22_X1 U10213 ( .A1(n8792), .A2(n8848), .B1(P2_REG2_REG_22__SCAN_IN), .B2(
        n9836), .ZN(n8793) );
  OAI21_X1 U10214 ( .B1(n4552), .B2(n8851), .A(n8793), .ZN(n8801) );
  INV_X1 U10215 ( .A(n8794), .ZN(n8796) );
  AOI21_X1 U10216 ( .B1(n8796), .B2(n8795), .A(n8825), .ZN(n8799) );
  AOI21_X1 U10217 ( .B1(n8799), .B2(n8798), .A(n8797), .ZN(n8906) );
  NOR2_X1 U10218 ( .A1(n8906), .A2(n9836), .ZN(n8800) );
  AOI211_X1 U10219 ( .C1(n8904), .C2(n8858), .A(n8801), .B(n8800), .ZN(n8802)
         );
  OAI21_X1 U10220 ( .B1(n8907), .B2(n8855), .A(n8802), .ZN(P2_U3274) );
  XNOR2_X1 U10221 ( .A(n8803), .B(n8806), .ZN(n8805) );
  AOI222_X1 U10222 ( .A1(n8843), .A2(n8805), .B1(n6444), .B2(n8840), .C1(n8804), .C2(n8838), .ZN(n8911) );
  XNOR2_X1 U10223 ( .A(n8807), .B(n8806), .ZN(n8912) );
  INV_X1 U10224 ( .A(n8912), .ZN(n8814) );
  XNOR2_X1 U10225 ( .A(n8811), .B(n8818), .ZN(n8909) );
  NAND2_X1 U10226 ( .A1(n8909), .A2(n8858), .ZN(n8810) );
  AOI22_X1 U10227 ( .A1(P2_REG2_REG_21__SCAN_IN), .A2(n9836), .B1(n8808), .B2(
        n8848), .ZN(n8809) );
  OAI211_X1 U10228 ( .C1(n8811), .C2(n8851), .A(n8810), .B(n8809), .ZN(n8812)
         );
  AOI21_X1 U10229 ( .B1(n8814), .B2(n8813), .A(n8812), .ZN(n8815) );
  OAI21_X1 U10230 ( .B1(n9836), .B2(n8911), .A(n8815), .ZN(P2_U3275) );
  XNOR2_X1 U10231 ( .A(n8816), .B(n8827), .ZN(n8917) );
  INV_X1 U10232 ( .A(n8817), .ZN(n8820) );
  INV_X1 U10233 ( .A(n8818), .ZN(n8819) );
  AOI21_X1 U10234 ( .B1(n8913), .B2(n8820), .A(n8819), .ZN(n8914) );
  INV_X1 U10235 ( .A(n8821), .ZN(n8822) );
  AOI22_X1 U10236 ( .A1(n9836), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8822), .B2(
        n8848), .ZN(n8823) );
  OAI21_X1 U10237 ( .B1(n8824), .B2(n8851), .A(n8823), .ZN(n8835) );
  AOI211_X1 U10238 ( .C1(n8827), .C2(n8826), .A(n8825), .B(n4434), .ZN(n8833)
         );
  OAI22_X1 U10239 ( .A1(n8831), .A2(n8830), .B1(n8829), .B2(n8828), .ZN(n8832)
         );
  NOR2_X1 U10240 ( .A1(n8833), .A2(n8832), .ZN(n8916) );
  NOR2_X1 U10241 ( .A1(n8916), .A2(n9836), .ZN(n8834) );
  AOI211_X1 U10242 ( .C1(n8914), .C2(n8858), .A(n8835), .B(n8834), .ZN(n8836)
         );
  OAI21_X1 U10243 ( .B1(n8855), .B2(n8917), .A(n8836), .ZN(P2_U3276) );
  XNOR2_X1 U10244 ( .A(n8837), .B(n8853), .ZN(n8842) );
  AOI222_X1 U10245 ( .A1(n8843), .A2(n8842), .B1(n8841), .B2(n8840), .C1(n8839), .C2(n8838), .ZN(n8926) );
  INV_X1 U10246 ( .A(n8844), .ZN(n8845) );
  AOI21_X1 U10247 ( .B1(n8923), .B2(n8846), .A(n8845), .ZN(n8924) );
  INV_X1 U10248 ( .A(n8847), .ZN(n8849) );
  AOI22_X1 U10249 ( .A1(n9836), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8849), .B2(
        n8848), .ZN(n8850) );
  OAI21_X1 U10250 ( .B1(n8852), .B2(n8851), .A(n8850), .ZN(n8857) );
  XNOR2_X1 U10251 ( .A(n8854), .B(n8853), .ZN(n8927) );
  NOR2_X1 U10252 ( .A1(n8927), .A2(n8855), .ZN(n8856) );
  AOI211_X1 U10253 ( .C1(n8924), .C2(n8858), .A(n8857), .B(n8856), .ZN(n8859)
         );
  OAI21_X1 U10254 ( .B1(n9836), .B2(n8926), .A(n8859), .ZN(P2_U3278) );
  NAND2_X1 U10255 ( .A1(n8860), .A2(n9882), .ZN(n8861) );
  OAI211_X1 U10256 ( .C1(n8862), .C2(n9901), .A(n8861), .B(n8865), .ZN(n8947)
         );
  MUX2_X1 U10257 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n8947), .S(n9996), .Z(
        P2_U3551) );
  NAND3_X1 U10258 ( .A1(n8864), .A2(n9883), .A3(n8863), .ZN(n8866) );
  OAI211_X1 U10259 ( .C1(n6196), .C2(n9899), .A(n8866), .B(n8865), .ZN(n8948)
         );
  MUX2_X1 U10260 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n8948), .S(n9996), .Z(
        P2_U3550) );
  MUX2_X1 U10261 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n8949), .S(n9996), .Z(
        P2_U3549) );
  AOI22_X1 U10262 ( .A1(n8872), .A2(n9883), .B1(n9882), .B2(n8871), .ZN(n8873)
         );
  OAI211_X1 U10263 ( .C1(n8875), .C2(n9532), .A(n8874), .B(n8873), .ZN(n8950)
         );
  MUX2_X1 U10264 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n8950), .S(n9996), .Z(
        P2_U3548) );
  AOI22_X1 U10265 ( .A1(n8877), .A2(n9883), .B1(n9882), .B2(n8876), .ZN(n8878)
         );
  OAI211_X1 U10266 ( .C1(n8880), .C2(n9532), .A(n8879), .B(n8878), .ZN(n8951)
         );
  MUX2_X1 U10267 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8951), .S(n9996), .Z(
        P2_U3547) );
  AOI211_X1 U10268 ( .C1(n9882), .C2(n8883), .A(n8882), .B(n8881), .ZN(n8884)
         );
  OAI21_X1 U10269 ( .B1(n8885), .B2(n9532), .A(n8884), .ZN(n8952) );
  MUX2_X1 U10270 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n8952), .S(n9996), .Z(
        P2_U3546) );
  AOI21_X1 U10271 ( .B1(n9882), .B2(n8887), .A(n8886), .ZN(n8888) );
  OAI211_X1 U10272 ( .C1(n8890), .C2(n9532), .A(n8889), .B(n8888), .ZN(n8953)
         );
  MUX2_X1 U10273 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8953), .S(n9996), .Z(
        P2_U3545) );
  AOI22_X1 U10274 ( .A1(n8892), .A2(n9883), .B1(n9882), .B2(n8891), .ZN(n8893)
         );
  OAI211_X1 U10275 ( .C1(n8895), .C2(n9532), .A(n8894), .B(n8893), .ZN(n8954)
         );
  MUX2_X1 U10276 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8954), .S(n9996), .Z(
        P2_U3544) );
  AOI22_X1 U10277 ( .A1(n8897), .A2(n9883), .B1(n9882), .B2(n8896), .ZN(n8901)
         );
  INV_X1 U10278 ( .A(n9532), .ZN(n9905) );
  NAND3_X1 U10279 ( .A1(n8899), .A2(n8898), .A3(n9905), .ZN(n8900) );
  NAND3_X1 U10280 ( .A1(n8902), .A2(n8901), .A3(n8900), .ZN(n8955) );
  MUX2_X1 U10281 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8955), .S(n9996), .Z(
        P2_U3543) );
  AOI22_X1 U10282 ( .A1(n8904), .A2(n9883), .B1(n9882), .B2(n8903), .ZN(n8905)
         );
  OAI211_X1 U10283 ( .C1(n8907), .C2(n9532), .A(n8906), .B(n8905), .ZN(n8956)
         );
  MUX2_X1 U10284 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n8956), .S(n9996), .Z(
        P2_U3542) );
  AOI22_X1 U10285 ( .A1(n8909), .A2(n9883), .B1(n9882), .B2(n8908), .ZN(n8910)
         );
  OAI211_X1 U10286 ( .C1(n8912), .C2(n9532), .A(n8911), .B(n8910), .ZN(n8957)
         );
  MUX2_X1 U10287 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n8957), .S(n9996), .Z(
        P2_U3541) );
  AOI22_X1 U10288 ( .A1(n8914), .A2(n9883), .B1(n9882), .B2(n8913), .ZN(n8915)
         );
  OAI211_X1 U10289 ( .C1(n8917), .C2(n9532), .A(n8916), .B(n8915), .ZN(n8958)
         );
  MUX2_X1 U10290 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n8958), .S(n9996), .Z(
        P2_U3540) );
  AOI211_X1 U10291 ( .C1(n9882), .C2(n8920), .A(n8919), .B(n8918), .ZN(n8921)
         );
  OAI21_X1 U10292 ( .B1(n9532), .B2(n8922), .A(n8921), .ZN(n8959) );
  MUX2_X1 U10293 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8959), .S(n9996), .Z(
        P2_U3539) );
  AOI22_X1 U10294 ( .A1(n8924), .A2(n9883), .B1(n9882), .B2(n8923), .ZN(n8925)
         );
  OAI211_X1 U10295 ( .C1(n8927), .C2(n9532), .A(n8926), .B(n8925), .ZN(n8960)
         );
  MUX2_X1 U10296 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n8960), .S(n9996), .Z(
        P2_U3538) );
  INV_X1 U10297 ( .A(n8928), .ZN(n8933) );
  AOI21_X1 U10298 ( .B1(n9882), .B2(n8930), .A(n8929), .ZN(n8931) );
  OAI211_X1 U10299 ( .C1(n8933), .C2(n9532), .A(n8932), .B(n8931), .ZN(n8961)
         );
  MUX2_X1 U10300 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8961), .S(n9996), .Z(
        P2_U3537) );
  OAI22_X1 U10301 ( .A1(n8935), .A2(n9901), .B1(n8934), .B2(n9899), .ZN(n8937)
         );
  AOI211_X1 U10302 ( .C1(n8938), .C2(n9905), .A(n8937), .B(n8936), .ZN(n8939)
         );
  INV_X1 U10303 ( .A(n8939), .ZN(n8962) );
  MUX2_X1 U10304 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8962), .S(n9996), .Z(
        P2_U3536) );
  OAI22_X1 U10305 ( .A1(n8941), .A2(n9901), .B1(n8940), .B2(n9899), .ZN(n8942)
         );
  INV_X1 U10306 ( .A(n8942), .ZN(n8943) );
  OAI21_X1 U10307 ( .B1(n8944), .B2(n9886), .A(n8943), .ZN(n8945) );
  OR2_X1 U10308 ( .A1(n8946), .A2(n8945), .ZN(n8963) );
  MUX2_X1 U10309 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n8963), .S(n9996), .Z(
        P2_U3533) );
  MUX2_X1 U10310 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n8947), .S(n9909), .Z(
        P2_U3519) );
  MUX2_X1 U10311 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n8948), .S(n9909), .Z(
        P2_U3518) );
  MUX2_X1 U10312 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n8950), .S(n9909), .Z(
        P2_U3516) );
  MUX2_X1 U10313 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8951), .S(n9909), .Z(
        P2_U3515) );
  MUX2_X1 U10314 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n8952), .S(n9909), .Z(
        P2_U3514) );
  MUX2_X1 U10315 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n8953), .S(n9909), .Z(
        P2_U3513) );
  MUX2_X1 U10316 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n8954), .S(n9909), .Z(
        P2_U3512) );
  MUX2_X1 U10317 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n8955), .S(n9909), .Z(
        P2_U3511) );
  MUX2_X1 U10318 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n8956), .S(n9909), .Z(
        P2_U3510) );
  MUX2_X1 U10319 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n8957), .S(n9909), .Z(
        P2_U3509) );
  MUX2_X1 U10320 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n8958), .S(n9909), .Z(
        P2_U3508) );
  MUX2_X1 U10321 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n8959), .S(n9909), .Z(
        P2_U3507) );
  MUX2_X1 U10322 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n8960), .S(n9909), .Z(
        P2_U3505) );
  MUX2_X1 U10323 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n8961), .S(n9909), .Z(
        P2_U3502) );
  MUX2_X1 U10324 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n8962), .S(n9909), .Z(
        P2_U3499) );
  MUX2_X1 U10325 ( .A(n8963), .B(P2_REG0_REG_13__SCAN_IN), .S(n9907), .Z(
        P2_U3490) );
  INV_X1 U10326 ( .A(n8964), .ZN(n9461) );
  INV_X1 U10327 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n10164) );
  NAND2_X1 U10328 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n10164), .ZN(n8966) );
  NOR3_X1 U10329 ( .A1(n8967), .A2(n8966), .A3(P2_U3152), .ZN(n8968) );
  AOI21_X1 U10330 ( .B1(n8970), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n8968), .ZN(
        n8969) );
  OAI21_X1 U10331 ( .B1(n9461), .B2(n8973), .A(n8969), .ZN(P2_U3327) );
  AOI22_X1 U10332 ( .A1(n8971), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n8970), .ZN(n8972) );
  OAI21_X1 U10333 ( .B1(n8974), .B2(n8973), .A(n8972), .ZN(P2_U3328) );
  INV_X1 U10334 ( .A(n8975), .ZN(n8976) );
  MUX2_X1 U10335 ( .A(n8976), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  NAND2_X1 U10336 ( .A1(n4487), .A2(n8977), .ZN(n8979) );
  XNOR2_X1 U10337 ( .A(n8979), .B(n8978), .ZN(n8984) );
  AOI22_X1 U10338 ( .A1(n9259), .A2(n9067), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3084), .ZN(n8981) );
  NAND2_X1 U10339 ( .A1(n9258), .A2(n9068), .ZN(n8980) );
  OAI211_X1 U10340 ( .C1(n9071), .C2(n9266), .A(n8981), .B(n8980), .ZN(n8982)
         );
  AOI21_X1 U10341 ( .B1(n9407), .B2(n9037), .A(n8982), .ZN(n8983) );
  OAI21_X1 U10342 ( .B1(n8984), .B2(n9075), .A(n8983), .ZN(P1_U3214) );
  XOR2_X1 U10343 ( .A(n8987), .B(n8986), .Z(n8988) );
  XNOR2_X1 U10344 ( .A(n8985), .B(n8988), .ZN(n8994) );
  NOR2_X1 U10345 ( .A1(n10119), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9102) );
  AOI21_X1 U10346 ( .B1(n9067), .B2(n9327), .A(n9102), .ZN(n8990) );
  NAND2_X1 U10347 ( .A1(n9049), .A2(n9319), .ZN(n8989) );
  OAI211_X1 U10348 ( .C1(n8991), .C2(n9058), .A(n8990), .B(n8989), .ZN(n8992)
         );
  AOI21_X1 U10349 ( .B1(n9425), .B2(n9037), .A(n8992), .ZN(n8993) );
  OAI21_X1 U10350 ( .B1(n8994), .B2(n9075), .A(n8993), .ZN(P1_U3217) );
  XOR2_X1 U10351 ( .A(n8996), .B(n8995), .Z(n9001) );
  AOI22_X1 U10352 ( .A1(n9068), .A2(n9327), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3084), .ZN(n8998) );
  NAND2_X1 U10353 ( .A1(n9049), .A2(n9295), .ZN(n8997) );
  OAI211_X1 U10354 ( .C1(n9291), .C2(n9014), .A(n8998), .B(n8997), .ZN(n8999)
         );
  AOI21_X1 U10355 ( .B1(n9417), .B2(n9037), .A(n8999), .ZN(n9000) );
  OAI21_X1 U10356 ( .B1(n9001), .B2(n9075), .A(n9000), .ZN(P1_U3221) );
  XOR2_X1 U10357 ( .A(n9003), .B(n9002), .Z(n9008) );
  NAND2_X1 U10358 ( .A1(n9232), .A2(n9067), .ZN(n9005) );
  AOI22_X1 U10359 ( .A1(n9259), .A2(n9068), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3084), .ZN(n9004) );
  OAI211_X1 U10360 ( .C1(n9071), .C2(n9225), .A(n9005), .B(n9004), .ZN(n9006)
         );
  AOI21_X1 U10361 ( .B1(n9395), .B2(n9073), .A(n9006), .ZN(n9007) );
  OAI21_X1 U10362 ( .B1(n9008), .B2(n9075), .A(n9007), .ZN(P1_U3223) );
  AOI21_X1 U10363 ( .B1(n9011), .B2(n9010), .A(n9009), .ZN(n9017) );
  AOI22_X1 U10364 ( .A1(n9280), .A2(n9068), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3084), .ZN(n9013) );
  NAND2_X1 U10365 ( .A1(n9247), .A2(n9049), .ZN(n9012) );
  OAI211_X1 U10366 ( .C1(n9245), .C2(n9014), .A(n9013), .B(n9012), .ZN(n9015)
         );
  AOI21_X1 U10367 ( .B1(n9402), .B2(n9037), .A(n9015), .ZN(n9016) );
  OAI21_X1 U10368 ( .B1(n9017), .B2(n9075), .A(n9016), .ZN(P1_U3227) );
  OAI21_X1 U10369 ( .B1(n9020), .B2(n9019), .A(n9018), .ZN(n9021) );
  NAND2_X1 U10370 ( .A1(n9021), .A2(n5747), .ZN(n9027) );
  NOR2_X1 U10371 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10215), .ZN(n9621) );
  AOI21_X1 U10372 ( .B1(n9037), .B2(n9022), .A(n9621), .ZN(n9026) );
  AOI22_X1 U10373 ( .A1(n9067), .A2(n9086), .B1(n9068), .B2(n9088), .ZN(n9025)
         );
  NAND2_X1 U10374 ( .A1(n9049), .A2(n9023), .ZN(n9024) );
  NAND4_X1 U10375 ( .A1(n9027), .A2(n9026), .A3(n9025), .A4(n9024), .ZN(
        P1_U3228) );
  INV_X1 U10376 ( .A(n9028), .ZN(n9033) );
  NAND2_X1 U10377 ( .A1(n4925), .A2(n9032), .ZN(n9030) );
  AOI22_X1 U10378 ( .A1(n9033), .A2(n9032), .B1(n9031), .B2(n9030), .ZN(n9039)
         );
  AOI22_X1 U10379 ( .A1(n9310), .A2(n9067), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3084), .ZN(n9035) );
  NAND2_X1 U10380 ( .A1(n9068), .A2(n9309), .ZN(n9034) );
  OAI211_X1 U10381 ( .C1(n9071), .C2(n9303), .A(n9035), .B(n9034), .ZN(n9036)
         );
  AOI21_X1 U10382 ( .B1(n9420), .B2(n9037), .A(n9036), .ZN(n9038) );
  OAI21_X1 U10383 ( .B1(n9039), .B2(n9075), .A(n9038), .ZN(P1_U3231) );
  INV_X1 U10384 ( .A(n9410), .ZN(n9277) );
  INV_X1 U10385 ( .A(n9043), .ZN(n9041) );
  NOR2_X1 U10386 ( .A1(n9040), .A2(n9041), .ZN(n9046) );
  AOI21_X1 U10387 ( .B1(n9044), .B2(n9043), .A(n9042), .ZN(n9045) );
  OAI21_X1 U10388 ( .B1(n9046), .B2(n9045), .A(n5747), .ZN(n9051) );
  AOI22_X1 U10389 ( .A1(n9280), .A2(n9067), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3084), .ZN(n9047) );
  OAI21_X1 U10390 ( .B1(n9124), .B2(n9058), .A(n9047), .ZN(n9048) );
  AOI21_X1 U10391 ( .B1(n9275), .B2(n9049), .A(n9048), .ZN(n9050) );
  OAI211_X1 U10392 ( .C1(n9277), .C2(n9063), .A(n9051), .B(n9050), .ZN(
        P1_U3233) );
  INV_X1 U10393 ( .A(n9432), .ZN(n9334) );
  AOI21_X1 U10394 ( .B1(n9055), .B2(n9054), .A(n9053), .ZN(n9056) );
  NOR2_X1 U10395 ( .A1(n9056), .A2(n9075), .ZN(n9057) );
  OAI21_X1 U10396 ( .B1(n4677), .B2(n9052), .A(n9057), .ZN(n9062) );
  NOR2_X1 U10397 ( .A1(n9071), .A2(n9335), .ZN(n9060) );
  NAND2_X1 U10398 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9683) );
  OAI21_X1 U10399 ( .B1(n9058), .B2(n9345), .A(n9683), .ZN(n9059) );
  AOI211_X1 U10400 ( .C1(n9067), .C2(n9309), .A(n9060), .B(n9059), .ZN(n9061)
         );
  OAI211_X1 U10401 ( .C1(n9334), .C2(n9063), .A(n9062), .B(n9061), .ZN(
        P1_U3236) );
  NAND2_X1 U10402 ( .A1(n4433), .A2(n9064), .ZN(n9065) );
  XNOR2_X1 U10403 ( .A(n9066), .B(n9065), .ZN(n9076) );
  NAND2_X1 U10404 ( .A1(n9217), .A2(n9067), .ZN(n9070) );
  AOI22_X1 U10405 ( .A1(n9216), .A2(n9068), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3084), .ZN(n9069) );
  OAI211_X1 U10406 ( .C1(n9071), .C2(n9207), .A(n9070), .B(n9069), .ZN(n9072)
         );
  AOI21_X1 U10407 ( .B1(n9391), .B2(n9073), .A(n9072), .ZN(n9074) );
  OAI21_X1 U10408 ( .B1(n9076), .B2(n9075), .A(n9074), .ZN(P1_U3238) );
  MUX2_X1 U10409 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9077), .S(P1_U4006), .Z(
        P1_U3585) );
  MUX2_X1 U10410 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9078), .S(P1_U4006), .Z(
        P1_U3584) );
  MUX2_X1 U10411 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9217), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U10412 ( .A(n9232), .B(P1_DATAO_REG_26__SCAN_IN), .S(n9089), .Z(
        P1_U3581) );
  MUX2_X1 U10413 ( .A(n9216), .B(P1_DATAO_REG_25__SCAN_IN), .S(n9089), .Z(
        P1_U3580) );
  MUX2_X1 U10414 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9259), .S(P1_U4006), .Z(
        P1_U3579) );
  MUX2_X1 U10415 ( .A(n9280), .B(P1_DATAO_REG_23__SCAN_IN), .S(n9089), .Z(
        P1_U3578) );
  MUX2_X1 U10416 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9258), .S(P1_U4006), .Z(
        P1_U3577) );
  MUX2_X1 U10417 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9310), .S(P1_U4006), .Z(
        P1_U3576) );
  MUX2_X1 U10418 ( .A(n9327), .B(P1_DATAO_REG_20__SCAN_IN), .S(n9089), .Z(
        P1_U3575) );
  MUX2_X1 U10419 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9309), .S(P1_U4006), .Z(
        P1_U3574) );
  MUX2_X1 U10420 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9362), .S(P1_U4006), .Z(
        P1_U3573) );
  MUX2_X1 U10421 ( .A(n9539), .B(P1_DATAO_REG_17__SCAN_IN), .S(n9089), .Z(
        P1_U3572) );
  MUX2_X1 U10422 ( .A(n9361), .B(P1_DATAO_REG_16__SCAN_IN), .S(n9089), .Z(
        P1_U3571) );
  MUX2_X1 U10423 ( .A(n9538), .B(P1_DATAO_REG_15__SCAN_IN), .S(n9089), .Z(
        P1_U3570) );
  MUX2_X1 U10424 ( .A(n9079), .B(P1_DATAO_REG_14__SCAN_IN), .S(n9089), .Z(
        P1_U3569) );
  MUX2_X1 U10425 ( .A(n9080), .B(P1_DATAO_REG_13__SCAN_IN), .S(n9089), .Z(
        P1_U3568) );
  MUX2_X1 U10426 ( .A(n9081), .B(P1_DATAO_REG_12__SCAN_IN), .S(n9089), .Z(
        P1_U3567) );
  MUX2_X1 U10427 ( .A(n9496), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9089), .Z(
        P1_U3566) );
  MUX2_X1 U10428 ( .A(n9082), .B(P1_DATAO_REG_10__SCAN_IN), .S(n9089), .Z(
        P1_U3565) );
  MUX2_X1 U10429 ( .A(n9497), .B(P1_DATAO_REG_9__SCAN_IN), .S(n9089), .Z(
        P1_U3564) );
  MUX2_X1 U10430 ( .A(n9083), .B(P1_DATAO_REG_8__SCAN_IN), .S(n9089), .Z(
        P1_U3563) );
  MUX2_X1 U10431 ( .A(n9084), .B(P1_DATAO_REG_7__SCAN_IN), .S(n9089), .Z(
        P1_U3562) );
  MUX2_X1 U10432 ( .A(n9085), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9089), .Z(
        P1_U3561) );
  MUX2_X1 U10433 ( .A(n9086), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9089), .Z(
        P1_U3560) );
  MUX2_X1 U10434 ( .A(n9087), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9089), .Z(
        P1_U3559) );
  MUX2_X1 U10435 ( .A(n9088), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9089), .Z(
        P1_U3558) );
  MUX2_X1 U10436 ( .A(n9712), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9089), .Z(
        P1_U3557) );
  MUX2_X1 U10437 ( .A(n5011), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9089), .Z(
        P1_U3556) );
  AOI21_X1 U10438 ( .B1(n9095), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9090), .ZN(
        n9689) );
  INV_X1 U10439 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n10013) );
  AOI22_X1 U10440 ( .A1(n9685), .A2(n10013), .B1(P1_REG2_REG_18__SCAN_IN), 
        .B2(n9092), .ZN(n9688) );
  NOR2_X1 U10441 ( .A1(n9689), .A2(n9688), .ZN(n9687) );
  AOI21_X1 U10442 ( .B1(P1_REG2_REG_18__SCAN_IN), .B2(n9685), .A(n9687), .ZN(
        n9091) );
  XNOR2_X1 U10443 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n9091), .ZN(n9101) );
  INV_X1 U10444 ( .A(n9101), .ZN(n9097) );
  INV_X1 U10445 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9093) );
  AOI22_X1 U10446 ( .A1(n9685), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n9093), .B2(
        n9092), .ZN(n9692) );
  AOI21_X1 U10447 ( .B1(n9095), .B2(P1_REG1_REG_17__SCAN_IN), .A(n9094), .ZN(
        n9691) );
  NAND2_X1 U10448 ( .A1(n9692), .A2(n9691), .ZN(n9690) );
  OAI21_X1 U10449 ( .B1(n9685), .B2(P1_REG1_REG_18__SCAN_IN), .A(n9690), .ZN(
        n9096) );
  XOR2_X1 U10450 ( .A(n9096), .B(P1_REG1_REG_19__SCAN_IN), .Z(n9098) );
  AOI21_X1 U10451 ( .B1(n9098), .B2(n9694), .A(n9686), .ZN(n9099) );
  INV_X1 U10452 ( .A(n9385), .ZN(n9194) );
  INV_X1 U10453 ( .A(n9395), .ZN(n9228) );
  NOR2_X1 U10454 ( .A1(n9547), .A2(n9544), .ZN(n9352) );
  NAND2_X1 U10455 ( .A1(n9352), .A2(n9358), .ZN(n9353) );
  INV_X1 U10456 ( .A(n9425), .ZN(n9321) );
  NAND2_X1 U10457 ( .A1(n9333), .A2(n9321), .ZN(n9316) );
  INV_X1 U10458 ( .A(n9417), .ZN(n9298) );
  NAND2_X1 U10459 ( .A1(n9302), .A2(n9298), .ZN(n9292) );
  NAND2_X1 U10460 ( .A1(n9194), .A2(n9206), .ZN(n9189) );
  NAND2_X1 U10461 ( .A1(n9161), .A2(n9178), .ZN(n9160) );
  NOR2_X1 U10462 ( .A1(n9111), .A2(n9160), .ZN(n9110) );
  XNOR2_X1 U10463 ( .A(n9107), .B(n9110), .ZN(n9372) );
  INV_X1 U10464 ( .A(P1_B_REG_SCAN_IN), .ZN(n9103) );
  NOR2_X1 U10465 ( .A1(n9104), .A2(n9103), .ZN(n9105) );
  OR2_X1 U10466 ( .A1(n9348), .A2(n9105), .ZN(n9159) );
  NOR2_X1 U10467 ( .A1(n9106), .A2(n9159), .ZN(n9369) );
  INV_X1 U10468 ( .A(n9369), .ZN(n9555) );
  NOR2_X1 U10469 ( .A1(n9728), .A2(n9555), .ZN(n9112) );
  NOR2_X1 U10470 ( .A1(n9107), .A2(n9357), .ZN(n9108) );
  AOI211_X1 U10471 ( .C1(n9728), .C2(P1_REG2_REG_31__SCAN_IN), .A(n9112), .B(
        n9108), .ZN(n9109) );
  OAI21_X1 U10472 ( .B1(n9372), .B2(n9166), .A(n9109), .ZN(P1_U3261) );
  INV_X1 U10473 ( .A(n9111), .ZN(n9556) );
  AOI21_X1 U10474 ( .B1(n9111), .B2(n9160), .A(n9110), .ZN(n9558) );
  NAND2_X1 U10475 ( .A1(n9558), .A2(n9366), .ZN(n9114) );
  AOI21_X1 U10476 ( .B1(n9728), .B2(P1_REG2_REG_30__SCAN_IN), .A(n9112), .ZN(
        n9113) );
  OAI211_X1 U10477 ( .C1(n9556), .C2(n9357), .A(n9114), .B(n9113), .ZN(
        P1_U3262) );
  INV_X1 U10478 ( .A(n9115), .ZN(n9118) );
  NOR2_X1 U10479 ( .A1(n9435), .A2(n9539), .ZN(n9120) );
  AOI22_X1 U10480 ( .A1(n9332), .A2(n9342), .B1(n9362), .B2(n9432), .ZN(n9315)
         );
  NOR2_X1 U10481 ( .A1(n9425), .A2(n9309), .ZN(n9121) );
  OAI22_X1 U10482 ( .A1(n9315), .A2(n9121), .B1(n9347), .B2(n9321), .ZN(n9301)
         );
  INV_X1 U10483 ( .A(n9420), .ZN(n9306) );
  NAND2_X1 U10484 ( .A1(n9277), .A2(n9291), .ZN(n9125) );
  NOR2_X1 U10485 ( .A1(n9407), .A2(n9280), .ZN(n9126) );
  INV_X1 U10486 ( .A(n9402), .ZN(n9250) );
  NAND2_X1 U10487 ( .A1(n9250), .A2(n9128), .ZN(n9130) );
  NAND2_X1 U10488 ( .A1(n9210), .A2(n9131), .ZN(n9132) );
  NAND2_X1 U10489 ( .A1(n9202), .A2(n9132), .ZN(n9187) );
  NAND2_X1 U10490 ( .A1(n9187), .A2(n9196), .ZN(n9186) );
  NAND2_X1 U10491 ( .A1(n9194), .A2(n9176), .ZN(n9133) );
  NAND2_X1 U10492 ( .A1(n9186), .A2(n9133), .ZN(n9170) );
  INV_X1 U10493 ( .A(n9170), .ZN(n9134) );
  NAND2_X1 U10494 ( .A1(n9179), .A2(n9197), .ZN(n9135) );
  NAND2_X1 U10495 ( .A1(n9172), .A2(n9135), .ZN(n9136) );
  XNOR2_X1 U10496 ( .A(n9136), .B(n9153), .ZN(n9373) );
  INV_X1 U10497 ( .A(n9373), .ZN(n9169) );
  INV_X1 U10498 ( .A(n9534), .ZN(n9137) );
  NAND2_X1 U10499 ( .A1(n9536), .A2(n9139), .ZN(n9360) );
  NAND2_X1 U10500 ( .A1(n9278), .A2(n9146), .ZN(n9257) );
  INV_X1 U10501 ( .A(n9153), .ZN(n9154) );
  XNOR2_X1 U10502 ( .A(n9155), .B(n9154), .ZN(n9156) );
  OAI222_X1 U10503 ( .A1(n9159), .A2(n9158), .B1(n9346), .B2(n9157), .C1(n9499), .C2(n9156), .ZN(n9375) );
  INV_X1 U10504 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n9162) );
  OAI22_X1 U10505 ( .A1(n9163), .A2(n9708), .B1(n9162), .B2(n9725), .ZN(n9164)
         );
  AOI21_X1 U10506 ( .B1(n9376), .B2(n9543), .A(n9164), .ZN(n9165) );
  OAI21_X1 U10507 ( .B1(n9374), .B2(n9166), .A(n9165), .ZN(n9167) );
  AOI21_X1 U10508 ( .B1(n9375), .B2(n9725), .A(n9167), .ZN(n9168) );
  OAI21_X1 U10509 ( .B1(n9169), .B2(n9368), .A(n9168), .ZN(P1_U3355) );
  NAND2_X1 U10510 ( .A1(n9170), .A2(n9173), .ZN(n9171) );
  INV_X1 U10511 ( .A(n9378), .ZN(n9185) );
  XNOR2_X1 U10512 ( .A(n9174), .B(n9173), .ZN(n9175) );
  OAI222_X1 U10513 ( .A1(n9348), .A2(n9177), .B1(n9346), .B2(n9176), .C1(n9499), .C2(n9175), .ZN(n9380) );
  INV_X1 U10514 ( .A(n9179), .ZN(n9379) );
  AOI21_X1 U10515 ( .B1(n9179), .B2(n9189), .A(n9178), .ZN(n9382) );
  NAND2_X1 U10516 ( .A1(n9382), .A2(n9366), .ZN(n9182) );
  AOI22_X1 U10517 ( .A1(n9180), .A2(n9541), .B1(P1_REG2_REG_28__SCAN_IN), .B2(
        n9728), .ZN(n9181) );
  OAI211_X1 U10518 ( .C1(n9379), .C2(n9357), .A(n9182), .B(n9181), .ZN(n9183)
         );
  AOI21_X1 U10519 ( .B1(n9380), .B2(n9725), .A(n9183), .ZN(n9184) );
  OAI21_X1 U10520 ( .B1(n9185), .B2(n9368), .A(n9184), .ZN(P1_U3263) );
  OAI21_X1 U10521 ( .B1(n9187), .B2(n9196), .A(n9186), .ZN(n9188) );
  INV_X1 U10522 ( .A(n9188), .ZN(n9389) );
  INV_X1 U10523 ( .A(n9206), .ZN(n9191) );
  INV_X1 U10524 ( .A(n9189), .ZN(n9190) );
  AOI21_X1 U10525 ( .B1(n9385), .B2(n9191), .A(n9190), .ZN(n9386) );
  AOI22_X1 U10526 ( .A1(n9192), .A2(n9541), .B1(P1_REG2_REG_27__SCAN_IN), .B2(
        n9728), .ZN(n9193) );
  OAI21_X1 U10527 ( .B1(n9194), .B2(n9357), .A(n9193), .ZN(n9200) );
  XOR2_X1 U10528 ( .A(n9196), .B(n9195), .Z(n9198) );
  AOI222_X1 U10529 ( .A1(n9717), .A2(n9198), .B1(n9197), .B2(n9711), .C1(n9232), .C2(n9713), .ZN(n9388) );
  NOR2_X1 U10530 ( .A1(n9388), .A2(n9728), .ZN(n9199) );
  AOI211_X1 U10531 ( .C1(n9386), .C2(n9366), .A(n9200), .B(n9199), .ZN(n9201)
         );
  OAI21_X1 U10532 ( .B1(n9389), .B2(n9368), .A(n9201), .ZN(P1_U3264) );
  OAI21_X1 U10533 ( .B1(n9204), .B2(n9203), .A(n9202), .ZN(n9205) );
  INV_X1 U10534 ( .A(n9205), .ZN(n9394) );
  AOI211_X1 U10535 ( .C1(n9391), .C2(n9223), .A(n9788), .B(n9206), .ZN(n9390)
         );
  NOR2_X1 U10536 ( .A1(n9728), .A2(n5505), .ZN(n9338) );
  INV_X1 U10537 ( .A(n9207), .ZN(n9208) );
  AOI22_X1 U10538 ( .A1(n9208), .A2(n9541), .B1(P1_REG2_REG_26__SCAN_IN), .B2(
        n9728), .ZN(n9209) );
  OAI21_X1 U10539 ( .B1(n9210), .B2(n9357), .A(n9209), .ZN(n9220) );
  AND2_X1 U10540 ( .A1(n9212), .A2(n9211), .ZN(n9215) );
  OAI21_X1 U10541 ( .B1(n9215), .B2(n9214), .A(n9213), .ZN(n9218) );
  AOI222_X1 U10542 ( .A1(n9717), .A2(n9218), .B1(n9217), .B2(n9711), .C1(n9216), .C2(n9713), .ZN(n9393) );
  NOR2_X1 U10543 ( .A1(n9393), .A2(n9728), .ZN(n9219) );
  AOI211_X1 U10544 ( .C1(n9390), .C2(n9338), .A(n9220), .B(n9219), .ZN(n9221)
         );
  OAI21_X1 U10545 ( .B1(n9394), .B2(n9368), .A(n9221), .ZN(P1_U3265) );
  XOR2_X1 U10546 ( .A(n9231), .B(n9222), .Z(n9399) );
  INV_X1 U10547 ( .A(n9223), .ZN(n9224) );
  AOI21_X1 U10548 ( .B1(n9395), .B2(n4531), .A(n9224), .ZN(n9396) );
  INV_X1 U10549 ( .A(n9225), .ZN(n9226) );
  AOI22_X1 U10550 ( .A1(n9226), .A2(n9541), .B1(P1_REG2_REG_25__SCAN_IN), .B2(
        n9728), .ZN(n9227) );
  OAI21_X1 U10551 ( .B1(n9228), .B2(n9357), .A(n9227), .ZN(n9235) );
  NAND2_X1 U10552 ( .A1(n9238), .A2(n9229), .ZN(n9230) );
  XOR2_X1 U10553 ( .A(n9231), .B(n9230), .Z(n9233) );
  AOI222_X1 U10554 ( .A1(n9717), .A2(n9233), .B1(n9232), .B2(n9711), .C1(n9259), .C2(n9713), .ZN(n9398) );
  NOR2_X1 U10555 ( .A1(n9398), .A2(n9728), .ZN(n9234) );
  AOI211_X1 U10556 ( .C1(n9396), .C2(n9366), .A(n9235), .B(n9234), .ZN(n9236)
         );
  OAI21_X1 U10557 ( .B1(n9399), .B2(n9368), .A(n9236), .ZN(P1_U3266) );
  XOR2_X1 U10558 ( .A(n9239), .B(n9237), .Z(n9404) );
  INV_X1 U10559 ( .A(n9238), .ZN(n9242) );
  AOI21_X1 U10560 ( .B1(n9254), .B2(n9240), .A(n9239), .ZN(n9241) );
  NOR2_X1 U10561 ( .A1(n9242), .A2(n9241), .ZN(n9243) );
  OAI222_X1 U10562 ( .A1(n9348), .A2(n9245), .B1(n9346), .B2(n9244), .C1(n9499), .C2(n9243), .ZN(n9400) );
  AOI211_X1 U10563 ( .C1(n9402), .C2(n9263), .A(n9788), .B(n9246), .ZN(n9401)
         );
  NAND2_X1 U10564 ( .A1(n9401), .A2(n9338), .ZN(n9249) );
  AOI22_X1 U10565 ( .A1(n9247), .A2(n9541), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n9728), .ZN(n9248) );
  OAI211_X1 U10566 ( .C1(n9250), .C2(n9357), .A(n9249), .B(n9248), .ZN(n9251)
         );
  AOI21_X1 U10567 ( .B1(n9400), .B2(n9725), .A(n9251), .ZN(n9252) );
  OAI21_X1 U10568 ( .B1(n9404), .B2(n9368), .A(n9252), .ZN(P1_U3267) );
  XNOR2_X1 U10569 ( .A(n9253), .B(n9255), .ZN(n9409) );
  NAND2_X1 U10570 ( .A1(n9254), .A2(n9717), .ZN(n9262) );
  AOI21_X1 U10571 ( .B1(n9257), .B2(n9256), .A(n9255), .ZN(n9261) );
  AOI22_X1 U10572 ( .A1(n9259), .A2(n9711), .B1(n9713), .B2(n9258), .ZN(n9260)
         );
  OAI21_X1 U10573 ( .B1(n9262), .B2(n9261), .A(n9260), .ZN(n9405) );
  INV_X1 U10574 ( .A(n9274), .ZN(n9265) );
  INV_X1 U10575 ( .A(n9263), .ZN(n9264) );
  AOI211_X1 U10576 ( .C1(n9407), .C2(n9265), .A(n9788), .B(n9264), .ZN(n9406)
         );
  NAND2_X1 U10577 ( .A1(n9406), .A2(n9338), .ZN(n9269) );
  INV_X1 U10578 ( .A(n9266), .ZN(n9267) );
  AOI22_X1 U10579 ( .A1(n9267), .A2(n9541), .B1(n9728), .B2(
        P1_REG2_REG_23__SCAN_IN), .ZN(n9268) );
  OAI211_X1 U10580 ( .C1(n9270), .C2(n9357), .A(n9269), .B(n9268), .ZN(n9271)
         );
  AOI21_X1 U10581 ( .B1(n9405), .B2(n9725), .A(n9271), .ZN(n9272) );
  OAI21_X1 U10582 ( .B1(n9409), .B2(n9368), .A(n9272), .ZN(P1_U3268) );
  XNOR2_X1 U10583 ( .A(n9273), .B(n9279), .ZN(n9414) );
  AOI21_X1 U10584 ( .B1(n9410), .B2(n9292), .A(n9274), .ZN(n9411) );
  AOI22_X1 U10585 ( .A1(n9728), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n9275), .B2(
        n9541), .ZN(n9276) );
  OAI21_X1 U10586 ( .B1(n9277), .B2(n9357), .A(n9276), .ZN(n9283) );
  XOR2_X1 U10587 ( .A(n9279), .B(n9278), .Z(n9281) );
  AOI222_X1 U10588 ( .A1(n9717), .A2(n9281), .B1(n9280), .B2(n9711), .C1(n9310), .C2(n9713), .ZN(n9413) );
  NOR2_X1 U10589 ( .A1(n9413), .A2(n9728), .ZN(n9282) );
  AOI211_X1 U10590 ( .C1(n9411), .C2(n9366), .A(n9283), .B(n9282), .ZN(n9284)
         );
  OAI21_X1 U10591 ( .B1(n9414), .B2(n9368), .A(n9284), .ZN(P1_U3269) );
  OAI21_X1 U10592 ( .B1(n9286), .B2(n9288), .A(n9285), .ZN(n9419) );
  XOR2_X1 U10593 ( .A(n9288), .B(n9287), .Z(n9289) );
  OAI222_X1 U10594 ( .A1(n9348), .A2(n9291), .B1(n9346), .B2(n9290), .C1(n9499), .C2(n9289), .ZN(n9415) );
  INV_X1 U10595 ( .A(n9302), .ZN(n9294) );
  INV_X1 U10596 ( .A(n9292), .ZN(n9293) );
  AOI211_X1 U10597 ( .C1(n9417), .C2(n9294), .A(n9788), .B(n9293), .ZN(n9416)
         );
  NAND2_X1 U10598 ( .A1(n9416), .A2(n9338), .ZN(n9297) );
  AOI22_X1 U10599 ( .A1(n9728), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n9295), .B2(
        n9541), .ZN(n9296) );
  OAI211_X1 U10600 ( .C1(n9298), .C2(n9357), .A(n9297), .B(n9296), .ZN(n9299)
         );
  AOI21_X1 U10601 ( .B1(n9415), .B2(n9725), .A(n9299), .ZN(n9300) );
  OAI21_X1 U10602 ( .B1(n9419), .B2(n9368), .A(n9300), .ZN(P1_U3270) );
  XOR2_X1 U10603 ( .A(n9307), .B(n9301), .Z(n9424) );
  AOI21_X1 U10604 ( .B1(n9420), .B2(n9316), .A(n9302), .ZN(n9421) );
  INV_X1 U10605 ( .A(n9303), .ZN(n9304) );
  AOI22_X1 U10606 ( .A1(n9728), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9304), .B2(
        n9541), .ZN(n9305) );
  OAI21_X1 U10607 ( .B1(n9306), .B2(n9357), .A(n9305), .ZN(n9313) );
  XNOR2_X1 U10608 ( .A(n9308), .B(n9307), .ZN(n9311) );
  AOI222_X1 U10609 ( .A1(n9717), .A2(n9311), .B1(n9310), .B2(n9711), .C1(n9309), .C2(n9713), .ZN(n9423) );
  NOR2_X1 U10610 ( .A1(n9423), .A2(n9728), .ZN(n9312) );
  AOI211_X1 U10611 ( .C1(n9421), .C2(n9366), .A(n9313), .B(n9312), .ZN(n9314)
         );
  OAI21_X1 U10612 ( .B1(n9424), .B2(n9368), .A(n9314), .ZN(P1_U3271) );
  XNOR2_X1 U10613 ( .A(n9315), .B(n9322), .ZN(n9429) );
  INV_X1 U10614 ( .A(n9333), .ZN(n9318) );
  INV_X1 U10615 ( .A(n9316), .ZN(n9317) );
  AOI21_X1 U10616 ( .B1(n9425), .B2(n9318), .A(n9317), .ZN(n9426) );
  AOI22_X1 U10617 ( .A1(n9728), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9319), .B2(
        n9541), .ZN(n9320) );
  OAI21_X1 U10618 ( .B1(n9321), .B2(n9357), .A(n9320), .ZN(n9330) );
  INV_X1 U10619 ( .A(n9322), .ZN(n9324) );
  NAND2_X1 U10620 ( .A1(n9324), .A2(n9323), .ZN(n9326) );
  OAI21_X1 U10621 ( .B1(n4383), .B2(n9326), .A(n9325), .ZN(n9328) );
  AOI222_X1 U10622 ( .A1(n9717), .A2(n9328), .B1(n9327), .B2(n9711), .C1(n9362), .C2(n9713), .ZN(n9428) );
  NOR2_X1 U10623 ( .A1(n9428), .A2(n9728), .ZN(n9329) );
  AOI211_X1 U10624 ( .C1(n9426), .C2(n9366), .A(n9330), .B(n9329), .ZN(n9331)
         );
  OAI21_X1 U10625 ( .B1(n9368), .B2(n9429), .A(n9331), .ZN(P1_U3272) );
  XNOR2_X1 U10626 ( .A(n9332), .B(n9342), .ZN(n9434) );
  AOI211_X1 U10627 ( .C1(n9432), .C2(n9353), .A(n9788), .B(n9333), .ZN(n9431)
         );
  NOR2_X1 U10628 ( .A1(n9334), .A2(n9357), .ZN(n9337) );
  OAI22_X1 U10629 ( .A1(n9725), .A2(n10013), .B1(n9335), .B2(n9708), .ZN(n9336) );
  AOI211_X1 U10630 ( .C1(n9431), .C2(n9338), .A(n9337), .B(n9336), .ZN(n9350)
         );
  INV_X1 U10631 ( .A(n9339), .ZN(n9340) );
  NOR2_X1 U10632 ( .A1(n9341), .A2(n9340), .ZN(n9343) );
  XNOR2_X1 U10633 ( .A(n9343), .B(n9342), .ZN(n9344) );
  OAI222_X1 U10634 ( .A1(n9348), .A2(n9347), .B1(n9346), .B2(n9345), .C1(n9499), .C2(n9344), .ZN(n9430) );
  NAND2_X1 U10635 ( .A1(n9430), .A2(n9725), .ZN(n9349) );
  OAI211_X1 U10636 ( .C1(n9434), .C2(n9368), .A(n9350), .B(n9349), .ZN(
        P1_U3273) );
  XNOR2_X1 U10637 ( .A(n9351), .B(n9359), .ZN(n9441) );
  INV_X1 U10638 ( .A(n9352), .ZN(n9548) );
  INV_X1 U10639 ( .A(n9353), .ZN(n9354) );
  AOI21_X1 U10640 ( .B1(n9435), .B2(n9548), .A(n9354), .ZN(n9437) );
  AOI22_X1 U10641 ( .A1(n9728), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9355), .B2(
        n9541), .ZN(n9356) );
  OAI21_X1 U10642 ( .B1(n9358), .B2(n9357), .A(n9356), .ZN(n9365) );
  XNOR2_X1 U10643 ( .A(n9360), .B(n9359), .ZN(n9363) );
  AOI222_X1 U10644 ( .A1(n9717), .A2(n9363), .B1(n9362), .B2(n9711), .C1(n9361), .C2(n9713), .ZN(n9439) );
  NOR2_X1 U10645 ( .A1(n9439), .A2(n9728), .ZN(n9364) );
  AOI211_X1 U10646 ( .C1(n9437), .C2(n9366), .A(n9365), .B(n9364), .ZN(n9367)
         );
  OAI21_X1 U10647 ( .B1(n9441), .B2(n9368), .A(n9367), .ZN(P1_U3274) );
  AOI21_X1 U10648 ( .B1(n9370), .B2(n9436), .A(n9369), .ZN(n9371) );
  OAI21_X1 U10649 ( .B1(n9372), .B2(n9788), .A(n9371), .ZN(n9442) );
  MUX2_X1 U10650 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9442), .S(n9806), .Z(
        P1_U3554) );
  NAND2_X1 U10651 ( .A1(n9373), .A2(n9783), .ZN(n9377) );
  MUX2_X1 U10652 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9443), .S(n9806), .Z(
        P1_U3552) );
  NAND2_X1 U10653 ( .A1(n9378), .A2(n9783), .ZN(n9384) );
  NOR2_X1 U10654 ( .A1(n9379), .A2(n9787), .ZN(n9381) );
  AOI211_X1 U10655 ( .C1(n9704), .C2(n9382), .A(n9381), .B(n9380), .ZN(n9383)
         );
  NAND2_X1 U10656 ( .A1(n9384), .A2(n9383), .ZN(n9444) );
  MUX2_X1 U10657 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9444), .S(n9806), .Z(
        P1_U3551) );
  AOI22_X1 U10658 ( .A1(n9386), .A2(n9704), .B1(n9436), .B2(n9385), .ZN(n9387)
         );
  OAI211_X1 U10659 ( .C1(n9389), .C2(n9440), .A(n9388), .B(n9387), .ZN(n9445)
         );
  MUX2_X1 U10660 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9445), .S(n9806), .Z(
        P1_U3550) );
  AOI21_X1 U10661 ( .B1(n9436), .B2(n9391), .A(n9390), .ZN(n9392) );
  OAI211_X1 U10662 ( .C1(n9394), .C2(n9440), .A(n9393), .B(n9392), .ZN(n9446)
         );
  MUX2_X1 U10663 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9446), .S(n9806), .Z(
        P1_U3549) );
  AOI22_X1 U10664 ( .A1(n9396), .A2(n9704), .B1(n9436), .B2(n9395), .ZN(n9397)
         );
  OAI211_X1 U10665 ( .C1(n9399), .C2(n9440), .A(n9398), .B(n9397), .ZN(n9447)
         );
  MUX2_X1 U10666 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9447), .S(n9806), .Z(
        P1_U3548) );
  AOI211_X1 U10667 ( .C1(n9436), .C2(n9402), .A(n9401), .B(n9400), .ZN(n9403)
         );
  OAI21_X1 U10668 ( .B1(n9404), .B2(n9440), .A(n9403), .ZN(n9448) );
  MUX2_X1 U10669 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9448), .S(n9806), .Z(
        P1_U3547) );
  AOI211_X1 U10670 ( .C1(n9436), .C2(n9407), .A(n9406), .B(n9405), .ZN(n9408)
         );
  OAI21_X1 U10671 ( .B1(n9409), .B2(n9440), .A(n9408), .ZN(n9449) );
  MUX2_X1 U10672 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9449), .S(n9806), .Z(
        P1_U3546) );
  AOI22_X1 U10673 ( .A1(n9411), .A2(n9704), .B1(n9436), .B2(n9410), .ZN(n9412)
         );
  OAI211_X1 U10674 ( .C1(n9414), .C2(n9440), .A(n9413), .B(n9412), .ZN(n9450)
         );
  MUX2_X1 U10675 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9450), .S(n9806), .Z(
        P1_U3545) );
  AOI211_X1 U10676 ( .C1(n9436), .C2(n9417), .A(n9416), .B(n9415), .ZN(n9418)
         );
  OAI21_X1 U10677 ( .B1(n9419), .B2(n9440), .A(n9418), .ZN(n9451) );
  MUX2_X1 U10678 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9451), .S(n9806), .Z(
        P1_U3544) );
  AOI22_X1 U10679 ( .A1(n9421), .A2(n9704), .B1(n9436), .B2(n9420), .ZN(n9422)
         );
  OAI211_X1 U10680 ( .C1(n9424), .C2(n9440), .A(n9423), .B(n9422), .ZN(n9452)
         );
  MUX2_X1 U10681 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9452), .S(n9806), .Z(
        P1_U3543) );
  AOI22_X1 U10682 ( .A1(n9426), .A2(n9704), .B1(n9436), .B2(n9425), .ZN(n9427)
         );
  OAI211_X1 U10683 ( .C1(n9429), .C2(n9440), .A(n9428), .B(n9427), .ZN(n9453)
         );
  MUX2_X1 U10684 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9453), .S(n9806), .Z(
        P1_U3542) );
  AOI211_X1 U10685 ( .C1(n9436), .C2(n9432), .A(n9431), .B(n9430), .ZN(n9433)
         );
  OAI21_X1 U10686 ( .B1(n9434), .B2(n9440), .A(n9433), .ZN(n9454) );
  MUX2_X1 U10687 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9454), .S(n9806), .Z(
        P1_U3541) );
  AOI22_X1 U10688 ( .A1(n9437), .A2(n9704), .B1(n9436), .B2(n9435), .ZN(n9438)
         );
  OAI211_X1 U10689 ( .C1(n9441), .C2(n9440), .A(n9439), .B(n9438), .ZN(n9455)
         );
  MUX2_X1 U10690 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9455), .S(n9806), .Z(
        P1_U3540) );
  MUX2_X1 U10691 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9442), .S(n9795), .Z(
        P1_U3522) );
  MUX2_X1 U10692 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9443), .S(n9795), .Z(
        P1_U3520) );
  MUX2_X1 U10693 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9444), .S(n9795), .Z(
        P1_U3519) );
  MUX2_X1 U10694 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9445), .S(n9795), .Z(
        P1_U3518) );
  MUX2_X1 U10695 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9446), .S(n9795), .Z(
        P1_U3517) );
  MUX2_X1 U10696 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9447), .S(n9795), .Z(
        P1_U3516) );
  MUX2_X1 U10697 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9448), .S(n9795), .Z(
        P1_U3515) );
  MUX2_X1 U10698 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9449), .S(n9795), .Z(
        P1_U3514) );
  MUX2_X1 U10699 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9450), .S(n9795), .Z(
        P1_U3513) );
  MUX2_X1 U10700 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9451), .S(n9795), .Z(
        P1_U3512) );
  MUX2_X1 U10701 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9452), .S(n9795), .Z(
        P1_U3511) );
  MUX2_X1 U10702 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9453), .S(n9795), .Z(
        P1_U3510) );
  MUX2_X1 U10703 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9454), .S(n9795), .Z(
        P1_U3508) );
  MUX2_X1 U10704 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9455), .S(n9795), .Z(
        P1_U3505) );
  NOR4_X1 U10705 ( .A1(n9457), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3084), .A4(
        n9456), .ZN(n9458) );
  AOI21_X1 U10706 ( .B1(n9459), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9458), .ZN(
        n9460) );
  OAI21_X1 U10707 ( .B1(n9461), .B2(n4370), .A(n9460), .ZN(P1_U3322) );
  AOI22_X1 U10708 ( .A1(n9813), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3152), .ZN(n9476) );
  INV_X1 U10709 ( .A(n9462), .ZN(n9466) );
  NAND2_X1 U10710 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n9463) );
  NAND2_X1 U10711 ( .A1(n9464), .A2(n9463), .ZN(n9465) );
  NAND3_X1 U10712 ( .A1(n9808), .A2(n9466), .A3(n9465), .ZN(n9472) );
  AOI21_X1 U10713 ( .B1(n9469), .B2(n9468), .A(n9467), .ZN(n9470) );
  NAND2_X1 U10714 ( .A1(n9807), .A2(n9470), .ZN(n9471) );
  OAI211_X1 U10715 ( .C1(n9809), .C2(n9473), .A(n9472), .B(n9471), .ZN(n9474)
         );
  INV_X1 U10716 ( .A(n9474), .ZN(n9475) );
  NAND2_X1 U10717 ( .A1(n9476), .A2(n9475), .ZN(P2_U3246) );
  AOI22_X1 U10718 ( .A1(n9813), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n9490) );
  AOI21_X1 U10719 ( .B1(n9479), .B2(n9478), .A(n9477), .ZN(n9480) );
  NAND2_X1 U10720 ( .A1(n9808), .A2(n9480), .ZN(n9486) );
  AOI21_X1 U10721 ( .B1(n9483), .B2(n9482), .A(n9481), .ZN(n9484) );
  NAND2_X1 U10722 ( .A1(n9807), .A2(n9484), .ZN(n9485) );
  OAI211_X1 U10723 ( .C1(n9809), .C2(n9487), .A(n9486), .B(n9485), .ZN(n9488)
         );
  INV_X1 U10724 ( .A(n9488), .ZN(n9489) );
  NAND2_X1 U10725 ( .A1(n9490), .A2(n9489), .ZN(P2_U3247) );
  XNOR2_X1 U10726 ( .A(n9491), .B(n9494), .ZN(n9518) );
  NAND2_X1 U10727 ( .A1(n9493), .A2(n9492), .ZN(n9495) );
  XNOR2_X1 U10728 ( .A(n9495), .B(n9494), .ZN(n9500) );
  AOI22_X1 U10729 ( .A1(n9713), .A2(n9497), .B1(n9496), .B2(n9711), .ZN(n9498)
         );
  OAI21_X1 U10730 ( .B1(n9500), .B2(n9499), .A(n9498), .ZN(n9501) );
  AOI21_X1 U10731 ( .B1(n9518), .B2(n9502), .A(n9501), .ZN(n9515) );
  AOI222_X1 U10732 ( .A1(n9504), .A2(n9543), .B1(n9503), .B2(n9541), .C1(
        P1_REG2_REG_10__SCAN_IN), .C2(n9728), .ZN(n9512) );
  INV_X1 U10733 ( .A(n9504), .ZN(n9514) );
  INV_X1 U10734 ( .A(n9505), .ZN(n9508) );
  INV_X1 U10735 ( .A(n9506), .ZN(n9507) );
  OAI211_X1 U10736 ( .C1(n9514), .C2(n9508), .A(n9507), .B(n9704), .ZN(n9513)
         );
  INV_X1 U10737 ( .A(n9513), .ZN(n9509) );
  AOI22_X1 U10738 ( .A1(n9518), .A2(n9510), .B1(n9550), .B2(n9509), .ZN(n9511)
         );
  OAI211_X1 U10739 ( .C1(n9728), .C2(n9515), .A(n9512), .B(n9511), .ZN(
        P1_U3281) );
  OAI21_X1 U10740 ( .B1(n9514), .B2(n9787), .A(n9513), .ZN(n9517) );
  INV_X1 U10741 ( .A(n9515), .ZN(n9516) );
  AOI211_X1 U10742 ( .C1(n9793), .C2(n9518), .A(n9517), .B(n9516), .ZN(n9520)
         );
  INV_X1 U10743 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n10228) );
  AOI22_X1 U10744 ( .A1(n9795), .A2(n9520), .B1(n10228), .B2(n9794), .ZN(
        P1_U3484) );
  AOI22_X1 U10745 ( .A1(n9806), .A2(n9520), .B1(n9519), .B2(n9803), .ZN(
        P1_U3533) );
  OAI22_X1 U10746 ( .A1(n9522), .A2(n9901), .B1(n4558), .B2(n9899), .ZN(n9524)
         );
  AOI211_X1 U10747 ( .C1(n9905), .C2(n9525), .A(n9524), .B(n9523), .ZN(n9527)
         );
  AOI22_X1 U10748 ( .A1(n9996), .A2(n9527), .B1(n6008), .B2(n9994), .ZN(
        P2_U3535) );
  INV_X1 U10749 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n9526) );
  AOI22_X1 U10750 ( .A1(n9909), .A2(n9527), .B1(n9526), .B2(n9907), .ZN(
        P2_U3496) );
  AOI22_X1 U10751 ( .A1(n9529), .A2(n9883), .B1(n9882), .B2(n9528), .ZN(n9530)
         );
  OAI211_X1 U10752 ( .C1(n9533), .C2(n9532), .A(n9531), .B(n9530), .ZN(n9995)
         );
  MUX2_X1 U10753 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n9995), .S(n9909), .Z(
        P2_U3493) );
  NAND2_X1 U10754 ( .A1(n9535), .A2(n9534), .ZN(n9537) );
  OAI21_X1 U10755 ( .B1(n9138), .B2(n9537), .A(n9536), .ZN(n9540) );
  AOI222_X1 U10756 ( .A1(n9717), .A2(n9540), .B1(n9539), .B2(n9711), .C1(n9538), .C2(n9713), .ZN(n9561) );
  AOI222_X1 U10757 ( .A1(n9544), .A2(n9543), .B1(P1_REG2_REG_16__SCAN_IN), 
        .B2(n9728), .C1(n9542), .C2(n9541), .ZN(n9554) );
  AOI21_X1 U10758 ( .B1(n9546), .B2(n9545), .A(n4436), .ZN(n9564) );
  INV_X1 U10759 ( .A(n9547), .ZN(n9549) );
  OAI211_X1 U10760 ( .C1(n9562), .C2(n9549), .A(n9548), .B(n9704), .ZN(n9560)
         );
  INV_X1 U10761 ( .A(n9560), .ZN(n9551) );
  AOI22_X1 U10762 ( .A1(n9564), .A2(n9552), .B1(n9551), .B2(n9550), .ZN(n9553)
         );
  OAI211_X1 U10763 ( .C1(n9728), .C2(n9561), .A(n9554), .B(n9553), .ZN(
        P1_U3275) );
  OAI21_X1 U10764 ( .B1(n9556), .B2(n9787), .A(n9555), .ZN(n9557) );
  AOI21_X1 U10765 ( .B1(n9558), .B2(n9704), .A(n9557), .ZN(n9590) );
  INV_X1 U10766 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9559) );
  AOI22_X1 U10767 ( .A1(n9806), .A2(n9590), .B1(n9559), .B2(n9803), .ZN(
        P1_U3553) );
  OAI211_X1 U10768 ( .C1(n9562), .C2(n9787), .A(n9561), .B(n9560), .ZN(n9563)
         );
  AOI21_X1 U10769 ( .B1(n9564), .B2(n9783), .A(n9563), .ZN(n9592) );
  AOI22_X1 U10770 ( .A1(n9806), .A2(n9592), .B1(n7893), .B2(n9803), .ZN(
        P1_U3539) );
  OAI22_X1 U10771 ( .A1(n9566), .A2(n9788), .B1(n9565), .B2(n9787), .ZN(n9568)
         );
  AOI211_X1 U10772 ( .C1(n9569), .C2(n9783), .A(n9568), .B(n9567), .ZN(n9593)
         );
  AOI22_X1 U10773 ( .A1(n9806), .A2(n9593), .B1(n9570), .B2(n9803), .ZN(
        P1_U3538) );
  OAI21_X1 U10774 ( .B1(n9572), .B2(n9787), .A(n9571), .ZN(n9573) );
  AOI211_X1 U10775 ( .C1(n9575), .C2(n9783), .A(n9574), .B(n9573), .ZN(n9595)
         );
  AOI22_X1 U10776 ( .A1(n9806), .A2(n9595), .B1(n7395), .B2(n9803), .ZN(
        P1_U3537) );
  OAI22_X1 U10777 ( .A1(n9577), .A2(n9788), .B1(n9576), .B2(n9787), .ZN(n9578)
         );
  AOI21_X1 U10778 ( .B1(n9579), .B2(n9793), .A(n9578), .ZN(n9580) );
  AND2_X1 U10779 ( .A1(n9581), .A2(n9580), .ZN(n9596) );
  AOI22_X1 U10780 ( .A1(n9806), .A2(n9596), .B1(n6966), .B2(n9803), .ZN(
        P1_U3536) );
  OAI22_X1 U10781 ( .A1(n9583), .A2(n9788), .B1(n9582), .B2(n9787), .ZN(n9584)
         );
  AOI21_X1 U10782 ( .B1(n9585), .B2(n9793), .A(n9584), .ZN(n9586) );
  AND2_X1 U10783 ( .A1(n9587), .A2(n9586), .ZN(n9598) );
  AOI22_X1 U10784 ( .A1(n9806), .A2(n9598), .B1(n9588), .B2(n9803), .ZN(
        P1_U3534) );
  INV_X1 U10785 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9589) );
  AOI22_X1 U10786 ( .A1(n9795), .A2(n9590), .B1(n9589), .B2(n9794), .ZN(
        P1_U3521) );
  INV_X1 U10787 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n9591) );
  AOI22_X1 U10788 ( .A1(n9795), .A2(n9592), .B1(n9591), .B2(n9794), .ZN(
        P1_U3502) );
  INV_X1 U10789 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n10200) );
  AOI22_X1 U10790 ( .A1(n9795), .A2(n9593), .B1(n10200), .B2(n9794), .ZN(
        P1_U3499) );
  INV_X1 U10791 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n9594) );
  AOI22_X1 U10792 ( .A1(n9795), .A2(n9595), .B1(n9594), .B2(n9794), .ZN(
        P1_U3496) );
  INV_X1 U10793 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n10199) );
  AOI22_X1 U10794 ( .A1(n9795), .A2(n9596), .B1(n10199), .B2(n9794), .ZN(
        P1_U3493) );
  INV_X1 U10795 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n9597) );
  AOI22_X1 U10796 ( .A1(n9795), .A2(n9598), .B1(n9597), .B2(n9794), .ZN(
        P1_U3487) );
  XNOR2_X1 U10797 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U10798 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  AOI21_X1 U10799 ( .B1(P1_REG1_REG_0__SCAN_IN), .B2(n4670), .A(n9599), .ZN(
        n9600) );
  NOR4_X1 U10800 ( .A1(n9603), .A2(n9602), .A3(n9601), .A4(n9600), .ZN(n9604)
         );
  AOI21_X1 U10801 ( .B1(n9668), .B2(P1_ADDR_REG_0__SCAN_IN), .A(n9604), .ZN(
        n9606) );
  NAND3_X1 U10802 ( .A1(n9694), .A2(n9949), .A3(n10055), .ZN(n9605) );
  OAI211_X1 U10803 ( .C1(P1_STATE_REG_SCAN_IN), .C2(n8218), .A(n9606), .B(
        n9605), .ZN(P1_U3241) );
  INV_X1 U10804 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9625) );
  INV_X1 U10805 ( .A(n9607), .ZN(n9611) );
  INV_X1 U10806 ( .A(n9608), .ZN(n9610) );
  OAI21_X1 U10807 ( .B1(n9611), .B2(n9610), .A(n9609), .ZN(n9614) );
  INV_X1 U10808 ( .A(n9612), .ZN(n9613) );
  AOI22_X1 U10809 ( .A1(n9695), .A2(n9614), .B1(n9686), .B2(n9613), .ZN(n9624)
         );
  NOR2_X1 U10810 ( .A1(n9616), .A2(n9615), .ZN(n9619) );
  OAI21_X1 U10811 ( .B1(n9619), .B2(n9618), .A(n9617), .ZN(n9622) );
  AOI211_X1 U10812 ( .C1(n9694), .C2(n9622), .A(n9621), .B(n9620), .ZN(n9623)
         );
  OAI211_X1 U10813 ( .C1(n9699), .C2(n9625), .A(n9624), .B(n9623), .ZN(
        P1_U3245) );
  OAI21_X1 U10814 ( .B1(n9628), .B2(n9627), .A(n9626), .ZN(n9638) );
  AND2_X1 U10815 ( .A1(n9630), .A2(n9629), .ZN(n9631) );
  OR2_X1 U10816 ( .A1(n9632), .A2(n9631), .ZN(n9635) );
  INV_X1 U10817 ( .A(n9633), .ZN(n9634) );
  OAI21_X1 U10818 ( .B1(n9636), .B2(n9635), .A(n9634), .ZN(n9637) );
  AOI21_X1 U10819 ( .B1(n9695), .B2(n9638), .A(n9637), .ZN(n9641) );
  AOI22_X1 U10820 ( .A1(n9668), .A2(P1_ADDR_REG_5__SCAN_IN), .B1(n9639), .B2(
        n9686), .ZN(n9640) );
  NAND2_X1 U10821 ( .A1(n9641), .A2(n9640), .ZN(P1_U3246) );
  NOR2_X1 U10822 ( .A1(n9643), .A2(n9642), .ZN(n9644) );
  OR3_X1 U10823 ( .A1(n9659), .A2(n9645), .A3(n9644), .ZN(n9651) );
  XNOR2_X1 U10824 ( .A(n9647), .B(n9646), .ZN(n9649) );
  AOI21_X1 U10825 ( .B1(n9694), .B2(n9649), .A(n9648), .ZN(n9650) );
  AND2_X1 U10826 ( .A1(n9651), .A2(n9650), .ZN(n9654) );
  AOI22_X1 U10827 ( .A1(n9668), .A2(P1_ADDR_REG_6__SCAN_IN), .B1(n9652), .B2(
        n9686), .ZN(n9653) );
  NAND2_X1 U10828 ( .A1(n9654), .A2(n9653), .ZN(P1_U3247) );
  NOR2_X1 U10829 ( .A1(n9656), .A2(n9655), .ZN(n9657) );
  OR3_X1 U10830 ( .A1(n9659), .A2(n9658), .A3(n9657), .ZN(n9666) );
  OAI21_X1 U10831 ( .B1(n9662), .B2(n9661), .A(n9660), .ZN(n9664) );
  AOI21_X1 U10832 ( .B1(n9694), .B2(n9664), .A(n9663), .ZN(n9665) );
  AND2_X1 U10833 ( .A1(n9666), .A2(n9665), .ZN(n9670) );
  AOI22_X1 U10834 ( .A1(n9668), .A2(P1_ADDR_REG_9__SCAN_IN), .B1(n9667), .B2(
        n9686), .ZN(n9669) );
  NAND2_X1 U10835 ( .A1(n9670), .A2(n9669), .ZN(P1_U3250) );
  INV_X1 U10836 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n9682) );
  AOI21_X1 U10837 ( .B1(n9686), .B2(n9672), .A(n9671), .ZN(n9681) );
  OAI21_X1 U10838 ( .B1(n9674), .B2(n4403), .A(n9673), .ZN(n9679) );
  OAI21_X1 U10839 ( .B1(n9677), .B2(n9676), .A(n9675), .ZN(n9678) );
  AOI22_X1 U10840 ( .A1(n9679), .A2(n9695), .B1(n9678), .B2(n9694), .ZN(n9680)
         );
  OAI211_X1 U10841 ( .C1(n9699), .C2(n9682), .A(n9681), .B(n9680), .ZN(
        P1_U3252) );
  INV_X1 U10842 ( .A(n9683), .ZN(n9684) );
  AOI21_X1 U10843 ( .B1(n9686), .B2(n9685), .A(n9684), .ZN(n9698) );
  AOI21_X1 U10844 ( .B1(n9689), .B2(n9688), .A(n9687), .ZN(n9696) );
  OAI21_X1 U10845 ( .B1(n9692), .B2(n9691), .A(n9690), .ZN(n9693) );
  AOI22_X1 U10846 ( .A1(n9696), .A2(n9695), .B1(n9694), .B2(n9693), .ZN(n9697)
         );
  OAI211_X1 U10847 ( .C1(n10083), .C2(n9699), .A(n9698), .B(n9697), .ZN(
        P1_U3259) );
  INV_X1 U10848 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n9727) );
  OAI21_X1 U10849 ( .B1(n9702), .B2(n9701), .A(n9700), .ZN(n9722) );
  INV_X1 U10850 ( .A(n9722), .ZN(n9760) );
  OAI211_X1 U10851 ( .C1(n9757), .C2(n9705), .A(n9704), .B(n9703), .ZN(n9756)
         );
  OAI22_X1 U10852 ( .A1(n9708), .A2(n9707), .B1(n9757), .B2(n9706), .ZN(n9709)
         );
  INV_X1 U10853 ( .A(n9709), .ZN(n9710) );
  OAI21_X1 U10854 ( .B1(n9756), .B2(n5505), .A(n9710), .ZN(n9723) );
  AOI22_X1 U10855 ( .A1(n9713), .A2(n6638), .B1(n9712), .B2(n9711), .ZN(n9720)
         );
  OAI21_X1 U10856 ( .B1(n4367), .B2(n9715), .A(n9714), .ZN(n9718) );
  NAND2_X1 U10857 ( .A1(n9718), .A2(n9717), .ZN(n9719) );
  OAI211_X1 U10858 ( .C1(n9722), .C2(n9721), .A(n9720), .B(n9719), .ZN(n9758)
         );
  AOI211_X1 U10859 ( .C1(n9724), .C2(n9760), .A(n9723), .B(n9758), .ZN(n9726)
         );
  AOI22_X1 U10860 ( .A1(n9728), .A2(n9727), .B1(n9726), .B2(n9725), .ZN(
        P1_U3290) );
  NOR2_X1 U10861 ( .A1(n9730), .A2(n9729), .ZN(n9751) );
  CLKBUF_X1 U10862 ( .A(n9751), .Z(n9744) );
  INV_X1 U10863 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n10193) );
  NOR2_X1 U10864 ( .A1(n9744), .A2(n10193), .ZN(P1_U3292) );
  INV_X1 U10865 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n9731) );
  NOR2_X1 U10866 ( .A1(n9744), .A2(n9731), .ZN(P1_U3293) );
  INV_X1 U10867 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n10137) );
  NOR2_X1 U10868 ( .A1(n9744), .A2(n10137), .ZN(P1_U3294) );
  INV_X1 U10869 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n9732) );
  NOR2_X1 U10870 ( .A1(n9744), .A2(n9732), .ZN(P1_U3295) );
  INV_X1 U10871 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n9733) );
  NOR2_X1 U10872 ( .A1(n9744), .A2(n9733), .ZN(P1_U3296) );
  NOR2_X1 U10873 ( .A1(n9744), .A2(n9734), .ZN(P1_U3297) );
  INV_X1 U10874 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n10143) );
  NOR2_X1 U10875 ( .A1(n9744), .A2(n10143), .ZN(P1_U3298) );
  INV_X1 U10876 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n9735) );
  NOR2_X1 U10877 ( .A1(n9744), .A2(n9735), .ZN(P1_U3299) );
  INV_X1 U10878 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n9736) );
  NOR2_X1 U10879 ( .A1(n9744), .A2(n9736), .ZN(P1_U3300) );
  NOR2_X1 U10880 ( .A1(n9744), .A2(n10158), .ZN(P1_U3301) );
  INV_X1 U10881 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n9737) );
  NOR2_X1 U10882 ( .A1(n9744), .A2(n9737), .ZN(P1_U3302) );
  INV_X1 U10883 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n9738) );
  NOR2_X1 U10884 ( .A1(n9744), .A2(n9738), .ZN(P1_U3303) );
  INV_X1 U10885 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n10117) );
  NOR2_X1 U10886 ( .A1(n9744), .A2(n10117), .ZN(P1_U3304) );
  INV_X1 U10887 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n9739) );
  NOR2_X1 U10888 ( .A1(n9744), .A2(n9739), .ZN(P1_U3305) );
  INV_X1 U10889 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n9740) );
  NOR2_X1 U10890 ( .A1(n9744), .A2(n9740), .ZN(P1_U3306) );
  INV_X1 U10891 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n9741) );
  NOR2_X1 U10892 ( .A1(n9744), .A2(n9741), .ZN(P1_U3307) );
  NOR2_X1 U10893 ( .A1(n9744), .A2(n10092), .ZN(P1_U3308) );
  INV_X1 U10894 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n9742) );
  NOR2_X1 U10895 ( .A1(n9744), .A2(n9742), .ZN(P1_U3309) );
  INV_X1 U10896 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n9743) );
  NOR2_X1 U10897 ( .A1(n9744), .A2(n9743), .ZN(P1_U3310) );
  NOR2_X1 U10898 ( .A1(n9751), .A2(n10040), .ZN(P1_U3311) );
  INV_X1 U10899 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n9745) );
  NOR2_X1 U10900 ( .A1(n9751), .A2(n9745), .ZN(P1_U3312) );
  INV_X1 U10901 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n9746) );
  NOR2_X1 U10902 ( .A1(n9751), .A2(n9746), .ZN(P1_U3313) );
  NOR2_X1 U10903 ( .A1(n9751), .A2(n10196), .ZN(P1_U3314) );
  INV_X1 U10904 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n9747) );
  NOR2_X1 U10905 ( .A1(n9751), .A2(n9747), .ZN(P1_U3315) );
  INV_X1 U10906 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n10103) );
  NOR2_X1 U10907 ( .A1(n9751), .A2(n10103), .ZN(P1_U3316) );
  INV_X1 U10908 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n10183) );
  NOR2_X1 U10909 ( .A1(n9751), .A2(n10183), .ZN(P1_U3317) );
  INV_X1 U10910 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n9748) );
  NOR2_X1 U10911 ( .A1(n9751), .A2(n9748), .ZN(P1_U3318) );
  INV_X1 U10912 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n9749) );
  NOR2_X1 U10913 ( .A1(n9751), .A2(n9749), .ZN(P1_U3319) );
  INV_X1 U10914 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n10026) );
  NOR2_X1 U10915 ( .A1(n9751), .A2(n10026), .ZN(P1_U3320) );
  INV_X1 U10916 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n9750) );
  NOR2_X1 U10917 ( .A1(n9751), .A2(n9750), .ZN(P1_U3321) );
  NAND2_X1 U10918 ( .A1(n9752), .A2(n9755), .ZN(n9753) );
  OAI21_X1 U10919 ( .B1(n9755), .B2(n9754), .A(n9753), .ZN(P1_U3441) );
  OAI21_X1 U10920 ( .B1(n9757), .B2(n9787), .A(n9756), .ZN(n9759) );
  AOI211_X1 U10921 ( .C1(n9793), .C2(n9760), .A(n9759), .B(n9758), .ZN(n9797)
         );
  INV_X1 U10922 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9761) );
  AOI22_X1 U10923 ( .A1(n9795), .A2(n9797), .B1(n9761), .B2(n9794), .ZN(
        P1_U3457) );
  OAI22_X1 U10924 ( .A1(n9763), .A2(n9788), .B1(n9762), .B2(n9787), .ZN(n9765)
         );
  AOI211_X1 U10925 ( .C1(n9793), .C2(n9766), .A(n9765), .B(n9764), .ZN(n9798)
         );
  INV_X1 U10926 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10004) );
  AOI22_X1 U10927 ( .A1(n9795), .A2(n9798), .B1(n10004), .B2(n9794), .ZN(
        P1_U3460) );
  OAI22_X1 U10928 ( .A1(n9768), .A2(n9788), .B1(n9767), .B2(n9787), .ZN(n9770)
         );
  AOI211_X1 U10929 ( .C1(n9793), .C2(n9771), .A(n9770), .B(n9769), .ZN(n9799)
         );
  INV_X1 U10930 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n9772) );
  AOI22_X1 U10931 ( .A1(n9795), .A2(n9799), .B1(n9772), .B2(n9794), .ZN(
        P1_U3466) );
  OAI22_X1 U10932 ( .A1(n9774), .A2(n9788), .B1(n9773), .B2(n9787), .ZN(n9776)
         );
  AOI211_X1 U10933 ( .C1(n9793), .C2(n9777), .A(n9776), .B(n9775), .ZN(n9801)
         );
  INV_X1 U10934 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9778) );
  AOI22_X1 U10935 ( .A1(n9795), .A2(n9801), .B1(n9778), .B2(n9794), .ZN(
        P1_U3472) );
  OAI22_X1 U10936 ( .A1(n9780), .A2(n9788), .B1(n9779), .B2(n9787), .ZN(n9782)
         );
  AOI211_X1 U10937 ( .C1(n9784), .C2(n9783), .A(n9782), .B(n9781), .ZN(n9802)
         );
  INV_X1 U10938 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9785) );
  AOI22_X1 U10939 ( .A1(n9795), .A2(n9802), .B1(n9785), .B2(n9794), .ZN(
        P1_U3478) );
  OAI22_X1 U10940 ( .A1(n9789), .A2(n9788), .B1(n4538), .B2(n9787), .ZN(n9791)
         );
  AOI211_X1 U10941 ( .C1(n9793), .C2(n9792), .A(n9791), .B(n9790), .ZN(n9805)
         );
  INV_X1 U10942 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10072) );
  AOI22_X1 U10943 ( .A1(n9795), .A2(n9805), .B1(n10072), .B2(n9794), .ZN(
        P1_U3481) );
  INV_X1 U10944 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n9796) );
  AOI22_X1 U10945 ( .A1(n9806), .A2(n9797), .B1(n9796), .B2(n9803), .ZN(
        P1_U3524) );
  INV_X1 U10946 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10187) );
  AOI22_X1 U10947 ( .A1(n9806), .A2(n9798), .B1(n10187), .B2(n9803), .ZN(
        P1_U3525) );
  AOI22_X1 U10948 ( .A1(n9806), .A2(n9799), .B1(n6714), .B2(n9803), .ZN(
        P1_U3527) );
  INV_X1 U10949 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n9800) );
  AOI22_X1 U10950 ( .A1(n9806), .A2(n9801), .B1(n9800), .B2(n9803), .ZN(
        P1_U3529) );
  AOI22_X1 U10951 ( .A1(n9806), .A2(n9802), .B1(n6720), .B2(n9803), .ZN(
        P1_U3531) );
  INV_X1 U10952 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n9804) );
  AOI22_X1 U10953 ( .A1(n9806), .A2(n9805), .B1(n9804), .B2(n9803), .ZN(
        P1_U3532) );
  AOI22_X1 U10954 ( .A1(n9808), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n9807), .ZN(n9817) );
  NAND2_X1 U10955 ( .A1(n9808), .A2(n10230), .ZN(n9810) );
  OAI211_X1 U10956 ( .C1(P2_REG1_REG_0__SCAN_IN), .C2(n9811), .A(n9810), .B(
        n9809), .ZN(n9812) );
  INV_X1 U10957 ( .A(n9812), .ZN(n9815) );
  AOI22_X1 U10958 ( .A1(n9813), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n9814) );
  OAI221_X1 U10959 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n9817), .C1(n9816), .C2(
        n9815), .A(n9814), .ZN(P2_U3245) );
  INV_X1 U10960 ( .A(n9819), .ZN(n9831) );
  INV_X1 U10961 ( .A(n9820), .ZN(n9830) );
  INV_X1 U10962 ( .A(n9821), .ZN(n9822) );
  OAI22_X1 U10963 ( .A1(n9825), .A2(n9824), .B1(n9823), .B2(n9822), .ZN(n9826)
         );
  AOI21_X1 U10964 ( .B1(n9828), .B2(n9827), .A(n9826), .ZN(n9829) );
  OAI211_X1 U10965 ( .C1(n9832), .C2(n9831), .A(n9830), .B(n9829), .ZN(n9833)
         );
  INV_X1 U10966 ( .A(n9833), .ZN(n9835) );
  AOI22_X1 U10967 ( .A1(n9836), .A2(n5872), .B1(n9835), .B2(n9834), .ZN(
        P2_U3291) );
  NOR2_X1 U10968 ( .A1(n9838), .A2(n9837), .ZN(n9839) );
  AND2_X1 U10969 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n9843), .ZN(P2_U3297) );
  INV_X1 U10970 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n10123) );
  NOR2_X1 U10971 ( .A1(n9839), .A2(n10123), .ZN(P2_U3298) );
  AND2_X1 U10972 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n9843), .ZN(P2_U3299) );
  AND2_X1 U10973 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n9843), .ZN(P2_U3300) );
  AND2_X1 U10974 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n9843), .ZN(P2_U3301) );
  AND2_X1 U10975 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n9843), .ZN(P2_U3302) );
  AND2_X1 U10976 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n9843), .ZN(P2_U3303) );
  INV_X1 U10977 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n10212) );
  NOR2_X1 U10978 ( .A1(n9839), .A2(n10212), .ZN(P2_U3304) );
  AND2_X1 U10979 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n9843), .ZN(P2_U3305) );
  AND2_X1 U10980 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n9843), .ZN(P2_U3306) );
  AND2_X1 U10981 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n9843), .ZN(P2_U3307) );
  AND2_X1 U10982 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n9843), .ZN(P2_U3308) );
  AND2_X1 U10983 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n9843), .ZN(P2_U3309) );
  AND2_X1 U10984 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n9843), .ZN(P2_U3310) );
  AND2_X1 U10985 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n9843), .ZN(P2_U3311) );
  AND2_X1 U10986 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n9843), .ZN(P2_U3312) );
  AND2_X1 U10987 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n9843), .ZN(P2_U3313) );
  INV_X1 U10988 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n10129) );
  NOR2_X1 U10989 ( .A1(n9839), .A2(n10129), .ZN(P2_U3314) );
  AND2_X1 U10990 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n9843), .ZN(P2_U3315) );
  INV_X1 U10991 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n10028) );
  NOR2_X1 U10992 ( .A1(n9839), .A2(n10028), .ZN(P2_U3316) );
  AND2_X1 U10993 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n9843), .ZN(P2_U3317) );
  AND2_X1 U10994 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n9843), .ZN(P2_U3318) );
  AND2_X1 U10995 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n9843), .ZN(P2_U3319) );
  INV_X1 U10996 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n10213) );
  NOR2_X1 U10997 ( .A1(n9839), .A2(n10213), .ZN(P2_U3320) );
  INV_X1 U10998 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n10045) );
  NOR2_X1 U10999 ( .A1(n9839), .A2(n10045), .ZN(P2_U3321) );
  AND2_X1 U11000 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n9843), .ZN(P2_U3322) );
  AND2_X1 U11001 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n9843), .ZN(P2_U3323) );
  AND2_X1 U11002 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n9843), .ZN(P2_U3324) );
  AND2_X1 U11003 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n9843), .ZN(P2_U3325) );
  AND2_X1 U11004 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n9843), .ZN(P2_U3326) );
  AOI22_X1 U11005 ( .A1(n9840), .A2(n9845), .B1(n10025), .B2(n9843), .ZN(
        P2_U3437) );
  NOR2_X1 U11006 ( .A1(n9842), .A2(n9841), .ZN(n9846) );
  AOI22_X1 U11007 ( .A1(n9846), .A2(n9845), .B1(n9844), .B2(n9843), .ZN(
        P2_U3438) );
  AOI22_X1 U11008 ( .A1(n9849), .A2(n9905), .B1(n9848), .B2(n9847), .ZN(n9850)
         );
  AND2_X1 U11009 ( .A1(n9851), .A2(n9850), .ZN(n9910) );
  AOI22_X1 U11010 ( .A1(n9909), .A2(n9910), .B1(n5838), .B2(n9907), .ZN(
        P2_U3451) );
  NAND3_X1 U11011 ( .A1(n9853), .A2(n9852), .A3(n9883), .ZN(n9854) );
  OAI21_X1 U11012 ( .B1(n6951), .B2(n9899), .A(n9854), .ZN(n9856) );
  AOI211_X1 U11013 ( .C1(n9905), .C2(n9857), .A(n9856), .B(n9855), .ZN(n9911)
         );
  AOI22_X1 U11014 ( .A1(n9909), .A2(n9911), .B1(n5849), .B2(n9907), .ZN(
        P2_U3454) );
  OAI22_X1 U11015 ( .A1(n9859), .A2(n9901), .B1(n9858), .B2(n9899), .ZN(n9862)
         );
  INV_X1 U11016 ( .A(n9860), .ZN(n9861) );
  AOI211_X1 U11017 ( .C1(n9905), .C2(n9863), .A(n9862), .B(n9861), .ZN(n9913)
         );
  AOI22_X1 U11018 ( .A1(n9909), .A2(n9913), .B1(n5827), .B2(n9907), .ZN(
        P2_U3457) );
  OAI22_X1 U11019 ( .A1(n9864), .A2(n9901), .B1(n5870), .B2(n9899), .ZN(n9865)
         );
  AOI21_X1 U11020 ( .B1(n9866), .B2(n9897), .A(n9865), .ZN(n9867) );
  AND2_X1 U11021 ( .A1(n9868), .A2(n9867), .ZN(n9914) );
  AOI22_X1 U11022 ( .A1(n9909), .A2(n9914), .B1(n5863), .B2(n9907), .ZN(
        P2_U3460) );
  OAI22_X1 U11023 ( .A1(n9870), .A2(n9901), .B1(n9869), .B2(n9899), .ZN(n9872)
         );
  AOI211_X1 U11024 ( .C1(n9905), .C2(n9873), .A(n9872), .B(n9871), .ZN(n9915)
         );
  AOI22_X1 U11025 ( .A1(n9909), .A2(n9915), .B1(n5887), .B2(n9907), .ZN(
        P2_U3463) );
  NAND2_X1 U11026 ( .A1(n9874), .A2(n9905), .ZN(n9880) );
  OAI22_X1 U11027 ( .A1(n9876), .A2(n9901), .B1(n9875), .B2(n9899), .ZN(n9877)
         );
  INV_X1 U11028 ( .A(n9877), .ZN(n9878) );
  AND3_X1 U11029 ( .A1(n9880), .A2(n9879), .A3(n9878), .ZN(n9916) );
  AOI22_X1 U11030 ( .A1(n9909), .A2(n9916), .B1(n5903), .B2(n9907), .ZN(
        P2_U3469) );
  AOI22_X1 U11031 ( .A1(n9884), .A2(n9883), .B1(n9882), .B2(n9881), .ZN(n9885)
         );
  OAI21_X1 U11032 ( .B1(n9887), .B2(n9886), .A(n9885), .ZN(n9888) );
  NOR2_X1 U11033 ( .A1(n9889), .A2(n9888), .ZN(n9917) );
  INV_X1 U11034 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10165) );
  AOI22_X1 U11035 ( .A1(n9909), .A2(n9917), .B1(n10165), .B2(n9907), .ZN(
        P2_U3475) );
  INV_X1 U11036 ( .A(n9890), .ZN(n9896) );
  INV_X1 U11037 ( .A(n9891), .ZN(n9892) );
  OAI22_X1 U11038 ( .A1(n9893), .A2(n9901), .B1(n9892), .B2(n9899), .ZN(n9895)
         );
  AOI211_X1 U11039 ( .C1(n9897), .C2(n9896), .A(n9895), .B(n9894), .ZN(n9918)
         );
  INV_X1 U11040 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n9898) );
  AOI22_X1 U11041 ( .A1(n9909), .A2(n9918), .B1(n9898), .B2(n9907), .ZN(
        P2_U3481) );
  OAI22_X1 U11042 ( .A1(n9902), .A2(n9901), .B1(n9900), .B2(n9899), .ZN(n9904)
         );
  AOI211_X1 U11043 ( .C1(n9906), .C2(n9905), .A(n9904), .B(n9903), .ZN(n9919)
         );
  INV_X1 U11044 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n9908) );
  AOI22_X1 U11045 ( .A1(n9909), .A2(n9919), .B1(n9908), .B2(n9907), .ZN(
        P2_U3487) );
  AOI22_X1 U11046 ( .A1(n9996), .A2(n9910), .B1(n5839), .B2(n9994), .ZN(
        P2_U3520) );
  AOI22_X1 U11047 ( .A1(n9996), .A2(n9911), .B1(n6551), .B2(n9994), .ZN(
        P2_U3521) );
  INV_X1 U11048 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n9912) );
  AOI22_X1 U11049 ( .A1(n9996), .A2(n9913), .B1(n9912), .B2(n9994), .ZN(
        P2_U3522) );
  AOI22_X1 U11050 ( .A1(n9996), .A2(n9914), .B1(n5861), .B2(n9994), .ZN(
        P2_U3523) );
  AOI22_X1 U11051 ( .A1(n9996), .A2(n9915), .B1(n5892), .B2(n9994), .ZN(
        P2_U3524) );
  AOI22_X1 U11052 ( .A1(n9996), .A2(n9916), .B1(n6590), .B2(n9994), .ZN(
        P2_U3526) );
  AOI22_X1 U11053 ( .A1(n9996), .A2(n9917), .B1(n5929), .B2(n9994), .ZN(
        P2_U3528) );
  AOI22_X1 U11054 ( .A1(n9996), .A2(n9918), .B1(n6924), .B2(n9994), .ZN(
        P2_U3530) );
  AOI22_X1 U11055 ( .A1(n9996), .A2(n9919), .B1(n7521), .B2(n9994), .ZN(
        P2_U3532) );
  OAI21_X1 U11056 ( .B1(n9922), .B2(n6671), .A(n9920), .ZN(n9921) );
  XNOR2_X1 U11057 ( .A(n9921), .B(P2_ADDR_REG_1__SCAN_IN), .ZN(ADD_1071_U5) );
  OAI21_X1 U11058 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(P2_ADDR_REG_0__SCAN_IN), 
        .A(n9922), .ZN(n9923) );
  INV_X1 U11059 ( .A(n9923), .ZN(ADD_1071_U46) );
  OAI21_X1 U11060 ( .B1(n9926), .B2(n9925), .A(n9924), .ZN(ADD_1071_U56) );
  OAI21_X1 U11061 ( .B1(n9929), .B2(n9928), .A(n9927), .ZN(ADD_1071_U57) );
  OAI21_X1 U11062 ( .B1(n9932), .B2(n9931), .A(n9930), .ZN(ADD_1071_U58) );
  OAI21_X1 U11063 ( .B1(n9935), .B2(n9934), .A(n9933), .ZN(ADD_1071_U59) );
  OAI21_X1 U11064 ( .B1(n9938), .B2(n9937), .A(n9936), .ZN(ADD_1071_U60) );
  OAI21_X1 U11065 ( .B1(n9941), .B2(n9940), .A(n9939), .ZN(ADD_1071_U61) );
  OAI21_X1 U11066 ( .B1(n9944), .B2(n9943), .A(n9942), .ZN(ADD_1071_U62) );
  OAI21_X1 U11067 ( .B1(n9947), .B2(n9946), .A(n9945), .ZN(ADD_1071_U63) );
  NAND4_X1 U11068 ( .A1(P1_D_REG_3__SCAN_IN), .A2(P2_DATAO_REG_29__SCAN_IN), 
        .A3(P2_REG2_REG_18__SCAN_IN), .A4(n10013), .ZN(n9948) );
  NOR3_X1 U11069 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P2_REG2_REG_29__SCAN_IN), 
        .A3(n9948), .ZN(n9958) );
  NOR4_X1 U11070 ( .A1(n9949), .A2(SI_23_), .A3(P1_DATAO_REG_20__SCAN_IN), 
        .A4(P2_REG3_REG_21__SCAN_IN), .ZN(n9950) );
  NAND3_X1 U11071 ( .A1(SI_27_), .A2(n9950), .A3(n10038), .ZN(n9956) );
  NOR4_X1 U11072 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(P1_DATAO_REG_25__SCAN_IN), 
        .A3(n10089), .A4(n10090), .ZN(n9954) );
  NOR4_X1 U11073 ( .A1(P1_REG3_REG_24__SCAN_IN), .A2(P1_REG0_REG_9__SCAN_IN), 
        .A3(n5710), .A4(n10076), .ZN(n9953) );
  NOR4_X1 U11074 ( .A1(P1_REG1_REG_17__SCAN_IN), .A2(P1_DATAO_REG_17__SCAN_IN), 
        .A3(P1_REG2_REG_0__SCAN_IN), .A4(n10117), .ZN(n9952) );
  NOR4_X1 U11075 ( .A1(P1_REG2_REG_29__SCAN_IN), .A2(P1_REG1_REG_8__SCAN_IN), 
        .A3(P2_REG0_REG_27__SCAN_IN), .A4(n10098), .ZN(n9951) );
  NAND4_X1 U11076 ( .A1(n9954), .A2(n9953), .A3(n9952), .A4(n9951), .ZN(n9955)
         );
  NOR4_X1 U11077 ( .A1(P1_REG1_REG_0__SCAN_IN), .A2(P1_U3084), .A3(n9956), 
        .A4(n9955), .ZN(n9957) );
  NAND4_X1 U11078 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P2_REG2_REG_19__SCAN_IN), 
        .A3(n9958), .A4(n9957), .ZN(n9969) );
  INV_X1 U11079 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n10225) );
  NAND4_X1 U11080 ( .A1(n9959), .A2(P1_REG0_REG_19__SCAN_IN), .A3(
        P2_REG2_REG_20__SCAN_IN), .A4(n10225), .ZN(n9968) );
  NAND4_X1 U11081 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_REG2_REG_7__SCAN_IN), 
        .A3(P2_REG1_REG_25__SCAN_IN), .A4(n10119), .ZN(n9960) );
  NOR3_X1 U11082 ( .A1(P1_REG2_REG_19__SCAN_IN), .A2(P1_REG0_REG_0__SCAN_IN), 
        .A3(n9960), .ZN(n9966) );
  NAND4_X1 U11083 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P2_REG3_REG_27__SCAN_IN), 
        .A3(n10187), .A4(n10186), .ZN(n9964) );
  NAND4_X1 U11084 ( .A1(SI_18_), .A2(P1_REG1_REG_24__SCAN_IN), .A3(n6163), 
        .A4(n10157), .ZN(n9963) );
  NAND4_X1 U11085 ( .A1(P1_D_REG_31__SCAN_IN), .A2(P2_REG1_REG_31__SCAN_IN), 
        .A3(P2_REG1_REG_16__SCAN_IN), .A4(n10215), .ZN(n9962) );
  NAND4_X1 U11086 ( .A1(P1_REG0_REG_13__SCAN_IN), .A2(P2_REG3_REG_16__SCAN_IN), 
        .A3(P2_REG1_REG_17__SCAN_IN), .A4(n10200), .ZN(n9961) );
  NOR4_X1 U11087 ( .A1(n9964), .A2(n9963), .A3(n9962), .A4(n9961), .ZN(n9965)
         );
  NAND4_X1 U11088 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P2_REG1_REG_29__SCAN_IN), 
        .A3(n9966), .A4(n9965), .ZN(n9967) );
  NOR4_X1 U11089 ( .A1(P1_REG0_REG_10__SCAN_IN), .A2(n9969), .A3(n9968), .A4(
        n9967), .ZN(n9993) );
  NOR4_X1 U11090 ( .A1(P2_REG2_REG_10__SCAN_IN), .A2(P2_REG0_REG_9__SCAN_IN), 
        .A3(n10223), .A4(n10164), .ZN(n9992) );
  NOR4_X1 U11091 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .A3(P2_ADDR_REG_2__SCAN_IN), .A4(n10194), .ZN(n9975) );
  NAND4_X1 U11092 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_12__SCAN_IN), .A3(
        P2_D_REG_7__SCAN_IN), .A4(n10025), .ZN(n9973) );
  NAND4_X1 U11093 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), 
        .A3(n10015), .A4(n10129), .ZN(n9972) );
  NAND4_X1 U11094 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n10029), .A3(n10082), 
        .A4(n10181), .ZN(n9971) );
  NAND4_X1 U11095 ( .A1(P1_DATAO_REG_11__SCAN_IN), .A2(n10216), .A3(n10150), 
        .A4(n10148), .ZN(n9970) );
  NOR4_X1 U11096 ( .A1(n9973), .A2(n9972), .A3(n9971), .A4(n9970), .ZN(n9974)
         );
  NAND4_X1 U11097 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(n9976), .A3(n9975), .A4(
        n9974), .ZN(n9990) );
  NAND4_X1 U11098 ( .A1(n5778), .A2(SI_7_), .A3(P2_DATAO_REG_0__SCAN_IN), .A4(
        P2_IR_REG_9__SCAN_IN), .ZN(n9980) );
  NOR4_X1 U11099 ( .A1(P2_REG1_REG_7__SCAN_IN), .A2(P2_REG2_REG_8__SCAN_IN), 
        .A3(P2_REG1_REG_8__SCAN_IN), .A4(n10165), .ZN(n9977) );
  INV_X1 U11100 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n10180) );
  NAND3_X1 U11101 ( .A1(n9978), .A2(n9977), .A3(n10180), .ZN(n9979) );
  NOR4_X1 U11102 ( .A1(n9980), .A2(n9979), .A3(P1_DATAO_REG_2__SCAN_IN), .A4(
        P1_DATAO_REG_1__SCAN_IN), .ZN(n9982) );
  NOR2_X1 U11103 ( .A1(n10122), .A2(n10147), .ZN(n9981) );
  NAND4_X1 U11104 ( .A1(n9982), .A2(P2_IR_REG_28__SCAN_IN), .A3(
        P2_IR_REG_2__SCAN_IN), .A4(n9981), .ZN(n9989) );
  NOR4_X1 U11105 ( .A1(P2_REG2_REG_0__SCAN_IN), .A2(P2_REG0_REG_0__SCAN_IN), 
        .A3(n5825), .A4(n10059), .ZN(n9986) );
  NOR4_X1 U11106 ( .A1(P2_REG2_REG_2__SCAN_IN), .A2(P2_REG1_REG_5__SCAN_IN), 
        .A3(n5861), .A4(n5889), .ZN(n9985) );
  NOR4_X1 U11107 ( .A1(P2_DATAO_REG_20__SCAN_IN), .A2(P1_REG0_REG_2__SCAN_IN), 
        .A3(P2_REG0_REG_25__SCAN_IN), .A4(P2_REG2_REG_21__SCAN_IN), .ZN(n9984)
         );
  INV_X1 U11108 ( .A(SI_30_), .ZN(n10000) );
  NOR4_X1 U11109 ( .A1(P1_REG3_REG_1__SCAN_IN), .A2(P2_REG0_REG_23__SCAN_IN), 
        .A3(P2_REG2_REG_15__SCAN_IN), .A4(n10000), .ZN(n9983) );
  NAND4_X1 U11110 ( .A1(n9986), .A2(n9985), .A3(n9984), .A4(n9983), .ZN(n9988)
         );
  NAND4_X1 U11111 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(P2_ADDR_REG_15__SCAN_IN), 
        .A3(P2_ADDR_REG_12__SCAN_IN), .A4(n10060), .ZN(n9987) );
  NOR4_X1 U11112 ( .A1(n9990), .A2(n9989), .A3(n9988), .A4(n9987), .ZN(n9991)
         );
  AND3_X1 U11113 ( .A1(n9993), .A2(n9992), .A3(n9991), .ZN(n10246) );
  AOI22_X1 U11114 ( .A1(n9996), .A2(n9995), .B1(P2_REG1_REG_14__SCAN_IN), .B2(
        n9994), .ZN(n10244) );
  AOI22_X1 U11115 ( .A1(n9998), .A2(keyinput12), .B1(keyinput53), .B2(n5825), 
        .ZN(n9997) );
  OAI221_X1 U11116 ( .B1(n9998), .B2(keyinput12), .C1(n5825), .C2(keyinput53), 
        .A(n9997), .ZN(n10010) );
  AOI22_X1 U11117 ( .A1(n10001), .A2(keyinput98), .B1(n10000), .B2(keyinput8), 
        .ZN(n9999) );
  OAI221_X1 U11118 ( .B1(n10001), .B2(keyinput98), .C1(n10000), .C2(keyinput8), 
        .A(n9999), .ZN(n10009) );
  AOI22_X1 U11119 ( .A1(n10003), .A2(keyinput120), .B1(n5949), .B2(keyinput123), .ZN(n10002) );
  OAI221_X1 U11120 ( .B1(n10003), .B2(keyinput120), .C1(n5949), .C2(
        keyinput123), .A(n10002), .ZN(n10008) );
  XOR2_X1 U11121 ( .A(n10004), .B(keyinput117), .Z(n10006) );
  XNOR2_X1 U11122 ( .A(P1_REG3_REG_1__SCAN_IN), .B(keyinput95), .ZN(n10005) );
  NAND2_X1 U11123 ( .A1(n10006), .A2(n10005), .ZN(n10007) );
  NOR4_X1 U11124 ( .A1(n10010), .A2(n10009), .A3(n10008), .A4(n10007), .ZN(
        n10053) );
  AOI22_X1 U11125 ( .A1(n6078), .A2(keyinput28), .B1(keyinput51), .B2(n5889), 
        .ZN(n10011) );
  OAI221_X1 U11126 ( .B1(n6078), .B2(keyinput28), .C1(n5889), .C2(keyinput51), 
        .A(n10011), .ZN(n10021) );
  AOI22_X1 U11127 ( .A1(n5920), .A2(keyinput96), .B1(n10013), .B2(keyinput55), 
        .ZN(n10012) );
  OAI221_X1 U11128 ( .B1(n5920), .B2(keyinput96), .C1(n10013), .C2(keyinput55), 
        .A(n10012), .ZN(n10020) );
  AOI22_X1 U11129 ( .A1(n5938), .A2(keyinput110), .B1(keyinput21), .B2(n10015), 
        .ZN(n10014) );
  OAI221_X1 U11130 ( .B1(n5938), .B2(keyinput110), .C1(n10015), .C2(keyinput21), .A(n10014), .ZN(n10019) );
  XOR2_X1 U11131 ( .A(n6175), .B(keyinput45), .Z(n10017) );
  XNOR2_X1 U11132 ( .A(P1_IR_REG_12__SCAN_IN), .B(keyinput13), .ZN(n10016) );
  NAND2_X1 U11133 ( .A1(n10017), .A2(n10016), .ZN(n10018) );
  NOR4_X1 U11134 ( .A1(n10021), .A2(n10020), .A3(n10019), .A4(n10018), .ZN(
        n10052) );
  AOI22_X1 U11135 ( .A1(n7617), .A2(keyinput74), .B1(n10023), .B2(keyinput67), 
        .ZN(n10022) );
  OAI221_X1 U11136 ( .B1(n7617), .B2(keyinput74), .C1(n10023), .C2(keyinput67), 
        .A(n10022), .ZN(n10036) );
  AOI22_X1 U11137 ( .A1(n10026), .A2(keyinput54), .B1(keyinput81), .B2(n10025), 
        .ZN(n10024) );
  OAI221_X1 U11138 ( .B1(n10026), .B2(keyinput54), .C1(n10025), .C2(keyinput81), .A(n10024), .ZN(n10035) );
  AOI22_X1 U11139 ( .A1(n10029), .A2(keyinput2), .B1(keyinput61), .B2(n10028), 
        .ZN(n10027) );
  OAI221_X1 U11140 ( .B1(n10029), .B2(keyinput2), .C1(n10028), .C2(keyinput61), 
        .A(n10027), .ZN(n10034) );
  INV_X1 U11141 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n10031) );
  AOI22_X1 U11142 ( .A1(n10032), .A2(keyinput10), .B1(n10031), .B2(keyinput77), 
        .ZN(n10030) );
  OAI221_X1 U11143 ( .B1(n10032), .B2(keyinput10), .C1(n10031), .C2(keyinput77), .A(n10030), .ZN(n10033) );
  NOR4_X1 U11144 ( .A1(n10036), .A2(n10035), .A3(n10034), .A4(n10033), .ZN(
        n10051) );
  AOI22_X1 U11145 ( .A1(n10038), .A2(keyinput25), .B1(keyinput18), .B2(n5826), 
        .ZN(n10037) );
  OAI221_X1 U11146 ( .B1(n10038), .B2(keyinput25), .C1(n5826), .C2(keyinput18), 
        .A(n10037), .ZN(n10049) );
  AOI22_X1 U11147 ( .A1(n10041), .A2(keyinput79), .B1(n10040), .B2(keyinput78), 
        .ZN(n10039) );
  OAI221_X1 U11148 ( .B1(n10041), .B2(keyinput79), .C1(n10040), .C2(keyinput78), .A(n10039), .ZN(n10048) );
  XOR2_X1 U11149 ( .A(n6057), .B(keyinput92), .Z(n10044) );
  XNOR2_X1 U11150 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(keyinput97), .ZN(n10043)
         );
  XNOR2_X1 U11151 ( .A(P1_IR_REG_9__SCAN_IN), .B(keyinput127), .ZN(n10042) );
  NAND3_X1 U11152 ( .A1(n10044), .A2(n10043), .A3(n10042), .ZN(n10047) );
  XNOR2_X1 U11153 ( .A(n10045), .B(keyinput100), .ZN(n10046) );
  NOR4_X1 U11154 ( .A1(n10049), .A2(n10048), .A3(n10047), .A4(n10046), .ZN(
        n10050) );
  NAND4_X1 U11155 ( .A1(n10053), .A2(n10052), .A3(n10051), .A4(n10050), .ZN(
        n10242) );
  AOI22_X1 U11156 ( .A1(n10055), .A2(keyinput50), .B1(P1_U3084), .B2(
        keyinput39), .ZN(n10054) );
  OAI221_X1 U11157 ( .B1(n10055), .B2(keyinput50), .C1(P1_U3084), .C2(
        keyinput39), .A(n10054), .ZN(n10067) );
  AOI22_X1 U11158 ( .A1(n4670), .A2(keyinput58), .B1(keyinput91), .B2(n10057), 
        .ZN(n10056) );
  OAI221_X1 U11159 ( .B1(n4670), .B2(keyinput58), .C1(n10057), .C2(keyinput91), 
        .A(n10056), .ZN(n10066) );
  AOI22_X1 U11160 ( .A1(n10060), .A2(keyinput94), .B1(n10059), .B2(keyinput27), 
        .ZN(n10058) );
  OAI221_X1 U11161 ( .B1(n10060), .B2(keyinput94), .C1(n10059), .C2(keyinput27), .A(n10058), .ZN(n10065) );
  AOI22_X1 U11162 ( .A1(n10063), .A2(keyinput63), .B1(keyinput35), .B2(n10062), 
        .ZN(n10061) );
  OAI221_X1 U11163 ( .B1(n10063), .B2(keyinput63), .C1(n10062), .C2(keyinput35), .A(n10061), .ZN(n10064) );
  NOR4_X1 U11164 ( .A1(n10067), .A2(n10066), .A3(n10065), .A4(n10064), .ZN(
        n10111) );
  AOI22_X1 U11165 ( .A1(n10069), .A2(keyinput70), .B1(keyinput115), .B2(n6560), 
        .ZN(n10068) );
  OAI221_X1 U11166 ( .B1(n10069), .B2(keyinput70), .C1(n6560), .C2(keyinput115), .A(n10068), .ZN(n10080) );
  AOI22_X1 U11167 ( .A1(n6406), .A2(keyinput34), .B1(n5710), .B2(keyinput0), 
        .ZN(n10070) );
  OAI221_X1 U11168 ( .B1(n6406), .B2(keyinput34), .C1(n5710), .C2(keyinput0), 
        .A(n10070), .ZN(n10079) );
  AOI22_X1 U11169 ( .A1(n10073), .A2(keyinput11), .B1(keyinput49), .B2(n10072), 
        .ZN(n10071) );
  OAI221_X1 U11170 ( .B1(n10073), .B2(keyinput11), .C1(n10072), .C2(keyinput49), .A(n10071), .ZN(n10078) );
  AOI22_X1 U11171 ( .A1(n10076), .A2(keyinput44), .B1(n10075), .B2(keyinput116), .ZN(n10074) );
  OAI221_X1 U11172 ( .B1(n10076), .B2(keyinput44), .C1(n10075), .C2(
        keyinput116), .A(n10074), .ZN(n10077) );
  NOR4_X1 U11173 ( .A1(n10080), .A2(n10079), .A3(n10078), .A4(n10077), .ZN(
        n10110) );
  AOI22_X1 U11174 ( .A1(n6720), .A2(keyinput111), .B1(n10082), .B2(keyinput105), .ZN(n10081) );
  OAI221_X1 U11175 ( .B1(n6720), .B2(keyinput111), .C1(n10082), .C2(
        keyinput105), .A(n10081), .ZN(n10087) );
  XNOR2_X1 U11176 ( .A(n10083), .B(keyinput30), .ZN(n10086) );
  XNOR2_X1 U11177 ( .A(n10084), .B(keyinput103), .ZN(n10085) );
  OR3_X1 U11178 ( .A1(n10087), .A2(n10086), .A3(n10085), .ZN(n10095) );
  AOI22_X1 U11179 ( .A1(n10090), .A2(keyinput84), .B1(n10089), .B2(keyinput41), 
        .ZN(n10088) );
  OAI221_X1 U11180 ( .B1(n10090), .B2(keyinput84), .C1(n10089), .C2(keyinput41), .A(n10088), .ZN(n10094) );
  AOI22_X1 U11181 ( .A1(n10092), .A2(keyinput122), .B1(keyinput52), .B2(n6822), 
        .ZN(n10091) );
  OAI221_X1 U11182 ( .B1(n10092), .B2(keyinput122), .C1(n6822), .C2(keyinput52), .A(n10091), .ZN(n10093) );
  NOR3_X1 U11183 ( .A1(n10095), .A2(n10094), .A3(n10093), .ZN(n10109) );
  AOI22_X1 U11184 ( .A1(n10098), .A2(keyinput9), .B1(keyinput101), .B2(n10097), 
        .ZN(n10096) );
  OAI221_X1 U11185 ( .B1(n10098), .B2(keyinput9), .C1(n10097), .C2(keyinput101), .A(n10096), .ZN(n10107) );
  INV_X1 U11186 ( .A(SI_7_), .ZN(n10100) );
  AOI22_X1 U11187 ( .A1(n10100), .A2(keyinput75), .B1(keyinput99), .B2(n5929), 
        .ZN(n10099) );
  OAI221_X1 U11188 ( .B1(n10100), .B2(keyinput75), .C1(n5929), .C2(keyinput99), 
        .A(n10099), .ZN(n10106) );
  AOI22_X1 U11189 ( .A1(n9162), .A2(keyinput16), .B1(keyinput56), .B2(n5838), 
        .ZN(n10101) );
  OAI221_X1 U11190 ( .B1(n9162), .B2(keyinput16), .C1(n5838), .C2(keyinput56), 
        .A(n10101), .ZN(n10105) );
  AOI22_X1 U11191 ( .A1(n10103), .A2(keyinput76), .B1(keyinput57), .B2(n7851), 
        .ZN(n10102) );
  OAI221_X1 U11192 ( .B1(n10103), .B2(keyinput76), .C1(n7851), .C2(keyinput57), 
        .A(n10102), .ZN(n10104) );
  NOR4_X1 U11193 ( .A1(n10107), .A2(n10106), .A3(n10105), .A4(n10104), .ZN(
        n10108) );
  NAND4_X1 U11194 ( .A1(n10111), .A2(n10110), .A3(n10109), .A4(n10108), .ZN(
        n10241) );
  AOI22_X1 U11195 ( .A1(n10114), .A2(keyinput69), .B1(n10113), .B2(keyinput114), .ZN(n10112) );
  OAI221_X1 U11196 ( .B1(n10114), .B2(keyinput69), .C1(n10113), .C2(
        keyinput114), .A(n10112), .ZN(n10127) );
  INV_X1 U11197 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n10116) );
  AOI22_X1 U11198 ( .A1(n10117), .A2(keyinput68), .B1(keyinput32), .B2(n10116), 
        .ZN(n10115) );
  OAI221_X1 U11199 ( .B1(n10117), .B2(keyinput68), .C1(n10116), .C2(keyinput32), .A(n10115), .ZN(n10126) );
  AOI22_X1 U11200 ( .A1(n10120), .A2(keyinput15), .B1(n10119), .B2(keyinput4), 
        .ZN(n10118) );
  OAI221_X1 U11201 ( .B1(n10120), .B2(keyinput15), .C1(n10119), .C2(keyinput4), 
        .A(n10118), .ZN(n10125) );
  AOI22_X1 U11202 ( .A1(n10123), .A2(keyinput48), .B1(n10122), .B2(keyinput125), .ZN(n10121) );
  OAI221_X1 U11203 ( .B1(n10123), .B2(keyinput48), .C1(n10122), .C2(
        keyinput125), .A(n10121), .ZN(n10124) );
  NOR4_X1 U11204 ( .A1(n10127), .A2(n10126), .A3(n10125), .A4(n10124), .ZN(
        n10175) );
  INV_X1 U11205 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n10130) );
  AOI22_X1 U11206 ( .A1(n10130), .A2(keyinput5), .B1(keyinput7), .B2(n10129), 
        .ZN(n10128) );
  OAI221_X1 U11207 ( .B1(n10130), .B2(keyinput5), .C1(n10129), .C2(keyinput7), 
        .A(n10128), .ZN(n10141) );
  AOI22_X1 U11208 ( .A1(n10133), .A2(keyinput23), .B1(n10132), .B2(keyinput108), .ZN(n10131) );
  OAI221_X1 U11209 ( .B1(n10133), .B2(keyinput23), .C1(n10132), .C2(
        keyinput108), .A(n10131), .ZN(n10140) );
  XNOR2_X1 U11210 ( .A(P2_IR_REG_28__SCAN_IN), .B(keyinput38), .ZN(n10136) );
  XNOR2_X1 U11211 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(keyinput17), .ZN(n10135)
         );
  XNOR2_X1 U11212 ( .A(keyinput86), .B(P2_REG1_REG_3__SCAN_IN), .ZN(n10134) );
  NAND3_X1 U11213 ( .A1(n10136), .A2(n10135), .A3(n10134), .ZN(n10139) );
  XNOR2_X1 U11214 ( .A(n10137), .B(keyinput62), .ZN(n10138) );
  NOR4_X1 U11215 ( .A1(n10141), .A2(n10140), .A3(n10139), .A4(n10138), .ZN(
        n10174) );
  AOI22_X1 U11216 ( .A1(n7290), .A2(keyinput126), .B1(n10143), .B2(keyinput40), 
        .ZN(n10142) );
  OAI221_X1 U11217 ( .B1(n7290), .B2(keyinput126), .C1(n10143), .C2(keyinput40), .A(n10142), .ZN(n10155) );
  INV_X1 U11218 ( .A(SI_18_), .ZN(n10145) );
  AOI22_X1 U11219 ( .A1(n10145), .A2(keyinput80), .B1(keyinput19), .B2(n6163), 
        .ZN(n10144) );
  OAI221_X1 U11220 ( .B1(n10145), .B2(keyinput80), .C1(n6163), .C2(keyinput19), 
        .A(n10144), .ZN(n10154) );
  AOI22_X1 U11221 ( .A1(n10148), .A2(keyinput46), .B1(keyinput1), .B2(n10147), 
        .ZN(n10146) );
  OAI221_X1 U11222 ( .B1(n10148), .B2(keyinput46), .C1(n10147), .C2(keyinput1), 
        .A(n10146), .ZN(n10153) );
  AOI22_X1 U11223 ( .A1(n10151), .A2(keyinput106), .B1(n10150), .B2(
        keyinput104), .ZN(n10149) );
  OAI221_X1 U11224 ( .B1(n10151), .B2(keyinput106), .C1(n10150), .C2(
        keyinput104), .A(n10149), .ZN(n10152) );
  NOR4_X1 U11225 ( .A1(n10155), .A2(n10154), .A3(n10153), .A4(n10152), .ZN(
        n10173) );
  AOI22_X1 U11226 ( .A1(n10158), .A2(keyinput66), .B1(keyinput121), .B2(n10157), .ZN(n10156) );
  OAI221_X1 U11227 ( .B1(n10158), .B2(keyinput66), .C1(n10157), .C2(
        keyinput121), .A(n10156), .ZN(n10171) );
  AOI22_X1 U11228 ( .A1(n10161), .A2(keyinput6), .B1(keyinput37), .B2(n10160), 
        .ZN(n10159) );
  OAI221_X1 U11229 ( .B1(n10161), .B2(keyinput6), .C1(n10160), .C2(keyinput37), 
        .A(n10159), .ZN(n10170) );
  INV_X1 U11230 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n10163) );
  AOI22_X1 U11231 ( .A1(n10164), .A2(keyinput42), .B1(keyinput64), .B2(n10163), 
        .ZN(n10162) );
  OAI221_X1 U11232 ( .B1(n10164), .B2(keyinput42), .C1(n10163), .C2(keyinput64), .A(n10162), .ZN(n10169) );
  XOR2_X1 U11233 ( .A(n10165), .B(keyinput31), .Z(n10167) );
  XNOR2_X1 U11234 ( .A(P2_IR_REG_4__SCAN_IN), .B(keyinput73), .ZN(n10166) );
  NAND2_X1 U11235 ( .A1(n10167), .A2(n10166), .ZN(n10168) );
  NOR4_X1 U11236 ( .A1(n10171), .A2(n10170), .A3(n10169), .A4(n10168), .ZN(
        n10172) );
  NAND4_X1 U11237 ( .A1(n10175), .A2(n10174), .A3(n10173), .A4(n10172), .ZN(
        n10240) );
  AOI22_X1 U11238 ( .A1(n10178), .A2(keyinput119), .B1(keyinput22), .B2(n10177), .ZN(n10176) );
  OAI221_X1 U11239 ( .B1(n10178), .B2(keyinput119), .C1(n10177), .C2(
        keyinput22), .A(n10176), .ZN(n10191) );
  AOI22_X1 U11240 ( .A1(n10181), .A2(keyinput124), .B1(keyinput26), .B2(n10180), .ZN(n10179) );
  OAI221_X1 U11241 ( .B1(n10181), .B2(keyinput124), .C1(n10180), .C2(
        keyinput26), .A(n10179), .ZN(n10190) );
  INV_X1 U11242 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n10184) );
  AOI22_X1 U11243 ( .A1(n10184), .A2(keyinput113), .B1(n10183), .B2(
        keyinput118), .ZN(n10182) );
  OAI221_X1 U11244 ( .B1(n10184), .B2(keyinput113), .C1(n10183), .C2(
        keyinput118), .A(n10182), .ZN(n10189) );
  AOI22_X1 U11245 ( .A1(n10187), .A2(keyinput65), .B1(n10186), .B2(keyinput24), 
        .ZN(n10185) );
  OAI221_X1 U11246 ( .B1(n10187), .B2(keyinput65), .C1(n10186), .C2(keyinput24), .A(n10185), .ZN(n10188) );
  NOR4_X1 U11247 ( .A1(n10191), .A2(n10190), .A3(n10189), .A4(n10188), .ZN(
        n10238) );
  AOI22_X1 U11248 ( .A1(n10194), .A2(keyinput109), .B1(n10193), .B2(keyinput88), .ZN(n10192) );
  OAI221_X1 U11249 ( .B1(n10194), .B2(keyinput109), .C1(n10193), .C2(
        keyinput88), .A(n10192), .ZN(n10206) );
  AOI22_X1 U11250 ( .A1(n10197), .A2(keyinput102), .B1(n10196), .B2(keyinput93), .ZN(n10195) );
  OAI221_X1 U11251 ( .B1(n10197), .B2(keyinput102), .C1(n10196), .C2(
        keyinput93), .A(n10195), .ZN(n10205) );
  AOI22_X1 U11252 ( .A1(n10200), .A2(keyinput33), .B1(n10199), .B2(keyinput90), 
        .ZN(n10198) );
  OAI221_X1 U11253 ( .B1(n10200), .B2(keyinput33), .C1(n10199), .C2(keyinput90), .A(n10198), .ZN(n10204) );
  XNOR2_X1 U11254 ( .A(P2_REG1_REG_17__SCAN_IN), .B(keyinput85), .ZN(n10202)
         );
  XNOR2_X1 U11255 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(keyinput72), .ZN(n10201)
         );
  NAND2_X1 U11256 ( .A1(n10202), .A2(n10201), .ZN(n10203) );
  NOR4_X1 U11257 ( .A1(n10206), .A2(n10205), .A3(n10204), .A4(n10203), .ZN(
        n10237) );
  AOI22_X1 U11258 ( .A1(n4970), .A2(keyinput47), .B1(keyinput83), .B2(n10208), 
        .ZN(n10207) );
  OAI221_X1 U11259 ( .B1(n4970), .B2(keyinput47), .C1(n10208), .C2(keyinput83), 
        .A(n10207), .ZN(n10220) );
  AOI22_X1 U11260 ( .A1(n10210), .A2(keyinput29), .B1(n6046), .B2(keyinput43), 
        .ZN(n10209) );
  OAI221_X1 U11261 ( .B1(n10210), .B2(keyinput29), .C1(n6046), .C2(keyinput43), 
        .A(n10209), .ZN(n10219) );
  AOI22_X1 U11262 ( .A1(n10213), .A2(keyinput112), .B1(n10212), .B2(
        keyinput107), .ZN(n10211) );
  OAI221_X1 U11263 ( .B1(n10213), .B2(keyinput112), .C1(n10212), .C2(
        keyinput107), .A(n10211), .ZN(n10218) );
  AOI22_X1 U11264 ( .A1(n10216), .A2(keyinput60), .B1(keyinput82), .B2(n10215), 
        .ZN(n10214) );
  OAI221_X1 U11265 ( .B1(n10216), .B2(keyinput60), .C1(n10215), .C2(keyinput82), .A(n10214), .ZN(n10217) );
  NOR4_X1 U11266 ( .A1(n10220), .A2(n10219), .A3(n10218), .A4(n10217), .ZN(
        n10236) );
  AOI22_X1 U11267 ( .A1(n10223), .A2(keyinput89), .B1(n10222), .B2(keyinput14), 
        .ZN(n10221) );
  OAI221_X1 U11268 ( .B1(n10223), .B2(keyinput89), .C1(n10222), .C2(keyinput14), .A(n10221), .ZN(n10234) );
  AOI22_X1 U11269 ( .A1(n10226), .A2(keyinput71), .B1(n10225), .B2(keyinput36), 
        .ZN(n10224) );
  OAI221_X1 U11270 ( .B1(n10226), .B2(keyinput71), .C1(n10225), .C2(keyinput36), .A(n10224), .ZN(n10233) );
  AOI22_X1 U11271 ( .A1(n10228), .A2(keyinput3), .B1(keyinput87), .B2(n6068), 
        .ZN(n10227) );
  OAI221_X1 U11272 ( .B1(n10228), .B2(keyinput3), .C1(n6068), .C2(keyinput87), 
        .A(n10227), .ZN(n10232) );
  AOI22_X1 U11273 ( .A1(n10230), .A2(keyinput20), .B1(n5421), .B2(keyinput59), 
        .ZN(n10229) );
  OAI221_X1 U11274 ( .B1(n10230), .B2(keyinput20), .C1(n5421), .C2(keyinput59), 
        .A(n10229), .ZN(n10231) );
  NOR4_X1 U11275 ( .A1(n10234), .A2(n10233), .A3(n10232), .A4(n10231), .ZN(
        n10235) );
  NAND4_X1 U11276 ( .A1(n10238), .A2(n10237), .A3(n10236), .A4(n10235), .ZN(
        n10239) );
  NOR4_X1 U11277 ( .A1(n10242), .A2(n10241), .A3(n10240), .A4(n10239), .ZN(
        n10243) );
  XOR2_X1 U11278 ( .A(n10244), .B(n10243), .Z(n10245) );
  XNOR2_X1 U11279 ( .A(n10246), .B(n10245), .ZN(P2_U3534) );
  OAI21_X1 U11280 ( .B1(n10249), .B2(n10248), .A(n10247), .ZN(ADD_1071_U48) );
  OAI21_X1 U11281 ( .B1(n10252), .B2(n10251), .A(n10250), .ZN(ADD_1071_U50) );
  OAI21_X1 U11282 ( .B1(n10255), .B2(n10254), .A(n10253), .ZN(ADD_1071_U51) );
  OAI21_X1 U11283 ( .B1(n10258), .B2(n10257), .A(n10256), .ZN(ADD_1071_U49) );
  OAI21_X1 U11284 ( .B1(n10261), .B2(n10260), .A(n10259), .ZN(ADD_1071_U55) );
  OAI21_X1 U11285 ( .B1(n10264), .B2(n10263), .A(n10262), .ZN(ADD_1071_U47) );
  AOI21_X1 U11286 ( .B1(n10267), .B2(n10266), .A(n10265), .ZN(ADD_1071_U54) );
  AOI21_X1 U11287 ( .B1(n10270), .B2(n10269), .A(n10268), .ZN(ADD_1071_U53) );
  OAI21_X1 U11288 ( .B1(n10273), .B2(n10272), .A(n10271), .ZN(ADD_1071_U52) );
  CLKBUF_X1 U4902 ( .A(n6050), .Z(n6206) );
  NOR2_X1 U4903 ( .A1(n4955), .A2(n4939), .ZN(n4940) );
  CLKBUF_X1 U4905 ( .A(n5037), .Z(n5758) );
  NAND2_X1 U4906 ( .A1(n5607), .A2(n5606), .ZN(n5629) );
  CLKBUF_X1 U5032 ( .A(n7655), .Z(n7656) );
  INV_X1 U5598 ( .A(n4973), .ZN(n5239) );
endmodule

