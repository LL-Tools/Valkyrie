

module b15_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, U3445, U3446, U3447, U3448, 
        U3213, U3212, U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, 
        U3203, U3202, U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, 
        U3193, U3192, U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, 
        U3183, U3182, U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, 
        U3175, U3174, U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, 
        U3165, U3164, U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, 
        U3155, U3154, U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, 
        U3146, U3145, U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, 
        U3136, U3135, U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, 
        U3126, U3125, U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, 
        U3116, U3115, U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, 
        U3106, U3105, U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, 
        U3096, U3095, U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, 
        U3086, U3085, U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, 
        U3076, U3075, U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, 
        U3066, U3065, U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, 
        U3056, U3055, U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, 
        U3046, U3045, U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, 
        U3036, U3035, U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, 
        U3026, U3025, U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, 
        U3460, U3461, U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, 
        U3015, U3014, U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, 
        U3005, U3004, U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, 
        U2995, U2994, U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, 
        U2985, U2984, U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, 
        U2975, U2974, U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, 
        U2965, U2964, U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, 
        U2955, U2954, U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, 
        U2945, U2944, U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, 
        U2935, U2934, U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, 
        U2925, U2924, U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, 
        U2915, U2914, U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, 
        U2905, U2904, U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, 
        U2895, U2894, U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, 
        U2885, U2884, U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, 
        U2875, U2874, U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, 
        U2865, U2864, U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, 
        U2855, U2854, U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, 
        U2845, U2844, U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, 
        U2835, U2834, U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, 
        U2825, U2824, U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, 
        U2815, U2814, U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, 
        U2805, U2804, U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, 
        U2795, U3468, U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, 
        U3473, U2790, U2789, U3474, U2788, keyinput0, keyinput1, keyinput2, 
        keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, 
        keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, 
        keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, 
        keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, 
        keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, 
        keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, 
        keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, 
        keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, 
        keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, 
        keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, 
        keyinput63 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1,
         keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7,
         keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13,
         keyinput14, keyinput15, keyinput16, keyinput17, keyinput18,
         keyinput19, keyinput20, keyinput21, keyinput22, keyinput23,
         keyinput24, keyinput25, keyinput26, keyinput27, keyinput28,
         keyinput29, keyinput30, keyinput31, keyinput32, keyinput33,
         keyinput34, keyinput35, keyinput36, keyinput37, keyinput38,
         keyinput39, keyinput40, keyinput41, keyinput42, keyinput43,
         keyinput44, keyinput45, keyinput46, keyinput47, keyinput48,
         keyinput49, keyinput50, keyinput51, keyinput52, keyinput53,
         keyinput54, keyinput55, keyinput56, keyinput57, keyinput58,
         keyinput59, keyinput60, keyinput61, keyinput62, keyinput63;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975,
         n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985,
         n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995,
         n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005,
         n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015,
         n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025,
         n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035,
         n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045,
         n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055,
         n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065,
         n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075,
         n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085,
         n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095,
         n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105,
         n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115,
         n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125,
         n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135,
         n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145,
         n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155,
         n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165,
         n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175,
         n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185,
         n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195,
         n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205,
         n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215,
         n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225,
         n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235,
         n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245,
         n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255,
         n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265,
         n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275,
         n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285,
         n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295,
         n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305,
         n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315,
         n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325,
         n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335,
         n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345,
         n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355,
         n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365,
         n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375,
         n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385,
         n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395,
         n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405,
         n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415,
         n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425,
         n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435,
         n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445,
         n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455,
         n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465,
         n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475,
         n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485,
         n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495,
         n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505,
         n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515,
         n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525,
         n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535,
         n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545,
         n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555,
         n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565,
         n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575,
         n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585,
         n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595,
         n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605,
         n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615,
         n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625,
         n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635,
         n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645,
         n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655,
         n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665,
         n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675,
         n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685,
         n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695,
         n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705,
         n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715,
         n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725,
         n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735,
         n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745,
         n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755,
         n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765,
         n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775,
         n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785,
         n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795,
         n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805,
         n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815,
         n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825,
         n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835,
         n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845,
         n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855,
         n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865,
         n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875,
         n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885,
         n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895,
         n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905,
         n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915,
         n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925,
         n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935,
         n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945,
         n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955,
         n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965,
         n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975,
         n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985,
         n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995,
         n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005,
         n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015,
         n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025,
         n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035,
         n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045,
         n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055,
         n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065,
         n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075,
         n4076, n4077, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086,
         n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096,
         n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106,
         n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116,
         n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126,
         n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136,
         n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146,
         n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156,
         n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166,
         n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176,
         n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186,
         n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196,
         n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206,
         n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216,
         n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226,
         n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236,
         n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246,
         n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256,
         n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266,
         n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276,
         n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286,
         n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296,
         n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306,
         n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316,
         n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326,
         n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336,
         n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346,
         n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356,
         n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366,
         n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376,
         n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386,
         n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396,
         n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406,
         n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416,
         n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426,
         n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436,
         n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446,
         n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456,
         n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466,
         n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476,
         n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486,
         n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496,
         n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506,
         n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516,
         n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526,
         n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536,
         n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546,
         n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556,
         n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
         n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576,
         n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586,
         n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596,
         n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606,
         n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616,
         n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626,
         n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636,
         n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646,
         n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656,
         n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666,
         n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676,
         n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686,
         n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696,
         n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706,
         n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716,
         n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726,
         n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736,
         n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746,
         n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756,
         n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766,
         n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776,
         n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786,
         n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796,
         n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806,
         n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816,
         n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826,
         n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836,
         n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846,
         n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856,
         n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866,
         n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876,
         n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886,
         n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896,
         n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906,
         n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916,
         n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926,
         n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936,
         n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946,
         n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956,
         n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966,
         n4967, n4968, n4969, n4971, n4972, n4973, n4974, n4975, n4976, n4977,
         n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987,
         n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997,
         n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007,
         n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017,
         n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027,
         n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037,
         n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047,
         n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057,
         n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067,
         n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077,
         n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087,
         n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097,
         n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107,
         n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117,
         n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127,
         n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137,
         n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147,
         n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157,
         n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167,
         n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177,
         n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187,
         n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197,
         n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207,
         n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217,
         n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227,
         n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237,
         n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247,
         n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257,
         n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267,
         n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277,
         n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287,
         n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297,
         n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307,
         n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317,
         n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327,
         n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337,
         n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347,
         n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357,
         n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367,
         n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377,
         n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387,
         n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397,
         n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407,
         n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417,
         n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427,
         n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437,
         n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447,
         n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457,
         n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467,
         n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477,
         n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487,
         n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497,
         n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5506, n5507, n5508,
         n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518,
         n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528,
         n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538,
         n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548,
         n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558,
         n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568,
         n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578,
         n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588,
         n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598,
         n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608,
         n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618,
         n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628,
         n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638,
         n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648,
         n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658,
         n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668,
         n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678,
         n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688,
         n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698,
         n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708,
         n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718,
         n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728,
         n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738,
         n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748,
         n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758,
         n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768,
         n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778,
         n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788,
         n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798,
         n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808,
         n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818,
         n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828,
         n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838,
         n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848,
         n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858,
         n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868,
         n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878,
         n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888,
         n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898,
         n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908,
         n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918,
         n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928,
         n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938,
         n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948,
         n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958,
         n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968,
         n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978,
         n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988,
         n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998,
         n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008,
         n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018,
         n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028,
         n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038,
         n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048,
         n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058,
         n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068,
         n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078,
         n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088,
         n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098,
         n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108,
         n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118,
         n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128,
         n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138,
         n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148,
         n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158,
         n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168,
         n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178,
         n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188,
         n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198,
         n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208,
         n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218,
         n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228,
         n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238,
         n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248,
         n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258,
         n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268,
         n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278,
         n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288,
         n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298,
         n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308,
         n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318,
         n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328,
         n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338,
         n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348,
         n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358,
         n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368,
         n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378,
         n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388,
         n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398,
         n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408,
         n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418,
         n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428,
         n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438,
         n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448,
         n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458,
         n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468,
         n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478,
         n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488,
         n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498,
         n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508,
         n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518,
         n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528,
         n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538,
         n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548,
         n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558,
         n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568,
         n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578,
         n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588,
         n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598,
         n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608,
         n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618,
         n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628,
         n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638,
         n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648,
         n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658,
         n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668,
         n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678,
         n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688,
         n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698,
         n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708,
         n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718,
         n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728,
         n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738,
         n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748,
         n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758,
         n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768,
         n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778,
         n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788,
         n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798,
         n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808,
         n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818,
         n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828,
         n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838,
         n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848,
         n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856;

  XNOR2_X1 U3414 ( .A(n3384), .B(n3383), .ZN(n3565) );
  CLKBUF_X2 U3415 ( .A(n3608), .Z(n4005) );
  CLKBUF_X2 U3416 ( .A(n3295), .Z(n3953) );
  CLKBUF_X2 U3417 ( .A(n3959), .Z(n3994) );
  INV_X1 U3418 ( .A(n3829), .ZN(n3980) );
  AND4_X2 U3419 ( .A1(n3245), .A2(n2987), .A3(n3244), .A4(n3243), .ZN(n4692)
         );
  AND4_X1 U3420 ( .A1(n3281), .A2(n3280), .A3(n3279), .A4(n3278), .ZN(n3282)
         );
  AND2_X2 U3421 ( .A1(n4542), .A2(n4517), .ZN(n3418) );
  CLKBUF_X1 U3422 ( .A(n6657), .Z(n2966) );
  NOR2_X1 U3423 ( .A1(n6610), .A2(n6678), .ZN(n6657) );
  CLKBUF_X3 U3425 ( .A(n3277), .Z(n3917) );
  AND2_X2 U3426 ( .A1(n4545), .A2(n4540), .ZN(n3827) );
  NAND2_X1 U3427 ( .A1(n4692), .A2(n4105), .ZN(n4340) );
  NAND2_X1 U3428 ( .A1(n3401), .A2(n3400), .ZN(n3541) );
  CLKBUF_X3 U3430 ( .A(n3262), .Z(n4099) );
  OR2_X1 U3431 ( .A1(n5755), .A2(n3075), .ZN(n3070) );
  NAND3_X1 U3432 ( .A1(n3565), .A2(n3568), .A3(n3439), .ZN(n3571) );
  BUF_X1 U3433 ( .A(n4263), .Z(n4326) );
  XOR2_X1 U3435 ( .A(n5233), .B(n5349), .Z(n5322) );
  XNOR2_X1 U3436 ( .A(n3045), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4391)
         );
  CLKBUF_X3 U3437 ( .A(n4685), .Z(n2976) );
  INV_X1 U3438 ( .A(n6183), .ZN(n6236) );
  NOR2_X1 U3439 ( .A1(n5563), .A2(n5564), .ZN(n5444) );
  NOR2_X1 U3440 ( .A1(n4220), .A2(n4337), .ZN(n2967) );
  AND4_X1 U3441 ( .A1(n3272), .A2(n3271), .A3(n3270), .A4(n3269), .ZN(n2968)
         );
  AND2_X4 U3442 ( .A1(n4536), .A2(n4517), .ZN(n4004) );
  NOR4_X2 U3443 ( .A1(n5794), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .A3(n5314), 
        .A4(n5641), .ZN(n4370) );
  NOR2_X4 U3444 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4541) );
  AND2_X1 U34450 ( .A1(n3067), .A2(n2991), .ZN(n4191) );
  CLKBUF_X1 U34460 ( .A(n5646), .Z(n5647) );
  NOR2_X1 U34480 ( .A1(n4809), .A2(n5987), .ZN(n6592) );
  NAND2_X1 U3449 ( .A1(n3043), .A2(n3571), .ZN(n5966) );
  CLKBUF_X1 U3450 ( .A(n3332), .Z(n4338) );
  INV_X4 U34510 ( .A(n4263), .ZN(n4490) );
  INV_X4 U34520 ( .A(n4234), .ZN(n2969) );
  INV_X1 U34530 ( .A(n4091), .ZN(n3467) );
  AND4_X1 U3454 ( .A1(n3177), .A2(n3176), .A3(n3175), .A4(n3174), .ZN(n2979)
         );
  AND4_X1 U34550 ( .A1(n3173), .A2(n3172), .A3(n3171), .A4(n3170), .ZN(n2986)
         );
  INV_X2 U34560 ( .A(n3424), .ZN(n3995) );
  BUF_X2 U3457 ( .A(n3880), .Z(n3997) );
  BUF_X2 U3458 ( .A(n3418), .Z(n3974) );
  CLKBUF_X2 U34590 ( .A(n4004), .Z(n3875) );
  XNOR2_X1 U34600 ( .A(n4191), .B(n4190), .ZN(n4376) );
  NOR2_X1 U34610 ( .A1(n5660), .A2(n5662), .ZN(n5663) );
  OR2_X1 U34620 ( .A1(n5311), .A2(n3065), .ZN(n5640) );
  AND2_X1 U34630 ( .A1(n3093), .A2(n3047), .ZN(n3074) );
  XNOR2_X1 U34640 ( .A(n4328), .B(n4327), .ZN(n5294) );
  AOI21_X1 U34650 ( .B1(n3095), .B2(n3097), .A(n2996), .ZN(n3094) );
  NAND2_X1 U3466 ( .A1(n2999), .A2(n3099), .ZN(n3097) );
  NAND2_X1 U3467 ( .A1(n3524), .A2(n3523), .ZN(n4829) );
  AND2_X2 U34680 ( .A1(n4121), .A2(n6354), .ZN(n4589) );
  OAI21_X1 U34690 ( .B1(n4142), .B2(n4164), .A(n4141), .ZN(n4143) );
  NAND2_X1 U34700 ( .A1(n4126), .A2(n4125), .ZN(n4127) );
  NAND2_X2 U34710 ( .A1(n4167), .A2(n4166), .ZN(n5760) );
  NAND2_X1 U34720 ( .A1(n3584), .A2(n3583), .ZN(n4167) );
  OAI21_X1 U34730 ( .B1(n5966), .B2(n4164), .A(n4117), .ZN(n4118) );
  NAND2_X1 U34740 ( .A1(n3463), .A2(n3462), .ZN(n3464) );
  CLKBUF_X1 U3475 ( .A(n4534), .Z(n6430) );
  NAND2_X1 U3476 ( .A1(n3144), .A2(n2997), .ZN(n3384) );
  NAND2_X1 U3477 ( .A1(n4262), .A2(n4261), .ZN(n5009) );
  NAND2_X1 U3478 ( .A1(n4448), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4459)
         );
  OAI21_X1 U3479 ( .B1(n5986), .B2(n4164), .A(n4108), .ZN(n4448) );
  NAND2_X2 U3480 ( .A1(n3554), .A2(n3553), .ZN(n5986) );
  CLKBUF_X1 U3481 ( .A(n3558), .Z(n6519) );
  NOR2_X1 U3482 ( .A1(n4642), .A2(n3129), .ZN(n4738) );
  NAND2_X1 U3483 ( .A1(n4241), .A2(n3166), .ZN(n4642) );
  NAND2_X1 U3484 ( .A1(n3416), .A2(n3414), .ZN(n3385) );
  INV_X1 U3485 ( .A(n3103), .ZN(n4509) );
  AND2_X1 U3486 ( .A1(n3056), .A2(n4074), .ZN(n3103) );
  NAND2_X1 U3487 ( .A1(n3347), .A2(n3346), .ZN(n4081) );
  NAND2_X1 U3488 ( .A1(n4230), .A2(n4229), .ZN(n4233) );
  AND2_X1 U3489 ( .A1(n3031), .A2(n3030), .ZN(n4071) );
  NAND2_X1 U3490 ( .A1(n3310), .A2(n3340), .ZN(n4342) );
  NOR2_X1 U3491 ( .A1(n3332), .A2(n4340), .ZN(n4080) );
  NAND2_X2 U3492 ( .A1(n5449), .A2(n4490), .ZN(n4312) );
  CLKBUF_X1 U3493 ( .A(n3319), .Z(n3724) );
  NAND2_X1 U3494 ( .A1(n3325), .A2(n3324), .ZN(n4209) );
  NAND2_X1 U3495 ( .A1(n4042), .A2(n3449), .ZN(n4073) );
  CLKBUF_X1 U3496 ( .A(n3351), .Z(n3352) );
  CLKBUF_X1 U3497 ( .A(n3324), .Z(n4709) );
  NAND2_X1 U3498 ( .A1(n3211), .A2(n4091), .ZN(n3312) );
  CLKBUF_X1 U3499 ( .A(n3326), .Z(n4339) );
  NAND2_X1 U3500 ( .A1(n3324), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3449) );
  NAND2_X1 U3501 ( .A1(n3467), .A2(n3313), .ZN(n4332) );
  NAND2_X1 U3502 ( .A1(n4105), .A2(n3326), .ZN(n4259) );
  INV_X1 U3503 ( .A(n3324), .ZN(n5277) );
  CLKBUF_X1 U3504 ( .A(n3311), .Z(n3333) );
  INV_X1 U3505 ( .A(n3313), .ZN(n4700) );
  NAND2_X2 U3506 ( .A1(n2986), .A2(n2979), .ZN(n4091) );
  NAND2_X2 U3507 ( .A1(n3188), .A2(n3187), .ZN(n3313) );
  NAND4_X2 U3508 ( .A1(n3210), .A2(n3209), .A3(n3208), .A4(n3207), .ZN(n3262)
         );
  AND4_X1 U3509 ( .A1(n3299), .A2(n3298), .A3(n3297), .A4(n3296), .ZN(n3305)
         );
  AND4_X1 U3510 ( .A1(n3229), .A2(n3228), .A3(n3227), .A4(n3226), .ZN(n3245)
         );
  AND4_X1 U3511 ( .A1(n3242), .A2(n3241), .A3(n3240), .A4(n3239), .ZN(n3243)
         );
  AND4_X1 U3512 ( .A1(n3202), .A2(n3201), .A3(n3200), .A4(n3199), .ZN(n3208)
         );
  AND4_X1 U3513 ( .A1(n3221), .A2(n3220), .A3(n3219), .A4(n3218), .ZN(n3222)
         );
  AND4_X1 U3514 ( .A1(n3186), .A2(n3185), .A3(n3184), .A4(n3183), .ZN(n3187)
         );
  AND4_X1 U3515 ( .A1(n3206), .A2(n3205), .A3(n3204), .A4(n3203), .ZN(n3207)
         );
  AND4_X1 U3516 ( .A1(n3276), .A2(n3275), .A3(n3274), .A4(n3273), .ZN(n3283)
         );
  AND4_X1 U3517 ( .A1(n3198), .A2(n3197), .A3(n3196), .A4(n3195), .ZN(n3209)
         );
  AND4_X1 U3518 ( .A1(n3238), .A2(n3237), .A3(n3236), .A4(n3235), .ZN(n3244)
         );
  AND4_X1 U3519 ( .A1(n3181), .A2(n3180), .A3(n3179), .A4(n3178), .ZN(n3188)
         );
  BUF_X2 U3520 ( .A(n3290), .Z(n3959) );
  BUF_X4 U3521 ( .A(n3246), .Z(n2970) );
  BUF_X2 U3522 ( .A(n3225), .Z(n3880) );
  BUF_X2 U3523 ( .A(n3253), .Z(n3931) );
  NAND2_X1 U3524 ( .A1(n3140), .A2(n3139), .ZN(n3374) );
  CLKBUF_X1 U3525 ( .A(n6515), .Z(n6524) );
  AND2_X1 U3526 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3139) );
  AND2_X2 U3527 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4540) );
  CLKBUF_X1 U3528 ( .A(n4588), .Z(n2971) );
  INV_X1 U3529 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n2972) );
  OAI21_X1 U3530 ( .B1(n5760), .B2(n5907), .A(n5903), .ZN(n2973) );
  XNOR2_X1 U3531 ( .A(n4127), .B(n4592), .ZN(n4588) );
  OAI21_X1 U3532 ( .B1(n5760), .B2(n5907), .A(n5903), .ZN(n5734) );
  AND2_X2 U3533 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4542) );
  AND2_X2 U3534 ( .A1(n3064), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4536)
         );
  NOR2_X1 U3535 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3140) );
  NOR2_X1 U3536 ( .A1(n3527), .A2(n3526), .ZN(n3525) );
  NAND2_X1 U3537 ( .A1(n4104), .A2(n4103), .ZN(n4494) );
  AND2_X2 U3538 ( .A1(n3070), .A2(n3074), .ZN(n2984) );
  NOR2_X2 U3539 ( .A1(n4361), .A2(n4495), .ZN(n6402) );
  AND2_X1 U3540 ( .A1(n4541), .A2(n4540), .ZN(n2975) );
  XNOR2_X1 U3541 ( .A(n3543), .B(n3567), .ZN(n4685) );
  NAND2_X1 U3542 ( .A1(n6603), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3030) );
  NAND2_X1 U3543 ( .A1(n4070), .A2(n4087), .ZN(n3031) );
  NAND2_X1 U3544 ( .A1(n4964), .A2(n2981), .ZN(n3040) );
  NAND2_X1 U3545 ( .A1(n5526), .A2(n5249), .ZN(n5523) );
  AND2_X1 U3546 ( .A1(n5248), .A2(n5247), .ZN(n5249) );
  NAND2_X1 U3547 ( .A1(n5235), .A2(n3100), .ZN(n5533) );
  NOR2_X1 U3548 ( .A1(n3101), .A2(n3013), .ZN(n3100) );
  INV_X1 U3549 ( .A(n5234), .ZN(n3101) );
  NOR2_X1 U3550 ( .A1(n4165), .A2(n4164), .ZN(n4166) );
  AOI21_X1 U3551 ( .B1(n3074), .B2(n3075), .A(n3072), .ZN(n3071) );
  INV_X1 U3552 ( .A(n4181), .ZN(n3072) );
  NAND2_X1 U3553 ( .A1(n3124), .A2(n5371), .ZN(n3123) );
  INV_X1 U3554 ( .A(n5361), .ZN(n3124) );
  NAND2_X1 U3555 ( .A1(n2977), .A2(n5395), .ZN(n5383) );
  AND2_X1 U3556 ( .A1(n3009), .A2(n3112), .ZN(n3111) );
  INV_X1 U3557 ( .A(n5206), .ZN(n3112) );
  INV_X1 U3558 ( .A(n3559), .ZN(n4018) );
  OR2_X1 U3559 ( .A1(n4132), .A2(n3623), .ZN(n3539) );
  AND2_X1 U3560 ( .A1(n5783), .A2(n4177), .ZN(n2978) );
  NOR2_X1 U3561 ( .A1(n4340), .A2(n4099), .ZN(n3341) );
  OR2_X1 U3562 ( .A1(n3411), .A2(n3410), .ZN(n4169) );
  INV_X1 U3563 ( .A(n4097), .ZN(n3413) );
  OR2_X1 U3564 ( .A1(n4042), .A2(n4169), .ZN(n3431) );
  NAND2_X1 U3565 ( .A1(n3320), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4042) );
  AND2_X1 U3566 ( .A1(n3333), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3049) );
  AOI22_X1 U3567 ( .A1(n4004), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3264), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3172) );
  AND4_X1 U3568 ( .A1(n3289), .A2(n3288), .A3(n3287), .A4(n3286), .ZN(n3307)
         );
  NAND2_X1 U3569 ( .A1(n6158), .A2(n3019), .ZN(n5504) );
  AND2_X1 U3570 ( .A1(n5533), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5526) );
  NAND2_X1 U3571 ( .A1(n3103), .A2(n3102), .ZN(n5235) );
  NOR2_X1 U3572 ( .A1(n4076), .A2(n6608), .ZN(n3102) );
  AND4_X1 U3573 ( .A1(n3268), .A2(n3267), .A3(n3266), .A4(n3265), .ZN(n3284)
         );
  AND2_X1 U3574 ( .A1(n6527), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4024) );
  INV_X2 U3575 ( .A(n4018), .ZN(n4025) );
  NAND2_X1 U3576 ( .A1(n3723), .A2(n3080), .ZN(n3772) );
  AND2_X1 U3577 ( .A1(n3081), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n3080)
         );
  NOR2_X1 U3578 ( .A1(n5797), .A2(n2994), .ZN(n5315) );
  AND2_X1 U3579 ( .A1(n5836), .A2(n4360), .ZN(n4396) );
  AND2_X1 U3580 ( .A1(n5437), .A2(n5436), .ZN(n5423) );
  NAND2_X1 U3581 ( .A1(n5693), .A2(n3164), .ZN(n5686) );
  NOR2_X1 U3582 ( .A1(n4349), .A2(n4348), .ZN(n4539) );
  NOR2_X1 U3583 ( .A1(n5892), .A2(n6392), .ZN(n5955) );
  CLKBUF_X1 U3584 ( .A(n4216), .Z(n4217) );
  NAND2_X1 U3585 ( .A1(n3103), .A2(n3050), .ZN(n3051) );
  AND2_X1 U3586 ( .A1(n2967), .A2(n4663), .ZN(n3050) );
  AND2_X1 U3587 ( .A1(n6427), .A2(n4917), .ZN(n6478) );
  INV_X1 U3588 ( .A(n5986), .ZN(n5987) );
  OR2_X1 U3589 ( .A1(n4217), .A2(n4098), .ZN(n4648) );
  NAND2_X1 U3590 ( .A1(n3109), .A2(n5293), .ZN(n3037) );
  INV_X1 U3591 ( .A(n3110), .ZN(n3109) );
  OAI21_X1 U3592 ( .B1(n5294), .B2(n6234), .A(n5292), .ZN(n3110) );
  OR2_X1 U3593 ( .A1(n5500), .A2(n5254), .ZN(n5455) );
  AND2_X1 U3594 ( .A1(n5271), .A2(n5270), .ZN(n6183) );
  NAND2_X1 U3595 ( .A1(n4536), .A2(n4516), .ZN(n3182) );
  INV_X1 U3596 ( .A(n3182), .ZN(n3954) );
  AND2_X1 U3597 ( .A1(n5345), .A2(n4044), .ZN(n4057) );
  OR2_X1 U3598 ( .A1(n4038), .A2(n4041), .ZN(n4031) );
  INV_X1 U3599 ( .A(n3827), .ZN(n3424) );
  BUF_X1 U3600 ( .A(n4006), .Z(n3916) );
  AND2_X1 U3601 ( .A1(n3464), .A2(n3127), .ZN(n3126) );
  NOR2_X1 U3602 ( .A1(n3526), .A2(n3128), .ZN(n3127) );
  INV_X1 U3603 ( .A(n3514), .ZN(n3128) );
  INV_X1 U3604 ( .A(n5754), .ZN(n3048) );
  INV_X1 U3605 ( .A(n3097), .ZN(n3096) );
  INV_X1 U3606 ( .A(n3098), .ZN(n3095) );
  AND2_X2 U3607 ( .A1(n4570), .A2(n4541), .ZN(n3277) );
  AOI22_X1 U3608 ( .A1(n3954), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4006), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3255) );
  AND2_X2 U3609 ( .A1(n4540), .A2(n4542), .ZN(n3224) );
  AOI22_X1 U3610 ( .A1(n3247), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3225), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3176) );
  AND2_X1 U3611 ( .A1(n3118), .A2(n3117), .ZN(n3116) );
  INV_X1 U3612 ( .A(n5421), .ZN(n3117) );
  NOR2_X1 U3613 ( .A1(n5469), .A2(n3086), .ZN(n3085) );
  OR2_X1 U3614 ( .A1(n5479), .A2(n5492), .ZN(n5459) );
  INV_X1 U3615 ( .A(n4954), .ZN(n3114) );
  NAND2_X1 U3616 ( .A1(n3581), .A2(n3582), .ZN(n4146) );
  NOR2_X2 U3617 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n4022) );
  NAND2_X1 U3618 ( .A1(n3073), .A2(n3071), .ZN(n4185) );
  INV_X1 U3619 ( .A(n5066), .ZN(n3068) );
  NAND2_X1 U3620 ( .A1(n3003), .A2(n2978), .ZN(n3147) );
  INV_X1 U3621 ( .A(n3149), .ZN(n3148) );
  AND2_X1 U3622 ( .A1(n4273), .A2(n4272), .ZN(n5931) );
  OR2_X1 U3623 ( .A1(n4347), .A2(n4505), .ZN(n4349) );
  INV_X1 U3624 ( .A(n5010), .ZN(n4261) );
  INV_X1 U3625 ( .A(n5008), .ZN(n4262) );
  NAND2_X1 U3626 ( .A1(n4249), .A2(n3130), .ZN(n3129) );
  INV_X1 U3627 ( .A(n4641), .ZN(n3130) );
  NAND2_X1 U3628 ( .A1(n4490), .A2(n2969), .ZN(n4322) );
  INV_X1 U3629 ( .A(n3449), .ZN(n3382) );
  OR2_X1 U3630 ( .A1(n3380), .A2(n3379), .ZN(n3381) );
  INV_X1 U3631 ( .A(n3571), .ZN(n3465) );
  NAND2_X1 U3632 ( .A1(n3448), .A2(n3447), .ZN(n5982) );
  OAI211_X1 U3633 ( .C1(n4061), .C2(n3053), .A(n3052), .B(n4072), .ZN(n3056)
         );
  OR2_X1 U3634 ( .A1(n4210), .A2(n4209), .ZN(n4423) );
  OR2_X1 U3635 ( .A1(n5427), .A2(n5265), .ZN(n5404) );
  NOR2_X1 U3636 ( .A1(n5515), .A2(n3107), .ZN(n6158) );
  NAND2_X1 U3637 ( .A1(n3108), .A2(REIP_REG_8__SCAN_IN), .ZN(n3107) );
  INV_X1 U3638 ( .A(n6192), .ZN(n3108) );
  NOR2_X1 U3639 ( .A1(n6192), .A2(n6734), .ZN(n3028) );
  OR2_X1 U3640 ( .A1(n3820), .A2(n6807), .ZN(n3845) );
  NOR2_X1 U3641 ( .A1(n3083), .A2(n3082), .ZN(n3081) );
  AND2_X1 U3642 ( .A1(n3702), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3723)
         );
  NOR2_X1 U3643 ( .A1(n3687), .A2(n6140), .ZN(n3702) );
  OR2_X1 U3644 ( .A1(n3625), .A2(n3620), .ZN(n3626) );
  INV_X1 U3645 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n6810) );
  NOR2_X1 U3646 ( .A1(n6810), .A2(n3626), .ZN(n3657) );
  AND2_X1 U3647 ( .A1(n4600), .A2(n4792), .ZN(n3580) );
  NAND2_X1 U3648 ( .A1(n3103), .A2(n4663), .ZN(n4652) );
  NAND2_X1 U3649 ( .A1(n5397), .A2(n3141), .ZN(n5242) );
  AND2_X1 U3650 ( .A1(n3012), .A2(n4318), .ZN(n3141) );
  NAND2_X1 U3651 ( .A1(n5397), .A2(n3142), .ZN(n5374) );
  NOR2_X1 U3652 ( .A1(n5372), .A2(n3143), .ZN(n3142) );
  NAND2_X1 U3653 ( .A1(n5397), .A2(n5385), .ZN(n5387) );
  XNOR2_X1 U3654 ( .A(n3008), .B(n3158), .ZN(n3157) );
  INV_X1 U3655 ( .A(n3152), .ZN(n5695) );
  AOI21_X1 U3656 ( .B1(n4378), .B2(n3155), .A(n4381), .ZN(n3153) );
  OR2_X1 U3657 ( .A1(n5709), .A2(n4379), .ZN(n3154) );
  AND2_X1 U3658 ( .A1(n4356), .A2(n3061), .ZN(n3057) );
  AND2_X1 U3659 ( .A1(n4292), .A2(n5466), .ZN(n5464) );
  NOR2_X1 U3660 ( .A1(n3135), .A2(n5467), .ZN(n3134) );
  INV_X1 U3661 ( .A(n5493), .ZN(n3135) );
  INV_X1 U3662 ( .A(n4259), .ZN(n5449) );
  INV_X1 U3663 ( .A(n5569), .ZN(n4284) );
  NAND2_X1 U3664 ( .A1(n5753), .A2(n3098), .ZN(n3046) );
  AND2_X1 U3665 ( .A1(n6392), .A2(n4351), .ZN(n3062) );
  NAND2_X1 U3666 ( .A1(n4174), .A2(n2989), .ZN(n3151) );
  NAND2_X1 U3667 ( .A1(n5067), .A2(n5066), .ZN(n4174) );
  OR2_X1 U3668 ( .A1(n3413), .A2(n4042), .ZN(n3400) );
  OAI211_X1 U3669 ( .C1(n3449), .C2(n3413), .A(n3431), .B(n3412), .ZN(n3540)
         );
  AND2_X1 U3670 ( .A1(n5083), .A2(n6430), .ZN(n6520) );
  XNOR2_X1 U3671 ( .A(n5983), .B(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6467)
         );
  NAND2_X1 U3672 ( .A1(n4582), .A2(n6603), .ZN(n5017) );
  NAND2_X1 U3673 ( .A1(n6605), .A2(n4581), .ZN(n4582) );
  AOI21_X1 U3674 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n6033), .A(n5017), .ZN(
        n6522) );
  AND2_X1 U3675 ( .A1(n4803), .A2(n2976), .ZN(n4751) );
  INV_X1 U3676 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6437) );
  INV_X1 U3677 ( .A(READY_N), .ZN(n6793) );
  OAI21_X1 U3678 ( .B1(n5318), .B2(n6234), .A(n5286), .ZN(n3035) );
  NOR2_X1 U3679 ( .A1(n5355), .A2(n5268), .ZN(n5284) );
  NAND2_X1 U3680 ( .A1(n5380), .A2(n5267), .ZN(n5355) );
  NOR2_X1 U3681 ( .A1(n5455), .A2(n3104), .ZN(n5259) );
  INV_X1 U3682 ( .A(n5256), .ZN(n3105) );
  NOR2_X1 U3683 ( .A1(n5404), .A2(n3032), .ZN(n5380) );
  NAND2_X1 U3684 ( .A1(REIP_REG_24__SCAN_IN), .A2(n5266), .ZN(n3032) );
  NAND2_X1 U3685 ( .A1(n6152), .A2(n3025), .ZN(n5472) );
  NAND2_X1 U3686 ( .A1(n6137), .A2(n5252), .ZN(n5500) );
  NAND2_X1 U3687 ( .A1(n6152), .A2(n5262), .ZN(n6123) );
  INV_X1 U3688 ( .A(n6197), .ZN(n6124) );
  NOR2_X1 U3689 ( .A1(n6616), .A2(n6218), .ZN(n5260) );
  INV_X1 U3690 ( .A(n5523), .ZN(n6216) );
  INV_X1 U3691 ( .A(n6202), .ZN(n6234) );
  INV_X1 U3692 ( .A(n6225), .ZN(n6232) );
  AOI21_X1 U3693 ( .B1(n5526), .B2(n5521), .A(n6197), .ZN(n6239) );
  OAI21_X1 U3694 ( .B1(n4473), .B2(n4092), .A(n4663), .ZN(n4093) );
  XNOR2_X1 U3695 ( .A(n4197), .B(n4196), .ZN(n5271) );
  OR2_X1 U3696 ( .A1(n4195), .A2(n5323), .ZN(n4197) );
  XNOR2_X1 U3697 ( .A(n4027), .B(n4026), .ZN(n5296) );
  AND2_X1 U3698 ( .A1(n5370), .A2(n3014), .ZN(n4027) );
  NAND2_X1 U3699 ( .A1(n3739), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3799)
         );
  NAND2_X1 U3700 ( .A1(n5812), .A2(n3010), .ZN(n5797) );
  INV_X1 U3701 ( .A(n5305), .ZN(n5831) );
  NAND2_X1 U3702 ( .A1(n5334), .A2(n4405), .ZN(n6398) );
  NAND2_X1 U3703 ( .A1(n4350), .A2(n4224), .ZN(n5961) );
  AND2_X1 U3704 ( .A1(n4350), .A2(n4330), .ZN(n6395) );
  INV_X1 U3705 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6033) );
  NAND2_X1 U3706 ( .A1(n3549), .A2(n3550), .ZN(n3554) );
  INV_X1 U3707 ( .A(n6519), .ZN(n5541) );
  INV_X1 U3708 ( .A(n6515), .ZN(n6428) );
  INV_X1 U3709 ( .A(n6430), .ZN(n6474) );
  NAND2_X1 U3710 ( .A1(n4747), .A2(n3442), .ZN(n4721) );
  OAI21_X1 U3711 ( .B1(n3063), .B2(n4339), .A(n3382), .ZN(n3160) );
  OAI211_X1 U3712 ( .C1(n3333), .C2(n3328), .A(n3313), .B(n3312), .ZN(n3332)
         );
  INV_X1 U3713 ( .A(n4070), .ZN(n4053) );
  AND2_X1 U3714 ( .A1(n4064), .A2(n4063), .ZN(n4066) );
  AOI21_X1 U3715 ( .B1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n3442), .A(n4066), 
        .ZN(n4062) );
  INV_X1 U3716 ( .A(n3374), .ZN(n3230) );
  NAND2_X1 U3717 ( .A1(n5760), .A2(n5912), .ZN(n3099) );
  OR2_X1 U3718 ( .A1(n3399), .A2(n3398), .ZN(n4097) );
  OR2_X1 U3719 ( .A1(n3461), .A2(n3460), .ZN(n4124) );
  AOI22_X1 U3720 ( .A1(n3246), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3224), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3174) );
  AOI22_X1 U3721 ( .A1(n3954), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3230), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3177) );
  AND2_X1 U3722 ( .A1(n4056), .A2(n4153), .ZN(n4070) );
  NAND2_X1 U3723 ( .A1(n3055), .A2(n4071), .ZN(n3052) );
  OAI21_X1 U3724 ( .B1(n4060), .B2(n4059), .A(n3001), .ZN(n3055) );
  NAND2_X1 U3725 ( .A1(n3054), .A2(n4071), .ZN(n3053) );
  INV_X1 U3726 ( .A(n4059), .ZN(n3054) );
  AOI221_X1 U3727 ( .B1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n4062), .C1(
        n4475), .C2(n4062), .A(n4036), .ZN(n4084) );
  NOR2_X1 U3728 ( .A1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n6409), .ZN(n4036)
         );
  NAND2_X1 U3729 ( .A1(n3343), .A2(n5277), .ZN(n4076) );
  INV_X1 U3730 ( .A(n4192), .ZN(n3325) );
  OR2_X1 U3731 ( .A1(n3856), .A2(n3855), .ZN(n3869) );
  AND2_X2 U3732 ( .A1(n4570), .A2(n4542), .ZN(n3225) );
  AOI22_X1 U3733 ( .A1(n3418), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3827), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3183) );
  OR2_X1 U3734 ( .A1(n3941), .A2(n3940), .ZN(n3951) );
  INV_X1 U3735 ( .A(n3988), .ZN(n4020) );
  NOR2_X1 U3736 ( .A1(n3845), .A2(n3844), .ZN(n3087) );
  AND2_X1 U3737 ( .A1(n3868), .A2(n3869), .ZN(n3901) );
  AND2_X1 U3738 ( .A1(n3803), .A2(n3119), .ZN(n3118) );
  OR2_X1 U3739 ( .A1(n4518), .A2(n6603), .ZN(n3988) );
  AND2_X1 U3740 ( .A1(n3508), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3517)
         );
  NOR2_X1 U3741 ( .A1(n3572), .A2(n3079), .ZN(n3508) );
  NAND2_X1 U3742 ( .A1(n3066), .A2(n4369), .ZN(n3065) );
  INV_X1 U3743 ( .A(n5668), .ZN(n3066) );
  INV_X1 U3744 ( .A(n5385), .ZN(n3143) );
  NOR2_X1 U3745 ( .A1(n5762), .A2(n4380), .ZN(n4381) );
  NOR2_X1 U3746 ( .A1(n3062), .A2(n3022), .ZN(n3061) );
  AOI21_X1 U3747 ( .B1(n3094), .B2(n3096), .A(n2993), .ZN(n3093) );
  NAND2_X1 U3748 ( .A1(n3048), .A2(n3094), .ZN(n3047) );
  INV_X1 U3749 ( .A(n3094), .ZN(n3075) );
  AND2_X1 U3750 ( .A1(n4178), .A2(n3099), .ZN(n3098) );
  NOR2_X1 U3751 ( .A1(n5784), .A2(n3150), .ZN(n3149) );
  INV_X1 U3752 ( .A(n4175), .ZN(n3150) );
  AND2_X1 U3753 ( .A1(n3326), .A2(n4099), .ZN(n4153) );
  INV_X1 U3754 ( .A(n4153), .ZN(n4164) );
  OR2_X1 U3755 ( .A1(n3417), .A2(n4042), .ZN(n4165) );
  OR2_X1 U3756 ( .A1(n3430), .A2(n3429), .ZN(n4106) );
  AND2_X2 U3757 ( .A1(n3036), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4517)
         );
  INV_X1 U3758 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3036) );
  NAND2_X1 U3759 ( .A1(n3724), .A2(n4099), .ZN(n4518) );
  INV_X1 U3760 ( .A(n2976), .ZN(n5979) );
  OR2_X2 U3762 ( .A1(n3259), .A2(n3258), .ZN(n4105) );
  INV_X1 U3763 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n5087) );
  NOR2_X1 U3764 ( .A1(n5246), .A2(n3326), .ZN(n3350) );
  INV_X1 U3765 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n3844) );
  NOR2_X1 U3766 ( .A1(n5264), .A2(n3026), .ZN(n3025) );
  INV_X1 U3767 ( .A(n5262), .ZN(n3026) );
  CLKBUF_X1 U3768 ( .A(n4113), .Z(n5273) );
  NOR2_X1 U3769 ( .A1(n3125), .A2(n3123), .ZN(n3122) );
  INV_X1 U3770 ( .A(n5350), .ZN(n3125) );
  INV_X1 U3771 ( .A(n5233), .ZN(n3120) );
  NOR2_X1 U3772 ( .A1(n3078), .A2(n3947), .ZN(n3076) );
  INV_X1 U3773 ( .A(n3123), .ZN(n3121) );
  AND2_X1 U3774 ( .A1(n3945), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n3946)
         );
  NAND2_X1 U3775 ( .A1(n3946), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n3990)
         );
  NAND2_X1 U3776 ( .A1(n3905), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n3944)
         );
  INV_X1 U3777 ( .A(n3907), .ZN(n3905) );
  NAND2_X1 U3778 ( .A1(n3087), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n3907)
         );
  INV_X1 U3779 ( .A(n3087), .ZN(n3873) );
  INV_X1 U3780 ( .A(n5297), .ZN(n3039) );
  AND2_X1 U3781 ( .A1(n3018), .A2(n3085), .ZN(n3084) );
  INV_X1 U3782 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5469) );
  NAND2_X1 U3783 ( .A1(n3739), .A2(n3085), .ZN(n3804) );
  INV_X1 U3784 ( .A(n3772), .ZN(n3739) );
  NAND2_X1 U3785 ( .A1(n3723), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3738)
         );
  AND2_X1 U3786 ( .A1(n3711), .A2(n3685), .ZN(n5750) );
  OR2_X1 U3787 ( .A1(n3671), .A2(n6150), .ZN(n3687) );
  AND3_X1 U3788 ( .A1(n3654), .A2(n3653), .A3(n3652), .ZN(n3655) );
  AND3_X1 U3789 ( .A1(n3639), .A2(n3638), .A3(n3637), .ZN(n3640) );
  INV_X1 U3790 ( .A(n4791), .ZN(n3041) );
  AND3_X1 U3791 ( .A1(n3607), .A2(n3606), .A3(n3605), .ZN(n4954) );
  NAND2_X1 U3792 ( .A1(n3588), .A2(n3007), .ZN(n3619) );
  NAND2_X1 U3793 ( .A1(n3513), .A2(n3512), .ZN(n4792) );
  AND2_X1 U3794 ( .A1(n3517), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3588)
         );
  NAND2_X1 U3795 ( .A1(n3516), .A2(n3711), .ZN(n3524) );
  NAND2_X1 U3796 ( .A1(PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n3572) );
  NAND2_X1 U3797 ( .A1(n4479), .A2(n3576), .ZN(n4604) );
  NAND2_X1 U3798 ( .A1(n5242), .A2(n2969), .ZN(n5240) );
  NAND2_X1 U3799 ( .A1(n5311), .A2(n5313), .ZN(n5639) );
  AND2_X1 U3800 ( .A1(n4315), .A2(n4314), .ZN(n5363) );
  NOR2_X1 U3801 ( .A1(n5760), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5667)
         );
  INV_X1 U3802 ( .A(n5311), .ZN(n5671) );
  AND2_X1 U3803 ( .A1(n5396), .A2(n4307), .ZN(n5397) );
  NOR2_X2 U3804 ( .A1(n5302), .A2(n5301), .ZN(n5396) );
  AND2_X1 U3805 ( .A1(n5570), .A2(n3132), .ZN(n5437) );
  NOR2_X1 U3806 ( .A1(n4295), .A2(n3133), .ZN(n3132) );
  INV_X1 U3807 ( .A(n3134), .ZN(n3133) );
  NOR2_X1 U3808 ( .A1(n5762), .A2(n4377), .ZN(n4378) );
  NOR2_X1 U3809 ( .A1(n2984), .A2(n5709), .ZN(n5708) );
  AND2_X1 U3810 ( .A1(n4288), .A2(n4287), .ZN(n5493) );
  AND3_X1 U3811 ( .A1(n4283), .A2(n4282), .A3(n4281), .ZN(n5569) );
  CLKBUF_X1 U3812 ( .A(n5577), .Z(n5587) );
  NAND2_X1 U3813 ( .A1(n2978), .A2(n2989), .ZN(n3089) );
  AND2_X1 U3814 ( .A1(n3147), .A2(n3069), .ZN(n3088) );
  NOR2_X2 U3815 ( .A1(n5009), .A2(n3136), .ZN(n5929) );
  NAND2_X1 U3816 ( .A1(n3138), .A2(n2980), .ZN(n3136) );
  OR2_X1 U3817 ( .A1(n5009), .A2(n3137), .ZN(n5934) );
  NAND2_X1 U3818 ( .A1(n4172), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4173)
         );
  CLKBUF_X1 U3819 ( .A(n5008), .Z(n5063) );
  CLKBUF_X1 U3820 ( .A(n4967), .Z(n4968) );
  XNOR2_X1 U3821 ( .A(n4161), .B(n6386), .ZN(n5158) );
  CLKBUF_X1 U3823 ( .A(n4738), .Z(n4795) );
  XNOR2_X1 U3824 ( .A(n4150), .B(n6780), .ZN(n4846) );
  INV_X1 U3825 ( .A(n4593), .ZN(n4241) );
  CLKBUF_X1 U3826 ( .A(n4593), .Z(n4607) );
  OR2_X1 U3827 ( .A1(n5918), .A2(n5922), .ZN(n5892) );
  INV_X1 U3828 ( .A(n5892), .ZN(n4361) );
  NAND2_X1 U3829 ( .A1(n4488), .A2(n4490), .ZN(n4489) );
  OR2_X1 U3830 ( .A1(n4208), .A2(n5345), .ZN(n4537) );
  AND2_X1 U3831 ( .A1(n4350), .A2(n4650), .ZN(n5918) );
  CLKBUF_X1 U3832 ( .A(n4514), .Z(n4515) );
  NAND2_X1 U3833 ( .A1(n3438), .A2(n3437), .ZN(n3568) );
  AND2_X2 U3834 ( .A1(n3169), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4516)
         );
  INV_X1 U3835 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3064) );
  CLKBUF_X1 U3836 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n4556) );
  AND2_X1 U3837 ( .A1(n4894), .A2(n6410), .ZN(n4895) );
  INV_X1 U3838 ( .A(n4105), .ZN(n3321) );
  OR2_X1 U3839 ( .A1(n5017), .A2(n6437), .ZN(n4720) );
  AND2_X1 U3840 ( .A1(n4629), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4075) );
  OR2_X1 U3841 ( .A1(n4208), .A2(n4192), .ZN(n4622) );
  INV_X1 U3842 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6527) );
  NAND2_X1 U3843 ( .A1(n5235), .A2(n5234), .ZN(n6679) );
  NOR2_X1 U3844 ( .A1(n5404), .A2(n6647), .ZN(n5403) );
  OR2_X1 U3845 ( .A1(n3027), .A2(n6643), .ZN(n5427) );
  OAI21_X1 U3846 ( .B1(n5504), .B2(n5250), .A(n6217), .ZN(n6137) );
  INV_X1 U3847 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n6140) );
  INV_X1 U3848 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n6150) );
  NOR2_X1 U3849 ( .A1(n6176), .A2(n5261), .ZN(n6152) );
  OR2_X1 U3850 ( .A1(n3029), .A2(n6623), .ZN(n6176) );
  INV_X1 U3851 ( .A(n6219), .ZN(n6181) );
  AND2_X1 U3852 ( .A1(n5291), .A2(n5245), .ZN(n6202) );
  AND2_X1 U3853 ( .A1(n5533), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6225) );
  NAND2_X1 U3854 ( .A1(n5523), .A2(n5533), .ZN(n6217) );
  INV_X1 U3855 ( .A(n5590), .ZN(n6248) );
  INV_X1 U3856 ( .A(n5588), .ZN(n6247) );
  INV_X1 U3857 ( .A(n6250), .ZN(n5595) );
  AND2_X1 U3858 ( .A1(n4487), .A2(n4663), .ZN(n6250) );
  INV_X1 U3859 ( .A(n6248), .ZN(n5597) );
  NOR2_X2 U3860 ( .A1(n6253), .A2(n3352), .ZN(n6251) );
  AND2_X1 U3861 ( .A1(n6261), .A2(n5341), .ZN(n6254) );
  AND2_X1 U3862 ( .A1(n6261), .A2(n4456), .ZN(n6257) );
  INV_X1 U3863 ( .A(n6257), .ZN(n4844) );
  NAND2_X1 U3864 ( .A1(n4653), .A2(n6603), .ZN(n6280) );
  OR2_X1 U3865 ( .A1(n6274), .A2(n6681), .ZN(n6281) );
  OR3_X1 U3866 ( .A1(n4652), .A2(n4651), .A3(n6082), .ZN(n6288) );
  INV_X2 U3867 ( .A(n6280), .ZN(n6681) );
  INV_X2 U3868 ( .A(n6281), .ZN(n6286) );
  OR2_X1 U3869 ( .A1(n5235), .A2(n4077), .ZN(n6307) );
  INV_X1 U3870 ( .A(n6348), .ZN(n6343) );
  INV_X1 U3871 ( .A(n6307), .ZN(n6346) );
  OR2_X1 U3872 ( .A1(n4652), .A2(n4648), .ZN(n6348) );
  OAI21_X1 U3873 ( .B1(n5348), .B2(n5350), .A(n5349), .ZN(n5645) );
  OAI21_X1 U3874 ( .B1(n3165), .B2(n5462), .A(n5461), .ZN(n5715) );
  NAND2_X1 U3875 ( .A1(n3723), .A2(n3081), .ZN(n3770) );
  NAND2_X1 U3876 ( .A1(n5775), .A2(n4457), .ZN(n6362) );
  OR2_X1 U3877 ( .A1(n4652), .A2(n4622), .ZN(n6092) );
  INV_X1 U3878 ( .A(n6362), .ZN(n5778) );
  INV_X2 U3879 ( .A(n5782), .ZN(n6358) );
  INV_X1 U3880 ( .A(n6398), .ZN(n6350) );
  NAND2_X1 U3881 ( .A1(n4406), .A2(n6524), .ZN(n5782) );
  INV_X1 U3882 ( .A(n5775), .ZN(n6351) );
  XNOR2_X1 U3883 ( .A(n3090), .B(n5314), .ZN(n5329) );
  NAND2_X1 U3884 ( .A1(n3092), .A2(n3091), .ZN(n3090) );
  NAND2_X1 U3885 ( .A1(n5639), .A2(n5641), .ZN(n3091) );
  NAND2_X1 U3886 ( .A1(n5640), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n3092) );
  NOR2_X1 U3887 ( .A1(n5831), .A2(n2995), .ZN(n5812) );
  OR2_X1 U3888 ( .A1(n4397), .A2(n4367), .ZN(n5828) );
  AND2_X1 U3889 ( .A1(n5886), .A2(n4365), .ZN(n5854) );
  AND2_X1 U3890 ( .A1(n4396), .A2(n4362), .ZN(n5305) );
  XNOR2_X1 U3891 ( .A(n3005), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n3159)
         );
  NAND2_X1 U3892 ( .A1(n4384), .A2(n4385), .ZN(n3045) );
  NAND2_X1 U3893 ( .A1(n4383), .A2(n5762), .ZN(n4384) );
  NAND2_X1 U3894 ( .A1(n5570), .A2(n3134), .ZN(n5448) );
  NOR2_X1 U3895 ( .A1(n5070), .A2(n3059), .ZN(n5881) );
  INV_X1 U3896 ( .A(n3062), .ZN(n3060) );
  AND2_X1 U3897 ( .A1(n6365), .A2(n4364), .ZN(n5886) );
  INV_X1 U3898 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5907) );
  NAND2_X1 U3899 ( .A1(n5924), .A2(n5946), .ZN(n6365) );
  NAND2_X1 U3900 ( .A1(n3151), .A2(n4175), .ZN(n5786) );
  INV_X1 U3901 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n5075) );
  AND2_X1 U3902 ( .A1(n4443), .A2(n4442), .ZN(n4496) );
  INV_X1 U3903 ( .A(n5961), .ZN(n6403) );
  INV_X1 U3904 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n4629) );
  CLKBUF_X1 U3905 ( .A(n4516), .Z(n4521) );
  AOI21_X1 U3906 ( .B1(n6603), .B2(STATE2_REG_3__SCAN_IN), .A(n4477), .ZN(
        n5977) );
  NOR2_X1 U3907 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n5334) );
  NAND4_X1 U3908 ( .A1(n4920), .A2(n6478), .A3(n6435), .A4(n4919), .ZN(n4946)
         );
  AND2_X1 U3909 ( .A1(n4921), .A2(n5987), .ZN(n5154) );
  INV_X1 U3910 ( .A(n6423), .ZN(n4914) );
  OR2_X1 U3911 ( .A1(n6439), .A2(n6438), .ZN(n6850) );
  OAI211_X1 U3912 ( .C1(n6515), .C2(n6032), .A(n6522), .B(n4691), .ZN(n4719)
         );
  INV_X1 U3913 ( .A(n6585), .ZN(n6001) );
  INV_X1 U3914 ( .A(n6846), .ZN(n6021) );
  AND2_X1 U3915 ( .A1(n5171), .A2(n5987), .ZN(n5202) );
  AOI22_X1 U3916 ( .A1(n5086), .A2(n6520), .B1(n5085), .B2(n6465), .ZN(n5117)
         );
  INV_X1 U3917 ( .A(n6530), .ZN(n5997) );
  INV_X1 U3918 ( .A(n6549), .ZN(n6009) );
  INV_X1 U3919 ( .A(n6556), .ZN(n6013) );
  INV_X1 U3920 ( .A(n6563), .ZN(n6017) );
  INV_X1 U3921 ( .A(n6592), .ZN(n5004) );
  INV_X1 U3922 ( .A(n6512), .ZN(n6470) );
  NOR2_X1 U3923 ( .A1(n4708), .A2(n5017), .ZN(n6530) );
  INV_X1 U3924 ( .A(n6534), .ZN(n6584) );
  NOR2_X1 U3925 ( .A1(n4704), .A2(n5017), .ZN(n6585) );
  INV_X1 U3926 ( .A(n6546), .ZN(n6489) );
  NOR2_X1 U3927 ( .A1(n6720), .A2(n5017), .ZN(n6549) );
  NOR2_X1 U3928 ( .A1(n4733), .A2(n5017), .ZN(n6556) );
  INV_X1 U3929 ( .A(n6560), .ZN(n6497) );
  NOR2_X1 U3930 ( .A1(n4841), .A2(n5017), .ZN(n6563) );
  INV_X1 U3931 ( .A(n6573), .ZN(n6504) );
  NOR2_X1 U3932 ( .A1(n4699), .A2(n5017), .ZN(n6578) );
  INV_X1 U3933 ( .A(n6513), .ZN(n6480) );
  INV_X1 U3934 ( .A(n6538), .ZN(n6586) );
  INV_X1 U3935 ( .A(n6539), .ZN(n6485) );
  NOR2_X1 U3936 ( .A1(n4687), .A2(n5017), .ZN(n6542) );
  INV_X1 U3937 ( .A(n6540), .ZN(n6486) );
  INV_X1 U3938 ( .A(n6547), .ZN(n6490) );
  INV_X1 U3939 ( .A(n6561), .ZN(n6498) );
  NAND2_X1 U3940 ( .A1(n6358), .A2(DATAI_30_), .ZN(n6854) );
  INV_X1 U3941 ( .A(n6567), .ZN(n6845) );
  NOR2_X1 U3942 ( .A1(n4843), .A2(n5017), .ZN(n6846) );
  INV_X1 U3943 ( .A(n6568), .ZN(n6849) );
  INV_X1 U3944 ( .A(n6582), .ZN(n6507) );
  OR2_X1 U3945 ( .A1(n4720), .A2(n4700), .ZN(n6573) );
  OAI211_X1 U3946 ( .C1(n4750), .C2(n4752), .A(n6522), .B(n4749), .ZN(n4784)
         );
  OR2_X1 U3947 ( .A1(n4509), .A2(n6437), .ZN(n6605) );
  AND3_X1 U3948 ( .A1(n6603), .A2(STATEBS16_REG_SCAN_IN), .A3(
        STATE2_REG_1__SCAN_IN), .ZN(n4406) );
  INV_X1 U3949 ( .A(n4658), .ZN(n4405) );
  NOR2_X1 U3950 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6683) );
  INV_X1 U3951 ( .A(n6669), .ZN(n6665) );
  NOR2_X2 U3952 ( .A1(STATE_REG_0__SCAN_IN), .A2(n6800), .ZN(n6688) );
  NAND2_X1 U3953 ( .A1(n3038), .A2(n2992), .ZN(U2796) );
  NAND2_X1 U3954 ( .A1(n5296), .A2(n6197), .ZN(n3038) );
  INV_X1 U3955 ( .A(n3035), .ZN(n3034) );
  NAND2_X1 U3956 ( .A1(n5322), .A2(n6197), .ZN(n3033) );
  INV_X1 U3957 ( .A(n5259), .ZN(n5367) );
  AND2_X1 U3958 ( .A1(n6216), .A2(n5260), .ZN(n6210) );
  AND2_X1 U3959 ( .A1(n4374), .A2(n4373), .ZN(n4375) );
  AND2_X2 U3960 ( .A1(n5444), .A2(n3011), .ZN(n2977) );
  NAND2_X1 U3961 ( .A1(n3113), .A2(n3009), .ZN(n5005) );
  INV_X1 U3962 ( .A(n4259), .ZN(n4234) );
  AND2_X2 U3963 ( .A1(n4570), .A2(n4536), .ZN(n3295) );
  NAND2_X1 U3964 ( .A1(n2974), .A2(n3118), .ZN(n5420) );
  INV_X2 U3965 ( .A(n3479), .ZN(n3455) );
  AND2_X1 U3966 ( .A1(n5930), .A2(n5931), .ZN(n2980) );
  AND2_X1 U3967 ( .A1(n3111), .A2(n3168), .ZN(n2981) );
  NAND2_X1 U3968 ( .A1(n2974), .A2(n3006), .ZN(n4386) );
  NAND2_X1 U3969 ( .A1(n3041), .A2(n4964), .ZN(n4953) );
  INV_X1 U3970 ( .A(n5258), .ZN(n3106) );
  OR2_X1 U3971 ( .A1(n3065), .A2(n3020), .ZN(n2982) );
  NAND2_X1 U3972 ( .A1(n3467), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3623) );
  INV_X1 U3973 ( .A(n3623), .ZN(n3711) );
  AND2_X1 U3974 ( .A1(n3025), .A2(n3021), .ZN(n2983) );
  NAND2_X1 U3976 ( .A1(n5570), .A2(n5493), .ZN(n5463) );
  OR2_X1 U3977 ( .A1(n5455), .A2(n5256), .ZN(n2985) );
  NAND2_X1 U3978 ( .A1(n2974), .A2(n3803), .ZN(n5433) );
  INV_X1 U3979 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n5338) );
  AND4_X1 U3980 ( .A1(n3234), .A2(n3233), .A3(n3232), .A4(n3231), .ZN(n2987)
         );
  OR2_X1 U3981 ( .A1(n5760), .A2(n6764), .ZN(n2988) );
  NAND2_X1 U3982 ( .A1(n5753), .A2(n4178), .ZN(n5744) );
  AND2_X1 U3983 ( .A1(n2988), .A2(n4173), .ZN(n2989) );
  NOR2_X1 U3984 ( .A1(n4953), .A2(n4954), .ZN(n4955) );
  AND2_X1 U3985 ( .A1(n2974), .A2(n3116), .ZN(n2990) );
  NOR2_X1 U3986 ( .A1(n5311), .A2(n5668), .ZN(n5660) );
  NAND2_X1 U3987 ( .A1(n5678), .A2(n4189), .ZN(n2991) );
  NOR2_X1 U3988 ( .A1(n5295), .A2(n3037), .ZN(n2992) );
  INV_X1 U3989 ( .A(n3042), .ZN(n3576) );
  OAI21_X1 U3990 ( .B1(n5966), .B2(n3623), .A(n3672), .ZN(n3042) );
  AND2_X1 U3991 ( .A1(n5716), .A2(n4180), .ZN(n2993) );
  AND2_X1 U3992 ( .A1(n5894), .A2(n5641), .ZN(n2994) );
  AND2_X1 U3993 ( .A1(n5894), .A2(n4368), .ZN(n2995) );
  AND2_X1 U3994 ( .A1(n5760), .A2(n4179), .ZN(n2996) );
  OR2_X1 U3995 ( .A1(n4112), .A2(n4042), .ZN(n2997) );
  NAND2_X1 U3996 ( .A1(n5769), .A2(n4176), .ZN(n2998) );
  AND2_X1 U3997 ( .A1(n5716), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n2999)
         );
  INV_X1 U3998 ( .A(n4953), .ZN(n3113) );
  OR2_X1 U3999 ( .A1(n5070), .A2(n3062), .ZN(n3000) );
  NAND2_X1 U4000 ( .A1(n4087), .A2(n4069), .ZN(n3001) );
  NAND2_X1 U4001 ( .A1(n3151), .A2(n3149), .ZN(n3002) );
  INV_X1 U4002 ( .A(n3138), .ZN(n3137) );
  NOR2_X1 U4003 ( .A1(n5209), .A2(n5230), .ZN(n3138) );
  OR2_X1 U4004 ( .A1(n2998), .A2(n3148), .ZN(n3003) );
  NOR2_X1 U4005 ( .A1(n5708), .A2(n4378), .ZN(n3004) );
  NAND2_X1 U4006 ( .A1(n3113), .A2(n3111), .ZN(n3115) );
  INV_X1 U4007 ( .A(n4379), .ZN(n3155) );
  NAND2_X1 U4008 ( .A1(n4474), .A2(n3369), .ZN(n4555) );
  AND2_X1 U4009 ( .A1(n4350), .A2(n4539), .ZN(n6392) );
  OR3_X1 U4010 ( .A1(n5716), .A2(n6786), .A3(n6783), .ZN(n3005) );
  OR2_X1 U4011 ( .A1(n5009), .A2(n5209), .ZN(n5210) );
  AND2_X1 U4012 ( .A1(n3116), .A2(n4387), .ZN(n3006) );
  AND2_X1 U4013 ( .A1(PHYADDRPOINTER_REG_6__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3007) );
  OR3_X1 U4014 ( .A1(n5762), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n3008) );
  NOR2_X1 U4015 ( .A1(n4496), .A2(n6392), .ZN(n5070) );
  INV_X1 U4016 ( .A(n5070), .ZN(n3058) );
  AND2_X1 U4017 ( .A1(n3114), .A2(n5006), .ZN(n3009) );
  OR2_X1 U4018 ( .A1(n5955), .A2(n4369), .ZN(n3010) );
  NAND2_X1 U4019 ( .A1(n6152), .A2(n2983), .ZN(n3027) );
  OR2_X1 U4020 ( .A1(n4642), .A2(n4641), .ZN(n3131) );
  AND2_X1 U4021 ( .A1(n3006), .A2(n3039), .ZN(n3011) );
  NAND2_X1 U4022 ( .A1(n4075), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6608) );
  NOR3_X1 U4023 ( .A1(n5372), .A2(n5363), .A3(n3143), .ZN(n3012) );
  NAND3_X1 U4024 ( .A1(n5237), .A2(n6398), .A3(n6599), .ZN(n3013) );
  NAND2_X1 U4025 ( .A1(n3946), .A2(n3076), .ZN(n3077) );
  AND2_X1 U4026 ( .A1(n3122), .A2(n3120), .ZN(n3014) );
  OR2_X1 U4027 ( .A1(n5523), .A2(n5267), .ZN(n3015) );
  AND2_X1 U4028 ( .A1(n3007), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3016)
         );
  INV_X2 U4029 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6603) );
  INV_X1 U4030 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3079) );
  INV_X1 U4031 ( .A(n5434), .ZN(n3119) );
  INV_X1 U4032 ( .A(n3264), .ZN(n3423) );
  AND2_X2 U4033 ( .A1(n5338), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4545)
         );
  AND2_X1 U4034 ( .A1(n3588), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3017)
         );
  AND2_X1 U4035 ( .A1(PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n3018) );
  INV_X1 U4036 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3082) );
  AND3_X1 U4037 ( .A1(REIP_REG_11__SCAN_IN), .A2(REIP_REG_9__SCAN_IN), .A3(
        REIP_REG_10__SCAN_IN), .ZN(n3019) );
  OR2_X1 U4038 ( .A1(n5314), .A2(n5641), .ZN(n3020) );
  AND2_X1 U4039 ( .A1(REIP_REG_20__SCAN_IN), .A2(REIP_REG_19__SCAN_IN), .ZN(
        n3021) );
  NAND2_X1 U4040 ( .A1(n4365), .A2(n5837), .ZN(n3022) );
  AND2_X1 U4041 ( .A1(n3076), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n3023)
         );
  INV_X1 U4042 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n3158) );
  INV_X1 U4043 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3086) );
  CLKBUF_X1 U4044 ( .A(n6847), .Z(n3024) );
  AND2_X4 U4045 ( .A1(n4570), .A2(n4545), .ZN(n3290) );
  NAND3_X1 U4046 ( .A1(n6216), .A2(n5260), .A3(REIP_REG_5__SCAN_IN), .ZN(n6194) );
  NAND3_X1 U4047 ( .A1(n6216), .A2(n5260), .A3(n3028), .ZN(n3029) );
  INV_X1 U4048 ( .A(n3029), .ZN(n6186) );
  NAND3_X1 U4049 ( .A1(n5285), .A2(n3034), .A3(n3033), .ZN(U2797) );
  NOR2_X2 U4050 ( .A1(n4791), .A2(n3040), .ZN(n5228) );
  NAND2_X1 U4051 ( .A1(n5228), .A2(n5591), .ZN(n5573) );
  NAND3_X1 U4052 ( .A1(n3570), .A2(n3569), .A3(n3566), .ZN(n3043) );
  AND2_X2 U4053 ( .A1(n4541), .A2(n4540), .ZN(n3253) );
  NAND2_X1 U4054 ( .A1(n3044), .A2(n3167), .ZN(U2963) );
  NAND2_X1 U4055 ( .A1(n4391), .A2(n4193), .ZN(n3044) );
  NAND2_X1 U4056 ( .A1(n5716), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5783) );
  NAND2_X1 U4057 ( .A1(n3046), .A2(n3097), .ZN(n5740) );
  NAND2_X1 U4058 ( .A1(n5755), .A2(n5754), .ZN(n5753) );
  NOR2_X4 U4059 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4570) );
  NAND2_X1 U4060 ( .A1(n5760), .A2(n4352), .ZN(n4178) );
  AND2_X2 U4061 ( .A1(n3049), .A2(n5277), .ZN(n4056) );
  AND2_X1 U4062 ( .A1(n4350), .A2(n4349), .ZN(n5922) );
  NAND2_X2 U4063 ( .A1(n4221), .A2(n3051), .ZN(n4350) );
  NAND2_X1 U4064 ( .A1(n3058), .A2(n3057), .ZN(n4358) );
  NAND2_X1 U4065 ( .A1(n4356), .A2(n3060), .ZN(n3059) );
  INV_X1 U4066 ( .A(n3063), .ZN(n3347) );
  OAI211_X1 U4067 ( .C1(n3263), .C2(n3319), .A(n3261), .B(n3260), .ZN(n3063)
         );
  INV_X1 U4068 ( .A(n3347), .ZN(n4210) );
  OR2_X2 U4069 ( .A1(n5311), .A2(n2982), .ZN(n3067) );
  NAND3_X1 U4070 ( .A1(n2989), .A2(n2978), .A3(n3068), .ZN(n3069) );
  NAND2_X1 U4071 ( .A1(n5755), .A2(n3074), .ZN(n3073) );
  NAND2_X1 U4072 ( .A1(n5760), .A2(n4171), .ZN(n4172) );
  NAND2_X1 U4073 ( .A1(n3946), .A2(n3023), .ZN(n4195) );
  INV_X1 U4074 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n3078) );
  NAND2_X1 U4075 ( .A1(n3588), .A2(n3016), .ZN(n3625) );
  INV_X1 U4076 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3083) );
  NAND2_X1 U4077 ( .A1(n3739), .A2(n3084), .ZN(n3820) );
  NOR2_X2 U4078 ( .A1(n5271), .A2(n5269), .ZN(n6197) );
  NAND2_X1 U4079 ( .A1(n3465), .A2(n3464), .ZN(n3527) );
  OAI21_X2 U4080 ( .B1(n5067), .B2(n3089), .A(n3088), .ZN(n5755) );
  NAND2_X2 U4081 ( .A1(n4163), .A2(n4162), .ZN(n5067) );
  NOR3_X1 U4082 ( .A1(n5455), .A2(n5256), .A3(n3106), .ZN(n5389) );
  NAND3_X1 U4083 ( .A1(n5258), .A2(n3105), .A3(n3015), .ZN(n3104) );
  NAND2_X1 U4084 ( .A1(n3313), .A2(n4091), .ZN(n3351) );
  INV_X1 U4085 ( .A(n3115), .ZN(n5205) );
  AND2_X1 U4086 ( .A1(n5370), .A2(n3121), .ZN(n5348) );
  NAND2_X1 U4087 ( .A1(n5370), .A2(n3122), .ZN(n5349) );
  NAND2_X1 U4088 ( .A1(n5370), .A2(n5371), .ZN(n5360) );
  NAND2_X1 U4089 ( .A1(n3465), .A2(n3126), .ZN(n3581) );
  INV_X1 U4090 ( .A(n3131), .ZN(n4737) );
  AND2_X1 U4091 ( .A1(n5397), .A2(n3012), .ZN(n5362) );
  NAND3_X1 U4092 ( .A1(n3440), .A2(n6603), .A3(n3369), .ZN(n3144) );
  NAND2_X1 U4093 ( .A1(n3145), .A2(n3146), .ZN(n3440) );
  INV_X1 U4094 ( .A(n3368), .ZN(n3145) );
  INV_X1 U4095 ( .A(n3367), .ZN(n3146) );
  NAND2_X1 U4096 ( .A1(n4174), .A2(n4173), .ZN(n5222) );
  NAND2_X1 U4097 ( .A1(n3290), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3195) );
  OAI21_X2 U4098 ( .B1(n2984), .B2(n3154), .A(n3153), .ZN(n3152) );
  NAND2_X1 U4099 ( .A1(n5686), .A2(n3157), .ZN(n3156) );
  OAI21_X1 U4100 ( .B1(n5686), .B2(n3159), .A(n3156), .ZN(n5310) );
  NAND3_X1 U4101 ( .A1(n3161), .A2(n3316), .A3(n3160), .ZN(n3363) );
  NAND2_X1 U4102 ( .A1(n3162), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3161) );
  NAND4_X1 U4103 ( .A1(n4080), .A2(n3314), .A3(n3336), .A4(n4342), .ZN(n3162)
         );
  NAND2_X1 U4104 ( .A1(n4113), .A2(n3340), .ZN(n3336) );
  NAND2_X2 U4105 ( .A1(n4187), .A2(n4186), .ZN(n5311) );
  NAND2_X1 U4106 ( .A1(n3362), .A2(n3386), .ZN(n3368) );
  NOR2_X1 U4107 ( .A1(n4332), .A2(n3320), .ZN(n3319) );
  NAND2_X1 U4108 ( .A1(n3328), .A2(n4105), .ZN(n3260) );
  INV_X1 U4109 ( .A(n3541), .ZN(n3438) );
  NOR2_X2 U4110 ( .A1(n5383), .A2(n5384), .ZN(n5370) );
  OAI21_X1 U4111 ( .B1(n5693), .B2(INSTADDRPOINTER_REG_22__SCAN_IN), .A(n5716), 
        .ZN(n4385) );
  NOR2_X1 U4112 ( .A1(n5966), .A2(n4684), .ZN(n5980) );
  AND2_X2 U4113 ( .A1(n3345), .A2(n5246), .ZN(n4113) );
  NOR2_X1 U4114 ( .A1(n4423), .A2(n3345), .ZN(n4650) );
  OR2_X1 U4115 ( .A1(n4518), .A2(n3345), .ZN(n4348) );
  AND2_X1 U4116 ( .A1(n4334), .A2(n3345), .ZN(n3346) );
  NAND2_X1 U4117 ( .A1(n5296), .A2(n4094), .ZN(n4096) );
  INV_X1 U4118 ( .A(n5635), .ZN(n6258) );
  NAND2_X2 U4119 ( .A1(n6261), .A2(n4455), .ZN(n5635) );
  OR2_X1 U4120 ( .A1(n3358), .A2(n4556), .ZN(n3163) );
  OR2_X1 U4121 ( .A1(n5716), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n3164)
         );
  NOR2_X1 U4122 ( .A1(n5565), .A2(n5459), .ZN(n3165) );
  AND2_X1 U4123 ( .A1(n4240), .A2(n4594), .ZN(n3166) );
  AND3_X1 U4124 ( .A1(n4265), .A2(n4282), .A3(n4264), .ZN(n5209) );
  INV_X1 U4125 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n4380) );
  INV_X1 U4126 ( .A(n4432), .ZN(n6298) );
  INV_X2 U4127 ( .A(n6688), .ZN(n6678) );
  INV_X2 U4128 ( .A(n3326), .ZN(n3345) );
  INV_X1 U4129 ( .A(n6092), .ZN(n4193) );
  AND2_X1 U4130 ( .A1(n4390), .A2(n4389), .ZN(n3167) );
  NAND2_X1 U4131 ( .A1(n3656), .A2(n3655), .ZN(n3168) );
  INV_X1 U4132 ( .A(n4042), .ZN(n3315) );
  INV_X1 U4133 ( .A(n3328), .ZN(n3329) );
  NAND2_X1 U4134 ( .A1(n4234), .A2(n3315), .ZN(n3316) );
  AND2_X1 U4135 ( .A1(n3337), .A2(n3336), .ZN(n3338) );
  INV_X1 U4136 ( .A(n4556), .ZN(n4028) );
  AOI22_X1 U4137 ( .A1(n3230), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3608), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3212) );
  NAND2_X1 U4138 ( .A1(n3354), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3360) );
  OR2_X1 U4139 ( .A1(n3485), .A2(n3484), .ZN(n4136) );
  NAND3_X1 U4140 ( .A1(n3361), .A2(n3360), .A3(n3359), .ZN(n3386) );
  INV_X1 U4141 ( .A(n5246), .ZN(n3324) );
  NAND2_X1 U4142 ( .A1(n3608), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3276) );
  OR2_X1 U4143 ( .A1(n3887), .A2(n3886), .ZN(n3902) );
  NOR2_X1 U4144 ( .A1(n3313), .A2(n6527), .ZN(n3559) );
  OR2_X1 U4145 ( .A1(n3507), .A2(n3506), .ZN(n4156) );
  AND4_X1 U4146 ( .A1(n3303), .A2(n3302), .A3(n3301), .A4(n3300), .ZN(n3304)
         );
  NAND2_X1 U4147 ( .A1(n4226), .A2(n4225), .ZN(n4230) );
  OR2_X1 U4148 ( .A1(n3866), .A2(n3865), .ZN(n3868) );
  INV_X1 U4149 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5495) );
  OR2_X1 U4150 ( .A1(n3495), .A2(n3494), .ZN(n4139) );
  INV_X1 U4151 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n6807) );
  INV_X1 U4152 ( .A(n4099), .ZN(n3348) );
  NOR2_X1 U4153 ( .A1(n5284), .A2(n5283), .ZN(n5285) );
  AND2_X1 U4154 ( .A1(n3641), .A2(n3640), .ZN(n5206) );
  AND2_X1 U4155 ( .A1(n4304), .A2(n4303), .ZN(n5301) );
  INV_X1 U4156 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3442) );
  XNOR2_X1 U4157 ( .A(n4474), .B(n5982), .ZN(n4534) );
  INV_X1 U4158 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n5983) );
  NAND2_X1 U4159 ( .A1(n4084), .A2(n4073), .ZN(n4074) );
  INV_X1 U4160 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4196) );
  AND2_X1 U4161 ( .A1(n5526), .A2(EBX_REG_31__SCAN_IN), .ZN(n5291) );
  NAND2_X1 U4162 ( .A1(n4089), .A2(n4088), .ZN(n4473) );
  OR2_X1 U4163 ( .A1(n5615), .A2(n5782), .ZN(n4390) );
  INV_X1 U4164 ( .A(n3786), .ZN(n5492) );
  INV_X1 U4165 ( .A(n4022), .ZN(n3971) );
  NAND2_X1 U4166 ( .A1(n3320), .A2(n4099), .ZN(n4192) );
  INV_X1 U4167 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5897) );
  INV_X1 U4168 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4502) );
  NOR2_X1 U4169 ( .A1(n4473), .A2(n4472), .ZN(n4612) );
  INV_X1 U4170 ( .A(n5122), .ZN(n5152) );
  AND2_X1 U4171 ( .A1(n4854), .A2(n5979), .ZN(n4921) );
  NOR2_X1 U4172 ( .A1(n4122), .A2(n4853), .ZN(n4854) );
  OR2_X1 U4173 ( .A1(n5988), .A2(n5987), .ZN(n6440) );
  NOR2_X1 U4174 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n6515) );
  INV_X1 U4175 ( .A(n6506), .ZN(n5200) );
  NAND2_X1 U4176 ( .A1(n3552), .A2(n3551), .ZN(n3553) );
  OR2_X1 U4177 ( .A1(n4720), .A2(n3345), .ZN(n6534) );
  OR2_X1 U4178 ( .A1(n4720), .A2(n3467), .ZN(n6567) );
  AND2_X1 U4179 ( .A1(n6261), .A2(n4700), .ZN(n4094) );
  INV_X2 U4180 ( .A(n6261), .ZN(n6253) );
  INV_X1 U4181 ( .A(n6288), .ZN(n6274) );
  NOR2_X1 U4182 ( .A1(n4650), .A2(n4649), .ZN(n4651) );
  INV_X1 U4183 ( .A(n6298), .ZN(n6332) );
  INV_X1 U4184 ( .A(n2974), .ZN(n5565) );
  AND2_X1 U4185 ( .A1(n3115), .A2(n5207), .ZN(n6164) );
  NAND2_X1 U4186 ( .A1(n6092), .A2(n4199), .ZN(n5775) );
  INV_X1 U4187 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4190) );
  NOR2_X1 U4188 ( .A1(n5828), .A2(n4368), .ZN(n5806) );
  OR2_X1 U4189 ( .A1(n5555), .A2(n6382), .ZN(n4402) );
  AND2_X1 U4190 ( .A1(n4297), .A2(n4296), .ZN(n5436) );
  AND2_X1 U4191 ( .A1(n4291), .A2(n4290), .ZN(n5467) );
  AND2_X1 U4192 ( .A1(n5936), .A2(n5935), .ZN(n6246) );
  NOR2_X1 U4193 ( .A1(n4922), .A2(n5987), .ZN(n5122) );
  OAI21_X1 U4194 ( .B1(n4921), .B2(n6428), .A(n6433), .ZN(n5125) );
  OAI21_X1 U4195 ( .B1(n4856), .B2(n4859), .A(n6036), .ZN(n4881) );
  OAI22_X1 U4196 ( .A1(n4899), .A2(n4895), .B1(n6527), .B2(n4896), .ZN(n6423)
         );
  INV_X1 U4197 ( .A(n6440), .ZN(n6848) );
  OAI211_X1 U4198 ( .C1(n6524), .C2(n5994), .A(n5993), .B(n6522), .ZN(n6024)
         );
  INV_X1 U4199 ( .A(n6511), .ZN(n6471) );
  AND2_X1 U4200 ( .A1(n5171), .A2(n5986), .ZN(n6506) );
  OAI211_X1 U4201 ( .C1(n5091), .C2(n6520), .A(n5090), .B(n6427), .ZN(n5114)
         );
  AND2_X1 U4202 ( .A1(n4915), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6465) );
  AND2_X1 U4203 ( .A1(n4122), .A2(n5966), .ZN(n5163) );
  INV_X1 U4204 ( .A(n6596), .ZN(n5001) );
  INV_X1 U4205 ( .A(n6553), .ZN(n6493) );
  INV_X1 U4206 ( .A(n6559), .ZN(n6494) );
  AND2_X1 U4207 ( .A1(n4751), .A2(n5986), .ZN(n5057) );
  INV_X1 U4208 ( .A(n6608), .ZN(n4663) );
  NOR2_X1 U4209 ( .A1(n4212), .A2(STATE_REG_0__SCAN_IN), .ZN(n4630) );
  INV_X1 U4210 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6610) );
  INV_X1 U4211 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6091) );
  NAND2_X1 U4212 ( .A1(n6250), .A2(n3313), .ZN(n5590) );
  INV_X1 U4213 ( .A(n6164), .ZN(n5214) );
  OR2_X1 U4214 ( .A1(n4830), .A2(n4730), .ZN(n6222) );
  NAND2_X1 U4215 ( .A1(n6307), .A2(n4093), .ZN(n6261) );
  OAI21_X1 U4216 ( .B1(n5435), .B2(n3119), .A(n5420), .ZN(n5700) );
  OAI21_X1 U4217 ( .B1(n5205), .B2(n3168), .A(n5593), .ZN(n5781) );
  AND2_X1 U4218 ( .A1(n4402), .A2(n4401), .ZN(n4403) );
  INV_X1 U4219 ( .A(n6395), .ZN(n6382) );
  INV_X1 U4220 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6409) );
  AOI22_X1 U4221 ( .A1(n5125), .A2(n5123), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5121), .ZN(n5156) );
  INV_X1 U4222 ( .A(n5154), .ZN(n4887) );
  OR2_X1 U4223 ( .A1(n4900), .A2(n5986), .ZN(n6853) );
  INV_X1 U4224 ( .A(n5985), .ZN(n6028) );
  INV_X1 U4225 ( .A(n6459), .ZN(n6074) );
  AOI22_X1 U4226 ( .A1(n4690), .A2(n4688), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6032), .ZN(n4725) );
  AOI22_X1 U4227 ( .A1(n5170), .A2(n5174), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5169), .ZN(n5204) );
  INV_X1 U4228 ( .A(n6542), .ZN(n6005) );
  INV_X1 U4229 ( .A(n6578), .ZN(n6027) );
  NAND2_X1 U4230 ( .A1(n5163), .A2(n5080), .ZN(n6575) );
  NAND2_X1 U4231 ( .A1(n5163), .A2(n4974), .ZN(n6596) );
  OR2_X1 U4232 ( .A1(n4809), .A2(n5986), .ZN(n5055) );
  AND2_X1 U4233 ( .A1(n5021), .A2(n5020), .ZN(n5060) );
  NAND2_X1 U4234 ( .A1(n4751), .A2(n5987), .ZN(n4952) );
  OR2_X1 U4235 ( .A1(n4659), .A2(n4658), .ZN(n5237) );
  NOR2_X1 U4236 ( .A1(n6688), .A2(n6089), .ZN(n6669) );
  INV_X1 U4237 ( .A(n4630), .ZN(n6082) );
  INV_X1 U4238 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6616) );
  INV_X1 U4239 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6647) );
  NAND2_X1 U4240 ( .A1(n6688), .A2(n6610), .ZN(n6659) );
  AOI22_X1 U4241 ( .A1(n3418), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3827), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3173) );
  AND2_X2 U4242 ( .A1(n4536), .A2(n4540), .ZN(n3264) );
  INV_X1 U4243 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3169) );
  AND2_X4 U4244 ( .A1(n4545), .A2(n4516), .ZN(n3608) );
  AND2_X2 U4245 ( .A1(n4516), .A2(n4542), .ZN(n3252) );
  AOI22_X1 U4246 ( .A1(n3608), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3252), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3171) );
  AOI22_X1 U4247 ( .A1(n3295), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3277), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3170) );
  AND2_X2 U4248 ( .A1(n4516), .A2(n4541), .ZN(n3247) );
  AOI22_X1 U4249 ( .A1(n3290), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n2975), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3175) );
  AND2_X2 U4250 ( .A1(n4517), .A2(n4541), .ZN(n3246) );
  AOI22_X1 U4251 ( .A1(n3230), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3608), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3181) );
  AOI22_X1 U4252 ( .A1(n3247), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3225), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3180) );
  AOI22_X1 U4253 ( .A1(n3295), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3246), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3179) );
  AOI22_X1 U4254 ( .A1(n3277), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3224), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3178) );
  INV_X2 U4255 ( .A(n3182), .ZN(n3975) );
  AOI22_X1 U4256 ( .A1(n3975), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3252), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3186) );
  AOI22_X1 U4257 ( .A1(n3264), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3290), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3185) );
  AOI22_X1 U4258 ( .A1(n4004), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3253), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3184) );
  INV_X1 U4259 ( .A(n4332), .ZN(n3555) );
  NAND2_X1 U4260 ( .A1(n3247), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3190) );
  NAND2_X1 U4261 ( .A1(n3608), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3189) );
  NAND2_X1 U4262 ( .A1(n3190), .A2(n3189), .ZN(n3194) );
  NAND2_X1 U4263 ( .A1(n3230), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3192)
         );
  NAND2_X1 U4264 ( .A1(n3225), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3191)
         );
  NAND2_X1 U4265 ( .A1(n3192), .A2(n3191), .ZN(n3193) );
  NOR2_X1 U4266 ( .A1(n3194), .A2(n3193), .ZN(n3210) );
  NAND2_X1 U4267 ( .A1(n3418), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3198)
         );
  NAND2_X1 U4268 ( .A1(n3264), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3197) );
  NAND2_X1 U4269 ( .A1(n3827), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3196)
         );
  NAND2_X1 U4270 ( .A1(n4004), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3202) );
  NAND2_X1 U4271 ( .A1(n3954), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3201) );
  NAND2_X1 U4272 ( .A1(n3252), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3200)
         );
  NAND2_X1 U4273 ( .A1(n3253), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3199) );
  NAND2_X1 U4274 ( .A1(n3246), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3206) );
  NAND2_X1 U4275 ( .A1(n3295), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3205) );
  NAND2_X1 U4276 ( .A1(n3277), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3204) );
  NAND2_X1 U4277 ( .A1(n3224), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3203)
         );
  INV_X1 U4278 ( .A(n3262), .ZN(n3211) );
  AOI22_X1 U4279 ( .A1(n3277), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n3224), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3214) );
  AOI22_X1 U4280 ( .A1(n3247), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3225), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3213) );
  NAND3_X1 U4281 ( .A1(n3214), .A2(n3213), .A3(n3212), .ZN(n3217) );
  AOI22_X1 U4282 ( .A1(n3295), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3246), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3215) );
  INV_X1 U4283 ( .A(n3215), .ZN(n3216) );
  NOR2_X1 U4284 ( .A1(n3217), .A2(n3216), .ZN(n3223) );
  AOI22_X1 U4285 ( .A1(n3418), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3827), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3221) );
  AOI22_X1 U4286 ( .A1(n3264), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3290), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3220) );
  AOI22_X1 U4287 ( .A1(n3975), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3252), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3219) );
  AOI22_X1 U4288 ( .A1(n4004), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3253), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3218) );
  NAND2_X1 U4289 ( .A1(n3223), .A2(n3222), .ZN(n3311) );
  INV_X2 U4290 ( .A(n3311), .ZN(n3320) );
  NAND2_X1 U4291 ( .A1(n3312), .A2(n3320), .ZN(n3308) );
  NAND2_X1 U4292 ( .A1(n3975), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3229) );
  NAND2_X1 U4293 ( .A1(n3608), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3228) );
  NAND2_X1 U4294 ( .A1(n3224), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3227)
         );
  NAND2_X1 U4295 ( .A1(n3880), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3226)
         );
  NAND2_X1 U4296 ( .A1(n3290), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3234) );
  INV_X2 U4297 ( .A(n3374), .ZN(n3285) );
  NAND2_X1 U4298 ( .A1(n3285), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3233)
         );
  NAND2_X1 U4299 ( .A1(n4006), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3232)
         );
  NAND2_X1 U4300 ( .A1(n3253), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3231) );
  NAND2_X1 U4301 ( .A1(n3418), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3238)
         );
  NAND2_X1 U4302 ( .A1(n4004), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3237) );
  NAND2_X1 U4303 ( .A1(n3264), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3236) );
  NAND2_X1 U4304 ( .A1(n3827), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3235)
         );
  NAND2_X1 U4305 ( .A1(n2970), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3242) );
  NAND2_X1 U4306 ( .A1(n3295), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3241) );
  NAND2_X1 U4307 ( .A1(n3247), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3240) );
  NAND2_X1 U4308 ( .A1(n3917), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3239) );
  INV_X2 U4309 ( .A(n4692), .ZN(n4337) );
  OAI21_X1 U4310 ( .B1(n3555), .B2(n3308), .A(n4337), .ZN(n3261) );
  NAND2_X2 U4311 ( .A1(n3467), .A2(n3262), .ZN(n3328) );
  AOI22_X1 U4312 ( .A1(n3285), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3608), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3251) );
  AOI22_X1 U4313 ( .A1(n3295), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n2970), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3250) );
  INV_X1 U4314 ( .A(n3247), .ZN(n3454) );
  AOI22_X1 U4315 ( .A1(n3247), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3880), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3249) );
  AOI22_X1 U4316 ( .A1(n3277), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3224), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3248) );
  NAND4_X1 U4317 ( .A1(n3251), .A2(n3250), .A3(n3249), .A4(n3248), .ZN(n3259)
         );
  AOI22_X1 U4318 ( .A1(n3418), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3827), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3257) );
  AOI22_X1 U4319 ( .A1(n3264), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3290), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3256) );
  BUF_X4 U4320 ( .A(n3252), .Z(n4006) );
  AOI22_X1 U4321 ( .A1(n4004), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3253), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3254) );
  NAND4_X1 U4322 ( .A1(n3257), .A2(n3256), .A3(n3255), .A4(n3254), .ZN(n3258)
         );
  OAI22_X1 U4323 ( .A1(n4700), .A2(n4692), .B1(n3351), .B2(n4099), .ZN(n3263)
         );
  NAND2_X1 U4324 ( .A1(n3418), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3268)
         );
  NAND2_X1 U4325 ( .A1(n3264), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3267) );
  NAND2_X1 U4326 ( .A1(n3827), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3266)
         );
  NAND2_X1 U4327 ( .A1(n3290), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3265) );
  NAND2_X1 U4328 ( .A1(n4004), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3272) );
  NAND2_X1 U4329 ( .A1(n3975), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3271) );
  NAND2_X1 U4330 ( .A1(n4006), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3270)
         );
  NAND2_X1 U4331 ( .A1(n3253), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3269) );
  NAND2_X1 U4332 ( .A1(n3285), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3275)
         );
  NAND2_X1 U4333 ( .A1(n3247), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3274) );
  NAND2_X1 U4334 ( .A1(n3880), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3273)
         );
  NAND2_X1 U4335 ( .A1(n3295), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3281) );
  NAND2_X1 U4336 ( .A1(n2970), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3280) );
  NAND2_X1 U4337 ( .A1(n3917), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3279) );
  NAND2_X1 U4338 ( .A1(n3224), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3278)
         );
  NAND4_X4 U4339 ( .A1(n3284), .A2(n2968), .A3(n3283), .A4(n3282), .ZN(n3326)
         );
  NAND2_X1 U4340 ( .A1(n4004), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3289) );
  NAND2_X1 U4341 ( .A1(n3264), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3288) );
  NAND2_X1 U4342 ( .A1(n3285), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3287)
         );
  NAND2_X1 U4343 ( .A1(n3253), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3286) );
  NAND2_X1 U4344 ( .A1(n3418), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3294)
         );
  NAND2_X1 U4345 ( .A1(n3975), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3293) );
  NAND2_X1 U4346 ( .A1(n3827), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3292)
         );
  NAND2_X1 U4347 ( .A1(n3959), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3291) );
  AND4_X2 U4348 ( .A1(n3294), .A2(n3293), .A3(n3292), .A4(n3291), .ZN(n3306)
         );
  NAND2_X1 U4349 ( .A1(n3295), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3299) );
  NAND2_X1 U4350 ( .A1(n2970), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3298) );
  NAND2_X1 U4351 ( .A1(n4006), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3297)
         );
  NAND2_X1 U4352 ( .A1(n3880), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3296)
         );
  NAND2_X1 U4353 ( .A1(n3608), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3303) );
  NAND2_X1 U4354 ( .A1(n3247), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3302) );
  NAND2_X1 U4355 ( .A1(n3917), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3301) );
  NAND2_X1 U4356 ( .A1(n3224), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3300)
         );
  NAND4_X4 U4357 ( .A1(n3307), .A2(n3306), .A3(n3305), .A4(n3304), .ZN(n5246)
         );
  INV_X1 U4358 ( .A(n3308), .ZN(n3309) );
  NAND2_X1 U4359 ( .A1(n3309), .A2(n3313), .ZN(n3340) );
  AND2_X1 U4360 ( .A1(n3328), .A2(n5246), .ZN(n3310) );
  XNOR2_X1 U4361 ( .A(STATE_REG_1__SCAN_IN), .B(STATE_REG_2__SCAN_IN), .ZN(
        n4212) );
  NAND2_X1 U4362 ( .A1(n3345), .A2(n4212), .ZN(n3344) );
  NAND2_X1 U4363 ( .A1(n3344), .A2(n3348), .ZN(n3314) );
  NAND2_X1 U4364 ( .A1(n3363), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3318) );
  NAND2_X1 U4365 ( .A1(n5334), .A2(n6603), .ZN(n4198) );
  MUX2_X1 U4366 ( .A(n4075), .B(n4198), .S(n6033), .Z(n3317) );
  NAND2_X1 U4367 ( .A1(n3318), .A2(n3317), .ZN(n3416) );
  NOR2_X2 U4368 ( .A1(n4105), .A2(n4337), .ZN(n3349) );
  NAND2_X1 U4369 ( .A1(n3724), .A2(n4483), .ZN(n3323) );
  INV_X1 U4370 ( .A(n5334), .ZN(n5975) );
  NOR2_X1 U4371 ( .A1(n5975), .A2(n6603), .ZN(n3322) );
  OR2_X1 U4372 ( .A1(n4192), .A2(n4259), .ZN(n4503) );
  NAND2_X2 U4373 ( .A1(n3321), .A2(n5246), .ZN(n4274) );
  NAND4_X1 U4374 ( .A1(n3323), .A2(n3322), .A3(n4503), .A4(n4274), .ZN(n3331)
         );
  INV_X1 U4375 ( .A(n3350), .ZN(n5345) );
  NAND2_X1 U4376 ( .A1(n4692), .A2(n5246), .ZN(n3327) );
  NAND3_X1 U4377 ( .A1(n4209), .A2(n5345), .A3(n3327), .ZN(n3330) );
  NAND2_X1 U4378 ( .A1(n3329), .A2(n4113), .ZN(n4206) );
  NAND2_X1 U4379 ( .A1(n3330), .A2(n4206), .ZN(n4336) );
  NOR2_X1 U4380 ( .A1(n3331), .A2(n4336), .ZN(n3339) );
  INV_X1 U4381 ( .A(n5345), .ZN(n5521) );
  NAND2_X1 U4382 ( .A1(n4210), .A2(n5521), .ZN(n4345) );
  NAND2_X1 U4383 ( .A1(n3328), .A2(n3333), .ZN(n3334) );
  NAND2_X1 U4384 ( .A1(n3334), .A2(n4105), .ZN(n3335) );
  OAI21_X1 U4385 ( .B1(n4338), .B2(n3335), .A(n3326), .ZN(n3337) );
  NAND3_X1 U4386 ( .A1(n3339), .A2(n4345), .A3(n3338), .ZN(n3414) );
  INV_X1 U4387 ( .A(n3340), .ZN(n3342) );
  NAND2_X1 U4388 ( .A1(n3342), .A2(n3341), .ZN(n4216) );
  INV_X1 U4389 ( .A(n4216), .ZN(n3343) );
  INV_X1 U4390 ( .A(n3344), .ZN(n3353) );
  INV_X1 U4391 ( .A(n4209), .ZN(n4334) );
  NAND3_X1 U4392 ( .A1(n3350), .A2(n3349), .A3(n3348), .ZN(n4090) );
  OR2_X2 U4393 ( .A1(n4090), .A2(n3352), .ZN(n4329) );
  OAI211_X1 U4394 ( .C1(n4076), .C2(n3353), .A(n4081), .B(n4329), .ZN(n3354)
         );
  INV_X1 U4395 ( .A(n3360), .ZN(n3357) );
  INV_X1 U4396 ( .A(n4198), .ZN(n3446) );
  NAND2_X1 U4397 ( .A1(n3446), .A2(n6467), .ZN(n3356) );
  INV_X1 U4398 ( .A(n4075), .ZN(n3445) );
  NAND2_X1 U4399 ( .A1(n3445), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3355) );
  NAND2_X1 U4400 ( .A1(n3356), .A2(n3355), .ZN(n3358) );
  NAND2_X1 U4401 ( .A1(n3357), .A2(n3163), .ZN(n3387) );
  NAND2_X1 U4402 ( .A1(n3385), .A2(n3387), .ZN(n3362) );
  NAND2_X1 U4403 ( .A1(n3363), .A2(n4556), .ZN(n3361) );
  INV_X1 U4404 ( .A(n3358), .ZN(n3359) );
  NAND3_X1 U4406 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), 
        .ZN(n3443) );
  NAND2_X1 U4407 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n3364) );
  NAND2_X1 U4408 ( .A1(n5087), .A2(n3364), .ZN(n3365) );
  NAND2_X1 U4409 ( .A1(n3443), .A2(n3365), .ZN(n4915) );
  OAI22_X1 U4410 ( .A1(n4198), .A2(n4915), .B1(n4075), .B2(n5087), .ZN(n3366)
         );
  AOI21_X1 U4411 ( .B1(n3441), .B2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n3366), 
        .ZN(n3367) );
  NAND2_X1 U4412 ( .A1(n3368), .A2(n3367), .ZN(n3369) );
  AOI22_X1 U4413 ( .A1(n3974), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3995), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3373) );
  AOI22_X1 U4414 ( .A1(n4002), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3994), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3372) );
  INV_X1 U4415 ( .A(n3975), .ZN(n3835) );
  INV_X2 U4416 ( .A(n3835), .ZN(n4003) );
  AOI22_X1 U4417 ( .A1(n4003), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4006), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3371) );
  AOI22_X1 U4418 ( .A1(n4004), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3931), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3370) );
  NAND4_X1 U4419 ( .A1(n3373), .A2(n3372), .A3(n3371), .A4(n3370), .ZN(n3380)
         );
  AOI22_X1 U4420 ( .A1(n3953), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n2970), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3378) );
  INV_X1 U4421 ( .A(n3285), .ZN(n3829) );
  AOI22_X1 U4422 ( .A1(n3980), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4005), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3377) );
  AOI22_X1 U4423 ( .A1(n3996), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3997), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3376) );
  INV_X1 U4424 ( .A(n3224), .ZN(n3479) );
  INV_X1 U4425 ( .A(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n6814) );
  AOI22_X1 U4426 ( .A1(n3881), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3455), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3375) );
  NAND4_X1 U4427 ( .A1(n3378), .A2(n3377), .A3(n3376), .A4(n3375), .ZN(n3379)
         );
  INV_X1 U4428 ( .A(n3381), .ZN(n4112) );
  AOI22_X1 U4429 ( .A1(n3382), .A2(n3381), .B1(n4056), .B2(
        INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3383) );
  INV_X1 U4430 ( .A(n3385), .ZN(n3389) );
  NAND2_X1 U4431 ( .A1(n3387), .A2(n3386), .ZN(n3388) );
  XNOR2_X1 U4432 ( .A(n3389), .B(n3388), .ZN(n4514) );
  NAND2_X1 U4433 ( .A1(n4514), .A2(n6603), .ZN(n3401) );
  AOI22_X1 U4434 ( .A1(n3974), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3995), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3393) );
  AOI22_X1 U4435 ( .A1(n4002), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3994), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3392) );
  AOI22_X1 U4436 ( .A1(n4003), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4006), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3391) );
  AOI22_X1 U4437 ( .A1(n4004), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3931), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3390) );
  NAND4_X1 U4438 ( .A1(n3393), .A2(n3392), .A3(n3391), .A4(n3390), .ZN(n3399)
         );
  AOI22_X1 U4439 ( .A1(n3953), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3806), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3397) );
  AOI22_X1 U4440 ( .A1(n3980), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4005), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3396) );
  AOI22_X1 U4441 ( .A1(n3996), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3997), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3395) );
  AOI22_X1 U4442 ( .A1(n3881), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3455), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3394) );
  NAND4_X1 U4443 ( .A1(n3397), .A2(n3396), .A3(n3395), .A4(n3394), .ZN(n3398)
         );
  AOI22_X1 U4444 ( .A1(n3974), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4002), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3405) );
  AOI22_X1 U4445 ( .A1(n4004), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3994), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3404) );
  AOI22_X1 U4446 ( .A1(n4003), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4006), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3403) );
  AOI22_X1 U4447 ( .A1(n3996), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3917), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3402) );
  NAND4_X1 U4448 ( .A1(n3405), .A2(n3404), .A3(n3403), .A4(n3402), .ZN(n3411)
         );
  AOI22_X1 U4449 ( .A1(n3980), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4005), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3409) );
  AOI22_X1 U4450 ( .A1(n3995), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3253), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3408) );
  AOI22_X1 U4451 ( .A1(n2970), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3997), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3407) );
  AOI22_X1 U4452 ( .A1(n3953), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3455), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3406) );
  NAND4_X1 U4453 ( .A1(n3409), .A2(n3408), .A3(n3407), .A4(n3406), .ZN(n3410)
         );
  NAND2_X1 U4454 ( .A1(n4056), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3412) );
  NAND2_X1 U4455 ( .A1(n3541), .A2(n3540), .ZN(n3566) );
  INV_X1 U4456 ( .A(n3414), .ZN(n3415) );
  XNOR2_X1 U4457 ( .A(n3416), .B(n3415), .ZN(n3558) );
  NAND2_X1 U4458 ( .A1(n3558), .A2(n6603), .ZN(n3432) );
  INV_X1 U4459 ( .A(n4169), .ZN(n3417) );
  AOI22_X1 U4460 ( .A1(n3974), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3994), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3422) );
  AOI22_X1 U4461 ( .A1(n4003), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4006), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3421) );
  AOI22_X1 U4462 ( .A1(n3953), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3996), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3420) );
  AOI22_X1 U4463 ( .A1(n3608), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3997), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3419) );
  NAND4_X1 U4464 ( .A1(n3422), .A2(n3421), .A3(n3420), .A4(n3419), .ZN(n3430)
         );
  AOI22_X1 U4465 ( .A1(n3285), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3806), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3428) );
  INV_X2 U4466 ( .A(n3423), .ZN(n4002) );
  AOI22_X1 U4467 ( .A1(n4002), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3995), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3427) );
  AOI22_X1 U4468 ( .A1(n3875), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3253), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3426) );
  AOI22_X1 U4469 ( .A1(n3881), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n3455), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3425) );
  NAND4_X1 U4470 ( .A1(n3428), .A2(n3427), .A3(n3426), .A4(n3425), .ZN(n3429)
         );
  MUX2_X1 U4471 ( .A(n4165), .B(n3431), .S(n4106), .Z(n3552) );
  NAND2_X1 U4472 ( .A1(n3432), .A2(n3552), .ZN(n3549) );
  INV_X1 U4473 ( .A(n4106), .ZN(n3435) );
  NAND2_X1 U4474 ( .A1(n4056), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3434) );
  AOI21_X1 U4475 ( .B1(n3320), .B2(n4169), .A(n6603), .ZN(n3433) );
  OAI211_X1 U4476 ( .C1(n3435), .C2(n5277), .A(n3434), .B(n3433), .ZN(n3550)
         );
  INV_X1 U4477 ( .A(n4165), .ZN(n3436) );
  AOI21_X1 U4478 ( .B1(n3549), .B2(n3550), .A(n3436), .ZN(n3542) );
  NAND2_X1 U4479 ( .A1(n3566), .A2(n3542), .ZN(n3439) );
  INV_X1 U4480 ( .A(n3540), .ZN(n3437) );
  BUF_X1 U4481 ( .A(n3440), .Z(n4474) );
  NAND2_X1 U4482 ( .A1(n3441), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3448) );
  INV_X1 U4483 ( .A(n3443), .ZN(n4747) );
  NAND2_X1 U4484 ( .A1(n3443), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3444) );
  NAND2_X1 U4485 ( .A1(n4721), .A2(n3444), .ZN(n6464) );
  AOI22_X1 U4486 ( .A1(n6464), .A2(n3446), .B1(n3445), .B2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3447) );
  NAND2_X1 U4487 ( .A1(n4534), .A2(n6603), .ZN(n3463) );
  AOI22_X1 U4488 ( .A1(n3974), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3995), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3453) );
  AOI22_X1 U4489 ( .A1(n4002), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3994), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3452) );
  AOI22_X1 U4490 ( .A1(n4003), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3916), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3451) );
  AOI22_X1 U4491 ( .A1(n3875), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3931), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3450) );
  NAND4_X1 U4492 ( .A1(n3453), .A2(n3452), .A3(n3451), .A4(n3450), .ZN(n3461)
         );
  AOI22_X1 U4493 ( .A1(n3953), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n2970), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3459) );
  AOI22_X1 U4494 ( .A1(n3980), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4005), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3458) );
  INV_X2 U4495 ( .A(n3454), .ZN(n3996) );
  AOI22_X1 U4496 ( .A1(n3996), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3997), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3457) );
  AOI22_X1 U4497 ( .A1(n3881), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3455), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3456) );
  NAND4_X1 U4498 ( .A1(n3459), .A2(n3458), .A3(n3457), .A4(n3456), .ZN(n3460)
         );
  AOI22_X1 U4499 ( .A1(n4073), .A2(n4124), .B1(n4056), .B2(
        INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3462) );
  INV_X1 U4500 ( .A(n3464), .ZN(n4683) );
  NAND2_X1 U4501 ( .A1(n3571), .A2(n4683), .ZN(n3466) );
  AND2_X2 U4502 ( .A1(n3466), .A2(n3527), .ZN(n4122) );
  NAND2_X1 U4503 ( .A1(n4122), .A2(n3711), .ZN(n3474) );
  INV_X1 U4504 ( .A(n3352), .ZN(n3468) );
  NAND2_X1 U4505 ( .A1(n3468), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3575) );
  INV_X1 U4506 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4554) );
  INV_X1 U4507 ( .A(n3508), .ZN(n3533) );
  NAND2_X1 U4508 ( .A1(n3079), .A2(n3572), .ZN(n3469) );
  NAND2_X1 U4509 ( .A1(n3533), .A2(n3469), .ZN(n6237) );
  AOI22_X1 U4510 ( .A1(n6237), .A2(n4022), .B1(n4024), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3471) );
  NAND2_X1 U4511 ( .A1(n4025), .A2(EAX_REG_3__SCAN_IN), .ZN(n3470) );
  OAI211_X1 U4512 ( .C1(n3575), .C2(n4554), .A(n3471), .B(n3470), .ZN(n3472)
         );
  INV_X1 U4513 ( .A(n3472), .ZN(n3473) );
  NAND2_X1 U4514 ( .A1(n3474), .A2(n3473), .ZN(n4600) );
  AOI22_X1 U4515 ( .A1(n3974), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3995), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3478) );
  AOI22_X1 U4516 ( .A1(INSTQUEUE_REG_6__4__SCAN_IN), .A2(n4003), .B1(n3994), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3477) );
  AOI22_X1 U4517 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n3806), .B1(n4005), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3476) );
  AOI22_X1 U4518 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n3980), .B1(n3916), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3475) );
  NAND4_X1 U4519 ( .A1(n3478), .A2(n3477), .A3(n3476), .A4(n3475), .ZN(n3485)
         );
  AOI22_X1 U4520 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n3875), .B1(n4002), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3483) );
  AOI22_X1 U4521 ( .A1(INSTQUEUE_REG_5__4__SCAN_IN), .A2(n3953), .B1(n3996), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3482) );
  AOI22_X1 U4522 ( .A1(n3931), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3997), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3481) );
  AOI22_X1 U4523 ( .A1(n3881), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3455), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3480) );
  NAND4_X1 U4524 ( .A1(n3483), .A2(n3482), .A3(n3481), .A4(n3480), .ZN(n3484)
         );
  AOI22_X1 U4525 ( .A1(n4073), .A2(n4136), .B1(n4056), .B2(
        INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3526) );
  AOI22_X1 U4526 ( .A1(n3974), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3995), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3489) );
  AOI22_X1 U4527 ( .A1(n4002), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3994), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3488) );
  AOI22_X1 U4528 ( .A1(n4003), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3916), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3487) );
  AOI22_X1 U4529 ( .A1(n3875), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3931), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3486) );
  NAND4_X1 U4530 ( .A1(n3489), .A2(n3488), .A3(n3487), .A4(n3486), .ZN(n3495)
         );
  AOI22_X1 U4531 ( .A1(n3953), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n2970), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3493) );
  AOI22_X1 U4532 ( .A1(n3980), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4005), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3492) );
  AOI22_X1 U4533 ( .A1(n3996), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3997), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3491) );
  AOI22_X1 U4534 ( .A1(n3881), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3455), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3490) );
  NAND4_X1 U4535 ( .A1(n3493), .A2(n3492), .A3(n3491), .A4(n3490), .ZN(n3494)
         );
  NAND2_X1 U4536 ( .A1(n4073), .A2(n4139), .ZN(n3497) );
  NAND2_X1 U4537 ( .A1(n4056), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3496) );
  NAND2_X1 U4538 ( .A1(n3497), .A2(n3496), .ZN(n3514) );
  AOI22_X1 U4539 ( .A1(n3995), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3994), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3501) );
  AOI22_X1 U4540 ( .A1(n4003), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4005), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3500) );
  AOI22_X1 U4541 ( .A1(n3806), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3996), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3499) );
  AOI22_X1 U4542 ( .A1(n3875), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3931), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3498) );
  NAND4_X1 U4543 ( .A1(n3501), .A2(n3500), .A3(n3499), .A4(n3498), .ZN(n3507)
         );
  AOI22_X1 U4544 ( .A1(n3974), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4002), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3505) );
  AOI22_X1 U4545 ( .A1(n3980), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3916), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3504) );
  AOI22_X1 U4546 ( .A1(n3953), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3997), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3503) );
  AOI22_X1 U4547 ( .A1(n3881), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3455), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3502) );
  NAND4_X1 U4548 ( .A1(n3505), .A2(n3504), .A3(n3503), .A4(n3502), .ZN(n3506)
         );
  AOI22_X1 U4549 ( .A1(n4073), .A2(n4156), .B1(n4056), .B2(
        INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3582) );
  NAND2_X1 U4550 ( .A1(n4146), .A2(n3711), .ZN(n3513) );
  XNOR2_X1 U4551 ( .A(n3588), .B(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n5511) );
  INV_X1 U4552 ( .A(EAX_REG_6__SCAN_IN), .ZN(n3510) );
  OAI21_X1 U4553 ( .B1(n6091), .B2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n6527), 
        .ZN(n3509) );
  OAI21_X1 U4554 ( .B1(n4018), .B2(n3510), .A(n3509), .ZN(n3511) );
  OAI21_X1 U4555 ( .B1(n3971), .B2(n5511), .A(n3511), .ZN(n3512) );
  OR2_X1 U4556 ( .A1(n3525), .A2(n3514), .ZN(n3515) );
  NAND2_X1 U4557 ( .A1(n3581), .A2(n3515), .ZN(n4142) );
  INV_X1 U4558 ( .A(n4142), .ZN(n3516) );
  INV_X1 U4559 ( .A(n3588), .ZN(n3519) );
  INV_X1 U4560 ( .A(n3517), .ZN(n3535) );
  INV_X1 U4561 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n6204) );
  NAND2_X1 U4562 ( .A1(n3535), .A2(n6204), .ZN(n3518) );
  NAND2_X1 U4563 ( .A1(n3519), .A2(n3518), .ZN(n6213) );
  NAND2_X1 U4564 ( .A1(n6213), .A2(n4022), .ZN(n3521) );
  NAND2_X1 U4565 ( .A1(n4024), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3520)
         );
  NAND2_X1 U4566 ( .A1(n3521), .A2(n3520), .ZN(n3522) );
  AOI21_X1 U4567 ( .B1(n4025), .B2(EAX_REG_5__SCAN_IN), .A(n3522), .ZN(n3523)
         );
  INV_X1 U4568 ( .A(n3525), .ZN(n3529) );
  NAND2_X1 U4569 ( .A1(n3527), .A2(n3526), .ZN(n3528) );
  NAND2_X1 U4570 ( .A1(n3529), .A2(n3528), .ZN(n4132) );
  INV_X1 U4571 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4475) );
  NAND2_X1 U4572 ( .A1(n6527), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3531)
         );
  NAND2_X1 U4573 ( .A1(n4025), .A2(EAX_REG_4__SCAN_IN), .ZN(n3530) );
  OAI211_X1 U4574 ( .C1(n3575), .C2(n4475), .A(n3531), .B(n3530), .ZN(n3536)
         );
  INV_X1 U4575 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3532) );
  NAND2_X1 U4576 ( .A1(n3533), .A2(n3532), .ZN(n3534) );
  NAND2_X1 U4577 ( .A1(n3535), .A2(n3534), .ZN(n6221) );
  MUX2_X1 U4578 ( .A(n3536), .B(n6221), .S(n4022), .Z(n3537) );
  INV_X1 U4579 ( .A(n3537), .ZN(n3538) );
  NAND2_X1 U4580 ( .A1(n3539), .A2(n3538), .ZN(n4727) );
  XNOR2_X1 U4581 ( .A(n3541), .B(n3540), .ZN(n3543) );
  INV_X1 U4582 ( .A(n3542), .ZN(n3567) );
  NAND2_X1 U4583 ( .A1(n2976), .A2(n3711), .ZN(n3548) );
  AOI22_X1 U4584 ( .A1(n4025), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n6527), .ZN(n3546) );
  INV_X1 U4585 ( .A(n3575), .ZN(n3544) );
  NAND2_X1 U4586 ( .A1(n3544), .A2(n4556), .ZN(n3545) );
  AND2_X1 U4587 ( .A1(n3546), .A2(n3545), .ZN(n3547) );
  NAND2_X1 U4588 ( .A1(n3548), .A2(n3547), .ZN(n4481) );
  INV_X1 U4589 ( .A(n3550), .ZN(n3551) );
  CLKBUF_X1 U4590 ( .A(n3555), .Z(n3556) );
  NAND2_X1 U4591 ( .A1(n5986), .A2(n3556), .ZN(n3557) );
  NAND2_X1 U4592 ( .A1(n3557), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4451) );
  NAND2_X1 U4593 ( .A1(n3559), .A2(EAX_REG_0__SCAN_IN), .ZN(n3561) );
  NAND2_X1 U4594 ( .A1(n6527), .A2(PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n3560)
         );
  OAI211_X1 U4595 ( .C1(n3575), .C2(n4502), .A(n3561), .B(n3560), .ZN(n3562)
         );
  AOI21_X1 U4596 ( .B1(n6519), .B2(n3711), .A(n3562), .ZN(n3563) );
  OR2_X1 U4597 ( .A1(n4451), .A2(n3563), .ZN(n4452) );
  INV_X1 U4598 ( .A(n3563), .ZN(n4453) );
  OR2_X1 U4599 ( .A1(n4453), .A2(n3971), .ZN(n3564) );
  NAND2_X1 U4600 ( .A1(n4452), .A2(n3564), .ZN(n4480) );
  NAND2_X1 U4601 ( .A1(n4481), .A2(n4480), .ZN(n4479) );
  INV_X1 U4602 ( .A(n3565), .ZN(n3570) );
  NAND2_X1 U4603 ( .A1(n3568), .A2(n3567), .ZN(n3569) );
  INV_X1 U4604 ( .A(n4024), .ZN(n3672) );
  OAI21_X1 U4605 ( .B1(PHYADDRPOINTER_REG_2__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_1__SCAN_IN), .A(n3572), .ZN(n6361) );
  AOI22_X1 U4606 ( .A1(n4022), .A2(n6361), .B1(n4024), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3574) );
  NAND2_X1 U4607 ( .A1(n4025), .A2(EAX_REG_2__SCAN_IN), .ZN(n3573) );
  OAI211_X1 U4608 ( .C1(n3575), .C2(n5338), .A(n3574), .B(n3573), .ZN(n4605)
         );
  NAND2_X1 U4609 ( .A1(n4604), .A2(n4605), .ZN(n3579) );
  INV_X1 U4610 ( .A(n4479), .ZN(n3577) );
  NAND2_X1 U4611 ( .A1(n3577), .A2(n3042), .ZN(n3578) );
  NAND2_X2 U4612 ( .A1(n3579), .A2(n3578), .ZN(n4599) );
  NAND4_X1 U4613 ( .A1(n3580), .A2(n4829), .A3(n4727), .A4(n4599), .ZN(n4791)
         );
  INV_X1 U4614 ( .A(n3581), .ZN(n3584) );
  INV_X1 U4615 ( .A(n3582), .ZN(n3583) );
  NAND2_X1 U4616 ( .A1(n4073), .A2(n4169), .ZN(n3586) );
  NAND2_X1 U4617 ( .A1(n4056), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3585) );
  NAND2_X1 U4618 ( .A1(n3586), .A2(n3585), .ZN(n3587) );
  XNOR2_X1 U4619 ( .A(n4167), .B(n3587), .ZN(n4154) );
  NAND2_X1 U4620 ( .A1(n4154), .A2(n3711), .ZN(n3593) );
  INV_X1 U4621 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3590) );
  OAI21_X1 U4622 ( .B1(PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n3017), .A(n3619), 
        .ZN(n6200) );
  NAND2_X1 U4623 ( .A1(n6200), .A2(n4022), .ZN(n3589) );
  OAI21_X1 U4624 ( .B1(n3590), .B2(n3672), .A(n3589), .ZN(n3591) );
  AOI21_X1 U4625 ( .B1(n4025), .B2(EAX_REG_7__SCAN_IN), .A(n3591), .ZN(n3592)
         );
  NAND2_X1 U4626 ( .A1(n3593), .A2(n3592), .ZN(n4964) );
  AOI22_X1 U4627 ( .A1(n3875), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3994), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3597) );
  AOI22_X1 U4628 ( .A1(n4003), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3980), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3596) );
  AOI22_X1 U4629 ( .A1(n3953), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3996), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3595) );
  AOI22_X1 U4630 ( .A1(n3881), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3455), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3594) );
  NAND4_X1 U4631 ( .A1(n3597), .A2(n3596), .A3(n3595), .A4(n3594), .ZN(n3603)
         );
  AOI22_X1 U4632 ( .A1(n3974), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n3995), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3601) );
  AOI22_X1 U4633 ( .A1(n4005), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3916), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3600) );
  AOI22_X1 U4634 ( .A1(n4002), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3931), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3599) );
  AOI22_X1 U4635 ( .A1(n2970), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3997), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3598) );
  NAND4_X1 U4636 ( .A1(n3601), .A2(n3600), .A3(n3599), .A4(n3598), .ZN(n3602)
         );
  OAI21_X1 U4637 ( .B1(n3603), .B2(n3602), .A(n3711), .ZN(n3607) );
  XNOR2_X1 U4638 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .B(n3619), .ZN(n6182) );
  INV_X1 U4639 ( .A(n6182), .ZN(n3604) );
  AOI22_X1 U4640 ( .A1(n4024), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .B1(n4022), 
        .B2(n3604), .ZN(n3606) );
  NAND2_X1 U4641 ( .A1(n4025), .A2(EAX_REG_8__SCAN_IN), .ZN(n3605) );
  AOI22_X1 U4642 ( .A1(n3974), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n3995), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3612) );
  AOI22_X1 U4643 ( .A1(n4002), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3994), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3611) );
  AOI22_X1 U4644 ( .A1(n3608), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3931), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3610) );
  AOI22_X1 U4645 ( .A1(n3953), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3455), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3609) );
  NAND4_X1 U4646 ( .A1(n3612), .A2(n3611), .A3(n3610), .A4(n3609), .ZN(n3618)
         );
  AOI22_X1 U4647 ( .A1(n3875), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3975), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3616) );
  AOI22_X1 U4648 ( .A1(n3980), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3916), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3615) );
  AOI22_X1 U4649 ( .A1(n3806), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3917), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3614) );
  AOI22_X1 U4650 ( .A1(n3996), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3997), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3613) );
  NAND4_X1 U4651 ( .A1(n3616), .A2(n3615), .A3(n3614), .A4(n3613), .ZN(n3617)
         );
  NOR2_X1 U4652 ( .A1(n3618), .A2(n3617), .ZN(n3624) );
  INV_X1 U4653 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3620) );
  XNOR2_X1 U4654 ( .A(n3625), .B(n3620), .ZN(n6171) );
  NAND2_X1 U4655 ( .A1(n6171), .A2(n4022), .ZN(n3622) );
  AOI22_X1 U4656 ( .A1(n4025), .A2(EAX_REG_9__SCAN_IN), .B1(n4024), .B2(
        PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3621) );
  OAI211_X1 U4657 ( .C1(n3624), .C2(n3623), .A(n3622), .B(n3621), .ZN(n5006)
         );
  AOI21_X1 U4658 ( .B1(n6810), .B2(n3626), .A(n3657), .ZN(n6163) );
  OR2_X1 U4659 ( .A1(n6163), .A2(n3971), .ZN(n3641) );
  AOI22_X1 U4660 ( .A1(n4003), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3980), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3630) );
  AOI22_X1 U4661 ( .A1(n3974), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3995), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3629) );
  AOI22_X1 U4662 ( .A1(n4005), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3917), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3628) );
  AOI22_X1 U4663 ( .A1(n4002), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3931), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3627) );
  NAND4_X1 U4664 ( .A1(n3630), .A2(n3629), .A3(n3628), .A4(n3627), .ZN(n3636)
         );
  AOI22_X1 U4665 ( .A1(n3875), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3994), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3634) );
  AOI22_X1 U4666 ( .A1(n3806), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3996), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3633) );
  AOI22_X1 U4667 ( .A1(n3916), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3997), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3632) );
  AOI22_X1 U4668 ( .A1(n3953), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3455), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3631) );
  NAND4_X1 U4669 ( .A1(n3634), .A2(n3633), .A3(n3632), .A4(n3631), .ZN(n3635)
         );
  OAI21_X1 U4670 ( .B1(n3636), .B2(n3635), .A(n3711), .ZN(n3639) );
  NAND2_X1 U4671 ( .A1(n4025), .A2(EAX_REG_10__SCAN_IN), .ZN(n3638) );
  NAND2_X1 U4672 ( .A1(n4024), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3637)
         );
  INV_X1 U4673 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n5774) );
  XNOR2_X1 U4674 ( .A(n3657), .B(n5774), .ZN(n5777) );
  OR2_X1 U4675 ( .A1(n5777), .A2(n3971), .ZN(n3656) );
  AOI22_X1 U4676 ( .A1(n3974), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3995), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3645) );
  AOI22_X1 U4677 ( .A1(n3875), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3975), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3644) );
  AOI22_X1 U4678 ( .A1(n4002), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3994), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3643) );
  AOI22_X1 U4679 ( .A1(n3916), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3455), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3642) );
  NAND4_X1 U4680 ( .A1(n3645), .A2(n3644), .A3(n3643), .A4(n3642), .ZN(n3651)
         );
  AOI22_X1 U4681 ( .A1(n3806), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3996), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3649) );
  AOI22_X1 U4682 ( .A1(n3980), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3931), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3648) );
  AOI22_X1 U4683 ( .A1(n3953), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3917), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3647) );
  AOI22_X1 U4684 ( .A1(n4005), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3997), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3646) );
  NAND4_X1 U4685 ( .A1(n3649), .A2(n3648), .A3(n3647), .A4(n3646), .ZN(n3650)
         );
  OAI21_X1 U4686 ( .B1(n3651), .B2(n3650), .A(n3711), .ZN(n3654) );
  NAND2_X1 U4687 ( .A1(n4025), .A2(EAX_REG_11__SCAN_IN), .ZN(n3653) );
  NAND2_X1 U4688 ( .A1(n4024), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3652)
         );
  NAND2_X1 U4689 ( .A1(n3657), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3671)
         );
  XNOR2_X1 U4690 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .B(n3671), .ZN(n6148)
         );
  AOI22_X1 U4691 ( .A1(n3959), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3916), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3661) );
  AOI22_X1 U4692 ( .A1(INSTQUEUE_REG_4__4__SCAN_IN), .A2(n3806), .B1(n3996), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3660) );
  AOI22_X1 U4693 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n4005), .B1(n3997), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3659) );
  AOI22_X1 U4694 ( .A1(n3953), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3455), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3658) );
  NAND4_X1 U4695 ( .A1(n3661), .A2(n3660), .A3(n3659), .A4(n3658), .ZN(n3667)
         );
  AOI22_X1 U4696 ( .A1(INSTQUEUE_REG_8__4__SCAN_IN), .A2(n3875), .B1(n4002), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3665) );
  AOI22_X1 U4697 ( .A1(n3974), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n3995), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3664) );
  AOI22_X1 U4698 ( .A1(n3980), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3881), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3663) );
  AOI22_X1 U4699 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n4003), .B1(n3931), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3662) );
  NAND4_X1 U4700 ( .A1(n3665), .A2(n3664), .A3(n3663), .A4(n3662), .ZN(n3666)
         );
  OR2_X1 U4701 ( .A1(n3667), .A2(n3666), .ZN(n3668) );
  AOI22_X1 U4702 ( .A1(n3711), .A2(n3668), .B1(n4024), .B2(
        PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3670) );
  NAND2_X1 U4703 ( .A1(n4025), .A2(EAX_REG_12__SCAN_IN), .ZN(n3669) );
  OAI211_X1 U4704 ( .C1(n6148), .C2(n3971), .A(n3670), .B(n3669), .ZN(n5591)
         );
  XNOR2_X1 U4705 ( .A(n3687), .B(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n6142)
         );
  NOR2_X1 U4706 ( .A1(n3672), .A2(n6140), .ZN(n3673) );
  AOI21_X1 U4707 ( .B1(n4025), .B2(EAX_REG_13__SCAN_IN), .A(n3673), .ZN(n3674)
         );
  OAI21_X1 U4708 ( .B1(n6142), .B2(n3971), .A(n3674), .ZN(n5574) );
  AOI22_X1 U4709 ( .A1(n3974), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3995), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3678) );
  AOI22_X1 U4710 ( .A1(n4002), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3994), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3677) );
  AOI22_X1 U4711 ( .A1(n4003), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3916), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3676) );
  AOI22_X1 U4712 ( .A1(n3875), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3931), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3675) );
  NAND4_X1 U4713 ( .A1(n3678), .A2(n3677), .A3(n3676), .A4(n3675), .ZN(n3684)
         );
  AOI22_X1 U4714 ( .A1(n3953), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3806), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3682) );
  AOI22_X1 U4715 ( .A1(n3980), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4005), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3681) );
  AOI22_X1 U4716 ( .A1(n3996), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n3997), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3680) );
  AOI22_X1 U4717 ( .A1(n3881), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3455), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3679) );
  NAND4_X1 U4718 ( .A1(n3682), .A2(n3681), .A3(n3680), .A4(n3679), .ZN(n3683)
         );
  OR2_X1 U4719 ( .A1(n3684), .A2(n3683), .ZN(n3685) );
  NAND2_X1 U4720 ( .A1(n5574), .A2(n5750), .ZN(n3686) );
  NAND2_X1 U4721 ( .A1(n5573), .A2(n3686), .ZN(n3722) );
  XNOR2_X1 U4722 ( .A(n3723), .B(n3082), .ZN(n6121) );
  AOI22_X1 U4723 ( .A1(n3974), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3995), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3691) );
  AOI22_X1 U4724 ( .A1(n3953), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3806), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3690) );
  AOI22_X1 U4725 ( .A1(n3994), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3916), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3689) );
  AOI22_X1 U4726 ( .A1(n3996), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3880), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3688) );
  NAND4_X1 U4727 ( .A1(n3691), .A2(n3690), .A3(n3689), .A4(n3688), .ZN(n3697)
         );
  AOI22_X1 U4728 ( .A1(n3875), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4002), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3695) );
  AOI22_X1 U4729 ( .A1(n3285), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4005), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3694) );
  AOI22_X1 U4730 ( .A1(n4003), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3931), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3693) );
  AOI22_X1 U4731 ( .A1(n3881), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3455), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3692) );
  NAND4_X1 U4732 ( .A1(n3695), .A2(n3694), .A3(n3693), .A4(n3692), .ZN(n3696)
         );
  OAI21_X1 U4733 ( .B1(n3697), .B2(n3696), .A(n3711), .ZN(n3700) );
  NAND2_X1 U4734 ( .A1(n4025), .A2(EAX_REG_15__SCAN_IN), .ZN(n3699) );
  NAND2_X1 U4735 ( .A1(n4024), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3698)
         );
  AND3_X1 U4736 ( .A1(n3700), .A2(n3699), .A3(n3698), .ZN(n3701) );
  OAI21_X1 U4737 ( .B1(n6121), .B2(n3971), .A(n3701), .ZN(n5576) );
  XNOR2_X1 U4738 ( .A(n3702), .B(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n6132)
         );
  NAND2_X1 U4739 ( .A1(n6132), .A2(n4022), .ZN(n3718) );
  AOI22_X1 U4740 ( .A1(n3974), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3995), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3706) );
  AOI22_X1 U4741 ( .A1(n4003), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3916), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3705) );
  AOI22_X1 U4742 ( .A1(n3806), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3996), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3704) );
  AOI22_X1 U4743 ( .A1(n3953), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3917), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3703) );
  NAND4_X1 U4744 ( .A1(n3706), .A2(n3705), .A3(n3704), .A4(n3703), .ZN(n3713)
         );
  AOI22_X1 U4745 ( .A1(n3285), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4005), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3710) );
  AOI22_X1 U4746 ( .A1(n4002), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3994), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3709) );
  AOI22_X1 U4747 ( .A1(n3875), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3931), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3708) );
  AOI22_X1 U4748 ( .A1(n3880), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3455), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3707) );
  NAND4_X1 U4749 ( .A1(n3710), .A2(n3709), .A3(n3708), .A4(n3707), .ZN(n3712)
         );
  OAI21_X1 U4750 ( .B1(n3713), .B2(n3712), .A(n3711), .ZN(n3716) );
  NAND2_X1 U4751 ( .A1(n4025), .A2(EAX_REG_14__SCAN_IN), .ZN(n3715) );
  NAND2_X1 U4752 ( .A1(n4024), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3714)
         );
  AND3_X1 U4753 ( .A1(n3716), .A2(n3715), .A3(n3714), .ZN(n3717) );
  NAND2_X1 U4754 ( .A1(n3718), .A2(n3717), .ZN(n5575) );
  OAI21_X1 U4755 ( .B1(n5750), .B2(n5574), .A(n5575), .ZN(n3719) );
  INV_X1 U4756 ( .A(n3719), .ZN(n3720) );
  AND2_X1 U4757 ( .A1(n5576), .A2(n3720), .ZN(n3721) );
  NAND2_X1 U4758 ( .A1(n3722), .A2(n3721), .ZN(n5563) );
  XNOR2_X1 U4759 ( .A(n3738), .B(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n6111)
         );
  INV_X1 U4760 ( .A(n6111), .ZN(n5735) );
  AOI22_X1 U4761 ( .A1(n4002), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3994), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3728) );
  AOI22_X1 U4762 ( .A1(n3875), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3285), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3727) );
  AOI22_X1 U4763 ( .A1(n3806), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3996), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3726) );
  AOI22_X1 U4764 ( .A1(n3881), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n3455), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3725) );
  NAND4_X1 U4765 ( .A1(n3728), .A2(n3727), .A3(n3726), .A4(n3725), .ZN(n3734)
         );
  AOI22_X1 U4766 ( .A1(n3974), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n3995), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3732) );
  AOI22_X1 U4767 ( .A1(n4005), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3916), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3731) );
  AOI22_X1 U4768 ( .A1(n4003), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3931), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3730) );
  AOI22_X1 U4769 ( .A1(n3953), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3880), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3729) );
  NAND4_X1 U4770 ( .A1(n3732), .A2(n3731), .A3(n3730), .A4(n3729), .ZN(n3733)
         );
  NOR2_X1 U4771 ( .A1(n3734), .A2(n3733), .ZN(n3736) );
  AOI22_X1 U4772 ( .A1(n4025), .A2(EAX_REG_16__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n4024), .ZN(n3735) );
  OAI21_X1 U4773 ( .B1(n3988), .B2(n3736), .A(n3735), .ZN(n3737) );
  AOI21_X1 U4774 ( .B1(n5735), .B2(n4022), .A(n3737), .ZN(n5564) );
  XNOR2_X1 U4775 ( .A(n3804), .B(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5706)
         );
  AOI22_X1 U4776 ( .A1(n4025), .A2(EAX_REG_20__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n6527), .ZN(n3753) );
  AOI22_X1 U4777 ( .A1(INSTQUEUE_REG_8__4__SCAN_IN), .A2(n4003), .B1(n3995), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3743) );
  AOI22_X1 U4778 ( .A1(n3875), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3806), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3742) );
  AOI22_X1 U4779 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n3285), .B1(n3994), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3741) );
  AOI22_X1 U4780 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n3953), .B1(n3916), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3740) );
  NAND4_X1 U4781 ( .A1(n3743), .A2(n3742), .A3(n3741), .A4(n3740), .ZN(n3751)
         );
  AOI22_X1 U4782 ( .A1(n3974), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n4005), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3749) );
  NAND2_X1 U4783 ( .A1(n4002), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3745)
         );
  NAND2_X1 U4784 ( .A1(n3917), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3744) );
  AND3_X1 U4785 ( .A1(n3745), .A2(n3971), .A3(n3744), .ZN(n3748) );
  AOI22_X1 U4786 ( .A1(n3996), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3931), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3747) );
  AOI22_X1 U4787 ( .A1(n3997), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3455), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3746) );
  NAND4_X1 U4788 ( .A1(n3749), .A2(n3748), .A3(n3747), .A4(n3746), .ZN(n3750)
         );
  NAND2_X1 U4789 ( .A1(n3988), .A2(n3971), .ZN(n3822) );
  OAI21_X1 U4790 ( .B1(n3751), .B2(n3750), .A(n3822), .ZN(n3752) );
  AOI22_X1 U4791 ( .A1(n5706), .A2(n4022), .B1(n3753), .B2(n3752), .ZN(n5446)
         );
  XNOR2_X1 U4792 ( .A(n3772), .B(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5720)
         );
  NAND2_X1 U4793 ( .A1(n5720), .A2(n4022), .ZN(n3769) );
  AOI22_X1 U4794 ( .A1(n4003), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3995), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3757) );
  AOI22_X1 U4795 ( .A1(n3953), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3959), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3756) );
  AOI22_X1 U4796 ( .A1(n3931), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3997), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3755) );
  AOI22_X1 U4797 ( .A1(n4005), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3455), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3754) );
  NAND4_X1 U4798 ( .A1(n3757), .A2(n3756), .A3(n3755), .A4(n3754), .ZN(n3765)
         );
  AOI22_X1 U4799 ( .A1(n3974), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3916), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3763) );
  AOI22_X1 U4800 ( .A1(n3980), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3806), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3762) );
  AOI22_X1 U4801 ( .A1(n3875), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3996), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3761) );
  NAND2_X1 U4802 ( .A1(n4002), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3759)
         );
  NAND2_X1 U4803 ( .A1(n3917), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3758) );
  AND3_X1 U4804 ( .A1(n3759), .A2(n3971), .A3(n3758), .ZN(n3760) );
  NAND4_X1 U4805 ( .A1(n3763), .A2(n3762), .A3(n3761), .A4(n3760), .ZN(n3764)
         );
  OAI21_X1 U4806 ( .B1(n3765), .B2(n3764), .A(n3822), .ZN(n3767) );
  AOI22_X1 U4807 ( .A1(n4025), .A2(EAX_REG_18__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n6527), .ZN(n3766) );
  NAND2_X1 U4808 ( .A1(n3767), .A2(n3766), .ZN(n3768) );
  NAND2_X1 U4809 ( .A1(n3769), .A2(n3768), .ZN(n5479) );
  NAND2_X1 U4810 ( .A1(n3770), .A2(n5495), .ZN(n3771) );
  NAND2_X1 U4811 ( .A1(n3772), .A2(n3771), .ZN(n5727) );
  AOI22_X1 U4812 ( .A1(n3974), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n4002), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3776) );
  AOI22_X1 U4813 ( .A1(n4005), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3916), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3775) );
  AOI22_X1 U4814 ( .A1(n3953), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3996), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3774) );
  AOI22_X1 U4815 ( .A1(n3881), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3455), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3773) );
  NAND4_X1 U4816 ( .A1(n3776), .A2(n3775), .A3(n3774), .A4(n3773), .ZN(n3782)
         );
  AOI22_X1 U4817 ( .A1(n4003), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3980), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3780) );
  AOI22_X1 U4818 ( .A1(n3995), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3994), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3779) );
  AOI22_X1 U4819 ( .A1(n3875), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3931), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3778) );
  AOI22_X1 U4820 ( .A1(n3806), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3997), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3777) );
  NAND4_X1 U4821 ( .A1(n3780), .A2(n3779), .A3(n3778), .A4(n3777), .ZN(n3781)
         );
  NOR2_X1 U4822 ( .A1(n3782), .A2(n3781), .ZN(n3784) );
  AOI22_X1 U4823 ( .A1(n4025), .A2(EAX_REG_17__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n6527), .ZN(n3783) );
  OAI21_X1 U4824 ( .B1(n3988), .B2(n3784), .A(n3783), .ZN(n3785) );
  MUX2_X1 U4825 ( .A(n5727), .B(n3785), .S(n3971), .Z(n3786) );
  AOI22_X1 U4826 ( .A1(n4002), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3995), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3790) );
  AOI22_X1 U4827 ( .A1(n3875), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3975), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3789) );
  AOI22_X1 U4828 ( .A1(n3953), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3996), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3788) );
  AOI22_X1 U4829 ( .A1(n3285), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3880), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3787) );
  NAND4_X1 U4830 ( .A1(n3790), .A2(n3789), .A3(n3788), .A4(n3787), .ZN(n3796)
         );
  AOI22_X1 U4831 ( .A1(n3806), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4005), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3794) );
  AOI22_X1 U4832 ( .A1(n3974), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3959), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3793) );
  AOI22_X1 U4833 ( .A1(n3916), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3931), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3792) );
  AOI22_X1 U4834 ( .A1(n3881), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n3455), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3791) );
  NAND4_X1 U4835 ( .A1(n3794), .A2(n3793), .A3(n3792), .A4(n3791), .ZN(n3795)
         );
  NOR2_X1 U4836 ( .A1(n3796), .A2(n3795), .ZN(n3798) );
  AOI22_X1 U4837 ( .A1(n4025), .A2(EAX_REG_19__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n6527), .ZN(n3797) );
  OAI21_X1 U4838 ( .B1(n3988), .B2(n3798), .A(n3797), .ZN(n3801) );
  NAND2_X1 U4839 ( .A1(n3799), .A2(n5469), .ZN(n3800) );
  NAND2_X1 U4840 ( .A1(n3804), .A2(n3800), .ZN(n5711) );
  MUX2_X1 U4841 ( .A(n3801), .B(n5711), .S(n4022), .Z(n5462) );
  INV_X1 U4842 ( .A(n5462), .ZN(n3802) );
  NOR2_X1 U4843 ( .A1(n5459), .A2(n3802), .ZN(n5445) );
  AND2_X1 U4844 ( .A1(n5446), .A2(n5445), .ZN(n3803) );
  INV_X1 U4845 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5702) );
  INV_X1 U4846 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n6811) );
  OAI21_X1 U4847 ( .B1(n3804), .B2(n5702), .A(n6811), .ZN(n3805) );
  NAND2_X1 U4848 ( .A1(n3805), .A2(n3820), .ZN(n5696) );
  INV_X1 U4849 ( .A(EAX_REG_21__SCAN_IN), .ZN(n6296) );
  AOI22_X1 U4850 ( .A1(n3875), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4002), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3810) );
  AOI22_X1 U4851 ( .A1(n4003), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3916), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3809) );
  AOI22_X1 U4852 ( .A1(n3806), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3881), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3808) );
  AOI22_X1 U4853 ( .A1(n3996), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3880), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3807) );
  NAND4_X1 U4854 ( .A1(n3810), .A2(n3809), .A3(n3808), .A4(n3807), .ZN(n3816)
         );
  AOI22_X1 U4855 ( .A1(n3285), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4005), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3814) );
  AOI22_X1 U4856 ( .A1(n3974), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3995), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3813) );
  AOI22_X1 U4857 ( .A1(n3959), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3931), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3812) );
  AOI22_X1 U4858 ( .A1(n3953), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3455), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3811) );
  NAND4_X1 U4859 ( .A1(n3814), .A2(n3813), .A3(n3812), .A4(n3811), .ZN(n3815)
         );
  OAI21_X1 U4860 ( .B1(n3816), .B2(n3815), .A(n4020), .ZN(n3818) );
  OAI21_X1 U4861 ( .B1(PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n6091), .A(n6527), 
        .ZN(n3817) );
  OAI211_X1 U4862 ( .C1(n4018), .C2(n6296), .A(n3818), .B(n3817), .ZN(n3819)
         );
  OAI21_X1 U4863 ( .B1(n5696), .B2(n3971), .A(n3819), .ZN(n5434) );
  NAND2_X1 U4864 ( .A1(n3820), .A2(n6807), .ZN(n3821) );
  NAND2_X1 U4865 ( .A1(n3845), .A2(n3821), .ZN(n5689) );
  INV_X1 U4866 ( .A(n3822), .ZN(n3842) );
  AOI22_X1 U4867 ( .A1(n4004), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3806), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3826) );
  AOI22_X1 U4868 ( .A1(n4005), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3994), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3825) );
  AOI22_X1 U4869 ( .A1(n3916), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3881), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3824) );
  AOI22_X1 U4870 ( .A1(n3974), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3931), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3823) );
  NAND4_X1 U4871 ( .A1(n3826), .A2(n3825), .A3(n3824), .A4(n3823), .ZN(n3839)
         );
  INV_X1 U4872 ( .A(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3828) );
  INV_X1 U4873 ( .A(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n5035) );
  OAI22_X1 U4874 ( .A1(n3829), .A2(n3828), .B1(n3424), .B2(n5035), .ZN(n3838)
         );
  INV_X1 U4875 ( .A(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3832) );
  AOI22_X1 U4876 ( .A1(n3953), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3997), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3831) );
  AOI21_X1 U4877 ( .B1(n4002), .B2(INSTQUEUE_REG_10__6__SCAN_IN), .A(n4022), 
        .ZN(n3830) );
  OAI211_X1 U4878 ( .C1(n3479), .C2(n3832), .A(n3831), .B(n3830), .ZN(n3837)
         );
  INV_X1 U4879 ( .A(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3834) );
  INV_X1 U4880 ( .A(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3833) );
  OAI22_X1 U4881 ( .A1(n3835), .A2(n3834), .B1(n3454), .B2(n3833), .ZN(n3836)
         );
  NOR4_X1 U4882 ( .A1(n3839), .A2(n3838), .A3(n3837), .A4(n3836), .ZN(n3841)
         );
  AOI22_X1 U4883 ( .A1(n4025), .A2(EAX_REG_22__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n6527), .ZN(n3840) );
  OAI21_X1 U4884 ( .B1(n3842), .B2(n3841), .A(n3840), .ZN(n3843) );
  OAI21_X1 U4885 ( .B1(n5689), .B2(n3971), .A(n3843), .ZN(n5421) );
  NAND2_X1 U4886 ( .A1(n3845), .A2(n3844), .ZN(n3846) );
  NAND2_X1 U4887 ( .A1(n3873), .A2(n3846), .ZN(n5414) );
  AOI22_X1 U4888 ( .A1(n3974), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3995), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3850) );
  AOI22_X1 U4889 ( .A1(n4002), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3994), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3849) );
  AOI22_X1 U4890 ( .A1(n3975), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3916), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3848) );
  AOI22_X1 U4891 ( .A1(n3875), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3931), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3847) );
  NAND4_X1 U4892 ( .A1(n3850), .A2(n3849), .A3(n3848), .A4(n3847), .ZN(n3856)
         );
  AOI22_X1 U4893 ( .A1(n3953), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3806), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3854) );
  AOI22_X1 U4894 ( .A1(n3980), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4005), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3853) );
  AOI22_X1 U4895 ( .A1(n3996), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3997), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3852) );
  AOI22_X1 U4896 ( .A1(n3881), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3455), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3851) );
  NAND4_X1 U4897 ( .A1(n3854), .A2(n3853), .A3(n3852), .A4(n3851), .ZN(n3855)
         );
  AOI22_X1 U4898 ( .A1(n3974), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3995), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3860) );
  AOI22_X1 U4899 ( .A1(n4002), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3994), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3859) );
  AOI22_X1 U4900 ( .A1(n3975), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3916), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3858) );
  AOI22_X1 U4901 ( .A1(n3875), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3931), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3857) );
  NAND4_X1 U4902 ( .A1(n3860), .A2(n3859), .A3(n3858), .A4(n3857), .ZN(n3866)
         );
  AOI22_X1 U4903 ( .A1(n3953), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3806), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3864) );
  AOI22_X1 U4904 ( .A1(n3285), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4005), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3863) );
  AOI22_X1 U4905 ( .A1(n3996), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3997), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3862) );
  AOI22_X1 U4906 ( .A1(n3881), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3455), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3861) );
  NAND4_X1 U4907 ( .A1(n3864), .A2(n3863), .A3(n3862), .A4(n3861), .ZN(n3865)
         );
  INV_X1 U4908 ( .A(n3901), .ZN(n3867) );
  OAI21_X1 U4909 ( .B1(n3869), .B2(n3868), .A(n3867), .ZN(n3871) );
  AOI22_X1 U4910 ( .A1(n4025), .A2(EAX_REG_23__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n6527), .ZN(n3870) );
  OAI21_X1 U4911 ( .B1(n3988), .B2(n3871), .A(n3870), .ZN(n3872) );
  MUX2_X1 U4912 ( .A(n5414), .B(n3872), .S(n3971), .Z(n4387) );
  INV_X1 U4913 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n6713) );
  NAND2_X1 U4914 ( .A1(n3873), .A2(n6713), .ZN(n3874) );
  NAND2_X1 U4915 ( .A1(n3907), .A2(n3874), .ZN(n5410) );
  AOI22_X1 U4916 ( .A1(n3974), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3995), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3879) );
  AOI22_X1 U4917 ( .A1(n4002), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3959), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3878) );
  AOI22_X1 U4918 ( .A1(n4003), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3916), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3877) );
  AOI22_X1 U4919 ( .A1(n3875), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3931), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3876) );
  NAND4_X1 U4920 ( .A1(n3879), .A2(n3878), .A3(n3877), .A4(n3876), .ZN(n3887)
         );
  AOI22_X1 U4921 ( .A1(n3953), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3806), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3885) );
  AOI22_X1 U4922 ( .A1(n3285), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4005), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3884) );
  AOI22_X1 U4923 ( .A1(n3996), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3880), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3883) );
  AOI22_X1 U4924 ( .A1(n3881), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3455), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3882) );
  NAND4_X1 U4925 ( .A1(n3885), .A2(n3884), .A3(n3883), .A4(n3882), .ZN(n3886)
         );
  XNOR2_X1 U4926 ( .A(n3901), .B(n3902), .ZN(n3889) );
  AOI22_X1 U4927 ( .A1(n4025), .A2(EAX_REG_24__SCAN_IN), .B1(n4024), .B2(
        PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n3888) );
  OAI21_X1 U4928 ( .B1(n3988), .B2(n3889), .A(n3888), .ZN(n3890) );
  AOI21_X1 U4929 ( .B1(n5410), .B2(n4022), .A(n3890), .ZN(n5297) );
  AOI22_X1 U4930 ( .A1(n3974), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3996), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3894) );
  AOI22_X1 U4931 ( .A1(n3875), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4003), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3893) );
  AOI22_X1 U4932 ( .A1(n4002), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3994), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3892) );
  AOI22_X1 U4933 ( .A1(n4005), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3916), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3891) );
  NAND4_X1 U4934 ( .A1(n3894), .A2(n3893), .A3(n3892), .A4(n3891), .ZN(n3900)
         );
  AOI22_X1 U4935 ( .A1(n3980), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3953), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3898) );
  AOI22_X1 U4936 ( .A1(n3995), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3881), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3897) );
  AOI22_X1 U4937 ( .A1(n3931), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3997), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3896) );
  AOI22_X1 U4938 ( .A1(n2970), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3455), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3895) );
  NAND4_X1 U4939 ( .A1(n3898), .A2(n3897), .A3(n3896), .A4(n3895), .ZN(n3899)
         );
  NOR2_X1 U4940 ( .A1(n3900), .A2(n3899), .ZN(n3910) );
  NAND2_X1 U4941 ( .A1(n3902), .A2(n3901), .ZN(n3911) );
  XNOR2_X1 U4942 ( .A(n3910), .B(n3911), .ZN(n3904) );
  AOI22_X1 U4943 ( .A1(n4025), .A2(EAX_REG_25__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n6527), .ZN(n3903) );
  OAI21_X1 U4944 ( .B1(n3988), .B2(n3904), .A(n3903), .ZN(n3909) );
  INV_X1 U4945 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n3906) );
  NAND2_X1 U4946 ( .A1(n3907), .A2(n3906), .ZN(n3908) );
  NAND2_X1 U4947 ( .A1(n3944), .A2(n3908), .ZN(n5682) );
  MUX2_X1 U4948 ( .A(n3909), .B(n5682), .S(n4022), .Z(n5395) );
  XOR2_X1 U4949 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .B(n3944), .Z(n5674) );
  INV_X1 U4950 ( .A(EAX_REG_26__SCAN_IN), .ZN(n3927) );
  OR2_X1 U4951 ( .A1(n3911), .A2(n3910), .ZN(n3929) );
  AOI22_X1 U4952 ( .A1(n3974), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n4002), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3915) );
  AOI22_X1 U4953 ( .A1(n3980), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3806), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3914) );
  AOI22_X1 U4954 ( .A1(n4003), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3931), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3913) );
  AOI22_X1 U4955 ( .A1(n3953), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3455), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3912) );
  NAND4_X1 U4956 ( .A1(n3915), .A2(n3914), .A3(n3913), .A4(n3912), .ZN(n3923)
         );
  AOI22_X1 U4957 ( .A1(n3995), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3994), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3921) );
  AOI22_X1 U4958 ( .A1(n3875), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3916), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3920) );
  AOI22_X1 U4959 ( .A1(n3996), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3917), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3919) );
  AOI22_X1 U4960 ( .A1(n4005), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3997), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3918) );
  NAND4_X1 U4961 ( .A1(n3921), .A2(n3920), .A3(n3919), .A4(n3918), .ZN(n3922)
         );
  NOR2_X1 U4962 ( .A1(n3923), .A2(n3922), .ZN(n3930) );
  XOR2_X1 U4963 ( .A(n3929), .B(n3930), .Z(n3924) );
  NAND2_X1 U4964 ( .A1(n3924), .A2(n4020), .ZN(n3926) );
  OAI21_X1 U4965 ( .B1(n6091), .B2(PHYADDRPOINTER_REG_26__SCAN_IN), .A(n6527), 
        .ZN(n3925) );
  OAI211_X1 U4966 ( .C1(n4018), .C2(n3927), .A(n3926), .B(n3925), .ZN(n3928)
         );
  OAI21_X1 U4967 ( .B1(n5674), .B2(n3971), .A(n3928), .ZN(n5384) );
  NOR2_X1 U4968 ( .A1(n3930), .A2(n3929), .ZN(n3952) );
  AOI22_X1 U4969 ( .A1(n3974), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3995), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3935) );
  AOI22_X1 U4970 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n4002), .B1(n3994), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3934) );
  AOI22_X1 U4971 ( .A1(n3975), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4006), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3933) );
  AOI22_X1 U4972 ( .A1(n3875), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3931), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3932) );
  NAND4_X1 U4973 ( .A1(n3935), .A2(n3934), .A3(n3933), .A4(n3932), .ZN(n3941)
         );
  AOI22_X1 U4974 ( .A1(INSTQUEUE_REG_8__4__SCAN_IN), .A2(n3953), .B1(n3806), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3939) );
  AOI22_X1 U4975 ( .A1(INSTQUEUE_REG_14__4__SCAN_IN), .A2(n3285), .B1(n4005), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3938) );
  AOI22_X1 U4976 ( .A1(INSTQUEUE_REG_5__4__SCAN_IN), .A2(n3996), .B1(n3997), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3937) );
  AOI22_X1 U4977 ( .A1(n3881), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3455), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3936) );
  NAND4_X1 U4978 ( .A1(n3939), .A2(n3938), .A3(n3937), .A4(n3936), .ZN(n3940)
         );
  XNOR2_X1 U4979 ( .A(n3952), .B(n3951), .ZN(n3943) );
  AOI22_X1 U4980 ( .A1(n4025), .A2(EAX_REG_27__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n6527), .ZN(n3942) );
  OAI21_X1 U4981 ( .B1(n3943), .B2(n3988), .A(n3942), .ZN(n3950) );
  INV_X1 U4982 ( .A(n3944), .ZN(n3945) );
  INV_X1 U4983 ( .A(n3946), .ZN(n3948) );
  INV_X1 U4984 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n3947) );
  NAND2_X1 U4985 ( .A1(n3948), .A2(n3947), .ZN(n3949) );
  NAND2_X1 U4986 ( .A1(n3990), .A2(n3949), .ZN(n5658) );
  MUX2_X1 U4987 ( .A(n3950), .B(n5658), .S(n4022), .Z(n5371) );
  XOR2_X1 U4988 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .B(n3990), .Z(n5654) );
  INV_X1 U4989 ( .A(EAX_REG_28__SCAN_IN), .ZN(n3969) );
  NAND2_X1 U4990 ( .A1(n3952), .A2(n3951), .ZN(n3972) );
  AOI22_X1 U4991 ( .A1(n3875), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3995), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3958) );
  AOI22_X1 U4992 ( .A1(n3953), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3996), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3957) );
  AOI22_X1 U4993 ( .A1(n3954), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3931), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3956) );
  AOI22_X1 U4994 ( .A1(n3285), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3997), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3955) );
  NAND4_X1 U4995 ( .A1(n3958), .A2(n3957), .A3(n3956), .A4(n3955), .ZN(n3965)
         );
  AOI22_X1 U4996 ( .A1(n3974), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n4002), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3963) );
  AOI22_X1 U4997 ( .A1(n2970), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4005), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3962) );
  AOI22_X1 U4998 ( .A1(n3959), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4006), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3961) );
  AOI22_X1 U4999 ( .A1(n3881), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3455), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3960) );
  NAND4_X1 U5000 ( .A1(n3963), .A2(n3962), .A3(n3961), .A4(n3960), .ZN(n3964)
         );
  NOR2_X1 U5001 ( .A1(n3965), .A2(n3964), .ZN(n3973) );
  XOR2_X1 U5002 ( .A(n3972), .B(n3973), .Z(n3966) );
  NAND2_X1 U5003 ( .A1(n3966), .A2(n4020), .ZN(n3968) );
  OAI21_X1 U5004 ( .B1(n6091), .B2(PHYADDRPOINTER_REG_28__SCAN_IN), .A(n6527), 
        .ZN(n3967) );
  OAI211_X1 U5005 ( .C1(n4018), .C2(n3969), .A(n3968), .B(n3967), .ZN(n3970)
         );
  OAI21_X1 U5006 ( .B1(n5654), .B2(n3971), .A(n3970), .ZN(n5361) );
  NOR2_X1 U5007 ( .A1(n3973), .A2(n3972), .ZN(n4014) );
  AOI22_X1 U5008 ( .A1(n3974), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3995), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3979) );
  AOI22_X1 U5009 ( .A1(n4002), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3994), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3978) );
  AOI22_X1 U5010 ( .A1(n3975), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4006), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3977) );
  AOI22_X1 U5011 ( .A1(n4004), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3931), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3976) );
  NAND4_X1 U5012 ( .A1(n3979), .A2(n3978), .A3(n3977), .A4(n3976), .ZN(n3986)
         );
  AOI22_X1 U5013 ( .A1(n3953), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n2970), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3984) );
  AOI22_X1 U5014 ( .A1(n3980), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4005), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3983) );
  AOI22_X1 U5015 ( .A1(n3996), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3997), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3982) );
  AOI22_X1 U5016 ( .A1(n3881), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3455), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3981) );
  NAND4_X1 U5017 ( .A1(n3984), .A2(n3983), .A3(n3982), .A4(n3981), .ZN(n3985)
         );
  OR2_X1 U5018 ( .A1(n3986), .A2(n3985), .ZN(n4013) );
  XNOR2_X1 U5019 ( .A(n4014), .B(n4013), .ZN(n3989) );
  AOI22_X1 U5020 ( .A1(n4025), .A2(EAX_REG_29__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n6527), .ZN(n3987) );
  OAI21_X1 U5021 ( .B1(n3989), .B2(n3988), .A(n3987), .ZN(n3993) );
  INV_X1 U5022 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n3991) );
  NAND2_X1 U5023 ( .A1(n3077), .A2(n3991), .ZN(n3992) );
  NAND2_X1 U5024 ( .A1(n4195), .A2(n3992), .ZN(n5637) );
  MUX2_X1 U5025 ( .A(n3993), .B(n5637), .S(n4022), .Z(n5350) );
  AOI22_X1 U5026 ( .A1(n3995), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3994), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4001) );
  AOI22_X1 U5027 ( .A1(n2970), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3996), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4000) );
  AOI22_X1 U5028 ( .A1(n3931), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3997), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3999) );
  AOI22_X1 U5029 ( .A1(n3881), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3455), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3998) );
  NAND4_X1 U5030 ( .A1(n4001), .A2(n4000), .A3(n3999), .A4(n3998), .ZN(n4012)
         );
  AOI22_X1 U5031 ( .A1(n3974), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n4002), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n4010) );
  AOI22_X1 U5032 ( .A1(n4004), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4003), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n4009) );
  AOI22_X1 U5033 ( .A1(n3953), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4005), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n4008) );
  AOI22_X1 U5034 ( .A1(n3285), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4006), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4007) );
  NAND4_X1 U5035 ( .A1(n4010), .A2(n4009), .A3(n4008), .A4(n4007), .ZN(n4011)
         );
  NOR2_X1 U5036 ( .A1(n4012), .A2(n4011), .ZN(n4016) );
  NAND2_X1 U5037 ( .A1(n4014), .A2(n4013), .ZN(n4015) );
  XOR2_X1 U5038 ( .A(n4016), .B(n4015), .Z(n4021) );
  INV_X1 U5039 ( .A(EAX_REG_30__SCAN_IN), .ZN(n4017) );
  INV_X1 U5040 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5323) );
  OAI22_X1 U5041 ( .A1(n4018), .A2(n4017), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5323), .ZN(n4019) );
  AOI21_X1 U5042 ( .B1(n4021), .B2(n4020), .A(n4019), .ZN(n4023) );
  XNOR2_X1 U5043 ( .A(n4195), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5326)
         );
  MUX2_X1 U5044 ( .A(n4023), .B(n5326), .S(n4022), .Z(n5233) );
  AOI22_X1 U5045 ( .A1(n4025), .A2(EAX_REG_31__SCAN_IN), .B1(n4024), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4026) );
  NAND2_X1 U5046 ( .A1(n5983), .A2(n4556), .ZN(n4030) );
  NAND2_X1 U5047 ( .A1(n4028), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4029) );
  NAND2_X1 U5048 ( .A1(n4030), .A2(n4029), .ZN(n4038) );
  NAND2_X1 U5049 ( .A1(n6033), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4041) );
  NAND2_X1 U5050 ( .A1(n4031), .A2(n4030), .ZN(n4055) );
  NAND2_X1 U5051 ( .A1(n5087), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4034) );
  NAND2_X1 U5052 ( .A1(n2972), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4032) );
  NAND2_X1 U5053 ( .A1(n4034), .A2(n4032), .ZN(n4054) );
  INV_X1 U5054 ( .A(n4054), .ZN(n4033) );
  NAND2_X1 U5055 ( .A1(n4055), .A2(n4033), .ZN(n4035) );
  NAND2_X1 U5056 ( .A1(n4035), .A2(n4034), .ZN(n4064) );
  MUX2_X1 U5057 ( .A(n3442), .B(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .S(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n4063) );
  NAND2_X1 U5058 ( .A1(n4084), .A2(n4070), .ZN(n4072) );
  INV_X1 U5059 ( .A(n4041), .ZN(n4037) );
  XNOR2_X1 U5060 ( .A(n4038), .B(n4037), .ZN(n4082) );
  NAND2_X1 U5061 ( .A1(n4073), .A2(n4339), .ZN(n4039) );
  NAND2_X1 U5062 ( .A1(n4039), .A2(n4099), .ZN(n4050) );
  NAND2_X1 U5063 ( .A1(n4502), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4040) );
  AND2_X1 U5064 ( .A1(n4041), .A2(n4040), .ZN(n4046) );
  OAI21_X1 U5065 ( .B1(n4042), .B2(n3348), .A(n4046), .ZN(n4043) );
  NAND2_X1 U5066 ( .A1(n4043), .A2(n5246), .ZN(n4045) );
  NAND2_X1 U5067 ( .A1(n3345), .A2(n4099), .ZN(n4044) );
  NAND2_X1 U5068 ( .A1(n4045), .A2(n4057), .ZN(n4049) );
  NAND2_X1 U5069 ( .A1(n4073), .A2(n4046), .ZN(n4047) );
  NAND2_X1 U5070 ( .A1(n4047), .A2(n4053), .ZN(n4048) );
  OAI211_X1 U5071 ( .C1(n4050), .C2(n4082), .A(n4049), .B(n4048), .ZN(n4052)
         );
  NAND3_X1 U5072 ( .A1(n4050), .A2(n4082), .A3(STATE2_REG_0__SCAN_IN), .ZN(
        n4051) );
  OAI211_X1 U5073 ( .C1(n4082), .C2(n4053), .A(n4052), .B(n4051), .ZN(n4061)
         );
  XNOR2_X1 U5074 ( .A(n4055), .B(n4054), .ZN(n4083) );
  INV_X1 U5075 ( .A(n4056), .ZN(n4069) );
  NAND2_X1 U5076 ( .A1(n4073), .A2(n4083), .ZN(n4058) );
  OAI211_X1 U5077 ( .C1(n4083), .C2(n4069), .A(n4058), .B(n4057), .ZN(n4060)
         );
  NOR2_X1 U5078 ( .A1(n4058), .A2(n4057), .ZN(n4059) );
  NAND3_X1 U5079 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n4062), .A3(n4475), .ZN(n4068) );
  NOR2_X1 U5080 ( .A1(n4064), .A2(n4063), .ZN(n4065) );
  NOR2_X1 U5081 ( .A1(n4066), .A2(n4065), .ZN(n4067) );
  NAND2_X1 U5082 ( .A1(n4068), .A2(n4067), .ZN(n4087) );
  NAND2_X1 U5083 ( .A1(n3326), .A2(n6793), .ZN(n4077) );
  NAND2_X1 U5084 ( .A1(n4518), .A2(n4709), .ZN(n4079) );
  NAND2_X1 U5085 ( .A1(n4080), .A2(n4079), .ZN(n4208) );
  OR2_X1 U5086 ( .A1(n4509), .A2(n4537), .ZN(n4089) );
  INV_X1 U5087 ( .A(n4081), .ZN(n4572) );
  NAND2_X1 U5088 ( .A1(n4083), .A2(n4082), .ZN(n4086) );
  INV_X1 U5089 ( .A(n4084), .ZN(n4085) );
  OAI21_X1 U5090 ( .B1(n4087), .B2(n4086), .A(n4085), .ZN(n4427) );
  NOR2_X1 U5091 ( .A1(READY_N), .A2(n4427), .ZN(n4213) );
  NAND2_X1 U5092 ( .A1(n4572), .A2(n4213), .ZN(n4088) );
  NAND3_X1 U5093 ( .A1(n4700), .A2(n3320), .A3(n4091), .ZN(n4482) );
  NOR2_X1 U5094 ( .A1(n4090), .A2(n4482), .ZN(n4092) );
  AOI22_X1 U5095 ( .A1(n6251), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n6253), .ZN(n4095) );
  NAND2_X1 U5096 ( .A1(n4096), .A2(n4095), .ZN(U2860) );
  NAND2_X1 U5097 ( .A1(n4685), .A2(n4153), .ZN(n4104) );
  NAND2_X1 U5098 ( .A1(n4097), .A2(n4106), .ZN(n4111) );
  OAI21_X1 U5099 ( .B1(n4106), .B2(n4097), .A(n4111), .ZN(n4101) );
  INV_X1 U5100 ( .A(n4113), .ZN(n4098) );
  INV_X1 U5101 ( .A(n4340), .ZN(n4100) );
  OAI211_X1 U5102 ( .C1(n4101), .C2(n4098), .A(n4100), .B(n4099), .ZN(n4102)
         );
  INV_X1 U5103 ( .A(n4102), .ZN(n4103) );
  NAND2_X1 U5104 ( .A1(n4709), .A2(n4105), .ZN(n4114) );
  OAI21_X1 U5105 ( .B1(n4098), .B2(n4106), .A(n4114), .ZN(n4107) );
  INV_X1 U5106 ( .A(n4107), .ZN(n4108) );
  XNOR2_X1 U5107 ( .A(n4459), .B(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4493)
         );
  NAND2_X1 U5108 ( .A1(n4494), .A2(n4493), .ZN(n4492) );
  INV_X1 U5109 ( .A(n4459), .ZN(n4109) );
  NAND2_X1 U5110 ( .A1(n4109), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4110)
         );
  AND2_X1 U5111 ( .A1(n4492), .A2(n4110), .ZN(n6356) );
  NAND2_X1 U5112 ( .A1(n4111), .A2(n4112), .ZN(n4123) );
  OAI21_X1 U5113 ( .B1(n4112), .B2(n4111), .A(n4123), .ZN(n4116) );
  INV_X1 U5114 ( .A(n4114), .ZN(n4115) );
  AOI21_X1 U5115 ( .B1(n4116), .B2(n5273), .A(n4115), .ZN(n4117) );
  NAND2_X1 U5116 ( .A1(n4118), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6353)
         );
  NAND2_X1 U5117 ( .A1(n6356), .A2(n6353), .ZN(n4121) );
  INV_X1 U5118 ( .A(n4118), .ZN(n4120) );
  INV_X1 U5119 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4119) );
  NAND2_X1 U5120 ( .A1(n4120), .A2(n4119), .ZN(n6354) );
  NAND2_X1 U5121 ( .A1(n4122), .A2(n4153), .ZN(n4126) );
  NAND2_X1 U5122 ( .A1(n4123), .A2(n4124), .ZN(n4138) );
  OAI211_X1 U5123 ( .C1(n4124), .C2(n4123), .A(n4138), .B(n5273), .ZN(n4125)
         );
  INV_X1 U5124 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4592) );
  NAND2_X1 U5125 ( .A1(n4589), .A2(n4588), .ZN(n4129) );
  NAND2_X1 U5126 ( .A1(n4127), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4128)
         );
  NAND2_X1 U5127 ( .A1(n4129), .A2(n4128), .ZN(n4637) );
  XNOR2_X1 U5128 ( .A(n4138), .B(n4136), .ZN(n4130) );
  NAND2_X1 U5129 ( .A1(n4130), .A2(n5273), .ZN(n4131) );
  OAI21_X1 U5130 ( .B1(n4132), .B2(n4164), .A(n4131), .ZN(n4133) );
  INV_X1 U5131 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4242) );
  XNOR2_X1 U5132 ( .A(n4133), .B(n4242), .ZN(n4636) );
  NAND2_X1 U5133 ( .A1(n4637), .A2(n4636), .ZN(n4135) );
  NAND2_X1 U5134 ( .A1(n4133), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4134)
         );
  NAND2_X1 U5135 ( .A1(n4135), .A2(n4134), .ZN(n4734) );
  INV_X1 U5136 ( .A(n4136), .ZN(n4137) );
  NOR2_X1 U5137 ( .A1(n4138), .A2(n4137), .ZN(n4140) );
  NAND2_X1 U5138 ( .A1(n4140), .A2(n4139), .ZN(n4155) );
  OAI211_X1 U5139 ( .C1(n4140), .C2(n4139), .A(n4155), .B(n5273), .ZN(n4141)
         );
  INV_X1 U5140 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4740) );
  XNOR2_X1 U5141 ( .A(n4143), .B(n4740), .ZN(n4735) );
  NAND2_X1 U5142 ( .A1(n4734), .A2(n4735), .ZN(n4145) );
  NAND2_X1 U5143 ( .A1(n4143), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4144)
         );
  NAND2_X1 U5144 ( .A1(n4145), .A2(n4144), .ZN(n4845) );
  NAND3_X1 U5145 ( .A1(n4167), .A2(n4146), .A3(n4153), .ZN(n4149) );
  XNOR2_X1 U5146 ( .A(n4155), .B(n4156), .ZN(n4147) );
  NAND2_X1 U5147 ( .A1(n4147), .A2(n5273), .ZN(n4148) );
  NAND2_X1 U5148 ( .A1(n4149), .A2(n4148), .ZN(n4150) );
  INV_X1 U5149 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n6780) );
  NAND2_X1 U5150 ( .A1(n4845), .A2(n4846), .ZN(n4152) );
  NAND2_X1 U5151 ( .A1(n4150), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4151)
         );
  NAND2_X1 U5152 ( .A1(n4152), .A2(n4151), .ZN(n5157) );
  NAND2_X1 U5153 ( .A1(n4154), .A2(n4153), .ZN(n4160) );
  INV_X1 U5154 ( .A(n4155), .ZN(n4157) );
  NAND2_X1 U5155 ( .A1(n4157), .A2(n4156), .ZN(n4168) );
  XNOR2_X1 U5156 ( .A(n4168), .B(n4169), .ZN(n4158) );
  NAND2_X1 U5157 ( .A1(n4158), .A2(n5273), .ZN(n4159) );
  NAND2_X1 U5158 ( .A1(n4160), .A2(n4159), .ZN(n4161) );
  INV_X1 U5159 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6386) );
  NAND2_X1 U5160 ( .A1(n5157), .A2(n5158), .ZN(n4163) );
  NAND2_X1 U5161 ( .A1(n4161), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4162)
         );
  INV_X1 U5162 ( .A(n4168), .ZN(n4170) );
  NAND3_X1 U5163 ( .A1(n4170), .A2(n5273), .A3(n4169), .ZN(n4171) );
  XNOR2_X1 U5164 ( .A(n4172), .B(n5075), .ZN(n5066) );
  INV_X1 U5165 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6764) );
  NAND2_X1 U5166 ( .A1(n5760), .A2(n6764), .ZN(n4175) );
  INV_X1 U5167 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5957) );
  AND2_X1 U5168 ( .A1(n5760), .A2(n5957), .ZN(n5784) );
  INV_X1 U5169 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6369) );
  NAND2_X1 U5170 ( .A1(n5760), .A2(n6369), .ZN(n5769) );
  INV_X1 U5171 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5761) );
  NAND2_X1 U5172 ( .A1(n5760), .A2(n5761), .ZN(n4176) );
  OAI21_X1 U5173 ( .B1(INSTADDRPOINTER_REG_11__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .A(n5716), .ZN(n4177) );
  INV_X4 U5174 ( .A(n5716), .ZN(n5762) );
  XNOR2_X1 U5175 ( .A(n5762), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5754)
         );
  INV_X1 U5176 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4352) );
  INV_X1 U5177 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5912) );
  NAND2_X1 U5178 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n4357) );
  NOR2_X1 U5179 ( .A1(n4357), .A2(n5897), .ZN(n4382) );
  NAND2_X1 U5180 ( .A1(n4382), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n4179) );
  INV_X1 U5181 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n6714) );
  INV_X1 U5182 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5885) );
  NAND4_X1 U5183 ( .A1(n5907), .A2(n6714), .A3(n5897), .A4(n5885), .ZN(n4180)
         );
  AND2_X1 U5184 ( .A1(INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5837) );
  AND2_X1 U5185 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5839) );
  NAND2_X1 U5186 ( .A1(n5837), .A2(n5839), .ZN(n4366) );
  NAND2_X1 U5187 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4367) );
  OAI21_X1 U5188 ( .B1(n4366), .B2(n4367), .A(n5762), .ZN(n4181) );
  NOR2_X1 U5189 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5838) );
  NOR2_X1 U5190 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4182) );
  INV_X1 U5191 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n4377) );
  NAND4_X1 U5192 ( .A1(n5838), .A2(n4182), .A3(n4380), .A4(n4377), .ZN(n4183)
         );
  NAND2_X1 U5193 ( .A1(n5716), .A2(n4183), .ZN(n4184) );
  NAND2_X1 U5194 ( .A1(n4185), .A2(n4184), .ZN(n5646) );
  INV_X1 U5195 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5648) );
  XNOR2_X1 U5196 ( .A(n5762), .B(n5648), .ZN(n5679) );
  OR2_X2 U5197 ( .A1(n5646), .A2(n5679), .ZN(n4187) );
  NAND2_X1 U5198 ( .A1(n5760), .A2(n5648), .ZN(n4186) );
  NAND2_X1 U5199 ( .A1(n5760), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5668) );
  AND2_X1 U5200 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4369) );
  INV_X1 U5201 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5641) );
  INV_X1 U5202 ( .A(n4187), .ZN(n5678) );
  NOR2_X1 U5203 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4188) );
  NAND2_X1 U5204 ( .A1(n5667), .A2(n4188), .ZN(n5312) );
  NOR3_X1 U5205 ( .A1(n5312), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4189) );
  INV_X1 U5206 ( .A(n4376), .ZN(n4194) );
  NAND2_X1 U5207 ( .A1(n4194), .A2(n4193), .ZN(n4204) );
  NAND2_X1 U5208 ( .A1(n6428), .A2(n4198), .ZN(n6680) );
  NAND2_X1 U5209 ( .A1(n6680), .A2(n6603), .ZN(n4199) );
  NAND2_X1 U5210 ( .A1(n6091), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4659) );
  NAND2_X1 U5211 ( .A1(n6603), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4200) );
  NAND2_X1 U5212 ( .A1(n4659), .A2(n4200), .ZN(n4457) );
  NAND2_X1 U5213 ( .A1(n6603), .A2(n6527), .ZN(n4658) );
  INV_X1 U5214 ( .A(REIP_REG_31__SCAN_IN), .ZN(n6813) );
  NOR2_X1 U5215 ( .A1(n6398), .A2(n6813), .ZN(n4371) );
  AOI21_X1 U5216 ( .B1(n6351), .B2(PHYADDRPOINTER_REG_31__SCAN_IN), .A(n4371), 
        .ZN(n4201) );
  OAI21_X1 U5217 ( .B1(n5271), .B2(n6362), .A(n4201), .ZN(n4202) );
  AOI21_X1 U5218 ( .B1(n5296), .B2(n6358), .A(n4202), .ZN(n4203) );
  NAND2_X1 U5219 ( .A1(n4204), .A2(n4203), .ZN(U2955) );
  INV_X1 U5220 ( .A(n4348), .ZN(n4205) );
  NAND2_X1 U5221 ( .A1(n4509), .A2(n4205), .ZN(n4465) );
  NAND2_X1 U5222 ( .A1(n4342), .A2(n4206), .ZN(n4207) );
  OR2_X1 U5223 ( .A1(n4208), .A2(n4207), .ZN(n4211) );
  NAND2_X1 U5224 ( .A1(n4211), .A2(n4423), .ZN(n4469) );
  OAI211_X1 U5225 ( .C1(n3345), .C2(n4630), .A(n4337), .B(n4213), .ZN(n4214)
         );
  NAND3_X1 U5226 ( .A1(n4465), .A2(n4469), .A3(n4214), .ZN(n4215) );
  NAND2_X1 U5227 ( .A1(n4215), .A2(n4663), .ZN(n4221) );
  OR2_X1 U5228 ( .A1(n3326), .A2(n4630), .ZN(n5248) );
  NAND2_X1 U5229 ( .A1(n5248), .A2(n6793), .ZN(n4218) );
  OAI211_X1 U5230 ( .C1(n4217), .C2(n4218), .A(n5246), .B(n3352), .ZN(n4219)
         );
  INV_X1 U5231 ( .A(n4219), .ZN(n4220) );
  NAND2_X2 U5232 ( .A1(n3326), .A2(n5246), .ZN(n4263) );
  OAI22_X1 U5233 ( .A1(n4217), .A2(n4263), .B1(n4329), .B2(n3320), .ZN(n4222)
         );
  INV_X1 U5234 ( .A(n4222), .ZN(n4223) );
  NAND4_X1 U5235 ( .A1(n4081), .A2(n4223), .A3(n4537), .A4(n4622), .ZN(n4224)
         );
  INV_X1 U5236 ( .A(n4312), .ZN(n4226) );
  INV_X1 U5237 ( .A(EBX_REG_1__SCAN_IN), .ZN(n4225) );
  INV_X1 U5238 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6400) );
  NAND2_X1 U5239 ( .A1(n4274), .A2(n6400), .ZN(n4228) );
  NAND2_X1 U5240 ( .A1(n4490), .A2(n4225), .ZN(n4227) );
  NAND3_X1 U5241 ( .A1(n4228), .A2(n2969), .A3(n4227), .ZN(n4229) );
  NAND2_X1 U5242 ( .A1(n4274), .A2(EBX_REG_0__SCAN_IN), .ZN(n4232) );
  INV_X1 U5243 ( .A(EBX_REG_0__SCAN_IN), .ZN(n5542) );
  NAND2_X1 U5244 ( .A1(n2969), .A2(n5542), .ZN(n4231) );
  NAND2_X1 U5245 ( .A1(n4232), .A2(n4231), .ZN(n4440) );
  XNOR2_X1 U5246 ( .A(n4233), .B(n4440), .ZN(n4488) );
  NAND2_X1 U5247 ( .A1(n4489), .A2(n4233), .ZN(n4593) );
  MUX2_X1 U5248 ( .A(n4322), .B(n2969), .S(EBX_REG_3__SCAN_IN), .Z(n4236) );
  NAND2_X2 U5249 ( .A1(n4274), .A2(n2969), .ZN(n4441) );
  OR2_X1 U5250 ( .A1(n4441), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4235)
         );
  NAND2_X1 U5251 ( .A1(n4236), .A2(n4235), .ZN(n4595) );
  INV_X1 U5252 ( .A(n4595), .ZN(n4240) );
  MUX2_X1 U5253 ( .A(n4312), .B(n4274), .S(EBX_REG_2__SCAN_IN), .Z(n4239) );
  OR2_X1 U5254 ( .A1(n4490), .A2(n4274), .ZN(n4282) );
  NAND2_X1 U5255 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n4326), .ZN(n4237)
         );
  AND2_X1 U5256 ( .A1(n4282), .A2(n4237), .ZN(n4238) );
  NAND2_X1 U5257 ( .A1(n4239), .A2(n4238), .ZN(n4594) );
  OR2_X1 U5258 ( .A1(n4312), .A2(EBX_REG_4__SCAN_IN), .ZN(n4247) );
  NAND2_X1 U5259 ( .A1(n4274), .A2(n4242), .ZN(n4245) );
  INV_X1 U5260 ( .A(EBX_REG_4__SCAN_IN), .ZN(n4243) );
  NAND2_X1 U5261 ( .A1(n4490), .A2(n4243), .ZN(n4244) );
  NAND3_X1 U5262 ( .A1(n4245), .A2(n2969), .A3(n4244), .ZN(n4246) );
  AND2_X1 U5263 ( .A1(n4247), .A2(n4246), .ZN(n4641) );
  MUX2_X1 U5264 ( .A(n4322), .B(n2969), .S(EBX_REG_5__SCAN_IN), .Z(n4248) );
  OAI21_X1 U5265 ( .B1(INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n4441), .A(n4248), 
        .ZN(n4739) );
  INV_X1 U5266 ( .A(n4739), .ZN(n4249) );
  OR2_X1 U5267 ( .A1(n4312), .A2(EBX_REG_6__SCAN_IN), .ZN(n4253) );
  NAND2_X1 U5268 ( .A1(n4274), .A2(n6780), .ZN(n4251) );
  INV_X1 U5269 ( .A(EBX_REG_6__SCAN_IN), .ZN(n5514) );
  NAND2_X1 U5270 ( .A1(n4490), .A2(n5514), .ZN(n4250) );
  NAND3_X1 U5271 ( .A1(n4251), .A2(n2969), .A3(n4250), .ZN(n4252) );
  NAND2_X1 U5272 ( .A1(n4253), .A2(n4252), .ZN(n4794) );
  NAND2_X1 U5273 ( .A1(n4738), .A2(n4794), .ZN(n4793) );
  MUX2_X1 U5274 ( .A(n4322), .B(n2969), .S(EBX_REG_7__SCAN_IN), .Z(n4254) );
  OAI21_X1 U5275 ( .B1(INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n4441), .A(n4254), 
        .ZN(n4969) );
  NOR2_X2 U5276 ( .A1(n4793), .A2(n4969), .ZN(n4967) );
  OR2_X1 U5277 ( .A1(n4312), .A2(EBX_REG_8__SCAN_IN), .ZN(n4258) );
  NAND2_X1 U5278 ( .A1(n4274), .A2(n5075), .ZN(n4256) );
  INV_X1 U5279 ( .A(EBX_REG_8__SCAN_IN), .ZN(n6179) );
  NAND2_X1 U5280 ( .A1(n4490), .A2(n6179), .ZN(n4255) );
  NAND3_X1 U5281 ( .A1(n4256), .A2(n2969), .A3(n4255), .ZN(n4257) );
  NAND2_X1 U5282 ( .A1(n4258), .A2(n4257), .ZN(n5061) );
  NAND2_X1 U5283 ( .A1(n4967), .A2(n5061), .ZN(n5008) );
  MUX2_X1 U5284 ( .A(n4322), .B(n4259), .S(EBX_REG_9__SCAN_IN), .Z(n4260) );
  OAI21_X1 U5285 ( .B1(INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n4441), .A(n4260), 
        .ZN(n5010) );
  MUX2_X1 U5286 ( .A(n4312), .B(n4274), .S(EBX_REG_10__SCAN_IN), .Z(n4265) );
  NAND2_X1 U5287 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n4326), .ZN(n4264) );
  NAND2_X1 U5288 ( .A1(n2969), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n4266) );
  OAI211_X1 U5289 ( .C1(n4326), .C2(EBX_REG_11__SCAN_IN), .A(n4274), .B(n4266), 
        .ZN(n4267) );
  OAI21_X1 U5290 ( .B1(n4322), .B2(EBX_REG_11__SCAN_IN), .A(n4267), .ZN(n5230)
         );
  MUX2_X1 U5291 ( .A(n4312), .B(n4274), .S(EBX_REG_12__SCAN_IN), .Z(n4270) );
  NAND2_X1 U5292 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n4326), .ZN(n4268) );
  AND2_X1 U5293 ( .A1(n4282), .A2(n4268), .ZN(n4269) );
  NAND2_X1 U5294 ( .A1(n4270), .A2(n4269), .ZN(n5930) );
  INV_X1 U5295 ( .A(n4322), .ZN(n4285) );
  INV_X1 U5296 ( .A(EBX_REG_13__SCAN_IN), .ZN(n6808) );
  NAND2_X1 U5297 ( .A1(n4285), .A2(n6808), .ZN(n4273) );
  NAND2_X1 U5298 ( .A1(n2969), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4271) );
  OAI211_X1 U5299 ( .C1(n4326), .C2(EBX_REG_13__SCAN_IN), .A(n4274), .B(n4271), 
        .ZN(n4272) );
  MUX2_X1 U5300 ( .A(n4312), .B(n4274), .S(EBX_REG_14__SCAN_IN), .Z(n4277) );
  NAND2_X1 U5301 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n4326), .ZN(n4275) );
  AND2_X1 U5302 ( .A1(n4282), .A2(n4275), .ZN(n4276) );
  NAND2_X1 U5303 ( .A1(n4277), .A2(n4276), .ZN(n5585) );
  NAND2_X1 U5304 ( .A1(n5929), .A2(n5585), .ZN(n5577) );
  NAND2_X1 U5305 ( .A1(n4441), .A2(EBX_REG_15__SCAN_IN), .ZN(n4279) );
  NAND2_X1 U5306 ( .A1(n4326), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n4278) );
  NAND2_X1 U5307 ( .A1(n4279), .A2(n4278), .ZN(n4280) );
  XNOR2_X1 U5308 ( .A(n4280), .B(n5449), .ZN(n5580) );
  NOR2_X2 U5309 ( .A1(n5577), .A2(n5580), .ZN(n5568) );
  MUX2_X1 U5310 ( .A(n4312), .B(n4274), .S(EBX_REG_16__SCAN_IN), .Z(n4283) );
  NAND2_X1 U5311 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n4326), .ZN(n4281) );
  AND2_X2 U5312 ( .A1(n5568), .A2(n4284), .ZN(n5570) );
  INV_X1 U5313 ( .A(EBX_REG_17__SCAN_IN), .ZN(n5562) );
  NAND2_X1 U5314 ( .A1(n4285), .A2(n5562), .ZN(n4288) );
  NAND2_X1 U5315 ( .A1(n2969), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n4286) );
  OAI211_X1 U5316 ( .C1(EBX_REG_17__SCAN_IN), .C2(n4326), .A(n4274), .B(n4286), 
        .ZN(n4287) );
  OR2_X1 U5317 ( .A1(n4312), .A2(EBX_REG_19__SCAN_IN), .ZN(n4291) );
  NAND2_X1 U5318 ( .A1(n4274), .A2(n4377), .ZN(n4289) );
  OAI211_X1 U5319 ( .C1(EBX_REG_19__SCAN_IN), .C2(n4326), .A(n4289), .B(n2969), 
        .ZN(n4290) );
  OR2_X1 U5320 ( .A1(n4441), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4292)
         );
  INV_X1 U5321 ( .A(EBX_REG_18__SCAN_IN), .ZN(n5483) );
  NAND2_X1 U5322 ( .A1(n4490), .A2(n5483), .ZN(n5466) );
  OAI22_X1 U5323 ( .A1(n4441), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        EBX_REG_20__SCAN_IN), .B2(n4326), .ZN(n5450) );
  NAND2_X1 U5324 ( .A1(n5464), .A2(n5450), .ZN(n4294) );
  NAND2_X1 U5325 ( .A1(n5449), .A2(EBX_REG_20__SCAN_IN), .ZN(n4293) );
  OAI211_X1 U5326 ( .C1(n5464), .C2(n5449), .A(n4294), .B(n4293), .ZN(n4295)
         );
  MUX2_X1 U5327 ( .A(n4322), .B(n2969), .S(EBX_REG_21__SCAN_IN), .Z(n4297) );
  OR2_X1 U5328 ( .A1(n4441), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n4296)
         );
  OR2_X1 U5329 ( .A1(n4312), .A2(EBX_REG_22__SCAN_IN), .ZN(n4300) );
  INV_X1 U5330 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n6783) );
  NAND2_X1 U5331 ( .A1(n4274), .A2(n6783), .ZN(n4298) );
  OAI211_X1 U5332 ( .C1(EBX_REG_22__SCAN_IN), .C2(n4326), .A(n4298), .B(n2969), 
        .ZN(n4299) );
  NAND2_X1 U5333 ( .A1(n4300), .A2(n4299), .ZN(n5422) );
  NAND2_X1 U5334 ( .A1(n5423), .A2(n5422), .ZN(n4392) );
  NAND2_X1 U5335 ( .A1(n2969), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4301) );
  OAI211_X1 U5336 ( .C1(EBX_REG_23__SCAN_IN), .C2(n4326), .A(n4274), .B(n4301), 
        .ZN(n4302) );
  OAI21_X1 U5337 ( .B1(n4322), .B2(EBX_REG_23__SCAN_IN), .A(n4302), .ZN(n4393)
         );
  OR2_X2 U5338 ( .A1(n4392), .A2(n4393), .ZN(n5302) );
  MUX2_X1 U5339 ( .A(n4312), .B(n4274), .S(EBX_REG_24__SCAN_IN), .Z(n4304) );
  NAND2_X1 U5340 ( .A1(n4326), .A2(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4303) );
  MUX2_X1 U5341 ( .A(n4322), .B(n2969), .S(EBX_REG_25__SCAN_IN), .Z(n4306) );
  OR2_X1 U5342 ( .A1(n4441), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n4305)
         );
  NAND2_X1 U5343 ( .A1(n4306), .A2(n4305), .ZN(n5399) );
  INV_X1 U5344 ( .A(n5399), .ZN(n4307) );
  OR2_X1 U5345 ( .A1(n4312), .A2(EBX_REG_26__SCAN_IN), .ZN(n4310) );
  INV_X1 U5346 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5650) );
  NAND2_X1 U5347 ( .A1(n4274), .A2(n5650), .ZN(n4308) );
  OAI211_X1 U5348 ( .C1(EBX_REG_26__SCAN_IN), .C2(n4326), .A(n4308), .B(n2969), 
        .ZN(n4309) );
  NAND2_X1 U5349 ( .A1(n4310), .A2(n4309), .ZN(n5385) );
  MUX2_X1 U5350 ( .A(n4322), .B(n2969), .S(EBX_REG_27__SCAN_IN), .Z(n4311) );
  OAI21_X1 U5351 ( .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n4441), .A(n4311), 
        .ZN(n5372) );
  OR2_X1 U5352 ( .A1(n4312), .A2(EBX_REG_28__SCAN_IN), .ZN(n4315) );
  INV_X1 U5353 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5802) );
  NAND2_X1 U5354 ( .A1(n4274), .A2(n5802), .ZN(n4313) );
  OAI211_X1 U5355 ( .C1(EBX_REG_28__SCAN_IN), .C2(n4326), .A(n4313), .B(n2969), 
        .ZN(n4314) );
  OR2_X1 U5356 ( .A1(n4441), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4320)
         );
  INV_X1 U5357 ( .A(EBX_REG_29__SCAN_IN), .ZN(n4316) );
  NAND2_X1 U5358 ( .A1(n4490), .A2(n4316), .ZN(n4317) );
  AND2_X1 U5359 ( .A1(n4320), .A2(n4317), .ZN(n4318) );
  AND2_X1 U5360 ( .A1(n4263), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4319)
         );
  AOI21_X1 U5361 ( .B1(n4441), .B2(EBX_REG_30__SCAN_IN), .A(n4319), .ZN(n5241)
         );
  INV_X1 U5362 ( .A(n4320), .ZN(n4321) );
  MUX2_X1 U5363 ( .A(EBX_REG_29__SCAN_IN), .B(n4321), .S(n2969), .Z(n4324) );
  NOR2_X1 U5364 ( .A1(n4322), .A2(EBX_REG_29__SCAN_IN), .ZN(n4323) );
  NOR2_X1 U5365 ( .A1(n4324), .A2(n4323), .ZN(n5351) );
  NAND3_X1 U5366 ( .A1(n5362), .A2(n5241), .A3(n5351), .ZN(n4325) );
  NAND2_X1 U5367 ( .A1(n5240), .A2(n4325), .ZN(n4328) );
  OAI22_X1 U5368 ( .A1(n4441), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        EBX_REG_31__SCAN_IN), .B2(n4326), .ZN(n4327) );
  INV_X1 U5369 ( .A(n5294), .ZN(n4331) );
  OAI21_X1 U5370 ( .B1(n4329), .B2(n3333), .A(n4648), .ZN(n4330) );
  NAND2_X1 U5371 ( .A1(n4331), .A2(n6395), .ZN(n4374) );
  INV_X1 U5372 ( .A(n4483), .ZN(n4333) );
  OR3_X1 U5373 ( .A1(n4333), .A2(n4518), .A3(n5246), .ZN(n4559) );
  NAND2_X1 U5374 ( .A1(n4334), .A2(n5449), .ZN(n4335) );
  OAI211_X1 U5375 ( .C1(n4090), .C2(n4332), .A(n4559), .B(n4335), .ZN(n4347)
         );
  INV_X1 U5376 ( .A(n4336), .ZN(n4344) );
  AOI22_X1 U5377 ( .A1(n4338), .A2(n5449), .B1(n4337), .B2(n3352), .ZN(n4343)
         );
  AND2_X1 U5378 ( .A1(n4709), .A2(n4339), .ZN(n5525) );
  AND2_X1 U5379 ( .A1(n5525), .A2(n4692), .ZN(n4467) );
  OAI21_X1 U5380 ( .B1(n4467), .B2(n4441), .A(n4340), .ZN(n4341) );
  AND4_X1 U5381 ( .A1(n4344), .A2(n4343), .A3(n4342), .A4(n4341), .ZN(n4346)
         );
  NAND2_X1 U5382 ( .A1(n4346), .A2(n4345), .ZN(n4505) );
  INV_X1 U5383 ( .A(n5955), .ZN(n5894) );
  NAND2_X1 U5384 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n4368) );
  OR2_X1 U5385 ( .A1(n4350), .A2(n6350), .ZN(n4443) );
  NOR2_X1 U5386 ( .A1(n6392), .A2(n5922), .ZN(n5920) );
  OR2_X1 U5387 ( .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n5920), .ZN(n4442)
         );
  NAND2_X1 U5388 ( .A1(n5955), .A2(n4496), .ZN(n4359) );
  INV_X1 U5389 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6389) );
  OAI21_X1 U5390 ( .B1(n6400), .B2(n6389), .A(n4119), .ZN(n6388) );
  NAND3_X1 U5391 ( .A1(INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_3__SCAN_IN), .A3(n6388), .ZN(n4736) );
  NOR2_X1 U5392 ( .A1(n4740), .A2(n4736), .ZN(n4848) );
  NAND2_X1 U5393 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n4848), .ZN(n5069)
         );
  NOR2_X1 U5394 ( .A1(n6386), .A2(n5075), .ZN(n5956) );
  NAND3_X1 U5395 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A3(n5956), .ZN(n4353) );
  NOR2_X1 U5396 ( .A1(n5069), .A2(n4353), .ZN(n4363) );
  INV_X1 U5397 ( .A(n4363), .ZN(n4351) );
  NAND2_X1 U5398 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5947) );
  NOR2_X1 U5399 ( .A1(n5947), .A2(n4352), .ZN(n5916) );
  NAND2_X1 U5400 ( .A1(n5916), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5895) );
  OR3_X1 U5401 ( .A1(n5895), .A2(n5907), .A3(n5897), .ZN(n4355) );
  NAND2_X1 U5402 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4638) );
  NAND2_X1 U5403 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6390) );
  NOR2_X1 U5404 ( .A1(n4638), .A2(n6390), .ZN(n4741) );
  NAND3_X1 U5405 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_6__SCAN_IN), .A3(n4741), .ZN(n5074) );
  NOR2_X1 U5406 ( .A1(n4353), .A2(n5074), .ZN(n5890) );
  INV_X1 U5407 ( .A(n4355), .ZN(n4364) );
  AOI21_X1 U5408 ( .B1(n5890), .B2(n4364), .A(n4361), .ZN(n4354) );
  AOI21_X1 U5409 ( .B1(n6392), .B2(n4355), .A(n4354), .ZN(n4356) );
  INV_X1 U5410 ( .A(n4357), .ZN(n4365) );
  NAND2_X1 U5411 ( .A1(n4359), .A2(n4358), .ZN(n5836) );
  OR2_X1 U5412 ( .A1(n5955), .A2(n5839), .ZN(n4360) );
  NOR2_X1 U5413 ( .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n5918), .ZN(n4495)
         );
  OR2_X1 U5414 ( .A1(n6392), .A2(n6402), .ZN(n5856) );
  NAND2_X1 U5415 ( .A1(n5856), .A2(n4367), .ZN(n4362) );
  OAI21_X1 U5416 ( .B1(n5955), .B2(INSTADDRPOINTER_REG_30__SCAN_IN), .A(n5315), 
        .ZN(n4372) );
  NAND2_X1 U5417 ( .A1(n6392), .A2(n4363), .ZN(n5924) );
  NAND2_X1 U5418 ( .A1(n5890), .A2(n6402), .ZN(n5946) );
  INV_X1 U5419 ( .A(n4366), .ZN(n5304) );
  NAND2_X1 U5420 ( .A1(n5854), .A2(n5304), .ZN(n4397) );
  NAND2_X1 U5421 ( .A1(n5806), .A2(n4369), .ZN(n5794) );
  AOI211_X1 U5422 ( .C1(n4372), .C2(INSTADDRPOINTER_REG_31__SCAN_IN), .A(n4371), .B(n4370), .ZN(n4373) );
  OAI21_X1 U5423 ( .B1(n4376), .B2(n5961), .A(n4375), .ZN(U2987) );
  XNOR2_X1 U5424 ( .A(n5762), .B(n4377), .ZN(n5709) );
  AND2_X1 U5425 ( .A1(n5760), .A2(n4380), .ZN(n4379) );
  XNOR2_X1 U5426 ( .A(n5762), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5694)
         );
  NAND2_X2 U5427 ( .A1(n5695), .A2(n5694), .ZN(n5693) );
  XNOR2_X1 U5428 ( .A(n5762), .B(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5739)
         );
  NAND2_X1 U5429 ( .A1(n5740), .A2(n5739), .ZN(n5903) );
  NAND3_X1 U5430 ( .A1(n5734), .A2(n4382), .A3(n5304), .ZN(n4383) );
  OAI21_X1 U5431 ( .B1(n2990), .B2(n4387), .A(n4386), .ZN(n5615) );
  AND2_X1 U5432 ( .A1(n6350), .A2(REIP_REG_23__SCAN_IN), .ZN(n4399) );
  NOR2_X1 U5433 ( .A1(n5414), .A2(n6362), .ZN(n4388) );
  AOI211_X1 U5434 ( .C1(PHYADDRPOINTER_REG_23__SCAN_IN), .C2(n6351), .A(n4399), 
        .B(n4388), .ZN(n4389) );
  NAND2_X1 U5435 ( .A1(n4391), .A2(n6403), .ZN(n4404) );
  INV_X1 U5436 ( .A(n4392), .ZN(n4395) );
  INV_X1 U5437 ( .A(n4393), .ZN(n4394) );
  OAI21_X1 U5438 ( .B1(n4395), .B2(n4394), .A(n5302), .ZN(n5555) );
  INV_X1 U5439 ( .A(n4396), .ZN(n4400) );
  NOR2_X1 U5440 ( .A1(n4397), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4398)
         );
  AOI211_X1 U5441 ( .C1(INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n4400), .A(n4399), .B(n4398), .ZN(n4401) );
  NAND2_X1 U5442 ( .A1(n4404), .A2(n4403), .ZN(U2995) );
  NAND2_X1 U5443 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATE2_REG_1__SCAN_IN), 
        .ZN(n4580) );
  INV_X1 U5444 ( .A(n4580), .ZN(n4653) );
  NAND2_X1 U5445 ( .A1(n4653), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4634) );
  INV_X1 U5446 ( .A(n4634), .ZN(n4578) );
  NOR2_X1 U5447 ( .A1(n6793), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4657) );
  NOR4_X1 U5448 ( .A1(n4578), .A2(n4657), .A3(n6683), .A4(n4405), .ZN(n4407)
         );
  OR2_X1 U5449 ( .A1(n4407), .A2(n4406), .ZN(U3150) );
  INV_X1 U5450 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6800) );
  NOR2_X1 U5451 ( .A1(n6793), .A2(n6800), .ZN(n6079) );
  AOI21_X1 U5452 ( .B1(HOLD), .B2(STATE_REG_2__SCAN_IN), .A(n6079), .ZN(n4416)
         );
  AND2_X1 U5453 ( .A1(STATE_REG_1__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n4415) );
  INV_X1 U5454 ( .A(n4415), .ZN(n4412) );
  INV_X1 U5455 ( .A(NA_N), .ZN(n6829) );
  AOI21_X1 U5456 ( .B1(n6829), .B2(READY_N), .A(n6800), .ZN(n4408) );
  INV_X1 U5457 ( .A(HOLD), .ZN(n6076) );
  AOI211_X1 U5458 ( .C1(REQUESTPENDING_REG_SCAN_IN), .C2(n6610), .A(n4408), 
        .B(n6076), .ZN(n4409) );
  INV_X1 U5459 ( .A(STATE_REG_0__SCAN_IN), .ZN(n6083) );
  OAI221_X1 U5460 ( .B1(n6610), .B2(NA_N), .C1(n6610), .C2(n6800), .A(n6083), 
        .ZN(n4413) );
  OAI21_X1 U5461 ( .B1(n4409), .B2(n6083), .A(n4413), .ZN(n4411) );
  NAND4_X1 U5462 ( .A1(STATE_REG_0__SCAN_IN), .A2(REQUESTPENDING_REG_SCAN_IN), 
        .A3(n6079), .A4(n6829), .ZN(n4410) );
  OAI211_X1 U5463 ( .C1(n4416), .C2(n4412), .A(n4411), .B(n4410), .ZN(U3183)
         );
  NOR2_X1 U5464 ( .A1(n6800), .A2(n6076), .ZN(n6077) );
  INV_X1 U5465 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6075) );
  OAI21_X1 U5466 ( .B1(n6077), .B2(n6075), .A(n6678), .ZN(n4414) );
  OAI211_X1 U5467 ( .C1(n4416), .C2(n4415), .A(n4414), .B(n4413), .ZN(U3181)
         );
  NOR2_X1 U5468 ( .A1(n4427), .A2(n4423), .ZN(n4419) );
  NAND2_X1 U5469 ( .A1(n4419), .A2(n4663), .ZN(n5234) );
  NAND2_X1 U5470 ( .A1(n6524), .A2(n4629), .ZN(n6087) );
  INV_X1 U5471 ( .A(n6087), .ZN(n5468) );
  INV_X1 U5472 ( .A(n5235), .ZN(n4431) );
  AOI211_X1 U5473 ( .C1(MEMORYFETCH_REG_SCAN_IN), .C2(n5234), .A(n5468), .B(
        n4431), .ZN(n4417) );
  INV_X1 U5474 ( .A(n4417), .ZN(U2788) );
  NAND2_X1 U5475 ( .A1(n4509), .A2(n5345), .ZN(n4421) );
  INV_X1 U5476 ( .A(n4076), .ZN(n4418) );
  OR2_X1 U5477 ( .A1(n4419), .A2(n4418), .ZN(n4420) );
  NAND2_X1 U5478 ( .A1(n4421), .A2(n4420), .ZN(n6085) );
  NAND3_X1 U5479 ( .A1(n5345), .A2(n6082), .A3(n4263), .ZN(n4422) );
  AND2_X1 U5480 ( .A1(n4422), .A2(n6793), .ZN(n6682) );
  NOR2_X1 U5481 ( .A1(n6085), .A2(n6682), .ZN(n4620) );
  OR2_X1 U5482 ( .A1(n4620), .A2(n6608), .ZN(n4428) );
  INV_X1 U5483 ( .A(n4428), .ZN(n6094) );
  INV_X1 U5484 ( .A(MORE_REG_SCAN_IN), .ZN(n4430) );
  INV_X1 U5485 ( .A(n4423), .ZN(n4426) );
  NAND3_X1 U5486 ( .A1(n4537), .A2(n4622), .A3(n4076), .ZN(n4424) );
  MUX2_X1 U5487 ( .A(n4539), .B(n4424), .S(n4509), .Z(n4425) );
  AOI21_X1 U5488 ( .B1(n4427), .B2(n4426), .A(n4425), .ZN(n4623) );
  OR2_X1 U5489 ( .A1(n4623), .A2(n4428), .ZN(n4429) );
  OAI21_X1 U5490 ( .B1(n6094), .B2(n4430), .A(n4429), .ZN(U3471) );
  INV_X1 U5491 ( .A(EAX_REG_13__SCAN_IN), .ZN(n6268) );
  INV_X1 U5492 ( .A(LWORD_REG_13__SCAN_IN), .ZN(n4433) );
  OAI21_X1 U5493 ( .B1(n5273), .B2(n6793), .A(n4431), .ZN(n4432) );
  INV_X1 U5494 ( .A(DATAI_13_), .ZN(n6716) );
  OAI222_X1 U5495 ( .A1(n6348), .A2(n6268), .B1(n4433), .B2(n6298), .C1(n6307), 
        .C2(n6716), .ZN(U2952) );
  INV_X1 U5496 ( .A(UWORD_REG_11__SCAN_IN), .ZN(n6718) );
  INV_X1 U5497 ( .A(DATAI_11_), .ZN(n4434) );
  NOR2_X1 U5498 ( .A1(n6307), .A2(n4434), .ZN(n6339) );
  INV_X1 U5499 ( .A(n6339), .ZN(n4436) );
  NAND2_X1 U5500 ( .A1(n6343), .A2(EAX_REG_27__SCAN_IN), .ZN(n4435) );
  OAI211_X1 U5501 ( .C1(n6298), .C2(n6718), .A(n4436), .B(n4435), .ZN(U2935)
         );
  INV_X1 U5502 ( .A(UWORD_REG_2__SCAN_IN), .ZN(n6823) );
  AND2_X1 U5503 ( .A1(n6346), .A2(DATAI_2_), .ZN(n6319) );
  INV_X1 U5504 ( .A(n6319), .ZN(n4438) );
  NAND2_X1 U5505 ( .A1(n6343), .A2(EAX_REG_18__SCAN_IN), .ZN(n4437) );
  OAI211_X1 U5506 ( .C1(n6298), .C2(n6823), .A(n4438), .B(n4437), .ZN(U2926)
         );
  INV_X1 U5507 ( .A(DATAI_7_), .ZN(n4699) );
  AOI22_X1 U5508 ( .A1(n6332), .A2(LWORD_REG_7__SCAN_IN), .B1(
        EAX_REG_7__SCAN_IN), .B2(n6343), .ZN(n4439) );
  OAI21_X1 U5509 ( .B1(n4699), .B2(n6307), .A(n4439), .ZN(U2946) );
  OAI21_X1 U5510 ( .B1(n4441), .B2(INSTADDRPOINTER_REG_0__SCAN_IN), .A(n4440), 
        .ZN(n5543) );
  INV_X1 U5511 ( .A(n5543), .ZN(n4447) );
  INV_X1 U5512 ( .A(REIP_REG_0__SCAN_IN), .ZN(n6675) );
  OAI21_X1 U5513 ( .B1(n6398), .B2(n6675), .A(n4442), .ZN(n4446) );
  INV_X1 U5514 ( .A(n5918), .ZN(n4444) );
  AOI21_X1 U5515 ( .B1(n4444), .B2(n4443), .A(n6389), .ZN(n4445) );
  AOI211_X1 U5516 ( .C1(n4447), .C2(n6395), .A(n4446), .B(n4445), .ZN(n4450)
         );
  OR2_X1 U5517 ( .A1(n4448), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4460)
         );
  NAND3_X1 U5518 ( .A1(n4460), .A2(n6403), .A3(n4459), .ZN(n4449) );
  NAND2_X1 U5519 ( .A1(n4450), .A2(n4449), .ZN(U3018) );
  INV_X1 U5520 ( .A(n4451), .ZN(n4454) );
  OAI21_X1 U5521 ( .B1(n4454), .B2(n4453), .A(n4452), .ZN(n5548) );
  NAND2_X1 U5522 ( .A1(n3328), .A2(n3313), .ZN(n4455) );
  INV_X1 U5523 ( .A(n4455), .ZN(n4456) );
  INV_X1 U5524 ( .A(DATAI_0_), .ZN(n4708) );
  INV_X1 U5525 ( .A(EAX_REG_0__SCAN_IN), .ZN(n6315) );
  OAI222_X1 U5526 ( .A1(n5548), .A2(n5635), .B1(n4844), .B2(n4708), .C1(n6261), 
        .C2(n6315), .ZN(U2891) );
  OR2_X1 U5527 ( .A1(n6351), .A2(n4457), .ZN(n4458) );
  AOI22_X1 U5528 ( .A1(n4458), .A2(PHYADDRPOINTER_REG_0__SCAN_IN), .B1(n6350), 
        .B2(REIP_REG_0__SCAN_IN), .ZN(n4462) );
  NAND3_X1 U5529 ( .A1(n4460), .A2(n4193), .A3(n4459), .ZN(n4461) );
  OAI211_X1 U5530 ( .C1(n5548), .C2(n5782), .A(n4462), .B(n4461), .ZN(U2986)
         );
  NAND2_X1 U5531 ( .A1(n4326), .A2(n6082), .ZN(n4463) );
  AOI22_X1 U5532 ( .A1(n4650), .A2(n4630), .B1(n3343), .B2(n4463), .ZN(n4464)
         );
  OR3_X1 U5533 ( .A1(n4509), .A2(READY_N), .A3(n4464), .ZN(n4471) );
  INV_X1 U5534 ( .A(n4465), .ZN(n4466) );
  NOR2_X1 U5535 ( .A1(n4467), .A2(n4466), .ZN(n4468) );
  AND2_X1 U5536 ( .A1(n4469), .A2(n4468), .ZN(n4470) );
  NAND2_X1 U5537 ( .A1(n4471), .A2(n4470), .ZN(n4472) );
  INV_X1 U5538 ( .A(FLUSH_REG_SCAN_IN), .ZN(n6093) );
  OAI22_X1 U5539 ( .A1(n4612), .A2(n6608), .B1(n6093), .B2(n4634), .ZN(n4477)
         );
  INV_X1 U5540 ( .A(n5977), .ZN(n4510) );
  INV_X1 U5541 ( .A(n5982), .ZN(n4975) );
  NOR2_X1 U5542 ( .A1(n4474), .A2(n4975), .ZN(n4476) );
  XNOR2_X1 U5543 ( .A(n4476), .B(n4475), .ZN(n6214) );
  NAND4_X1 U5544 ( .A1(n4477), .A2(n5334), .A3(n4572), .A4(n6214), .ZN(n4478)
         );
  OAI21_X1 U5545 ( .B1(n4475), .B2(n4510), .A(n4478), .ZN(U3455) );
  OAI21_X1 U5546 ( .B1(n4481), .B2(n4480), .A(n4479), .ZN(n5540) );
  NAND2_X1 U5547 ( .A1(n4509), .A2(n4539), .ZN(n4486) );
  INV_X1 U5548 ( .A(n4482), .ZN(n4484) );
  NAND4_X1 U5549 ( .A1(n4484), .A2(n3348), .A3(n4483), .A4(n4490), .ZN(n4485)
         );
  NAND2_X1 U5550 ( .A1(n4486), .A2(n4485), .ZN(n4487) );
  NAND2_X1 U5551 ( .A1(n6250), .A2(n4700), .ZN(n5588) );
  OAI21_X1 U5552 ( .B1(n4488), .B2(n4490), .A(n4489), .ZN(n4500) );
  AOI22_X1 U5553 ( .A1(n6247), .A2(n4500), .B1(EBX_REG_1__SCAN_IN), .B2(n5595), 
        .ZN(n4491) );
  OAI21_X1 U5554 ( .B1(n5540), .B2(n5590), .A(n4491), .ZN(U2858) );
  OAI222_X1 U5555 ( .A1(n5543), .A2(n5588), .B1(n5542), .B2(n6250), .C1(n5548), 
        .C2(n5597), .ZN(U2859) );
  OAI21_X1 U5556 ( .B1(n4494), .B2(n4493), .A(n4492), .ZN(n4533) );
  INV_X1 U5557 ( .A(REIP_REG_1__SCAN_IN), .ZN(n5522) );
  NOR2_X1 U5558 ( .A1(n6398), .A2(n5522), .ZN(n4529) );
  NOR2_X1 U5559 ( .A1(n5955), .A2(n4495), .ZN(n4498) );
  INV_X1 U5560 ( .A(n4496), .ZN(n4497) );
  MUX2_X1 U5561 ( .A(n4498), .B(n4497), .S(INSTADDRPOINTER_REG_1__SCAN_IN), 
        .Z(n4499) );
  AOI211_X1 U5562 ( .C1(n6395), .C2(n4500), .A(n4529), .B(n4499), .ZN(n4501)
         );
  OAI21_X1 U5563 ( .B1(n5961), .B2(n4533), .A(n4501), .ZN(U3017) );
  INV_X1 U5564 ( .A(n4650), .ZN(n4550) );
  NOR2_X1 U5565 ( .A1(n4550), .A2(n4502), .ZN(n4609) );
  INV_X1 U5566 ( .A(n4609), .ZN(n4513) );
  NAND3_X1 U5567 ( .A1(n4217), .A2(n4090), .A3(n4503), .ZN(n4504) );
  OR2_X1 U5568 ( .A1(n4505), .A2(n4504), .ZN(n4506) );
  NOR2_X1 U5569 ( .A1(n4572), .A2(n4506), .ZN(n4564) );
  OAI22_X1 U5570 ( .A1(n5541), .A2(n4564), .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n4518), .ZN(n4610) );
  INV_X1 U5571 ( .A(n4610), .ZN(n4507) );
  NOR2_X1 U5572 ( .A1(n4507), .A2(STATE2_REG_3__SCAN_IN), .ZN(n4508) );
  MUX2_X1 U5573 ( .A(n6389), .B(n4508), .S(n4629), .Z(n4511) );
  OAI21_X1 U5574 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6605), .A(n4510), 
        .ZN(n4524) );
  OAI22_X1 U5575 ( .A1(n4511), .A2(n4524), .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n4510), .ZN(n4512) );
  OAI21_X1 U5576 ( .B1(n4513), .B2(n5975), .A(n4512), .ZN(U3461) );
  INV_X1 U5577 ( .A(n4564), .ZN(n4553) );
  NOR2_X1 U5578 ( .A1(n4517), .A2(n4521), .ZN(n4519) );
  OAI22_X1 U5579 ( .A1(n4550), .A2(n4556), .B1(n4519), .B2(n4518), .ZN(n4520)
         );
  AOI21_X1 U5580 ( .B1(n4515), .B2(n4553), .A(n4520), .ZN(n4611) );
  INV_X1 U5581 ( .A(n4611), .ZN(n4523) );
  AOI22_X1 U5582 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n4190), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n6400), .ZN(n5330) );
  NAND2_X1 U5583 ( .A1(STATE2_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5331) );
  INV_X1 U5584 ( .A(n5331), .ZN(n4522) );
  INV_X1 U5585 ( .A(n6605), .ZN(n5337) );
  AOI222_X1 U5586 ( .A1(n4523), .A2(n5334), .B1(n5330), .B2(n4522), .C1(n4521), 
        .C2(n5337), .ZN(n4526) );
  INV_X1 U5587 ( .A(n4524), .ZN(n4525) );
  OAI22_X1 U5588 ( .A1(n4526), .A2(n5977), .B1(n4028), .B2(n4525), .ZN(U3460)
         );
  INV_X1 U5589 ( .A(n5540), .ZN(n4527) );
  NAND2_X1 U5590 ( .A1(n4527), .A2(n6358), .ZN(n4532) );
  INV_X1 U5591 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n4530) );
  AND2_X1 U5592 ( .A1(n6351), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n4528)
         );
  AOI211_X1 U5593 ( .C1(n4530), .C2(n5778), .A(n4529), .B(n4528), .ZN(n4531)
         );
  OAI211_X1 U5594 ( .C1(n4533), .C2(n6092), .A(n4532), .B(n4531), .ZN(U2985)
         );
  NAND2_X1 U5595 ( .A1(n4556), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4535) );
  AOI22_X1 U5596 ( .A1(n4536), .A2(n4556), .B1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n4535), .ZN(n4551) );
  INV_X1 U5597 ( .A(n4537), .ZN(n4538) );
  OR2_X1 U5598 ( .A1(n4539), .A2(n4538), .ZN(n4562) );
  MUX2_X1 U5599 ( .A(n4541), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n4540), 
        .Z(n4543) );
  NOR2_X1 U5600 ( .A1(n4543), .A2(n4542), .ZN(n4544) );
  NAND2_X1 U5601 ( .A1(n4562), .A2(n4544), .ZN(n4549) );
  INV_X1 U5602 ( .A(n4559), .ZN(n4547) );
  INV_X1 U5603 ( .A(n4540), .ZN(n5336) );
  AOI21_X1 U5604 ( .B1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n5336), .A(n4545), 
        .ZN(n4546) );
  NAND2_X1 U5605 ( .A1(n3423), .A2(n4546), .ZN(n5973) );
  NAND2_X1 U5606 ( .A1(n4547), .A2(n5973), .ZN(n4548) );
  OAI211_X1 U5607 ( .C1(n4551), .C2(n4550), .A(n4549), .B(n4548), .ZN(n4552)
         );
  AOI21_X1 U5608 ( .B1(n6430), .B2(n4553), .A(n4552), .ZN(n5976) );
  INV_X1 U5609 ( .A(n4612), .ZN(n4565) );
  MUX2_X1 U5610 ( .A(n4554), .B(n5976), .S(n4565), .Z(n4619) );
  INV_X1 U5611 ( .A(n4619), .ZN(n4566) );
  XNOR2_X1 U5612 ( .A(n4540), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4561)
         );
  XNOR2_X1 U5613 ( .A(n2972), .B(n4556), .ZN(n4557) );
  NAND2_X1 U5614 ( .A1(n4650), .A2(n4557), .ZN(n4558) );
  OAI21_X1 U5615 ( .B1(n4561), .B2(n4559), .A(n4558), .ZN(n4560) );
  AOI21_X1 U5616 ( .B1(n4562), .B2(n4561), .A(n4560), .ZN(n4563) );
  OAI21_X1 U5617 ( .B1(n4555), .B2(n4564), .A(n4563), .ZN(n5335) );
  MUX2_X1 U5618 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n5335), .S(n4565), 
        .Z(n4616) );
  NAND3_X1 U5619 ( .A1(n4566), .A2(n4629), .A3(n4616), .ZN(n4569) );
  NAND2_X1 U5620 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6093), .ZN(n4575) );
  INV_X1 U5621 ( .A(n4575), .ZN(n4567) );
  NAND2_X1 U5622 ( .A1(n4542), .A2(n4567), .ZN(n4568) );
  NAND2_X1 U5623 ( .A1(n4569), .A2(n4568), .ZN(n4626) );
  INV_X1 U5624 ( .A(n4570), .ZN(n4571) );
  NAND2_X1 U5625 ( .A1(n4626), .A2(n4571), .ZN(n4584) );
  NAND2_X1 U5626 ( .A1(n6214), .A2(n4572), .ZN(n4574) );
  NAND2_X1 U5627 ( .A1(n4612), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4573) );
  NAND2_X1 U5628 ( .A1(n4574), .A2(n4573), .ZN(n4577) );
  NOR2_X1 U5629 ( .A1(n4575), .A2(n4475), .ZN(n4576) );
  AOI21_X1 U5630 ( .B1(n4577), .B2(n4629), .A(n4576), .ZN(n4624) );
  NAND3_X1 U5631 ( .A1(n4584), .A2(n4624), .A3(n6093), .ZN(n4579) );
  NAND2_X1 U5632 ( .A1(n4579), .A2(n4578), .ZN(n4583) );
  INV_X1 U5633 ( .A(n6683), .ZN(n6604) );
  NAND2_X1 U5634 ( .A1(n6604), .A2(n4580), .ZN(n4581) );
  NAND2_X1 U5635 ( .A1(n4583), .A2(n5017), .ZN(n6408) );
  NAND3_X1 U5636 ( .A1(n4584), .A2(n4653), .A3(n4624), .ZN(n6597) );
  INV_X1 U5637 ( .A(n6597), .ZN(n4586) );
  NOR2_X1 U5638 ( .A1(n4629), .A2(STATE2_REG_3__SCAN_IN), .ZN(n5970) );
  OAI22_X1 U5639 ( .A1(n5986), .A2(n6428), .B1(n5970), .B2(n5541), .ZN(n4585)
         );
  OAI21_X1 U5640 ( .B1(n4586), .B2(n4585), .A(n6408), .ZN(n4587) );
  OAI21_X1 U5641 ( .B1(n6408), .B2(n6033), .A(n4587), .ZN(U3465) );
  XNOR2_X1 U5642 ( .A(n2971), .B(n4589), .ZN(n4682) );
  INV_X1 U5643 ( .A(n6392), .ZN(n5071) );
  AOI21_X1 U5644 ( .B1(n5892), .B2(n6390), .A(n5070), .ZN(n6407) );
  OAI21_X1 U5645 ( .B1(n5071), .B2(n6388), .A(n6407), .ZN(n4646) );
  INV_X1 U5646 ( .A(n6388), .ZN(n4591) );
  INV_X1 U5647 ( .A(n6390), .ZN(n4590) );
  AOI21_X1 U5648 ( .B1(n4590), .B2(n6402), .A(n6392), .ZN(n5068) );
  NOR2_X1 U5649 ( .A1(n4591), .A2(n5068), .ZN(n4639) );
  AOI22_X1 U5650 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n4646), .B1(n4639), 
        .B2(n4592), .ZN(n4598) );
  INV_X1 U5651 ( .A(n4594), .ZN(n4606) );
  OAI21_X1 U5652 ( .B1(n4607), .B2(n4606), .A(n4595), .ZN(n4596) );
  AND2_X1 U5653 ( .A1(n4596), .A2(n4642), .ZN(n6231) );
  INV_X1 U5654 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6614) );
  NOR2_X1 U5655 ( .A1(n6398), .A2(n6614), .ZN(n4677) );
  AOI21_X1 U5656 ( .B1(n6395), .B2(n6231), .A(n4677), .ZN(n4597) );
  OAI211_X1 U5657 ( .C1(n4682), .C2(n5961), .A(n4598), .B(n4597), .ZN(U3015)
         );
  NAND2_X1 U5658 ( .A1(n4599), .A2(n4600), .ZN(n4729) );
  OR2_X1 U5659 ( .A1(n4599), .A2(n4600), .ZN(n4601) );
  NAND2_X1 U5660 ( .A1(n4729), .A2(n4601), .ZN(n6238) );
  AOI22_X1 U5661 ( .A1(n6247), .A2(n6231), .B1(EBX_REG_3__SCAN_IN), .B2(n5595), 
        .ZN(n4602) );
  OAI21_X1 U5662 ( .B1(n6238), .B2(n5590), .A(n4602), .ZN(U2856) );
  INV_X1 U5663 ( .A(DATAI_1_), .ZN(n4704) );
  INV_X1 U5664 ( .A(EAX_REG_1__SCAN_IN), .ZN(n6318) );
  OAI222_X1 U5665 ( .A1(n5540), .A2(n5635), .B1(n4844), .B2(n4704), .C1(n6261), 
        .C2(n6318), .ZN(U2890) );
  INV_X1 U5666 ( .A(n4599), .ZN(n4603) );
  OAI21_X1 U5667 ( .B1(n4605), .B2(n4604), .A(n4603), .ZN(n6352) );
  INV_X1 U5668 ( .A(DATAI_2_), .ZN(n4687) );
  INV_X1 U5669 ( .A(EAX_REG_2__SCAN_IN), .ZN(n6321) );
  OAI222_X1 U5670 ( .A1(n6352), .A2(n5635), .B1(n4844), .B2(n4687), .C1(n6261), 
        .C2(n6321), .ZN(U2889) );
  INV_X1 U5671 ( .A(DATAI_3_), .ZN(n6720) );
  INV_X1 U5672 ( .A(EAX_REG_3__SCAN_IN), .ZN(n6324) );
  OAI222_X1 U5673 ( .A1(n6238), .A2(n5635), .B1(n4844), .B2(n6720), .C1(n6261), 
        .C2(n6324), .ZN(U2888) );
  INV_X1 U5674 ( .A(EBX_REG_2__SCAN_IN), .ZN(n4608) );
  XNOR2_X1 U5675 ( .A(n4607), .B(n4606), .ZN(n6393) );
  OAI222_X1 U5676 ( .A1(n5597), .A2(n6352), .B1(n4608), .B2(n6250), .C1(n5588), 
        .C2(n6393), .ZN(U2857) );
  NOR3_X1 U5677 ( .A1(n4610), .A2(n4609), .A3(n6033), .ZN(n4613) );
  NOR2_X1 U5678 ( .A1(n4613), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4615)
         );
  AOI211_X1 U5679 ( .C1(n4613), .C2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(n4612), .B(n4611), .ZN(n4614) );
  AOI211_X1 U5680 ( .C1(n5087), .C2(n4616), .A(n4615), .B(n4614), .ZN(n4618)
         );
  NOR2_X1 U5681 ( .A1(n4616), .A2(n5087), .ZN(n4617) );
  OAI22_X1 U5682 ( .A1(n4618), .A2(n4617), .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n4619), .ZN(n4628) );
  AOI21_X1 U5683 ( .B1(n4619), .B2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n4627) );
  OAI21_X1 U5684 ( .B1(FLUSH_REG_SCAN_IN), .B2(MORE_REG_SCAN_IN), .A(n4620), 
        .ZN(n4621) );
  NAND4_X1 U5685 ( .A1(n4624), .A2(n4623), .A3(n4622), .A4(n4621), .ZN(n4625)
         );
  AOI211_X1 U5686 ( .C1(n4628), .C2(n4627), .A(n4626), .B(n4625), .ZN(n6609)
         );
  AOI21_X1 U5687 ( .B1(n6609), .B2(n4629), .A(n6603), .ZN(n4633) );
  NOR2_X1 U5688 ( .A1(READY_N), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5274) );
  NAND2_X1 U5689 ( .A1(n4630), .A2(n5274), .ZN(n5272) );
  AOI21_X1 U5690 ( .B1(STATE2_REG_1__SCAN_IN), .B2(READY_N), .A(
        STATE2_REG_0__SCAN_IN), .ZN(n4631) );
  INV_X1 U5691 ( .A(n4631), .ZN(n4632) );
  OAI211_X1 U5692 ( .C1(n4648), .C2(n5272), .A(STATE2_REG_2__SCAN_IN), .B(
        n4632), .ZN(n6602) );
  NOR2_X1 U5693 ( .A1(n4633), .A2(n6602), .ZN(n4660) );
  OAI21_X1 U5694 ( .B1(n4660), .B2(n6603), .A(STATE2_REG_3__SCAN_IN), .ZN(
        n4635) );
  NAND2_X1 U5695 ( .A1(n4635), .A2(n4634), .ZN(U3453) );
  XNOR2_X1 U5696 ( .A(n4636), .B(n4637), .ZN(n4802) );
  OAI211_X1 U5697 ( .C1(INSTADDRPOINTER_REG_3__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A(n4639), .B(n4638), .ZN(n4640) );
  INV_X1 U5698 ( .A(n4640), .ZN(n4645) );
  AND2_X1 U5699 ( .A1(n4642), .A2(n4641), .ZN(n4643) );
  OR2_X1 U5700 ( .A1(n4643), .A2(n4737), .ZN(n6228) );
  OAI22_X1 U5701 ( .A1(n6382), .A2(n6228), .B1(n6616), .B2(n6398), .ZN(n4644)
         );
  AOI211_X1 U5702 ( .C1(n4646), .C2(INSTADDRPOINTER_REG_4__SCAN_IN), .A(n4645), 
        .B(n4644), .ZN(n4647) );
  OAI21_X1 U5703 ( .B1(n5961), .B2(n4802), .A(n4647), .ZN(U3014) );
  INV_X1 U5704 ( .A(DATAO_REG_24__SCAN_IN), .ZN(n4656) );
  INV_X1 U5705 ( .A(n4648), .ZN(n4649) );
  NOR2_X2 U5706 ( .A1(n6288), .A2(n4709), .ZN(n6263) );
  INV_X1 U5707 ( .A(n6263), .ZN(n4655) );
  INV_X1 U5708 ( .A(EAX_REG_24__SCAN_IN), .ZN(n6736) );
  INV_X1 U5709 ( .A(UWORD_REG_8__SCAN_IN), .ZN(n4654) );
  OAI222_X1 U5710 ( .A1(n4656), .A2(n6281), .B1(n4655), .B2(n6736), .C1(n6280), 
        .C2(n4654), .ZN(U2899) );
  NOR2_X1 U5711 ( .A1(n4660), .A2(n4657), .ZN(n6598) );
  NAND2_X1 U5712 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n4658), .ZN(n4665) );
  NOR3_X1 U5713 ( .A1(n5975), .A2(READY_N), .A3(n6603), .ZN(n4662) );
  INV_X1 U5714 ( .A(n4660), .ZN(n4661) );
  OAI21_X1 U5715 ( .B1(n4663), .B2(n4662), .A(n4661), .ZN(n4664) );
  OAI211_X1 U5716 ( .C1(n6598), .C2(n4665), .A(n5237), .B(n4664), .ZN(U3149)
         );
  AOI222_X1 U5717 ( .A1(EAX_REG_30__SCAN_IN), .A2(n6263), .B1(n6286), .B2(
        DATAO_REG_30__SCAN_IN), .C1(n6681), .C2(UWORD_REG_14__SCAN_IN), .ZN(
        n4666) );
  INV_X1 U5718 ( .A(n4666), .ZN(U2893) );
  AOI222_X1 U5719 ( .A1(EAX_REG_16__SCAN_IN), .A2(n6263), .B1(n6286), .B2(
        DATAO_REG_16__SCAN_IN), .C1(n6681), .C2(UWORD_REG_0__SCAN_IN), .ZN(
        n4667) );
  INV_X1 U5720 ( .A(n4667), .ZN(U2907) );
  AOI222_X1 U5721 ( .A1(EAX_REG_17__SCAN_IN), .A2(n6263), .B1(n6286), .B2(
        DATAO_REG_17__SCAN_IN), .C1(n6681), .C2(UWORD_REG_1__SCAN_IN), .ZN(
        n4668) );
  INV_X1 U5722 ( .A(n4668), .ZN(U2906) );
  AOI222_X1 U5723 ( .A1(EAX_REG_27__SCAN_IN), .A2(n6263), .B1(n6286), .B2(
        DATAO_REG_27__SCAN_IN), .C1(n6681), .C2(UWORD_REG_11__SCAN_IN), .ZN(
        n4669) );
  INV_X1 U5724 ( .A(n4669), .ZN(U2896) );
  AOI222_X1 U5725 ( .A1(EAX_REG_26__SCAN_IN), .A2(n6263), .B1(n6286), .B2(
        DATAO_REG_26__SCAN_IN), .C1(n6681), .C2(UWORD_REG_10__SCAN_IN), .ZN(
        n4670) );
  INV_X1 U5726 ( .A(n4670), .ZN(U2897) );
  AOI222_X1 U5727 ( .A1(EAX_REG_23__SCAN_IN), .A2(n6263), .B1(n6286), .B2(
        DATAO_REG_23__SCAN_IN), .C1(n6681), .C2(UWORD_REG_7__SCAN_IN), .ZN(
        n4671) );
  INV_X1 U5728 ( .A(n4671), .ZN(U2900) );
  AOI222_X1 U5729 ( .A1(EAX_REG_22__SCAN_IN), .A2(n6263), .B1(n6286), .B2(
        DATAO_REG_22__SCAN_IN), .C1(n6681), .C2(UWORD_REG_6__SCAN_IN), .ZN(
        n4672) );
  INV_X1 U5730 ( .A(n4672), .ZN(U2901) );
  AOI222_X1 U5731 ( .A1(EAX_REG_29__SCAN_IN), .A2(n6263), .B1(n6286), .B2(
        DATAO_REG_29__SCAN_IN), .C1(n6681), .C2(UWORD_REG_13__SCAN_IN), .ZN(
        n4673) );
  INV_X1 U5732 ( .A(n4673), .ZN(U2894) );
  AOI222_X1 U5733 ( .A1(EAX_REG_28__SCAN_IN), .A2(n6263), .B1(n6286), .B2(
        DATAO_REG_28__SCAN_IN), .C1(n6681), .C2(UWORD_REG_12__SCAN_IN), .ZN(
        n4674) );
  INV_X1 U5734 ( .A(n4674), .ZN(U2895) );
  AOI222_X1 U5735 ( .A1(EAX_REG_20__SCAN_IN), .A2(n6263), .B1(n6286), .B2(
        DATAO_REG_20__SCAN_IN), .C1(n6681), .C2(UWORD_REG_4__SCAN_IN), .ZN(
        n4675) );
  INV_X1 U5736 ( .A(n4675), .ZN(U2903) );
  AOI222_X1 U5737 ( .A1(EAX_REG_19__SCAN_IN), .A2(n6263), .B1(n6286), .B2(
        DATAO_REG_19__SCAN_IN), .C1(n6681), .C2(UWORD_REG_3__SCAN_IN), .ZN(
        n4676) );
  INV_X1 U5738 ( .A(n4676), .ZN(U2904) );
  INV_X1 U5739 ( .A(n6238), .ZN(n4680) );
  AOI21_X1 U5740 ( .B1(n6351), .B2(PHYADDRPOINTER_REG_3__SCAN_IN), .A(n4677), 
        .ZN(n4678) );
  OAI21_X1 U5741 ( .B1(n6237), .B2(n6362), .A(n4678), .ZN(n4679) );
  AOI21_X1 U5742 ( .B1(n4680), .B2(n6358), .A(n4679), .ZN(n4681) );
  OAI21_X1 U5743 ( .B1(n4682), .B2(n6092), .A(n4681), .ZN(U2983) );
  INV_X1 U5744 ( .A(n4683), .ZN(n4684) );
  INV_X1 U5745 ( .A(n5980), .ZN(n4686) );
  NAND2_X1 U5746 ( .A1(n2976), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6516) );
  NOR2_X1 U5747 ( .A1(n4686), .A2(n6516), .ZN(n4889) );
  NOR2_X1 U5748 ( .A1(n4889), .A2(n6428), .ZN(n4690) );
  INV_X1 U5749 ( .A(n4555), .ZN(n5527) );
  NAND2_X1 U5750 ( .A1(n5527), .A2(n4515), .ZN(n5015) );
  OR2_X1 U5751 ( .A1(n5015), .A2(n5982), .ZN(n6030) );
  OAI21_X1 U5752 ( .B1(n6030), .B2(n5541), .A(n4721), .ZN(n4688) );
  AND3_X1 U5753 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n3442), .ZN(n6032) );
  INV_X1 U5754 ( .A(n4688), .ZN(n4689) );
  NAND2_X1 U5755 ( .A1(n4690), .A2(n4689), .ZN(n4691) );
  NAND2_X1 U5756 ( .A1(n4719), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4695) );
  NAND2_X1 U5757 ( .A1(n6358), .A2(DATAI_18_), .ZN(n6540) );
  NAND3_X1 U5758 ( .A1(n5980), .A2(n2976), .A3(n5987), .ZN(n6511) );
  NAND3_X1 U5759 ( .A1(n5980), .A2(n5986), .A3(n2976), .ZN(n6462) );
  NAND2_X1 U5760 ( .A1(n6358), .A2(DATAI_26_), .ZN(n6545) );
  OR2_X1 U5761 ( .A1(n4720), .A2(n4692), .ZN(n6539) );
  OAI22_X1 U5762 ( .A1(n6462), .A2(n6545), .B1(n4721), .B2(n6539), .ZN(n4693)
         );
  AOI21_X1 U5763 ( .B1(n6486), .B2(n6471), .A(n4693), .ZN(n4694) );
  OAI211_X1 U5764 ( .C1(n4725), .C2(n6005), .A(n4695), .B(n4694), .ZN(U3078)
         );
  INV_X1 U5765 ( .A(DATAI_6_), .ZN(n4843) );
  NAND2_X1 U5766 ( .A1(n4719), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4698) );
  NAND2_X1 U5767 ( .A1(n6358), .A2(DATAI_22_), .ZN(n6568) );
  OAI22_X1 U5768 ( .A1(n6462), .A2(n6854), .B1(n4721), .B2(n6567), .ZN(n4696)
         );
  AOI21_X1 U5769 ( .B1(n6849), .B2(n6471), .A(n4696), .ZN(n4697) );
  OAI211_X1 U5770 ( .C1(n4725), .C2(n6021), .A(n4698), .B(n4697), .ZN(U3082)
         );
  NAND2_X1 U5771 ( .A1(n4719), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4703) );
  NAND2_X1 U5772 ( .A1(n6358), .A2(DATAI_23_), .ZN(n6582) );
  NAND2_X1 U5773 ( .A1(n6358), .A2(DATAI_31_), .ZN(n6574) );
  OAI22_X1 U5774 ( .A1(n6462), .A2(n6574), .B1(n4721), .B2(n6573), .ZN(n4701)
         );
  AOI21_X1 U5775 ( .B1(n6507), .B2(n6471), .A(n4701), .ZN(n4702) );
  OAI211_X1 U5776 ( .C1(n4725), .C2(n6027), .A(n4703), .B(n4702), .ZN(U3083)
         );
  NAND2_X1 U5777 ( .A1(n4719), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4707) );
  NAND2_X1 U5778 ( .A1(n6358), .A2(DATAI_17_), .ZN(n6538) );
  NAND2_X1 U5779 ( .A1(n6358), .A2(DATAI_25_), .ZN(n6589) );
  OAI22_X1 U5780 ( .A1(n6462), .A2(n6589), .B1(n4721), .B2(n6534), .ZN(n4705)
         );
  AOI21_X1 U5781 ( .B1(n6586), .B2(n6471), .A(n4705), .ZN(n4706) );
  OAI211_X1 U5782 ( .C1(n4725), .C2(n6001), .A(n4707), .B(n4706), .ZN(U3077)
         );
  NAND2_X1 U5783 ( .A1(n4719), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4712) );
  NAND2_X1 U5784 ( .A1(n6358), .A2(DATAI_16_), .ZN(n6513) );
  NAND2_X1 U5785 ( .A1(n6358), .A2(DATAI_24_), .ZN(n6533) );
  OR2_X1 U5786 ( .A1(n4720), .A2(n4709), .ZN(n6512) );
  OAI22_X1 U5787 ( .A1(n6462), .A2(n6533), .B1(n4721), .B2(n6512), .ZN(n4710)
         );
  AOI21_X1 U5788 ( .B1(n6480), .B2(n6471), .A(n4710), .ZN(n4711) );
  OAI211_X1 U5789 ( .C1(n4725), .C2(n5997), .A(n4712), .B(n4711), .ZN(U3076)
         );
  INV_X1 U5790 ( .A(DATAI_5_), .ZN(n4841) );
  NAND2_X1 U5791 ( .A1(n4719), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4715) );
  NAND2_X1 U5792 ( .A1(n6358), .A2(DATAI_21_), .ZN(n6561) );
  NAND2_X1 U5793 ( .A1(n6358), .A2(DATAI_29_), .ZN(n6566) );
  OR2_X1 U5794 ( .A1(n4720), .A2(n3348), .ZN(n6560) );
  OAI22_X1 U5795 ( .A1(n6462), .A2(n6566), .B1(n4721), .B2(n6560), .ZN(n4713)
         );
  AOI21_X1 U5796 ( .B1(n6498), .B2(n6471), .A(n4713), .ZN(n4714) );
  OAI211_X1 U5797 ( .C1(n4725), .C2(n6017), .A(n4715), .B(n4714), .ZN(U3081)
         );
  INV_X1 U5798 ( .A(DATAI_4_), .ZN(n4733) );
  NAND2_X1 U5799 ( .A1(n4719), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4718) );
  NAND2_X1 U5800 ( .A1(n6358), .A2(DATAI_20_), .ZN(n6559) );
  NAND2_X1 U5801 ( .A1(n6358), .A2(DATAI_28_), .ZN(n6554) );
  OR2_X1 U5802 ( .A1(n4720), .A2(n3320), .ZN(n6553) );
  OAI22_X1 U5803 ( .A1(n6462), .A2(n6554), .B1(n4721), .B2(n6553), .ZN(n4716)
         );
  AOI21_X1 U5804 ( .B1(n6494), .B2(n6471), .A(n4716), .ZN(n4717) );
  OAI211_X1 U5805 ( .C1(n4725), .C2(n6013), .A(n4718), .B(n4717), .ZN(U3080)
         );
  NAND2_X1 U5806 ( .A1(n4719), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4724) );
  NAND2_X1 U5807 ( .A1(n6358), .A2(DATAI_19_), .ZN(n6547) );
  NAND2_X1 U5808 ( .A1(n6358), .A2(DATAI_27_), .ZN(n6552) );
  OR2_X1 U5809 ( .A1(n4720), .A2(n3321), .ZN(n6546) );
  OAI22_X1 U5810 ( .A1(n6462), .A2(n6552), .B1(n4721), .B2(n6546), .ZN(n4722)
         );
  AOI21_X1 U5811 ( .B1(n6490), .B2(n6471), .A(n4722), .ZN(n4723) );
  OAI211_X1 U5812 ( .C1(n4725), .C2(n6009), .A(n4724), .B(n4723), .ZN(U3079)
         );
  AOI222_X1 U5813 ( .A1(n6286), .A2(DATAO_REG_21__SCAN_IN), .B1(n6263), .B2(
        EAX_REG_21__SCAN_IN), .C1(n6681), .C2(UWORD_REG_5__SCAN_IN), .ZN(n4726) );
  INV_X1 U5814 ( .A(n4726), .ZN(U2902) );
  INV_X1 U5815 ( .A(n4727), .ZN(n4728) );
  NOR2_X1 U5816 ( .A1(n4729), .A2(n4728), .ZN(n4830) );
  AND2_X1 U5817 ( .A1(n4729), .A2(n4728), .ZN(n4730) );
  INV_X1 U5818 ( .A(n6228), .ZN(n4731) );
  AOI22_X1 U5819 ( .A1(n6247), .A2(n4731), .B1(EBX_REG_4__SCAN_IN), .B2(n5595), 
        .ZN(n4732) );
  OAI21_X1 U5820 ( .B1(n6222), .B2(n5590), .A(n4732), .ZN(U2855) );
  INV_X1 U5821 ( .A(EAX_REG_4__SCAN_IN), .ZN(n6327) );
  OAI222_X1 U5822 ( .A1(n6222), .A2(n5635), .B1(n4844), .B2(n4733), .C1(n6261), 
        .C2(n6327), .ZN(U2887) );
  XNOR2_X1 U5823 ( .A(n4734), .B(n4735), .ZN(n4838) );
  OAI21_X1 U5824 ( .B1(n5955), .B2(n4848), .A(n6407), .ZN(n4849) );
  OAI21_X1 U5825 ( .B1(n5071), .B2(n4736), .A(n4740), .ZN(n4744) );
  AOI21_X1 U5826 ( .B1(n4739), .B2(n3131), .A(n4795), .ZN(n6201) );
  INV_X1 U5827 ( .A(n6201), .ZN(n4839) );
  NAND3_X1 U5828 ( .A1(n4741), .A2(n6402), .A3(n4740), .ZN(n4742) );
  INV_X1 U5829 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6734) );
  OR2_X1 U5830 ( .A1(n6734), .A2(n6398), .ZN(n4835) );
  OAI211_X1 U5831 ( .C1(n6382), .C2(n4839), .A(n4742), .B(n4835), .ZN(n4743)
         );
  AOI21_X1 U5832 ( .B1(n4849), .B2(n4744), .A(n4743), .ZN(n4745) );
  OAI21_X1 U5833 ( .B1(n5961), .B2(n4838), .A(n4745), .ZN(U3013) );
  NOR2_X1 U5834 ( .A1(n5966), .A2(n4683), .ZN(n4803) );
  INV_X1 U5835 ( .A(n4751), .ZN(n4746) );
  NAND2_X1 U5836 ( .A1(n6524), .A2(n6091), .ZN(n6433) );
  INV_X1 U5837 ( .A(n6433), .ZN(n4976) );
  AOI21_X1 U5838 ( .B1(n4746), .B2(n6358), .A(n4976), .ZN(n4750) );
  INV_X1 U5839 ( .A(n5015), .ZN(n6038) );
  AND2_X1 U5840 ( .A1(n6430), .A2(n6519), .ZN(n5166) );
  NAND2_X1 U5841 ( .A1(n6038), .A2(n5166), .ZN(n4748) );
  NAND2_X1 U5842 ( .A1(n4747), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4787) );
  NAND2_X1 U5843 ( .A1(n4748), .A2(n4787), .ZN(n4752) );
  NAND3_X1 U5844 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n5016) );
  NAND2_X1 U5845 ( .A1(n6428), .A2(n5016), .ZN(n4749) );
  NAND2_X1 U5846 ( .A1(n4784), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4759)
         );
  INV_X1 U5847 ( .A(n6552), .ZN(n6054) );
  NAND2_X1 U5848 ( .A1(n4752), .A2(n6524), .ZN(n4755) );
  INV_X1 U5849 ( .A(n5016), .ZN(n4753) );
  NAND2_X1 U5850 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n4753), .ZN(n4754) );
  NAND2_X1 U5851 ( .A1(n4755), .A2(n4754), .ZN(n4785) );
  NAND2_X1 U5852 ( .A1(n4785), .A2(n6549), .ZN(n4756) );
  OAI21_X1 U5853 ( .B1(n4787), .B2(n6546), .A(n4756), .ZN(n4757) );
  AOI21_X1 U5854 ( .B1(n5057), .B2(n6054), .A(n4757), .ZN(n4758) );
  OAI211_X1 U5855 ( .C1(n4952), .C2(n6547), .A(n4759), .B(n4758), .ZN(U3143)
         );
  NAND2_X1 U5856 ( .A1(n4784), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4763)
         );
  INV_X1 U5857 ( .A(n6545), .ZN(n6411) );
  NAND2_X1 U5858 ( .A1(n4785), .A2(n6542), .ZN(n4760) );
  OAI21_X1 U5859 ( .B1(n4787), .B2(n6539), .A(n4760), .ZN(n4761) );
  AOI21_X1 U5860 ( .B1(n5057), .B2(n6411), .A(n4761), .ZN(n4762) );
  OAI211_X1 U5861 ( .C1(n4952), .C2(n6540), .A(n4763), .B(n4762), .ZN(U3142)
         );
  NAND2_X1 U5862 ( .A1(n4784), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4767)
         );
  INV_X1 U5863 ( .A(n6589), .ZN(n6045) );
  NAND2_X1 U5864 ( .A1(n4785), .A2(n6585), .ZN(n4764) );
  OAI21_X1 U5865 ( .B1(n4787), .B2(n6534), .A(n4764), .ZN(n4765) );
  AOI21_X1 U5866 ( .B1(n5057), .B2(n6045), .A(n4765), .ZN(n4766) );
  OAI211_X1 U5867 ( .C1(n4952), .C2(n6538), .A(n4767), .B(n4766), .ZN(U3141)
         );
  NAND2_X1 U5868 ( .A1(n4784), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4771)
         );
  INV_X1 U5869 ( .A(n6574), .ZN(n6421) );
  NAND2_X1 U5870 ( .A1(n4785), .A2(n6578), .ZN(n4768) );
  OAI21_X1 U5871 ( .B1(n4787), .B2(n6573), .A(n4768), .ZN(n4769) );
  AOI21_X1 U5872 ( .B1(n5057), .B2(n6421), .A(n4769), .ZN(n4770) );
  OAI211_X1 U5873 ( .C1(n4952), .C2(n6582), .A(n4771), .B(n4770), .ZN(U3147)
         );
  NAND2_X1 U5874 ( .A1(n4784), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4775)
         );
  INV_X1 U5875 ( .A(n6854), .ZN(n6067) );
  NAND2_X1 U5876 ( .A1(n4785), .A2(n6846), .ZN(n4772) );
  OAI21_X1 U5877 ( .B1(n4787), .B2(n6567), .A(n4772), .ZN(n4773) );
  AOI21_X1 U5878 ( .B1(n5057), .B2(n6067), .A(n4773), .ZN(n4774) );
  OAI211_X1 U5879 ( .C1(n4952), .C2(n6568), .A(n4775), .B(n4774), .ZN(U3146)
         );
  NAND2_X1 U5880 ( .A1(n4784), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4779)
         );
  INV_X1 U5881 ( .A(n6566), .ZN(n6417) );
  NAND2_X1 U5882 ( .A1(n4785), .A2(n6563), .ZN(n4776) );
  OAI21_X1 U5883 ( .B1(n4787), .B2(n6560), .A(n4776), .ZN(n4777) );
  AOI21_X1 U5884 ( .B1(n5057), .B2(n6417), .A(n4777), .ZN(n4778) );
  OAI211_X1 U5885 ( .C1(n4952), .C2(n6561), .A(n4779), .B(n4778), .ZN(U3145)
         );
  NAND2_X1 U5886 ( .A1(n4784), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4783)
         );
  INV_X1 U5887 ( .A(n6554), .ZN(n6414) );
  NAND2_X1 U5888 ( .A1(n4785), .A2(n6556), .ZN(n4780) );
  OAI21_X1 U5889 ( .B1(n4787), .B2(n6553), .A(n4780), .ZN(n4781) );
  AOI21_X1 U5890 ( .B1(n5057), .B2(n6414), .A(n4781), .ZN(n4782) );
  OAI211_X1 U5891 ( .C1(n4952), .C2(n6559), .A(n4783), .B(n4782), .ZN(U3144)
         );
  NAND2_X1 U5892 ( .A1(n4784), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4790)
         );
  INV_X1 U5893 ( .A(n6533), .ZN(n6458) );
  NAND2_X1 U5894 ( .A1(n4785), .A2(n6530), .ZN(n4786) );
  OAI21_X1 U5895 ( .B1(n4787), .B2(n6512), .A(n4786), .ZN(n4788) );
  AOI21_X1 U5896 ( .B1(n5057), .B2(n6458), .A(n4788), .ZN(n4789) );
  OAI211_X1 U5897 ( .C1(n4952), .C2(n6513), .A(n4790), .B(n4789), .ZN(U3140)
         );
  AND2_X1 U5898 ( .A1(n4830), .A2(n4829), .ZN(n4831) );
  OAI21_X1 U5899 ( .B1(n4831), .B2(n4792), .A(n4791), .ZN(n5520) );
  OAI21_X1 U5900 ( .B1(n4795), .B2(n4794), .A(n4793), .ZN(n4796) );
  INV_X1 U5901 ( .A(n4796), .ZN(n5512) );
  AOI22_X1 U5902 ( .A1(n6247), .A2(n5512), .B1(EBX_REG_6__SCAN_IN), .B2(n5595), 
        .ZN(n4797) );
  OAI21_X1 U5903 ( .B1(n5520), .B2(n5590), .A(n4797), .ZN(U2853) );
  INV_X1 U5904 ( .A(n6222), .ZN(n4800) );
  AOI22_X1 U5905 ( .A1(n6351), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .B1(n6350), 
        .B2(REIP_REG_4__SCAN_IN), .ZN(n4798) );
  OAI21_X1 U5906 ( .B1(n6221), .B2(n6362), .A(n4798), .ZN(n4799) );
  AOI21_X1 U5907 ( .B1(n4800), .B2(n6358), .A(n4799), .ZN(n4801) );
  OAI21_X1 U5908 ( .B1(n6092), .B2(n4802), .A(n4801), .ZN(U2982) );
  NAND2_X1 U5909 ( .A1(n4803), .A2(n5979), .ZN(n4809) );
  INV_X1 U5910 ( .A(n4515), .ZN(n5964) );
  NAND2_X1 U5911 ( .A1(n5527), .A2(n5964), .ZN(n6429) );
  INV_X1 U5912 ( .A(n6429), .ZN(n4983) );
  NAND3_X1 U5913 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n5983), .ZN(n4978) );
  NOR2_X1 U5914 ( .A1(n6033), .A2(n4978), .ZN(n4826) );
  AOI21_X1 U5915 ( .B1(n4983), .B2(n5166), .A(n4826), .ZN(n4808) );
  INV_X1 U5916 ( .A(n4808), .ZN(n4806) );
  INV_X1 U5917 ( .A(n4809), .ZN(n4804) );
  NAND2_X1 U5918 ( .A1(n4804), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4888) );
  NAND2_X1 U5919 ( .A1(n6524), .A2(n4888), .ZN(n4807) );
  NAND2_X1 U5920 ( .A1(n6428), .A2(n4978), .ZN(n4805) );
  OAI211_X1 U5921 ( .C1(n4806), .C2(n4807), .A(n6522), .B(n4805), .ZN(n4825)
         );
  OAI22_X1 U5922 ( .A1(n4808), .A2(n4807), .B1(n6527), .B2(n4978), .ZN(n4824)
         );
  AOI22_X1 U5923 ( .A1(INSTQUEUE_REG_13__6__SCAN_IN), .A2(n4825), .B1(n6846), 
        .B2(n4824), .ZN(n4811) );
  AOI22_X1 U5924 ( .A1(n6592), .A2(n6067), .B1(n4826), .B2(n6845), .ZN(n4810)
         );
  OAI211_X1 U5925 ( .C1(n5055), .C2(n6568), .A(n4811), .B(n4810), .ZN(U3130)
         );
  AOI22_X1 U5926 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n4825), .B1(n6578), 
        .B2(n4824), .ZN(n4813) );
  AOI22_X1 U5927 ( .A1(n6592), .A2(n6421), .B1(n4826), .B2(n6504), .ZN(n4812)
         );
  OAI211_X1 U5928 ( .C1(n5055), .C2(n6582), .A(n4813), .B(n4812), .ZN(U3131)
         );
  AOI22_X1 U5929 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(n4825), .B1(n6563), 
        .B2(n4824), .ZN(n4815) );
  AOI22_X1 U5930 ( .A1(n6592), .A2(n6417), .B1(n4826), .B2(n6497), .ZN(n4814)
         );
  OAI211_X1 U5931 ( .C1(n5055), .C2(n6561), .A(n4815), .B(n4814), .ZN(U3129)
         );
  AOI22_X1 U5932 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n4825), .B1(n6556), 
        .B2(n4824), .ZN(n4817) );
  AOI22_X1 U5933 ( .A1(n6592), .A2(n6414), .B1(n4826), .B2(n6493), .ZN(n4816)
         );
  OAI211_X1 U5934 ( .C1(n5055), .C2(n6559), .A(n4817), .B(n4816), .ZN(U3128)
         );
  AOI22_X1 U5935 ( .A1(INSTQUEUE_REG_13__2__SCAN_IN), .A2(n4825), .B1(n6542), 
        .B2(n4824), .ZN(n4819) );
  AOI22_X1 U5936 ( .A1(n6592), .A2(n6411), .B1(n4826), .B2(n6485), .ZN(n4818)
         );
  OAI211_X1 U5937 ( .C1(n5055), .C2(n6540), .A(n4819), .B(n4818), .ZN(U3126)
         );
  AOI22_X1 U5938 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n4825), .B1(n6585), 
        .B2(n4824), .ZN(n4821) );
  AOI22_X1 U5939 ( .A1(n6592), .A2(n6045), .B1(n4826), .B2(n6584), .ZN(n4820)
         );
  OAI211_X1 U5940 ( .C1(n5055), .C2(n6538), .A(n4821), .B(n4820), .ZN(U3125)
         );
  AOI22_X1 U5941 ( .A1(INSTQUEUE_REG_13__3__SCAN_IN), .A2(n4825), .B1(n6549), 
        .B2(n4824), .ZN(n4823) );
  AOI22_X1 U5942 ( .A1(n6592), .A2(n6054), .B1(n4826), .B2(n6489), .ZN(n4822)
         );
  OAI211_X1 U5943 ( .C1(n5055), .C2(n6547), .A(n4823), .B(n4822), .ZN(U3127)
         );
  AOI22_X1 U5944 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n4825), .B1(n6530), 
        .B2(n4824), .ZN(n4828) );
  AOI22_X1 U5945 ( .A1(n6592), .A2(n6458), .B1(n6470), .B2(n4826), .ZN(n4827)
         );
  OAI211_X1 U5946 ( .C1(n5055), .C2(n6513), .A(n4828), .B(n4827), .ZN(U3124)
         );
  INV_X1 U5947 ( .A(n4829), .ZN(n4833) );
  INV_X1 U5948 ( .A(n4830), .ZN(n4832) );
  AOI21_X1 U5949 ( .B1(n4833), .B2(n4832), .A(n4831), .ZN(n6206) );
  NAND2_X1 U5950 ( .A1(n6351), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n4834)
         );
  OAI211_X1 U5951 ( .C1(n6362), .C2(n6213), .A(n4835), .B(n4834), .ZN(n4836)
         );
  AOI21_X1 U5952 ( .B1(n6206), .B2(n6358), .A(n4836), .ZN(n4837) );
  OAI21_X1 U5953 ( .B1(n6092), .B2(n4838), .A(n4837), .ZN(U2981) );
  INV_X1 U5954 ( .A(n6206), .ZN(n4842) );
  INV_X1 U5955 ( .A(EBX_REG_5__SCAN_IN), .ZN(n4840) );
  OAI222_X1 U5956 ( .A1(n4842), .A2(n5590), .B1(n4840), .B2(n6250), .C1(n5588), 
        .C2(n4839), .ZN(U2854) );
  INV_X1 U5957 ( .A(EAX_REG_5__SCAN_IN), .ZN(n6826) );
  OAI222_X1 U5958 ( .A1(n4842), .A2(n5635), .B1(n4844), .B2(n4841), .C1(n6261), 
        .C2(n6826), .ZN(U2886) );
  OAI222_X1 U5959 ( .A1(n5520), .A2(n5635), .B1(n4844), .B2(n4843), .C1(n6261), 
        .C2(n3510), .ZN(U2885) );
  XNOR2_X1 U5960 ( .A(n4845), .B(n4846), .ZN(n4963) );
  NOR2_X1 U5961 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n5068), .ZN(n4847)
         );
  AOI22_X1 U5962 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n4849), .B1(n4848), 
        .B2(n4847), .ZN(n4852) );
  INV_X1 U5963 ( .A(REIP_REG_6__SCAN_IN), .ZN(n4850) );
  NOR2_X1 U5964 ( .A1(n6398), .A2(n4850), .ZN(n4958) );
  AOI21_X1 U5965 ( .B1(n6395), .B2(n5512), .A(n4958), .ZN(n4851) );
  OAI211_X1 U5966 ( .C1(n5961), .C2(n4963), .A(n4852), .B(n4851), .ZN(U3012)
         );
  INV_X1 U5967 ( .A(n5966), .ZN(n4853) );
  NAND2_X1 U5968 ( .A1(n4854), .A2(n2976), .ZN(n4900) );
  NOR2_X2 U5969 ( .A1(n4900), .A2(n5987), .ZN(n6422) );
  OAI21_X1 U5970 ( .B1(n6422), .B2(n5154), .A(n6433), .ZN(n4855) );
  AND2_X1 U5971 ( .A1(n4555), .A2(n4515), .ZN(n5083) );
  NAND2_X1 U5972 ( .A1(n6474), .A2(n5083), .ZN(n4893) );
  AOI21_X1 U5973 ( .B1(n4855), .B2(n4893), .A(STATE2_REG_3__SCAN_IN), .ZN(
        n4856) );
  NOR2_X1 U5974 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4918) );
  NAND2_X1 U5975 ( .A1(n4918), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4896) );
  NOR2_X1 U5976 ( .A1(n4896), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4859)
         );
  NAND2_X1 U5977 ( .A1(n6467), .A2(n3442), .ZN(n6039) );
  AOI21_X1 U5978 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6039), .A(n5017), .ZN(
        n6036) );
  NAND2_X1 U5979 ( .A1(n4881), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4862) );
  INV_X1 U5980 ( .A(n4893), .ZN(n4858) );
  INV_X1 U5981 ( .A(n6039), .ZN(n4857) );
  AOI22_X1 U5982 ( .A1(n4858), .A2(n6515), .B1(n6465), .B2(n4857), .ZN(n4883)
         );
  INV_X1 U5983 ( .A(n4859), .ZN(n4882) );
  OAI22_X1 U5984 ( .A1(n4883), .A2(n6017), .B1(n6560), .B2(n4882), .ZN(n4860)
         );
  AOI21_X1 U5985 ( .B1(n6422), .B2(n6498), .A(n4860), .ZN(n4861) );
  OAI211_X1 U5986 ( .C1(n4887), .C2(n6566), .A(n4862), .B(n4861), .ZN(U3041)
         );
  NAND2_X1 U5987 ( .A1(n4881), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4865) );
  OAI22_X1 U5988 ( .A1(n4883), .A2(n6013), .B1(n6553), .B2(n4882), .ZN(n4863)
         );
  AOI21_X1 U5989 ( .B1(n6422), .B2(n6494), .A(n4863), .ZN(n4864) );
  OAI211_X1 U5990 ( .C1(n4887), .C2(n6554), .A(n4865), .B(n4864), .ZN(U3040)
         );
  NAND2_X1 U5991 ( .A1(n4881), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4868) );
  OAI22_X1 U5992 ( .A1(n4883), .A2(n6009), .B1(n6546), .B2(n4882), .ZN(n4866)
         );
  AOI21_X1 U5993 ( .B1(n6422), .B2(n6490), .A(n4866), .ZN(n4867) );
  OAI211_X1 U5994 ( .C1(n4887), .C2(n6552), .A(n4868), .B(n4867), .ZN(U3039)
         );
  NAND2_X1 U5995 ( .A1(n4881), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4871) );
  OAI22_X1 U5996 ( .A1(n4883), .A2(n6005), .B1(n6539), .B2(n4882), .ZN(n4869)
         );
  AOI21_X1 U5997 ( .B1(n6422), .B2(n6486), .A(n4869), .ZN(n4870) );
  OAI211_X1 U5998 ( .C1(n4887), .C2(n6545), .A(n4871), .B(n4870), .ZN(U3038)
         );
  NAND2_X1 U5999 ( .A1(n4881), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4874) );
  OAI22_X1 U6000 ( .A1(n4883), .A2(n6001), .B1(n6534), .B2(n4882), .ZN(n4872)
         );
  AOI21_X1 U6001 ( .B1(n6422), .B2(n6586), .A(n4872), .ZN(n4873) );
  OAI211_X1 U6002 ( .C1(n4887), .C2(n6589), .A(n4874), .B(n4873), .ZN(U3037)
         );
  NAND2_X1 U6003 ( .A1(n4881), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4877) );
  OAI22_X1 U6004 ( .A1(n4883), .A2(n6027), .B1(n6573), .B2(n4882), .ZN(n4875)
         );
  AOI21_X1 U6005 ( .B1(n6422), .B2(n6507), .A(n4875), .ZN(n4876) );
  OAI211_X1 U6006 ( .C1(n4887), .C2(n6574), .A(n4877), .B(n4876), .ZN(U3043)
         );
  NAND2_X1 U6007 ( .A1(n4881), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4880) );
  OAI22_X1 U6008 ( .A1(n4883), .A2(n6021), .B1(n6567), .B2(n4882), .ZN(n4878)
         );
  AOI21_X1 U6009 ( .B1(n6422), .B2(n6849), .A(n4878), .ZN(n4879) );
  OAI211_X1 U6010 ( .C1(n4887), .C2(n6854), .A(n4880), .B(n4879), .ZN(U3042)
         );
  NAND2_X1 U6011 ( .A1(n4881), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4886) );
  OAI22_X1 U6012 ( .A1(n4883), .A2(n5997), .B1(n6512), .B2(n4882), .ZN(n4884)
         );
  AOI21_X1 U6013 ( .B1(n6422), .B2(n6480), .A(n4884), .ZN(n4885) );
  OAI211_X1 U6014 ( .C1(n4887), .C2(n6533), .A(n4886), .B(n4885), .ZN(U3036)
         );
  INV_X1 U6015 ( .A(n4888), .ZN(n4890) );
  NOR3_X1 U6016 ( .A1(n4890), .A2(n4889), .A3(n5163), .ZN(n5969) );
  INV_X1 U6017 ( .A(n6516), .ZN(n4891) );
  NAND3_X1 U6018 ( .A1(n5969), .A2(n4891), .A3(n5966), .ZN(n4892) );
  NAND2_X1 U6019 ( .A1(n4892), .A2(n6524), .ZN(n4899) );
  OR2_X1 U6020 ( .A1(n4893), .A2(n5541), .ZN(n4894) );
  OR2_X1 U6021 ( .A1(n4896), .A2(n6033), .ZN(n6410) );
  INV_X1 U6022 ( .A(n4895), .ZN(n4898) );
  NAND2_X1 U6023 ( .A1(n6428), .A2(n4896), .ZN(n4897) );
  OAI211_X1 U6024 ( .C1(n4899), .C2(n4898), .A(n6522), .B(n4897), .ZN(n6424)
         );
  NOR2_X1 U6025 ( .A1(n6853), .A2(n6547), .ZN(n4902) );
  INV_X1 U6026 ( .A(n6422), .ZN(n4910) );
  OAI22_X1 U6027 ( .A1(n4910), .A2(n6552), .B1(n6546), .B2(n6410), .ZN(n4901)
         );
  AOI211_X1 U6028 ( .C1(n6424), .C2(INSTQUEUE_REG_3__3__SCAN_IN), .A(n4902), 
        .B(n4901), .ZN(n4903) );
  OAI21_X1 U6029 ( .B1(n4914), .B2(n6009), .A(n4903), .ZN(U3047) );
  NOR2_X1 U6030 ( .A1(n6853), .A2(n6568), .ZN(n4905) );
  OAI22_X1 U6031 ( .A1(n4910), .A2(n6854), .B1(n6567), .B2(n6410), .ZN(n4904)
         );
  AOI211_X1 U6032 ( .C1(n6424), .C2(INSTQUEUE_REG_3__6__SCAN_IN), .A(n4905), 
        .B(n4904), .ZN(n4906) );
  OAI21_X1 U6033 ( .B1(n4914), .B2(n6021), .A(n4906), .ZN(U3050) );
  NOR2_X1 U6034 ( .A1(n6853), .A2(n6538), .ZN(n4908) );
  OAI22_X1 U6035 ( .A1(n4910), .A2(n6589), .B1(n6534), .B2(n6410), .ZN(n4907)
         );
  AOI211_X1 U6036 ( .C1(n6424), .C2(INSTQUEUE_REG_3__1__SCAN_IN), .A(n4908), 
        .B(n4907), .ZN(n4909) );
  OAI21_X1 U6037 ( .B1(n4914), .B2(n6001), .A(n4909), .ZN(U3045) );
  NOR2_X1 U6038 ( .A1(n6853), .A2(n6513), .ZN(n4912) );
  OAI22_X1 U6039 ( .A1(n4910), .A2(n6533), .B1(n6512), .B2(n6410), .ZN(n4911)
         );
  AOI211_X1 U6040 ( .C1(n6424), .C2(INSTQUEUE_REG_3__0__SCAN_IN), .A(n4912), 
        .B(n4911), .ZN(n4913) );
  OAI21_X1 U6041 ( .B1(n4914), .B2(n5997), .A(n4913), .ZN(U3044) );
  NAND2_X1 U6042 ( .A1(n5964), .A2(n4555), .ZN(n6473) );
  INV_X1 U6043 ( .A(n6473), .ZN(n5165) );
  NAND2_X1 U6044 ( .A1(n6474), .A2(n5165), .ZN(n5118) );
  OAI211_X1 U6045 ( .C1(n4976), .C2(n4952), .A(n5125), .B(n5118), .ZN(n4920)
         );
  INV_X1 U6046 ( .A(n4915), .ZN(n4916) );
  NAND2_X1 U6047 ( .A1(n4916), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6427) );
  AOI21_X1 U6048 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6467), .A(n5017), .ZN(
        n4917) );
  NAND2_X1 U6049 ( .A1(n6464), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6435) );
  NAND2_X1 U6050 ( .A1(n4918), .A2(n5983), .ZN(n5124) );
  OR2_X1 U6051 ( .A1(n5124), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4947)
         );
  NAND2_X1 U6052 ( .A1(n4947), .A2(STATE2_REG_3__SCAN_IN), .ZN(n4919) );
  NAND2_X1 U6053 ( .A1(n4946), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4927) );
  INV_X1 U6054 ( .A(n4921), .ZN(n4922) );
  INV_X1 U6055 ( .A(n5118), .ZN(n4924) );
  INV_X1 U6056 ( .A(n6465), .ZN(n6035) );
  NOR3_X1 U6057 ( .A1(n6035), .A2(n6464), .A3(n6467), .ZN(n4923) );
  AOI21_X1 U6058 ( .B1(n4924), .B2(n6515), .A(n4923), .ZN(n4948) );
  OAI22_X1 U6059 ( .A1(n4948), .A2(n6021), .B1(n6567), .B2(n4947), .ZN(n4925)
         );
  AOI21_X1 U6060 ( .B1(n5122), .B2(n6849), .A(n4925), .ZN(n4926) );
  OAI211_X1 U6061 ( .C1(n4952), .C2(n6854), .A(n4927), .B(n4926), .ZN(U3026)
         );
  NAND2_X1 U6062 ( .A1(n4946), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4930) );
  OAI22_X1 U6063 ( .A1(n4948), .A2(n5997), .B1(n6512), .B2(n4947), .ZN(n4928)
         );
  AOI21_X1 U6064 ( .B1(n5122), .B2(n6480), .A(n4928), .ZN(n4929) );
  OAI211_X1 U6065 ( .C1(n4952), .C2(n6533), .A(n4930), .B(n4929), .ZN(U3020)
         );
  NAND2_X1 U6066 ( .A1(n4946), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4933) );
  OAI22_X1 U6067 ( .A1(n4948), .A2(n6009), .B1(n6546), .B2(n4947), .ZN(n4931)
         );
  AOI21_X1 U6068 ( .B1(n5122), .B2(n6490), .A(n4931), .ZN(n4932) );
  OAI211_X1 U6069 ( .C1(n4952), .C2(n6552), .A(n4933), .B(n4932), .ZN(U3023)
         );
  NAND2_X1 U6070 ( .A1(n4946), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4936) );
  OAI22_X1 U6071 ( .A1(n4948), .A2(n6013), .B1(n6553), .B2(n4947), .ZN(n4934)
         );
  AOI21_X1 U6072 ( .B1(n5122), .B2(n6494), .A(n4934), .ZN(n4935) );
  OAI211_X1 U6073 ( .C1(n4952), .C2(n6554), .A(n4936), .B(n4935), .ZN(U3024)
         );
  NAND2_X1 U6074 ( .A1(n4946), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4939) );
  OAI22_X1 U6075 ( .A1(n4948), .A2(n6017), .B1(n6560), .B2(n4947), .ZN(n4937)
         );
  AOI21_X1 U6076 ( .B1(n5122), .B2(n6498), .A(n4937), .ZN(n4938) );
  OAI211_X1 U6077 ( .C1(n4952), .C2(n6566), .A(n4939), .B(n4938), .ZN(U3025)
         );
  NAND2_X1 U6078 ( .A1(n4946), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4942) );
  OAI22_X1 U6079 ( .A1(n4948), .A2(n6027), .B1(n6573), .B2(n4947), .ZN(n4940)
         );
  AOI21_X1 U6080 ( .B1(n5122), .B2(n6507), .A(n4940), .ZN(n4941) );
  OAI211_X1 U6081 ( .C1(n4952), .C2(n6574), .A(n4942), .B(n4941), .ZN(U3027)
         );
  NAND2_X1 U6082 ( .A1(n4946), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4945) );
  OAI22_X1 U6083 ( .A1(n4948), .A2(n6005), .B1(n6539), .B2(n4947), .ZN(n4943)
         );
  AOI21_X1 U6084 ( .B1(n5122), .B2(n6486), .A(n4943), .ZN(n4944) );
  OAI211_X1 U6085 ( .C1(n4952), .C2(n6545), .A(n4945), .B(n4944), .ZN(U3022)
         );
  NAND2_X1 U6086 ( .A1(n4946), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4951) );
  OAI22_X1 U6087 ( .A1(n4948), .A2(n6001), .B1(n6534), .B2(n4947), .ZN(n4949)
         );
  AOI21_X1 U6088 ( .B1(n5122), .B2(n6586), .A(n4949), .ZN(n4950) );
  OAI211_X1 U6089 ( .C1(n4952), .C2(n6589), .A(n4951), .B(n4950), .ZN(U3021)
         );
  AND2_X1 U6090 ( .A1(n4953), .A2(n4954), .ZN(n4956) );
  OR2_X1 U6091 ( .A1(n4956), .A2(n4955), .ZN(n5217) );
  AOI22_X1 U6092 ( .A1(n6257), .A2(DATAI_8_), .B1(n6253), .B2(
        EAX_REG_8__SCAN_IN), .ZN(n4957) );
  OAI21_X1 U6093 ( .B1(n5217), .B2(n5635), .A(n4957), .ZN(U2883) );
  INV_X1 U6094 ( .A(n5520), .ZN(n4961) );
  AOI21_X1 U6095 ( .B1(n6351), .B2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n4958), 
        .ZN(n4959) );
  OAI21_X1 U6096 ( .B1(n5511), .B2(n6362), .A(n4959), .ZN(n4960) );
  AOI21_X1 U6097 ( .B1(n4961), .B2(n6358), .A(n4960), .ZN(n4962) );
  OAI21_X1 U6098 ( .B1(n6092), .B2(n4963), .A(n4962), .ZN(U2980) );
  INV_X1 U6099 ( .A(n4964), .ZN(n4965) );
  AOI21_X1 U6100 ( .B1(n4965), .B2(n4791), .A(n3113), .ZN(n6198) );
  INV_X1 U6101 ( .A(n6198), .ZN(n4973) );
  AOI22_X1 U6102 ( .A1(n6257), .A2(DATAI_7_), .B1(n6253), .B2(
        EAX_REG_7__SCAN_IN), .ZN(n4966) );
  OAI21_X1 U6103 ( .B1(n4973), .B2(n5635), .A(n4966), .ZN(U2884) );
  INV_X1 U6104 ( .A(EBX_REG_7__SCAN_IN), .ZN(n4972) );
  AND2_X1 U6105 ( .A1(n4793), .A2(n4969), .ZN(n4971) );
  OR2_X1 U6106 ( .A1(n4968), .A2(n4971), .ZN(n6381) );
  OAI222_X1 U6107 ( .A1(n4973), .A2(n5597), .B1(n4972), .B2(n6250), .C1(n5588), 
        .C2(n6381), .ZN(U2852) );
  AND2_X1 U6108 ( .A1(n2976), .A2(n5987), .ZN(n4974) );
  NOR3_X1 U6109 ( .A1(n5001), .A2(n6592), .A3(n6428), .ZN(n4977) );
  OAI22_X1 U6110 ( .A1(n4977), .A2(n4976), .B1(n4975), .B2(n6429), .ZN(n4980)
         );
  AOI211_X1 U6111 ( .C1(n6467), .C2(STATE2_REG_2__SCAN_IN), .A(n6465), .B(
        n5017), .ZN(n6436) );
  OR2_X1 U6112 ( .A1(n6464), .A2(n6527), .ZN(n6477) );
  NOR2_X1 U6113 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4978), .ZN(n6590)
         );
  INV_X1 U6114 ( .A(n6590), .ZN(n4999) );
  NAND2_X1 U6115 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n4999), .ZN(n4979) );
  NAND4_X1 U6116 ( .A1(n4980), .A2(n6436), .A3(n6477), .A4(n4979), .ZN(n6593)
         );
  NAND2_X1 U6117 ( .A1(n6593), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4986)
         );
  AND2_X1 U6118 ( .A1(n6430), .A2(n6515), .ZN(n6463) );
  INV_X1 U6119 ( .A(n6464), .ZN(n4981) );
  NOR3_X1 U6120 ( .A1(n4981), .A2(n6427), .A3(n6467), .ZN(n4982) );
  AOI21_X1 U6121 ( .B1(n4983), .B2(n6463), .A(n4982), .ZN(n6583) );
  OAI22_X1 U6122 ( .A1(n6583), .A2(n6027), .B1(n6573), .B2(n4999), .ZN(n4984)
         );
  AOI21_X1 U6123 ( .B1(n5001), .B2(n6421), .A(n4984), .ZN(n4985) );
  OAI211_X1 U6124 ( .C1(n6582), .C2(n5004), .A(n4986), .B(n4985), .ZN(U3123)
         );
  NAND2_X1 U6125 ( .A1(n6593), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4989)
         );
  OAI22_X1 U6126 ( .A1(n6583), .A2(n6013), .B1(n6553), .B2(n4999), .ZN(n4987)
         );
  AOI21_X1 U6127 ( .B1(n5001), .B2(n6414), .A(n4987), .ZN(n4988) );
  OAI211_X1 U6128 ( .C1(n6559), .C2(n5004), .A(n4989), .B(n4988), .ZN(U3120)
         );
  NAND2_X1 U6129 ( .A1(n6593), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n4992)
         );
  OAI22_X1 U6130 ( .A1(n6583), .A2(n5997), .B1(n6512), .B2(n4999), .ZN(n4990)
         );
  AOI21_X1 U6131 ( .B1(n5001), .B2(n6458), .A(n4990), .ZN(n4991) );
  OAI211_X1 U6132 ( .C1(n5004), .C2(n6513), .A(n4992), .B(n4991), .ZN(U3116)
         );
  NAND2_X1 U6133 ( .A1(n6593), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4995)
         );
  OAI22_X1 U6134 ( .A1(n6583), .A2(n6009), .B1(n6546), .B2(n4999), .ZN(n4993)
         );
  AOI21_X1 U6135 ( .B1(n5001), .B2(n6054), .A(n4993), .ZN(n4994) );
  OAI211_X1 U6136 ( .C1(n6547), .C2(n5004), .A(n4995), .B(n4994), .ZN(U3119)
         );
  NAND2_X1 U6137 ( .A1(n6593), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4998)
         );
  OAI22_X1 U6138 ( .A1(n6583), .A2(n6017), .B1(n6560), .B2(n4999), .ZN(n4996)
         );
  AOI21_X1 U6139 ( .B1(n5001), .B2(n6417), .A(n4996), .ZN(n4997) );
  OAI211_X1 U6140 ( .C1(n6561), .C2(n5004), .A(n4998), .B(n4997), .ZN(U3121)
         );
  NAND2_X1 U6141 ( .A1(n6593), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n5003)
         );
  OAI22_X1 U6142 ( .A1(n6583), .A2(n6005), .B1(n6539), .B2(n4999), .ZN(n5000)
         );
  AOI21_X1 U6143 ( .B1(n5001), .B2(n6411), .A(n5000), .ZN(n5002) );
  OAI211_X1 U6144 ( .C1(n6540), .C2(n5004), .A(n5003), .B(n5002), .ZN(U3118)
         );
  OR2_X1 U6145 ( .A1(n4955), .A2(n5006), .ZN(n5007) );
  NAND2_X1 U6146 ( .A1(n5005), .A2(n5007), .ZN(n6170) );
  INV_X1 U6147 ( .A(n5009), .ZN(n5212) );
  AOI21_X1 U6148 ( .B1(n5010), .B2(n5063), .A(n5212), .ZN(n6372) );
  AOI22_X1 U6149 ( .A1(n6372), .A2(n6247), .B1(EBX_REG_9__SCAN_IN), .B2(n5595), 
        .ZN(n5011) );
  OAI21_X1 U6150 ( .B1(n6170), .B2(n5590), .A(n5011), .ZN(U2850) );
  AOI22_X1 U6151 ( .A1(n6257), .A2(DATAI_9_), .B1(n6253), .B2(
        EAX_REG_9__SCAN_IN), .ZN(n5012) );
  OAI21_X1 U6152 ( .B1(n6170), .B2(n5635), .A(n5012), .ZN(U2882) );
  INV_X1 U6153 ( .A(n5055), .ZN(n5013) );
  OAI21_X1 U6154 ( .B1(n5013), .B2(n5057), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5014) );
  OAI211_X1 U6155 ( .C1(n6474), .C2(n5015), .A(n5014), .B(n6524), .ZN(n5021)
         );
  NOR2_X1 U6156 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5016), .ZN(n5052)
         );
  INV_X1 U6157 ( .A(n5052), .ZN(n5019) );
  NAND2_X1 U6158 ( .A1(n6467), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5084) );
  AOI21_X1 U6159 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5084), .A(n5017), .ZN(
        n5018) );
  INV_X1 U6160 ( .A(n5018), .ZN(n5089) );
  AOI211_X1 U6161 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5019), .A(n5089), .B(
        n6465), .ZN(n5020) );
  INV_X1 U6162 ( .A(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n5027) );
  NAND2_X1 U6163 ( .A1(n6038), .A2(n6463), .ZN(n5023) );
  OR2_X1 U6164 ( .A1(n6427), .A2(n5084), .ZN(n5022) );
  NAND2_X1 U6165 ( .A1(n5023), .A2(n5022), .ZN(n5053) );
  AOI22_X1 U6166 ( .A1(n5053), .A2(n6549), .B1(n6489), .B2(n5052), .ZN(n5024)
         );
  OAI21_X1 U6167 ( .B1(n5055), .B2(n6552), .A(n5024), .ZN(n5025) );
  AOI21_X1 U6168 ( .B1(n6490), .B2(n5057), .A(n5025), .ZN(n5026) );
  OAI21_X1 U6169 ( .B1(n5060), .B2(n5027), .A(n5026), .ZN(U3135) );
  INV_X1 U6170 ( .A(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n5031) );
  AOI22_X1 U6171 ( .A1(n5053), .A2(n6542), .B1(n6485), .B2(n5052), .ZN(n5028)
         );
  OAI21_X1 U6172 ( .B1(n5055), .B2(n6545), .A(n5028), .ZN(n5029) );
  AOI21_X1 U6173 ( .B1(n6486), .B2(n5057), .A(n5029), .ZN(n5030) );
  OAI21_X1 U6174 ( .B1(n5060), .B2(n5031), .A(n5030), .ZN(U3134) );
  AOI22_X1 U6175 ( .A1(n5053), .A2(n6846), .B1(n6845), .B2(n5052), .ZN(n5032)
         );
  OAI21_X1 U6176 ( .B1(n5055), .B2(n6854), .A(n5032), .ZN(n5033) );
  AOI21_X1 U6177 ( .B1(n6849), .B2(n5057), .A(n5033), .ZN(n5034) );
  OAI21_X1 U6178 ( .B1(n5060), .B2(n5035), .A(n5034), .ZN(U3138) );
  INV_X1 U6179 ( .A(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n5039) );
  AOI22_X1 U6180 ( .A1(n5053), .A2(n6578), .B1(n6504), .B2(n5052), .ZN(n5036)
         );
  OAI21_X1 U6181 ( .B1(n5055), .B2(n6574), .A(n5036), .ZN(n5037) );
  AOI21_X1 U6182 ( .B1(n6507), .B2(n5057), .A(n5037), .ZN(n5038) );
  OAI21_X1 U6183 ( .B1(n5060), .B2(n5039), .A(n5038), .ZN(U3139) );
  INV_X1 U6184 ( .A(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n5043) );
  AOI22_X1 U6185 ( .A1(n5053), .A2(n6556), .B1(n6493), .B2(n5052), .ZN(n5040)
         );
  OAI21_X1 U6186 ( .B1(n5055), .B2(n6554), .A(n5040), .ZN(n5041) );
  AOI21_X1 U6187 ( .B1(n6494), .B2(n5057), .A(n5041), .ZN(n5042) );
  OAI21_X1 U6188 ( .B1(n5060), .B2(n5043), .A(n5042), .ZN(U3136) );
  INV_X1 U6189 ( .A(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n5047) );
  AOI22_X1 U6190 ( .A1(n5053), .A2(n6530), .B1(n6470), .B2(n5052), .ZN(n5044)
         );
  OAI21_X1 U6191 ( .B1(n5055), .B2(n6533), .A(n5044), .ZN(n5045) );
  AOI21_X1 U6192 ( .B1(n6480), .B2(n5057), .A(n5045), .ZN(n5046) );
  OAI21_X1 U6193 ( .B1(n5060), .B2(n5047), .A(n5046), .ZN(U3132) );
  INV_X1 U6194 ( .A(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n5051) );
  AOI22_X1 U6195 ( .A1(n5053), .A2(n6585), .B1(n6584), .B2(n5052), .ZN(n5048)
         );
  OAI21_X1 U6196 ( .B1(n5055), .B2(n6589), .A(n5048), .ZN(n5049) );
  AOI21_X1 U6197 ( .B1(n6586), .B2(n5057), .A(n5049), .ZN(n5050) );
  OAI21_X1 U6198 ( .B1(n5060), .B2(n5051), .A(n5050), .ZN(U3133) );
  INV_X1 U6199 ( .A(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n5059) );
  AOI22_X1 U6200 ( .A1(n5053), .A2(n6563), .B1(n6497), .B2(n5052), .ZN(n5054)
         );
  OAI21_X1 U6201 ( .B1(n5055), .B2(n6566), .A(n5054), .ZN(n5056) );
  AOI21_X1 U6202 ( .B1(n6498), .B2(n5057), .A(n5056), .ZN(n5058) );
  OAI21_X1 U6203 ( .B1(n5060), .B2(n5059), .A(n5058), .ZN(U3137) );
  INV_X1 U6204 ( .A(n5217), .ZN(n6184) );
  OR2_X1 U6205 ( .A1(n4968), .A2(n5061), .ZN(n5062) );
  NAND2_X1 U6206 ( .A1(n5063), .A2(n5062), .ZN(n6177) );
  OAI22_X1 U6207 ( .A1(n6177), .A2(n5588), .B1(n6179), .B2(n6250), .ZN(n5064)
         );
  AOI21_X1 U6208 ( .B1(n6184), .B2(n6248), .A(n5064), .ZN(n5065) );
  INV_X1 U6209 ( .A(n5065), .ZN(U2851) );
  XNOR2_X1 U6210 ( .A(n5066), .B(n5067), .ZN(n5221) );
  NOR2_X1 U6211 ( .A1(n5069), .A2(n5068), .ZN(n6378) );
  AOI21_X1 U6212 ( .B1(n6386), .B2(n5075), .A(n5956), .ZN(n5078) );
  NAND2_X1 U6213 ( .A1(n6350), .A2(REIP_REG_8__SCAN_IN), .ZN(n5215) );
  OAI21_X1 U6214 ( .B1(n6177), .B2(n6382), .A(n5215), .ZN(n5077) );
  INV_X1 U6215 ( .A(n5069), .ZN(n5072) );
  OAI21_X1 U6216 ( .B1(n5072), .B2(n5071), .A(n3058), .ZN(n5073) );
  AOI21_X1 U6217 ( .B1(n5892), .B2(n5074), .A(n5073), .ZN(n6387) );
  NOR2_X1 U6218 ( .A1(n6387), .A2(n5075), .ZN(n5076) );
  AOI211_X1 U6219 ( .C1(n6378), .C2(n5078), .A(n5077), .B(n5076), .ZN(n5079)
         );
  OAI21_X1 U6220 ( .B1(n5961), .B2(n5221), .A(n5079), .ZN(U3010) );
  INV_X1 U6221 ( .A(n5163), .ZN(n6517) );
  NOR2_X1 U6222 ( .A1(n6517), .A2(n2976), .ZN(n5171) );
  AND2_X1 U6223 ( .A1(n2976), .A2(n5986), .ZN(n5080) );
  INV_X1 U6224 ( .A(n6575), .ZN(n5081) );
  OAI21_X1 U6225 ( .B1(n5202), .B2(n5081), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5082) );
  NAND2_X1 U6226 ( .A1(n5082), .A2(n6524), .ZN(n5091) );
  INV_X1 U6227 ( .A(n5091), .ZN(n5086) );
  INV_X1 U6228 ( .A(n5084), .ZN(n5085) );
  AND3_X1 U6229 ( .A1(n5087), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6525) );
  NAND2_X1 U6230 ( .A1(n6525), .A2(n6033), .ZN(n5112) );
  OAI22_X1 U6231 ( .A1(n6575), .A2(n6540), .B1(n6539), .B2(n5112), .ZN(n5088)
         );
  AOI21_X1 U6232 ( .B1(n6411), .B2(n5202), .A(n5088), .ZN(n5093) );
  AOI21_X1 U6233 ( .B1(n5112), .B2(STATE2_REG_3__SCAN_IN), .A(n5089), .ZN(
        n5090) );
  NAND2_X1 U6234 ( .A1(n5114), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n5092)
         );
  OAI211_X1 U6235 ( .C1(n5117), .C2(n6005), .A(n5093), .B(n5092), .ZN(U3102)
         );
  OAI22_X1 U6236 ( .A1(n6575), .A2(n6568), .B1(n6567), .B2(n5112), .ZN(n5094)
         );
  AOI21_X1 U6237 ( .B1(n6067), .B2(n5202), .A(n5094), .ZN(n5096) );
  NAND2_X1 U6238 ( .A1(n5114), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n5095)
         );
  OAI211_X1 U6239 ( .C1(n5117), .C2(n6021), .A(n5096), .B(n5095), .ZN(U3106)
         );
  OAI22_X1 U6240 ( .A1(n6575), .A2(n6559), .B1(n6553), .B2(n5112), .ZN(n5097)
         );
  AOI21_X1 U6241 ( .B1(n6414), .B2(n5202), .A(n5097), .ZN(n5099) );
  NAND2_X1 U6242 ( .A1(n5114), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n5098)
         );
  OAI211_X1 U6243 ( .C1(n5117), .C2(n6013), .A(n5099), .B(n5098), .ZN(U3104)
         );
  OAI22_X1 U6244 ( .A1(n6575), .A2(n6547), .B1(n6546), .B2(n5112), .ZN(n5100)
         );
  AOI21_X1 U6245 ( .B1(n6054), .B2(n5202), .A(n5100), .ZN(n5102) );
  NAND2_X1 U6246 ( .A1(n5114), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n5101)
         );
  OAI211_X1 U6247 ( .C1(n5117), .C2(n6009), .A(n5102), .B(n5101), .ZN(U3103)
         );
  OAI22_X1 U6248 ( .A1(n6575), .A2(n6513), .B1(n6512), .B2(n5112), .ZN(n5103)
         );
  AOI21_X1 U6249 ( .B1(n6458), .B2(n5202), .A(n5103), .ZN(n5105) );
  NAND2_X1 U6250 ( .A1(n5114), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n5104)
         );
  OAI211_X1 U6251 ( .C1(n5117), .C2(n5997), .A(n5105), .B(n5104), .ZN(U3100)
         );
  OAI22_X1 U6252 ( .A1(n6575), .A2(n6538), .B1(n6534), .B2(n5112), .ZN(n5106)
         );
  AOI21_X1 U6253 ( .B1(n6045), .B2(n5202), .A(n5106), .ZN(n5108) );
  NAND2_X1 U6254 ( .A1(n5114), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n5107)
         );
  OAI211_X1 U6255 ( .C1(n5117), .C2(n6001), .A(n5108), .B(n5107), .ZN(U3101)
         );
  OAI22_X1 U6256 ( .A1(n6575), .A2(n6582), .B1(n6573), .B2(n5112), .ZN(n5109)
         );
  AOI21_X1 U6257 ( .B1(n6421), .B2(n5202), .A(n5109), .ZN(n5111) );
  NAND2_X1 U6258 ( .A1(n5114), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n5110)
         );
  OAI211_X1 U6259 ( .C1(n5117), .C2(n6027), .A(n5111), .B(n5110), .ZN(U3107)
         );
  OAI22_X1 U6260 ( .A1(n6575), .A2(n6561), .B1(n6560), .B2(n5112), .ZN(n5113)
         );
  AOI21_X1 U6261 ( .B1(n6417), .B2(n5202), .A(n5113), .ZN(n5116) );
  NAND2_X1 U6262 ( .A1(n5114), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n5115)
         );
  OAI211_X1 U6263 ( .C1(n5117), .C2(n6017), .A(n5116), .B(n5115), .ZN(U3105)
         );
  OR2_X1 U6264 ( .A1(n5118), .A2(n5541), .ZN(n5120) );
  NOR2_X1 U6265 ( .A1(n5124), .A2(n6033), .ZN(n5150) );
  INV_X1 U6266 ( .A(n5150), .ZN(n5119) );
  NAND2_X1 U6267 ( .A1(n5120), .A2(n5119), .ZN(n5123) );
  INV_X1 U6268 ( .A(n5124), .ZN(n5121) );
  INV_X1 U6269 ( .A(n5123), .ZN(n5126) );
  AOI22_X1 U6270 ( .A1(n5126), .A2(n5125), .B1(n6428), .B2(n5124), .ZN(n5127)
         );
  NAND2_X1 U6271 ( .A1(n6522), .A2(n5127), .ZN(n5149) );
  AOI22_X1 U6272 ( .A1(n6504), .A2(n5150), .B1(INSTQUEUE_REG_1__7__SCAN_IN), 
        .B2(n5149), .ZN(n5128) );
  OAI21_X1 U6273 ( .B1(n5152), .B2(n6574), .A(n5128), .ZN(n5129) );
  AOI21_X1 U6274 ( .B1(n6507), .B2(n5154), .A(n5129), .ZN(n5130) );
  OAI21_X1 U6275 ( .B1(n5156), .B2(n6027), .A(n5130), .ZN(U3035) );
  AOI22_X1 U6276 ( .A1(n6493), .A2(n5150), .B1(INSTQUEUE_REG_1__4__SCAN_IN), 
        .B2(n5149), .ZN(n5131) );
  OAI21_X1 U6277 ( .B1(n5152), .B2(n6554), .A(n5131), .ZN(n5132) );
  AOI21_X1 U6278 ( .B1(n6494), .B2(n5154), .A(n5132), .ZN(n5133) );
  OAI21_X1 U6279 ( .B1(n5156), .B2(n6013), .A(n5133), .ZN(U3032) );
  AOI22_X1 U6280 ( .A1(n6497), .A2(n5150), .B1(INSTQUEUE_REG_1__5__SCAN_IN), 
        .B2(n5149), .ZN(n5134) );
  OAI21_X1 U6281 ( .B1(n5152), .B2(n6566), .A(n5134), .ZN(n5135) );
  AOI21_X1 U6282 ( .B1(n6498), .B2(n5154), .A(n5135), .ZN(n5136) );
  OAI21_X1 U6283 ( .B1(n5156), .B2(n6017), .A(n5136), .ZN(U3033) );
  AOI22_X1 U6284 ( .A1(n6485), .A2(n5150), .B1(INSTQUEUE_REG_1__2__SCAN_IN), 
        .B2(n5149), .ZN(n5137) );
  OAI21_X1 U6285 ( .B1(n5152), .B2(n6545), .A(n5137), .ZN(n5138) );
  AOI21_X1 U6286 ( .B1(n6486), .B2(n5154), .A(n5138), .ZN(n5139) );
  OAI21_X1 U6287 ( .B1(n5156), .B2(n6005), .A(n5139), .ZN(U3030) );
  AOI22_X1 U6288 ( .A1(n6489), .A2(n5150), .B1(INSTQUEUE_REG_1__3__SCAN_IN), 
        .B2(n5149), .ZN(n5140) );
  OAI21_X1 U6289 ( .B1(n5152), .B2(n6552), .A(n5140), .ZN(n5141) );
  AOI21_X1 U6290 ( .B1(n6490), .B2(n5154), .A(n5141), .ZN(n5142) );
  OAI21_X1 U6291 ( .B1(n5156), .B2(n6009), .A(n5142), .ZN(U3031) );
  AOI22_X1 U6292 ( .A1(n6470), .A2(n5150), .B1(INSTQUEUE_REG_1__0__SCAN_IN), 
        .B2(n5149), .ZN(n5143) );
  OAI21_X1 U6293 ( .B1(n5152), .B2(n6533), .A(n5143), .ZN(n5144) );
  AOI21_X1 U6294 ( .B1(n6480), .B2(n5154), .A(n5144), .ZN(n5145) );
  OAI21_X1 U6295 ( .B1(n5156), .B2(n5997), .A(n5145), .ZN(U3028) );
  AOI22_X1 U6296 ( .A1(n6584), .A2(n5150), .B1(INSTQUEUE_REG_1__1__SCAN_IN), 
        .B2(n5149), .ZN(n5146) );
  OAI21_X1 U6297 ( .B1(n5152), .B2(n6589), .A(n5146), .ZN(n5147) );
  AOI21_X1 U6298 ( .B1(n6586), .B2(n5154), .A(n5147), .ZN(n5148) );
  OAI21_X1 U6299 ( .B1(n5156), .B2(n6001), .A(n5148), .ZN(U3029) );
  AOI22_X1 U6300 ( .A1(n6845), .A2(n5150), .B1(INSTQUEUE_REG_1__6__SCAN_IN), 
        .B2(n5149), .ZN(n5151) );
  OAI21_X1 U6301 ( .B1(n5152), .B2(n6854), .A(n5151), .ZN(n5153) );
  AOI21_X1 U6302 ( .B1(n6849), .B2(n5154), .A(n5153), .ZN(n5155) );
  OAI21_X1 U6303 ( .B1(n5156), .B2(n6021), .A(n5155), .ZN(U3034) );
  XOR2_X1 U6304 ( .A(n5158), .B(n5157), .Z(n6384) );
  INV_X1 U6305 ( .A(n6384), .ZN(n5162) );
  NAND2_X1 U6306 ( .A1(n6350), .A2(REIP_REG_7__SCAN_IN), .ZN(n6379) );
  NAND2_X1 U6307 ( .A1(n6351), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n5159)
         );
  OAI211_X1 U6308 ( .C1(n6362), .C2(n6200), .A(n6379), .B(n5159), .ZN(n5160)
         );
  AOI21_X1 U6309 ( .B1(n6198), .B2(n6358), .A(n5160), .ZN(n5161) );
  OAI21_X1 U6310 ( .B1(n5162), .B2(n6092), .A(n5161), .ZN(U2979) );
  NAND3_X1 U6311 ( .A1(n5163), .A2(n5979), .A3(STATEBS16_REG_SCAN_IN), .ZN(
        n5164) );
  NAND2_X1 U6312 ( .A1(n5164), .A2(n6524), .ZN(n5175) );
  INV_X1 U6313 ( .A(n5175), .ZN(n5170) );
  NAND2_X1 U6314 ( .A1(n5166), .A2(n5165), .ZN(n5168) );
  NOR2_X1 U6315 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n5167) );
  NAND2_X1 U6316 ( .A1(n5167), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6469) );
  OR2_X1 U6317 ( .A1(n6469), .A2(n6033), .ZN(n5172) );
  NAND2_X1 U6318 ( .A1(n5168), .A2(n5172), .ZN(n5174) );
  INV_X1 U6319 ( .A(n6469), .ZN(n5169) );
  INV_X1 U6320 ( .A(n5172), .ZN(n5198) );
  NAND2_X1 U6321 ( .A1(n6428), .A2(n6469), .ZN(n5173) );
  OAI211_X1 U6322 ( .C1(n5175), .C2(n5174), .A(n6522), .B(n5173), .ZN(n5197)
         );
  AOI22_X1 U6323 ( .A1(n6845), .A2(n5198), .B1(INSTQUEUE_REG_9__6__SCAN_IN), 
        .B2(n5197), .ZN(n5176) );
  OAI21_X1 U6324 ( .B1(n5200), .B2(n6854), .A(n5176), .ZN(n5177) );
  AOI21_X1 U6325 ( .B1(n6849), .B2(n5202), .A(n5177), .ZN(n5178) );
  OAI21_X1 U6326 ( .B1(n5204), .B2(n6021), .A(n5178), .ZN(U3098) );
  AOI22_X1 U6327 ( .A1(n6584), .A2(n5198), .B1(INSTQUEUE_REG_9__1__SCAN_IN), 
        .B2(n5197), .ZN(n5179) );
  OAI21_X1 U6328 ( .B1(n5200), .B2(n6589), .A(n5179), .ZN(n5180) );
  AOI21_X1 U6329 ( .B1(n6586), .B2(n5202), .A(n5180), .ZN(n5181) );
  OAI21_X1 U6330 ( .B1(n5204), .B2(n6001), .A(n5181), .ZN(U3093) );
  AOI22_X1 U6331 ( .A1(n6497), .A2(n5198), .B1(INSTQUEUE_REG_9__5__SCAN_IN), 
        .B2(n5197), .ZN(n5182) );
  OAI21_X1 U6332 ( .B1(n5200), .B2(n6566), .A(n5182), .ZN(n5183) );
  AOI21_X1 U6333 ( .B1(n6498), .B2(n5202), .A(n5183), .ZN(n5184) );
  OAI21_X1 U6334 ( .B1(n5204), .B2(n6017), .A(n5184), .ZN(U3097) );
  AOI22_X1 U6335 ( .A1(n6485), .A2(n5198), .B1(INSTQUEUE_REG_9__2__SCAN_IN), 
        .B2(n5197), .ZN(n5185) );
  OAI21_X1 U6336 ( .B1(n5200), .B2(n6545), .A(n5185), .ZN(n5186) );
  AOI21_X1 U6337 ( .B1(n6486), .B2(n5202), .A(n5186), .ZN(n5187) );
  OAI21_X1 U6338 ( .B1(n5204), .B2(n6005), .A(n5187), .ZN(U3094) );
  AOI22_X1 U6339 ( .A1(n6493), .A2(n5198), .B1(INSTQUEUE_REG_9__4__SCAN_IN), 
        .B2(n5197), .ZN(n5188) );
  OAI21_X1 U6340 ( .B1(n5200), .B2(n6554), .A(n5188), .ZN(n5189) );
  AOI21_X1 U6341 ( .B1(n6494), .B2(n5202), .A(n5189), .ZN(n5190) );
  OAI21_X1 U6342 ( .B1(n5204), .B2(n6013), .A(n5190), .ZN(U3096) );
  AOI22_X1 U6343 ( .A1(n6504), .A2(n5198), .B1(INSTQUEUE_REG_9__7__SCAN_IN), 
        .B2(n5197), .ZN(n5191) );
  OAI21_X1 U6344 ( .B1(n5200), .B2(n6574), .A(n5191), .ZN(n5192) );
  AOI21_X1 U6345 ( .B1(n6507), .B2(n5202), .A(n5192), .ZN(n5193) );
  OAI21_X1 U6346 ( .B1(n5204), .B2(n6027), .A(n5193), .ZN(U3099) );
  AOI22_X1 U6347 ( .A1(n6489), .A2(n5198), .B1(INSTQUEUE_REG_9__3__SCAN_IN), 
        .B2(n5197), .ZN(n5194) );
  OAI21_X1 U6348 ( .B1(n5200), .B2(n6552), .A(n5194), .ZN(n5195) );
  AOI21_X1 U6349 ( .B1(n6490), .B2(n5202), .A(n5195), .ZN(n5196) );
  OAI21_X1 U6350 ( .B1(n5204), .B2(n6009), .A(n5196), .ZN(U3095) );
  AOI22_X1 U6351 ( .A1(n6470), .A2(n5198), .B1(INSTQUEUE_REG_9__0__SCAN_IN), 
        .B2(n5197), .ZN(n5199) );
  OAI21_X1 U6352 ( .B1(n5200), .B2(n6533), .A(n5199), .ZN(n5201) );
  AOI21_X1 U6353 ( .B1(n6480), .B2(n5202), .A(n5201), .ZN(n5203) );
  OAI21_X1 U6354 ( .B1(n5204), .B2(n5997), .A(n5203), .ZN(U3092) );
  NAND2_X1 U6355 ( .A1(n5005), .A2(n5206), .ZN(n5207) );
  AOI22_X1 U6356 ( .A1(n6257), .A2(DATAI_10_), .B1(n6253), .B2(
        EAX_REG_10__SCAN_IN), .ZN(n5208) );
  OAI21_X1 U6357 ( .B1(n5214), .B2(n5635), .A(n5208), .ZN(U2881) );
  INV_X1 U6358 ( .A(EBX_REG_10__SCAN_IN), .ZN(n5213) );
  INV_X1 U6359 ( .A(n5209), .ZN(n5211) );
  OAI21_X1 U6360 ( .B1(n5212), .B2(n5211), .A(n5210), .ZN(n6161) );
  OAI222_X1 U6361 ( .A1(n5214), .A2(n5597), .B1(n5213), .B2(n6250), .C1(n5588), 
        .C2(n6161), .ZN(U2849) );
  INV_X1 U6362 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n5216) );
  OAI21_X1 U6363 ( .B1(n5775), .B2(n5216), .A(n5215), .ZN(n5219) );
  NOR2_X1 U6364 ( .A1(n5217), .A2(n5782), .ZN(n5218) );
  AOI211_X1 U6365 ( .C1(n5778), .C2(n6182), .A(n5219), .B(n5218), .ZN(n5220)
         );
  OAI21_X1 U6366 ( .B1(n6092), .B2(n5221), .A(n5220), .ZN(U2978) );
  XNOR2_X1 U6367 ( .A(n5762), .B(n6764), .ZN(n5223) );
  XNOR2_X1 U6368 ( .A(n5222), .B(n5223), .ZN(n6374) );
  NAND2_X1 U6369 ( .A1(n6374), .A2(n4193), .ZN(n5227) );
  INV_X1 U6370 ( .A(REIP_REG_9__SCAN_IN), .ZN(n5224) );
  NOR2_X1 U6371 ( .A1(n6398), .A2(n5224), .ZN(n6371) );
  NOR2_X1 U6372 ( .A1(n6362), .A2(n6171), .ZN(n5225) );
  AOI211_X1 U6373 ( .C1(n6351), .C2(PHYADDRPOINTER_REG_9__SCAN_IN), .A(n6371), 
        .B(n5225), .ZN(n5226) );
  OAI211_X1 U6374 ( .C1(n5782), .C2(n6170), .A(n5227), .B(n5226), .ZN(U2977)
         );
  INV_X1 U6375 ( .A(n5228), .ZN(n5593) );
  INV_X1 U6376 ( .A(n5934), .ZN(n5229) );
  AOI21_X1 U6377 ( .B1(n5230), .B2(n5210), .A(n5229), .ZN(n6364) );
  AOI22_X1 U6378 ( .A1(n6364), .A2(n6247), .B1(EBX_REG_11__SCAN_IN), .B2(n5595), .ZN(n5231) );
  OAI21_X1 U6379 ( .B1(n5781), .B2(n5597), .A(n5231), .ZN(U2848) );
  AOI22_X1 U6380 ( .A1(n6257), .A2(DATAI_11_), .B1(n6253), .B2(
        EAX_REG_11__SCAN_IN), .ZN(n5232) );
  OAI21_X1 U6381 ( .B1(n5781), .B2(n5635), .A(n5232), .ZN(U2880) );
  AND2_X1 U6382 ( .A1(STATE2_REG_0__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n5236) );
  NAND2_X1 U6383 ( .A1(n6683), .A2(n5236), .ZN(n6599) );
  NAND2_X1 U6384 ( .A1(n5533), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5269) );
  INV_X1 U6385 ( .A(n5241), .ZN(n5239) );
  NAND2_X1 U6386 ( .A1(n5242), .A2(n5362), .ZN(n5238) );
  NAND3_X1 U6387 ( .A1(n5240), .A2(n5239), .A3(n5238), .ZN(n5244) );
  OAI211_X1 U6388 ( .C1(n5362), .C2(n2969), .A(n5242), .B(n5241), .ZN(n5243)
         );
  NAND2_X1 U6389 ( .A1(n5244), .A2(n5243), .ZN(n5318) );
  NOR2_X1 U6390 ( .A1(n4263), .A2(n5274), .ZN(n5245) );
  AND2_X1 U6391 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n5267) );
  AND2_X1 U6392 ( .A1(n5246), .A2(n5274), .ZN(n5247) );
  INV_X1 U6393 ( .A(REIP_REG_8__SCAN_IN), .ZN(n6623) );
  NAND2_X1 U6394 ( .A1(REIP_REG_7__SCAN_IN), .A2(REIP_REG_6__SCAN_IN), .ZN(
        n6192) );
  NAND4_X1 U6395 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_3__SCAN_IN), .A3(
        REIP_REG_2__SCAN_IN), .A4(n5533), .ZN(n6218) );
  NAND2_X1 U6396 ( .A1(REIP_REG_5__SCAN_IN), .A2(n5260), .ZN(n5515) );
  NAND3_X1 U6397 ( .A1(REIP_REG_14__SCAN_IN), .A2(REIP_REG_13__SCAN_IN), .A3(
        REIP_REG_12__SCAN_IN), .ZN(n5250) );
  NAND2_X1 U6398 ( .A1(REIP_REG_15__SCAN_IN), .A2(REIP_REG_16__SCAN_IN), .ZN(
        n6110) );
  INV_X1 U6399 ( .A(n6110), .ZN(n5251) );
  AND2_X1 U6400 ( .A1(REIP_REG_17__SCAN_IN), .A2(n5251), .ZN(n5263) );
  INV_X1 U6401 ( .A(n5263), .ZN(n5476) );
  NAND2_X1 U6402 ( .A1(n6217), .A2(n5476), .ZN(n5252) );
  NAND2_X1 U6403 ( .A1(n3021), .A2(REIP_REG_18__SCAN_IN), .ZN(n5253) );
  AND2_X1 U6404 ( .A1(n6217), .A2(n5253), .ZN(n5254) );
  INV_X1 U6405 ( .A(REIP_REG_23__SCAN_IN), .ZN(n6644) );
  INV_X1 U6406 ( .A(REIP_REG_22__SCAN_IN), .ZN(n6645) );
  INV_X1 U6407 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6643) );
  OR3_X1 U6408 ( .A1(n6644), .A2(n6645), .A3(n6643), .ZN(n5255) );
  AND2_X1 U6409 ( .A1(n6217), .A2(n5255), .ZN(n5256) );
  AND2_X1 U6410 ( .A1(REIP_REG_26__SCAN_IN), .A2(REIP_REG_25__SCAN_IN), .ZN(
        n5266) );
  INV_X1 U6411 ( .A(n5266), .ZN(n5257) );
  OAI21_X1 U6412 ( .B1(n5257), .B2(n6647), .A(n6217), .ZN(n5258) );
  NAND2_X1 U6413 ( .A1(n5259), .A2(REIP_REG_29__SCAN_IN), .ZN(n5356) );
  NAND2_X1 U6414 ( .A1(n5389), .A2(n5523), .ZN(n5289) );
  NAND3_X1 U6415 ( .A1(n5356), .A2(REIP_REG_30__SCAN_IN), .A3(n5289), .ZN(
        n5286) );
  NAND3_X1 U6416 ( .A1(REIP_REG_11__SCAN_IN), .A2(REIP_REG_10__SCAN_IN), .A3(
        REIP_REG_9__SCAN_IN), .ZN(n5261) );
  AND3_X1 U6417 ( .A1(REIP_REG_12__SCAN_IN), .A2(REIP_REG_14__SCAN_IN), .A3(
        REIP_REG_13__SCAN_IN), .ZN(n5262) );
  NAND2_X1 U6418 ( .A1(n5263), .A2(REIP_REG_18__SCAN_IN), .ZN(n5264) );
  NAND2_X1 U6419 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .ZN(
        n5265) );
  INV_X1 U6420 ( .A(REIP_REG_30__SCAN_IN), .ZN(n6663) );
  NAND2_X1 U6421 ( .A1(n6663), .A2(REIP_REG_29__SCAN_IN), .ZN(n5268) );
  INV_X1 U6422 ( .A(n5269), .ZN(n5270) );
  NAND2_X1 U6423 ( .A1(n6183), .A2(n5326), .ZN(n5282) );
  AND2_X1 U6424 ( .A1(n5273), .A2(n5272), .ZN(n5290) );
  INV_X1 U6425 ( .A(n5290), .ZN(n5279) );
  INV_X1 U6426 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5276) );
  INV_X1 U6427 ( .A(n5274), .ZN(n5275) );
  NAND3_X1 U6428 ( .A1(n5277), .A2(n5276), .A3(n5275), .ZN(n5278) );
  NAND2_X1 U6429 ( .A1(n5279), .A2(n5278), .ZN(n5280) );
  AND2_X2 U6430 ( .A1(n5526), .A2(n5280), .ZN(n6242) );
  AOI22_X1 U6431 ( .A1(n6242), .A2(EBX_REG_30__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n6225), .ZN(n5281) );
  NAND2_X1 U6432 ( .A1(n5282), .A2(n5281), .ZN(n5283) );
  OAI22_X1 U6433 ( .A1(n5294), .A2(n5588), .B1(n6250), .B2(n5276), .ZN(U2828)
         );
  INV_X1 U6434 ( .A(n5322), .ZN(n5344) );
  INV_X1 U6435 ( .A(EBX_REG_30__SCAN_IN), .ZN(n5287) );
  OAI222_X1 U6436 ( .A1(n5588), .A2(n5318), .B1(n5597), .B2(n5344), .C1(n5287), 
        .C2(n6250), .ZN(U2829) );
  NAND3_X1 U6437 ( .A1(n6813), .A2(REIP_REG_30__SCAN_IN), .A3(
        REIP_REG_29__SCAN_IN), .ZN(n5288) );
  NOR2_X1 U6438 ( .A1(n5355), .A2(n5288), .ZN(n5295) );
  OAI211_X1 U6439 ( .C1(n5356), .C2(n6663), .A(REIP_REG_31__SCAN_IN), .B(n5289), .ZN(n5293) );
  AOI22_X1 U6440 ( .A1(n5291), .A2(n5290), .B1(PHYADDRPOINTER_REG_31__SCAN_IN), 
        .B2(n6225), .ZN(n5292) );
  INV_X1 U6441 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n6786) );
  AOI21_X1 U6442 ( .B1(n5297), .B2(n4386), .A(n2977), .ZN(n5407) );
  NOR2_X1 U6443 ( .A1(n6398), .A2(n6647), .ZN(n5308) );
  AOI21_X1 U6444 ( .B1(n6351), .B2(PHYADDRPOINTER_REG_24__SCAN_IN), .A(n5308), 
        .ZN(n5298) );
  OAI21_X1 U6445 ( .B1(n5410), .B2(n6362), .A(n5298), .ZN(n5299) );
  AOI21_X1 U6446 ( .B1(n5407), .B2(n6358), .A(n5299), .ZN(n5300) );
  OAI21_X1 U6447 ( .B1(n5310), .B2(n6092), .A(n5300), .ZN(U2962) );
  AND2_X1 U6448 ( .A1(n5302), .A2(n5301), .ZN(n5303) );
  NOR2_X1 U6449 ( .A1(n5396), .A2(n5303), .ZN(n5553) );
  NAND3_X1 U6450 ( .A1(n5854), .A2(n5304), .A3(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5306) );
  AOI21_X1 U6451 ( .B1(n3158), .B2(n5306), .A(n5305), .ZN(n5307) );
  AOI211_X1 U6452 ( .C1(n5553), .C2(n6395), .A(n5308), .B(n5307), .ZN(n5309)
         );
  OAI21_X1 U6453 ( .B1(n5310), .B2(n5961), .A(n5309), .ZN(U2994) );
  INV_X1 U6454 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5314) );
  INV_X1 U6455 ( .A(n5312), .ZN(n5313) );
  INV_X1 U6456 ( .A(n5315), .ZN(n5317) );
  NOR2_X1 U6457 ( .A1(n6398), .A2(n6663), .ZN(n5325) );
  NOR3_X1 U6458 ( .A1(n5794), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(n5641), 
        .ZN(n5316) );
  AOI211_X1 U6459 ( .C1(n5317), .C2(INSTADDRPOINTER_REG_30__SCAN_IN), .A(n5325), .B(n5316), .ZN(n5321) );
  INV_X1 U6460 ( .A(n5318), .ZN(n5319) );
  NAND2_X1 U6461 ( .A1(n5319), .A2(n6395), .ZN(n5320) );
  OAI211_X1 U6462 ( .C1(n5329), .C2(n5961), .A(n5321), .B(n5320), .ZN(U2988)
         );
  NAND2_X1 U6463 ( .A1(n5322), .A2(n6358), .ZN(n5328) );
  NOR2_X1 U6464 ( .A1(n5775), .A2(n5323), .ZN(n5324) );
  AOI211_X1 U6465 ( .C1(n5326), .C2(n5778), .A(n5325), .B(n5324), .ZN(n5327)
         );
  OAI211_X1 U6466 ( .C1(n5329), .C2(n6092), .A(n5328), .B(n5327), .ZN(U2956)
         );
  NOR2_X1 U6467 ( .A1(n5331), .A2(n5330), .ZN(n5333) );
  NOR3_X1 U6468 ( .A1(n6605), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n5336), 
        .ZN(n5332) );
  AOI211_X1 U6469 ( .C1(n5335), .C2(n5334), .A(n5333), .B(n5332), .ZN(n5340)
         );
  AOI21_X1 U6470 ( .B1(n5337), .B2(n5336), .A(n5977), .ZN(n5339) );
  OAI22_X1 U6471 ( .A1(n5340), .A2(n5977), .B1(n5339), .B2(n5338), .ZN(U3459)
         );
  AOI22_X1 U6472 ( .A1(n6251), .A2(DATAI_30_), .B1(EAX_REG_30__SCAN_IN), .B2(
        n6253), .ZN(n5343) );
  AND2_X1 U6473 ( .A1(n3348), .A2(n3313), .ZN(n5341) );
  NAND2_X1 U6474 ( .A1(n6254), .A2(DATAI_14_), .ZN(n5342) );
  OAI211_X1 U6475 ( .C1(n5344), .C2(n5635), .A(n5343), .B(n5342), .ZN(U2861)
         );
  OR2_X1 U6476 ( .A1(n5468), .A2(READREQUEST_REG_SCAN_IN), .ZN(n5347) );
  NAND2_X1 U6477 ( .A1(n5345), .A2(n4263), .ZN(n5346) );
  MUX2_X1 U6478 ( .A(n5347), .B(n5346), .S(n6679), .Z(U3474) );
  INV_X1 U6479 ( .A(n5362), .ZN(n5352) );
  XNOR2_X1 U6480 ( .A(n5352), .B(n5351), .ZN(n5792) );
  AOI22_X1 U6481 ( .A1(n6242), .A2(EBX_REG_29__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n6225), .ZN(n5353) );
  OAI21_X1 U6482 ( .B1(n6236), .B2(n5637), .A(n5353), .ZN(n5354) );
  AOI21_X1 U6483 ( .B1(n5792), .B2(n6202), .A(n5354), .ZN(n5359) );
  INV_X1 U6484 ( .A(n5355), .ZN(n5357) );
  OAI21_X1 U6485 ( .B1(n5357), .B2(REIP_REG_29__SCAN_IN), .A(n5356), .ZN(n5358) );
  OAI211_X1 U6486 ( .C1(n5645), .C2(n6124), .A(n5359), .B(n5358), .ZN(U2798)
         );
  AOI21_X1 U6487 ( .B1(n5361), .B2(n5360), .A(n5348), .ZN(n5656) );
  INV_X1 U6488 ( .A(n5656), .ZN(n5602) );
  AOI21_X1 U6489 ( .B1(n5363), .B2(n5374), .A(n5362), .ZN(n5807) );
  NAND2_X1 U6490 ( .A1(n5807), .A2(n6202), .ZN(n5365) );
  AOI22_X1 U6491 ( .A1(n6242), .A2(EBX_REG_28__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n6225), .ZN(n5364) );
  OAI211_X1 U6492 ( .C1(n6236), .C2(n5654), .A(n5365), .B(n5364), .ZN(n5366)
         );
  AOI21_X1 U6493 ( .B1(REIP_REG_28__SCAN_IN), .B2(n5367), .A(n5366), .ZN(n5369) );
  INV_X1 U6494 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6654) );
  NAND3_X1 U6495 ( .A1(n5380), .A2(REIP_REG_27__SCAN_IN), .A3(n6654), .ZN(
        n5368) );
  OAI211_X1 U6496 ( .C1(n5602), .C2(n6124), .A(n5369), .B(n5368), .ZN(U2799)
         );
  OAI21_X1 U6497 ( .B1(n5370), .B2(n5371), .A(n5360), .ZN(n5666) );
  INV_X1 U6498 ( .A(n5389), .ZN(n5379) );
  NAND2_X1 U6499 ( .A1(n5387), .A2(n5372), .ZN(n5373) );
  NAND2_X1 U6500 ( .A1(n5374), .A2(n5373), .ZN(n5819) );
  AOI22_X1 U6501 ( .A1(n6242), .A2(EBX_REG_27__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n6225), .ZN(n5377) );
  INV_X1 U6502 ( .A(n5658), .ZN(n5375) );
  NAND2_X1 U6503 ( .A1(n6183), .A2(n5375), .ZN(n5376) );
  OAI211_X1 U6504 ( .C1(n5819), .C2(n6234), .A(n5377), .B(n5376), .ZN(n5378)
         );
  AOI21_X1 U6505 ( .B1(n5379), .B2(REIP_REG_27__SCAN_IN), .A(n5378), .ZN(n5382) );
  INV_X1 U6506 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6652) );
  NAND2_X1 U6507 ( .A1(n5380), .A2(n6652), .ZN(n5381) );
  OAI211_X1 U6508 ( .C1(n5666), .C2(n6124), .A(n5382), .B(n5381), .ZN(U2800)
         );
  AOI21_X1 U6509 ( .B1(n5384), .B2(n5383), .A(n5370), .ZN(n5676) );
  INV_X1 U6510 ( .A(n5676), .ZN(n5607) );
  OR2_X1 U6511 ( .A1(n5397), .A2(n5385), .ZN(n5386) );
  NAND2_X1 U6512 ( .A1(n5387), .A2(n5386), .ZN(n5824) );
  INV_X1 U6513 ( .A(n5824), .ZN(n5393) );
  AOI22_X1 U6514 ( .A1(n6242), .A2(EBX_REG_26__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n6225), .ZN(n5388) );
  OAI21_X1 U6515 ( .B1(n6236), .B2(n5674), .A(n5388), .ZN(n5392) );
  AOI21_X1 U6516 ( .B1(n5403), .B2(REIP_REG_25__SCAN_IN), .A(
        REIP_REG_26__SCAN_IN), .ZN(n5390) );
  NOR2_X1 U6517 ( .A1(n5390), .A2(n5389), .ZN(n5391) );
  AOI211_X1 U6518 ( .C1(n6202), .C2(n5393), .A(n5392), .B(n5391), .ZN(n5394)
         );
  OAI21_X1 U6519 ( .B1(n5607), .B2(n6124), .A(n5394), .ZN(U2801) );
  OAI21_X1 U6520 ( .B1(n2977), .B2(n5395), .A(n5383), .ZN(n5680) );
  INV_X1 U6521 ( .A(REIP_REG_25__SCAN_IN), .ZN(n6650) );
  INV_X1 U6522 ( .A(n5396), .ZN(n5398) );
  AOI21_X1 U6523 ( .B1(n5399), .B2(n5398), .A(n5397), .ZN(n5832) );
  NAND2_X1 U6524 ( .A1(n5832), .A2(n6202), .ZN(n5401) );
  AOI22_X1 U6525 ( .A1(n6242), .A2(EBX_REG_25__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n6225), .ZN(n5400) );
  OAI211_X1 U6526 ( .C1(n6236), .C2(n5682), .A(n5401), .B(n5400), .ZN(n5402)
         );
  AOI21_X1 U6527 ( .B1(n5403), .B2(n6650), .A(n5402), .ZN(n5406) );
  NOR2_X1 U6528 ( .A1(n5404), .A2(REIP_REG_24__SCAN_IN), .ZN(n5411) );
  OAI21_X1 U6529 ( .B1(n5411), .B2(n2985), .A(REIP_REG_25__SCAN_IN), .ZN(n5405) );
  OAI211_X1 U6530 ( .C1(n5680), .C2(n6124), .A(n5406), .B(n5405), .ZN(U2802)
         );
  INV_X1 U6531 ( .A(n5407), .ZN(n5612) );
  NAND2_X1 U6532 ( .A1(n5553), .A2(n6202), .ZN(n5409) );
  AOI22_X1 U6533 ( .A1(n6242), .A2(EBX_REG_24__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n6225), .ZN(n5408) );
  OAI211_X1 U6534 ( .C1(n6236), .C2(n5410), .A(n5409), .B(n5408), .ZN(n5412)
         );
  AOI211_X1 U6535 ( .C1(REIP_REG_24__SCAN_IN), .C2(n2985), .A(n5412), .B(n5411), .ZN(n5413) );
  OAI21_X1 U6536 ( .B1(n5612), .B2(n6124), .A(n5413), .ZN(U2803) );
  OAI21_X1 U6537 ( .B1(n5427), .B2(n6645), .A(n6644), .ZN(n5418) );
  NOR2_X1 U6538 ( .A1(n6236), .A2(n5414), .ZN(n5417) );
  AOI22_X1 U6539 ( .A1(n6242), .A2(EBX_REG_23__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n6225), .ZN(n5415) );
  OAI21_X1 U6540 ( .B1(n5555), .B2(n6234), .A(n5415), .ZN(n5416) );
  AOI211_X1 U6541 ( .C1(n5418), .C2(n2985), .A(n5417), .B(n5416), .ZN(n5419)
         );
  OAI21_X1 U6542 ( .B1(n5615), .B2(n6124), .A(n5419), .ZN(U2804) );
  AOI21_X1 U6543 ( .B1(n5421), .B2(n5420), .A(n2990), .ZN(n5691) );
  INV_X1 U6544 ( .A(n5691), .ZN(n5618) );
  INV_X1 U6545 ( .A(n5689), .ZN(n5430) );
  OR2_X1 U6546 ( .A1(n5423), .A2(n5422), .ZN(n5424) );
  AND2_X1 U6547 ( .A1(n4392), .A2(n5424), .ZN(n5842) );
  NAND2_X1 U6548 ( .A1(n5842), .A2(n6202), .ZN(n5426) );
  AOI22_X1 U6549 ( .A1(n6242), .A2(EBX_REG_22__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n6225), .ZN(n5425) );
  NAND2_X1 U6550 ( .A1(n5426), .A2(n5425), .ZN(n5429) );
  NOR2_X1 U6551 ( .A1(n5427), .A2(REIP_REG_22__SCAN_IN), .ZN(n5428) );
  AOI211_X1 U6552 ( .C1(n6183), .C2(n5430), .A(n5429), .B(n5428), .ZN(n5432)
         );
  NOR2_X1 U6553 ( .A1(n3027), .A2(REIP_REG_21__SCAN_IN), .ZN(n5441) );
  OAI21_X1 U6554 ( .B1(n5441), .B2(n5455), .A(REIP_REG_22__SCAN_IN), .ZN(n5431) );
  OAI211_X1 U6555 ( .C1(n5618), .C2(n6124), .A(n5432), .B(n5431), .ZN(U2805)
         );
  INV_X1 U6556 ( .A(n5433), .ZN(n5435) );
  XNOR2_X1 U6557 ( .A(n5437), .B(n5436), .ZN(n5853) );
  INV_X1 U6558 ( .A(n5696), .ZN(n5438) );
  NAND2_X1 U6559 ( .A1(n6183), .A2(n5438), .ZN(n5440) );
  AOI22_X1 U6560 ( .A1(n6242), .A2(EBX_REG_21__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n6225), .ZN(n5439) );
  OAI211_X1 U6561 ( .C1(n5853), .C2(n6234), .A(n5440), .B(n5439), .ZN(n5442)
         );
  AOI211_X1 U6562 ( .C1(REIP_REG_21__SCAN_IN), .C2(n5455), .A(n5442), .B(n5441), .ZN(n5443) );
  OAI21_X1 U6563 ( .B1(n5700), .B2(n6124), .A(n5443), .ZN(U2806) );
  AND2_X1 U6564 ( .A1(n2974), .A2(n5445), .ZN(n5460) );
  OR2_X1 U6565 ( .A1(n5460), .A2(n5446), .ZN(n5447) );
  NAND2_X1 U6566 ( .A1(n5433), .A2(n5447), .ZN(n5703) );
  MUX2_X1 U6567 ( .A(n5464), .B(n5449), .S(n5448), .Z(n5451) );
  XNOR2_X1 U6568 ( .A(n5451), .B(n5450), .ZN(n5861) );
  INV_X1 U6569 ( .A(n5706), .ZN(n5453) );
  AOI22_X1 U6570 ( .A1(n6242), .A2(EBX_REG_20__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n6225), .ZN(n5452) );
  OAI21_X1 U6571 ( .B1(n6236), .B2(n5453), .A(n5452), .ZN(n5454) );
  AOI21_X1 U6572 ( .B1(n6202), .B2(n5861), .A(n5454), .ZN(n5458) );
  INV_X1 U6573 ( .A(REIP_REG_19__SCAN_IN), .ZN(n5710) );
  NOR2_X1 U6574 ( .A1(n5472), .A2(n5710), .ZN(n5456) );
  OAI21_X1 U6575 ( .B1(n5456), .B2(REIP_REG_20__SCAN_IN), .A(n5455), .ZN(n5457) );
  OAI211_X1 U6576 ( .C1(n5703), .C2(n6124), .A(n5458), .B(n5457), .ZN(U2807)
         );
  INV_X1 U6577 ( .A(n5460), .ZN(n5461) );
  INV_X1 U6578 ( .A(n5711), .ZN(n5475) );
  INV_X1 U6579 ( .A(n5464), .ZN(n5465) );
  MUX2_X1 U6580 ( .A(n5466), .B(n5465), .S(n2969), .Z(n5481) );
  NOR2_X1 U6581 ( .A1(n5463), .A2(n5481), .ZN(n5480) );
  XOR2_X1 U6582 ( .A(n5467), .B(n5480), .Z(n5872) );
  NAND2_X1 U6583 ( .A1(n5533), .A2(n5468), .ZN(n6219) );
  OAI21_X1 U6584 ( .B1(n6232), .B2(n5469), .A(n6219), .ZN(n5470) );
  AOI21_X1 U6585 ( .B1(n6242), .B2(EBX_REG_19__SCAN_IN), .A(n5470), .ZN(n5471)
         );
  OAI21_X1 U6586 ( .B1(n5872), .B2(n6234), .A(n5471), .ZN(n5474) );
  NOR2_X1 U6587 ( .A1(n5472), .A2(REIP_REG_19__SCAN_IN), .ZN(n5473) );
  AOI211_X1 U6588 ( .C1(n6183), .C2(n5475), .A(n5474), .B(n5473), .ZN(n5478)
         );
  NOR3_X1 U6589 ( .A1(n6123), .A2(REIP_REG_18__SCAN_IN), .A3(n5476), .ZN(n5487) );
  OAI21_X1 U6590 ( .B1(n5487), .B2(n5500), .A(REIP_REG_19__SCAN_IN), .ZN(n5477) );
  OAI211_X1 U6591 ( .C1(n5715), .C2(n6124), .A(n5478), .B(n5477), .ZN(U2808)
         );
  OR2_X1 U6592 ( .A1(n5565), .A2(n5492), .ZN(n5490) );
  AOI21_X1 U6593 ( .B1(n5479), .B2(n5490), .A(n3165), .ZN(n5723) );
  INV_X1 U6594 ( .A(n5723), .ZN(n5627) );
  INV_X1 U6595 ( .A(n5720), .ZN(n5486) );
  AOI21_X1 U6596 ( .B1(n5463), .B2(n5481), .A(n5480), .ZN(n5877) );
  INV_X1 U6597 ( .A(n6242), .ZN(n6178) );
  AOI21_X1 U6598 ( .B1(n6225), .B2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n6181), 
        .ZN(n5482) );
  OAI21_X1 U6599 ( .B1(n6178), .B2(n5483), .A(n5482), .ZN(n5484) );
  AOI21_X1 U6600 ( .B1(n5877), .B2(n6202), .A(n5484), .ZN(n5485) );
  OAI21_X1 U6601 ( .B1(n6236), .B2(n5486), .A(n5485), .ZN(n5488) );
  AOI211_X1 U6602 ( .C1(REIP_REG_18__SCAN_IN), .C2(n5500), .A(n5488), .B(n5487), .ZN(n5489) );
  OAI21_X1 U6603 ( .B1(n5627), .B2(n6124), .A(n5489), .ZN(U2809) );
  INV_X1 U6604 ( .A(n5490), .ZN(n5491) );
  AOI21_X1 U6605 ( .B1(n5492), .B2(n5565), .A(n5491), .ZN(n5729) );
  INV_X1 U6606 ( .A(n5729), .ZN(n5630) );
  INV_X1 U6607 ( .A(n5727), .ZN(n5499) );
  OR2_X1 U6608 ( .A1(n5570), .A2(n5493), .ZN(n5494) );
  NAND2_X1 U6609 ( .A1(n5463), .A2(n5494), .ZN(n5882) );
  OAI21_X1 U6610 ( .B1(n6232), .B2(n5495), .A(n6219), .ZN(n5496) );
  AOI21_X1 U6611 ( .B1(n6242), .B2(EBX_REG_17__SCAN_IN), .A(n5496), .ZN(n5497)
         );
  OAI21_X1 U6612 ( .B1(n5882), .B2(n6234), .A(n5497), .ZN(n5498) );
  AOI21_X1 U6613 ( .B1(n6183), .B2(n5499), .A(n5498), .ZN(n5503) );
  NOR2_X1 U6614 ( .A1(n6123), .A2(n6110), .ZN(n5501) );
  OAI21_X1 U6615 ( .B1(n5501), .B2(REIP_REG_17__SCAN_IN), .A(n5500), .ZN(n5502) );
  OAI211_X1 U6616 ( .C1(n5630), .C2(n6124), .A(n5503), .B(n5502), .ZN(U2810)
         );
  NAND2_X1 U6618 ( .A1(n6217), .A2(n5504), .ZN(n6156) );
  INV_X1 U6619 ( .A(REIP_REG_11__SCAN_IN), .ZN(n6627) );
  NAND2_X1 U6620 ( .A1(REIP_REG_10__SCAN_IN), .A2(REIP_REG_9__SCAN_IN), .ZN(
        n6157) );
  OAI33_X1 U6621 ( .A1(1'b0), .A2(n6156), .A3(n6627), .B1(REIP_REG_11__SCAN_IN), .B2(n6176), .B3(n6157), .ZN(n5506) );
  INV_X1 U6622 ( .A(n5506), .ZN(n5510) );
  AOI22_X1 U6623 ( .A1(n5777), .A2(n6183), .B1(n6202), .B2(n6364), .ZN(n5507)
         );
  OAI211_X1 U6624 ( .C1(n6232), .C2(n5774), .A(n5507), .B(n6219), .ZN(n5508)
         );
  AOI21_X1 U6625 ( .B1(n6242), .B2(EBX_REG_11__SCAN_IN), .A(n5508), .ZN(n5509)
         );
  OAI211_X1 U6626 ( .C1(n5781), .C2(n6124), .A(n5510), .B(n5509), .ZN(U2816)
         );
  INV_X1 U6627 ( .A(n5511), .ZN(n5518) );
  AOI22_X1 U6628 ( .A1(PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n6225), .B1(n6202), 
        .B2(n5512), .ZN(n5513) );
  OAI211_X1 U6629 ( .C1(n6178), .C2(n5514), .A(n5513), .B(n6219), .ZN(n5517)
         );
  NAND2_X1 U6630 ( .A1(n6217), .A2(n5515), .ZN(n6208) );
  AOI22_X1 U6631 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6208), .B1(n6194), .B2(n4850), .ZN(n5516) );
  AOI211_X1 U6632 ( .C1(n6183), .C2(n5518), .A(n5517), .B(n5516), .ZN(n5519)
         );
  OAI21_X1 U6633 ( .B1(n6124), .B2(n5520), .A(n5519), .ZN(U2821) );
  NAND2_X1 U6634 ( .A1(n6216), .A2(n5522), .ZN(n5535) );
  NAND2_X1 U6635 ( .A1(n5535), .A2(n5533), .ZN(n6229) );
  NOR3_X1 U6636 ( .A1(n5523), .A2(REIP_REG_2__SCAN_IN), .A3(n5522), .ZN(n5524)
         );
  AOI21_X1 U6637 ( .B1(n6225), .B2(PHYADDRPOINTER_REG_2__SCAN_IN), .A(n5524), 
        .ZN(n5529) );
  AND2_X1 U6638 ( .A1(n5526), .A2(n5525), .ZN(n6215) );
  AOI22_X1 U6639 ( .A1(n6242), .A2(EBX_REG_2__SCAN_IN), .B1(n6215), .B2(n5527), 
        .ZN(n5528) );
  OAI211_X1 U6640 ( .C1(n6393), .C2(n6234), .A(n5529), .B(n5528), .ZN(n5531)
         );
  NOR2_X1 U6641 ( .A1(n6236), .A2(n6361), .ZN(n5530) );
  AOI211_X1 U6642 ( .C1(REIP_REG_2__SCAN_IN), .C2(n6229), .A(n5531), .B(n5530), 
        .ZN(n5532) );
  OAI21_X1 U6643 ( .B1(n6239), .B2(n6352), .A(n5532), .ZN(U2825) );
  INV_X1 U6644 ( .A(n5533), .ZN(n5534) );
  AOI22_X1 U6645 ( .A1(n6215), .A2(n4515), .B1(n5534), .B2(REIP_REG_1__SCAN_IN), .ZN(n5536) );
  OAI211_X1 U6646 ( .C1(n6178), .C2(n4225), .A(n5536), .B(n5535), .ZN(n5537)
         );
  AOI21_X1 U6647 ( .B1(n6202), .B2(n4488), .A(n5537), .ZN(n5539) );
  MUX2_X1 U6648 ( .A(n6236), .B(n6232), .S(PHYADDRPOINTER_REG_1__SCAN_IN), .Z(
        n5538) );
  OAI211_X1 U6649 ( .C1(n6239), .C2(n5540), .A(n5539), .B(n5538), .ZN(U2826)
         );
  INV_X1 U6650 ( .A(n6215), .ZN(n6233) );
  OAI22_X1 U6651 ( .A1(n5542), .A2(n6178), .B1(n6233), .B2(n5541), .ZN(n5545)
         );
  NOR2_X1 U6652 ( .A1(n6234), .A2(n5543), .ZN(n5544) );
  AOI211_X1 U6653 ( .C1(REIP_REG_0__SCAN_IN), .C2(n6217), .A(n5545), .B(n5544), 
        .ZN(n5547) );
  OAI21_X1 U6654 ( .B1(n6183), .B2(n6225), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n5546) );
  OAI211_X1 U6655 ( .C1(n6239), .C2(n5548), .A(n5547), .B(n5546), .ZN(U2827)
         );
  AOI22_X1 U6656 ( .A1(n5792), .A2(n6247), .B1(EBX_REG_29__SCAN_IN), .B2(n5595), .ZN(n5549) );
  OAI21_X1 U6657 ( .B1(n5645), .B2(n5590), .A(n5549), .ZN(U2830) );
  AOI22_X1 U6658 ( .A1(n5807), .A2(n6247), .B1(EBX_REG_28__SCAN_IN), .B2(n5595), .ZN(n5550) );
  OAI21_X1 U6659 ( .B1(n5602), .B2(n5597), .A(n5550), .ZN(U2831) );
  INV_X1 U6660 ( .A(EBX_REG_27__SCAN_IN), .ZN(n5551) );
  OAI222_X1 U6661 ( .A1(n5597), .A2(n5666), .B1(n5551), .B2(n6250), .C1(n5819), 
        .C2(n5588), .ZN(U2832) );
  INV_X1 U6662 ( .A(EBX_REG_26__SCAN_IN), .ZN(n6801) );
  OAI222_X1 U6663 ( .A1(n5597), .A2(n5607), .B1(n6801), .B2(n6250), .C1(n5824), 
        .C2(n5588), .ZN(U2833) );
  AOI22_X1 U6664 ( .A1(n5832), .A2(n6247), .B1(EBX_REG_25__SCAN_IN), .B2(n5595), .ZN(n5552) );
  OAI21_X1 U6665 ( .B1(n5680), .B2(n5597), .A(n5552), .ZN(U2834) );
  AOI22_X1 U6666 ( .A1(n5553), .A2(n6247), .B1(EBX_REG_24__SCAN_IN), .B2(n5595), .ZN(n5554) );
  OAI21_X1 U6667 ( .B1(n5612), .B2(n5597), .A(n5554), .ZN(U2835) );
  INV_X1 U6668 ( .A(EBX_REG_23__SCAN_IN), .ZN(n5556) );
  OAI222_X1 U6669 ( .A1(n5597), .A2(n5615), .B1(n5556), .B2(n6250), .C1(n5555), 
        .C2(n5588), .ZN(U2836) );
  AOI22_X1 U6670 ( .A1(n5842), .A2(n6247), .B1(EBX_REG_22__SCAN_IN), .B2(n5595), .ZN(n5557) );
  OAI21_X1 U6671 ( .B1(n5618), .B2(n5597), .A(n5557), .ZN(U2837) );
  INV_X1 U6672 ( .A(EBX_REG_21__SCAN_IN), .ZN(n5558) );
  OAI222_X1 U6673 ( .A1(n5700), .A2(n5590), .B1(n5558), .B2(n6250), .C1(n5853), 
        .C2(n5588), .ZN(U2838) );
  AOI22_X1 U6674 ( .A1(n5861), .A2(n6247), .B1(EBX_REG_20__SCAN_IN), .B2(n5595), .ZN(n5559) );
  OAI21_X1 U6675 ( .B1(n5703), .B2(n5597), .A(n5559), .ZN(U2839) );
  INV_X1 U6676 ( .A(EBX_REG_19__SCAN_IN), .ZN(n5560) );
  OAI222_X1 U6677 ( .A1(n5715), .A2(n5590), .B1(n5560), .B2(n6250), .C1(n5588), 
        .C2(n5872), .ZN(U2840) );
  INV_X1 U6678 ( .A(n5877), .ZN(n5561) );
  OAI222_X1 U6679 ( .A1(n5597), .A2(n5627), .B1(n6250), .B2(n5483), .C1(n5561), 
        .C2(n5588), .ZN(U2841) );
  OAI222_X1 U6680 ( .A1(n5597), .A2(n5630), .B1(n5562), .B2(n6250), .C1(n5882), 
        .C2(n5588), .ZN(U2842) );
  INV_X1 U6681 ( .A(n5563), .ZN(n5567) );
  INV_X1 U6682 ( .A(n5564), .ZN(n5566) );
  OAI21_X1 U6683 ( .B1(n5567), .B2(n5566), .A(n5565), .ZN(n6115) );
  INV_X1 U6684 ( .A(EBX_REG_16__SCAN_IN), .ZN(n5572) );
  INV_X1 U6685 ( .A(n5568), .ZN(n5578) );
  AND2_X1 U6686 ( .A1(n5578), .A2(n5569), .ZN(n5571) );
  OR2_X1 U6687 ( .A1(n5571), .A2(n5570), .ZN(n6113) );
  OAI222_X1 U6688 ( .A1(n6115), .A2(n5597), .B1(n6250), .B2(n5572), .C1(n6113), 
        .C2(n5588), .ZN(U2843) );
  XNOR2_X1 U6689 ( .A(n5573), .B(n5574), .ZN(n5752) );
  INV_X1 U6690 ( .A(n5573), .ZN(n5592) );
  AOI22_X1 U6691 ( .A1(n5752), .A2(n5750), .B1(n5592), .B2(n5574), .ZN(n5584)
         );
  INV_X1 U6692 ( .A(n5575), .ZN(n5583) );
  NOR2_X1 U6693 ( .A1(n5584), .A2(n5583), .ZN(n5582) );
  OAI21_X1 U6694 ( .B1(n5582), .B2(n5576), .A(n5563), .ZN(n6125) );
  INV_X1 U6695 ( .A(n5578), .ZN(n5579) );
  AOI21_X1 U6696 ( .B1(n5580), .B2(n5587), .A(n5579), .ZN(n6120) );
  AOI22_X1 U6697 ( .A1(n6120), .A2(n6247), .B1(EBX_REG_15__SCAN_IN), .B2(n5595), .ZN(n5581) );
  OAI21_X1 U6698 ( .B1(n6125), .B2(n5597), .A(n5581), .ZN(U2844) );
  AOI21_X1 U6699 ( .B1(n5584), .B2(n5583), .A(n5582), .ZN(n6134) );
  INV_X1 U6700 ( .A(n6134), .ZN(n5633) );
  INV_X1 U6701 ( .A(EBX_REG_14__SCAN_IN), .ZN(n5589) );
  OR2_X1 U6702 ( .A1(n5929), .A2(n5585), .ZN(n5586) );
  NAND2_X1 U6703 ( .A1(n5587), .A2(n5586), .ZN(n6129) );
  OAI222_X1 U6704 ( .A1(n5633), .A2(n5590), .B1(n6250), .B2(n5589), .C1(n6129), 
        .C2(n5588), .ZN(U2845) );
  INV_X1 U6705 ( .A(n5591), .ZN(n5594) );
  AOI21_X1 U6706 ( .B1(n5594), .B2(n5593), .A(n5592), .ZN(n6153) );
  INV_X1 U6707 ( .A(n6153), .ZN(n5636) );
  XNOR2_X1 U6708 ( .A(n5934), .B(n5930), .ZN(n6147) );
  AOI22_X1 U6709 ( .A1(n6147), .A2(n6247), .B1(EBX_REG_12__SCAN_IN), .B2(n5595), .ZN(n5596) );
  OAI21_X1 U6710 ( .B1(n5636), .B2(n5597), .A(n5596), .ZN(U2847) );
  AOI22_X1 U6711 ( .A1(n6251), .A2(DATAI_29_), .B1(EAX_REG_29__SCAN_IN), .B2(
        n6253), .ZN(n5599) );
  NAND2_X1 U6712 ( .A1(n6254), .A2(DATAI_13_), .ZN(n5598) );
  OAI211_X1 U6713 ( .C1(n5645), .C2(n5635), .A(n5599), .B(n5598), .ZN(U2862)
         );
  AOI22_X1 U6714 ( .A1(n6251), .A2(DATAI_28_), .B1(EAX_REG_28__SCAN_IN), .B2(
        n6253), .ZN(n5601) );
  NAND2_X1 U6715 ( .A1(n6254), .A2(DATAI_12_), .ZN(n5600) );
  OAI211_X1 U6716 ( .C1(n5602), .C2(n5635), .A(n5601), .B(n5600), .ZN(U2863)
         );
  AOI22_X1 U6717 ( .A1(n6251), .A2(DATAI_27_), .B1(EAX_REG_27__SCAN_IN), .B2(
        n6253), .ZN(n5604) );
  NAND2_X1 U6718 ( .A1(n6254), .A2(DATAI_11_), .ZN(n5603) );
  OAI211_X1 U6719 ( .C1(n5666), .C2(n5635), .A(n5604), .B(n5603), .ZN(U2864)
         );
  AOI22_X1 U6720 ( .A1(n6251), .A2(DATAI_26_), .B1(EAX_REG_26__SCAN_IN), .B2(
        n6253), .ZN(n5606) );
  NAND2_X1 U6721 ( .A1(n6254), .A2(DATAI_10_), .ZN(n5605) );
  OAI211_X1 U6722 ( .C1(n5607), .C2(n5635), .A(n5606), .B(n5605), .ZN(U2865)
         );
  AOI22_X1 U6723 ( .A1(n6251), .A2(DATAI_25_), .B1(EAX_REG_25__SCAN_IN), .B2(
        n6253), .ZN(n5609) );
  NAND2_X1 U6724 ( .A1(n6254), .A2(DATAI_9_), .ZN(n5608) );
  OAI211_X1 U6725 ( .C1(n5680), .C2(n5635), .A(n5609), .B(n5608), .ZN(U2866)
         );
  AOI22_X1 U6726 ( .A1(n6251), .A2(DATAI_24_), .B1(EAX_REG_24__SCAN_IN), .B2(
        n6253), .ZN(n5611) );
  NAND2_X1 U6727 ( .A1(n6254), .A2(DATAI_8_), .ZN(n5610) );
  OAI211_X1 U6728 ( .C1(n5612), .C2(n5635), .A(n5611), .B(n5610), .ZN(U2867)
         );
  AOI22_X1 U6729 ( .A1(n6251), .A2(DATAI_23_), .B1(EAX_REG_23__SCAN_IN), .B2(
        n6253), .ZN(n5614) );
  NAND2_X1 U6730 ( .A1(n6254), .A2(DATAI_7_), .ZN(n5613) );
  OAI211_X1 U6731 ( .C1(n5615), .C2(n5635), .A(n5614), .B(n5613), .ZN(U2868)
         );
  AOI22_X1 U6732 ( .A1(n6251), .A2(DATAI_22_), .B1(EAX_REG_22__SCAN_IN), .B2(
        n6253), .ZN(n5617) );
  NAND2_X1 U6733 ( .A1(n6254), .A2(DATAI_6_), .ZN(n5616) );
  OAI211_X1 U6734 ( .C1(n5618), .C2(n5635), .A(n5617), .B(n5616), .ZN(U2869)
         );
  AOI22_X1 U6735 ( .A1(n6251), .A2(DATAI_21_), .B1(EAX_REG_21__SCAN_IN), .B2(
        n6253), .ZN(n5620) );
  NAND2_X1 U6736 ( .A1(n6254), .A2(DATAI_5_), .ZN(n5619) );
  OAI211_X1 U6737 ( .C1(n5700), .C2(n5635), .A(n5620), .B(n5619), .ZN(U2870)
         );
  AOI22_X1 U6738 ( .A1(n6251), .A2(DATAI_20_), .B1(EAX_REG_20__SCAN_IN), .B2(
        n6253), .ZN(n5622) );
  NAND2_X1 U6739 ( .A1(n6254), .A2(DATAI_4_), .ZN(n5621) );
  OAI211_X1 U6740 ( .C1(n5703), .C2(n5635), .A(n5622), .B(n5621), .ZN(U2871)
         );
  AOI22_X1 U6741 ( .A1(n6251), .A2(DATAI_19_), .B1(EAX_REG_19__SCAN_IN), .B2(
        n6253), .ZN(n5624) );
  NAND2_X1 U6742 ( .A1(n6254), .A2(DATAI_3_), .ZN(n5623) );
  OAI211_X1 U6743 ( .C1(n5715), .C2(n5635), .A(n5624), .B(n5623), .ZN(U2872)
         );
  AOI22_X1 U6744 ( .A1(n6251), .A2(DATAI_18_), .B1(EAX_REG_18__SCAN_IN), .B2(
        n6253), .ZN(n5626) );
  NAND2_X1 U6745 ( .A1(n6254), .A2(DATAI_2_), .ZN(n5625) );
  OAI211_X1 U6746 ( .C1(n5627), .C2(n5635), .A(n5626), .B(n5625), .ZN(U2873)
         );
  AOI22_X1 U6747 ( .A1(n6251), .A2(DATAI_17_), .B1(EAX_REG_17__SCAN_IN), .B2(
        n6253), .ZN(n5629) );
  NAND2_X1 U6748 ( .A1(n6254), .A2(DATAI_1_), .ZN(n5628) );
  OAI211_X1 U6749 ( .C1(n5630), .C2(n5635), .A(n5629), .B(n5628), .ZN(U2874)
         );
  AOI22_X1 U6750 ( .A1(n6257), .A2(DATAI_15_), .B1(n6253), .B2(
        EAX_REG_15__SCAN_IN), .ZN(n5631) );
  OAI21_X1 U6751 ( .B1(n6125), .B2(n5635), .A(n5631), .ZN(U2876) );
  AOI22_X1 U6752 ( .A1(n6257), .A2(DATAI_14_), .B1(n6253), .B2(
        EAX_REG_14__SCAN_IN), .ZN(n5632) );
  OAI21_X1 U6753 ( .B1(n5633), .B2(n5635), .A(n5632), .ZN(U2877) );
  AOI22_X1 U6754 ( .A1(n6257), .A2(DATAI_12_), .B1(n6253), .B2(
        EAX_REG_12__SCAN_IN), .ZN(n5634) );
  OAI21_X1 U6755 ( .B1(n5636), .B2(n5635), .A(n5634), .ZN(U2879) );
  INV_X1 U6756 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6656) );
  NOR2_X1 U6757 ( .A1(n6398), .A2(n6656), .ZN(n5796) );
  NOR2_X1 U6758 ( .A1(n5637), .A2(n6362), .ZN(n5638) );
  AOI211_X1 U6759 ( .C1(PHYADDRPOINTER_REG_29__SCAN_IN), .C2(n6351), .A(n5796), 
        .B(n5638), .ZN(n5644) );
  NAND2_X1 U6760 ( .A1(n5640), .A2(n5639), .ZN(n5642) );
  XNOR2_X1 U6761 ( .A(n5642), .B(n5641), .ZN(n5793) );
  NAND2_X1 U6762 ( .A1(n5793), .A2(n4193), .ZN(n5643) );
  OAI211_X1 U6763 ( .C1(n5645), .C2(n5782), .A(n5644), .B(n5643), .ZN(U2957)
         );
  NAND3_X1 U6764 ( .A1(n5671), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .A3(n5760), .ZN(n5651) );
  INV_X1 U6765 ( .A(n5647), .ZN(n5649) );
  NAND3_X1 U6766 ( .A1(n5649), .A2(n5667), .A3(n5648), .ZN(n5661) );
  AOI22_X1 U6767 ( .A1(n5651), .A2(n5661), .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n5650), .ZN(n5652) );
  XNOR2_X1 U6768 ( .A(n5652), .B(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5810)
         );
  NOR2_X1 U6769 ( .A1(n6398), .A2(n6654), .ZN(n5804) );
  AOI21_X1 U6770 ( .B1(n6351), .B2(PHYADDRPOINTER_REG_28__SCAN_IN), .A(n5804), 
        .ZN(n5653) );
  OAI21_X1 U6771 ( .B1(n5654), .B2(n6362), .A(n5653), .ZN(n5655) );
  AOI21_X1 U6772 ( .B1(n5656), .B2(n6358), .A(n5655), .ZN(n5657) );
  OAI21_X1 U6773 ( .B1(n6092), .B2(n5810), .A(n5657), .ZN(U2958) );
  NOR2_X1 U6774 ( .A1(n6398), .A2(n6652), .ZN(n5814) );
  NOR2_X1 U6775 ( .A1(n5658), .A2(n6362), .ZN(n5659) );
  AOI211_X1 U6776 ( .C1(PHYADDRPOINTER_REG_27__SCAN_IN), .C2(n6351), .A(n5814), 
        .B(n5659), .ZN(n5665) );
  INV_X1 U6777 ( .A(n5661), .ZN(n5662) );
  XNOR2_X1 U6778 ( .A(n5663), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5811)
         );
  NAND2_X1 U6779 ( .A1(n5811), .A2(n4193), .ZN(n5664) );
  OAI211_X1 U6780 ( .C1(n5666), .C2(n5782), .A(n5665), .B(n5664), .ZN(U2959)
         );
  INV_X1 U6781 ( .A(n5667), .ZN(n5669) );
  NAND2_X1 U6782 ( .A1(n5669), .A2(n5668), .ZN(n5670) );
  XNOR2_X1 U6783 ( .A(n5671), .B(n5670), .ZN(n5827) );
  INV_X1 U6784 ( .A(REIP_REG_26__SCAN_IN), .ZN(n5672) );
  NOR2_X1 U6785 ( .A1(n6398), .A2(n5672), .ZN(n5820) );
  AOI21_X1 U6786 ( .B1(n6351), .B2(PHYADDRPOINTER_REG_26__SCAN_IN), .A(n5820), 
        .ZN(n5673) );
  OAI21_X1 U6787 ( .B1(n5674), .B2(n6362), .A(n5673), .ZN(n5675) );
  AOI21_X1 U6788 ( .B1(n5676), .B2(n6358), .A(n5675), .ZN(n5677) );
  OAI21_X1 U6789 ( .B1(n5827), .B2(n6092), .A(n5677), .ZN(U2960) );
  AOI21_X1 U6790 ( .B1(n5679), .B2(n5647), .A(n5678), .ZN(n5835) );
  INV_X1 U6791 ( .A(n5680), .ZN(n5684) );
  NOR2_X1 U6792 ( .A1(n6398), .A2(n6650), .ZN(n5830) );
  AOI21_X1 U6793 ( .B1(n6351), .B2(PHYADDRPOINTER_REG_25__SCAN_IN), .A(n5830), 
        .ZN(n5681) );
  OAI21_X1 U6794 ( .B1(n5682), .B2(n6362), .A(n5681), .ZN(n5683) );
  AOI21_X1 U6795 ( .B1(n5684), .B2(n6358), .A(n5683), .ZN(n5685) );
  OAI21_X1 U6796 ( .B1(n5835), .B2(n6092), .A(n5685), .ZN(U2961) );
  XNOR2_X1 U6797 ( .A(n5762), .B(n6783), .ZN(n5687) );
  XNOR2_X1 U6798 ( .A(n5686), .B(n5687), .ZN(n5845) );
  NOR2_X1 U6799 ( .A1(n6398), .A2(n6645), .ZN(n5841) );
  AOI21_X1 U6800 ( .B1(n6351), .B2(PHYADDRPOINTER_REG_22__SCAN_IN), .A(n5841), 
        .ZN(n5688) );
  OAI21_X1 U6801 ( .B1(n5689), .B2(n6362), .A(n5688), .ZN(n5690) );
  AOI21_X1 U6802 ( .B1(n5691), .B2(n6358), .A(n5690), .ZN(n5692) );
  OAI21_X1 U6803 ( .B1(n5845), .B2(n6092), .A(n5692), .ZN(U2964) );
  OAI21_X1 U6804 ( .B1(n5695), .B2(n5694), .A(n5693), .ZN(n5846) );
  NAND2_X1 U6805 ( .A1(n5846), .A2(n4193), .ZN(n5699) );
  NOR2_X1 U6806 ( .A1(n6398), .A2(n6643), .ZN(n5849) );
  NOR2_X1 U6807 ( .A1(n5696), .A2(n6362), .ZN(n5697) );
  AOI211_X1 U6808 ( .C1(n6351), .C2(PHYADDRPOINTER_REG_21__SCAN_IN), .A(n5849), 
        .B(n5697), .ZN(n5698) );
  OAI211_X1 U6809 ( .C1(n5782), .C2(n5700), .A(n5699), .B(n5698), .ZN(U2965)
         );
  XNOR2_X1 U6810 ( .A(n5762), .B(n4380), .ZN(n5701) );
  XNOR2_X1 U6811 ( .A(n3004), .B(n5701), .ZN(n5863) );
  NAND2_X1 U6812 ( .A1(n6350), .A2(REIP_REG_20__SCAN_IN), .ZN(n5857) );
  OAI21_X1 U6813 ( .B1(n5775), .B2(n5702), .A(n5857), .ZN(n5705) );
  NOR2_X1 U6814 ( .A1(n5703), .A2(n5782), .ZN(n5704) );
  AOI211_X1 U6815 ( .C1(n5778), .C2(n5706), .A(n5705), .B(n5704), .ZN(n5707)
         );
  OAI21_X1 U6816 ( .B1(n5863), .B2(n6092), .A(n5707), .ZN(U2966) );
  INV_X1 U6817 ( .A(n5708), .ZN(n5865) );
  NAND2_X1 U6818 ( .A1(n2984), .A2(n5709), .ZN(n5864) );
  NAND3_X1 U6819 ( .A1(n5865), .A2(n4193), .A3(n5864), .ZN(n5714) );
  NOR2_X1 U6820 ( .A1(n6398), .A2(n5710), .ZN(n5868) );
  NOR2_X1 U6821 ( .A1(n5711), .A2(n6362), .ZN(n5712) );
  AOI211_X1 U6822 ( .C1(n6351), .C2(PHYADDRPOINTER_REG_19__SCAN_IN), .A(n5868), 
        .B(n5712), .ZN(n5713) );
  OAI211_X1 U6823 ( .C1(n5782), .C2(n5715), .A(n5714), .B(n5713), .ZN(U2967)
         );
  NOR2_X1 U6824 ( .A1(n5762), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5731)
         );
  NAND2_X1 U6825 ( .A1(n5731), .A2(n5885), .ZN(n5718) );
  NOR2_X1 U6826 ( .A1(n5716), .A2(n5897), .ZN(n5732) );
  NAND2_X1 U6827 ( .A1(n5732), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5717) );
  MUX2_X1 U6828 ( .A(n5718), .B(n5717), .S(n5734), .Z(n5719) );
  XNOR2_X1 U6829 ( .A(n5719), .B(n6714), .ZN(n5879) );
  NAND2_X1 U6830 ( .A1(n5778), .A2(n5720), .ZN(n5721) );
  NAND2_X1 U6831 ( .A1(n6350), .A2(REIP_REG_18__SCAN_IN), .ZN(n5874) );
  OAI211_X1 U6832 ( .C1(n5775), .C2(n3086), .A(n5721), .B(n5874), .ZN(n5722)
         );
  AOI21_X1 U6833 ( .B1(n5723), .B2(n6358), .A(n5722), .ZN(n5724) );
  OAI21_X1 U6834 ( .B1(n5879), .B2(n6092), .A(n5724), .ZN(U2968) );
  MUX2_X1 U6835 ( .A(n5731), .B(n5732), .S(n2973), .Z(n5725) );
  XNOR2_X1 U6836 ( .A(n5725), .B(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5888)
         );
  NAND2_X1 U6837 ( .A1(n6350), .A2(REIP_REG_17__SCAN_IN), .ZN(n5880) );
  NAND2_X1 U6838 ( .A1(n6351), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5726)
         );
  OAI211_X1 U6839 ( .C1(n6362), .C2(n5727), .A(n5880), .B(n5726), .ZN(n5728)
         );
  AOI21_X1 U6840 ( .B1(n5729), .B2(n6358), .A(n5728), .ZN(n5730) );
  OAI21_X1 U6841 ( .B1(n5888), .B2(n6092), .A(n5730), .ZN(U2969) );
  NOR2_X1 U6842 ( .A1(n5732), .A2(n5731), .ZN(n5733) );
  XNOR2_X1 U6843 ( .A(n2973), .B(n5733), .ZN(n5889) );
  NAND2_X1 U6844 ( .A1(n5889), .A2(n4193), .ZN(n5738) );
  AND2_X1 U6845 ( .A1(n6350), .A2(REIP_REG_16__SCAN_IN), .ZN(n5899) );
  NOR2_X1 U6846 ( .A1(n6362), .A2(n5735), .ZN(n5736) );
  AOI211_X1 U6847 ( .C1(n6351), .C2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n5899), 
        .B(n5736), .ZN(n5737) );
  OAI211_X1 U6848 ( .C1(n5782), .C2(n6115), .A(n5738), .B(n5737), .ZN(U2970)
         );
  OR2_X1 U6849 ( .A1(n5740), .A2(n5739), .ZN(n5904) );
  NAND3_X1 U6850 ( .A1(n5904), .A2(n5903), .A3(n4193), .ZN(n5743) );
  NAND2_X1 U6851 ( .A1(n6350), .A2(REIP_REG_15__SCAN_IN), .ZN(n5905) );
  OAI21_X1 U6852 ( .B1(n5775), .B2(n3082), .A(n5905), .ZN(n5741) );
  AOI21_X1 U6853 ( .B1(n5778), .B2(n6121), .A(n5741), .ZN(n5742) );
  OAI211_X1 U6854 ( .C1(n5782), .C2(n6125), .A(n5743), .B(n5742), .ZN(U2971)
         );
  XNOR2_X1 U6855 ( .A(n5762), .B(n5912), .ZN(n5745) );
  XNOR2_X1 U6856 ( .A(n5744), .B(n5745), .ZN(n5928) );
  INV_X1 U6857 ( .A(REIP_REG_14__SCAN_IN), .ZN(n5746) );
  OR2_X1 U6858 ( .A1(n6398), .A2(n5746), .ZN(n5914) );
  NAND2_X1 U6859 ( .A1(n6351), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5747)
         );
  OAI211_X1 U6860 ( .C1(n6362), .C2(n6132), .A(n5914), .B(n5747), .ZN(n5748)
         );
  AOI21_X1 U6861 ( .B1(n6134), .B2(n6358), .A(n5748), .ZN(n5749) );
  OAI21_X1 U6862 ( .B1(n6092), .B2(n5928), .A(n5749), .ZN(U2972) );
  INV_X1 U6863 ( .A(n5750), .ZN(n5751) );
  XNOR2_X1 U6864 ( .A(n5752), .B(n5751), .ZN(n6259) );
  INV_X1 U6865 ( .A(n6259), .ZN(n5759) );
  OAI21_X1 U6866 ( .B1(n5755), .B2(n5754), .A(n5753), .ZN(n5937) );
  NAND2_X1 U6867 ( .A1(n5937), .A2(n4193), .ZN(n5758) );
  NAND2_X1 U6868 ( .A1(n6350), .A2(REIP_REG_13__SCAN_IN), .ZN(n5938) );
  OAI21_X1 U6869 ( .B1(n5775), .B2(n6140), .A(n5938), .ZN(n5756) );
  AOI21_X1 U6870 ( .B1(n5778), .B2(n6142), .A(n5756), .ZN(n5757) );
  OAI211_X1 U6871 ( .C1(n5759), .C2(n5782), .A(n5758), .B(n5757), .ZN(U2973)
         );
  NAND2_X1 U6872 ( .A1(n3002), .A2(n5783), .ZN(n5772) );
  NOR2_X1 U6873 ( .A1(n5760), .A2(n6369), .ZN(n5771) );
  AOI21_X1 U6874 ( .B1(n5772), .B2(n5769), .A(n5771), .ZN(n5764) );
  XNOR2_X1 U6875 ( .A(n5762), .B(n5761), .ZN(n5763) );
  XNOR2_X1 U6876 ( .A(n5764), .B(n5763), .ZN(n5954) );
  INV_X1 U6877 ( .A(n6148), .ZN(n5766) );
  AND2_X1 U6878 ( .A1(n6350), .A2(REIP_REG_12__SCAN_IN), .ZN(n5952) );
  AOI21_X1 U6879 ( .B1(n6351), .B2(PHYADDRPOINTER_REG_12__SCAN_IN), .A(n5952), 
        .ZN(n5765) );
  OAI21_X1 U6880 ( .B1(n5766), .B2(n6362), .A(n5765), .ZN(n5767) );
  AOI21_X1 U6881 ( .B1(n6153), .B2(n6358), .A(n5767), .ZN(n5768) );
  OAI21_X1 U6882 ( .B1(n5954), .B2(n6092), .A(n5768), .ZN(U2974) );
  INV_X1 U6883 ( .A(n5769), .ZN(n5770) );
  NOR2_X1 U6884 ( .A1(n5771), .A2(n5770), .ZN(n5773) );
  XOR2_X1 U6885 ( .A(n5773), .B(n5772), .Z(n6366) );
  NAND2_X1 U6886 ( .A1(n6366), .A2(n4193), .ZN(n5780) );
  NOR2_X1 U6887 ( .A1(n6398), .A2(n6627), .ZN(n6363) );
  NOR2_X1 U6888 ( .A1(n5775), .A2(n5774), .ZN(n5776) );
  AOI211_X1 U6889 ( .C1(n5778), .C2(n5777), .A(n6363), .B(n5776), .ZN(n5779)
         );
  OAI211_X1 U6890 ( .C1(n5782), .C2(n5781), .A(n5780), .B(n5779), .ZN(U2975)
         );
  INV_X1 U6891 ( .A(n5783), .ZN(n5785) );
  NOR2_X1 U6892 ( .A1(n5785), .A2(n5784), .ZN(n5787) );
  XOR2_X1 U6893 ( .A(n5787), .B(n5786), .Z(n5962) );
  INV_X1 U6894 ( .A(n6163), .ZN(n5789) );
  AOI22_X1 U6895 ( .A1(n6351), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .B1(n6350), 
        .B2(REIP_REG_10__SCAN_IN), .ZN(n5788) );
  OAI21_X1 U6896 ( .B1(n6362), .B2(n5789), .A(n5788), .ZN(n5790) );
  AOI21_X1 U6897 ( .B1(n6164), .B2(n6358), .A(n5790), .ZN(n5791) );
  OAI21_X1 U6898 ( .B1(n5962), .B2(n6092), .A(n5791), .ZN(U2976) );
  INV_X1 U6899 ( .A(n5792), .ZN(n5800) );
  NAND2_X1 U6900 ( .A1(n5793), .A2(n6403), .ZN(n5799) );
  NOR2_X1 U6901 ( .A1(n5794), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5795)
         );
  AOI211_X1 U6902 ( .C1(n5797), .C2(INSTADDRPOINTER_REG_29__SCAN_IN), .A(n5796), .B(n5795), .ZN(n5798) );
  OAI211_X1 U6903 ( .C1(n6382), .C2(n5800), .A(n5799), .B(n5798), .ZN(U2989)
         );
  INV_X1 U6904 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5801) );
  NOR2_X1 U6905 ( .A1(n5801), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5805)
         );
  NAND2_X1 U6906 ( .A1(n5806), .A2(n5801), .ZN(n5813) );
  AOI21_X1 U6907 ( .B1(n5812), .B2(n5813), .A(n5802), .ZN(n5803) );
  AOI211_X1 U6908 ( .C1(n5806), .C2(n5805), .A(n5804), .B(n5803), .ZN(n5809)
         );
  NAND2_X1 U6909 ( .A1(n5807), .A2(n6395), .ZN(n5808) );
  OAI211_X1 U6910 ( .C1(n5810), .C2(n5961), .A(n5809), .B(n5808), .ZN(U2990)
         );
  NAND2_X1 U6911 ( .A1(n5811), .A2(n6403), .ZN(n5818) );
  INV_X1 U6912 ( .A(n5812), .ZN(n5816) );
  INV_X1 U6913 ( .A(n5813), .ZN(n5815) );
  AOI211_X1 U6914 ( .C1(n5816), .C2(INSTADDRPOINTER_REG_27__SCAN_IN), .A(n5815), .B(n5814), .ZN(n5817) );
  OAI211_X1 U6915 ( .C1(n6382), .C2(n5819), .A(n5818), .B(n5817), .ZN(U2991)
         );
  XNOR2_X1 U6916 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .B(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5822) );
  INV_X1 U6917 ( .A(n5820), .ZN(n5821) );
  OAI21_X1 U6918 ( .B1(n5828), .B2(n5822), .A(n5821), .ZN(n5823) );
  AOI21_X1 U6919 ( .B1(n5831), .B2(INSTADDRPOINTER_REG_26__SCAN_IN), .A(n5823), 
        .ZN(n5826) );
  OR2_X1 U6920 ( .A1(n5824), .A2(n6382), .ZN(n5825) );
  OAI211_X1 U6921 ( .C1(n5827), .C2(n5961), .A(n5826), .B(n5825), .ZN(U2992)
         );
  NOR2_X1 U6922 ( .A1(n5828), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5829)
         );
  AOI211_X1 U6923 ( .C1(INSTADDRPOINTER_REG_25__SCAN_IN), .C2(n5831), .A(n5830), .B(n5829), .ZN(n5834) );
  NAND2_X1 U6924 ( .A1(n5832), .A2(n6395), .ZN(n5833) );
  OAI211_X1 U6925 ( .C1(n5835), .C2(n5961), .A(n5834), .B(n5833), .ZN(U2993)
         );
  INV_X1 U6926 ( .A(n5836), .ZN(n5850) );
  NAND2_X1 U6927 ( .A1(n5854), .A2(n5837), .ZN(n5847) );
  NOR3_X1 U6928 ( .A1(n5847), .A2(n5839), .A3(n5838), .ZN(n5840) );
  AOI211_X1 U6929 ( .C1(n5850), .C2(INSTADDRPOINTER_REG_22__SCAN_IN), .A(n5841), .B(n5840), .ZN(n5844) );
  NAND2_X1 U6930 ( .A1(n5842), .A2(n6395), .ZN(n5843) );
  OAI211_X1 U6931 ( .C1(n5845), .C2(n5961), .A(n5844), .B(n5843), .ZN(U2996)
         );
  NAND2_X1 U6932 ( .A1(n5846), .A2(n6403), .ZN(n5852) );
  NOR2_X1 U6933 ( .A1(n5847), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5848)
         );
  AOI211_X1 U6934 ( .C1(n5850), .C2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n5849), .B(n5848), .ZN(n5851) );
  OAI211_X1 U6935 ( .C1(n6382), .C2(n5853), .A(n5852), .B(n5851), .ZN(U2997)
         );
  INV_X1 U6936 ( .A(n5854), .ZN(n5866) );
  XNOR2_X1 U6937 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .B(
        INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5859) );
  INV_X1 U6938 ( .A(n5881), .ZN(n5855) );
  AOI21_X1 U6939 ( .B1(n5885), .B2(n5856), .A(n5855), .ZN(n5875) );
  OAI21_X1 U6940 ( .B1(INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n5955), .A(n5875), 
        .ZN(n5869) );
  NAND2_X1 U6941 ( .A1(n5869), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5858) );
  OAI211_X1 U6942 ( .C1(n5866), .C2(n5859), .A(n5858), .B(n5857), .ZN(n5860)
         );
  AOI21_X1 U6943 ( .B1(n5861), .B2(n6395), .A(n5860), .ZN(n5862) );
  OAI21_X1 U6944 ( .B1(n5863), .B2(n5961), .A(n5862), .ZN(U2998) );
  NAND3_X1 U6945 ( .A1(n5865), .A2(n6403), .A3(n5864), .ZN(n5871) );
  NOR2_X1 U6946 ( .A1(n5866), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5867)
         );
  AOI211_X1 U6947 ( .C1(n5869), .C2(INSTADDRPOINTER_REG_19__SCAN_IN), .A(n5868), .B(n5867), .ZN(n5870) );
  OAI211_X1 U6948 ( .C1(n5872), .C2(n6382), .A(n5871), .B(n5870), .ZN(U2999)
         );
  NAND3_X1 U6949 ( .A1(n5886), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .A3(n6714), .ZN(n5873) );
  OAI211_X1 U6950 ( .C1(n5875), .C2(n6714), .A(n5874), .B(n5873), .ZN(n5876)
         );
  AOI21_X1 U6951 ( .B1(n5877), .B2(n6395), .A(n5876), .ZN(n5878) );
  OAI21_X1 U6952 ( .B1(n5879), .B2(n5961), .A(n5878), .ZN(U3000) );
  OAI21_X1 U6953 ( .B1(n5881), .B2(n5885), .A(n5880), .ZN(n5884) );
  NOR2_X1 U6954 ( .A1(n5882), .A2(n6382), .ZN(n5883) );
  AOI211_X1 U6955 ( .C1(n5886), .C2(n5885), .A(n5884), .B(n5883), .ZN(n5887)
         );
  OAI21_X1 U6956 ( .B1(n5888), .B2(n5961), .A(n5887), .ZN(U3001) );
  NAND2_X1 U6957 ( .A1(n5889), .A2(n6403), .ZN(n5902) );
  NOR3_X1 U6958 ( .A1(n5895), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .A3(n5907), 
        .ZN(n5900) );
  INV_X1 U6959 ( .A(n5890), .ZN(n5891) );
  AOI21_X1 U6960 ( .B1(n5892), .B2(n5891), .A(n3000), .ZN(n6370) );
  INV_X1 U6961 ( .A(n6370), .ZN(n5893) );
  AOI21_X1 U6962 ( .B1(n5895), .B2(n5894), .A(n5893), .ZN(n5908) );
  NOR2_X1 U6963 ( .A1(n5895), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5896)
         );
  NAND2_X1 U6964 ( .A1(n6365), .A2(n5896), .ZN(n5906) );
  AOI21_X1 U6965 ( .B1(n5908), .B2(n5906), .A(n5897), .ZN(n5898) );
  AOI211_X1 U6966 ( .C1(n5900), .C2(n6365), .A(n5899), .B(n5898), .ZN(n5901)
         );
  OAI211_X1 U6967 ( .C1(n6382), .C2(n6113), .A(n5902), .B(n5901), .ZN(U3002)
         );
  NAND3_X1 U6968 ( .A1(n5904), .A2(n5903), .A3(n6403), .ZN(n5911) );
  OAI211_X1 U6969 ( .C1(n5908), .C2(n5907), .A(n5906), .B(n5905), .ZN(n5909)
         );
  AOI21_X1 U6970 ( .B1(n6395), .B2(n6120), .A(n5909), .ZN(n5910) );
  NAND2_X1 U6971 ( .A1(n5911), .A2(n5910), .ZN(U3003) );
  NAND3_X1 U6972 ( .A1(n6365), .A2(n5916), .A3(n5912), .ZN(n5913) );
  OAI211_X1 U6973 ( .C1(n6129), .C2(n6382), .A(n5914), .B(n5913), .ZN(n5915)
         );
  INV_X1 U6974 ( .A(n5915), .ZN(n5927) );
  INV_X1 U6975 ( .A(n5947), .ZN(n5921) );
  INV_X1 U6976 ( .A(n5916), .ZN(n5917) );
  NAND2_X1 U6977 ( .A1(n5918), .A2(n5917), .ZN(n5919) );
  OAI211_X1 U6978 ( .C1(n5921), .C2(n5920), .A(n6370), .B(n5919), .ZN(n5942)
         );
  INV_X1 U6979 ( .A(n5922), .ZN(n5923) );
  AOI21_X1 U6980 ( .B1(n5924), .B2(n5923), .A(INSTADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n5925) );
  OAI21_X1 U6981 ( .B1(n5942), .B2(n5925), .A(INSTADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n5926) );
  OAI211_X1 U6982 ( .C1(n5928), .C2(n5961), .A(n5927), .B(n5926), .ZN(U3004)
         );
  INV_X1 U6983 ( .A(n5929), .ZN(n5936) );
  INV_X1 U6984 ( .A(n5930), .ZN(n5933) );
  INV_X1 U6985 ( .A(n5931), .ZN(n5932) );
  OAI21_X1 U6986 ( .B1(n5934), .B2(n5933), .A(n5932), .ZN(n5935) );
  INV_X1 U6987 ( .A(n6246), .ZN(n5945) );
  NAND2_X1 U6988 ( .A1(n5937), .A2(n6403), .ZN(n5944) );
  INV_X1 U6989 ( .A(n5938), .ZN(n5941) );
  INV_X1 U6990 ( .A(n6365), .ZN(n5939) );
  NOR3_X1 U6991 ( .A1(n5939), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .A3(n5947), 
        .ZN(n5940) );
  AOI211_X1 U6992 ( .C1(n5942), .C2(INSTADDRPOINTER_REG_13__SCAN_IN), .A(n5941), .B(n5940), .ZN(n5943) );
  OAI211_X1 U6993 ( .C1(n6382), .C2(n5945), .A(n5944), .B(n5943), .ZN(U3005)
         );
  INV_X1 U6994 ( .A(n5946), .ZN(n5948) );
  OAI21_X1 U6995 ( .B1(n6392), .B2(n5948), .A(n5947), .ZN(n5950) );
  AOI21_X1 U6996 ( .B1(n6365), .B2(INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5949) );
  AOI21_X1 U6997 ( .B1(n6370), .B2(n5950), .A(n5949), .ZN(n5951) );
  AOI211_X1 U6998 ( .C1(n6395), .C2(n6147), .A(n5952), .B(n5951), .ZN(n5953)
         );
  OAI21_X1 U6999 ( .B1(n5954), .B2(n5961), .A(n5953), .ZN(U3006) );
  OAI21_X1 U7000 ( .B1(n5955), .B2(n5956), .A(n6387), .ZN(n6373) );
  INV_X1 U7001 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6625) );
  OAI22_X1 U7002 ( .A1(n6161), .A2(n6382), .B1(n6625), .B2(n6398), .ZN(n5959)
         );
  NAND2_X1 U7003 ( .A1(n5956), .A2(n6378), .ZN(n6377) );
  AOI221_X1 U7004 ( .B1(INSTADDRPOINTER_REG_9__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .C1(n6764), .C2(n5957), .A(n6377), 
        .ZN(n5958) );
  AOI211_X1 U7005 ( .C1(INSTADDRPOINTER_REG_10__SCAN_IN), .C2(n6373), .A(n5959), .B(n5958), .ZN(n5960) );
  OAI21_X1 U7006 ( .B1(n5962), .B2(n5961), .A(n5960), .ZN(U3008) );
  OAI211_X1 U7007 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n2976), .A(n6516), .B(
        n6524), .ZN(n5963) );
  OAI21_X1 U7008 ( .B1(n5970), .B2(n5964), .A(n5963), .ZN(n5965) );
  MUX2_X1 U7009 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n5965), .S(n6408), 
        .Z(U3464) );
  XNOR2_X1 U7010 ( .A(n6516), .B(n5966), .ZN(n5967) );
  OAI22_X1 U7011 ( .A1(n5967), .A2(n6428), .B1(n5970), .B2(n4555), .ZN(n5968)
         );
  MUX2_X1 U7012 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n5968), .S(n6408), 
        .Z(U3463) );
  INV_X1 U7013 ( .A(n4122), .ZN(n5971) );
  OAI222_X1 U7014 ( .A1(n6433), .A2(n5971), .B1(n6474), .B2(n5970), .C1(n6428), 
        .C2(n5969), .ZN(n5972) );
  MUX2_X1 U7015 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n5972), .S(n6408), 
        .Z(U3462) );
  INV_X1 U7016 ( .A(n5973), .ZN(n5974) );
  OAI22_X1 U7017 ( .A1(n5976), .A2(n5975), .B1(n5974), .B2(n6605), .ZN(n5978)
         );
  MUX2_X1 U7018 ( .A(n5978), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n5977), 
        .Z(U3456) );
  NAND2_X1 U7019 ( .A1(n5980), .A2(n5979), .ZN(n5988) );
  INV_X1 U7020 ( .A(n5988), .ZN(n5981) );
  AOI21_X1 U7021 ( .B1(n5981), .B2(STATEBS16_REG_SCAN_IN), .A(n6428), .ZN(
        n5992) );
  INV_X1 U7022 ( .A(n5992), .ZN(n5984) );
  NOR2_X1 U7023 ( .A1(n6429), .A2(n5982), .ZN(n6432) );
  NAND3_X1 U7024 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n3442), .A3(n5983), .ZN(n6431) );
  NOR2_X1 U7025 ( .A1(n6033), .A2(n6431), .ZN(n5989) );
  AOI21_X1 U7026 ( .B1(n6432), .B2(n6519), .A(n5989), .ZN(n5991) );
  OAI22_X1 U7027 ( .A1(n5984), .A2(n5991), .B1(n6431), .B2(n6527), .ZN(n5985)
         );
  NOR2_X2 U7028 ( .A1(n5988), .A2(n5986), .ZN(n6457) );
  INV_X1 U7029 ( .A(n5989), .ZN(n6022) );
  OAI22_X1 U7030 ( .A1(n6440), .A2(n6533), .B1(n6512), .B2(n6022), .ZN(n5990)
         );
  AOI21_X1 U7031 ( .B1(n6480), .B2(n6457), .A(n5990), .ZN(n5996) );
  INV_X1 U7032 ( .A(n6431), .ZN(n5994) );
  NAND2_X1 U7033 ( .A1(n5992), .A2(n5991), .ZN(n5993) );
  NAND2_X1 U7034 ( .A1(n6024), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n5995) );
  OAI211_X1 U7035 ( .C1(n6028), .C2(n5997), .A(n5996), .B(n5995), .ZN(U3060)
         );
  OAI22_X1 U7036 ( .A1(n6440), .A2(n6589), .B1(n6534), .B2(n6022), .ZN(n5998)
         );
  AOI21_X1 U7037 ( .B1(n6586), .B2(n6457), .A(n5998), .ZN(n6000) );
  NAND2_X1 U7038 ( .A1(n6024), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n5999) );
  OAI211_X1 U7039 ( .C1(n6028), .C2(n6001), .A(n6000), .B(n5999), .ZN(U3061)
         );
  OAI22_X1 U7040 ( .A1(n6440), .A2(n6545), .B1(n6539), .B2(n6022), .ZN(n6002)
         );
  AOI21_X1 U7041 ( .B1(n6486), .B2(n6457), .A(n6002), .ZN(n6004) );
  NAND2_X1 U7042 ( .A1(n6024), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n6003) );
  OAI211_X1 U7043 ( .C1(n6028), .C2(n6005), .A(n6004), .B(n6003), .ZN(U3062)
         );
  OAI22_X1 U7044 ( .A1(n6440), .A2(n6552), .B1(n6546), .B2(n6022), .ZN(n6006)
         );
  AOI21_X1 U7045 ( .B1(n6490), .B2(n6457), .A(n6006), .ZN(n6008) );
  NAND2_X1 U7046 ( .A1(n6024), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n6007) );
  OAI211_X1 U7047 ( .C1(n6028), .C2(n6009), .A(n6008), .B(n6007), .ZN(U3063)
         );
  OAI22_X1 U7048 ( .A1(n6440), .A2(n6554), .B1(n6553), .B2(n6022), .ZN(n6010)
         );
  AOI21_X1 U7049 ( .B1(n6494), .B2(n6457), .A(n6010), .ZN(n6012) );
  NAND2_X1 U7050 ( .A1(n6024), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n6011) );
  OAI211_X1 U7051 ( .C1(n6028), .C2(n6013), .A(n6012), .B(n6011), .ZN(U3064)
         );
  OAI22_X1 U7052 ( .A1(n6440), .A2(n6566), .B1(n6560), .B2(n6022), .ZN(n6014)
         );
  AOI21_X1 U7053 ( .B1(n6498), .B2(n6457), .A(n6014), .ZN(n6016) );
  NAND2_X1 U7054 ( .A1(n6024), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n6015) );
  OAI211_X1 U7055 ( .C1(n6028), .C2(n6017), .A(n6016), .B(n6015), .ZN(U3065)
         );
  OAI22_X1 U7056 ( .A1(n6440), .A2(n6854), .B1(n6567), .B2(n6022), .ZN(n6018)
         );
  AOI21_X1 U7057 ( .B1(n6849), .B2(n6457), .A(n6018), .ZN(n6020) );
  NAND2_X1 U7058 ( .A1(n6024), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n6019) );
  OAI211_X1 U7059 ( .C1(n6028), .C2(n6021), .A(n6020), .B(n6019), .ZN(U3066)
         );
  OAI22_X1 U7060 ( .A1(n6440), .A2(n6574), .B1(n6573), .B2(n6022), .ZN(n6023)
         );
  AOI21_X1 U7061 ( .B1(n6507), .B2(n6457), .A(n6023), .ZN(n6026) );
  NAND2_X1 U7062 ( .A1(n6024), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n6025) );
  OAI211_X1 U7063 ( .C1(n6028), .C2(n6027), .A(n6026), .B(n6025), .ZN(U3067)
         );
  INV_X1 U7064 ( .A(n6462), .ZN(n6029) );
  OAI21_X1 U7065 ( .B1(n6457), .B2(n6029), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n6031) );
  NAND3_X1 U7066 ( .A1(n6031), .A2(n6524), .A3(n6030), .ZN(n6037) );
  NAND2_X1 U7067 ( .A1(n6033), .A2(n6032), .ZN(n6042) );
  NAND2_X1 U7068 ( .A1(n6042), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6034) );
  NAND4_X1 U7069 ( .A1(n6037), .A2(n6036), .A3(n6035), .A4(n6034), .ZN(n6459)
         );
  INV_X1 U7070 ( .A(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n6047) );
  NAND3_X1 U7071 ( .A1(n6038), .A2(n6474), .A3(n6515), .ZN(n6041) );
  OR2_X1 U7072 ( .A1(n6427), .A2(n6039), .ZN(n6040) );
  NAND2_X1 U7073 ( .A1(n6041), .A2(n6040), .ZN(n6456) );
  INV_X1 U7074 ( .A(n6042), .ZN(n6455) );
  AOI22_X1 U7075 ( .A1(n6456), .A2(n6585), .B1(n6584), .B2(n6455), .ZN(n6043)
         );
  OAI21_X1 U7076 ( .B1(n6462), .B2(n6538), .A(n6043), .ZN(n6044) );
  AOI21_X1 U7077 ( .B1(n6045), .B2(n6457), .A(n6044), .ZN(n6046) );
  OAI21_X1 U7078 ( .B1(n6074), .B2(n6047), .A(n6046), .ZN(U3069) );
  INV_X1 U7079 ( .A(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n6051) );
  AOI22_X1 U7080 ( .A1(n6456), .A2(n6542), .B1(n6485), .B2(n6455), .ZN(n6048)
         );
  OAI21_X1 U7081 ( .B1(n6462), .B2(n6540), .A(n6048), .ZN(n6049) );
  AOI21_X1 U7082 ( .B1(n6411), .B2(n6457), .A(n6049), .ZN(n6050) );
  OAI21_X1 U7083 ( .B1(n6074), .B2(n6051), .A(n6050), .ZN(U3070) );
  INV_X1 U7084 ( .A(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n6056) );
  AOI22_X1 U7085 ( .A1(n6456), .A2(n6549), .B1(n6489), .B2(n6455), .ZN(n6052)
         );
  OAI21_X1 U7086 ( .B1(n6462), .B2(n6547), .A(n6052), .ZN(n6053) );
  AOI21_X1 U7087 ( .B1(n6054), .B2(n6457), .A(n6053), .ZN(n6055) );
  OAI21_X1 U7088 ( .B1(n6074), .B2(n6056), .A(n6055), .ZN(U3071) );
  INV_X1 U7089 ( .A(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n6060) );
  AOI22_X1 U7090 ( .A1(n6456), .A2(n6556), .B1(n6493), .B2(n6455), .ZN(n6057)
         );
  OAI21_X1 U7091 ( .B1(n6462), .B2(n6559), .A(n6057), .ZN(n6058) );
  AOI21_X1 U7092 ( .B1(n6414), .B2(n6457), .A(n6058), .ZN(n6059) );
  OAI21_X1 U7093 ( .B1(n6074), .B2(n6060), .A(n6059), .ZN(U3072) );
  INV_X1 U7094 ( .A(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n6064) );
  AOI22_X1 U7095 ( .A1(n6456), .A2(n6563), .B1(n6497), .B2(n6455), .ZN(n6061)
         );
  OAI21_X1 U7096 ( .B1(n6462), .B2(n6561), .A(n6061), .ZN(n6062) );
  AOI21_X1 U7097 ( .B1(n6417), .B2(n6457), .A(n6062), .ZN(n6063) );
  OAI21_X1 U7098 ( .B1(n6074), .B2(n6064), .A(n6063), .ZN(U3073) );
  INV_X1 U7099 ( .A(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n6069) );
  AOI22_X1 U7100 ( .A1(n6456), .A2(n6846), .B1(n6845), .B2(n6455), .ZN(n6065)
         );
  OAI21_X1 U7101 ( .B1(n6462), .B2(n6568), .A(n6065), .ZN(n6066) );
  AOI21_X1 U7102 ( .B1(n6067), .B2(n6457), .A(n6066), .ZN(n6068) );
  OAI21_X1 U7103 ( .B1(n6074), .B2(n6069), .A(n6068), .ZN(U3074) );
  INV_X1 U7104 ( .A(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n6073) );
  AOI22_X1 U7105 ( .A1(n6456), .A2(n6578), .B1(n6504), .B2(n6455), .ZN(n6070)
         );
  OAI21_X1 U7106 ( .B1(n6462), .B2(n6582), .A(n6070), .ZN(n6071) );
  AOI21_X1 U7107 ( .B1(n6421), .B2(n6457), .A(n6071), .ZN(n6072) );
  OAI21_X1 U7108 ( .B1(n6074), .B2(n6073), .A(n6072), .ZN(U3075) );
  NOR2_X1 U7109 ( .A1(n6083), .A2(n6075), .ZN(n6078) );
  OAI22_X1 U7110 ( .A1(n6078), .A2(n6077), .B1(n6610), .B2(n6076), .ZN(n6081)
         );
  INV_X1 U7111 ( .A(n6079), .ZN(n6080) );
  NAND3_X1 U7112 ( .A1(n6082), .A2(n6081), .A3(n6080), .ZN(U3182) );
  AND2_X1 U7113 ( .A1(n6286), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  AOI21_X1 U7114 ( .B1(STATE_REG_1__SCAN_IN), .B2(n6610), .A(n6083), .ZN(n6089) );
  INV_X1 U7115 ( .A(ADS_N_REG_SCAN_IN), .ZN(n6084) );
  AOI21_X1 U7116 ( .B1(n6089), .B2(n6084), .A(n6688), .ZN(U2789) );
  OAI21_X1 U7117 ( .B1(n6085), .B2(n6608), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n6086) );
  OAI21_X1 U7118 ( .B1(n6087), .B2(n6603), .A(n6086), .ZN(U2790) );
  NOR2_X1 U7119 ( .A1(STATE_REG_2__SCAN_IN), .A2(STATE_REG_0__SCAN_IN), .ZN(
        n6090) );
  OAI21_X1 U7120 ( .B1(D_C_N_REG_SCAN_IN), .B2(n6090), .A(n6678), .ZN(n6088)
         );
  OAI21_X1 U7121 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n6678), .A(n6088), .ZN(
        U2791) );
  OAI21_X1 U7122 ( .B1(n6090), .B2(BS16_N), .A(n6669), .ZN(n6667) );
  OAI21_X1 U7123 ( .B1(n6669), .B2(n6091), .A(n6667), .ZN(U2792) );
  OAI21_X1 U7124 ( .B1(n6094), .B2(n6093), .A(n6092), .ZN(U2793) );
  NOR4_X1 U7125 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(
        DATAWIDTH_REG_19__SCAN_IN), .A3(DATAWIDTH_REG_20__SCAN_IN), .A4(
        DATAWIDTH_REG_21__SCAN_IN), .ZN(n6098) );
  NOR4_X1 U7126 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(
        DATAWIDTH_REG_15__SCAN_IN), .A3(DATAWIDTH_REG_16__SCAN_IN), .A4(
        DATAWIDTH_REG_17__SCAN_IN), .ZN(n6097) );
  NOR4_X1 U7127 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(
        DATAWIDTH_REG_28__SCAN_IN), .A3(DATAWIDTH_REG_29__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n6096) );
  NOR4_X1 U7128 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(
        DATAWIDTH_REG_23__SCAN_IN), .A3(DATAWIDTH_REG_25__SCAN_IN), .A4(
        DATAWIDTH_REG_26__SCAN_IN), .ZN(n6095) );
  NAND4_X1 U7129 ( .A1(n6098), .A2(n6097), .A3(n6096), .A4(n6095), .ZN(n6104)
         );
  NOR4_X1 U7130 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(
        DATAWIDTH_REG_10__SCAN_IN), .A3(DATAWIDTH_REG_2__SCAN_IN), .A4(
        DATAWIDTH_REG_3__SCAN_IN), .ZN(n6102) );
  AOI211_X1 U7131 ( .C1(DATAWIDTH_REG_1__SCAN_IN), .C2(
        DATAWIDTH_REG_0__SCAN_IN), .A(DATAWIDTH_REG_7__SCAN_IN), .B(
        DATAWIDTH_REG_30__SCAN_IN), .ZN(n6101) );
  NOR4_X1 U7132 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(DATAWIDTH_REG_11__SCAN_IN), .A3(DATAWIDTH_REG_12__SCAN_IN), .A4(DATAWIDTH_REG_13__SCAN_IN), .ZN(n6100)
         );
  NOR4_X1 U7133 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(DATAWIDTH_REG_5__SCAN_IN), 
        .A3(DATAWIDTH_REG_6__SCAN_IN), .A4(DATAWIDTH_REG_8__SCAN_IN), .ZN(
        n6099) );
  NAND4_X1 U7134 ( .A1(n6102), .A2(n6101), .A3(n6100), .A4(n6099), .ZN(n6103)
         );
  NOR2_X1 U7135 ( .A1(n6104), .A2(n6103), .ZN(n6673) );
  INV_X1 U7136 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n6106) );
  NOR3_X1 U7137 ( .A1(REIP_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .A3(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6107) );
  OAI21_X1 U7138 ( .B1(REIP_REG_1__SCAN_IN), .B2(n6107), .A(n6673), .ZN(n6105)
         );
  OAI21_X1 U7139 ( .B1(n6673), .B2(n6106), .A(n6105), .ZN(U2794) );
  INV_X1 U7140 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6668) );
  AOI21_X1 U7141 ( .B1(n5522), .B2(n6668), .A(n6107), .ZN(n6109) );
  INV_X1 U7142 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n6108) );
  INV_X1 U7143 ( .A(n6673), .ZN(n6676) );
  AOI22_X1 U7144 ( .A1(n6673), .A2(n6109), .B1(n6108), .B2(n6676), .ZN(U2795)
         );
  OAI21_X1 U7145 ( .B1(REIP_REG_15__SCAN_IN), .B2(REIP_REG_16__SCAN_IN), .A(
        n6110), .ZN(n6119) );
  AOI22_X1 U7146 ( .A1(EBX_REG_16__SCAN_IN), .A2(n6242), .B1(n6111), .B2(n6183), .ZN(n6112) );
  OAI21_X1 U7147 ( .B1(n6234), .B2(n6113), .A(n6112), .ZN(n6114) );
  AOI211_X1 U7148 ( .C1(n6225), .C2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n6181), 
        .B(n6114), .ZN(n6118) );
  INV_X1 U7149 ( .A(n6115), .ZN(n6252) );
  INV_X1 U7150 ( .A(n6137), .ZN(n6116) );
  AOI22_X1 U7151 ( .A1(n6252), .A2(n6197), .B1(n6116), .B2(
        REIP_REG_16__SCAN_IN), .ZN(n6117) );
  OAI211_X1 U7152 ( .C1(n6123), .C2(n6119), .A(n6118), .B(n6117), .ZN(U2811)
         );
  INV_X1 U7153 ( .A(REIP_REG_15__SCAN_IN), .ZN(n6751) );
  AOI22_X1 U7154 ( .A1(n6121), .A2(n6183), .B1(n6202), .B2(n6120), .ZN(n6122)
         );
  OAI211_X1 U7155 ( .C1(n6232), .C2(n3082), .A(n6122), .B(n6219), .ZN(n6127)
         );
  OAI22_X1 U7156 ( .A1(n6125), .A2(n6124), .B1(REIP_REG_15__SCAN_IN), .B2(
        n6123), .ZN(n6126) );
  AOI211_X1 U7157 ( .C1(EBX_REG_15__SCAN_IN), .C2(n6242), .A(n6127), .B(n6126), 
        .ZN(n6128) );
  OAI21_X1 U7158 ( .B1(n6751), .B2(n6137), .A(n6128), .ZN(U2812) );
  INV_X1 U7159 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6632) );
  INV_X1 U7160 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6629) );
  NOR2_X1 U7161 ( .A1(n6632), .A2(n6629), .ZN(n6143) );
  AOI21_X1 U7162 ( .B1(n6152), .B2(n6143), .A(REIP_REG_14__SCAN_IN), .ZN(n6138) );
  INV_X1 U7163 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n6130) );
  OAI22_X1 U7164 ( .A1(n6130), .A2(n6232), .B1(n6234), .B2(n6129), .ZN(n6131)
         );
  AOI211_X1 U7165 ( .C1(n6242), .C2(EBX_REG_14__SCAN_IN), .A(n6181), .B(n6131), 
        .ZN(n6136) );
  INV_X1 U7166 ( .A(n6132), .ZN(n6133) );
  AOI22_X1 U7167 ( .A1(n6134), .A2(n6197), .B1(n6133), .B2(n6183), .ZN(n6135)
         );
  OAI211_X1 U7168 ( .C1(n6138), .C2(n6137), .A(n6136), .B(n6135), .ZN(U2813)
         );
  AOI22_X1 U7169 ( .A1(EBX_REG_13__SCAN_IN), .A2(n6242), .B1(n6202), .B2(n6246), .ZN(n6139) );
  OAI211_X1 U7170 ( .C1(n6232), .C2(n6140), .A(n6139), .B(n6219), .ZN(n6141)
         );
  AOI21_X1 U7171 ( .B1(n6142), .B2(n6183), .A(n6141), .ZN(n6146) );
  AOI21_X1 U7172 ( .B1(n6632), .B2(n6629), .A(n6143), .ZN(n6144) );
  AOI22_X1 U7173 ( .A1(n6259), .A2(n6197), .B1(n6152), .B2(n6144), .ZN(n6145)
         );
  OAI211_X1 U7174 ( .C1(n6632), .C2(n6156), .A(n6146), .B(n6145), .ZN(U2814)
         );
  AOI22_X1 U7175 ( .A1(n6148), .A2(n6183), .B1(n6202), .B2(n6147), .ZN(n6149)
         );
  OAI211_X1 U7176 ( .C1(n6232), .C2(n6150), .A(n6149), .B(n6219), .ZN(n6151)
         );
  AOI21_X1 U7177 ( .B1(EBX_REG_12__SCAN_IN), .B2(n6242), .A(n6151), .ZN(n6155)
         );
  AOI22_X1 U7178 ( .A1(n6153), .A2(n6197), .B1(n6152), .B2(n6629), .ZN(n6154)
         );
  OAI211_X1 U7179 ( .C1(n6629), .C2(n6156), .A(n6155), .B(n6154), .ZN(U2815)
         );
  OAI21_X1 U7180 ( .B1(REIP_REG_10__SCAN_IN), .B2(REIP_REG_9__SCAN_IN), .A(
        n6157), .ZN(n6167) );
  INV_X1 U7181 ( .A(n6217), .ZN(n6159) );
  NOR2_X1 U7182 ( .A1(n6159), .A2(n6158), .ZN(n6185) );
  AOI22_X1 U7183 ( .A1(EBX_REG_10__SCAN_IN), .A2(n6242), .B1(
        REIP_REG_10__SCAN_IN), .B2(n6185), .ZN(n6160) );
  OAI21_X1 U7184 ( .B1(n6234), .B2(n6161), .A(n6160), .ZN(n6162) );
  AOI211_X1 U7185 ( .C1(n6225), .C2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n6181), 
        .B(n6162), .ZN(n6166) );
  AOI22_X1 U7186 ( .A1(n6164), .A2(n6197), .B1(n6183), .B2(n6163), .ZN(n6165)
         );
  OAI211_X1 U7187 ( .C1(n6176), .C2(n6167), .A(n6166), .B(n6165), .ZN(U2817)
         );
  AOI22_X1 U7188 ( .A1(EBX_REG_9__SCAN_IN), .A2(n6242), .B1(n6202), .B2(n6372), 
        .ZN(n6168) );
  OAI211_X1 U7189 ( .C1(n6232), .C2(n3620), .A(n6168), .B(n6219), .ZN(n6169)
         );
  AOI21_X1 U7190 ( .B1(REIP_REG_9__SCAN_IN), .B2(n6185), .A(n6169), .ZN(n6175)
         );
  INV_X1 U7191 ( .A(n6170), .ZN(n6173) );
  INV_X1 U7192 ( .A(n6171), .ZN(n6172) );
  AOI22_X1 U7193 ( .A1(n6173), .A2(n6197), .B1(n6183), .B2(n6172), .ZN(n6174)
         );
  OAI211_X1 U7194 ( .C1(REIP_REG_9__SCAN_IN), .C2(n6176), .A(n6175), .B(n6174), 
        .ZN(U2818) );
  OAI22_X1 U7195 ( .A1(n6179), .A2(n6178), .B1(n6234), .B2(n6177), .ZN(n6180)
         );
  AOI211_X1 U7196 ( .C1(n6225), .C2(PHYADDRPOINTER_REG_8__SCAN_IN), .A(n6181), 
        .B(n6180), .ZN(n6189) );
  AOI22_X1 U7197 ( .A1(n6197), .A2(n6184), .B1(n6183), .B2(n6182), .ZN(n6188)
         );
  OAI21_X1 U7198 ( .B1(REIP_REG_8__SCAN_IN), .B2(n6186), .A(n6185), .ZN(n6187)
         );
  NAND3_X1 U7199 ( .A1(n6189), .A2(n6188), .A3(n6187), .ZN(U2819) );
  INV_X1 U7200 ( .A(n6381), .ZN(n6190) );
  AOI22_X1 U7201 ( .A1(EBX_REG_7__SCAN_IN), .A2(n6242), .B1(n6202), .B2(n6190), 
        .ZN(n6191) );
  OAI211_X1 U7202 ( .C1(n6232), .C2(n3590), .A(n6191), .B(n6219), .ZN(n6196)
         );
  OAI21_X1 U7203 ( .B1(REIP_REG_7__SCAN_IN), .B2(REIP_REG_6__SCAN_IN), .A(
        n6192), .ZN(n6193) );
  INV_X1 U7204 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6620) );
  OAI22_X1 U7205 ( .A1(n6194), .A2(n6193), .B1(n6620), .B2(n6208), .ZN(n6195)
         );
  AOI211_X1 U7206 ( .C1(n6198), .C2(n6197), .A(n6196), .B(n6195), .ZN(n6199)
         );
  OAI21_X1 U7207 ( .B1(n6200), .B2(n6236), .A(n6199), .ZN(U2820) );
  INV_X1 U7208 ( .A(n6239), .ZN(n6207) );
  AOI22_X1 U7209 ( .A1(EBX_REG_5__SCAN_IN), .A2(n6242), .B1(n6202), .B2(n6201), 
        .ZN(n6203) );
  OAI211_X1 U7210 ( .C1(n6232), .C2(n6204), .A(n6203), .B(n6219), .ZN(n6205)
         );
  AOI21_X1 U7211 ( .B1(n6207), .B2(n6206), .A(n6205), .ZN(n6212) );
  INV_X1 U7212 ( .A(n6208), .ZN(n6209) );
  OAI21_X1 U7213 ( .B1(REIP_REG_5__SCAN_IN), .B2(n6210), .A(n6209), .ZN(n6211)
         );
  OAI211_X1 U7214 ( .C1(n6236), .C2(n6213), .A(n6212), .B(n6211), .ZN(U2822)
         );
  AOI22_X1 U7215 ( .A1(n6242), .A2(EBX_REG_4__SCAN_IN), .B1(n6215), .B2(n6214), 
        .ZN(n6227) );
  NAND4_X1 U7216 ( .A1(n6216), .A2(REIP_REG_1__SCAN_IN), .A3(
        REIP_REG_2__SCAN_IN), .A4(REIP_REG_3__SCAN_IN), .ZN(n6220) );
  NAND2_X1 U7217 ( .A1(n6218), .A2(n6217), .ZN(n6245) );
  OAI221_X1 U7218 ( .B1(REIP_REG_4__SCAN_IN), .B2(n6220), .C1(n6616), .C2(
        n6245), .A(n6219), .ZN(n6224) );
  OAI22_X1 U7219 ( .A1(n6239), .A2(n6222), .B1(n6221), .B2(n6236), .ZN(n6223)
         );
  AOI211_X1 U7220 ( .C1(PHYADDRPOINTER_REG_4__SCAN_IN), .C2(n6225), .A(n6224), 
        .B(n6223), .ZN(n6226) );
  OAI211_X1 U7221 ( .C1(n6234), .C2(n6228), .A(n6227), .B(n6226), .ZN(U2823)
         );
  INV_X1 U7222 ( .A(n6229), .ZN(n6230) );
  NAND2_X1 U7223 ( .A1(n6230), .A2(REIP_REG_2__SCAN_IN), .ZN(n6244) );
  INV_X1 U7224 ( .A(n6231), .ZN(n6235) );
  OAI222_X1 U7225 ( .A1(n6235), .A2(n6234), .B1(n6233), .B2(n6474), .C1(n6232), 
        .C2(n3079), .ZN(n6241) );
  OAI22_X1 U7226 ( .A1(n6239), .A2(n6238), .B1(n6237), .B2(n6236), .ZN(n6240)
         );
  AOI211_X1 U7227 ( .C1(EBX_REG_3__SCAN_IN), .C2(n6242), .A(n6241), .B(n6240), 
        .ZN(n6243) );
  OAI221_X1 U7228 ( .B1(n6245), .B2(n6614), .C1(n6245), .C2(n6244), .A(n6243), 
        .ZN(U2824) );
  AOI22_X1 U7229 ( .A1(n6259), .A2(n6248), .B1(n6247), .B2(n6246), .ZN(n6249)
         );
  OAI21_X1 U7230 ( .B1(n6250), .B2(n6808), .A(n6249), .ZN(U2846) );
  AOI22_X1 U7231 ( .A1(n6252), .A2(n6258), .B1(n6251), .B2(DATAI_16_), .ZN(
        n6256) );
  AOI22_X1 U7232 ( .A1(n6254), .A2(DATAI_0_), .B1(n6253), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n6255) );
  NAND2_X1 U7233 ( .A1(n6256), .A2(n6255), .ZN(U2875) );
  AOI22_X1 U7234 ( .A1(n6259), .A2(n6258), .B1(DATAI_13_), .B2(n6257), .ZN(
        n6260) );
  OAI21_X1 U7235 ( .B1(n6268), .B2(n6261), .A(n6260), .ZN(U2878) );
  INV_X1 U7236 ( .A(DATAO_REG_25__SCAN_IN), .ZN(n6743) );
  AOI22_X1 U7237 ( .A1(n6263), .A2(EAX_REG_25__SCAN_IN), .B1(n6681), .B2(
        UWORD_REG_9__SCAN_IN), .ZN(n6262) );
  OAI21_X1 U7238 ( .B1(n6743), .B2(n6281), .A(n6262), .ZN(U2898) );
  AOI22_X1 U7239 ( .A1(n6286), .A2(DATAO_REG_18__SCAN_IN), .B1(
        EAX_REG_18__SCAN_IN), .B2(n6263), .ZN(n6264) );
  OAI21_X1 U7240 ( .B1(n6823), .B2(n6280), .A(n6264), .ZN(U2905) );
  INV_X1 U7241 ( .A(EAX_REG_15__SCAN_IN), .ZN(n6349) );
  AOI22_X1 U7242 ( .A1(n6681), .A2(LWORD_REG_15__SCAN_IN), .B1(n6286), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6265) );
  OAI21_X1 U7243 ( .B1(n6349), .B2(n6288), .A(n6265), .ZN(U2908) );
  INV_X1 U7244 ( .A(DATAO_REG_14__SCAN_IN), .ZN(n6762) );
  AOI22_X1 U7245 ( .A1(EAX_REG_14__SCAN_IN), .A2(n6274), .B1(n6681), .B2(
        LWORD_REG_14__SCAN_IN), .ZN(n6266) );
  OAI21_X1 U7246 ( .B1(n6762), .B2(n6281), .A(n6266), .ZN(U2909) );
  AOI22_X1 U7247 ( .A1(n6681), .A2(LWORD_REG_13__SCAN_IN), .B1(n6286), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n6267) );
  OAI21_X1 U7248 ( .B1(n6268), .B2(n6288), .A(n6267), .ZN(U2910) );
  INV_X1 U7249 ( .A(EAX_REG_12__SCAN_IN), .ZN(n6765) );
  AOI22_X1 U7250 ( .A1(n6681), .A2(LWORD_REG_12__SCAN_IN), .B1(n6286), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6269) );
  OAI21_X1 U7251 ( .B1(n6765), .B2(n6288), .A(n6269), .ZN(U2911) );
  INV_X1 U7252 ( .A(EAX_REG_11__SCAN_IN), .ZN(n6753) );
  AOI22_X1 U7253 ( .A1(n6681), .A2(LWORD_REG_11__SCAN_IN), .B1(n6286), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n6270) );
  OAI21_X1 U7254 ( .B1(n6753), .B2(n6288), .A(n6270), .ZN(U2912) );
  INV_X1 U7255 ( .A(EAX_REG_10__SCAN_IN), .ZN(n6272) );
  AOI22_X1 U7256 ( .A1(n6681), .A2(LWORD_REG_10__SCAN_IN), .B1(n6286), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n6271) );
  OAI21_X1 U7257 ( .B1(n6272), .B2(n6288), .A(n6271), .ZN(U2913) );
  INV_X1 U7258 ( .A(LWORD_REG_9__SCAN_IN), .ZN(n6750) );
  AOI22_X1 U7259 ( .A1(EAX_REG_9__SCAN_IN), .A2(n6274), .B1(n6286), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n6273) );
  OAI21_X1 U7260 ( .B1(n6750), .B2(n6280), .A(n6273), .ZN(U2914) );
  INV_X1 U7261 ( .A(DATAO_REG_8__SCAN_IN), .ZN(n6737) );
  AOI22_X1 U7262 ( .A1(EAX_REG_8__SCAN_IN), .A2(n6274), .B1(n6681), .B2(
        LWORD_REG_8__SCAN_IN), .ZN(n6275) );
  OAI21_X1 U7263 ( .B1(n6737), .B2(n6281), .A(n6275), .ZN(U2915) );
  INV_X1 U7264 ( .A(EAX_REG_7__SCAN_IN), .ZN(n6277) );
  AOI22_X1 U7265 ( .A1(n6681), .A2(LWORD_REG_7__SCAN_IN), .B1(n6286), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n6276) );
  OAI21_X1 U7266 ( .B1(n6277), .B2(n6288), .A(n6276), .ZN(U2916) );
  AOI22_X1 U7267 ( .A1(n6681), .A2(LWORD_REG_6__SCAN_IN), .B1(n6286), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n6278) );
  OAI21_X1 U7268 ( .B1(n3510), .B2(n6288), .A(n6278), .ZN(U2917) );
  INV_X1 U7269 ( .A(DATAO_REG_5__SCAN_IN), .ZN(n6745) );
  INV_X1 U7270 ( .A(LWORD_REG_5__SCAN_IN), .ZN(n6279) );
  OAI222_X1 U7271 ( .A1(n6281), .A2(n6745), .B1(n6288), .B2(n6826), .C1(n6280), 
        .C2(n6279), .ZN(U2918) );
  AOI22_X1 U7272 ( .A1(n6681), .A2(LWORD_REG_4__SCAN_IN), .B1(n6286), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n6282) );
  OAI21_X1 U7273 ( .B1(n6327), .B2(n6288), .A(n6282), .ZN(U2919) );
  AOI22_X1 U7274 ( .A1(n6681), .A2(LWORD_REG_3__SCAN_IN), .B1(n6286), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n6283) );
  OAI21_X1 U7275 ( .B1(n6324), .B2(n6288), .A(n6283), .ZN(U2920) );
  AOI22_X1 U7276 ( .A1(n6681), .A2(LWORD_REG_2__SCAN_IN), .B1(n6286), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n6284) );
  OAI21_X1 U7277 ( .B1(n6321), .B2(n6288), .A(n6284), .ZN(U2921) );
  AOI22_X1 U7278 ( .A1(n6681), .A2(LWORD_REG_1__SCAN_IN), .B1(n6286), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n6285) );
  OAI21_X1 U7279 ( .B1(n6318), .B2(n6288), .A(n6285), .ZN(U2922) );
  AOI22_X1 U7280 ( .A1(n6681), .A2(LWORD_REG_0__SCAN_IN), .B1(n6286), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n6287) );
  OAI21_X1 U7281 ( .B1(n6315), .B2(n6288), .A(n6287), .ZN(U2923) );
  INV_X1 U7282 ( .A(EAX_REG_16__SCAN_IN), .ZN(n6744) );
  AND2_X1 U7283 ( .A1(n6346), .A2(DATAI_0_), .ZN(n6313) );
  AOI21_X1 U7284 ( .B1(UWORD_REG_0__SCAN_IN), .B2(n6332), .A(n6313), .ZN(n6289) );
  OAI21_X1 U7285 ( .B1(n6744), .B2(n6348), .A(n6289), .ZN(U2924) );
  INV_X1 U7286 ( .A(EAX_REG_17__SCAN_IN), .ZN(n6291) );
  AND2_X1 U7287 ( .A1(n6346), .A2(DATAI_1_), .ZN(n6316) );
  AOI21_X1 U7288 ( .B1(UWORD_REG_1__SCAN_IN), .B2(n6332), .A(n6316), .ZN(n6290) );
  OAI21_X1 U7289 ( .B1(n6291), .B2(n6348), .A(n6290), .ZN(U2925) );
  INV_X1 U7290 ( .A(EAX_REG_19__SCAN_IN), .ZN(n6792) );
  AND2_X1 U7291 ( .A1(n6346), .A2(DATAI_3_), .ZN(n6322) );
  AOI21_X1 U7292 ( .B1(UWORD_REG_3__SCAN_IN), .B2(n6332), .A(n6322), .ZN(n6292) );
  OAI21_X1 U7293 ( .B1(n6792), .B2(n6348), .A(n6292), .ZN(U2927) );
  INV_X1 U7294 ( .A(EAX_REG_20__SCAN_IN), .ZN(n6294) );
  AND2_X1 U7295 ( .A1(n6346), .A2(DATAI_4_), .ZN(n6325) );
  AOI21_X1 U7296 ( .B1(UWORD_REG_4__SCAN_IN), .B2(n6332), .A(n6325), .ZN(n6293) );
  OAI21_X1 U7297 ( .B1(n6294), .B2(n6348), .A(n6293), .ZN(U2928) );
  AND2_X1 U7298 ( .A1(n6346), .A2(DATAI_5_), .ZN(n6328) );
  AOI21_X1 U7299 ( .B1(UWORD_REG_5__SCAN_IN), .B2(n6332), .A(n6328), .ZN(n6295) );
  OAI21_X1 U7300 ( .B1(n6296), .B2(n6348), .A(n6295), .ZN(U2929) );
  INV_X1 U7301 ( .A(EAX_REG_22__SCAN_IN), .ZN(n6795) );
  AND2_X1 U7302 ( .A1(n6346), .A2(DATAI_6_), .ZN(n6330) );
  AOI21_X1 U7303 ( .B1(UWORD_REG_6__SCAN_IN), .B2(n6332), .A(n6330), .ZN(n6297) );
  OAI21_X1 U7304 ( .B1(n6795), .B2(n6348), .A(n6297), .ZN(U2930) );
  INV_X1 U7305 ( .A(EAX_REG_23__SCAN_IN), .ZN(n6300) );
  AOI22_X1 U7306 ( .A1(UWORD_REG_7__SCAN_IN), .A2(n4432), .B1(n6346), .B2(
        DATAI_7_), .ZN(n6299) );
  OAI21_X1 U7307 ( .B1(n6300), .B2(n6348), .A(n6299), .ZN(U2931) );
  NAND2_X1 U7308 ( .A1(n6346), .A2(DATAI_8_), .ZN(n6333) );
  INV_X1 U7309 ( .A(n6333), .ZN(n6301) );
  AOI21_X1 U7310 ( .B1(UWORD_REG_8__SCAN_IN), .B2(n6332), .A(n6301), .ZN(n6302) );
  OAI21_X1 U7311 ( .B1(n6736), .B2(n6348), .A(n6302), .ZN(U2932) );
  AOI22_X1 U7312 ( .A1(n6332), .A2(UWORD_REG_9__SCAN_IN), .B1(
        EAX_REG_25__SCAN_IN), .B2(n6343), .ZN(n6303) );
  NAND2_X1 U7313 ( .A1(n6346), .A2(DATAI_9_), .ZN(n6335) );
  NAND2_X1 U7314 ( .A1(n6303), .A2(n6335), .ZN(U2933) );
  NAND2_X1 U7315 ( .A1(n6346), .A2(DATAI_10_), .ZN(n6337) );
  INV_X1 U7316 ( .A(n6337), .ZN(n6304) );
  AOI21_X1 U7317 ( .B1(UWORD_REG_10__SCAN_IN), .B2(n6332), .A(n6304), .ZN(
        n6305) );
  OAI21_X1 U7318 ( .B1(n3927), .B2(n6348), .A(n6305), .ZN(U2934) );
  INV_X1 U7319 ( .A(DATAI_12_), .ZN(n6306) );
  NOR2_X1 U7320 ( .A1(n6307), .A2(n6306), .ZN(n6341) );
  AOI21_X1 U7321 ( .B1(UWORD_REG_12__SCAN_IN), .B2(n6332), .A(n6341), .ZN(
        n6308) );
  OAI21_X1 U7322 ( .B1(n3969), .B2(n6348), .A(n6308), .ZN(U2936) );
  INV_X1 U7323 ( .A(EAX_REG_29__SCAN_IN), .ZN(n6310) );
  AOI22_X1 U7324 ( .A1(UWORD_REG_13__SCAN_IN), .A2(n4432), .B1(n6346), .B2(
        DATAI_13_), .ZN(n6309) );
  OAI21_X1 U7325 ( .B1(n6310), .B2(n6348), .A(n6309), .ZN(U2937) );
  NAND2_X1 U7326 ( .A1(n6346), .A2(DATAI_14_), .ZN(n6344) );
  INV_X1 U7327 ( .A(n6344), .ZN(n6311) );
  AOI21_X1 U7328 ( .B1(UWORD_REG_14__SCAN_IN), .B2(n6332), .A(n6311), .ZN(
        n6312) );
  OAI21_X1 U7329 ( .B1(n4017), .B2(n6348), .A(n6312), .ZN(U2938) );
  AOI21_X1 U7330 ( .B1(LWORD_REG_0__SCAN_IN), .B2(n4432), .A(n6313), .ZN(n6314) );
  OAI21_X1 U7331 ( .B1(n6315), .B2(n6348), .A(n6314), .ZN(U2939) );
  AOI21_X1 U7332 ( .B1(LWORD_REG_1__SCAN_IN), .B2(n4432), .A(n6316), .ZN(n6317) );
  OAI21_X1 U7333 ( .B1(n6318), .B2(n6348), .A(n6317), .ZN(U2940) );
  AOI21_X1 U7334 ( .B1(LWORD_REG_2__SCAN_IN), .B2(n4432), .A(n6319), .ZN(n6320) );
  OAI21_X1 U7335 ( .B1(n6321), .B2(n6348), .A(n6320), .ZN(U2941) );
  AOI21_X1 U7336 ( .B1(LWORD_REG_3__SCAN_IN), .B2(n4432), .A(n6322), .ZN(n6323) );
  OAI21_X1 U7337 ( .B1(n6324), .B2(n6348), .A(n6323), .ZN(U2942) );
  AOI21_X1 U7338 ( .B1(LWORD_REG_4__SCAN_IN), .B2(n4432), .A(n6325), .ZN(n6326) );
  OAI21_X1 U7339 ( .B1(n6327), .B2(n6348), .A(n6326), .ZN(U2943) );
  AOI21_X1 U7340 ( .B1(LWORD_REG_5__SCAN_IN), .B2(n6332), .A(n6328), .ZN(n6329) );
  OAI21_X1 U7341 ( .B1(n6826), .B2(n6348), .A(n6329), .ZN(U2944) );
  AOI21_X1 U7342 ( .B1(LWORD_REG_6__SCAN_IN), .B2(n6332), .A(n6330), .ZN(n6331) );
  OAI21_X1 U7343 ( .B1(n3510), .B2(n6348), .A(n6331), .ZN(U2945) );
  AOI22_X1 U7344 ( .A1(n6332), .A2(LWORD_REG_8__SCAN_IN), .B1(
        EAX_REG_8__SCAN_IN), .B2(n6343), .ZN(n6334) );
  NAND2_X1 U7345 ( .A1(n6334), .A2(n6333), .ZN(U2947) );
  AOI22_X1 U7346 ( .A1(n6332), .A2(LWORD_REG_9__SCAN_IN), .B1(
        EAX_REG_9__SCAN_IN), .B2(n6343), .ZN(n6336) );
  NAND2_X1 U7347 ( .A1(n6336), .A2(n6335), .ZN(U2948) );
  AOI22_X1 U7348 ( .A1(n6332), .A2(LWORD_REG_10__SCAN_IN), .B1(
        EAX_REG_10__SCAN_IN), .B2(n6343), .ZN(n6338) );
  NAND2_X1 U7349 ( .A1(n6338), .A2(n6337), .ZN(U2949) );
  AOI21_X1 U7350 ( .B1(LWORD_REG_11__SCAN_IN), .B2(n4432), .A(n6339), .ZN(
        n6340) );
  OAI21_X1 U7351 ( .B1(n6753), .B2(n6348), .A(n6340), .ZN(U2950) );
  AOI21_X1 U7352 ( .B1(LWORD_REG_12__SCAN_IN), .B2(n4432), .A(n6341), .ZN(
        n6342) );
  OAI21_X1 U7353 ( .B1(n6765), .B2(n6348), .A(n6342), .ZN(U2951) );
  AOI22_X1 U7354 ( .A1(n6332), .A2(LWORD_REG_14__SCAN_IN), .B1(
        EAX_REG_14__SCAN_IN), .B2(n6343), .ZN(n6345) );
  NAND2_X1 U7355 ( .A1(n6345), .A2(n6344), .ZN(U2953) );
  AOI22_X1 U7356 ( .A1(LWORD_REG_15__SCAN_IN), .A2(n4432), .B1(n6346), .B2(
        DATAI_15_), .ZN(n6347) );
  OAI21_X1 U7357 ( .B1(n6349), .B2(n6348), .A(n6347), .ZN(U2954) );
  AOI22_X1 U7358 ( .A1(n6351), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .B1(n6350), 
        .B2(REIP_REG_2__SCAN_IN), .ZN(n6360) );
  INV_X1 U7359 ( .A(n6352), .ZN(n6357) );
  NAND2_X1 U7360 ( .A1(n6354), .A2(n6353), .ZN(n6355) );
  XOR2_X1 U7361 ( .A(n6356), .B(n6355), .Z(n6404) );
  AOI22_X1 U7362 ( .A1(n6358), .A2(n6357), .B1(n6404), .B2(n4193), .ZN(n6359)
         );
  OAI211_X1 U7363 ( .C1(n6362), .C2(n6361), .A(n6360), .B(n6359), .ZN(U2984)
         );
  AOI21_X1 U7364 ( .B1(n6364), .B2(n6395), .A(n6363), .ZN(n6368) );
  AOI22_X1 U7365 ( .A1(n6366), .A2(n6403), .B1(n6369), .B2(n6365), .ZN(n6367)
         );
  OAI211_X1 U7366 ( .C1(n6370), .C2(n6369), .A(n6368), .B(n6367), .ZN(U3007)
         );
  AOI21_X1 U7367 ( .B1(n6372), .B2(n6395), .A(n6371), .ZN(n6376) );
  AOI22_X1 U7368 ( .A1(n6374), .A2(n6403), .B1(INSTADDRPOINTER_REG_9__SCAN_IN), 
        .B2(n6373), .ZN(n6375) );
  OAI211_X1 U7369 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n6377), .A(n6376), 
        .B(n6375), .ZN(U3009) );
  NAND2_X1 U7370 ( .A1(n6378), .A2(n6386), .ZN(n6380) );
  OAI211_X1 U7371 ( .C1(n6382), .C2(n6381), .A(n6380), .B(n6379), .ZN(n6383)
         );
  AOI21_X1 U7372 ( .B1(n6384), .B2(n6403), .A(n6383), .ZN(n6385) );
  OAI21_X1 U7373 ( .B1(n6387), .B2(n6386), .A(n6385), .ZN(U3011) );
  INV_X1 U7374 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6612) );
  OAI21_X1 U7375 ( .B1(n6390), .B2(n6389), .A(n6388), .ZN(n6391) );
  NAND2_X1 U7376 ( .A1(n6392), .A2(n6391), .ZN(n6397) );
  INV_X1 U7377 ( .A(n6393), .ZN(n6394) );
  NAND2_X1 U7378 ( .A1(n6395), .A2(n6394), .ZN(n6396) );
  OAI211_X1 U7379 ( .C1(n6612), .C2(n6398), .A(n6397), .B(n6396), .ZN(n6399)
         );
  INV_X1 U7380 ( .A(n6399), .ZN(n6406) );
  NOR2_X1 U7381 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n6400), .ZN(n6401)
         );
  AOI22_X1 U7382 ( .A1(n6404), .A2(n6403), .B1(n6402), .B2(n6401), .ZN(n6405)
         );
  OAI211_X1 U7383 ( .C1(n6407), .C2(n4119), .A(n6406), .B(n6405), .ZN(U3016)
         );
  NOR2_X1 U7384 ( .A1(n6409), .A2(n6408), .ZN(U3019) );
  INV_X1 U7385 ( .A(n6410), .ZN(n6420) );
  AOI22_X1 U7386 ( .A1(n6422), .A2(n6411), .B1(n6485), .B2(n6420), .ZN(n6413)
         );
  AOI22_X1 U7387 ( .A1(INSTQUEUE_REG_3__2__SCAN_IN), .A2(n6424), .B1(n6542), 
        .B2(n6423), .ZN(n6412) );
  OAI211_X1 U7388 ( .C1(n6540), .C2(n6853), .A(n6413), .B(n6412), .ZN(U3046)
         );
  AOI22_X1 U7389 ( .A1(n6422), .A2(n6414), .B1(n6493), .B2(n6420), .ZN(n6416)
         );
  AOI22_X1 U7390 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n6424), .B1(n6556), 
        .B2(n6423), .ZN(n6415) );
  OAI211_X1 U7391 ( .C1(n6559), .C2(n6853), .A(n6416), .B(n6415), .ZN(U3048)
         );
  AOI22_X1 U7392 ( .A1(n6422), .A2(n6417), .B1(n6497), .B2(n6420), .ZN(n6419)
         );
  AOI22_X1 U7393 ( .A1(INSTQUEUE_REG_3__5__SCAN_IN), .A2(n6424), .B1(n6563), 
        .B2(n6423), .ZN(n6418) );
  OAI211_X1 U7394 ( .C1(n6561), .C2(n6853), .A(n6419), .B(n6418), .ZN(U3049)
         );
  AOI22_X1 U7395 ( .A1(n6422), .A2(n6421), .B1(n6504), .B2(n6420), .ZN(n6426)
         );
  AOI22_X1 U7396 ( .A1(INSTQUEUE_REG_3__7__SCAN_IN), .A2(n6424), .B1(n6578), 
        .B2(n6423), .ZN(n6425) );
  OAI211_X1 U7397 ( .C1(n6582), .C2(n6853), .A(n6426), .B(n6425), .ZN(U3051)
         );
  OAI33_X1 U7398 ( .A1(n6430), .A2(n6429), .A3(n6428), .B1(n6464), .B2(n6427), 
        .B3(n6467), .ZN(n6847) );
  NOR2_X1 U7399 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6431), .ZN(n6844)
         );
  AOI22_X1 U7400 ( .A1(n3024), .A2(n6530), .B1(n6470), .B2(n6844), .ZN(n6442)
         );
  NAND3_X1 U7401 ( .A1(n6853), .A2(n6524), .A3(n6440), .ZN(n6434) );
  AOI21_X1 U7402 ( .B1(n6434), .B2(n6433), .A(n6432), .ZN(n6439) );
  OAI211_X1 U7403 ( .C1(n6844), .C2(n6437), .A(n6436), .B(n6435), .ZN(n6438)
         );
  AOI22_X1 U7404 ( .A1(n6850), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n6480), 
        .B2(n6848), .ZN(n6441) );
  OAI211_X1 U7405 ( .C1(n6533), .C2(n6853), .A(n6442), .B(n6441), .ZN(U3052)
         );
  AOI22_X1 U7406 ( .A1(n3024), .A2(n6585), .B1(n6584), .B2(n6844), .ZN(n6444)
         );
  AOI22_X1 U7407 ( .A1(n6850), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n6586), 
        .B2(n6848), .ZN(n6443) );
  OAI211_X1 U7408 ( .C1(n6589), .C2(n6853), .A(n6444), .B(n6443), .ZN(U3053)
         );
  AOI22_X1 U7409 ( .A1(n3024), .A2(n6542), .B1(n6485), .B2(n6844), .ZN(n6446)
         );
  AOI22_X1 U7410 ( .A1(n6850), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n6486), 
        .B2(n6848), .ZN(n6445) );
  OAI211_X1 U7411 ( .C1(n6545), .C2(n6853), .A(n6446), .B(n6445), .ZN(U3054)
         );
  AOI22_X1 U7412 ( .A1(n3024), .A2(n6549), .B1(n6489), .B2(n6844), .ZN(n6448)
         );
  AOI22_X1 U7413 ( .A1(n6850), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n6490), 
        .B2(n6848), .ZN(n6447) );
  OAI211_X1 U7414 ( .C1(n6552), .C2(n6853), .A(n6448), .B(n6447), .ZN(U3055)
         );
  AOI22_X1 U7415 ( .A1(n3024), .A2(n6556), .B1(n6493), .B2(n6844), .ZN(n6450)
         );
  AOI22_X1 U7416 ( .A1(n6850), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n6494), 
        .B2(n6848), .ZN(n6449) );
  OAI211_X1 U7417 ( .C1(n6554), .C2(n6853), .A(n6450), .B(n6449), .ZN(U3056)
         );
  AOI22_X1 U7418 ( .A1(n3024), .A2(n6563), .B1(n6497), .B2(n6844), .ZN(n6452)
         );
  AOI22_X1 U7419 ( .A1(n6850), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n6498), 
        .B2(n6848), .ZN(n6451) );
  OAI211_X1 U7420 ( .C1(n6566), .C2(n6853), .A(n6452), .B(n6451), .ZN(U3057)
         );
  AOI22_X1 U7421 ( .A1(n3024), .A2(n6578), .B1(n6504), .B2(n6844), .ZN(n6454)
         );
  AOI22_X1 U7422 ( .A1(n6850), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n6507), 
        .B2(n6848), .ZN(n6453) );
  OAI211_X1 U7423 ( .C1(n6574), .C2(n6853), .A(n6454), .B(n6453), .ZN(U3059)
         );
  AOI22_X1 U7424 ( .A1(n6456), .A2(n6530), .B1(n6470), .B2(n6455), .ZN(n6461)
         );
  AOI22_X1 U7425 ( .A1(n6459), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n6458), 
        .B2(n6457), .ZN(n6460) );
  OAI211_X1 U7426 ( .C1(n6513), .C2(n6462), .A(n6461), .B(n6460), .ZN(U3068)
         );
  INV_X1 U7427 ( .A(n6463), .ZN(n6468) );
  NAND2_X1 U7428 ( .A1(n6465), .A2(n6464), .ZN(n6466) );
  OAI22_X1 U7429 ( .A1(n6468), .A2(n6473), .B1(n6467), .B2(n6466), .ZN(n6505)
         );
  OR2_X1 U7430 ( .A1(n6469), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6475)
         );
  INV_X1 U7431 ( .A(n6475), .ZN(n6503) );
  AOI22_X1 U7432 ( .A1(n6505), .A2(n6530), .B1(n6470), .B2(n6503), .ZN(n6482)
         );
  OAI21_X1 U7433 ( .B1(n6506), .B2(n6471), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n6472) );
  OAI211_X1 U7434 ( .C1(n6474), .C2(n6473), .A(n6472), .B(n6515), .ZN(n6479)
         );
  NAND2_X1 U7435 ( .A1(n6475), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6476) );
  NAND4_X1 U7436 ( .A1(n6479), .A2(n6478), .A3(n6477), .A4(n6476), .ZN(n6508)
         );
  AOI22_X1 U7437 ( .A1(n6508), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n6480), 
        .B2(n6506), .ZN(n6481) );
  OAI211_X1 U7438 ( .C1(n6533), .C2(n6511), .A(n6482), .B(n6481), .ZN(U3084)
         );
  AOI22_X1 U7439 ( .A1(n6505), .A2(n6585), .B1(n6584), .B2(n6503), .ZN(n6484)
         );
  AOI22_X1 U7440 ( .A1(n6508), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n6586), 
        .B2(n6506), .ZN(n6483) );
  OAI211_X1 U7441 ( .C1(n6589), .C2(n6511), .A(n6484), .B(n6483), .ZN(U3085)
         );
  AOI22_X1 U7442 ( .A1(n6505), .A2(n6542), .B1(n6485), .B2(n6503), .ZN(n6488)
         );
  AOI22_X1 U7443 ( .A1(n6508), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n6486), 
        .B2(n6506), .ZN(n6487) );
  OAI211_X1 U7444 ( .C1(n6545), .C2(n6511), .A(n6488), .B(n6487), .ZN(U3086)
         );
  AOI22_X1 U7445 ( .A1(n6505), .A2(n6549), .B1(n6489), .B2(n6503), .ZN(n6492)
         );
  AOI22_X1 U7446 ( .A1(n6508), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n6490), 
        .B2(n6506), .ZN(n6491) );
  OAI211_X1 U7447 ( .C1(n6552), .C2(n6511), .A(n6492), .B(n6491), .ZN(U3087)
         );
  AOI22_X1 U7448 ( .A1(n6505), .A2(n6556), .B1(n6493), .B2(n6503), .ZN(n6496)
         );
  AOI22_X1 U7449 ( .A1(n6508), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n6494), 
        .B2(n6506), .ZN(n6495) );
  OAI211_X1 U7450 ( .C1(n6554), .C2(n6511), .A(n6496), .B(n6495), .ZN(U3088)
         );
  AOI22_X1 U7451 ( .A1(n6505), .A2(n6563), .B1(n6497), .B2(n6503), .ZN(n6500)
         );
  AOI22_X1 U7452 ( .A1(n6508), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n6498), 
        .B2(n6506), .ZN(n6499) );
  OAI211_X1 U7453 ( .C1(n6566), .C2(n6511), .A(n6500), .B(n6499), .ZN(U3089)
         );
  AOI22_X1 U7454 ( .A1(n6505), .A2(n6846), .B1(n6845), .B2(n6503), .ZN(n6502)
         );
  AOI22_X1 U7455 ( .A1(n6508), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n6849), 
        .B2(n6506), .ZN(n6501) );
  OAI211_X1 U7456 ( .C1(n6854), .C2(n6511), .A(n6502), .B(n6501), .ZN(U3090)
         );
  AOI22_X1 U7457 ( .A1(n6505), .A2(n6578), .B1(n6504), .B2(n6503), .ZN(n6510)
         );
  AOI22_X1 U7458 ( .A1(n6508), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n6507), 
        .B2(n6506), .ZN(n6509) );
  OAI211_X1 U7459 ( .C1(n6574), .C2(n6511), .A(n6510), .B(n6509), .ZN(U3091)
         );
  NAND2_X1 U7460 ( .A1(n6525), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6572) );
  OAI22_X1 U7461 ( .A1(n6596), .A2(n6513), .B1(n6512), .B2(n6572), .ZN(n6514)
         );
  INV_X1 U7462 ( .A(n6514), .ZN(n6532) );
  OAI21_X1 U7463 ( .B1(n6517), .B2(n6516), .A(n6515), .ZN(n6529) );
  INV_X1 U7464 ( .A(n6529), .ZN(n6521) );
  INV_X1 U7465 ( .A(n6572), .ZN(n6518) );
  AOI21_X1 U7466 ( .B1(n6520), .B2(n6519), .A(n6518), .ZN(n6528) );
  NAND2_X1 U7467 ( .A1(n6521), .A2(n6528), .ZN(n6523) );
  OAI211_X1 U7468 ( .C1(n6524), .C2(n6525), .A(n6523), .B(n6522), .ZN(n6579)
         );
  INV_X1 U7469 ( .A(n6525), .ZN(n6526) );
  OAI22_X1 U7470 ( .A1(n6529), .A2(n6528), .B1(n6527), .B2(n6526), .ZN(n6577)
         );
  AOI22_X1 U7471 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6579), .B1(n6530), 
        .B2(n6577), .ZN(n6531) );
  OAI211_X1 U7472 ( .C1(n6533), .C2(n6575), .A(n6532), .B(n6531), .ZN(U3108)
         );
  OAI22_X1 U7473 ( .A1(n6575), .A2(n6589), .B1(n6534), .B2(n6572), .ZN(n6535)
         );
  INV_X1 U7474 ( .A(n6535), .ZN(n6537) );
  AOI22_X1 U7475 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6579), .B1(n6585), 
        .B2(n6577), .ZN(n6536) );
  OAI211_X1 U7476 ( .C1(n6538), .C2(n6596), .A(n6537), .B(n6536), .ZN(U3109)
         );
  OAI22_X1 U7477 ( .A1(n6596), .A2(n6540), .B1(n6539), .B2(n6572), .ZN(n6541)
         );
  INV_X1 U7478 ( .A(n6541), .ZN(n6544) );
  AOI22_X1 U7479 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6579), .B1(n6542), 
        .B2(n6577), .ZN(n6543) );
  OAI211_X1 U7480 ( .C1(n6545), .C2(n6575), .A(n6544), .B(n6543), .ZN(U3110)
         );
  OAI22_X1 U7481 ( .A1(n6596), .A2(n6547), .B1(n6546), .B2(n6572), .ZN(n6548)
         );
  INV_X1 U7482 ( .A(n6548), .ZN(n6551) );
  AOI22_X1 U7483 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6579), .B1(n6549), 
        .B2(n6577), .ZN(n6550) );
  OAI211_X1 U7484 ( .C1(n6552), .C2(n6575), .A(n6551), .B(n6550), .ZN(U3111)
         );
  OAI22_X1 U7485 ( .A1(n6575), .A2(n6554), .B1(n6553), .B2(n6572), .ZN(n6555)
         );
  INV_X1 U7486 ( .A(n6555), .ZN(n6558) );
  AOI22_X1 U7487 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6579), .B1(n6556), 
        .B2(n6577), .ZN(n6557) );
  OAI211_X1 U7488 ( .C1(n6559), .C2(n6596), .A(n6558), .B(n6557), .ZN(U3112)
         );
  OAI22_X1 U7489 ( .A1(n6596), .A2(n6561), .B1(n6560), .B2(n6572), .ZN(n6562)
         );
  INV_X1 U7490 ( .A(n6562), .ZN(n6565) );
  AOI22_X1 U7491 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6579), .B1(n6563), 
        .B2(n6577), .ZN(n6564) );
  OAI211_X1 U7492 ( .C1(n6566), .C2(n6575), .A(n6565), .B(n6564), .ZN(U3113)
         );
  OAI22_X1 U7493 ( .A1(n6596), .A2(n6568), .B1(n6567), .B2(n6572), .ZN(n6569)
         );
  INV_X1 U7494 ( .A(n6569), .ZN(n6571) );
  AOI22_X1 U7495 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6579), .B1(n6846), 
        .B2(n6577), .ZN(n6570) );
  OAI211_X1 U7496 ( .C1(n6854), .C2(n6575), .A(n6571), .B(n6570), .ZN(U3114)
         );
  OAI22_X1 U7497 ( .A1(n6575), .A2(n6574), .B1(n6573), .B2(n6572), .ZN(n6576)
         );
  INV_X1 U7498 ( .A(n6576), .ZN(n6581) );
  AOI22_X1 U7499 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6579), .B1(n6578), 
        .B2(n6577), .ZN(n6580) );
  OAI211_X1 U7500 ( .C1(n6582), .C2(n6596), .A(n6581), .B(n6580), .ZN(U3115)
         );
  INV_X1 U7501 ( .A(n6583), .ZN(n6591) );
  AOI22_X1 U7502 ( .A1(n6591), .A2(n6585), .B1(n6584), .B2(n6590), .ZN(n6588)
         );
  AOI22_X1 U7503 ( .A1(n6593), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n6592), 
        .B2(n6586), .ZN(n6587) );
  OAI211_X1 U7504 ( .C1(n6589), .C2(n6596), .A(n6588), .B(n6587), .ZN(U3117)
         );
  AOI22_X1 U7505 ( .A1(n6591), .A2(n6846), .B1(n6845), .B2(n6590), .ZN(n6595)
         );
  AOI22_X1 U7506 ( .A1(n6593), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n6592), 
        .B2(n6849), .ZN(n6594) );
  OAI211_X1 U7507 ( .C1(n6854), .C2(n6596), .A(n6595), .B(n6594), .ZN(U3122)
         );
  AOI21_X1 U7508 ( .B1(n6598), .B2(n6597), .A(n6603), .ZN(n6601) );
  INV_X1 U7509 ( .A(n6599), .ZN(n6600) );
  NOR2_X1 U7510 ( .A1(n6601), .A2(n6600), .ZN(n6607) );
  OAI211_X1 U7511 ( .C1(n6605), .C2(n6604), .A(n6603), .B(n6602), .ZN(n6606)
         );
  OAI211_X1 U7512 ( .C1(n6609), .C2(n6608), .A(n6607), .B(n6606), .ZN(U3148)
         );
  AND2_X1 U7513 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6665), .ZN(U3151) );
  INV_X1 U7514 ( .A(DATAWIDTH_REG_30__SCAN_IN), .ZN(n6733) );
  NOR2_X1 U7515 ( .A1(n6669), .A2(n6733), .ZN(U3152) );
  AND2_X1 U7516 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6665), .ZN(U3153) );
  AND2_X1 U7517 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6665), .ZN(U3154) );
  AND2_X1 U7518 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6665), .ZN(U3155) );
  AND2_X1 U7519 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6665), .ZN(U3156) );
  AND2_X1 U7520 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6665), .ZN(U3157) );
  INV_X1 U7521 ( .A(DATAWIDTH_REG_24__SCAN_IN), .ZN(n6754) );
  NOR2_X1 U7522 ( .A1(n6669), .A2(n6754), .ZN(U3158) );
  AND2_X1 U7523 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n6665), .ZN(U3159) );
  AND2_X1 U7524 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6665), .ZN(U3160) );
  AND2_X1 U7525 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6665), .ZN(U3161) );
  AND2_X1 U7526 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6665), .ZN(U3162) );
  AND2_X1 U7527 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6665), .ZN(U3163) );
  AND2_X1 U7528 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6665), .ZN(U3164) );
  AND2_X1 U7529 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6665), .ZN(U3165) );
  AND2_X1 U7530 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6665), .ZN(U3166) );
  AND2_X1 U7531 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n6665), .ZN(U3167) );
  AND2_X1 U7532 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6665), .ZN(U3168) );
  AND2_X1 U7533 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6665), .ZN(U3169) );
  AND2_X1 U7534 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n6665), .ZN(U3170) );
  AND2_X1 U7535 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6665), .ZN(U3171) );
  INV_X1 U7536 ( .A(DATAWIDTH_REG_10__SCAN_IN), .ZN(n6761) );
  NOR2_X1 U7537 ( .A1(n6669), .A2(n6761), .ZN(U3172) );
  AND2_X1 U7538 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6665), .ZN(U3173) );
  AND2_X1 U7539 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n6665), .ZN(U3174) );
  INV_X1 U7540 ( .A(DATAWIDTH_REG_7__SCAN_IN), .ZN(n6728) );
  NOR2_X1 U7541 ( .A1(n6669), .A2(n6728), .ZN(U3175) );
  AND2_X1 U7542 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6665), .ZN(U3176) );
  AND2_X1 U7543 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n6665), .ZN(U3177) );
  AND2_X1 U7544 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6665), .ZN(U3178) );
  AND2_X1 U7545 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6665), .ZN(U3179) );
  AND2_X1 U7546 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6665), .ZN(U3180) );
  AOI22_X1 U7547 ( .A1(REIP_REG_1__SCAN_IN), .A2(n2966), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n6678), .ZN(n6611) );
  OAI21_X1 U7548 ( .B1(n6612), .B2(n6659), .A(n6611), .ZN(U3184) );
  AOI22_X1 U7549 ( .A1(REIP_REG_2__SCAN_IN), .A2(n2966), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6678), .ZN(n6613) );
  OAI21_X1 U7550 ( .B1(n6614), .B2(n6659), .A(n6613), .ZN(U3185) );
  AOI22_X1 U7551 ( .A1(REIP_REG_3__SCAN_IN), .A2(n2966), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6678), .ZN(n6615) );
  OAI21_X1 U7552 ( .B1(n6616), .B2(n6659), .A(n6615), .ZN(U3186) );
  AOI22_X1 U7553 ( .A1(REIP_REG_4__SCAN_IN), .A2(n2966), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6678), .ZN(n6617) );
  OAI21_X1 U7554 ( .B1(n6734), .B2(n6659), .A(n6617), .ZN(U3187) );
  AOI22_X1 U7555 ( .A1(REIP_REG_5__SCAN_IN), .A2(n2966), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6678), .ZN(n6618) );
  OAI21_X1 U7556 ( .B1(n4850), .B2(n6659), .A(n6618), .ZN(U3188) );
  AOI22_X1 U7557 ( .A1(REIP_REG_6__SCAN_IN), .A2(n2966), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6678), .ZN(n6619) );
  OAI21_X1 U7558 ( .B1(n6620), .B2(n6659), .A(n6619), .ZN(U3189) );
  AOI22_X1 U7559 ( .A1(REIP_REG_7__SCAN_IN), .A2(n2966), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n6678), .ZN(n6621) );
  OAI21_X1 U7560 ( .B1(n6623), .B2(n6659), .A(n6621), .ZN(U3190) );
  INV_X1 U7561 ( .A(n2966), .ZN(n6662) );
  INV_X1 U7562 ( .A(n6659), .ZN(n6660) );
  AOI22_X1 U7563 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6660), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n6678), .ZN(n6622) );
  OAI21_X1 U7564 ( .B1(n6623), .B2(n6662), .A(n6622), .ZN(U3191) );
  AOI22_X1 U7565 ( .A1(REIP_REG_9__SCAN_IN), .A2(n2966), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n6678), .ZN(n6624) );
  OAI21_X1 U7566 ( .B1(n6625), .B2(n6659), .A(n6624), .ZN(U3192) );
  AOI22_X1 U7567 ( .A1(REIP_REG_10__SCAN_IN), .A2(n2966), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n6678), .ZN(n6626) );
  OAI21_X1 U7568 ( .B1(n6627), .B2(n6659), .A(n6626), .ZN(U3193) );
  AOI22_X1 U7569 ( .A1(REIP_REG_11__SCAN_IN), .A2(n2966), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6678), .ZN(n6628) );
  OAI21_X1 U7570 ( .B1(n6629), .B2(n6659), .A(n6628), .ZN(U3194) );
  AOI22_X1 U7571 ( .A1(REIP_REG_12__SCAN_IN), .A2(n2966), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n6678), .ZN(n6630) );
  OAI21_X1 U7572 ( .B1(n6632), .B2(n6659), .A(n6630), .ZN(U3195) );
  AOI22_X1 U7573 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6660), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6678), .ZN(n6631) );
  OAI21_X1 U7574 ( .B1(n6632), .B2(n6662), .A(n6631), .ZN(U3196) );
  AOI22_X1 U7575 ( .A1(REIP_REG_14__SCAN_IN), .A2(n2966), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6678), .ZN(n6633) );
  OAI21_X1 U7576 ( .B1(n6751), .B2(n6659), .A(n6633), .ZN(U3197) );
  AOI22_X1 U7577 ( .A1(REIP_REG_16__SCAN_IN), .A2(n6660), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n6678), .ZN(n6634) );
  OAI21_X1 U7578 ( .B1(n6751), .B2(n6662), .A(n6634), .ZN(U3198) );
  INV_X1 U7579 ( .A(REIP_REG_17__SCAN_IN), .ZN(n6637) );
  AOI22_X1 U7580 ( .A1(REIP_REG_16__SCAN_IN), .A2(n2966), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6678), .ZN(n6635) );
  OAI21_X1 U7581 ( .B1(n6637), .B2(n6659), .A(n6635), .ZN(U3199) );
  AOI22_X1 U7582 ( .A1(REIP_REG_18__SCAN_IN), .A2(n6660), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6678), .ZN(n6636) );
  OAI21_X1 U7583 ( .B1(n6637), .B2(n6662), .A(n6636), .ZN(U3200) );
  INV_X1 U7584 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6639) );
  AOI22_X1 U7585 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6660), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n6678), .ZN(n6638) );
  OAI21_X1 U7586 ( .B1(n6639), .B2(n6662), .A(n6638), .ZN(U3201) );
  INV_X1 U7587 ( .A(REIP_REG_20__SCAN_IN), .ZN(n6641) );
  AOI22_X1 U7588 ( .A1(REIP_REG_19__SCAN_IN), .A2(n2966), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6678), .ZN(n6640) );
  OAI21_X1 U7589 ( .B1(n6641), .B2(n6659), .A(n6640), .ZN(U3202) );
  INV_X1 U7590 ( .A(ADDRESS_REG_19__SCAN_IN), .ZN(n6721) );
  OAI222_X1 U7591 ( .A1(n6662), .A2(n6641), .B1(n6721), .B2(n6688), .C1(n6643), 
        .C2(n6659), .ZN(U3203) );
  AOI22_X1 U7592 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6660), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n6678), .ZN(n6642) );
  OAI21_X1 U7593 ( .B1(n6643), .B2(n6662), .A(n6642), .ZN(U3204) );
  INV_X1 U7594 ( .A(ADDRESS_REG_21__SCAN_IN), .ZN(n6731) );
  OAI222_X1 U7595 ( .A1(n6662), .A2(n6645), .B1(n6731), .B2(n6688), .C1(n6644), 
        .C2(n6659), .ZN(U3205) );
  AOI22_X1 U7596 ( .A1(REIP_REG_23__SCAN_IN), .A2(n2966), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6678), .ZN(n6646) );
  OAI21_X1 U7597 ( .B1(n6647), .B2(n6659), .A(n6646), .ZN(U3206) );
  AOI22_X1 U7598 ( .A1(REIP_REG_24__SCAN_IN), .A2(n2966), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n6678), .ZN(n6648) );
  OAI21_X1 U7599 ( .B1(n6650), .B2(n6659), .A(n6648), .ZN(U3207) );
  AOI22_X1 U7600 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6660), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6678), .ZN(n6649) );
  OAI21_X1 U7601 ( .B1(n6650), .B2(n6662), .A(n6649), .ZN(U3208) );
  AOI22_X1 U7602 ( .A1(REIP_REG_26__SCAN_IN), .A2(n2966), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6678), .ZN(n6651) );
  OAI21_X1 U7603 ( .B1(n6652), .B2(n6659), .A(n6651), .ZN(U3209) );
  AOI22_X1 U7604 ( .A1(REIP_REG_27__SCAN_IN), .A2(n2966), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n6678), .ZN(n6653) );
  OAI21_X1 U7605 ( .B1(n6654), .B2(n6659), .A(n6653), .ZN(U3210) );
  AOI22_X1 U7606 ( .A1(REIP_REG_28__SCAN_IN), .A2(n2966), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n6678), .ZN(n6655) );
  OAI21_X1 U7607 ( .B1(n6656), .B2(n6659), .A(n6655), .ZN(U3211) );
  AOI22_X1 U7608 ( .A1(REIP_REG_29__SCAN_IN), .A2(n2966), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n6678), .ZN(n6658) );
  OAI21_X1 U7609 ( .B1(n6663), .B2(n6659), .A(n6658), .ZN(U3212) );
  AOI22_X1 U7610 ( .A1(REIP_REG_31__SCAN_IN), .A2(n6660), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6678), .ZN(n6661) );
  OAI21_X1 U7611 ( .B1(n6663), .B2(n6662), .A(n6661), .ZN(U3213) );
  MUX2_X1 U7612 ( .A(BE_N_REG_3__SCAN_IN), .B(BYTEENABLE_REG_3__SCAN_IN), .S(
        n6688), .Z(U3445) );
  MUX2_X1 U7613 ( .A(BE_N_REG_2__SCAN_IN), .B(BYTEENABLE_REG_2__SCAN_IN), .S(
        n6688), .Z(U3446) );
  MUX2_X1 U7614 ( .A(BE_N_REG_1__SCAN_IN), .B(BYTEENABLE_REG_1__SCAN_IN), .S(
        n6688), .Z(U3447) );
  MUX2_X1 U7615 ( .A(BE_N_REG_0__SCAN_IN), .B(BYTEENABLE_REG_0__SCAN_IN), .S(
        n6688), .Z(U3448) );
  INV_X1 U7616 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6666) );
  INV_X1 U7617 ( .A(n6667), .ZN(n6664) );
  AOI21_X1 U7618 ( .B1(n6666), .B2(n6665), .A(n6664), .ZN(U3451) );
  OAI21_X1 U7619 ( .B1(n6669), .B2(n6668), .A(n6667), .ZN(U3452) );
  AOI21_X1 U7620 ( .B1(REIP_REG_0__SCAN_IN), .B2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6670) );
  AOI22_X1 U7621 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .B1(
        n6670), .B2(n5522), .ZN(n6672) );
  INV_X1 U7622 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6671) );
  AOI22_X1 U7623 ( .A1(n6673), .A2(n6672), .B1(n6671), .B2(n6676), .ZN(U3468)
         );
  INV_X1 U7624 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6677) );
  NOR2_X1 U7625 ( .A1(n6676), .A2(REIP_REG_1__SCAN_IN), .ZN(n6674) );
  AOI22_X1 U7626 ( .A1(n6677), .A2(n6676), .B1(n6675), .B2(n6674), .ZN(U3469)
         );
  INV_X1 U7627 ( .A(W_R_N_REG_SCAN_IN), .ZN(n6822) );
  AOI22_X1 U7628 ( .A1(n6688), .A2(READREQUEST_REG_SCAN_IN), .B1(n6822), .B2(
        n6678), .ZN(U3470) );
  AOI211_X1 U7629 ( .C1(n6681), .C2(n6793), .A(n6680), .B(n6679), .ZN(n6687)
         );
  OAI211_X1 U7630 ( .C1(n4098), .C2(STATEBS16_REG_SCAN_IN), .A(n6682), .B(
        STATE2_REG_2__SCAN_IN), .ZN(n6684) );
  AOI21_X1 U7631 ( .B1(n6684), .B2(STATE2_REG_0__SCAN_IN), .A(n6683), .ZN(
        n6686) );
  NAND2_X1 U7632 ( .A1(n6687), .A2(REQUESTPENDING_REG_SCAN_IN), .ZN(n6685) );
  OAI21_X1 U7633 ( .B1(n6687), .B2(n6686), .A(n6685), .ZN(U3472) );
  MUX2_X1 U7634 ( .A(M_IO_N_REG_SCAN_IN), .B(MEMORYFETCH_REG_SCAN_IN), .S(
        n6688), .Z(U3473) );
  INV_X1 U7635 ( .A(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n6796) );
  NAND4_X1 U7636 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(
        INSTQUEUE_REG_9__4__SCAN_IN), .A3(INSTQUEUE_REG_7__7__SCAN_IN), .A4(
        n6796), .ZN(n6694) );
  INV_X1 U7637 ( .A(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n6730) );
  INV_X1 U7638 ( .A(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n6781) );
  NAND4_X1 U7639 ( .A1(INSTQUEUE_REG_14__2__SCAN_IN), .A2(
        INSTQUEUE_REG_0__2__SCAN_IN), .A3(n6730), .A4(n6781), .ZN(n6693) );
  NAND4_X1 U7640 ( .A1(INSTQUEUE_REG_2__3__SCAN_IN), .A2(STATE_REG_1__SCAN_IN), 
        .A3(INSTADDRPOINTER_REG_18__SCAN_IN), .A4(
        PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n6689) );
  INV_X1 U7641 ( .A(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n6798) );
  NOR3_X1 U7642 ( .A1(INSTQUEUE_REG_12__5__SCAN_IN), .A2(n6689), .A3(
        INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n6691) );
  INV_X1 U7643 ( .A(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n6690) );
  NAND3_X1 U7644 ( .A1(n6691), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .A3(n6690), 
        .ZN(n6692) );
  NOR3_X1 U7645 ( .A1(n6694), .A2(n6693), .A3(n6692), .ZN(n6843) );
  NAND4_X1 U7646 ( .A1(DATAI_13_), .A2(EAX_REG_6__SCAN_IN), .A3(
        ADDRESS_REG_19__SCAN_IN), .A4(n6718), .ZN(n6711) );
  NAND4_X1 U7647 ( .A1(DATAO_REG_5__SCAN_IN), .A2(DATAO_REG_25__SCAN_IN), .A3(
        n6753), .A4(n6744), .ZN(n6710) );
  NOR3_X1 U7648 ( .A1(REIP_REG_5__SCAN_IN), .A2(DATAI_3_), .A3(
        ADDRESS_REG_21__SCAN_IN), .ZN(n6696) );
  NOR3_X1 U7649 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(DATAO_REG_8__SCAN_IN), 
        .A3(n6736), .ZN(n6695) );
  NAND4_X1 U7650 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6696), .A3(
        DATAWIDTH_REG_24__SCAN_IN), .A4(n6695), .ZN(n6709) );
  INV_X1 U7651 ( .A(DATAI_23_), .ZN(n6697) );
  NAND4_X1 U7652 ( .A1(DATAO_REG_14__SCAN_IN), .A2(n6751), .A3(n6697), .A4(
        n6750), .ZN(n6701) );
  NAND4_X1 U7653 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        EAX_REG_12__SCAN_IN), .A3(DATAI_31_), .A4(DATAWIDTH_REG_10__SCAN_IN), 
        .ZN(n6700) );
  NAND4_X1 U7654 ( .A1(EAX_REG_19__SCAN_IN), .A2(EAX_REG_22__SCAN_IN), .A3(
        n6793), .A4(n3947), .ZN(n6699) );
  NAND4_X1 U7655 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(D_C_N_REG_SCAN_IN), 
        .A3(n6801), .A4(n5746), .ZN(n6698) );
  NOR4_X1 U7656 ( .A1(n6701), .A2(n6700), .A3(n6699), .A4(n6698), .ZN(n6707)
         );
  NOR3_X1 U7657 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        DATAO_REG_24__SCAN_IN), .A3(n6786), .ZN(n6706) );
  NAND4_X1 U7658 ( .A1(EAX_REG_27__SCAN_IN), .A2(UWORD_REG_2__SCAN_IN), .A3(
        W_R_N_REG_SCAN_IN), .A4(n6826), .ZN(n6704) );
  NAND3_X1 U7659 ( .A1(EAX_REG_26__SCAN_IN), .A2(REIP_REG_31__SCAN_IN), .A3(
        DATAI_28_), .ZN(n6703) );
  NAND4_X1 U7660 ( .A1(PHYADDRPOINTER_REG_22__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_10__SCAN_IN), .A3(n6808), .A4(n6811), .ZN(n6702) );
  NOR4_X1 U7661 ( .A1(NA_N), .A2(n6704), .A3(n6703), .A4(n6702), .ZN(n6705) );
  NAND4_X1 U7662 ( .A1(EBX_REG_15__SCAN_IN), .A2(n6707), .A3(n6706), .A4(n6705), .ZN(n6708) );
  NOR4_X1 U7663 ( .A1(n6711), .A2(n6710), .A3(n6709), .A4(n6708), .ZN(n6842)
         );
  AOI22_X1 U7664 ( .A1(n6714), .A2(keyinput44), .B1(keyinput58), .B2(n6713), 
        .ZN(n6712) );
  OAI221_X1 U7665 ( .B1(n6714), .B2(keyinput44), .C1(n6713), .C2(keyinput58), 
        .A(n6712), .ZN(n6725) );
  AOI22_X1 U7666 ( .A1(n6716), .A2(keyinput27), .B1(n3510), .B2(keyinput12), 
        .ZN(n6715) );
  OAI221_X1 U7667 ( .B1(n6716), .B2(keyinput27), .C1(n3510), .C2(keyinput12), 
        .A(n6715), .ZN(n6724) );
  AOI22_X1 U7668 ( .A1(n6718), .A2(keyinput38), .B1(n5031), .B2(keyinput63), 
        .ZN(n6717) );
  OAI221_X1 U7669 ( .B1(n6718), .B2(keyinput38), .C1(n5031), .C2(keyinput63), 
        .A(n6717), .ZN(n6723) );
  AOI22_X1 U7670 ( .A1(n6721), .A2(keyinput9), .B1(n6720), .B2(keyinput40), 
        .ZN(n6719) );
  OAI221_X1 U7671 ( .B1(n6721), .B2(keyinput9), .C1(n6720), .C2(keyinput40), 
        .A(n6719), .ZN(n6722) );
  NOR4_X1 U7672 ( .A1(n6725), .A2(n6724), .A3(n6723), .A4(n6722), .ZN(n6775)
         );
  INV_X1 U7673 ( .A(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n6727) );
  AOI22_X1 U7674 ( .A1(n6728), .A2(keyinput23), .B1(n6727), .B2(keyinput4), 
        .ZN(n6726) );
  OAI221_X1 U7675 ( .B1(n6728), .B2(keyinput23), .C1(n6727), .C2(keyinput4), 
        .A(n6726), .ZN(n6741) );
  AOI22_X1 U7676 ( .A1(n6731), .A2(keyinput61), .B1(n6730), .B2(keyinput22), 
        .ZN(n6729) );
  OAI221_X1 U7677 ( .B1(n6731), .B2(keyinput61), .C1(n6730), .C2(keyinput22), 
        .A(n6729), .ZN(n6740) );
  AOI22_X1 U7678 ( .A1(n6734), .A2(keyinput0), .B1(keyinput21), .B2(n6733), 
        .ZN(n6732) );
  OAI221_X1 U7679 ( .B1(n6734), .B2(keyinput0), .C1(n6733), .C2(keyinput21), 
        .A(n6732), .ZN(n6739) );
  AOI22_X1 U7680 ( .A1(n6737), .A2(keyinput60), .B1(n6736), .B2(keyinput6), 
        .ZN(n6735) );
  OAI221_X1 U7681 ( .B1(n6737), .B2(keyinput60), .C1(n6736), .C2(keyinput6), 
        .A(n6735), .ZN(n6738) );
  NOR4_X1 U7682 ( .A1(n6741), .A2(n6740), .A3(n6739), .A4(n6738), .ZN(n6774)
         );
  AOI22_X1 U7683 ( .A1(n6744), .A2(keyinput15), .B1(keyinput26), .B2(n6743), 
        .ZN(n6742) );
  OAI221_X1 U7684 ( .B1(n6744), .B2(keyinput15), .C1(n6743), .C2(keyinput26), 
        .A(n6742), .ZN(n6748) );
  XOR2_X1 U7685 ( .A(INSTQUEUE_REG_9__3__SCAN_IN), .B(keyinput35), .Z(n6747)
         );
  XNOR2_X1 U7686 ( .A(n6745), .B(keyinput1), .ZN(n6746) );
  OR3_X1 U7687 ( .A1(n6748), .A2(n6747), .A3(n6746), .ZN(n6757) );
  AOI22_X1 U7688 ( .A1(n6751), .A2(keyinput56), .B1(keyinput42), .B2(n6750), 
        .ZN(n6749) );
  OAI221_X1 U7689 ( .B1(n6751), .B2(keyinput56), .C1(n6750), .C2(keyinput42), 
        .A(n6749), .ZN(n6756) );
  AOI22_X1 U7690 ( .A1(n6754), .A2(keyinput55), .B1(n6753), .B2(keyinput59), 
        .ZN(n6752) );
  OAI221_X1 U7691 ( .B1(n6754), .B2(keyinput55), .C1(n6753), .C2(keyinput59), 
        .A(n6752), .ZN(n6755) );
  NOR3_X1 U7692 ( .A1(n6757), .A2(n6756), .A3(n6755), .ZN(n6773) );
  INV_X1 U7693 ( .A(DATAI_31_), .ZN(n6759) );
  AOI22_X1 U7694 ( .A1(n6759), .A2(keyinput37), .B1(n3947), .B2(keyinput28), 
        .ZN(n6758) );
  OAI221_X1 U7695 ( .B1(n6759), .B2(keyinput37), .C1(n3947), .C2(keyinput28), 
        .A(n6758), .ZN(n6771) );
  AOI22_X1 U7696 ( .A1(n6762), .A2(keyinput24), .B1(keyinput54), .B2(n6761), 
        .ZN(n6760) );
  OAI221_X1 U7697 ( .B1(n6762), .B2(keyinput24), .C1(n6761), .C2(keyinput54), 
        .A(n6760), .ZN(n6770) );
  AOI22_X1 U7698 ( .A1(n6765), .A2(keyinput16), .B1(n6764), .B2(keyinput62), 
        .ZN(n6763) );
  OAI221_X1 U7699 ( .B1(n6765), .B2(keyinput16), .C1(n6764), .C2(keyinput62), 
        .A(n6763), .ZN(n6769) );
  XNOR2_X1 U7700 ( .A(INSTQUEUE_REG_12__5__SCAN_IN), .B(keyinput11), .ZN(n6767) );
  XNOR2_X1 U7701 ( .A(keyinput57), .B(DATAI_23_), .ZN(n6766) );
  NAND2_X1 U7702 ( .A1(n6767), .A2(n6766), .ZN(n6768) );
  NOR4_X1 U7703 ( .A1(n6771), .A2(n6770), .A3(n6769), .A4(n6768), .ZN(n6772)
         );
  NAND4_X1 U7704 ( .A1(n6775), .A2(n6774), .A3(n6773), .A4(n6772), .ZN(n6841)
         );
  INV_X1 U7705 ( .A(D_C_N_REG_SCAN_IN), .ZN(n6778) );
  INV_X1 U7706 ( .A(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n6777) );
  AOI22_X1 U7707 ( .A1(n6778), .A2(keyinput29), .B1(n6777), .B2(keyinput53), 
        .ZN(n6776) );
  OAI221_X1 U7708 ( .B1(n6778), .B2(keyinput29), .C1(n6777), .C2(keyinput53), 
        .A(n6776), .ZN(n6790) );
  AOI22_X1 U7709 ( .A1(n6781), .A2(keyinput50), .B1(keyinput18), .B2(n6780), 
        .ZN(n6779) );
  OAI221_X1 U7710 ( .B1(n6781), .B2(keyinput50), .C1(n6780), .C2(keyinput18), 
        .A(n6779), .ZN(n6789) );
  AOI22_X1 U7711 ( .A1(n4656), .A2(keyinput17), .B1(n6783), .B2(keyinput30), 
        .ZN(n6782) );
  OAI221_X1 U7712 ( .B1(n4656), .B2(keyinput17), .C1(n6783), .C2(keyinput30), 
        .A(n6782), .ZN(n6788) );
  INV_X1 U7713 ( .A(EBX_REG_15__SCAN_IN), .ZN(n6785) );
  AOI22_X1 U7714 ( .A1(n6786), .A2(keyinput25), .B1(keyinput43), .B2(n6785), 
        .ZN(n6784) );
  OAI221_X1 U7715 ( .B1(n6786), .B2(keyinput25), .C1(n6785), .C2(keyinput43), 
        .A(n6784), .ZN(n6787) );
  NOR4_X1 U7716 ( .A1(n6790), .A2(n6789), .A3(n6788), .A4(n6787), .ZN(n6839)
         );
  AOI22_X1 U7717 ( .A1(n6793), .A2(keyinput31), .B1(keyinput36), .B2(n6792), 
        .ZN(n6791) );
  OAI221_X1 U7718 ( .B1(n6793), .B2(keyinput31), .C1(n6792), .C2(keyinput36), 
        .A(n6791), .ZN(n6805) );
  AOI22_X1 U7719 ( .A1(n6796), .A2(keyinput5), .B1(keyinput13), .B2(n6795), 
        .ZN(n6794) );
  OAI221_X1 U7720 ( .B1(n6796), .B2(keyinput5), .C1(n6795), .C2(keyinput13), 
        .A(n6794), .ZN(n6804) );
  AOI22_X1 U7721 ( .A1(n5746), .A2(keyinput7), .B1(n6798), .B2(keyinput47), 
        .ZN(n6797) );
  OAI221_X1 U7722 ( .B1(n5746), .B2(keyinput7), .C1(n6798), .C2(keyinput47), 
        .A(n6797), .ZN(n6803) );
  AOI22_X1 U7723 ( .A1(n6801), .A2(keyinput48), .B1(n6800), .B2(keyinput34), 
        .ZN(n6799) );
  OAI221_X1 U7724 ( .B1(n6801), .B2(keyinput48), .C1(n6800), .C2(keyinput34), 
        .A(n6799), .ZN(n6802) );
  NOR4_X1 U7725 ( .A1(n6805), .A2(n6804), .A3(n6803), .A4(n6802), .ZN(n6838)
         );
  AOI22_X1 U7726 ( .A1(n6808), .A2(keyinput46), .B1(keyinput19), .B2(n6807), 
        .ZN(n6806) );
  OAI221_X1 U7727 ( .B1(n6808), .B2(keyinput46), .C1(n6807), .C2(keyinput19), 
        .A(n6806), .ZN(n6820) );
  AOI22_X1 U7728 ( .A1(n6811), .A2(keyinput45), .B1(keyinput14), .B2(n6810), 
        .ZN(n6809) );
  OAI221_X1 U7729 ( .B1(n6811), .B2(keyinput45), .C1(n6810), .C2(keyinput14), 
        .A(n6809), .ZN(n6819) );
  AOI22_X1 U7730 ( .A1(n6814), .A2(keyinput8), .B1(keyinput3), .B2(n6813), 
        .ZN(n6812) );
  OAI221_X1 U7731 ( .B1(n6814), .B2(keyinput8), .C1(n6813), .C2(keyinput3), 
        .A(n6812), .ZN(n6818) );
  XNOR2_X1 U7732 ( .A(INSTQUEUE_REG_7__7__SCAN_IN), .B(keyinput33), .ZN(n6816)
         );
  XNOR2_X1 U7733 ( .A(keyinput32), .B(EAX_REG_26__SCAN_IN), .ZN(n6815) );
  NAND2_X1 U7734 ( .A1(n6816), .A2(n6815), .ZN(n6817) );
  NOR4_X1 U7735 ( .A1(n6820), .A2(n6819), .A3(n6818), .A4(n6817), .ZN(n6837)
         );
  AOI22_X1 U7736 ( .A1(n6823), .A2(keyinput49), .B1(keyinput51), .B2(n6822), 
        .ZN(n6821) );
  OAI221_X1 U7737 ( .B1(n6823), .B2(keyinput49), .C1(n6822), .C2(keyinput51), 
        .A(n6821), .ZN(n6835) );
  INV_X1 U7738 ( .A(EAX_REG_27__SCAN_IN), .ZN(n6825) );
  AOI22_X1 U7739 ( .A1(n6826), .A2(keyinput2), .B1(keyinput39), .B2(n6825), 
        .ZN(n6824) );
  OAI221_X1 U7740 ( .B1(n6826), .B2(keyinput2), .C1(n6825), .C2(keyinput39), 
        .A(n6824), .ZN(n6834) );
  INV_X1 U7741 ( .A(DATAI_28_), .ZN(n6828) );
  AOI22_X1 U7742 ( .A1(n6829), .A2(keyinput10), .B1(n6828), .B2(keyinput20), 
        .ZN(n6827) );
  OAI221_X1 U7743 ( .B1(n6829), .B2(keyinput10), .C1(n6828), .C2(keyinput20), 
        .A(n6827), .ZN(n6833) );
  XNOR2_X1 U7744 ( .A(INSTQUEUE_REG_9__4__SCAN_IN), .B(keyinput52), .ZN(n6831)
         );
  XNOR2_X1 U7745 ( .A(keyinput41), .B(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n6830)
         );
  NAND2_X1 U7746 ( .A1(n6831), .A2(n6830), .ZN(n6832) );
  NOR4_X1 U7747 ( .A1(n6835), .A2(n6834), .A3(n6833), .A4(n6832), .ZN(n6836)
         );
  NAND4_X1 U7748 ( .A1(n6839), .A2(n6838), .A3(n6837), .A4(n6836), .ZN(n6840)
         );
  AOI211_X1 U7749 ( .C1(n6843), .C2(n6842), .A(n6841), .B(n6840), .ZN(n6856)
         );
  AOI22_X1 U7750 ( .A1(n3024), .A2(n6846), .B1(n6845), .B2(n6844), .ZN(n6852)
         );
  AOI22_X1 U7751 ( .A1(n6850), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n6849), 
        .B2(n6848), .ZN(n6851) );
  OAI211_X1 U7752 ( .C1(n6854), .C2(n6853), .A(n6852), .B(n6851), .ZN(n6855)
         );
  XOR2_X1 U7753 ( .A(n6856), .B(n6855), .Z(U3058) );
  CLKBUF_X1 U3424 ( .A(n3917), .Z(n3881) );
  CLKBUF_X1 U3429 ( .A(n2970), .Z(n3806) );
  CLKBUF_X1 U3434 ( .A(n3363), .Z(n3441) );
  CLKBUF_X1 U34470 ( .A(n3349), .Z(n4483) );
  INV_X2 U3761 ( .A(n5760), .ZN(n5716) );
  CLKBUF_X1 U3822 ( .A(n5444), .Z(n2974) );
endmodule

